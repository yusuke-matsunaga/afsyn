module affine2(
  input clock,
  input reset,
  input start,
  output busy,
  output [1:0] imem00_bank,
  output imem00_rd,
  input [127:0] imem00_in,
  output [1:0] imem01_bank,
  output imem01_rd,
  input [127:0] imem01_in,
  output [1:0] imem02_bank,
  output imem02_rd,
  input [127:0] imem02_in,
  output [1:0] imem03_bank,
  output imem03_rd,
  input [127:0] imem03_in,
  output [1:0] imem04_bank,
  output imem04_rd,
  input [127:0] imem04_in,
  output [1:0] imem05_bank,
  output imem05_rd,
  input [127:0] imem05_in,
  output [1:0] imem06_bank,
  output imem06_rd,
  input [127:0] imem06_in,
  output [1:0] imem07_bank,
  output imem07_rd,
  input [127:0] imem07_in,
  output [5:0] omem00_bank,
  output omem00_wr,
  output [8:0] omem00_out,
  output [5:0] omem01_bank,
  output omem01_wr,
  output [8:0] omem01_out,
  output [5:0] omem02_bank,
  output omem02_wr,
  output [8:0] omem02_out,
  output [5:0] omem03_bank,
  output omem03_wr,
  output [8:0] omem03_out,
  output [5:0] omem04_bank,
  output omem04_wr,
  output [8:0] omem04_out);


  // 0 番目の OP1
  reg [3:0] op1_00_in00;
  reg       op1_00_inv00;
  reg [3:0] op1_00_in01;
  reg       op1_00_inv01;
  reg [3:0] op1_00_in02;
  reg       op1_00_inv02;
  reg [3:0] op1_00_in03;
  reg       op1_00_inv03;
  reg [3:0] op1_00_in04;
  reg       op1_00_inv04;
  reg [3:0] op1_00_in05;
  reg       op1_00_inv05;
  reg [3:0] op1_00_in06;
  reg       op1_00_inv06;
  reg [3:0] op1_00_in07;
  reg       op1_00_inv07;
  reg [3:0] op1_00_in08;
  reg       op1_00_inv08;
  reg [3:0] op1_00_in09;
  reg       op1_00_inv09;
  reg [3:0] op1_00_in10;
  reg       op1_00_inv10;
  reg [3:0] op1_00_in11;
  reg       op1_00_inv11;
  reg [3:0] op1_00_in12;
  reg       op1_00_inv12;
  reg [3:0] op1_00_in13;
  reg       op1_00_inv13;
  reg [3:0] op1_00_in14;
  reg       op1_00_inv14;
  reg [3:0] op1_00_in15;
  reg       op1_00_inv15;
  reg [3:0] op1_00_in16;
  reg       op1_00_inv16;
  reg [3:0] op1_00_in17;
  reg       op1_00_inv17;
  reg [3:0] op1_00_in18;
  reg       op1_00_inv18;
  reg [3:0] op1_00_in19;
  reg       op1_00_inv19;
  reg [3:0] op1_00_in20;
  reg       op1_00_inv20;
  reg [3:0] op1_00_in21;
  reg       op1_00_inv21;
  reg [3:0] op1_00_in22;
  reg       op1_00_inv22;
  reg [3:0] op1_00_in23;
  reg       op1_00_inv23;
  reg [3:0] op1_00_in24;
  reg       op1_00_inv24;
  reg [3:0] op1_00_in25;
  reg       op1_00_inv25;
  reg [3:0] op1_00_in26;
  reg       op1_00_inv26;
  reg [3:0] op1_00_in27;
  reg       op1_00_inv27;
  reg [3:0] op1_00_in28;
  reg       op1_00_inv28;
  reg [3:0] op1_00_in29;
  reg       op1_00_inv29;
  reg [3:0] op1_00_in30;
  reg       op1_00_inv30;
  reg [3:0] op1_00_in31;
  reg       op1_00_inv31;
  wire [8:0] op1_00_out;
  affine2_op1 op1_00(
    .data0_in(op1_00_in00),
    .inv0_in(op1_00_inv00),
    .data1_in(op1_00_in01),
    .inv1_in(op1_00_inv01),
    .data2_in(op1_00_in02),
    .inv2_in(op1_00_inv02),
    .data3_in(op1_00_in03),
    .inv3_in(op1_00_inv03),
    .data4_in(op1_00_in04),
    .inv4_in(op1_00_inv04),
    .data5_in(op1_00_in05),
    .inv5_in(op1_00_inv05),
    .data6_in(op1_00_in06),
    .inv6_in(op1_00_inv06),
    .data7_in(op1_00_in07),
    .inv7_in(op1_00_inv07),
    .data8_in(op1_00_in08),
    .inv8_in(op1_00_inv08),
    .data9_in(op1_00_in09),
    .inv9_in(op1_00_inv09),
    .data10_in(op1_00_in10),
    .inv10_in(op1_00_inv10),
    .data11_in(op1_00_in11),
    .inv11_in(op1_00_inv11),
    .data12_in(op1_00_in12),
    .inv12_in(op1_00_inv12),
    .data13_in(op1_00_in13),
    .inv13_in(op1_00_inv13),
    .data14_in(op1_00_in14),
    .inv14_in(op1_00_inv14),
    .data15_in(op1_00_in15),
    .inv15_in(op1_00_inv15),
    .data16_in(op1_00_in16),
    .inv16_in(op1_00_inv16),
    .data17_in(op1_00_in17),
    .inv17_in(op1_00_inv17),
    .data18_in(op1_00_in18),
    .inv18_in(op1_00_inv18),
    .data19_in(op1_00_in19),
    .inv19_in(op1_00_inv19),
    .data20_in(op1_00_in20),
    .inv20_in(op1_00_inv20),
    .data21_in(op1_00_in21),
    .inv21_in(op1_00_inv21),
    .data22_in(op1_00_in22),
    .inv22_in(op1_00_inv22),
    .data23_in(op1_00_in23),
    .inv23_in(op1_00_inv23),
    .data24_in(op1_00_in24),
    .inv24_in(op1_00_inv24),
    .data25_in(op1_00_in25),
    .inv25_in(op1_00_inv25),
    .data26_in(op1_00_in26),
    .inv26_in(op1_00_inv26),
    .data27_in(op1_00_in27),
    .inv27_in(op1_00_inv27),
    .data28_in(op1_00_in28),
    .inv28_in(op1_00_inv28),
    .data29_in(op1_00_in29),
    .inv29_in(op1_00_inv29),
    .data30_in(op1_00_in30),
    .inv30_in(op1_00_inv30),
    .data31_in(op1_00_in31),
    .inv31_in(op1_00_inv31),
    .data_out(op1_00_out));

  // 1 番目の OP1
  reg [3:0] op1_01_in00;
  reg       op1_01_inv00;
  reg [3:0] op1_01_in01;
  reg       op1_01_inv01;
  reg [3:0] op1_01_in02;
  reg       op1_01_inv02;
  reg [3:0] op1_01_in03;
  reg       op1_01_inv03;
  reg [3:0] op1_01_in04;
  reg       op1_01_inv04;
  reg [3:0] op1_01_in05;
  reg       op1_01_inv05;
  reg [3:0] op1_01_in06;
  reg       op1_01_inv06;
  reg [3:0] op1_01_in07;
  reg       op1_01_inv07;
  reg [3:0] op1_01_in08;
  reg       op1_01_inv08;
  reg [3:0] op1_01_in09;
  reg       op1_01_inv09;
  reg [3:0] op1_01_in10;
  reg       op1_01_inv10;
  reg [3:0] op1_01_in11;
  reg       op1_01_inv11;
  reg [3:0] op1_01_in12;
  reg       op1_01_inv12;
  reg [3:0] op1_01_in13;
  reg       op1_01_inv13;
  reg [3:0] op1_01_in14;
  reg       op1_01_inv14;
  reg [3:0] op1_01_in15;
  reg       op1_01_inv15;
  reg [3:0] op1_01_in16;
  reg       op1_01_inv16;
  reg [3:0] op1_01_in17;
  reg       op1_01_inv17;
  reg [3:0] op1_01_in18;
  reg       op1_01_inv18;
  reg [3:0] op1_01_in19;
  reg       op1_01_inv19;
  reg [3:0] op1_01_in20;
  reg       op1_01_inv20;
  reg [3:0] op1_01_in21;
  reg       op1_01_inv21;
  reg [3:0] op1_01_in22;
  reg       op1_01_inv22;
  reg [3:0] op1_01_in23;
  reg       op1_01_inv23;
  reg [3:0] op1_01_in24;
  reg       op1_01_inv24;
  reg [3:0] op1_01_in25;
  reg       op1_01_inv25;
  reg [3:0] op1_01_in26;
  reg       op1_01_inv26;
  reg [3:0] op1_01_in27;
  reg       op1_01_inv27;
  reg [3:0] op1_01_in28;
  reg       op1_01_inv28;
  reg [3:0] op1_01_in29;
  reg       op1_01_inv29;
  reg [3:0] op1_01_in30;
  reg       op1_01_inv30;
  reg [3:0] op1_01_in31;
  reg       op1_01_inv31;
  wire [8:0] op1_01_out;
  affine2_op1 op1_01(
    .data0_in(op1_01_in00),
    .inv0_in(op1_01_inv00),
    .data1_in(op1_01_in01),
    .inv1_in(op1_01_inv01),
    .data2_in(op1_01_in02),
    .inv2_in(op1_01_inv02),
    .data3_in(op1_01_in03),
    .inv3_in(op1_01_inv03),
    .data4_in(op1_01_in04),
    .inv4_in(op1_01_inv04),
    .data5_in(op1_01_in05),
    .inv5_in(op1_01_inv05),
    .data6_in(op1_01_in06),
    .inv6_in(op1_01_inv06),
    .data7_in(op1_01_in07),
    .inv7_in(op1_01_inv07),
    .data8_in(op1_01_in08),
    .inv8_in(op1_01_inv08),
    .data9_in(op1_01_in09),
    .inv9_in(op1_01_inv09),
    .data10_in(op1_01_in10),
    .inv10_in(op1_01_inv10),
    .data11_in(op1_01_in11),
    .inv11_in(op1_01_inv11),
    .data12_in(op1_01_in12),
    .inv12_in(op1_01_inv12),
    .data13_in(op1_01_in13),
    .inv13_in(op1_01_inv13),
    .data14_in(op1_01_in14),
    .inv14_in(op1_01_inv14),
    .data15_in(op1_01_in15),
    .inv15_in(op1_01_inv15),
    .data16_in(op1_01_in16),
    .inv16_in(op1_01_inv16),
    .data17_in(op1_01_in17),
    .inv17_in(op1_01_inv17),
    .data18_in(op1_01_in18),
    .inv18_in(op1_01_inv18),
    .data19_in(op1_01_in19),
    .inv19_in(op1_01_inv19),
    .data20_in(op1_01_in20),
    .inv20_in(op1_01_inv20),
    .data21_in(op1_01_in21),
    .inv21_in(op1_01_inv21),
    .data22_in(op1_01_in22),
    .inv22_in(op1_01_inv22),
    .data23_in(op1_01_in23),
    .inv23_in(op1_01_inv23),
    .data24_in(op1_01_in24),
    .inv24_in(op1_01_inv24),
    .data25_in(op1_01_in25),
    .inv25_in(op1_01_inv25),
    .data26_in(op1_01_in26),
    .inv26_in(op1_01_inv26),
    .data27_in(op1_01_in27),
    .inv27_in(op1_01_inv27),
    .data28_in(op1_01_in28),
    .inv28_in(op1_01_inv28),
    .data29_in(op1_01_in29),
    .inv29_in(op1_01_inv29),
    .data30_in(op1_01_in30),
    .inv30_in(op1_01_inv30),
    .data31_in(op1_01_in31),
    .inv31_in(op1_01_inv31),
    .data_out(op1_01_out));

  // 2 番目の OP1
  reg [3:0] op1_02_in00;
  reg       op1_02_inv00;
  reg [3:0] op1_02_in01;
  reg       op1_02_inv01;
  reg [3:0] op1_02_in02;
  reg       op1_02_inv02;
  reg [3:0] op1_02_in03;
  reg       op1_02_inv03;
  reg [3:0] op1_02_in04;
  reg       op1_02_inv04;
  reg [3:0] op1_02_in05;
  reg       op1_02_inv05;
  reg [3:0] op1_02_in06;
  reg       op1_02_inv06;
  reg [3:0] op1_02_in07;
  reg       op1_02_inv07;
  reg [3:0] op1_02_in08;
  reg       op1_02_inv08;
  reg [3:0] op1_02_in09;
  reg       op1_02_inv09;
  reg [3:0] op1_02_in10;
  reg       op1_02_inv10;
  reg [3:0] op1_02_in11;
  reg       op1_02_inv11;
  reg [3:0] op1_02_in12;
  reg       op1_02_inv12;
  reg [3:0] op1_02_in13;
  reg       op1_02_inv13;
  reg [3:0] op1_02_in14;
  reg       op1_02_inv14;
  reg [3:0] op1_02_in15;
  reg       op1_02_inv15;
  reg [3:0] op1_02_in16;
  reg       op1_02_inv16;
  reg [3:0] op1_02_in17;
  reg       op1_02_inv17;
  reg [3:0] op1_02_in18;
  reg       op1_02_inv18;
  reg [3:0] op1_02_in19;
  reg       op1_02_inv19;
  reg [3:0] op1_02_in20;
  reg       op1_02_inv20;
  reg [3:0] op1_02_in21;
  reg       op1_02_inv21;
  reg [3:0] op1_02_in22;
  reg       op1_02_inv22;
  reg [3:0] op1_02_in23;
  reg       op1_02_inv23;
  reg [3:0] op1_02_in24;
  reg       op1_02_inv24;
  reg [3:0] op1_02_in25;
  reg       op1_02_inv25;
  reg [3:0] op1_02_in26;
  reg       op1_02_inv26;
  reg [3:0] op1_02_in27;
  reg       op1_02_inv27;
  reg [3:0] op1_02_in28;
  reg       op1_02_inv28;
  reg [3:0] op1_02_in29;
  reg       op1_02_inv29;
  reg [3:0] op1_02_in30;
  reg       op1_02_inv30;
  reg [3:0] op1_02_in31;
  reg       op1_02_inv31;
  wire [8:0] op1_02_out;
  affine2_op1 op1_02(
    .data0_in(op1_02_in00),
    .inv0_in(op1_02_inv00),
    .data1_in(op1_02_in01),
    .inv1_in(op1_02_inv01),
    .data2_in(op1_02_in02),
    .inv2_in(op1_02_inv02),
    .data3_in(op1_02_in03),
    .inv3_in(op1_02_inv03),
    .data4_in(op1_02_in04),
    .inv4_in(op1_02_inv04),
    .data5_in(op1_02_in05),
    .inv5_in(op1_02_inv05),
    .data6_in(op1_02_in06),
    .inv6_in(op1_02_inv06),
    .data7_in(op1_02_in07),
    .inv7_in(op1_02_inv07),
    .data8_in(op1_02_in08),
    .inv8_in(op1_02_inv08),
    .data9_in(op1_02_in09),
    .inv9_in(op1_02_inv09),
    .data10_in(op1_02_in10),
    .inv10_in(op1_02_inv10),
    .data11_in(op1_02_in11),
    .inv11_in(op1_02_inv11),
    .data12_in(op1_02_in12),
    .inv12_in(op1_02_inv12),
    .data13_in(op1_02_in13),
    .inv13_in(op1_02_inv13),
    .data14_in(op1_02_in14),
    .inv14_in(op1_02_inv14),
    .data15_in(op1_02_in15),
    .inv15_in(op1_02_inv15),
    .data16_in(op1_02_in16),
    .inv16_in(op1_02_inv16),
    .data17_in(op1_02_in17),
    .inv17_in(op1_02_inv17),
    .data18_in(op1_02_in18),
    .inv18_in(op1_02_inv18),
    .data19_in(op1_02_in19),
    .inv19_in(op1_02_inv19),
    .data20_in(op1_02_in20),
    .inv20_in(op1_02_inv20),
    .data21_in(op1_02_in21),
    .inv21_in(op1_02_inv21),
    .data22_in(op1_02_in22),
    .inv22_in(op1_02_inv22),
    .data23_in(op1_02_in23),
    .inv23_in(op1_02_inv23),
    .data24_in(op1_02_in24),
    .inv24_in(op1_02_inv24),
    .data25_in(op1_02_in25),
    .inv25_in(op1_02_inv25),
    .data26_in(op1_02_in26),
    .inv26_in(op1_02_inv26),
    .data27_in(op1_02_in27),
    .inv27_in(op1_02_inv27),
    .data28_in(op1_02_in28),
    .inv28_in(op1_02_inv28),
    .data29_in(op1_02_in29),
    .inv29_in(op1_02_inv29),
    .data30_in(op1_02_in30),
    .inv30_in(op1_02_inv30),
    .data31_in(op1_02_in31),
    .inv31_in(op1_02_inv31),
    .data_out(op1_02_out));

  // 3 番目の OP1
  reg [3:0] op1_03_in00;
  reg       op1_03_inv00;
  reg [3:0] op1_03_in01;
  reg       op1_03_inv01;
  reg [3:0] op1_03_in02;
  reg       op1_03_inv02;
  reg [3:0] op1_03_in03;
  reg       op1_03_inv03;
  reg [3:0] op1_03_in04;
  reg       op1_03_inv04;
  reg [3:0] op1_03_in05;
  reg       op1_03_inv05;
  reg [3:0] op1_03_in06;
  reg       op1_03_inv06;
  reg [3:0] op1_03_in07;
  reg       op1_03_inv07;
  reg [3:0] op1_03_in08;
  reg       op1_03_inv08;
  reg [3:0] op1_03_in09;
  reg       op1_03_inv09;
  reg [3:0] op1_03_in10;
  reg       op1_03_inv10;
  reg [3:0] op1_03_in11;
  reg       op1_03_inv11;
  reg [3:0] op1_03_in12;
  reg       op1_03_inv12;
  reg [3:0] op1_03_in13;
  reg       op1_03_inv13;
  reg [3:0] op1_03_in14;
  reg       op1_03_inv14;
  reg [3:0] op1_03_in15;
  reg       op1_03_inv15;
  reg [3:0] op1_03_in16;
  reg       op1_03_inv16;
  reg [3:0] op1_03_in17;
  reg       op1_03_inv17;
  reg [3:0] op1_03_in18;
  reg       op1_03_inv18;
  reg [3:0] op1_03_in19;
  reg       op1_03_inv19;
  reg [3:0] op1_03_in20;
  reg       op1_03_inv20;
  reg [3:0] op1_03_in21;
  reg       op1_03_inv21;
  reg [3:0] op1_03_in22;
  reg       op1_03_inv22;
  reg [3:0] op1_03_in23;
  reg       op1_03_inv23;
  reg [3:0] op1_03_in24;
  reg       op1_03_inv24;
  reg [3:0] op1_03_in25;
  reg       op1_03_inv25;
  reg [3:0] op1_03_in26;
  reg       op1_03_inv26;
  reg [3:0] op1_03_in27;
  reg       op1_03_inv27;
  reg [3:0] op1_03_in28;
  reg       op1_03_inv28;
  reg [3:0] op1_03_in29;
  reg       op1_03_inv29;
  reg [3:0] op1_03_in30;
  reg       op1_03_inv30;
  reg [3:0] op1_03_in31;
  reg       op1_03_inv31;
  wire [8:0] op1_03_out;
  affine2_op1 op1_03(
    .data0_in(op1_03_in00),
    .inv0_in(op1_03_inv00),
    .data1_in(op1_03_in01),
    .inv1_in(op1_03_inv01),
    .data2_in(op1_03_in02),
    .inv2_in(op1_03_inv02),
    .data3_in(op1_03_in03),
    .inv3_in(op1_03_inv03),
    .data4_in(op1_03_in04),
    .inv4_in(op1_03_inv04),
    .data5_in(op1_03_in05),
    .inv5_in(op1_03_inv05),
    .data6_in(op1_03_in06),
    .inv6_in(op1_03_inv06),
    .data7_in(op1_03_in07),
    .inv7_in(op1_03_inv07),
    .data8_in(op1_03_in08),
    .inv8_in(op1_03_inv08),
    .data9_in(op1_03_in09),
    .inv9_in(op1_03_inv09),
    .data10_in(op1_03_in10),
    .inv10_in(op1_03_inv10),
    .data11_in(op1_03_in11),
    .inv11_in(op1_03_inv11),
    .data12_in(op1_03_in12),
    .inv12_in(op1_03_inv12),
    .data13_in(op1_03_in13),
    .inv13_in(op1_03_inv13),
    .data14_in(op1_03_in14),
    .inv14_in(op1_03_inv14),
    .data15_in(op1_03_in15),
    .inv15_in(op1_03_inv15),
    .data16_in(op1_03_in16),
    .inv16_in(op1_03_inv16),
    .data17_in(op1_03_in17),
    .inv17_in(op1_03_inv17),
    .data18_in(op1_03_in18),
    .inv18_in(op1_03_inv18),
    .data19_in(op1_03_in19),
    .inv19_in(op1_03_inv19),
    .data20_in(op1_03_in20),
    .inv20_in(op1_03_inv20),
    .data21_in(op1_03_in21),
    .inv21_in(op1_03_inv21),
    .data22_in(op1_03_in22),
    .inv22_in(op1_03_inv22),
    .data23_in(op1_03_in23),
    .inv23_in(op1_03_inv23),
    .data24_in(op1_03_in24),
    .inv24_in(op1_03_inv24),
    .data25_in(op1_03_in25),
    .inv25_in(op1_03_inv25),
    .data26_in(op1_03_in26),
    .inv26_in(op1_03_inv26),
    .data27_in(op1_03_in27),
    .inv27_in(op1_03_inv27),
    .data28_in(op1_03_in28),
    .inv28_in(op1_03_inv28),
    .data29_in(op1_03_in29),
    .inv29_in(op1_03_inv29),
    .data30_in(op1_03_in30),
    .inv30_in(op1_03_inv30),
    .data31_in(op1_03_in31),
    .inv31_in(op1_03_inv31),
    .data_out(op1_03_out));

  // 4 番目の OP1
  reg [3:0] op1_04_in00;
  reg       op1_04_inv00;
  reg [3:0] op1_04_in01;
  reg       op1_04_inv01;
  reg [3:0] op1_04_in02;
  reg       op1_04_inv02;
  reg [3:0] op1_04_in03;
  reg       op1_04_inv03;
  reg [3:0] op1_04_in04;
  reg       op1_04_inv04;
  reg [3:0] op1_04_in05;
  reg       op1_04_inv05;
  reg [3:0] op1_04_in06;
  reg       op1_04_inv06;
  reg [3:0] op1_04_in07;
  reg       op1_04_inv07;
  reg [3:0] op1_04_in08;
  reg       op1_04_inv08;
  reg [3:0] op1_04_in09;
  reg       op1_04_inv09;
  reg [3:0] op1_04_in10;
  reg       op1_04_inv10;
  reg [3:0] op1_04_in11;
  reg       op1_04_inv11;
  reg [3:0] op1_04_in12;
  reg       op1_04_inv12;
  reg [3:0] op1_04_in13;
  reg       op1_04_inv13;
  reg [3:0] op1_04_in14;
  reg       op1_04_inv14;
  reg [3:0] op1_04_in15;
  reg       op1_04_inv15;
  reg [3:0] op1_04_in16;
  reg       op1_04_inv16;
  reg [3:0] op1_04_in17;
  reg       op1_04_inv17;
  reg [3:0] op1_04_in18;
  reg       op1_04_inv18;
  reg [3:0] op1_04_in19;
  reg       op1_04_inv19;
  reg [3:0] op1_04_in20;
  reg       op1_04_inv20;
  reg [3:0] op1_04_in21;
  reg       op1_04_inv21;
  reg [3:0] op1_04_in22;
  reg       op1_04_inv22;
  reg [3:0] op1_04_in23;
  reg       op1_04_inv23;
  reg [3:0] op1_04_in24;
  reg       op1_04_inv24;
  reg [3:0] op1_04_in25;
  reg       op1_04_inv25;
  reg [3:0] op1_04_in26;
  reg       op1_04_inv26;
  reg [3:0] op1_04_in27;
  reg       op1_04_inv27;
  reg [3:0] op1_04_in28;
  reg       op1_04_inv28;
  reg [3:0] op1_04_in29;
  reg       op1_04_inv29;
  reg [3:0] op1_04_in30;
  reg       op1_04_inv30;
  reg [3:0] op1_04_in31;
  reg       op1_04_inv31;
  wire [8:0] op1_04_out;
  affine2_op1 op1_04(
    .data0_in(op1_04_in00),
    .inv0_in(op1_04_inv00),
    .data1_in(op1_04_in01),
    .inv1_in(op1_04_inv01),
    .data2_in(op1_04_in02),
    .inv2_in(op1_04_inv02),
    .data3_in(op1_04_in03),
    .inv3_in(op1_04_inv03),
    .data4_in(op1_04_in04),
    .inv4_in(op1_04_inv04),
    .data5_in(op1_04_in05),
    .inv5_in(op1_04_inv05),
    .data6_in(op1_04_in06),
    .inv6_in(op1_04_inv06),
    .data7_in(op1_04_in07),
    .inv7_in(op1_04_inv07),
    .data8_in(op1_04_in08),
    .inv8_in(op1_04_inv08),
    .data9_in(op1_04_in09),
    .inv9_in(op1_04_inv09),
    .data10_in(op1_04_in10),
    .inv10_in(op1_04_inv10),
    .data11_in(op1_04_in11),
    .inv11_in(op1_04_inv11),
    .data12_in(op1_04_in12),
    .inv12_in(op1_04_inv12),
    .data13_in(op1_04_in13),
    .inv13_in(op1_04_inv13),
    .data14_in(op1_04_in14),
    .inv14_in(op1_04_inv14),
    .data15_in(op1_04_in15),
    .inv15_in(op1_04_inv15),
    .data16_in(op1_04_in16),
    .inv16_in(op1_04_inv16),
    .data17_in(op1_04_in17),
    .inv17_in(op1_04_inv17),
    .data18_in(op1_04_in18),
    .inv18_in(op1_04_inv18),
    .data19_in(op1_04_in19),
    .inv19_in(op1_04_inv19),
    .data20_in(op1_04_in20),
    .inv20_in(op1_04_inv20),
    .data21_in(op1_04_in21),
    .inv21_in(op1_04_inv21),
    .data22_in(op1_04_in22),
    .inv22_in(op1_04_inv22),
    .data23_in(op1_04_in23),
    .inv23_in(op1_04_inv23),
    .data24_in(op1_04_in24),
    .inv24_in(op1_04_inv24),
    .data25_in(op1_04_in25),
    .inv25_in(op1_04_inv25),
    .data26_in(op1_04_in26),
    .inv26_in(op1_04_inv26),
    .data27_in(op1_04_in27),
    .inv27_in(op1_04_inv27),
    .data28_in(op1_04_in28),
    .inv28_in(op1_04_inv28),
    .data29_in(op1_04_in29),
    .inv29_in(op1_04_inv29),
    .data30_in(op1_04_in30),
    .inv30_in(op1_04_inv30),
    .data31_in(op1_04_in31),
    .inv31_in(op1_04_inv31),
    .data_out(op1_04_out));

  // 5 番目の OP1
  reg [3:0] op1_05_in00;
  reg       op1_05_inv00;
  reg [3:0] op1_05_in01;
  reg       op1_05_inv01;
  reg [3:0] op1_05_in02;
  reg       op1_05_inv02;
  reg [3:0] op1_05_in03;
  reg       op1_05_inv03;
  reg [3:0] op1_05_in04;
  reg       op1_05_inv04;
  reg [3:0] op1_05_in05;
  reg       op1_05_inv05;
  reg [3:0] op1_05_in06;
  reg       op1_05_inv06;
  reg [3:0] op1_05_in07;
  reg       op1_05_inv07;
  reg [3:0] op1_05_in08;
  reg       op1_05_inv08;
  reg [3:0] op1_05_in09;
  reg       op1_05_inv09;
  reg [3:0] op1_05_in10;
  reg       op1_05_inv10;
  reg [3:0] op1_05_in11;
  reg       op1_05_inv11;
  reg [3:0] op1_05_in12;
  reg       op1_05_inv12;
  reg [3:0] op1_05_in13;
  reg       op1_05_inv13;
  reg [3:0] op1_05_in14;
  reg       op1_05_inv14;
  reg [3:0] op1_05_in15;
  reg       op1_05_inv15;
  reg [3:0] op1_05_in16;
  reg       op1_05_inv16;
  reg [3:0] op1_05_in17;
  reg       op1_05_inv17;
  reg [3:0] op1_05_in18;
  reg       op1_05_inv18;
  reg [3:0] op1_05_in19;
  reg       op1_05_inv19;
  reg [3:0] op1_05_in20;
  reg       op1_05_inv20;
  reg [3:0] op1_05_in21;
  reg       op1_05_inv21;
  reg [3:0] op1_05_in22;
  reg       op1_05_inv22;
  reg [3:0] op1_05_in23;
  reg       op1_05_inv23;
  reg [3:0] op1_05_in24;
  reg       op1_05_inv24;
  reg [3:0] op1_05_in25;
  reg       op1_05_inv25;
  reg [3:0] op1_05_in26;
  reg       op1_05_inv26;
  reg [3:0] op1_05_in27;
  reg       op1_05_inv27;
  reg [3:0] op1_05_in28;
  reg       op1_05_inv28;
  reg [3:0] op1_05_in29;
  reg       op1_05_inv29;
  reg [3:0] op1_05_in30;
  reg       op1_05_inv30;
  reg [3:0] op1_05_in31;
  reg       op1_05_inv31;
  wire [8:0] op1_05_out;
  affine2_op1 op1_05(
    .data0_in(op1_05_in00),
    .inv0_in(op1_05_inv00),
    .data1_in(op1_05_in01),
    .inv1_in(op1_05_inv01),
    .data2_in(op1_05_in02),
    .inv2_in(op1_05_inv02),
    .data3_in(op1_05_in03),
    .inv3_in(op1_05_inv03),
    .data4_in(op1_05_in04),
    .inv4_in(op1_05_inv04),
    .data5_in(op1_05_in05),
    .inv5_in(op1_05_inv05),
    .data6_in(op1_05_in06),
    .inv6_in(op1_05_inv06),
    .data7_in(op1_05_in07),
    .inv7_in(op1_05_inv07),
    .data8_in(op1_05_in08),
    .inv8_in(op1_05_inv08),
    .data9_in(op1_05_in09),
    .inv9_in(op1_05_inv09),
    .data10_in(op1_05_in10),
    .inv10_in(op1_05_inv10),
    .data11_in(op1_05_in11),
    .inv11_in(op1_05_inv11),
    .data12_in(op1_05_in12),
    .inv12_in(op1_05_inv12),
    .data13_in(op1_05_in13),
    .inv13_in(op1_05_inv13),
    .data14_in(op1_05_in14),
    .inv14_in(op1_05_inv14),
    .data15_in(op1_05_in15),
    .inv15_in(op1_05_inv15),
    .data16_in(op1_05_in16),
    .inv16_in(op1_05_inv16),
    .data17_in(op1_05_in17),
    .inv17_in(op1_05_inv17),
    .data18_in(op1_05_in18),
    .inv18_in(op1_05_inv18),
    .data19_in(op1_05_in19),
    .inv19_in(op1_05_inv19),
    .data20_in(op1_05_in20),
    .inv20_in(op1_05_inv20),
    .data21_in(op1_05_in21),
    .inv21_in(op1_05_inv21),
    .data22_in(op1_05_in22),
    .inv22_in(op1_05_inv22),
    .data23_in(op1_05_in23),
    .inv23_in(op1_05_inv23),
    .data24_in(op1_05_in24),
    .inv24_in(op1_05_inv24),
    .data25_in(op1_05_in25),
    .inv25_in(op1_05_inv25),
    .data26_in(op1_05_in26),
    .inv26_in(op1_05_inv26),
    .data27_in(op1_05_in27),
    .inv27_in(op1_05_inv27),
    .data28_in(op1_05_in28),
    .inv28_in(op1_05_inv28),
    .data29_in(op1_05_in29),
    .inv29_in(op1_05_inv29),
    .data30_in(op1_05_in30),
    .inv30_in(op1_05_inv30),
    .data31_in(op1_05_in31),
    .inv31_in(op1_05_inv31),
    .data_out(op1_05_out));

  // 6 番目の OP1
  reg [3:0] op1_06_in00;
  reg       op1_06_inv00;
  reg [3:0] op1_06_in01;
  reg       op1_06_inv01;
  reg [3:0] op1_06_in02;
  reg       op1_06_inv02;
  reg [3:0] op1_06_in03;
  reg       op1_06_inv03;
  reg [3:0] op1_06_in04;
  reg       op1_06_inv04;
  reg [3:0] op1_06_in05;
  reg       op1_06_inv05;
  reg [3:0] op1_06_in06;
  reg       op1_06_inv06;
  reg [3:0] op1_06_in07;
  reg       op1_06_inv07;
  reg [3:0] op1_06_in08;
  reg       op1_06_inv08;
  reg [3:0] op1_06_in09;
  reg       op1_06_inv09;
  reg [3:0] op1_06_in10;
  reg       op1_06_inv10;
  reg [3:0] op1_06_in11;
  reg       op1_06_inv11;
  reg [3:0] op1_06_in12;
  reg       op1_06_inv12;
  reg [3:0] op1_06_in13;
  reg       op1_06_inv13;
  reg [3:0] op1_06_in14;
  reg       op1_06_inv14;
  reg [3:0] op1_06_in15;
  reg       op1_06_inv15;
  reg [3:0] op1_06_in16;
  reg       op1_06_inv16;
  reg [3:0] op1_06_in17;
  reg       op1_06_inv17;
  reg [3:0] op1_06_in18;
  reg       op1_06_inv18;
  reg [3:0] op1_06_in19;
  reg       op1_06_inv19;
  reg [3:0] op1_06_in20;
  reg       op1_06_inv20;
  reg [3:0] op1_06_in21;
  reg       op1_06_inv21;
  reg [3:0] op1_06_in22;
  reg       op1_06_inv22;
  reg [3:0] op1_06_in23;
  reg       op1_06_inv23;
  reg [3:0] op1_06_in24;
  reg       op1_06_inv24;
  reg [3:0] op1_06_in25;
  reg       op1_06_inv25;
  reg [3:0] op1_06_in26;
  reg       op1_06_inv26;
  reg [3:0] op1_06_in27;
  reg       op1_06_inv27;
  reg [3:0] op1_06_in28;
  reg       op1_06_inv28;
  reg [3:0] op1_06_in29;
  reg       op1_06_inv29;
  reg [3:0] op1_06_in30;
  reg       op1_06_inv30;
  reg [3:0] op1_06_in31;
  reg       op1_06_inv31;
  wire [8:0] op1_06_out;
  affine2_op1 op1_06(
    .data0_in(op1_06_in00),
    .inv0_in(op1_06_inv00),
    .data1_in(op1_06_in01),
    .inv1_in(op1_06_inv01),
    .data2_in(op1_06_in02),
    .inv2_in(op1_06_inv02),
    .data3_in(op1_06_in03),
    .inv3_in(op1_06_inv03),
    .data4_in(op1_06_in04),
    .inv4_in(op1_06_inv04),
    .data5_in(op1_06_in05),
    .inv5_in(op1_06_inv05),
    .data6_in(op1_06_in06),
    .inv6_in(op1_06_inv06),
    .data7_in(op1_06_in07),
    .inv7_in(op1_06_inv07),
    .data8_in(op1_06_in08),
    .inv8_in(op1_06_inv08),
    .data9_in(op1_06_in09),
    .inv9_in(op1_06_inv09),
    .data10_in(op1_06_in10),
    .inv10_in(op1_06_inv10),
    .data11_in(op1_06_in11),
    .inv11_in(op1_06_inv11),
    .data12_in(op1_06_in12),
    .inv12_in(op1_06_inv12),
    .data13_in(op1_06_in13),
    .inv13_in(op1_06_inv13),
    .data14_in(op1_06_in14),
    .inv14_in(op1_06_inv14),
    .data15_in(op1_06_in15),
    .inv15_in(op1_06_inv15),
    .data16_in(op1_06_in16),
    .inv16_in(op1_06_inv16),
    .data17_in(op1_06_in17),
    .inv17_in(op1_06_inv17),
    .data18_in(op1_06_in18),
    .inv18_in(op1_06_inv18),
    .data19_in(op1_06_in19),
    .inv19_in(op1_06_inv19),
    .data20_in(op1_06_in20),
    .inv20_in(op1_06_inv20),
    .data21_in(op1_06_in21),
    .inv21_in(op1_06_inv21),
    .data22_in(op1_06_in22),
    .inv22_in(op1_06_inv22),
    .data23_in(op1_06_in23),
    .inv23_in(op1_06_inv23),
    .data24_in(op1_06_in24),
    .inv24_in(op1_06_inv24),
    .data25_in(op1_06_in25),
    .inv25_in(op1_06_inv25),
    .data26_in(op1_06_in26),
    .inv26_in(op1_06_inv26),
    .data27_in(op1_06_in27),
    .inv27_in(op1_06_inv27),
    .data28_in(op1_06_in28),
    .inv28_in(op1_06_inv28),
    .data29_in(op1_06_in29),
    .inv29_in(op1_06_inv29),
    .data30_in(op1_06_in30),
    .inv30_in(op1_06_inv30),
    .data31_in(op1_06_in31),
    .inv31_in(op1_06_inv31),
    .data_out(op1_06_out));

  // 7 番目の OP1
  reg [3:0] op1_07_in00;
  reg       op1_07_inv00;
  reg [3:0] op1_07_in01;
  reg       op1_07_inv01;
  reg [3:0] op1_07_in02;
  reg       op1_07_inv02;
  reg [3:0] op1_07_in03;
  reg       op1_07_inv03;
  reg [3:0] op1_07_in04;
  reg       op1_07_inv04;
  reg [3:0] op1_07_in05;
  reg       op1_07_inv05;
  reg [3:0] op1_07_in06;
  reg       op1_07_inv06;
  reg [3:0] op1_07_in07;
  reg       op1_07_inv07;
  reg [3:0] op1_07_in08;
  reg       op1_07_inv08;
  reg [3:0] op1_07_in09;
  reg       op1_07_inv09;
  reg [3:0] op1_07_in10;
  reg       op1_07_inv10;
  reg [3:0] op1_07_in11;
  reg       op1_07_inv11;
  reg [3:0] op1_07_in12;
  reg       op1_07_inv12;
  reg [3:0] op1_07_in13;
  reg       op1_07_inv13;
  reg [3:0] op1_07_in14;
  reg       op1_07_inv14;
  reg [3:0] op1_07_in15;
  reg       op1_07_inv15;
  reg [3:0] op1_07_in16;
  reg       op1_07_inv16;
  reg [3:0] op1_07_in17;
  reg       op1_07_inv17;
  reg [3:0] op1_07_in18;
  reg       op1_07_inv18;
  reg [3:0] op1_07_in19;
  reg       op1_07_inv19;
  reg [3:0] op1_07_in20;
  reg       op1_07_inv20;
  reg [3:0] op1_07_in21;
  reg       op1_07_inv21;
  reg [3:0] op1_07_in22;
  reg       op1_07_inv22;
  reg [3:0] op1_07_in23;
  reg       op1_07_inv23;
  reg [3:0] op1_07_in24;
  reg       op1_07_inv24;
  reg [3:0] op1_07_in25;
  reg       op1_07_inv25;
  reg [3:0] op1_07_in26;
  reg       op1_07_inv26;
  reg [3:0] op1_07_in27;
  reg       op1_07_inv27;
  reg [3:0] op1_07_in28;
  reg       op1_07_inv28;
  reg [3:0] op1_07_in29;
  reg       op1_07_inv29;
  reg [3:0] op1_07_in30;
  reg       op1_07_inv30;
  reg [3:0] op1_07_in31;
  reg       op1_07_inv31;
  wire [8:0] op1_07_out;
  affine2_op1 op1_07(
    .data0_in(op1_07_in00),
    .inv0_in(op1_07_inv00),
    .data1_in(op1_07_in01),
    .inv1_in(op1_07_inv01),
    .data2_in(op1_07_in02),
    .inv2_in(op1_07_inv02),
    .data3_in(op1_07_in03),
    .inv3_in(op1_07_inv03),
    .data4_in(op1_07_in04),
    .inv4_in(op1_07_inv04),
    .data5_in(op1_07_in05),
    .inv5_in(op1_07_inv05),
    .data6_in(op1_07_in06),
    .inv6_in(op1_07_inv06),
    .data7_in(op1_07_in07),
    .inv7_in(op1_07_inv07),
    .data8_in(op1_07_in08),
    .inv8_in(op1_07_inv08),
    .data9_in(op1_07_in09),
    .inv9_in(op1_07_inv09),
    .data10_in(op1_07_in10),
    .inv10_in(op1_07_inv10),
    .data11_in(op1_07_in11),
    .inv11_in(op1_07_inv11),
    .data12_in(op1_07_in12),
    .inv12_in(op1_07_inv12),
    .data13_in(op1_07_in13),
    .inv13_in(op1_07_inv13),
    .data14_in(op1_07_in14),
    .inv14_in(op1_07_inv14),
    .data15_in(op1_07_in15),
    .inv15_in(op1_07_inv15),
    .data16_in(op1_07_in16),
    .inv16_in(op1_07_inv16),
    .data17_in(op1_07_in17),
    .inv17_in(op1_07_inv17),
    .data18_in(op1_07_in18),
    .inv18_in(op1_07_inv18),
    .data19_in(op1_07_in19),
    .inv19_in(op1_07_inv19),
    .data20_in(op1_07_in20),
    .inv20_in(op1_07_inv20),
    .data21_in(op1_07_in21),
    .inv21_in(op1_07_inv21),
    .data22_in(op1_07_in22),
    .inv22_in(op1_07_inv22),
    .data23_in(op1_07_in23),
    .inv23_in(op1_07_inv23),
    .data24_in(op1_07_in24),
    .inv24_in(op1_07_inv24),
    .data25_in(op1_07_in25),
    .inv25_in(op1_07_inv25),
    .data26_in(op1_07_in26),
    .inv26_in(op1_07_inv26),
    .data27_in(op1_07_in27),
    .inv27_in(op1_07_inv27),
    .data28_in(op1_07_in28),
    .inv28_in(op1_07_inv28),
    .data29_in(op1_07_in29),
    .inv29_in(op1_07_inv29),
    .data30_in(op1_07_in30),
    .inv30_in(op1_07_inv30),
    .data31_in(op1_07_in31),
    .inv31_in(op1_07_inv31),
    .data_out(op1_07_out));

  // 8 番目の OP1
  reg [3:0] op1_08_in00;
  reg       op1_08_inv00;
  reg [3:0] op1_08_in01;
  reg       op1_08_inv01;
  reg [3:0] op1_08_in02;
  reg       op1_08_inv02;
  reg [3:0] op1_08_in03;
  reg       op1_08_inv03;
  reg [3:0] op1_08_in04;
  reg       op1_08_inv04;
  reg [3:0] op1_08_in05;
  reg       op1_08_inv05;
  reg [3:0] op1_08_in06;
  reg       op1_08_inv06;
  reg [3:0] op1_08_in07;
  reg       op1_08_inv07;
  reg [3:0] op1_08_in08;
  reg       op1_08_inv08;
  reg [3:0] op1_08_in09;
  reg       op1_08_inv09;
  reg [3:0] op1_08_in10;
  reg       op1_08_inv10;
  reg [3:0] op1_08_in11;
  reg       op1_08_inv11;
  reg [3:0] op1_08_in12;
  reg       op1_08_inv12;
  reg [3:0] op1_08_in13;
  reg       op1_08_inv13;
  reg [3:0] op1_08_in14;
  reg       op1_08_inv14;
  reg [3:0] op1_08_in15;
  reg       op1_08_inv15;
  reg [3:0] op1_08_in16;
  reg       op1_08_inv16;
  reg [3:0] op1_08_in17;
  reg       op1_08_inv17;
  reg [3:0] op1_08_in18;
  reg       op1_08_inv18;
  reg [3:0] op1_08_in19;
  reg       op1_08_inv19;
  reg [3:0] op1_08_in20;
  reg       op1_08_inv20;
  reg [3:0] op1_08_in21;
  reg       op1_08_inv21;
  reg [3:0] op1_08_in22;
  reg       op1_08_inv22;
  reg [3:0] op1_08_in23;
  reg       op1_08_inv23;
  reg [3:0] op1_08_in24;
  reg       op1_08_inv24;
  reg [3:0] op1_08_in25;
  reg       op1_08_inv25;
  reg [3:0] op1_08_in26;
  reg       op1_08_inv26;
  reg [3:0] op1_08_in27;
  reg       op1_08_inv27;
  reg [3:0] op1_08_in28;
  reg       op1_08_inv28;
  reg [3:0] op1_08_in29;
  reg       op1_08_inv29;
  reg [3:0] op1_08_in30;
  reg       op1_08_inv30;
  reg [3:0] op1_08_in31;
  reg       op1_08_inv31;
  wire [8:0] op1_08_out;
  affine2_op1 op1_08(
    .data0_in(op1_08_in00),
    .inv0_in(op1_08_inv00),
    .data1_in(op1_08_in01),
    .inv1_in(op1_08_inv01),
    .data2_in(op1_08_in02),
    .inv2_in(op1_08_inv02),
    .data3_in(op1_08_in03),
    .inv3_in(op1_08_inv03),
    .data4_in(op1_08_in04),
    .inv4_in(op1_08_inv04),
    .data5_in(op1_08_in05),
    .inv5_in(op1_08_inv05),
    .data6_in(op1_08_in06),
    .inv6_in(op1_08_inv06),
    .data7_in(op1_08_in07),
    .inv7_in(op1_08_inv07),
    .data8_in(op1_08_in08),
    .inv8_in(op1_08_inv08),
    .data9_in(op1_08_in09),
    .inv9_in(op1_08_inv09),
    .data10_in(op1_08_in10),
    .inv10_in(op1_08_inv10),
    .data11_in(op1_08_in11),
    .inv11_in(op1_08_inv11),
    .data12_in(op1_08_in12),
    .inv12_in(op1_08_inv12),
    .data13_in(op1_08_in13),
    .inv13_in(op1_08_inv13),
    .data14_in(op1_08_in14),
    .inv14_in(op1_08_inv14),
    .data15_in(op1_08_in15),
    .inv15_in(op1_08_inv15),
    .data16_in(op1_08_in16),
    .inv16_in(op1_08_inv16),
    .data17_in(op1_08_in17),
    .inv17_in(op1_08_inv17),
    .data18_in(op1_08_in18),
    .inv18_in(op1_08_inv18),
    .data19_in(op1_08_in19),
    .inv19_in(op1_08_inv19),
    .data20_in(op1_08_in20),
    .inv20_in(op1_08_inv20),
    .data21_in(op1_08_in21),
    .inv21_in(op1_08_inv21),
    .data22_in(op1_08_in22),
    .inv22_in(op1_08_inv22),
    .data23_in(op1_08_in23),
    .inv23_in(op1_08_inv23),
    .data24_in(op1_08_in24),
    .inv24_in(op1_08_inv24),
    .data25_in(op1_08_in25),
    .inv25_in(op1_08_inv25),
    .data26_in(op1_08_in26),
    .inv26_in(op1_08_inv26),
    .data27_in(op1_08_in27),
    .inv27_in(op1_08_inv27),
    .data28_in(op1_08_in28),
    .inv28_in(op1_08_inv28),
    .data29_in(op1_08_in29),
    .inv29_in(op1_08_inv29),
    .data30_in(op1_08_in30),
    .inv30_in(op1_08_inv30),
    .data31_in(op1_08_in31),
    .inv31_in(op1_08_inv31),
    .data_out(op1_08_out));

  // 9 番目の OP1
  reg [3:0] op1_09_in00;
  reg       op1_09_inv00;
  reg [3:0] op1_09_in01;
  reg       op1_09_inv01;
  reg [3:0] op1_09_in02;
  reg       op1_09_inv02;
  reg [3:0] op1_09_in03;
  reg       op1_09_inv03;
  reg [3:0] op1_09_in04;
  reg       op1_09_inv04;
  reg [3:0] op1_09_in05;
  reg       op1_09_inv05;
  reg [3:0] op1_09_in06;
  reg       op1_09_inv06;
  reg [3:0] op1_09_in07;
  reg       op1_09_inv07;
  reg [3:0] op1_09_in08;
  reg       op1_09_inv08;
  reg [3:0] op1_09_in09;
  reg       op1_09_inv09;
  reg [3:0] op1_09_in10;
  reg       op1_09_inv10;
  reg [3:0] op1_09_in11;
  reg       op1_09_inv11;
  reg [3:0] op1_09_in12;
  reg       op1_09_inv12;
  reg [3:0] op1_09_in13;
  reg       op1_09_inv13;
  reg [3:0] op1_09_in14;
  reg       op1_09_inv14;
  reg [3:0] op1_09_in15;
  reg       op1_09_inv15;
  reg [3:0] op1_09_in16;
  reg       op1_09_inv16;
  reg [3:0] op1_09_in17;
  reg       op1_09_inv17;
  reg [3:0] op1_09_in18;
  reg       op1_09_inv18;
  reg [3:0] op1_09_in19;
  reg       op1_09_inv19;
  reg [3:0] op1_09_in20;
  reg       op1_09_inv20;
  reg [3:0] op1_09_in21;
  reg       op1_09_inv21;
  reg [3:0] op1_09_in22;
  reg       op1_09_inv22;
  reg [3:0] op1_09_in23;
  reg       op1_09_inv23;
  reg [3:0] op1_09_in24;
  reg       op1_09_inv24;
  reg [3:0] op1_09_in25;
  reg       op1_09_inv25;
  reg [3:0] op1_09_in26;
  reg       op1_09_inv26;
  reg [3:0] op1_09_in27;
  reg       op1_09_inv27;
  reg [3:0] op1_09_in28;
  reg       op1_09_inv28;
  reg [3:0] op1_09_in29;
  reg       op1_09_inv29;
  reg [3:0] op1_09_in30;
  reg       op1_09_inv30;
  reg [3:0] op1_09_in31;
  reg       op1_09_inv31;
  wire [8:0] op1_09_out;
  affine2_op1 op1_09(
    .data0_in(op1_09_in00),
    .inv0_in(op1_09_inv00),
    .data1_in(op1_09_in01),
    .inv1_in(op1_09_inv01),
    .data2_in(op1_09_in02),
    .inv2_in(op1_09_inv02),
    .data3_in(op1_09_in03),
    .inv3_in(op1_09_inv03),
    .data4_in(op1_09_in04),
    .inv4_in(op1_09_inv04),
    .data5_in(op1_09_in05),
    .inv5_in(op1_09_inv05),
    .data6_in(op1_09_in06),
    .inv6_in(op1_09_inv06),
    .data7_in(op1_09_in07),
    .inv7_in(op1_09_inv07),
    .data8_in(op1_09_in08),
    .inv8_in(op1_09_inv08),
    .data9_in(op1_09_in09),
    .inv9_in(op1_09_inv09),
    .data10_in(op1_09_in10),
    .inv10_in(op1_09_inv10),
    .data11_in(op1_09_in11),
    .inv11_in(op1_09_inv11),
    .data12_in(op1_09_in12),
    .inv12_in(op1_09_inv12),
    .data13_in(op1_09_in13),
    .inv13_in(op1_09_inv13),
    .data14_in(op1_09_in14),
    .inv14_in(op1_09_inv14),
    .data15_in(op1_09_in15),
    .inv15_in(op1_09_inv15),
    .data16_in(op1_09_in16),
    .inv16_in(op1_09_inv16),
    .data17_in(op1_09_in17),
    .inv17_in(op1_09_inv17),
    .data18_in(op1_09_in18),
    .inv18_in(op1_09_inv18),
    .data19_in(op1_09_in19),
    .inv19_in(op1_09_inv19),
    .data20_in(op1_09_in20),
    .inv20_in(op1_09_inv20),
    .data21_in(op1_09_in21),
    .inv21_in(op1_09_inv21),
    .data22_in(op1_09_in22),
    .inv22_in(op1_09_inv22),
    .data23_in(op1_09_in23),
    .inv23_in(op1_09_inv23),
    .data24_in(op1_09_in24),
    .inv24_in(op1_09_inv24),
    .data25_in(op1_09_in25),
    .inv25_in(op1_09_inv25),
    .data26_in(op1_09_in26),
    .inv26_in(op1_09_inv26),
    .data27_in(op1_09_in27),
    .inv27_in(op1_09_inv27),
    .data28_in(op1_09_in28),
    .inv28_in(op1_09_inv28),
    .data29_in(op1_09_in29),
    .inv29_in(op1_09_inv29),
    .data30_in(op1_09_in30),
    .inv30_in(op1_09_inv30),
    .data31_in(op1_09_in31),
    .inv31_in(op1_09_inv31),
    .data_out(op1_09_out));

  // 10 番目の OP1
  reg [3:0] op1_10_in00;
  reg       op1_10_inv00;
  reg [3:0] op1_10_in01;
  reg       op1_10_inv01;
  reg [3:0] op1_10_in02;
  reg       op1_10_inv02;
  reg [3:0] op1_10_in03;
  reg       op1_10_inv03;
  reg [3:0] op1_10_in04;
  reg       op1_10_inv04;
  reg [3:0] op1_10_in05;
  reg       op1_10_inv05;
  reg [3:0] op1_10_in06;
  reg       op1_10_inv06;
  reg [3:0] op1_10_in07;
  reg       op1_10_inv07;
  reg [3:0] op1_10_in08;
  reg       op1_10_inv08;
  reg [3:0] op1_10_in09;
  reg       op1_10_inv09;
  reg [3:0] op1_10_in10;
  reg       op1_10_inv10;
  reg [3:0] op1_10_in11;
  reg       op1_10_inv11;
  reg [3:0] op1_10_in12;
  reg       op1_10_inv12;
  reg [3:0] op1_10_in13;
  reg       op1_10_inv13;
  reg [3:0] op1_10_in14;
  reg       op1_10_inv14;
  reg [3:0] op1_10_in15;
  reg       op1_10_inv15;
  reg [3:0] op1_10_in16;
  reg       op1_10_inv16;
  reg [3:0] op1_10_in17;
  reg       op1_10_inv17;
  reg [3:0] op1_10_in18;
  reg       op1_10_inv18;
  reg [3:0] op1_10_in19;
  reg       op1_10_inv19;
  reg [3:0] op1_10_in20;
  reg       op1_10_inv20;
  reg [3:0] op1_10_in21;
  reg       op1_10_inv21;
  reg [3:0] op1_10_in22;
  reg       op1_10_inv22;
  reg [3:0] op1_10_in23;
  reg       op1_10_inv23;
  reg [3:0] op1_10_in24;
  reg       op1_10_inv24;
  reg [3:0] op1_10_in25;
  reg       op1_10_inv25;
  reg [3:0] op1_10_in26;
  reg       op1_10_inv26;
  reg [3:0] op1_10_in27;
  reg       op1_10_inv27;
  reg [3:0] op1_10_in28;
  reg       op1_10_inv28;
  reg [3:0] op1_10_in29;
  reg       op1_10_inv29;
  reg [3:0] op1_10_in30;
  reg       op1_10_inv30;
  reg [3:0] op1_10_in31;
  reg       op1_10_inv31;
  wire [8:0] op1_10_out;
  affine2_op1 op1_10(
    .data0_in(op1_10_in00),
    .inv0_in(op1_10_inv00),
    .data1_in(op1_10_in01),
    .inv1_in(op1_10_inv01),
    .data2_in(op1_10_in02),
    .inv2_in(op1_10_inv02),
    .data3_in(op1_10_in03),
    .inv3_in(op1_10_inv03),
    .data4_in(op1_10_in04),
    .inv4_in(op1_10_inv04),
    .data5_in(op1_10_in05),
    .inv5_in(op1_10_inv05),
    .data6_in(op1_10_in06),
    .inv6_in(op1_10_inv06),
    .data7_in(op1_10_in07),
    .inv7_in(op1_10_inv07),
    .data8_in(op1_10_in08),
    .inv8_in(op1_10_inv08),
    .data9_in(op1_10_in09),
    .inv9_in(op1_10_inv09),
    .data10_in(op1_10_in10),
    .inv10_in(op1_10_inv10),
    .data11_in(op1_10_in11),
    .inv11_in(op1_10_inv11),
    .data12_in(op1_10_in12),
    .inv12_in(op1_10_inv12),
    .data13_in(op1_10_in13),
    .inv13_in(op1_10_inv13),
    .data14_in(op1_10_in14),
    .inv14_in(op1_10_inv14),
    .data15_in(op1_10_in15),
    .inv15_in(op1_10_inv15),
    .data16_in(op1_10_in16),
    .inv16_in(op1_10_inv16),
    .data17_in(op1_10_in17),
    .inv17_in(op1_10_inv17),
    .data18_in(op1_10_in18),
    .inv18_in(op1_10_inv18),
    .data19_in(op1_10_in19),
    .inv19_in(op1_10_inv19),
    .data20_in(op1_10_in20),
    .inv20_in(op1_10_inv20),
    .data21_in(op1_10_in21),
    .inv21_in(op1_10_inv21),
    .data22_in(op1_10_in22),
    .inv22_in(op1_10_inv22),
    .data23_in(op1_10_in23),
    .inv23_in(op1_10_inv23),
    .data24_in(op1_10_in24),
    .inv24_in(op1_10_inv24),
    .data25_in(op1_10_in25),
    .inv25_in(op1_10_inv25),
    .data26_in(op1_10_in26),
    .inv26_in(op1_10_inv26),
    .data27_in(op1_10_in27),
    .inv27_in(op1_10_inv27),
    .data28_in(op1_10_in28),
    .inv28_in(op1_10_inv28),
    .data29_in(op1_10_in29),
    .inv29_in(op1_10_inv29),
    .data30_in(op1_10_in30),
    .inv30_in(op1_10_inv30),
    .data31_in(op1_10_in31),
    .inv31_in(op1_10_inv31),
    .data_out(op1_10_out));

  // 11 番目の OP1
  reg [3:0] op1_11_in00;
  reg       op1_11_inv00;
  reg [3:0] op1_11_in01;
  reg       op1_11_inv01;
  reg [3:0] op1_11_in02;
  reg       op1_11_inv02;
  reg [3:0] op1_11_in03;
  reg       op1_11_inv03;
  reg [3:0] op1_11_in04;
  reg       op1_11_inv04;
  reg [3:0] op1_11_in05;
  reg       op1_11_inv05;
  reg [3:0] op1_11_in06;
  reg       op1_11_inv06;
  reg [3:0] op1_11_in07;
  reg       op1_11_inv07;
  reg [3:0] op1_11_in08;
  reg       op1_11_inv08;
  reg [3:0] op1_11_in09;
  reg       op1_11_inv09;
  reg [3:0] op1_11_in10;
  reg       op1_11_inv10;
  reg [3:0] op1_11_in11;
  reg       op1_11_inv11;
  reg [3:0] op1_11_in12;
  reg       op1_11_inv12;
  reg [3:0] op1_11_in13;
  reg       op1_11_inv13;
  reg [3:0] op1_11_in14;
  reg       op1_11_inv14;
  reg [3:0] op1_11_in15;
  reg       op1_11_inv15;
  reg [3:0] op1_11_in16;
  reg       op1_11_inv16;
  reg [3:0] op1_11_in17;
  reg       op1_11_inv17;
  reg [3:0] op1_11_in18;
  reg       op1_11_inv18;
  reg [3:0] op1_11_in19;
  reg       op1_11_inv19;
  reg [3:0] op1_11_in20;
  reg       op1_11_inv20;
  reg [3:0] op1_11_in21;
  reg       op1_11_inv21;
  reg [3:0] op1_11_in22;
  reg       op1_11_inv22;
  reg [3:0] op1_11_in23;
  reg       op1_11_inv23;
  reg [3:0] op1_11_in24;
  reg       op1_11_inv24;
  reg [3:0] op1_11_in25;
  reg       op1_11_inv25;
  reg [3:0] op1_11_in26;
  reg       op1_11_inv26;
  reg [3:0] op1_11_in27;
  reg       op1_11_inv27;
  reg [3:0] op1_11_in28;
  reg       op1_11_inv28;
  reg [3:0] op1_11_in29;
  reg       op1_11_inv29;
  reg [3:0] op1_11_in30;
  reg       op1_11_inv30;
  reg [3:0] op1_11_in31;
  reg       op1_11_inv31;
  wire [8:0] op1_11_out;
  affine2_op1 op1_11(
    .data0_in(op1_11_in00),
    .inv0_in(op1_11_inv00),
    .data1_in(op1_11_in01),
    .inv1_in(op1_11_inv01),
    .data2_in(op1_11_in02),
    .inv2_in(op1_11_inv02),
    .data3_in(op1_11_in03),
    .inv3_in(op1_11_inv03),
    .data4_in(op1_11_in04),
    .inv4_in(op1_11_inv04),
    .data5_in(op1_11_in05),
    .inv5_in(op1_11_inv05),
    .data6_in(op1_11_in06),
    .inv6_in(op1_11_inv06),
    .data7_in(op1_11_in07),
    .inv7_in(op1_11_inv07),
    .data8_in(op1_11_in08),
    .inv8_in(op1_11_inv08),
    .data9_in(op1_11_in09),
    .inv9_in(op1_11_inv09),
    .data10_in(op1_11_in10),
    .inv10_in(op1_11_inv10),
    .data11_in(op1_11_in11),
    .inv11_in(op1_11_inv11),
    .data12_in(op1_11_in12),
    .inv12_in(op1_11_inv12),
    .data13_in(op1_11_in13),
    .inv13_in(op1_11_inv13),
    .data14_in(op1_11_in14),
    .inv14_in(op1_11_inv14),
    .data15_in(op1_11_in15),
    .inv15_in(op1_11_inv15),
    .data16_in(op1_11_in16),
    .inv16_in(op1_11_inv16),
    .data17_in(op1_11_in17),
    .inv17_in(op1_11_inv17),
    .data18_in(op1_11_in18),
    .inv18_in(op1_11_inv18),
    .data19_in(op1_11_in19),
    .inv19_in(op1_11_inv19),
    .data20_in(op1_11_in20),
    .inv20_in(op1_11_inv20),
    .data21_in(op1_11_in21),
    .inv21_in(op1_11_inv21),
    .data22_in(op1_11_in22),
    .inv22_in(op1_11_inv22),
    .data23_in(op1_11_in23),
    .inv23_in(op1_11_inv23),
    .data24_in(op1_11_in24),
    .inv24_in(op1_11_inv24),
    .data25_in(op1_11_in25),
    .inv25_in(op1_11_inv25),
    .data26_in(op1_11_in26),
    .inv26_in(op1_11_inv26),
    .data27_in(op1_11_in27),
    .inv27_in(op1_11_inv27),
    .data28_in(op1_11_in28),
    .inv28_in(op1_11_inv28),
    .data29_in(op1_11_in29),
    .inv29_in(op1_11_inv29),
    .data30_in(op1_11_in30),
    .inv30_in(op1_11_inv30),
    .data31_in(op1_11_in31),
    .inv31_in(op1_11_inv31),
    .data_out(op1_11_out));

  // 12 番目の OP1
  reg [3:0] op1_12_in00;
  reg       op1_12_inv00;
  reg [3:0] op1_12_in01;
  reg       op1_12_inv01;
  reg [3:0] op1_12_in02;
  reg       op1_12_inv02;
  reg [3:0] op1_12_in03;
  reg       op1_12_inv03;
  reg [3:0] op1_12_in04;
  reg       op1_12_inv04;
  reg [3:0] op1_12_in05;
  reg       op1_12_inv05;
  reg [3:0] op1_12_in06;
  reg       op1_12_inv06;
  reg [3:0] op1_12_in07;
  reg       op1_12_inv07;
  reg [3:0] op1_12_in08;
  reg       op1_12_inv08;
  reg [3:0] op1_12_in09;
  reg       op1_12_inv09;
  reg [3:0] op1_12_in10;
  reg       op1_12_inv10;
  reg [3:0] op1_12_in11;
  reg       op1_12_inv11;
  reg [3:0] op1_12_in12;
  reg       op1_12_inv12;
  reg [3:0] op1_12_in13;
  reg       op1_12_inv13;
  reg [3:0] op1_12_in14;
  reg       op1_12_inv14;
  reg [3:0] op1_12_in15;
  reg       op1_12_inv15;
  reg [3:0] op1_12_in16;
  reg       op1_12_inv16;
  reg [3:0] op1_12_in17;
  reg       op1_12_inv17;
  reg [3:0] op1_12_in18;
  reg       op1_12_inv18;
  reg [3:0] op1_12_in19;
  reg       op1_12_inv19;
  reg [3:0] op1_12_in20;
  reg       op1_12_inv20;
  reg [3:0] op1_12_in21;
  reg       op1_12_inv21;
  reg [3:0] op1_12_in22;
  reg       op1_12_inv22;
  reg [3:0] op1_12_in23;
  reg       op1_12_inv23;
  reg [3:0] op1_12_in24;
  reg       op1_12_inv24;
  reg [3:0] op1_12_in25;
  reg       op1_12_inv25;
  reg [3:0] op1_12_in26;
  reg       op1_12_inv26;
  reg [3:0] op1_12_in27;
  reg       op1_12_inv27;
  reg [3:0] op1_12_in28;
  reg       op1_12_inv28;
  reg [3:0] op1_12_in29;
  reg       op1_12_inv29;
  reg [3:0] op1_12_in30;
  reg       op1_12_inv30;
  reg [3:0] op1_12_in31;
  reg       op1_12_inv31;
  wire [8:0] op1_12_out;
  affine2_op1 op1_12(
    .data0_in(op1_12_in00),
    .inv0_in(op1_12_inv00),
    .data1_in(op1_12_in01),
    .inv1_in(op1_12_inv01),
    .data2_in(op1_12_in02),
    .inv2_in(op1_12_inv02),
    .data3_in(op1_12_in03),
    .inv3_in(op1_12_inv03),
    .data4_in(op1_12_in04),
    .inv4_in(op1_12_inv04),
    .data5_in(op1_12_in05),
    .inv5_in(op1_12_inv05),
    .data6_in(op1_12_in06),
    .inv6_in(op1_12_inv06),
    .data7_in(op1_12_in07),
    .inv7_in(op1_12_inv07),
    .data8_in(op1_12_in08),
    .inv8_in(op1_12_inv08),
    .data9_in(op1_12_in09),
    .inv9_in(op1_12_inv09),
    .data10_in(op1_12_in10),
    .inv10_in(op1_12_inv10),
    .data11_in(op1_12_in11),
    .inv11_in(op1_12_inv11),
    .data12_in(op1_12_in12),
    .inv12_in(op1_12_inv12),
    .data13_in(op1_12_in13),
    .inv13_in(op1_12_inv13),
    .data14_in(op1_12_in14),
    .inv14_in(op1_12_inv14),
    .data15_in(op1_12_in15),
    .inv15_in(op1_12_inv15),
    .data16_in(op1_12_in16),
    .inv16_in(op1_12_inv16),
    .data17_in(op1_12_in17),
    .inv17_in(op1_12_inv17),
    .data18_in(op1_12_in18),
    .inv18_in(op1_12_inv18),
    .data19_in(op1_12_in19),
    .inv19_in(op1_12_inv19),
    .data20_in(op1_12_in20),
    .inv20_in(op1_12_inv20),
    .data21_in(op1_12_in21),
    .inv21_in(op1_12_inv21),
    .data22_in(op1_12_in22),
    .inv22_in(op1_12_inv22),
    .data23_in(op1_12_in23),
    .inv23_in(op1_12_inv23),
    .data24_in(op1_12_in24),
    .inv24_in(op1_12_inv24),
    .data25_in(op1_12_in25),
    .inv25_in(op1_12_inv25),
    .data26_in(op1_12_in26),
    .inv26_in(op1_12_inv26),
    .data27_in(op1_12_in27),
    .inv27_in(op1_12_inv27),
    .data28_in(op1_12_in28),
    .inv28_in(op1_12_inv28),
    .data29_in(op1_12_in29),
    .inv29_in(op1_12_inv29),
    .data30_in(op1_12_in30),
    .inv30_in(op1_12_inv30),
    .data31_in(op1_12_in31),
    .inv31_in(op1_12_inv31),
    .data_out(op1_12_out));

  // 13 番目の OP1
  reg [3:0] op1_13_in00;
  reg       op1_13_inv00;
  reg [3:0] op1_13_in01;
  reg       op1_13_inv01;
  reg [3:0] op1_13_in02;
  reg       op1_13_inv02;
  reg [3:0] op1_13_in03;
  reg       op1_13_inv03;
  reg [3:0] op1_13_in04;
  reg       op1_13_inv04;
  reg [3:0] op1_13_in05;
  reg       op1_13_inv05;
  reg [3:0] op1_13_in06;
  reg       op1_13_inv06;
  reg [3:0] op1_13_in07;
  reg       op1_13_inv07;
  reg [3:0] op1_13_in08;
  reg       op1_13_inv08;
  reg [3:0] op1_13_in09;
  reg       op1_13_inv09;
  reg [3:0] op1_13_in10;
  reg       op1_13_inv10;
  reg [3:0] op1_13_in11;
  reg       op1_13_inv11;
  reg [3:0] op1_13_in12;
  reg       op1_13_inv12;
  reg [3:0] op1_13_in13;
  reg       op1_13_inv13;
  reg [3:0] op1_13_in14;
  reg       op1_13_inv14;
  reg [3:0] op1_13_in15;
  reg       op1_13_inv15;
  reg [3:0] op1_13_in16;
  reg       op1_13_inv16;
  reg [3:0] op1_13_in17;
  reg       op1_13_inv17;
  reg [3:0] op1_13_in18;
  reg       op1_13_inv18;
  reg [3:0] op1_13_in19;
  reg       op1_13_inv19;
  reg [3:0] op1_13_in20;
  reg       op1_13_inv20;
  reg [3:0] op1_13_in21;
  reg       op1_13_inv21;
  reg [3:0] op1_13_in22;
  reg       op1_13_inv22;
  reg [3:0] op1_13_in23;
  reg       op1_13_inv23;
  reg [3:0] op1_13_in24;
  reg       op1_13_inv24;
  reg [3:0] op1_13_in25;
  reg       op1_13_inv25;
  reg [3:0] op1_13_in26;
  reg       op1_13_inv26;
  reg [3:0] op1_13_in27;
  reg       op1_13_inv27;
  reg [3:0] op1_13_in28;
  reg       op1_13_inv28;
  reg [3:0] op1_13_in29;
  reg       op1_13_inv29;
  reg [3:0] op1_13_in30;
  reg       op1_13_inv30;
  reg [3:0] op1_13_in31;
  reg       op1_13_inv31;
  wire [8:0] op1_13_out;
  affine2_op1 op1_13(
    .data0_in(op1_13_in00),
    .inv0_in(op1_13_inv00),
    .data1_in(op1_13_in01),
    .inv1_in(op1_13_inv01),
    .data2_in(op1_13_in02),
    .inv2_in(op1_13_inv02),
    .data3_in(op1_13_in03),
    .inv3_in(op1_13_inv03),
    .data4_in(op1_13_in04),
    .inv4_in(op1_13_inv04),
    .data5_in(op1_13_in05),
    .inv5_in(op1_13_inv05),
    .data6_in(op1_13_in06),
    .inv6_in(op1_13_inv06),
    .data7_in(op1_13_in07),
    .inv7_in(op1_13_inv07),
    .data8_in(op1_13_in08),
    .inv8_in(op1_13_inv08),
    .data9_in(op1_13_in09),
    .inv9_in(op1_13_inv09),
    .data10_in(op1_13_in10),
    .inv10_in(op1_13_inv10),
    .data11_in(op1_13_in11),
    .inv11_in(op1_13_inv11),
    .data12_in(op1_13_in12),
    .inv12_in(op1_13_inv12),
    .data13_in(op1_13_in13),
    .inv13_in(op1_13_inv13),
    .data14_in(op1_13_in14),
    .inv14_in(op1_13_inv14),
    .data15_in(op1_13_in15),
    .inv15_in(op1_13_inv15),
    .data16_in(op1_13_in16),
    .inv16_in(op1_13_inv16),
    .data17_in(op1_13_in17),
    .inv17_in(op1_13_inv17),
    .data18_in(op1_13_in18),
    .inv18_in(op1_13_inv18),
    .data19_in(op1_13_in19),
    .inv19_in(op1_13_inv19),
    .data20_in(op1_13_in20),
    .inv20_in(op1_13_inv20),
    .data21_in(op1_13_in21),
    .inv21_in(op1_13_inv21),
    .data22_in(op1_13_in22),
    .inv22_in(op1_13_inv22),
    .data23_in(op1_13_in23),
    .inv23_in(op1_13_inv23),
    .data24_in(op1_13_in24),
    .inv24_in(op1_13_inv24),
    .data25_in(op1_13_in25),
    .inv25_in(op1_13_inv25),
    .data26_in(op1_13_in26),
    .inv26_in(op1_13_inv26),
    .data27_in(op1_13_in27),
    .inv27_in(op1_13_inv27),
    .data28_in(op1_13_in28),
    .inv28_in(op1_13_inv28),
    .data29_in(op1_13_in29),
    .inv29_in(op1_13_inv29),
    .data30_in(op1_13_in30),
    .inv30_in(op1_13_inv30),
    .data31_in(op1_13_in31),
    .inv31_in(op1_13_inv31),
    .data_out(op1_13_out));

  // 14 番目の OP1
  reg [3:0] op1_14_in00;
  reg       op1_14_inv00;
  reg [3:0] op1_14_in01;
  reg       op1_14_inv01;
  reg [3:0] op1_14_in02;
  reg       op1_14_inv02;
  reg [3:0] op1_14_in03;
  reg       op1_14_inv03;
  reg [3:0] op1_14_in04;
  reg       op1_14_inv04;
  reg [3:0] op1_14_in05;
  reg       op1_14_inv05;
  reg [3:0] op1_14_in06;
  reg       op1_14_inv06;
  reg [3:0] op1_14_in07;
  reg       op1_14_inv07;
  reg [3:0] op1_14_in08;
  reg       op1_14_inv08;
  reg [3:0] op1_14_in09;
  reg       op1_14_inv09;
  reg [3:0] op1_14_in10;
  reg       op1_14_inv10;
  reg [3:0] op1_14_in11;
  reg       op1_14_inv11;
  reg [3:0] op1_14_in12;
  reg       op1_14_inv12;
  reg [3:0] op1_14_in13;
  reg       op1_14_inv13;
  reg [3:0] op1_14_in14;
  reg       op1_14_inv14;
  reg [3:0] op1_14_in15;
  reg       op1_14_inv15;
  reg [3:0] op1_14_in16;
  reg       op1_14_inv16;
  reg [3:0] op1_14_in17;
  reg       op1_14_inv17;
  reg [3:0] op1_14_in18;
  reg       op1_14_inv18;
  reg [3:0] op1_14_in19;
  reg       op1_14_inv19;
  reg [3:0] op1_14_in20;
  reg       op1_14_inv20;
  reg [3:0] op1_14_in21;
  reg       op1_14_inv21;
  reg [3:0] op1_14_in22;
  reg       op1_14_inv22;
  reg [3:0] op1_14_in23;
  reg       op1_14_inv23;
  reg [3:0] op1_14_in24;
  reg       op1_14_inv24;
  reg [3:0] op1_14_in25;
  reg       op1_14_inv25;
  reg [3:0] op1_14_in26;
  reg       op1_14_inv26;
  reg [3:0] op1_14_in27;
  reg       op1_14_inv27;
  reg [3:0] op1_14_in28;
  reg       op1_14_inv28;
  reg [3:0] op1_14_in29;
  reg       op1_14_inv29;
  reg [3:0] op1_14_in30;
  reg       op1_14_inv30;
  reg [3:0] op1_14_in31;
  reg       op1_14_inv31;
  wire [8:0] op1_14_out;
  affine2_op1 op1_14(
    .data0_in(op1_14_in00),
    .inv0_in(op1_14_inv00),
    .data1_in(op1_14_in01),
    .inv1_in(op1_14_inv01),
    .data2_in(op1_14_in02),
    .inv2_in(op1_14_inv02),
    .data3_in(op1_14_in03),
    .inv3_in(op1_14_inv03),
    .data4_in(op1_14_in04),
    .inv4_in(op1_14_inv04),
    .data5_in(op1_14_in05),
    .inv5_in(op1_14_inv05),
    .data6_in(op1_14_in06),
    .inv6_in(op1_14_inv06),
    .data7_in(op1_14_in07),
    .inv7_in(op1_14_inv07),
    .data8_in(op1_14_in08),
    .inv8_in(op1_14_inv08),
    .data9_in(op1_14_in09),
    .inv9_in(op1_14_inv09),
    .data10_in(op1_14_in10),
    .inv10_in(op1_14_inv10),
    .data11_in(op1_14_in11),
    .inv11_in(op1_14_inv11),
    .data12_in(op1_14_in12),
    .inv12_in(op1_14_inv12),
    .data13_in(op1_14_in13),
    .inv13_in(op1_14_inv13),
    .data14_in(op1_14_in14),
    .inv14_in(op1_14_inv14),
    .data15_in(op1_14_in15),
    .inv15_in(op1_14_inv15),
    .data16_in(op1_14_in16),
    .inv16_in(op1_14_inv16),
    .data17_in(op1_14_in17),
    .inv17_in(op1_14_inv17),
    .data18_in(op1_14_in18),
    .inv18_in(op1_14_inv18),
    .data19_in(op1_14_in19),
    .inv19_in(op1_14_inv19),
    .data20_in(op1_14_in20),
    .inv20_in(op1_14_inv20),
    .data21_in(op1_14_in21),
    .inv21_in(op1_14_inv21),
    .data22_in(op1_14_in22),
    .inv22_in(op1_14_inv22),
    .data23_in(op1_14_in23),
    .inv23_in(op1_14_inv23),
    .data24_in(op1_14_in24),
    .inv24_in(op1_14_inv24),
    .data25_in(op1_14_in25),
    .inv25_in(op1_14_inv25),
    .data26_in(op1_14_in26),
    .inv26_in(op1_14_inv26),
    .data27_in(op1_14_in27),
    .inv27_in(op1_14_inv27),
    .data28_in(op1_14_in28),
    .inv28_in(op1_14_inv28),
    .data29_in(op1_14_in29),
    .inv29_in(op1_14_inv29),
    .data30_in(op1_14_in30),
    .inv30_in(op1_14_inv30),
    .data31_in(op1_14_in31),
    .inv31_in(op1_14_inv31),
    .data_out(op1_14_out));

  // 15 番目の OP1
  reg [3:0] op1_15_in00;
  reg       op1_15_inv00;
  reg [3:0] op1_15_in01;
  reg       op1_15_inv01;
  reg [3:0] op1_15_in02;
  reg       op1_15_inv02;
  reg [3:0] op1_15_in03;
  reg       op1_15_inv03;
  reg [3:0] op1_15_in04;
  reg       op1_15_inv04;
  reg [3:0] op1_15_in05;
  reg       op1_15_inv05;
  reg [3:0] op1_15_in06;
  reg       op1_15_inv06;
  reg [3:0] op1_15_in07;
  reg       op1_15_inv07;
  reg [3:0] op1_15_in08;
  reg       op1_15_inv08;
  reg [3:0] op1_15_in09;
  reg       op1_15_inv09;
  reg [3:0] op1_15_in10;
  reg       op1_15_inv10;
  reg [3:0] op1_15_in11;
  reg       op1_15_inv11;
  reg [3:0] op1_15_in12;
  reg       op1_15_inv12;
  reg [3:0] op1_15_in13;
  reg       op1_15_inv13;
  reg [3:0] op1_15_in14;
  reg       op1_15_inv14;
  reg [3:0] op1_15_in15;
  reg       op1_15_inv15;
  reg [3:0] op1_15_in16;
  reg       op1_15_inv16;
  reg [3:0] op1_15_in17;
  reg       op1_15_inv17;
  reg [3:0] op1_15_in18;
  reg       op1_15_inv18;
  reg [3:0] op1_15_in19;
  reg       op1_15_inv19;
  reg [3:0] op1_15_in20;
  reg       op1_15_inv20;
  reg [3:0] op1_15_in21;
  reg       op1_15_inv21;
  reg [3:0] op1_15_in22;
  reg       op1_15_inv22;
  reg [3:0] op1_15_in23;
  reg       op1_15_inv23;
  reg [3:0] op1_15_in24;
  reg       op1_15_inv24;
  reg [3:0] op1_15_in25;
  reg       op1_15_inv25;
  reg [3:0] op1_15_in26;
  reg       op1_15_inv26;
  reg [3:0] op1_15_in27;
  reg       op1_15_inv27;
  reg [3:0] op1_15_in28;
  reg       op1_15_inv28;
  reg [3:0] op1_15_in29;
  reg       op1_15_inv29;
  reg [3:0] op1_15_in30;
  reg       op1_15_inv30;
  reg [3:0] op1_15_in31;
  reg       op1_15_inv31;
  wire [8:0] op1_15_out;
  affine2_op1 op1_15(
    .data0_in(op1_15_in00),
    .inv0_in(op1_15_inv00),
    .data1_in(op1_15_in01),
    .inv1_in(op1_15_inv01),
    .data2_in(op1_15_in02),
    .inv2_in(op1_15_inv02),
    .data3_in(op1_15_in03),
    .inv3_in(op1_15_inv03),
    .data4_in(op1_15_in04),
    .inv4_in(op1_15_inv04),
    .data5_in(op1_15_in05),
    .inv5_in(op1_15_inv05),
    .data6_in(op1_15_in06),
    .inv6_in(op1_15_inv06),
    .data7_in(op1_15_in07),
    .inv7_in(op1_15_inv07),
    .data8_in(op1_15_in08),
    .inv8_in(op1_15_inv08),
    .data9_in(op1_15_in09),
    .inv9_in(op1_15_inv09),
    .data10_in(op1_15_in10),
    .inv10_in(op1_15_inv10),
    .data11_in(op1_15_in11),
    .inv11_in(op1_15_inv11),
    .data12_in(op1_15_in12),
    .inv12_in(op1_15_inv12),
    .data13_in(op1_15_in13),
    .inv13_in(op1_15_inv13),
    .data14_in(op1_15_in14),
    .inv14_in(op1_15_inv14),
    .data15_in(op1_15_in15),
    .inv15_in(op1_15_inv15),
    .data16_in(op1_15_in16),
    .inv16_in(op1_15_inv16),
    .data17_in(op1_15_in17),
    .inv17_in(op1_15_inv17),
    .data18_in(op1_15_in18),
    .inv18_in(op1_15_inv18),
    .data19_in(op1_15_in19),
    .inv19_in(op1_15_inv19),
    .data20_in(op1_15_in20),
    .inv20_in(op1_15_inv20),
    .data21_in(op1_15_in21),
    .inv21_in(op1_15_inv21),
    .data22_in(op1_15_in22),
    .inv22_in(op1_15_inv22),
    .data23_in(op1_15_in23),
    .inv23_in(op1_15_inv23),
    .data24_in(op1_15_in24),
    .inv24_in(op1_15_inv24),
    .data25_in(op1_15_in25),
    .inv25_in(op1_15_inv25),
    .data26_in(op1_15_in26),
    .inv26_in(op1_15_inv26),
    .data27_in(op1_15_in27),
    .inv27_in(op1_15_inv27),
    .data28_in(op1_15_in28),
    .inv28_in(op1_15_inv28),
    .data29_in(op1_15_in29),
    .inv29_in(op1_15_inv29),
    .data30_in(op1_15_in30),
    .inv30_in(op1_15_inv30),
    .data31_in(op1_15_in31),
    .inv31_in(op1_15_inv31),
    .data_out(op1_15_out));

  // 0 番目の OP2
  reg [8:0] op2_00_in00;
  reg [8:0] op2_00_in01;
  reg [8:0] op2_00_in02;
  reg [8:0] op2_00_in03;
  reg [8:0] op2_00_in04;
  reg [8:0] op2_00_in05;
  reg [8:0] op2_00_in06;
  reg [8:0] op2_00_in07;
  reg [8:0] op2_00_in08;
  reg [8:0] op2_00_in09;
  reg [8:0] op2_00_in10;
  reg [8:0] op2_00_in11;
  reg [8:0] op2_00_in12;
  reg [8:0] op2_00_in13;
  reg [8:0] op2_00_in14;
  reg [8:0] op2_00_in15;
  reg [8:0] op2_00_in16;
  reg [8:0] op2_00_in17;
  reg [8:0] op2_00_in18;
  reg [8:0] op2_00_in19;
  reg [8:0] op2_00_in20;
  reg [8:0] op2_00_in21;
  reg [8:0] op2_00_in22;
  reg [8:0] op2_00_in23;
  reg [8:0] op2_00_in24;
  reg [8:0] op2_00_in25;
  reg [8:0] op2_00_in26;
  reg [8:0] op2_00_in27;
  reg [8:0] op2_00_in28;
  reg [8:0] op2_00_in29;
  reg [8:0] op2_00_in30;
  reg [8:0] op2_00_bias;
  wire [8:0] op2_00_out;
  affine2_op2 op2_00(
    .data0_in(op2_00_in00),
    .data1_in(op2_00_in01),
    .data2_in(op2_00_in02),
    .data3_in(op2_00_in03),
    .data4_in(op2_00_in04),
    .data5_in(op2_00_in05),
    .data6_in(op2_00_in06),
    .data7_in(op2_00_in07),
    .data8_in(op2_00_in08),
    .data9_in(op2_00_in09),
    .data10_in(op2_00_in10),
    .data11_in(op2_00_in11),
    .data12_in(op2_00_in12),
    .data13_in(op2_00_in13),
    .data14_in(op2_00_in14),
    .data15_in(op2_00_in15),
    .data16_in(op2_00_in16),
    .data17_in(op2_00_in17),
    .data18_in(op2_00_in18),
    .data19_in(op2_00_in19),
    .data20_in(op2_00_in20),
    .data21_in(op2_00_in21),
    .data22_in(op2_00_in22),
    .data23_in(op2_00_in23),
    .data24_in(op2_00_in24),
    .data25_in(op2_00_in25),
    .data26_in(op2_00_in26),
    .data27_in(op2_00_in27),
    .data28_in(op2_00_in28),
    .data29_in(op2_00_in29),
    .data30_in(op2_00_in30),
    .data31_in(op2_00_bias),
    .data_out(op2_00_out));

  // 1 番目の OP2
  reg [8:0] op2_01_in00;
  reg [8:0] op2_01_in01;
  reg [8:0] op2_01_in02;
  reg [8:0] op2_01_in03;
  reg [8:0] op2_01_in04;
  reg [8:0] op2_01_in05;
  reg [8:0] op2_01_in06;
  reg [8:0] op2_01_in07;
  reg [8:0] op2_01_in08;
  reg [8:0] op2_01_in09;
  reg [8:0] op2_01_in10;
  reg [8:0] op2_01_in11;
  reg [8:0] op2_01_in12;
  reg [8:0] op2_01_in13;
  reg [8:0] op2_01_in14;
  reg [8:0] op2_01_in15;
  reg [8:0] op2_01_in16;
  reg [8:0] op2_01_in17;
  reg [8:0] op2_01_in18;
  reg [8:0] op2_01_in19;
  reg [8:0] op2_01_in20;
  reg [8:0] op2_01_in21;
  reg [8:0] op2_01_in22;
  reg [8:0] op2_01_in23;
  reg [8:0] op2_01_in24;
  reg [8:0] op2_01_in25;
  reg [8:0] op2_01_in26;
  reg [8:0] op2_01_in27;
  reg [8:0] op2_01_in28;
  reg [8:0] op2_01_in29;
  reg [8:0] op2_01_in30;
  reg [8:0] op2_01_bias;
  wire [8:0] op2_01_out;
  affine2_op2 op2_01(
    .data0_in(op2_01_in00),
    .data1_in(op2_01_in01),
    .data2_in(op2_01_in02),
    .data3_in(op2_01_in03),
    .data4_in(op2_01_in04),
    .data5_in(op2_01_in05),
    .data6_in(op2_01_in06),
    .data7_in(op2_01_in07),
    .data8_in(op2_01_in08),
    .data9_in(op2_01_in09),
    .data10_in(op2_01_in10),
    .data11_in(op2_01_in11),
    .data12_in(op2_01_in12),
    .data13_in(op2_01_in13),
    .data14_in(op2_01_in14),
    .data15_in(op2_01_in15),
    .data16_in(op2_01_in16),
    .data17_in(op2_01_in17),
    .data18_in(op2_01_in18),
    .data19_in(op2_01_in19),
    .data20_in(op2_01_in20),
    .data21_in(op2_01_in21),
    .data22_in(op2_01_in22),
    .data23_in(op2_01_in23),
    .data24_in(op2_01_in24),
    .data25_in(op2_01_in25),
    .data26_in(op2_01_in26),
    .data27_in(op2_01_in27),
    .data28_in(op2_01_in28),
    .data29_in(op2_01_in29),
    .data30_in(op2_01_in30),
    .data31_in(op2_01_bias),
    .data_out(op2_01_out));

  // 2 番目の OP2
  reg [8:0] op2_02_in00;
  reg [8:0] op2_02_in01;
  reg [8:0] op2_02_in02;
  reg [8:0] op2_02_in03;
  reg [8:0] op2_02_in04;
  reg [8:0] op2_02_in05;
  reg [8:0] op2_02_in06;
  reg [8:0] op2_02_in07;
  reg [8:0] op2_02_in08;
  reg [8:0] op2_02_in09;
  reg [8:0] op2_02_in10;
  reg [8:0] op2_02_in11;
  reg [8:0] op2_02_in12;
  reg [8:0] op2_02_in13;
  reg [8:0] op2_02_in14;
  reg [8:0] op2_02_in15;
  reg [8:0] op2_02_in16;
  reg [8:0] op2_02_in17;
  reg [8:0] op2_02_in18;
  reg [8:0] op2_02_in19;
  reg [8:0] op2_02_in20;
  reg [8:0] op2_02_in21;
  reg [8:0] op2_02_in22;
  reg [8:0] op2_02_in23;
  reg [8:0] op2_02_in24;
  reg [8:0] op2_02_in25;
  reg [8:0] op2_02_in26;
  reg [8:0] op2_02_in27;
  reg [8:0] op2_02_in28;
  reg [8:0] op2_02_in29;
  reg [8:0] op2_02_in30;
  reg [8:0] op2_02_bias;
  wire [8:0] op2_02_out;
  affine2_op2 op2_02(
    .data0_in(op2_02_in00),
    .data1_in(op2_02_in01),
    .data2_in(op2_02_in02),
    .data3_in(op2_02_in03),
    .data4_in(op2_02_in04),
    .data5_in(op2_02_in05),
    .data6_in(op2_02_in06),
    .data7_in(op2_02_in07),
    .data8_in(op2_02_in08),
    .data9_in(op2_02_in09),
    .data10_in(op2_02_in10),
    .data11_in(op2_02_in11),
    .data12_in(op2_02_in12),
    .data13_in(op2_02_in13),
    .data14_in(op2_02_in14),
    .data15_in(op2_02_in15),
    .data16_in(op2_02_in16),
    .data17_in(op2_02_in17),
    .data18_in(op2_02_in18),
    .data19_in(op2_02_in19),
    .data20_in(op2_02_in20),
    .data21_in(op2_02_in21),
    .data22_in(op2_02_in22),
    .data23_in(op2_02_in23),
    .data24_in(op2_02_in24),
    .data25_in(op2_02_in25),
    .data26_in(op2_02_in26),
    .data27_in(op2_02_in27),
    .data28_in(op2_02_in28),
    .data29_in(op2_02_in29),
    .data30_in(op2_02_in30),
    .data31_in(op2_02_bias),
    .data_out(op2_02_out));

  // 3 番目の OP2
  reg [8:0] op2_03_in00;
  reg [8:0] op2_03_in01;
  reg [8:0] op2_03_in02;
  reg [8:0] op2_03_in03;
  reg [8:0] op2_03_in04;
  reg [8:0] op2_03_in05;
  reg [8:0] op2_03_in06;
  reg [8:0] op2_03_in07;
  reg [8:0] op2_03_in08;
  reg [8:0] op2_03_in09;
  reg [8:0] op2_03_in10;
  reg [8:0] op2_03_in11;
  reg [8:0] op2_03_in12;
  reg [8:0] op2_03_in13;
  reg [8:0] op2_03_in14;
  reg [8:0] op2_03_in15;
  reg [8:0] op2_03_in16;
  reg [8:0] op2_03_in17;
  reg [8:0] op2_03_in18;
  reg [8:0] op2_03_in19;
  reg [8:0] op2_03_in20;
  reg [8:0] op2_03_in21;
  reg [8:0] op2_03_in22;
  reg [8:0] op2_03_in23;
  reg [8:0] op2_03_in24;
  reg [8:0] op2_03_in25;
  reg [8:0] op2_03_in26;
  reg [8:0] op2_03_in27;
  reg [8:0] op2_03_in28;
  reg [8:0] op2_03_in29;
  reg [8:0] op2_03_in30;
  reg [8:0] op2_03_bias;
  wire [8:0] op2_03_out;
  affine2_op2 op2_03(
    .data0_in(op2_03_in00),
    .data1_in(op2_03_in01),
    .data2_in(op2_03_in02),
    .data3_in(op2_03_in03),
    .data4_in(op2_03_in04),
    .data5_in(op2_03_in05),
    .data6_in(op2_03_in06),
    .data7_in(op2_03_in07),
    .data8_in(op2_03_in08),
    .data9_in(op2_03_in09),
    .data10_in(op2_03_in10),
    .data11_in(op2_03_in11),
    .data12_in(op2_03_in12),
    .data13_in(op2_03_in13),
    .data14_in(op2_03_in14),
    .data15_in(op2_03_in15),
    .data16_in(op2_03_in16),
    .data17_in(op2_03_in17),
    .data18_in(op2_03_in18),
    .data19_in(op2_03_in19),
    .data20_in(op2_03_in20),
    .data21_in(op2_03_in21),
    .data22_in(op2_03_in22),
    .data23_in(op2_03_in23),
    .data24_in(op2_03_in24),
    .data25_in(op2_03_in25),
    .data26_in(op2_03_in26),
    .data27_in(op2_03_in27),
    .data28_in(op2_03_in28),
    .data29_in(op2_03_in29),
    .data30_in(op2_03_in30),
    .data31_in(op2_03_bias),
    .data_out(op2_03_out));

  // 中間レジスタ
  reg [8:0] reg_0000;
  reg [8:0] reg_0001;
  reg [8:0] reg_0002;
  reg [8:0] reg_0003;
  reg [8:0] reg_0004;
  reg [8:0] reg_0005;
  reg [8:0] reg_0006;
  reg [8:0] reg_0007;
  reg [8:0] reg_0008;
  reg [8:0] reg_0009;
  reg [8:0] reg_0010;
  reg [8:0] reg_0011;
  reg [8:0] reg_0012;
  reg [8:0] reg_0013;
  reg [8:0] reg_0014;
  reg [8:0] reg_0015;
  reg [8:0] reg_0016;
  reg [8:0] reg_0017;
  reg [8:0] reg_0018;
  reg [8:0] reg_0019;
  reg [8:0] reg_0020;
  reg [8:0] reg_0021;
  reg [8:0] reg_0022;
  reg [8:0] reg_0023;
  reg [8:0] reg_0024;
  reg [8:0] reg_0025;
  reg [8:0] reg_0026;
  reg [8:0] reg_0027;
  reg [8:0] reg_0028;
  reg [8:0] reg_0029;
  reg [8:0] reg_0030;
  reg [8:0] reg_0031;
  reg [8:0] reg_0032;
  reg [8:0] reg_0033;
  reg [8:0] reg_0034;
  reg [8:0] reg_0035;
  reg [8:0] reg_0036;
  reg [8:0] reg_0037;
  reg [8:0] reg_0038;
  reg [8:0] reg_0039;
  reg [8:0] reg_0040;
  reg [8:0] reg_0041;
  reg [8:0] reg_0042;
  reg [8:0] reg_0043;
  reg [8:0] reg_0044;
  reg [8:0] reg_0045;
  reg [8:0] reg_0046;
  reg [8:0] reg_0047;
  reg [8:0] reg_0048;
  reg [8:0] reg_0049;
  reg [8:0] reg_0050;
  reg [8:0] reg_0051;
  reg [8:0] reg_0052;
  reg [8:0] reg_0053;
  reg [8:0] reg_0054;
  reg [8:0] reg_0055;
  reg [8:0] reg_0056;
  reg [8:0] reg_0057;
  reg [8:0] reg_0058;
  reg [8:0] reg_0059;
  reg [8:0] reg_0060;
  reg [8:0] reg_0061;
  reg [8:0] reg_0062;
  reg [8:0] reg_0063;
  reg [8:0] reg_0064;
  reg [8:0] reg_0065;
  reg [8:0] reg_0066;
  reg [8:0] reg_0067;
  reg [8:0] reg_0068;
  reg [8:0] reg_0069;
  reg [8:0] reg_0070;
  reg [8:0] reg_0071;
  reg [8:0] reg_0072;
  reg [8:0] reg_0073;
  reg [8:0] reg_0074;
  reg [8:0] reg_0075;
  reg [8:0] reg_0076;
  reg [8:0] reg_0077;
  reg [8:0] reg_0078;
  reg [8:0] reg_0079;
  reg [8:0] reg_0080;
  reg [8:0] reg_0081;
  reg [8:0] reg_0082;
  reg [8:0] reg_0083;
  reg [8:0] reg_0084;
  reg [8:0] reg_0085;
  reg [8:0] reg_0086;
  reg [8:0] reg_0087;
  reg [8:0] reg_0088;
  reg [8:0] reg_0089;
  reg [8:0] reg_0090;
  reg [8:0] reg_0091;
  reg [8:0] reg_0092;
  reg [8:0] reg_0093;
  reg [8:0] reg_0094;
  reg [8:0] reg_0095;
  reg [8:0] reg_0096;
  reg [8:0] reg_0097;
  reg [8:0] reg_0098;
  reg [8:0] reg_0099;
  reg [8:0] reg_0100;
  reg [8:0] reg_0101;
  reg [8:0] reg_0102;
  reg [8:0] reg_0103;
  reg [8:0] reg_0104;
  reg [8:0] reg_0105;
  reg [8:0] reg_0106;
  reg [8:0] reg_0107;
  reg [8:0] reg_0108;
  reg [8:0] reg_0109;
  reg [8:0] reg_0110;
  reg [8:0] reg_0111;
  reg [8:0] reg_0112;
  reg [8:0] reg_0113;
  reg [8:0] reg_0114;
  reg [8:0] reg_0115;
  reg [8:0] reg_0116;
  reg [8:0] reg_0117;
  reg [8:0] reg_0118;
  reg [8:0] reg_0119;
  reg [8:0] reg_0120;
  reg [8:0] reg_0121;
  reg [8:0] reg_0122;
  reg [8:0] reg_0123;
  reg [8:0] reg_0124;
  reg [8:0] reg_0125;
  reg [8:0] reg_0126;
  reg [8:0] reg_0127;
  reg [8:0] reg_0128;
  reg [8:0] reg_0129;
  reg [8:0] reg_0130;
  reg [8:0] reg_0131;
  reg [8:0] reg_0132;
  reg [8:0] reg_0133;
  reg [8:0] reg_0134;
  reg [8:0] reg_0135;
  reg [8:0] reg_0136;
  reg [8:0] reg_0137;
  reg [8:0] reg_0138;
  reg [8:0] reg_0139;
  reg [8:0] reg_0140;
  reg [8:0] reg_0141;
  reg [8:0] reg_0142;
  reg [8:0] reg_0143;
  reg [8:0] reg_0144;
  reg [8:0] reg_0145;
  reg [8:0] reg_0146;
  reg [8:0] reg_0147;
  reg [8:0] reg_0148;
  reg [8:0] reg_0149;
  reg [8:0] reg_0150;
  reg [8:0] reg_0151;
  reg [8:0] reg_0152;
  reg [8:0] reg_0153;
  reg [8:0] reg_0154;
  reg [8:0] reg_0155;
  reg [8:0] reg_0156;
  reg [8:0] reg_0157;
  reg [8:0] reg_0158;
  reg [8:0] reg_0159;
  reg [8:0] reg_0160;
  reg [8:0] reg_0161;
  reg [8:0] reg_0162;
  reg [8:0] reg_0163;
  reg [8:0] reg_0164;
  reg [8:0] reg_0165;
  reg [8:0] reg_0166;
  reg [8:0] reg_0167;
  reg [8:0] reg_0168;
  reg [8:0] reg_0169;
  reg [8:0] reg_0170;
  reg [8:0] reg_0171;
  reg [8:0] reg_0172;
  reg [8:0] reg_0173;
  reg [8:0] reg_0174;
  reg [8:0] reg_0175;
  reg [8:0] reg_0176;
  reg [8:0] reg_0177;
  reg [8:0] reg_0178;
  reg [8:0] reg_0179;
  reg [8:0] reg_0180;
  reg [8:0] reg_0181;
  reg [8:0] reg_0182;
  reg [8:0] reg_0183;
  reg [8:0] reg_0184;
  reg [8:0] reg_0185;
  reg [8:0] reg_0186;
  reg [8:0] reg_0187;
  reg [8:0] reg_0188;
  reg [8:0] reg_0189;
  reg [8:0] reg_0190;
  reg [8:0] reg_0191;
  reg [8:0] reg_0192;
  reg [8:0] reg_0193;
  reg [8:0] reg_0194;
  reg [8:0] reg_0195;
  reg [8:0] reg_0196;
  reg [8:0] reg_0197;
  reg [8:0] reg_0198;
  reg [8:0] reg_0199;
  reg [8:0] reg_0200;
  reg [8:0] reg_0201;
  reg [8:0] reg_0202;
  reg [8:0] reg_0203;
  reg [8:0] reg_0204;
  reg [8:0] reg_0205;
  reg [8:0] reg_0206;
  reg [8:0] reg_0207;
  reg [8:0] reg_0208;
  reg [8:0] reg_0209;
  reg [8:0] reg_0210;
  reg [8:0] reg_0211;
  reg [8:0] reg_0212;
  reg [8:0] reg_0213;
  reg [8:0] reg_0214;
  reg [8:0] reg_0215;
  reg [8:0] reg_0216;
  reg [8:0] reg_0217;
  reg [8:0] reg_0218;
  reg [8:0] reg_0219;
  reg [8:0] reg_0220;
  reg [8:0] reg_0221;
  reg [8:0] reg_0222;
  reg [8:0] reg_0223;
  reg [8:0] reg_0224;
  reg [8:0] reg_0225;
  reg [8:0] reg_0226;
  reg [8:0] reg_0227;
  reg [8:0] reg_0228;
  reg [8:0] reg_0229;
  reg [8:0] reg_0230;
  reg [8:0] reg_0231;
  reg [8:0] reg_0232;
  reg [8:0] reg_0233;
  reg [8:0] reg_0234;
  reg [8:0] reg_0235;
  reg [8:0] reg_0236;
  reg [8:0] reg_0237;
  reg [8:0] reg_0238;
  reg [8:0] reg_0239;
  reg [8:0] reg_0240;
  reg [8:0] reg_0241;
  reg [8:0] reg_0242;
  reg [8:0] reg_0243;
  reg [8:0] reg_0244;
  reg [8:0] reg_0245;
  reg [8:0] reg_0246;
  reg [8:0] reg_0247;
  reg [8:0] reg_0248;
  reg [8:0] reg_0249;
  reg [8:0] reg_0250;
  reg [8:0] reg_0251;
  reg [8:0] reg_0252;
  reg [8:0] reg_0253;
  reg [8:0] reg_0254;
  reg [8:0] reg_0255;
  reg [8:0] reg_0256;
  reg [8:0] reg_0257;
  reg [8:0] reg_0258;
  reg [8:0] reg_0259;
  reg [8:0] reg_0260;
  reg [8:0] reg_0261;
  reg [8:0] reg_0262;
  reg [8:0] reg_0263;
  reg [8:0] reg_0264;
  reg [8:0] reg_0265;
  reg [8:0] reg_0266;
  reg [8:0] reg_0267;
  reg [8:0] reg_0268;
  reg [8:0] reg_0269;
  reg [8:0] reg_0270;
  reg [8:0] reg_0271;
  reg [8:0] reg_0272;
  reg [8:0] reg_0273;
  reg [8:0] reg_0274;
  reg [8:0] reg_0275;
  reg [8:0] reg_0276;
  reg [8:0] reg_0277;
  reg [8:0] reg_0278;
  reg [8:0] reg_0279;
  reg [8:0] reg_0280;
  reg [8:0] reg_0281;
  reg [8:0] reg_0282;
  reg [8:0] reg_0283;
  reg [8:0] reg_0284;
  reg [8:0] reg_0285;
  reg [8:0] reg_0286;
  reg [8:0] reg_0287;
  reg [8:0] reg_0288;
  reg [8:0] reg_0289;
  reg [8:0] reg_0290;
  reg [8:0] reg_0291;
  reg [8:0] reg_0292;
  reg [8:0] reg_0293;
  reg [8:0] reg_0294;
  reg [8:0] reg_0295;
  reg [8:0] reg_0296;
  reg [8:0] reg_0297;
  reg [8:0] reg_0298;
  reg [8:0] reg_0299;
  reg [8:0] reg_0300;
  reg [8:0] reg_0301;
  reg [8:0] reg_0302;
  reg [8:0] reg_0303;
  reg [8:0] reg_0304;
  reg [8:0] reg_0305;
  reg [8:0] reg_0306;
  reg [8:0] reg_0307;
  reg [8:0] reg_0308;
  reg [8:0] reg_0309;
  reg [8:0] reg_0310;
  reg [8:0] reg_0311;
  reg [8:0] reg_0312;
  reg [8:0] reg_0313;
  reg [8:0] reg_0314;
  reg [8:0] reg_0315;
  reg [8:0] reg_0316;
  reg [8:0] reg_0317;
  reg [8:0] reg_0318;
  reg [8:0] reg_0319;
  reg [8:0] reg_0320;
  reg [8:0] reg_0321;
  reg [8:0] reg_0322;
  reg [8:0] reg_0323;
  reg [8:0] reg_0324;
  reg [8:0] reg_0325;
  reg [8:0] reg_0326;
  reg [8:0] reg_0327;
  reg [8:0] reg_0328;
  reg [8:0] reg_0329;
  reg [8:0] reg_0330;
  reg [8:0] reg_0331;
  reg [8:0] reg_0332;
  reg [8:0] reg_0333;
  reg [8:0] reg_0334;
  reg [8:0] reg_0335;
  reg [8:0] reg_0336;
  reg [8:0] reg_0337;
  reg [8:0] reg_0338;
  reg [8:0] reg_0339;
  reg [8:0] reg_0340;
  reg [8:0] reg_0341;
  reg [8:0] reg_0342;
  reg [8:0] reg_0343;
  reg [8:0] reg_0344;
  reg [8:0] reg_0345;
  reg [8:0] reg_0346;
  reg [8:0] reg_0347;
  reg [8:0] reg_0348;
  reg [8:0] reg_0349;
  reg [8:0] reg_0350;
  reg [8:0] reg_0351;
  reg [8:0] reg_0352;
  reg [8:0] reg_0353;
  reg [8:0] reg_0354;
  reg [8:0] reg_0355;
  reg [8:0] reg_0356;
  reg [8:0] reg_0357;
  reg [8:0] reg_0358;
  reg [8:0] reg_0359;
  reg [8:0] reg_0360;
  reg [8:0] reg_0361;
  reg [8:0] reg_0362;
  reg [8:0] reg_0363;
  reg [8:0] reg_0364;
  reg [8:0] reg_0365;
  reg [8:0] reg_0366;
  reg [8:0] reg_0367;
  reg [8:0] reg_0368;
  reg [8:0] reg_0369;
  reg [8:0] reg_0370;
  reg [8:0] reg_0371;
  reg [8:0] reg_0372;
  reg [8:0] reg_0373;
  reg [8:0] reg_0374;
  reg [8:0] reg_0375;
  reg [8:0] reg_0376;
  reg [8:0] reg_0377;
  reg [8:0] reg_0378;
  reg [8:0] reg_0379;
  reg [8:0] reg_0380;
  reg [8:0] reg_0381;
  reg [8:0] reg_0382;
  reg [8:0] reg_0383;
  reg [8:0] reg_0384;
  reg [8:0] reg_0385;
  reg [8:0] reg_0386;
  reg [8:0] reg_0387;
  reg [8:0] reg_0388;
  reg [8:0] reg_0389;
  reg [8:0] reg_0390;
  reg [8:0] reg_0391;
  reg [8:0] reg_0392;
  reg [8:0] reg_0393;
  reg [8:0] reg_0394;
  reg [8:0] reg_0395;
  reg [8:0] reg_0396;
  reg [8:0] reg_0397;
  reg [8:0] reg_0398;
  reg [8:0] reg_0399;
  reg [8:0] reg_0400;
  reg [8:0] reg_0401;
  reg [8:0] reg_0402;
  reg [8:0] reg_0403;
  reg [8:0] reg_0404;
  reg [8:0] reg_0405;
  reg [8:0] reg_0406;
  reg [8:0] reg_0407;
  reg [8:0] reg_0408;
  reg [8:0] reg_0409;
  reg [8:0] reg_0410;
  reg [8:0] reg_0411;
  reg [8:0] reg_0412;
  reg [8:0] reg_0413;
  reg [8:0] reg_0414;
  reg [8:0] reg_0415;
  reg [8:0] reg_0416;
  reg [8:0] reg_0417;
  reg [8:0] reg_0418;
  reg [8:0] reg_0419;
  reg [8:0] reg_0420;
  reg [8:0] reg_0421;
  reg [8:0] reg_0422;
  reg [8:0] reg_0423;
  reg [8:0] reg_0424;
  reg [8:0] reg_0425;
  reg [8:0] reg_0426;
  reg [8:0] reg_0427;
  reg [8:0] reg_0428;
  reg [8:0] reg_0429;
  reg [8:0] reg_0430;
  reg [8:0] reg_0431;
  reg [8:0] reg_0432;
  reg [8:0] reg_0433;
  reg [8:0] reg_0434;
  reg [8:0] reg_0435;
  reg [8:0] reg_0436;
  reg [8:0] reg_0437;
  reg [8:0] reg_0438;
  reg [8:0] reg_0439;
  reg [8:0] reg_0440;
  reg [8:0] reg_0441;
  reg [8:0] reg_0442;
  reg [8:0] reg_0443;
  reg [8:0] reg_0444;
  reg [8:0] reg_0445;
  reg [8:0] reg_0446;
  reg [8:0] reg_0447;
  reg [8:0] reg_0448;
  reg [8:0] reg_0449;
  reg [8:0] reg_0450;
  reg [8:0] reg_0451;
  reg [8:0] reg_0452;
  reg [8:0] reg_0453;
  reg [8:0] reg_0454;
  reg [8:0] reg_0455;
  reg [8:0] reg_0456;
  reg [8:0] reg_0457;
  reg [8:0] reg_0458;
  reg [8:0] reg_0459;
  reg [8:0] reg_0460;
  reg [8:0] reg_0461;
  reg [8:0] reg_0462;
  reg [8:0] reg_0463;
  reg [8:0] reg_0464;
  reg [8:0] reg_0465;
  reg [8:0] reg_0466;
  reg [8:0] reg_0467;
  reg [8:0] reg_0468;
  reg [8:0] reg_0469;
  reg [8:0] reg_0470;
  reg [8:0] reg_0471;
  reg [8:0] reg_0472;
  reg [8:0] reg_0473;
  reg [8:0] reg_0474;
  reg [8:0] reg_0475;
  reg [8:0] reg_0476;
  reg [8:0] reg_0477;
  reg [8:0] reg_0478;
  reg [8:0] reg_0479;
  reg [8:0] reg_0480;
  reg [8:0] reg_0481;
  reg [8:0] reg_0482;
  reg [8:0] reg_0483;
  reg [8:0] reg_0484;
  reg [8:0] reg_0485;
  reg [8:0] reg_0486;
  reg [8:0] reg_0487;
  reg [8:0] reg_0488;
  reg [8:0] reg_0489;
  reg [8:0] reg_0490;
  reg [8:0] reg_0491;
  reg [8:0] reg_0492;
  reg [8:0] reg_0493;
  reg [8:0] reg_0494;
  reg [8:0] reg_0495;
  reg [8:0] reg_0496;
  reg [8:0] reg_0497;
  reg [8:0] reg_0498;
  reg [8:0] reg_0499;
  reg [8:0] reg_0500;
  reg [8:0] reg_0501;
  reg [8:0] reg_0502;
  reg [8:0] reg_0503;
  reg [8:0] reg_0504;
  reg [8:0] reg_0505;
  reg [8:0] reg_0506;
  reg [8:0] reg_0507;
  reg [8:0] reg_0508;
  reg [8:0] reg_0509;
  reg [8:0] reg_0510;
  reg [8:0] reg_0511;
  reg [8:0] reg_0512;
  reg [8:0] reg_0513;
  reg [8:0] reg_0514;
  reg [8:0] reg_0515;
  reg [8:0] reg_0516;
  reg [8:0] reg_0517;
  reg [8:0] reg_0518;
  reg [8:0] reg_0519;
  reg [8:0] reg_0520;
  reg [8:0] reg_0521;
  reg [8:0] reg_0522;
  reg [8:0] reg_0523;
  reg [8:0] reg_0524;
  reg [8:0] reg_0525;
  reg [8:0] reg_0526;
  reg [8:0] reg_0527;
  reg [8:0] reg_0528;
  reg [8:0] reg_0529;
  reg [8:0] reg_0530;
  reg [8:0] reg_0531;
  reg [8:0] reg_0532;
  reg [8:0] reg_0533;
  reg [8:0] reg_0534;
  reg [8:0] reg_0535;
  reg [8:0] reg_0536;
  reg [8:0] reg_0537;
  reg [8:0] reg_0538;
  reg [8:0] reg_0539;
  reg [8:0] reg_0540;
  reg [8:0] reg_0541;
  reg [8:0] reg_0542;
  reg [8:0] reg_0543;
  reg [8:0] reg_0544;
  reg [8:0] reg_0545;
  reg [8:0] reg_0546;
  reg [8:0] reg_0547;
  reg [8:0] reg_0548;
  reg [8:0] reg_0549;
  reg [8:0] reg_0550;
  reg [8:0] reg_0551;
  reg [8:0] reg_0552;
  reg [8:0] reg_0553;
  reg [8:0] reg_0554;
  reg [8:0] reg_0555;
  reg [8:0] reg_0556;
  reg [8:0] reg_0557;
  reg [8:0] reg_0558;
  reg [8:0] reg_0559;
  reg [8:0] reg_0560;
  reg [8:0] reg_0561;
  reg [8:0] reg_0562;
  reg [8:0] reg_0563;
  reg [8:0] reg_0564;
  reg [8:0] reg_0565;
  reg [8:0] reg_0566;
  reg [8:0] reg_0567;
  reg [8:0] reg_0568;
  reg [8:0] reg_0569;
  reg [8:0] reg_0570;
  reg [8:0] reg_0571;
  reg [8:0] reg_0572;
  reg [8:0] reg_0573;
  reg [8:0] reg_0574;
  reg [8:0] reg_0575;
  reg [8:0] reg_0576;
  reg [8:0] reg_0577;
  reg [8:0] reg_0578;
  reg [8:0] reg_0579;
  reg [8:0] reg_0580;
  reg [8:0] reg_0581;
  reg [8:0] reg_0582;
  reg [8:0] reg_0583;
  reg [8:0] reg_0584;
  reg [8:0] reg_0585;
  reg [8:0] reg_0586;
  reg [8:0] reg_0587;
  reg [8:0] reg_0588;
  reg [8:0] reg_0589;
  reg [8:0] reg_0590;
  reg [8:0] reg_0591;
  reg [8:0] reg_0592;
  reg [8:0] reg_0593;
  reg [8:0] reg_0594;
  reg [8:0] reg_0595;
  reg [8:0] reg_0596;
  reg [8:0] reg_0597;
  reg [8:0] reg_0598;
  reg [8:0] reg_0599;
  reg [8:0] reg_0600;
  reg [8:0] reg_0601;
  reg [8:0] reg_0602;
  reg [8:0] reg_0603;
  reg [8:0] reg_0604;
  reg [8:0] reg_0605;
  reg [8:0] reg_0606;
  reg [8:0] reg_0607;
  reg [8:0] reg_0608;
  reg [8:0] reg_0609;
  reg [8:0] reg_0610;
  reg [8:0] reg_0611;
  reg [8:0] reg_0612;
  reg [8:0] reg_0613;
  reg [8:0] reg_0614;
  reg [8:0] reg_0615;
  reg [8:0] reg_0616;
  reg [8:0] reg_0617;
  reg [8:0] reg_0618;
  reg [8:0] reg_0619;
  reg [8:0] reg_0620;
  reg [8:0] reg_0621;
  reg [8:0] reg_0622;
  reg [8:0] reg_0623;
  reg [8:0] reg_0624;
  reg [8:0] reg_0625;
  reg [8:0] reg_0626;
  reg [8:0] reg_0627;
  reg [8:0] reg_0628;
  reg [8:0] reg_0629;
  reg [8:0] reg_0630;
  reg [8:0] reg_0631;
  reg [8:0] reg_0632;
  reg [8:0] reg_0633;
  reg [8:0] reg_0634;
  reg [8:0] reg_0635;
  reg [8:0] reg_0636;
  reg [8:0] reg_0637;
  reg [8:0] reg_0638;
  reg [8:0] reg_0639;
  reg [8:0] reg_0640;
  reg [8:0] reg_0641;
  reg [8:0] reg_0642;
  reg [8:0] reg_0643;
  reg [8:0] reg_0644;
  reg [8:0] reg_0645;
  reg [8:0] reg_0646;
  reg [8:0] reg_0647;
  reg [8:0] reg_0648;
  reg [8:0] reg_0649;
  reg [8:0] reg_0650;
  reg [8:0] reg_0651;
  reg [8:0] reg_0652;
  reg [8:0] reg_0653;
  reg [8:0] reg_0654;
  reg [8:0] reg_0655;
  reg [8:0] reg_0656;
  reg [8:0] reg_0657;
  reg [8:0] reg_0658;
  reg [8:0] reg_0659;
  reg [8:0] reg_0660;
  reg [8:0] reg_0661;
  reg [8:0] reg_0662;
  reg [8:0] reg_0663;
  reg [8:0] reg_0664;
  reg [8:0] reg_0665;
  reg [8:0] reg_0666;
  reg [8:0] reg_0667;
  reg [8:0] reg_0668;
  reg [8:0] reg_0669;
  reg [8:0] reg_0670;
  reg [8:0] reg_0671;
  reg [8:0] reg_0672;
  reg [8:0] reg_0673;
  reg [8:0] reg_0674;
  reg [8:0] reg_0675;
  reg [8:0] reg_0676;
  reg [8:0] reg_0677;
  reg [8:0] reg_0678;
  reg [8:0] reg_0679;
  reg [8:0] reg_0680;
  reg [8:0] reg_0681;
  reg [8:0] reg_0682;
  reg [8:0] reg_0683;
  reg [8:0] reg_0684;
  reg [8:0] reg_0685;
  reg [8:0] reg_0686;
  reg [8:0] reg_0687;
  reg [8:0] reg_0688;
  reg [8:0] reg_0689;
  reg [8:0] reg_0690;
  reg [8:0] reg_0691;
  reg [8:0] reg_0692;
  reg [8:0] reg_0693;
  reg [8:0] reg_0694;
  reg [8:0] reg_0695;
  reg [8:0] reg_0696;
  reg [8:0] reg_0697;
  reg [8:0] reg_0698;
  reg [8:0] reg_0699;
  reg [8:0] reg_0700;
  reg [8:0] reg_0701;
  reg [8:0] reg_0702;
  reg [8:0] reg_0703;
  reg [8:0] reg_0704;
  reg [8:0] reg_0705;
  reg [8:0] reg_0706;
  reg [8:0] reg_0707;
  reg [8:0] reg_0708;
  reg [8:0] reg_0709;
  reg [8:0] reg_0710;
  reg [8:0] reg_0711;
  reg [8:0] reg_0712;
  reg [8:0] reg_0713;
  reg [8:0] reg_0714;
  reg [8:0] reg_0715;
  reg [8:0] reg_0716;
  reg [8:0] reg_0717;
  reg [8:0] reg_0718;
  reg [8:0] reg_0719;
  reg [8:0] reg_0720;
  reg [8:0] reg_0721;
  reg [8:0] reg_0722;
  reg [8:0] reg_0723;
  reg [8:0] reg_0724;
  reg [8:0] reg_0725;
  reg [8:0] reg_0726;
  reg [8:0] reg_0727;
  reg [8:0] reg_0728;
  reg [8:0] reg_0729;
  reg [8:0] reg_0730;
  reg [8:0] reg_0731;
  reg [8:0] reg_0732;
  reg [8:0] reg_0733;
  reg [8:0] reg_0734;
  reg [8:0] reg_0735;
  reg [8:0] reg_0736;
  reg [8:0] reg_0737;
  reg [8:0] reg_0738;
  reg [8:0] reg_0739;
  reg [8:0] reg_0740;
  reg [8:0] reg_0741;
  reg [8:0] reg_0742;
  reg [8:0] reg_0743;
  reg [8:0] reg_0744;
  reg [8:0] reg_0745;
  reg [8:0] reg_0746;
  reg [8:0] reg_0747;
  reg [8:0] reg_0748;
  reg [8:0] reg_0749;
  reg [8:0] reg_0750;
  reg [8:0] reg_0751;
  reg [8:0] reg_0752;
  reg [8:0] reg_0753;
  reg [8:0] reg_0754;
  reg [8:0] reg_0755;
  reg [8:0] reg_0756;
  reg [8:0] reg_0757;
  reg [8:0] reg_0758;
  reg [8:0] reg_0759;
  reg [8:0] reg_0760;
  reg [8:0] reg_0761;
  reg [8:0] reg_0762;
  reg [8:0] reg_0763;
  reg [8:0] reg_0764;
  reg [8:0] reg_0765;
  reg [8:0] reg_0766;
  reg [8:0] reg_0767;
  reg [8:0] reg_0768;
  reg [8:0] reg_0769;
  reg [8:0] reg_0770;
  reg [8:0] reg_0771;
  reg [8:0] reg_0772;
  reg [8:0] reg_0773;
  reg [8:0] reg_0774;
  reg [8:0] reg_0775;
  reg [8:0] reg_0776;
  reg [8:0] reg_0777;
  reg [8:0] reg_0778;
  reg [8:0] reg_0779;
  reg [8:0] reg_0780;
  reg [8:0] reg_0781;
  reg [8:0] reg_0782;
  reg [8:0] reg_0783;
  reg [8:0] reg_0784;
  reg [8:0] reg_0785;
  reg [8:0] reg_0786;
  reg [8:0] reg_0787;
  reg [8:0] reg_0788;
  reg [8:0] reg_0789;
  reg [8:0] reg_0790;
  reg [8:0] reg_0791;
  reg [8:0] reg_0792;
  reg [8:0] reg_0793;
  reg [8:0] reg_0794;
  reg [8:0] reg_0795;
  reg [8:0] reg_0796;
  reg [8:0] reg_0797;
  reg [8:0] reg_0798;
  reg [8:0] reg_0799;
  reg [8:0] reg_0800;
  reg [8:0] reg_0801;
  reg [8:0] reg_0802;
  reg [8:0] reg_0803;
  reg [8:0] reg_0804;
  reg [8:0] reg_0805;
  reg [8:0] reg_0806;
  reg [8:0] reg_0807;
  reg [8:0] reg_0808;
  reg [8:0] reg_0809;
  reg [8:0] reg_0810;
  reg [8:0] reg_0811;
  reg [8:0] reg_0812;
  reg [8:0] reg_0813;
  reg [8:0] reg_0814;
  reg [8:0] reg_0815;
  reg [8:0] reg_0816;
  reg [8:0] reg_0817;
  reg [8:0] reg_0818;
  reg [8:0] reg_0819;
  reg [8:0] reg_0820;
  reg [8:0] reg_0821;
  reg [8:0] reg_0822;
  reg [8:0] reg_0823;
  reg [8:0] reg_0824;
  reg [8:0] reg_0825;
  reg [8:0] reg_0826;
  reg [8:0] reg_0827;
  reg [8:0] reg_0828;
  reg [8:0] reg_0829;
  reg [8:0] reg_0830;
  reg [8:0] reg_0831;
  reg [8:0] reg_0832;
  reg [8:0] reg_0833;
  reg [8:0] reg_0834;
  reg [8:0] reg_0835;
  reg [8:0] reg_0836;
  reg [8:0] reg_0837;
  reg [8:0] reg_0838;
  reg [8:0] reg_0839;
  reg [8:0] reg_0840;
  reg [8:0] reg_0841;
  reg [8:0] reg_0842;
  reg [8:0] reg_0843;
  reg [8:0] reg_0844;
  reg [8:0] reg_0845;
  reg [8:0] reg_0846;
  reg [8:0] reg_0847;
  reg [8:0] reg_0848;
  reg [8:0] reg_0849;
  reg [8:0] reg_0850;
  reg [8:0] reg_0851;
  reg [8:0] reg_0852;
  reg [8:0] reg_0853;
  reg [8:0] reg_0854;
  reg [8:0] reg_0855;
  reg [8:0] reg_0856;
  reg [8:0] reg_0857;
  reg [8:0] reg_0858;
  reg [8:0] reg_0859;
  reg [8:0] reg_0860;
  reg [8:0] reg_0861;
  reg [8:0] reg_0862;
  reg [8:0] reg_0863;
  reg [8:0] reg_0864;
  reg [8:0] reg_0865;
  reg [8:0] reg_0866;
  reg [8:0] reg_0867;
  reg [8:0] reg_0868;
  reg [8:0] reg_0869;
  reg [8:0] reg_0870;
  reg [8:0] reg_0871;
  reg [8:0] reg_0872;
  reg [8:0] reg_0873;
  reg [8:0] reg_0874;
  reg [8:0] reg_0875;
  reg [8:0] reg_0876;
  reg [8:0] reg_0877;
  reg [8:0] reg_0878;
  reg [8:0] reg_0879;
  reg [8:0] reg_0880;
  reg [8:0] reg_0881;
  reg [8:0] reg_0882;
  reg [8:0] reg_0883;
  reg [8:0] reg_0884;
  reg [8:0] reg_0885;
  reg [8:0] reg_0886;
  reg [8:0] reg_0887;
  reg [8:0] reg_0888;
  reg [8:0] reg_0889;
  reg [8:0] reg_0890;
  reg [8:0] reg_0891;
  reg [8:0] reg_0892;
  reg [8:0] reg_0893;
  reg [8:0] reg_0894;
  reg [8:0] reg_0895;
  reg [8:0] reg_0896;
  reg [8:0] reg_0897;
  reg [8:0] reg_0898;
  reg [8:0] reg_0899;
  reg [8:0] reg_0900;
  reg [8:0] reg_0901;
  reg [8:0] reg_0902;
  reg [8:0] reg_0903;
  reg [8:0] reg_0904;
  reg [8:0] reg_0905;
  reg [8:0] reg_0906;
  reg [8:0] reg_0907;
  reg [8:0] reg_0908;
  reg [8:0] reg_0909;
  reg [8:0] reg_0910;
  reg [8:0] reg_0911;
  reg [8:0] reg_0912;
  reg [8:0] reg_0913;
  reg [8:0] reg_0914;
  reg [8:0] reg_0915;
  reg [8:0] reg_0916;
  reg [8:0] reg_0917;
  reg [8:0] reg_0918;
  reg [8:0] reg_0919;
  reg [8:0] reg_0920;
  reg [8:0] reg_0921;
  reg [8:0] reg_0922;
  reg [8:0] reg_0923;
  reg [8:0] reg_0924;
  reg [8:0] reg_0925;
  reg [8:0] reg_0926;
  reg [8:0] reg_0927;
  reg [8:0] reg_0928;
  reg [8:0] reg_0929;
  reg [8:0] reg_0930;
  reg [8:0] reg_0931;
  reg [8:0] reg_0932;
  reg [8:0] reg_0933;
  reg [8:0] reg_0934;
  reg [8:0] reg_0935;
  reg [8:0] reg_0936;
  reg [8:0] reg_0937;
  reg [8:0] reg_0938;
  reg [8:0] reg_0939;
  reg [8:0] reg_0940;
  reg [8:0] reg_0941;
  reg [8:0] reg_0942;
  reg [8:0] reg_0943;
  reg [8:0] reg_0944;
  reg [8:0] reg_0945;
  reg [8:0] reg_0946;
  reg [8:0] reg_0947;
  reg [8:0] reg_0948;
  reg [8:0] reg_0949;
  reg [8:0] reg_0950;
  reg [8:0] reg_0951;
  reg [8:0] reg_0952;
  reg [8:0] reg_0953;
  reg [8:0] reg_0954;
  reg [8:0] reg_0955;
  reg [8:0] reg_0956;
  reg [8:0] reg_0957;
  reg [8:0] reg_0958;
  reg [8:0] reg_0959;
  reg [8:0] reg_0960;
  reg [8:0] reg_0961;
  reg [8:0] reg_0962;
  reg [8:0] reg_0963;
  reg [8:0] reg_0964;
  reg [8:0] reg_0965;
  reg [8:0] reg_0966;
  reg [8:0] reg_0967;
  reg [8:0] reg_0968;
  reg [8:0] reg_0969;
  reg [8:0] reg_0970;
  reg [8:0] reg_0971;
  reg [8:0] reg_0972;
  reg [8:0] reg_0973;
  reg [8:0] reg_0974;
  reg [8:0] reg_0975;
  reg [8:0] reg_0976;
  reg [8:0] reg_0977;
  reg [8:0] reg_0978;
  reg [8:0] reg_0979;
  reg [8:0] reg_0980;
  reg [8:0] reg_0981;
  reg [8:0] reg_0982;
  reg [8:0] reg_0983;
  reg [8:0] reg_0984;
  reg [8:0] reg_0985;
  reg [8:0] reg_0986;
  reg [8:0] reg_0987;
  reg [8:0] reg_0988;
  reg [8:0] reg_0989;
  reg [8:0] reg_0990;
  reg [8:0] reg_0991;
  reg [8:0] reg_0992;
  reg [8:0] reg_0993;
  reg [8:0] reg_0994;
  reg [8:0] reg_0995;
  reg [8:0] reg_0996;
  reg [8:0] reg_0997;
  reg [8:0] reg_0998;
  reg [8:0] reg_0999;
  reg [8:0] reg_1000;
  reg [8:0] reg_1001;
  reg [8:0] reg_1002;
  reg [8:0] reg_1003;
  reg [8:0] reg_1004;
  reg [8:0] reg_1005;
  reg [8:0] reg_1006;
  reg [8:0] reg_1007;
  reg [8:0] reg_1008;
  reg [8:0] reg_1009;
  reg [8:0] reg_1010;
  reg [8:0] reg_1011;
  reg [8:0] reg_1012;
  reg [8:0] reg_1013;
  reg [8:0] reg_1014;
  reg [8:0] reg_1015;
  reg [8:0] reg_1016;
  reg [8:0] reg_1017;
  reg [8:0] reg_1018;
  reg [8:0] reg_1019;
  reg [8:0] reg_1020;
  reg [8:0] reg_1021;
  reg [8:0] reg_1022;
  reg [8:0] reg_1023;
  reg [8:0] reg_1024;
  reg [8:0] reg_1025;
  reg [8:0] reg_1026;
  reg [8:0] reg_1027;
  reg [8:0] reg_1028;
  reg [8:0] reg_1029;
  reg [8:0] reg_1030;
  reg [8:0] reg_1031;
  reg [8:0] reg_1032;
  reg [8:0] reg_1033;
  reg [8:0] reg_1034;
  reg [8:0] reg_1035;
  reg [8:0] reg_1036;
  reg [8:0] reg_1037;
  reg [8:0] reg_1038;
  reg [8:0] reg_1039;
  reg [8:0] reg_1040;
  reg [8:0] reg_1041;
  reg [8:0] reg_1042;
  reg [8:0] reg_1043;
  reg [8:0] reg_1044;
  reg [8:0] reg_1045;
  reg [8:0] reg_1046;
  reg [8:0] reg_1047;
  reg [8:0] reg_1048;
  reg [8:0] reg_1049;
  reg [8:0] reg_1050;
  reg [8:0] reg_1051;
  reg [8:0] reg_1052;
  reg [8:0] reg_1053;
  reg [8:0] reg_1054;
  reg [8:0] reg_1055;
  reg [8:0] reg_1056;
  reg [8:0] reg_1057;

  // 制御マシンの状態
  reg [7:0] state;
  reg _busy;
  assign busy = _busy;
  // 制御マシンの動作
  always @ ( posedge clock or negedge reset ) begin
    if ( !reset ) begin
      _busy <= 0;
      state <= 0;
    end
    else if ( _busy ) begin
      if ( state < 138 ) begin
        state <= state + 1;
      end
      else begin
        _busy <= 0;
        state <= 0;
      end
    end
    else if ( start ) begin
      _busy <= 1;
    end
  end

  // 0番目の入力用メモリブロックの制御
  reg [1:0] _imem00_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem00_bank = 0;
    2: _imem00_bank = 1;
    1: _imem00_bank = 2;
    0: _imem00_bank = 3;
    4: _imem00_bank = 0;
    5: _imem00_bank = 0;
    6: _imem00_bank = 0;
    7: _imem00_bank = 0;
    8: _imem00_bank = 0;
    9: _imem00_bank = 0;
    10: _imem00_bank = 0;
    11: _imem00_bank = 0;
    12: _imem00_bank = 0;
    13: _imem00_bank = 0;
    14: _imem00_bank = 0;
    15: _imem00_bank = 0;
    16: _imem00_bank = 0;
    17: _imem00_bank = 0;
    18: _imem00_bank = 0;
    19: _imem00_bank = 0;
    20: _imem00_bank = 0;
    21: _imem00_bank = 0;
    22: _imem00_bank = 0;
    23: _imem00_bank = 0;
    24: _imem00_bank = 0;
    25: _imem00_bank = 0;
    26: _imem00_bank = 0;
    27: _imem00_bank = 0;
    28: _imem00_bank = 0;
    29: _imem00_bank = 0;
    30: _imem00_bank = 0;
    31: _imem00_bank = 0;
    32: _imem00_bank = 0;
    33: _imem00_bank = 0;
    34: _imem00_bank = 0;
    35: _imem00_bank = 0;
    36: _imem00_bank = 0;
    37: _imem00_bank = 0;
    38: _imem00_bank = 0;
    39: _imem00_bank = 0;
    40: _imem00_bank = 0;
    41: _imem00_bank = 0;
    42: _imem00_bank = 0;
    43: _imem00_bank = 0;
    44: _imem00_bank = 0;
    45: _imem00_bank = 0;
    46: _imem00_bank = 0;
    47: _imem00_bank = 0;
    48: _imem00_bank = 0;
    49: _imem00_bank = 0;
    50: _imem00_bank = 0;
    51: _imem00_bank = 0;
    52: _imem00_bank = 0;
    53: _imem00_bank = 1;
    54: _imem00_bank = 0;
    55: _imem00_bank = 0;
    56: _imem00_bank = 0;
    57: _imem00_bank = 0;
    58: _imem00_bank = 0;
    59: _imem00_bank = 0;
    60: _imem00_bank = 0;
    61: _imem00_bank = 0;
    62: _imem00_bank = 0;
    63: _imem00_bank = 0;
    64: _imem00_bank = 0;
    65: _imem00_bank = 0;
    66: _imem00_bank = 0;
    67: _imem00_bank = 0;
    68: _imem00_bank = 0;
    69: _imem00_bank = 0;
    70: _imem00_bank = 0;
    71: _imem00_bank = 0;
    72: _imem00_bank = 0;
    73: _imem00_bank = 0;
    74: _imem00_bank = 0;
    75: _imem00_bank = 0;
    76: _imem00_bank = 0;
    77: _imem00_bank = 0;
    78: _imem00_bank = 0;
    79: _imem00_bank = 0;
    80: _imem00_bank = 0;
    81: _imem00_bank = 0;
    82: _imem00_bank = 0;
    83: _imem00_bank = 0;
    84: _imem00_bank = 0;
    85: _imem00_bank = 0;
    86: _imem00_bank = 0;
    87: _imem00_bank = 0;
    88: _imem00_bank = 0;
    89: _imem00_bank = 1;
    90: _imem00_bank = 0;
    91: _imem00_bank = 0;
    92: _imem00_bank = 0;
    93: _imem00_bank = 0;
    94: _imem00_bank = 0;
    95: _imem00_bank = 0;
    default: _imem00_bank = 0;
    endcase
  end // always @ ( * )
  assign imem00_bank = _imem00_bank;
  reg _imem00_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem00_rd = 1;
    2: _imem00_rd = 1;
    1: _imem00_rd = 1;
    0: _imem00_rd = 1;
    4: _imem00_rd = 1;
    5: _imem00_rd = 1;
    6: _imem00_rd = 1;
    7: _imem00_rd = 1;
    8: _imem00_rd = 1;
    9: _imem00_rd = 1;
    10: _imem00_rd = 1;
    11: _imem00_rd = 1;
    12: _imem00_rd = 1;
    13: _imem00_rd = 1;
    14: _imem00_rd = 1;
    15: _imem00_rd = 1;
    16: _imem00_rd = 1;
    17: _imem00_rd = 1;
    18: _imem00_rd = 1;
    19: _imem00_rd = 1;
    20: _imem00_rd = 1;
    21: _imem00_rd = 1;
    22: _imem00_rd = 1;
    23: _imem00_rd = 1;
    24: _imem00_rd = 1;
    25: _imem00_rd = 1;
    26: _imem00_rd = 1;
    27: _imem00_rd = 1;
    28: _imem00_rd = 1;
    29: _imem00_rd = 1;
    30: _imem00_rd = 1;
    31: _imem00_rd = 1;
    32: _imem00_rd = 1;
    33: _imem00_rd = 1;
    34: _imem00_rd = 1;
    35: _imem00_rd = 1;
    36: _imem00_rd = 1;
    37: _imem00_rd = 1;
    38: _imem00_rd = 1;
    39: _imem00_rd = 1;
    40: _imem00_rd = 1;
    41: _imem00_rd = 1;
    42: _imem00_rd = 1;
    43: _imem00_rd = 1;
    44: _imem00_rd = 1;
    45: _imem00_rd = 1;
    46: _imem00_rd = 1;
    47: _imem00_rd = 1;
    48: _imem00_rd = 1;
    49: _imem00_rd = 1;
    50: _imem00_rd = 1;
    51: _imem00_rd = 1;
    52: _imem00_rd = 1;
    53: _imem00_rd = 1;
    54: _imem00_rd = 1;
    55: _imem00_rd = 1;
    56: _imem00_rd = 1;
    57: _imem00_rd = 1;
    58: _imem00_rd = 1;
    59: _imem00_rd = 1;
    60: _imem00_rd = 1;
    61: _imem00_rd = 1;
    62: _imem00_rd = 1;
    63: _imem00_rd = 1;
    64: _imem00_rd = 1;
    65: _imem00_rd = 1;
    66: _imem00_rd = 1;
    67: _imem00_rd = 1;
    68: _imem00_rd = 1;
    69: _imem00_rd = 1;
    70: _imem00_rd = 1;
    71: _imem00_rd = 1;
    72: _imem00_rd = 1;
    73: _imem00_rd = 1;
    74: _imem00_rd = 1;
    75: _imem00_rd = 1;
    76: _imem00_rd = 1;
    77: _imem00_rd = 1;
    78: _imem00_rd = 1;
    79: _imem00_rd = 1;
    80: _imem00_rd = 1;
    81: _imem00_rd = 1;
    82: _imem00_rd = 1;
    83: _imem00_rd = 1;
    84: _imem00_rd = 1;
    85: _imem00_rd = 1;
    86: _imem00_rd = 1;
    87: _imem00_rd = 1;
    88: _imem00_rd = 1;
    89: _imem00_rd = 1;
    90: _imem00_rd = 1;
    91: _imem00_rd = 1;
    92: _imem00_rd = 1;
    93: _imem00_rd = 1;
    94: _imem00_rd = 1;
    95: _imem00_rd = 1;
    default: _imem00_rd = 0;
    endcase
  end // always @ ( * )
  assign imem00_rd = _imem00_rd;

  // 1番目の入力用メモリブロックの制御
  reg [1:0] _imem01_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem01_bank = 0;
    2: _imem01_bank = 1;
    1: _imem01_bank = 2;
    0: _imem01_bank = 3;
    4: _imem01_bank = 0;
    5: _imem01_bank = 0;
    6: _imem01_bank = 0;
    7: _imem01_bank = 0;
    8: _imem01_bank = 2;
    9: _imem01_bank = 1;
    10: _imem01_bank = 0;
    11: _imem01_bank = 0;
    12: _imem01_bank = 0;
    13: _imem01_bank = 0;
    14: _imem01_bank = 0;
    15: _imem01_bank = 0;
    16: _imem01_bank = 0;
    17: _imem01_bank = 0;
    18: _imem01_bank = 0;
    19: _imem01_bank = 0;
    20: _imem01_bank = 0;
    21: _imem01_bank = 0;
    22: _imem01_bank = 0;
    23: _imem01_bank = 1;
    24: _imem01_bank = 0;
    25: _imem01_bank = 0;
    26: _imem01_bank = 0;
    27: _imem01_bank = 0;
    28: _imem01_bank = 0;
    29: _imem01_bank = 0;
    30: _imem01_bank = 0;
    31: _imem01_bank = 0;
    32: _imem01_bank = 0;
    33: _imem01_bank = 0;
    34: _imem01_bank = 0;
    35: _imem01_bank = 0;
    36: _imem01_bank = 0;
    37: _imem01_bank = 0;
    38: _imem01_bank = 2;
    39: _imem01_bank = 2;
    40: _imem01_bank = 0;
    41: _imem01_bank = 0;
    42: _imem01_bank = 0;
    43: _imem01_bank = 0;
    44: _imem01_bank = 0;
    45: _imem01_bank = 0;
    46: _imem01_bank = 1;
    47: _imem01_bank = 1;
    48: _imem01_bank = 0;
    49: _imem01_bank = 0;
    50: _imem01_bank = 0;
    51: _imem01_bank = 3;
    52: _imem01_bank = 0;
    53: _imem01_bank = 0;
    54: _imem01_bank = 0;
    55: _imem01_bank = 0;
    56: _imem01_bank = 0;
    57: _imem01_bank = 0;
    58: _imem01_bank = 0;
    59: _imem01_bank = 0;
    60: _imem01_bank = 0;
    61: _imem01_bank = 0;
    62: _imem01_bank = 0;
    63: _imem01_bank = 0;
    64: _imem01_bank = 0;
    65: _imem01_bank = 0;
    66: _imem01_bank = 0;
    67: _imem01_bank = 1;
    68: _imem01_bank = 0;
    69: _imem01_bank = 0;
    70: _imem01_bank = 0;
    71: _imem01_bank = 0;
    72: _imem01_bank = 0;
    73: _imem01_bank = 0;
    74: _imem01_bank = 0;
    75: _imem01_bank = 0;
    76: _imem01_bank = 0;
    77: _imem01_bank = 0;
    78: _imem01_bank = 0;
    79: _imem01_bank = 0;
    80: _imem01_bank = 0;
    81: _imem01_bank = 0;
    82: _imem01_bank = 0;
    83: _imem01_bank = 0;
    84: _imem01_bank = 0;
    85: _imem01_bank = 0;
    86: _imem01_bank = 0;
    87: _imem01_bank = 0;
    88: _imem01_bank = 0;
    89: _imem01_bank = 0;
    90: _imem01_bank = 0;
    91: _imem01_bank = 2;
    92: _imem01_bank = 1;
    93: _imem01_bank = 2;
    94: _imem01_bank = 1;
    95: _imem01_bank = 0;
    default: _imem01_bank = 0;
    endcase
  end // always @ ( * )
  assign imem01_bank = _imem01_bank;
  reg _imem01_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem01_rd = 1;
    2: _imem01_rd = 1;
    1: _imem01_rd = 1;
    0: _imem01_rd = 1;
    4: _imem01_rd = 1;
    5: _imem01_rd = 1;
    6: _imem01_rd = 1;
    7: _imem01_rd = 1;
    8: _imem01_rd = 1;
    9: _imem01_rd = 1;
    10: _imem01_rd = 1;
    11: _imem01_rd = 1;
    12: _imem01_rd = 1;
    13: _imem01_rd = 1;
    14: _imem01_rd = 1;
    15: _imem01_rd = 1;
    16: _imem01_rd = 1;
    17: _imem01_rd = 1;
    18: _imem01_rd = 1;
    19: _imem01_rd = 1;
    20: _imem01_rd = 1;
    21: _imem01_rd = 1;
    22: _imem01_rd = 1;
    23: _imem01_rd = 1;
    24: _imem01_rd = 1;
    25: _imem01_rd = 1;
    26: _imem01_rd = 1;
    27: _imem01_rd = 1;
    28: _imem01_rd = 1;
    29: _imem01_rd = 1;
    30: _imem01_rd = 1;
    31: _imem01_rd = 1;
    32: _imem01_rd = 1;
    33: _imem01_rd = 1;
    34: _imem01_rd = 1;
    35: _imem01_rd = 1;
    36: _imem01_rd = 1;
    37: _imem01_rd = 1;
    38: _imem01_rd = 1;
    39: _imem01_rd = 1;
    40: _imem01_rd = 1;
    41: _imem01_rd = 1;
    42: _imem01_rd = 1;
    43: _imem01_rd = 1;
    44: _imem01_rd = 1;
    45: _imem01_rd = 1;
    46: _imem01_rd = 1;
    47: _imem01_rd = 1;
    48: _imem01_rd = 1;
    49: _imem01_rd = 1;
    50: _imem01_rd = 1;
    51: _imem01_rd = 1;
    52: _imem01_rd = 1;
    53: _imem01_rd = 1;
    54: _imem01_rd = 1;
    55: _imem01_rd = 1;
    56: _imem01_rd = 1;
    57: _imem01_rd = 1;
    58: _imem01_rd = 1;
    59: _imem01_rd = 1;
    60: _imem01_rd = 1;
    61: _imem01_rd = 1;
    62: _imem01_rd = 1;
    63: _imem01_rd = 1;
    64: _imem01_rd = 1;
    65: _imem01_rd = 1;
    66: _imem01_rd = 1;
    67: _imem01_rd = 1;
    68: _imem01_rd = 1;
    69: _imem01_rd = 1;
    70: _imem01_rd = 1;
    71: _imem01_rd = 1;
    72: _imem01_rd = 1;
    73: _imem01_rd = 1;
    74: _imem01_rd = 1;
    75: _imem01_rd = 1;
    76: _imem01_rd = 1;
    77: _imem01_rd = 1;
    78: _imem01_rd = 1;
    79: _imem01_rd = 1;
    80: _imem01_rd = 1;
    81: _imem01_rd = 1;
    82: _imem01_rd = 1;
    83: _imem01_rd = 1;
    84: _imem01_rd = 1;
    85: _imem01_rd = 1;
    86: _imem01_rd = 1;
    87: _imem01_rd = 1;
    88: _imem01_rd = 1;
    89: _imem01_rd = 1;
    90: _imem01_rd = 1;
    91: _imem01_rd = 1;
    92: _imem01_rd = 1;
    93: _imem01_rd = 1;
    94: _imem01_rd = 1;
    95: _imem01_rd = 1;
    default: _imem01_rd = 0;
    endcase
  end // always @ ( * )
  assign imem01_rd = _imem01_rd;

  // 2番目の入力用メモリブロックの制御
  reg [1:0] _imem02_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem02_bank = 0;
    2: _imem02_bank = 1;
    1: _imem02_bank = 2;
    0: _imem02_bank = 3;
    4: _imem02_bank = 0;
    5: _imem02_bank = 0;
    6: _imem02_bank = 0;
    7: _imem02_bank = 0;
    8: _imem02_bank = 0;
    9: _imem02_bank = 0;
    10: _imem02_bank = 0;
    11: _imem02_bank = 0;
    12: _imem02_bank = 0;
    13: _imem02_bank = 0;
    14: _imem02_bank = 0;
    15: _imem02_bank = 0;
    16: _imem02_bank = 0;
    17: _imem02_bank = 0;
    18: _imem02_bank = 0;
    19: _imem02_bank = 3;
    20: _imem02_bank = 0;
    21: _imem02_bank = 0;
    22: _imem02_bank = 0;
    23: _imem02_bank = 0;
    24: _imem02_bank = 2;
    25: _imem02_bank = 0;
    26: _imem02_bank = 0;
    27: _imem02_bank = 0;
    28: _imem02_bank = 0;
    29: _imem02_bank = 0;
    30: _imem02_bank = 0;
    31: _imem02_bank = 0;
    32: _imem02_bank = 0;
    33: _imem02_bank = 0;
    34: _imem02_bank = 0;
    35: _imem02_bank = 0;
    36: _imem02_bank = 0;
    37: _imem02_bank = 0;
    38: _imem02_bank = 0;
    39: _imem02_bank = 0;
    40: _imem02_bank = 0;
    41: _imem02_bank = 0;
    42: _imem02_bank = 0;
    43: _imem02_bank = 1;
    44: _imem02_bank = 0;
    45: _imem02_bank = 0;
    46: _imem02_bank = 0;
    47: _imem02_bank = 0;
    48: _imem02_bank = 0;
    49: _imem02_bank = 0;
    50: _imem02_bank = 2;
    51: _imem02_bank = 0;
    52: _imem02_bank = 0;
    53: _imem02_bank = 0;
    54: _imem02_bank = 0;
    55: _imem02_bank = 0;
    56: _imem02_bank = 0;
    57: _imem02_bank = 0;
    58: _imem02_bank = 0;
    59: _imem02_bank = 0;
    60: _imem02_bank = 0;
    61: _imem02_bank = 1;
    62: _imem02_bank = 0;
    63: _imem02_bank = 0;
    64: _imem02_bank = 0;
    65: _imem02_bank = 0;
    66: _imem02_bank = 0;
    67: _imem02_bank = 0;
    68: _imem02_bank = 0;
    69: _imem02_bank = 0;
    70: _imem02_bank = 1;
    71: _imem02_bank = 0;
    72: _imem02_bank = 0;
    73: _imem02_bank = 0;
    74: _imem02_bank = 0;
    75: _imem02_bank = 0;
    76: _imem02_bank = 0;
    77: _imem02_bank = 0;
    78: _imem02_bank = 0;
    79: _imem02_bank = 0;
    80: _imem02_bank = 0;
    81: _imem02_bank = 0;
    82: _imem02_bank = 1;
    83: _imem02_bank = 3;
    84: _imem02_bank = 0;
    85: _imem02_bank = 0;
    86: _imem02_bank = 0;
    87: _imem02_bank = 0;
    88: _imem02_bank = 0;
    89: _imem02_bank = 0;
    90: _imem02_bank = 0;
    91: _imem02_bank = 0;
    92: _imem02_bank = 0;
    93: _imem02_bank = 0;
    94: _imem02_bank = 0;
    95: _imem02_bank = 0;
    default: _imem02_bank = 0;
    endcase
  end // always @ ( * )
  assign imem02_bank = _imem02_bank;
  reg _imem02_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem02_rd = 1;
    2: _imem02_rd = 1;
    1: _imem02_rd = 1;
    0: _imem02_rd = 1;
    4: _imem02_rd = 1;
    5: _imem02_rd = 1;
    6: _imem02_rd = 1;
    7: _imem02_rd = 1;
    8: _imem02_rd = 1;
    9: _imem02_rd = 1;
    10: _imem02_rd = 1;
    11: _imem02_rd = 1;
    12: _imem02_rd = 1;
    13: _imem02_rd = 1;
    14: _imem02_rd = 1;
    15: _imem02_rd = 1;
    16: _imem02_rd = 1;
    17: _imem02_rd = 1;
    18: _imem02_rd = 1;
    19: _imem02_rd = 1;
    20: _imem02_rd = 1;
    21: _imem02_rd = 1;
    22: _imem02_rd = 1;
    23: _imem02_rd = 1;
    24: _imem02_rd = 1;
    25: _imem02_rd = 1;
    26: _imem02_rd = 1;
    27: _imem02_rd = 1;
    28: _imem02_rd = 1;
    29: _imem02_rd = 1;
    30: _imem02_rd = 1;
    31: _imem02_rd = 1;
    32: _imem02_rd = 1;
    33: _imem02_rd = 1;
    34: _imem02_rd = 1;
    35: _imem02_rd = 1;
    36: _imem02_rd = 1;
    37: _imem02_rd = 1;
    38: _imem02_rd = 1;
    39: _imem02_rd = 1;
    40: _imem02_rd = 1;
    41: _imem02_rd = 1;
    42: _imem02_rd = 1;
    43: _imem02_rd = 1;
    44: _imem02_rd = 1;
    45: _imem02_rd = 1;
    46: _imem02_rd = 1;
    47: _imem02_rd = 1;
    48: _imem02_rd = 1;
    49: _imem02_rd = 1;
    50: _imem02_rd = 1;
    51: _imem02_rd = 1;
    52: _imem02_rd = 1;
    53: _imem02_rd = 1;
    54: _imem02_rd = 1;
    55: _imem02_rd = 1;
    56: _imem02_rd = 1;
    57: _imem02_rd = 1;
    58: _imem02_rd = 1;
    59: _imem02_rd = 1;
    60: _imem02_rd = 1;
    61: _imem02_rd = 1;
    62: _imem02_rd = 1;
    63: _imem02_rd = 1;
    64: _imem02_rd = 1;
    65: _imem02_rd = 1;
    66: _imem02_rd = 1;
    67: _imem02_rd = 1;
    68: _imem02_rd = 1;
    69: _imem02_rd = 1;
    70: _imem02_rd = 1;
    71: _imem02_rd = 1;
    72: _imem02_rd = 1;
    73: _imem02_rd = 1;
    74: _imem02_rd = 1;
    75: _imem02_rd = 1;
    76: _imem02_rd = 1;
    77: _imem02_rd = 1;
    78: _imem02_rd = 1;
    79: _imem02_rd = 1;
    80: _imem02_rd = 1;
    81: _imem02_rd = 1;
    82: _imem02_rd = 1;
    83: _imem02_rd = 1;
    84: _imem02_rd = 1;
    85: _imem02_rd = 1;
    86: _imem02_rd = 1;
    87: _imem02_rd = 1;
    88: _imem02_rd = 1;
    89: _imem02_rd = 1;
    90: _imem02_rd = 1;
    91: _imem02_rd = 1;
    92: _imem02_rd = 1;
    93: _imem02_rd = 1;
    94: _imem02_rd = 1;
    95: _imem02_rd = 1;
    default: _imem02_rd = 0;
    endcase
  end // always @ ( * )
  assign imem02_rd = _imem02_rd;

  // 3番目の入力用メモリブロックの制御
  reg [1:0] _imem03_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem03_bank = 0;
    2: _imem03_bank = 1;
    1: _imem03_bank = 2;
    0: _imem03_bank = 3;
    4: _imem03_bank = 3;
    5: _imem03_bank = 0;
    6: _imem03_bank = 0;
    7: _imem03_bank = 0;
    8: _imem03_bank = 0;
    9: _imem03_bank = 0;
    10: _imem03_bank = 0;
    11: _imem03_bank = 0;
    12: _imem03_bank = 0;
    13: _imem03_bank = 0;
    14: _imem03_bank = 0;
    15: _imem03_bank = 0;
    16: _imem03_bank = 0;
    17: _imem03_bank = 0;
    18: _imem03_bank = 0;
    19: _imem03_bank = 0;
    20: _imem03_bank = 0;
    21: _imem03_bank = 0;
    22: _imem03_bank = 0;
    23: _imem03_bank = 0;
    24: _imem03_bank = 0;
    25: _imem03_bank = 0;
    26: _imem03_bank = 2;
    27: _imem03_bank = 0;
    28: _imem03_bank = 0;
    29: _imem03_bank = 1;
    30: _imem03_bank = 0;
    31: _imem03_bank = 0;
    32: _imem03_bank = 0;
    33: _imem03_bank = 0;
    34: _imem03_bank = 0;
    35: _imem03_bank = 0;
    36: _imem03_bank = 0;
    37: _imem03_bank = 0;
    38: _imem03_bank = 0;
    39: _imem03_bank = 0;
    40: _imem03_bank = 0;
    41: _imem03_bank = 0;
    42: _imem03_bank = 0;
    43: _imem03_bank = 0;
    44: _imem03_bank = 0;
    45: _imem03_bank = 0;
    46: _imem03_bank = 0;
    47: _imem03_bank = 0;
    48: _imem03_bank = 0;
    49: _imem03_bank = 0;
    50: _imem03_bank = 0;
    51: _imem03_bank = 0;
    52: _imem03_bank = 1;
    53: _imem03_bank = 1;
    54: _imem03_bank = 0;
    55: _imem03_bank = 0;
    56: _imem03_bank = 0;
    57: _imem03_bank = 0;
    58: _imem03_bank = 0;
    59: _imem03_bank = 0;
    60: _imem03_bank = 0;
    61: _imem03_bank = 0;
    62: _imem03_bank = 0;
    63: _imem03_bank = 0;
    64: _imem03_bank = 0;
    65: _imem03_bank = 0;
    66: _imem03_bank = 0;
    67: _imem03_bank = 0;
    68: _imem03_bank = 2;
    69: _imem03_bank = 0;
    70: _imem03_bank = 0;
    71: _imem03_bank = 0;
    72: _imem03_bank = 0;
    73: _imem03_bank = 0;
    74: _imem03_bank = 0;
    75: _imem03_bank = 0;
    76: _imem03_bank = 0;
    77: _imem03_bank = 0;
    78: _imem03_bank = 0;
    79: _imem03_bank = 0;
    80: _imem03_bank = 0;
    81: _imem03_bank = 0;
    82: _imem03_bank = 0;
    83: _imem03_bank = 0;
    84: _imem03_bank = 0;
    85: _imem03_bank = 0;
    86: _imem03_bank = 1;
    87: _imem03_bank = 0;
    88: _imem03_bank = 3;
    89: _imem03_bank = 0;
    90: _imem03_bank = 0;
    91: _imem03_bank = 0;
    92: _imem03_bank = 0;
    93: _imem03_bank = 0;
    94: _imem03_bank = 0;
    95: _imem03_bank = 0;
    default: _imem03_bank = 0;
    endcase
  end // always @ ( * )
  assign imem03_bank = _imem03_bank;
  reg _imem03_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem03_rd = 1;
    2: _imem03_rd = 1;
    1: _imem03_rd = 1;
    0: _imem03_rd = 1;
    4: _imem03_rd = 1;
    5: _imem03_rd = 1;
    6: _imem03_rd = 1;
    7: _imem03_rd = 1;
    8: _imem03_rd = 1;
    9: _imem03_rd = 1;
    10: _imem03_rd = 1;
    11: _imem03_rd = 1;
    12: _imem03_rd = 1;
    13: _imem03_rd = 1;
    14: _imem03_rd = 1;
    15: _imem03_rd = 1;
    16: _imem03_rd = 1;
    17: _imem03_rd = 1;
    18: _imem03_rd = 1;
    19: _imem03_rd = 1;
    20: _imem03_rd = 1;
    21: _imem03_rd = 1;
    22: _imem03_rd = 1;
    23: _imem03_rd = 1;
    24: _imem03_rd = 1;
    25: _imem03_rd = 1;
    26: _imem03_rd = 1;
    27: _imem03_rd = 1;
    28: _imem03_rd = 1;
    29: _imem03_rd = 1;
    30: _imem03_rd = 1;
    31: _imem03_rd = 1;
    32: _imem03_rd = 1;
    33: _imem03_rd = 1;
    34: _imem03_rd = 1;
    35: _imem03_rd = 1;
    36: _imem03_rd = 1;
    37: _imem03_rd = 1;
    38: _imem03_rd = 1;
    39: _imem03_rd = 1;
    40: _imem03_rd = 1;
    41: _imem03_rd = 1;
    42: _imem03_rd = 1;
    43: _imem03_rd = 1;
    44: _imem03_rd = 1;
    45: _imem03_rd = 1;
    46: _imem03_rd = 1;
    47: _imem03_rd = 1;
    48: _imem03_rd = 1;
    49: _imem03_rd = 1;
    50: _imem03_rd = 1;
    51: _imem03_rd = 1;
    52: _imem03_rd = 1;
    53: _imem03_rd = 1;
    54: _imem03_rd = 1;
    55: _imem03_rd = 1;
    56: _imem03_rd = 1;
    57: _imem03_rd = 1;
    58: _imem03_rd = 1;
    59: _imem03_rd = 1;
    60: _imem03_rd = 1;
    61: _imem03_rd = 1;
    62: _imem03_rd = 1;
    63: _imem03_rd = 1;
    64: _imem03_rd = 1;
    65: _imem03_rd = 1;
    66: _imem03_rd = 1;
    67: _imem03_rd = 1;
    68: _imem03_rd = 1;
    69: _imem03_rd = 1;
    70: _imem03_rd = 1;
    71: _imem03_rd = 1;
    72: _imem03_rd = 1;
    73: _imem03_rd = 1;
    74: _imem03_rd = 1;
    75: _imem03_rd = 1;
    76: _imem03_rd = 1;
    77: _imem03_rd = 1;
    78: _imem03_rd = 1;
    79: _imem03_rd = 1;
    80: _imem03_rd = 1;
    81: _imem03_rd = 1;
    82: _imem03_rd = 1;
    83: _imem03_rd = 1;
    84: _imem03_rd = 1;
    85: _imem03_rd = 1;
    86: _imem03_rd = 1;
    87: _imem03_rd = 1;
    88: _imem03_rd = 1;
    89: _imem03_rd = 1;
    90: _imem03_rd = 1;
    91: _imem03_rd = 1;
    92: _imem03_rd = 1;
    93: _imem03_rd = 1;
    94: _imem03_rd = 1;
    95: _imem03_rd = 1;
    default: _imem03_rd = 0;
    endcase
  end // always @ ( * )
  assign imem03_rd = _imem03_rd;

  // 4番目の入力用メモリブロックの制御
  reg [1:0] _imem04_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem04_bank = 0;
    2: _imem04_bank = 1;
    1: _imem04_bank = 2;
    0: _imem04_bank = 3;
    4: _imem04_bank = 0;
    5: _imem04_bank = 0;
    6: _imem04_bank = 0;
    7: _imem04_bank = 0;
    8: _imem04_bank = 0;
    9: _imem04_bank = 0;
    10: _imem04_bank = 0;
    11: _imem04_bank = 0;
    12: _imem04_bank = 0;
    13: _imem04_bank = 0;
    14: _imem04_bank = 0;
    15: _imem04_bank = 0;
    16: _imem04_bank = 3;
    17: _imem04_bank = 2;
    18: _imem04_bank = 0;
    19: _imem04_bank = 0;
    20: _imem04_bank = 1;
    21: _imem04_bank = 0;
    22: _imem04_bank = 1;
    23: _imem04_bank = 0;
    24: _imem04_bank = 0;
    25: _imem04_bank = 0;
    26: _imem04_bank = 0;
    27: _imem04_bank = 0;
    28: _imem04_bank = 0;
    29: _imem04_bank = 0;
    30: _imem04_bank = 0;
    31: _imem04_bank = 0;
    32: _imem04_bank = 0;
    33: _imem04_bank = 0;
    34: _imem04_bank = 0;
    35: _imem04_bank = 0;
    36: _imem04_bank = 0;
    37: _imem04_bank = 0;
    38: _imem04_bank = 0;
    39: _imem04_bank = 0;
    40: _imem04_bank = 2;
    41: _imem04_bank = 0;
    42: _imem04_bank = 0;
    43: _imem04_bank = 0;
    44: _imem04_bank = 3;
    45: _imem04_bank = 0;
    46: _imem04_bank = 0;
    47: _imem04_bank = 3;
    48: _imem04_bank = 0;
    49: _imem04_bank = 0;
    50: _imem04_bank = 0;
    51: _imem04_bank = 0;
    52: _imem04_bank = 0;
    53: _imem04_bank = 0;
    54: _imem04_bank = 0;
    55: _imem04_bank = 0;
    56: _imem04_bank = 0;
    57: _imem04_bank = 3;
    58: _imem04_bank = 0;
    59: _imem04_bank = 0;
    60: _imem04_bank = 0;
    61: _imem04_bank = 0;
    62: _imem04_bank = 0;
    63: _imem04_bank = 0;
    64: _imem04_bank = 0;
    65: _imem04_bank = 0;
    66: _imem04_bank = 0;
    67: _imem04_bank = 0;
    68: _imem04_bank = 0;
    69: _imem04_bank = 0;
    70: _imem04_bank = 0;
    71: _imem04_bank = 0;
    72: _imem04_bank = 0;
    73: _imem04_bank = 0;
    74: _imem04_bank = 0;
    75: _imem04_bank = 0;
    76: _imem04_bank = 0;
    77: _imem04_bank = 0;
    78: _imem04_bank = 0;
    79: _imem04_bank = 0;
    80: _imem04_bank = 0;
    81: _imem04_bank = 1;
    82: _imem04_bank = 0;
    83: _imem04_bank = 0;
    84: _imem04_bank = 0;
    85: _imem04_bank = 0;
    86: _imem04_bank = 0;
    87: _imem04_bank = 0;
    88: _imem04_bank = 0;
    89: _imem04_bank = 0;
    90: _imem04_bank = 0;
    91: _imem04_bank = 0;
    92: _imem04_bank = 0;
    93: _imem04_bank = 0;
    94: _imem04_bank = 0;
    95: _imem04_bank = 0;
    default: _imem04_bank = 0;
    endcase
  end // always @ ( * )
  assign imem04_bank = _imem04_bank;
  reg _imem04_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem04_rd = 1;
    2: _imem04_rd = 1;
    1: _imem04_rd = 1;
    0: _imem04_rd = 1;
    4: _imem04_rd = 1;
    5: _imem04_rd = 1;
    6: _imem04_rd = 1;
    7: _imem04_rd = 1;
    8: _imem04_rd = 1;
    9: _imem04_rd = 1;
    10: _imem04_rd = 1;
    11: _imem04_rd = 1;
    12: _imem04_rd = 1;
    13: _imem04_rd = 1;
    14: _imem04_rd = 1;
    15: _imem04_rd = 1;
    16: _imem04_rd = 1;
    17: _imem04_rd = 1;
    18: _imem04_rd = 1;
    19: _imem04_rd = 1;
    20: _imem04_rd = 1;
    21: _imem04_rd = 1;
    22: _imem04_rd = 1;
    23: _imem04_rd = 1;
    24: _imem04_rd = 1;
    25: _imem04_rd = 1;
    26: _imem04_rd = 1;
    27: _imem04_rd = 1;
    28: _imem04_rd = 1;
    29: _imem04_rd = 1;
    30: _imem04_rd = 1;
    31: _imem04_rd = 1;
    32: _imem04_rd = 1;
    33: _imem04_rd = 1;
    34: _imem04_rd = 1;
    35: _imem04_rd = 1;
    36: _imem04_rd = 1;
    37: _imem04_rd = 1;
    38: _imem04_rd = 1;
    39: _imem04_rd = 1;
    40: _imem04_rd = 1;
    41: _imem04_rd = 1;
    42: _imem04_rd = 1;
    43: _imem04_rd = 1;
    44: _imem04_rd = 1;
    45: _imem04_rd = 1;
    46: _imem04_rd = 1;
    47: _imem04_rd = 1;
    48: _imem04_rd = 1;
    49: _imem04_rd = 1;
    50: _imem04_rd = 1;
    51: _imem04_rd = 1;
    52: _imem04_rd = 1;
    53: _imem04_rd = 1;
    54: _imem04_rd = 1;
    55: _imem04_rd = 1;
    56: _imem04_rd = 1;
    57: _imem04_rd = 1;
    58: _imem04_rd = 1;
    59: _imem04_rd = 1;
    60: _imem04_rd = 1;
    61: _imem04_rd = 1;
    62: _imem04_rd = 1;
    63: _imem04_rd = 1;
    64: _imem04_rd = 1;
    65: _imem04_rd = 1;
    66: _imem04_rd = 1;
    67: _imem04_rd = 1;
    68: _imem04_rd = 1;
    69: _imem04_rd = 1;
    70: _imem04_rd = 1;
    71: _imem04_rd = 1;
    72: _imem04_rd = 1;
    73: _imem04_rd = 1;
    74: _imem04_rd = 1;
    75: _imem04_rd = 1;
    76: _imem04_rd = 1;
    77: _imem04_rd = 1;
    78: _imem04_rd = 1;
    79: _imem04_rd = 1;
    80: _imem04_rd = 1;
    81: _imem04_rd = 1;
    82: _imem04_rd = 1;
    83: _imem04_rd = 1;
    84: _imem04_rd = 1;
    85: _imem04_rd = 1;
    86: _imem04_rd = 1;
    87: _imem04_rd = 1;
    88: _imem04_rd = 1;
    89: _imem04_rd = 1;
    90: _imem04_rd = 1;
    91: _imem04_rd = 1;
    92: _imem04_rd = 1;
    93: _imem04_rd = 1;
    94: _imem04_rd = 1;
    95: _imem04_rd = 1;
    default: _imem04_rd = 0;
    endcase
  end // always @ ( * )
  assign imem04_rd = _imem04_rd;

  // 5番目の入力用メモリブロックの制御
  reg [1:0] _imem05_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem05_bank = 0;
    2: _imem05_bank = 1;
    1: _imem05_bank = 2;
    0: _imem05_bank = 3;
    4: _imem05_bank = 1;
    5: _imem05_bank = 0;
    6: _imem05_bank = 0;
    7: _imem05_bank = 0;
    8: _imem05_bank = 0;
    9: _imem05_bank = 0;
    10: _imem05_bank = 2;
    11: _imem05_bank = 0;
    12: _imem05_bank = 0;
    13: _imem05_bank = 0;
    14: _imem05_bank = 0;
    15: _imem05_bank = 0;
    16: _imem05_bank = 0;
    17: _imem05_bank = 0;
    18: _imem05_bank = 2;
    19: _imem05_bank = 0;
    20: _imem05_bank = 0;
    21: _imem05_bank = 0;
    22: _imem05_bank = 0;
    23: _imem05_bank = 0;
    24: _imem05_bank = 0;
    25: _imem05_bank = 0;
    26: _imem05_bank = 0;
    27: _imem05_bank = 0;
    28: _imem05_bank = 0;
    29: _imem05_bank = 0;
    30: _imem05_bank = 0;
    31: _imem05_bank = 0;
    32: _imem05_bank = 0;
    33: _imem05_bank = 0;
    34: _imem05_bank = 0;
    35: _imem05_bank = 0;
    36: _imem05_bank = 0;
    37: _imem05_bank = 0;
    38: _imem05_bank = 0;
    39: _imem05_bank = 0;
    40: _imem05_bank = 0;
    41: _imem05_bank = 0;
    42: _imem05_bank = 0;
    43: _imem05_bank = 0;
    44: _imem05_bank = 0;
    45: _imem05_bank = 0;
    46: _imem05_bank = 0;
    47: _imem05_bank = 0;
    48: _imem05_bank = 2;
    49: _imem05_bank = 0;
    50: _imem05_bank = 0;
    51: _imem05_bank = 0;
    52: _imem05_bank = 0;
    53: _imem05_bank = 0;
    54: _imem05_bank = 1;
    55: _imem05_bank = 0;
    56: _imem05_bank = 0;
    57: _imem05_bank = 0;
    58: _imem05_bank = 0;
    59: _imem05_bank = 1;
    60: _imem05_bank = 0;
    61: _imem05_bank = 0;
    62: _imem05_bank = 0;
    63: _imem05_bank = 1;
    64: _imem05_bank = 2;
    65: _imem05_bank = 0;
    66: _imem05_bank = 1;
    67: _imem05_bank = 0;
    68: _imem05_bank = 0;
    69: _imem05_bank = 0;
    70: _imem05_bank = 0;
    71: _imem05_bank = 1;
    72: _imem05_bank = 3;
    73: _imem05_bank = 0;
    74: _imem05_bank = 0;
    75: _imem05_bank = 0;
    76: _imem05_bank = 0;
    77: _imem05_bank = 2;
    78: _imem05_bank = 0;
    79: _imem05_bank = 0;
    80: _imem05_bank = 0;
    81: _imem05_bank = 0;
    82: _imem05_bank = 0;
    83: _imem05_bank = 0;
    84: _imem05_bank = 0;
    85: _imem05_bank = 2;
    86: _imem05_bank = 0;
    87: _imem05_bank = 0;
    88: _imem05_bank = 0;
    89: _imem05_bank = 0;
    90: _imem05_bank = 0;
    91: _imem05_bank = 0;
    92: _imem05_bank = 0;
    93: _imem05_bank = 0;
    94: _imem05_bank = 0;
    95: _imem05_bank = 0;
    default: _imem05_bank = 0;
    endcase
  end // always @ ( * )
  assign imem05_bank = _imem05_bank;
  reg _imem05_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem05_rd = 1;
    2: _imem05_rd = 1;
    1: _imem05_rd = 1;
    0: _imem05_rd = 1;
    4: _imem05_rd = 1;
    5: _imem05_rd = 1;
    6: _imem05_rd = 1;
    7: _imem05_rd = 1;
    8: _imem05_rd = 1;
    9: _imem05_rd = 1;
    10: _imem05_rd = 1;
    11: _imem05_rd = 1;
    12: _imem05_rd = 1;
    13: _imem05_rd = 1;
    14: _imem05_rd = 1;
    15: _imem05_rd = 1;
    16: _imem05_rd = 1;
    17: _imem05_rd = 1;
    18: _imem05_rd = 1;
    19: _imem05_rd = 1;
    20: _imem05_rd = 1;
    21: _imem05_rd = 1;
    22: _imem05_rd = 1;
    23: _imem05_rd = 1;
    24: _imem05_rd = 1;
    25: _imem05_rd = 1;
    26: _imem05_rd = 1;
    27: _imem05_rd = 1;
    28: _imem05_rd = 1;
    29: _imem05_rd = 1;
    30: _imem05_rd = 1;
    31: _imem05_rd = 1;
    32: _imem05_rd = 1;
    33: _imem05_rd = 1;
    34: _imem05_rd = 1;
    35: _imem05_rd = 1;
    36: _imem05_rd = 1;
    37: _imem05_rd = 1;
    38: _imem05_rd = 1;
    39: _imem05_rd = 1;
    40: _imem05_rd = 1;
    41: _imem05_rd = 1;
    42: _imem05_rd = 1;
    43: _imem05_rd = 1;
    44: _imem05_rd = 1;
    45: _imem05_rd = 1;
    46: _imem05_rd = 1;
    47: _imem05_rd = 1;
    48: _imem05_rd = 1;
    49: _imem05_rd = 1;
    50: _imem05_rd = 1;
    51: _imem05_rd = 1;
    52: _imem05_rd = 1;
    53: _imem05_rd = 1;
    54: _imem05_rd = 1;
    55: _imem05_rd = 1;
    56: _imem05_rd = 1;
    57: _imem05_rd = 1;
    58: _imem05_rd = 1;
    59: _imem05_rd = 1;
    60: _imem05_rd = 1;
    61: _imem05_rd = 1;
    62: _imem05_rd = 1;
    63: _imem05_rd = 1;
    64: _imem05_rd = 1;
    65: _imem05_rd = 1;
    66: _imem05_rd = 1;
    67: _imem05_rd = 1;
    68: _imem05_rd = 1;
    69: _imem05_rd = 1;
    70: _imem05_rd = 1;
    71: _imem05_rd = 1;
    72: _imem05_rd = 1;
    73: _imem05_rd = 1;
    74: _imem05_rd = 1;
    75: _imem05_rd = 1;
    76: _imem05_rd = 1;
    77: _imem05_rd = 1;
    78: _imem05_rd = 1;
    79: _imem05_rd = 1;
    80: _imem05_rd = 1;
    81: _imem05_rd = 1;
    82: _imem05_rd = 1;
    83: _imem05_rd = 1;
    84: _imem05_rd = 1;
    85: _imem05_rd = 1;
    86: _imem05_rd = 1;
    87: _imem05_rd = 1;
    88: _imem05_rd = 1;
    89: _imem05_rd = 1;
    90: _imem05_rd = 1;
    91: _imem05_rd = 1;
    92: _imem05_rd = 1;
    93: _imem05_rd = 1;
    94: _imem05_rd = 1;
    95: _imem05_rd = 1;
    default: _imem05_rd = 0;
    endcase
  end // always @ ( * )
  assign imem05_rd = _imem05_rd;

  // 6番目の入力用メモリブロックの制御
  reg [1:0] _imem06_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem06_bank = 0;
    2: _imem06_bank = 1;
    1: _imem06_bank = 2;
    0: _imem06_bank = 3;
    4: _imem06_bank = 0;
    5: _imem06_bank = 0;
    6: _imem06_bank = 0;
    7: _imem06_bank = 3;
    8: _imem06_bank = 0;
    9: _imem06_bank = 0;
    10: _imem06_bank = 0;
    11: _imem06_bank = 0;
    12: _imem06_bank = 0;
    13: _imem06_bank = 0;
    14: _imem06_bank = 0;
    15: _imem06_bank = 0;
    16: _imem06_bank = 0;
    17: _imem06_bank = 0;
    18: _imem06_bank = 0;
    19: _imem06_bank = 0;
    20: _imem06_bank = 0;
    21: _imem06_bank = 0;
    22: _imem06_bank = 0;
    23: _imem06_bank = 0;
    24: _imem06_bank = 0;
    25: _imem06_bank = 0;
    26: _imem06_bank = 0;
    27: _imem06_bank = 2;
    28: _imem06_bank = 0;
    29: _imem06_bank = 0;
    30: _imem06_bank = 3;
    31: _imem06_bank = 0;
    32: _imem06_bank = 0;
    33: _imem06_bank = 0;
    34: _imem06_bank = 1;
    35: _imem06_bank = 3;
    36: _imem06_bank = 0;
    37: _imem06_bank = 1;
    38: _imem06_bank = 0;
    39: _imem06_bank = 0;
    40: _imem06_bank = 0;
    41: _imem06_bank = 0;
    42: _imem06_bank = 0;
    43: _imem06_bank = 0;
    44: _imem06_bank = 0;
    45: _imem06_bank = 0;
    46: _imem06_bank = 0;
    47: _imem06_bank = 0;
    48: _imem06_bank = 0;
    49: _imem06_bank = 0;
    50: _imem06_bank = 0;
    51: _imem06_bank = 0;
    52: _imem06_bank = 0;
    53: _imem06_bank = 0;
    54: _imem06_bank = 0;
    55: _imem06_bank = 1;
    56: _imem06_bank = 2;
    57: _imem06_bank = 0;
    58: _imem06_bank = 0;
    59: _imem06_bank = 3;
    60: _imem06_bank = 0;
    61: _imem06_bank = 0;
    62: _imem06_bank = 0;
    63: _imem06_bank = 0;
    64: _imem06_bank = 0;
    65: _imem06_bank = 0;
    66: _imem06_bank = 0;
    67: _imem06_bank = 0;
    68: _imem06_bank = 0;
    69: _imem06_bank = 3;
    70: _imem06_bank = 0;
    71: _imem06_bank = 0;
    72: _imem06_bank = 0;
    73: _imem06_bank = 0;
    74: _imem06_bank = 0;
    75: _imem06_bank = 0;
    76: _imem06_bank = 0;
    77: _imem06_bank = 0;
    78: _imem06_bank = 0;
    79: _imem06_bank = 0;
    80: _imem06_bank = 0;
    81: _imem06_bank = 0;
    82: _imem06_bank = 0;
    83: _imem06_bank = 0;
    84: _imem06_bank = 2;
    85: _imem06_bank = 0;
    86: _imem06_bank = 0;
    87: _imem06_bank = 3;
    88: _imem06_bank = 0;
    89: _imem06_bank = 0;
    90: _imem06_bank = 0;
    91: _imem06_bank = 0;
    92: _imem06_bank = 0;
    93: _imem06_bank = 0;
    94: _imem06_bank = 0;
    95: _imem06_bank = 0;
    default: _imem06_bank = 0;
    endcase
  end // always @ ( * )
  assign imem06_bank = _imem06_bank;
  reg _imem06_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem06_rd = 1;
    2: _imem06_rd = 1;
    1: _imem06_rd = 1;
    0: _imem06_rd = 1;
    4: _imem06_rd = 1;
    5: _imem06_rd = 1;
    6: _imem06_rd = 1;
    7: _imem06_rd = 1;
    8: _imem06_rd = 1;
    9: _imem06_rd = 1;
    10: _imem06_rd = 1;
    11: _imem06_rd = 1;
    12: _imem06_rd = 1;
    13: _imem06_rd = 1;
    14: _imem06_rd = 1;
    15: _imem06_rd = 1;
    16: _imem06_rd = 1;
    17: _imem06_rd = 1;
    18: _imem06_rd = 1;
    19: _imem06_rd = 1;
    20: _imem06_rd = 1;
    21: _imem06_rd = 1;
    22: _imem06_rd = 1;
    23: _imem06_rd = 1;
    24: _imem06_rd = 1;
    25: _imem06_rd = 1;
    26: _imem06_rd = 1;
    27: _imem06_rd = 1;
    28: _imem06_rd = 1;
    29: _imem06_rd = 1;
    30: _imem06_rd = 1;
    31: _imem06_rd = 1;
    32: _imem06_rd = 1;
    33: _imem06_rd = 1;
    34: _imem06_rd = 1;
    35: _imem06_rd = 1;
    36: _imem06_rd = 1;
    37: _imem06_rd = 1;
    38: _imem06_rd = 1;
    39: _imem06_rd = 1;
    40: _imem06_rd = 1;
    41: _imem06_rd = 1;
    42: _imem06_rd = 1;
    43: _imem06_rd = 1;
    44: _imem06_rd = 1;
    45: _imem06_rd = 1;
    46: _imem06_rd = 1;
    47: _imem06_rd = 1;
    48: _imem06_rd = 1;
    49: _imem06_rd = 1;
    50: _imem06_rd = 1;
    51: _imem06_rd = 1;
    52: _imem06_rd = 1;
    53: _imem06_rd = 1;
    54: _imem06_rd = 1;
    55: _imem06_rd = 1;
    56: _imem06_rd = 1;
    57: _imem06_rd = 1;
    58: _imem06_rd = 1;
    59: _imem06_rd = 1;
    60: _imem06_rd = 1;
    61: _imem06_rd = 1;
    62: _imem06_rd = 1;
    63: _imem06_rd = 1;
    64: _imem06_rd = 1;
    65: _imem06_rd = 1;
    66: _imem06_rd = 1;
    67: _imem06_rd = 1;
    68: _imem06_rd = 1;
    69: _imem06_rd = 1;
    70: _imem06_rd = 1;
    71: _imem06_rd = 1;
    72: _imem06_rd = 1;
    73: _imem06_rd = 1;
    74: _imem06_rd = 1;
    75: _imem06_rd = 1;
    76: _imem06_rd = 1;
    77: _imem06_rd = 1;
    78: _imem06_rd = 1;
    79: _imem06_rd = 1;
    80: _imem06_rd = 1;
    81: _imem06_rd = 1;
    82: _imem06_rd = 1;
    83: _imem06_rd = 1;
    84: _imem06_rd = 1;
    85: _imem06_rd = 1;
    86: _imem06_rd = 1;
    87: _imem06_rd = 1;
    88: _imem06_rd = 1;
    89: _imem06_rd = 1;
    90: _imem06_rd = 1;
    91: _imem06_rd = 1;
    92: _imem06_rd = 1;
    93: _imem06_rd = 1;
    94: _imem06_rd = 1;
    95: _imem06_rd = 1;
    default: _imem06_rd = 0;
    endcase
  end // always @ ( * )
  assign imem06_rd = _imem06_rd;

  // 7番目の入力用メモリブロックの制御
  reg [1:0] _imem07_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem07_bank = 0;
    2: _imem07_bank = 1;
    1: _imem07_bank = 2;
    0: _imem07_bank = 3;
    4: _imem07_bank = 0;
    5: _imem07_bank = 0;
    6: _imem07_bank = 0;
    7: _imem07_bank = 0;
    8: _imem07_bank = 0;
    9: _imem07_bank = 0;
    10: _imem07_bank = 0;
    11: _imem07_bank = 0;
    12: _imem07_bank = 0;
    13: _imem07_bank = 0;
    14: _imem07_bank = 0;
    15: _imem07_bank = 0;
    16: _imem07_bank = 0;
    17: _imem07_bank = 0;
    18: _imem07_bank = 0;
    19: _imem07_bank = 0;
    20: _imem07_bank = 0;
    21: _imem07_bank = 0;
    22: _imem07_bank = 0;
    23: _imem07_bank = 0;
    24: _imem07_bank = 0;
    25: _imem07_bank = 0;
    26: _imem07_bank = 0;
    27: _imem07_bank = 0;
    28: _imem07_bank = 0;
    29: _imem07_bank = 0;
    30: _imem07_bank = 0;
    31: _imem07_bank = 0;
    32: _imem07_bank = 0;
    33: _imem07_bank = 0;
    34: _imem07_bank = 0;
    35: _imem07_bank = 0;
    36: _imem07_bank = 0;
    37: _imem07_bank = 0;
    38: _imem07_bank = 0;
    39: _imem07_bank = 0;
    40: _imem07_bank = 0;
    41: _imem07_bank = 2;
    42: _imem07_bank = 0;
    43: _imem07_bank = 0;
    44: _imem07_bank = 0;
    45: _imem07_bank = 0;
    46: _imem07_bank = 0;
    47: _imem07_bank = 0;
    48: _imem07_bank = 0;
    49: _imem07_bank = 0;
    50: _imem07_bank = 0;
    51: _imem07_bank = 0;
    52: _imem07_bank = 0;
    53: _imem07_bank = 0;
    54: _imem07_bank = 0;
    55: _imem07_bank = 0;
    56: _imem07_bank = 0;
    57: _imem07_bank = 0;
    58: _imem07_bank = 0;
    59: _imem07_bank = 0;
    60: _imem07_bank = 0;
    61: _imem07_bank = 0;
    62: _imem07_bank = 0;
    63: _imem07_bank = 0;
    64: _imem07_bank = 0;
    65: _imem07_bank = 0;
    66: _imem07_bank = 0;
    67: _imem07_bank = 0;
    68: _imem07_bank = 0;
    69: _imem07_bank = 0;
    70: _imem07_bank = 0;
    71: _imem07_bank = 0;
    72: _imem07_bank = 0;
    73: _imem07_bank = 1;
    74: _imem07_bank = 0;
    75: _imem07_bank = 0;
    76: _imem07_bank = 0;
    77: _imem07_bank = 1;
    78: _imem07_bank = 0;
    79: _imem07_bank = 3;
    80: _imem07_bank = 3;
    81: _imem07_bank = 0;
    82: _imem07_bank = 0;
    83: _imem07_bank = 0;
    84: _imem07_bank = 0;
    85: _imem07_bank = 0;
    86: _imem07_bank = 0;
    87: _imem07_bank = 0;
    88: _imem07_bank = 0;
    89: _imem07_bank = 0;
    90: _imem07_bank = 0;
    91: _imem07_bank = 0;
    92: _imem07_bank = 0;
    93: _imem07_bank = 0;
    94: _imem07_bank = 0;
    95: _imem07_bank = 0;
    default: _imem07_bank = 0;
    endcase
  end // always @ ( * )
  assign imem07_bank = _imem07_bank;
  reg _imem07_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem07_rd = 1;
    2: _imem07_rd = 1;
    1: _imem07_rd = 1;
    0: _imem07_rd = 1;
    4: _imem07_rd = 1;
    5: _imem07_rd = 1;
    6: _imem07_rd = 1;
    7: _imem07_rd = 1;
    8: _imem07_rd = 1;
    9: _imem07_rd = 1;
    10: _imem07_rd = 1;
    11: _imem07_rd = 1;
    12: _imem07_rd = 1;
    13: _imem07_rd = 1;
    14: _imem07_rd = 1;
    15: _imem07_rd = 1;
    16: _imem07_rd = 1;
    17: _imem07_rd = 1;
    18: _imem07_rd = 1;
    19: _imem07_rd = 1;
    20: _imem07_rd = 1;
    21: _imem07_rd = 1;
    22: _imem07_rd = 1;
    23: _imem07_rd = 1;
    24: _imem07_rd = 1;
    25: _imem07_rd = 1;
    26: _imem07_rd = 1;
    27: _imem07_rd = 1;
    28: _imem07_rd = 1;
    29: _imem07_rd = 1;
    30: _imem07_rd = 1;
    31: _imem07_rd = 1;
    32: _imem07_rd = 1;
    33: _imem07_rd = 1;
    34: _imem07_rd = 1;
    35: _imem07_rd = 1;
    36: _imem07_rd = 1;
    37: _imem07_rd = 1;
    38: _imem07_rd = 1;
    39: _imem07_rd = 1;
    40: _imem07_rd = 1;
    41: _imem07_rd = 1;
    42: _imem07_rd = 1;
    43: _imem07_rd = 1;
    44: _imem07_rd = 1;
    45: _imem07_rd = 1;
    46: _imem07_rd = 1;
    47: _imem07_rd = 1;
    48: _imem07_rd = 1;
    49: _imem07_rd = 1;
    50: _imem07_rd = 1;
    51: _imem07_rd = 1;
    52: _imem07_rd = 1;
    53: _imem07_rd = 1;
    54: _imem07_rd = 1;
    55: _imem07_rd = 1;
    56: _imem07_rd = 1;
    57: _imem07_rd = 1;
    58: _imem07_rd = 1;
    59: _imem07_rd = 1;
    60: _imem07_rd = 1;
    61: _imem07_rd = 1;
    62: _imem07_rd = 1;
    63: _imem07_rd = 1;
    64: _imem07_rd = 1;
    65: _imem07_rd = 1;
    66: _imem07_rd = 1;
    67: _imem07_rd = 1;
    68: _imem07_rd = 1;
    69: _imem07_rd = 1;
    70: _imem07_rd = 1;
    71: _imem07_rd = 1;
    72: _imem07_rd = 1;
    73: _imem07_rd = 1;
    74: _imem07_rd = 1;
    75: _imem07_rd = 1;
    76: _imem07_rd = 1;
    77: _imem07_rd = 1;
    78: _imem07_rd = 1;
    79: _imem07_rd = 1;
    80: _imem07_rd = 1;
    81: _imem07_rd = 1;
    82: _imem07_rd = 1;
    83: _imem07_rd = 1;
    84: _imem07_rd = 1;
    85: _imem07_rd = 1;
    86: _imem07_rd = 1;
    87: _imem07_rd = 1;
    88: _imem07_rd = 1;
    89: _imem07_rd = 1;
    90: _imem07_rd = 1;
    91: _imem07_rd = 1;
    92: _imem07_rd = 1;
    93: _imem07_rd = 1;
    94: _imem07_rd = 1;
    95: _imem07_rd = 1;
    default: _imem07_rd = 0;
    endcase
  end // always @ ( * )
  assign imem07_rd = _imem07_rd;

  // 0番目の出力用メモリブロックの制御
  reg [5:0] _omem00_bank;
  always @ ( * ) begin
    case ( state )
    7: _omem00_bank = 0;
    8: _omem00_bank = 1;
    9: _omem00_bank = 2;
    10: _omem00_bank = 3;
    11: _omem00_bank = 4;
    12: _omem00_bank = 5;
    13: _omem00_bank = 6;
    14: _omem00_bank = 7;
    15: _omem00_bank = 8;
    16: _omem00_bank = 9;
    17: _omem00_bank = 10;
    18: _omem00_bank = 11;
    19: _omem00_bank = 12;
    20: _omem00_bank = 13;
    21: _omem00_bank = 14;
    22: _omem00_bank = 15;
    23: _omem00_bank = 16;
    24: _omem00_bank = 17;
    25: _omem00_bank = 18;
    26: _omem00_bank = 19;
    27: _omem00_bank = 20;
    28: _omem00_bank = 21;
    29: _omem00_bank = 22;
    30: _omem00_bank = 23;
    31: _omem00_bank = 24;
    32: _omem00_bank = 25;
    33: _omem00_bank = 26;
    34: _omem00_bank = 27;
    35: _omem00_bank = 28;
    36: _omem00_bank = 29;
    37: _omem00_bank = 30;
    38: _omem00_bank = 31;
    39: _omem00_bank = 32;
    40: _omem00_bank = 33;
    41: _omem00_bank = 34;
    42: _omem00_bank = 35;
    43: _omem00_bank = 36;
    44: _omem00_bank = 37;
    45: _omem00_bank = 38;
    46: _omem00_bank = 39;
    47: _omem00_bank = 40;
    48: _omem00_bank = 41;
    49: _omem00_bank = 42;
    50: _omem00_bank = 43;
    51: _omem00_bank = 44;
    52: _omem00_bank = 45;
    53: _omem00_bank = 46;
    54: _omem00_bank = 47;
    55: _omem00_bank = 48;
    56: _omem00_bank = 49;
    57: _omem00_bank = 50;
    58: _omem00_bank = 51;
    59: _omem00_bank = 52;
    60: _omem00_bank = 53;
    61: _omem00_bank = 54;
    62: _omem00_bank = 55;
    63: _omem00_bank = 56;
    64: _omem00_bank = 57;
    65: _omem00_bank = 58;
    66: _omem00_bank = 59;
    default: _omem00_bank = 0;
    endcase
  end // always @ ( * )
  assign omem00_bank = _omem00_bank;
  reg _omem00_wr;
  always @ ( * ) begin
    case ( state )
    7: _omem00_wr = 1;
    8: _omem00_wr = 1;
    9: _omem00_wr = 1;
    10: _omem00_wr = 1;
    11: _omem00_wr = 1;
    12: _omem00_wr = 1;
    13: _omem00_wr = 1;
    14: _omem00_wr = 1;
    15: _omem00_wr = 1;
    16: _omem00_wr = 1;
    17: _omem00_wr = 1;
    18: _omem00_wr = 1;
    19: _omem00_wr = 1;
    20: _omem00_wr = 1;
    21: _omem00_wr = 1;
    22: _omem00_wr = 1;
    23: _omem00_wr = 1;
    24: _omem00_wr = 1;
    25: _omem00_wr = 1;
    26: _omem00_wr = 1;
    27: _omem00_wr = 1;
    28: _omem00_wr = 1;
    29: _omem00_wr = 1;
    30: _omem00_wr = 1;
    31: _omem00_wr = 1;
    32: _omem00_wr = 1;
    33: _omem00_wr = 1;
    34: _omem00_wr = 1;
    35: _omem00_wr = 1;
    36: _omem00_wr = 1;
    37: _omem00_wr = 1;
    38: _omem00_wr = 1;
    39: _omem00_wr = 1;
    40: _omem00_wr = 1;
    41: _omem00_wr = 1;
    42: _omem00_wr = 1;
    43: _omem00_wr = 1;
    44: _omem00_wr = 1;
    45: _omem00_wr = 1;
    46: _omem00_wr = 1;
    47: _omem00_wr = 1;
    48: _omem00_wr = 1;
    49: _omem00_wr = 1;
    50: _omem00_wr = 1;
    51: _omem00_wr = 1;
    52: _omem00_wr = 1;
    53: _omem00_wr = 1;
    54: _omem00_wr = 1;
    55: _omem00_wr = 1;
    56: _omem00_wr = 1;
    57: _omem00_wr = 1;
    58: _omem00_wr = 1;
    59: _omem00_wr = 1;
    60: _omem00_wr = 1;
    61: _omem00_wr = 1;
    62: _omem00_wr = 1;
    63: _omem00_wr = 1;
    64: _omem00_wr = 1;
    65: _omem00_wr = 1;
    66: _omem00_wr = 1;
    default: _omem00_wr = 0;
    endcase
  end // always @ ( * )
  assign omem00_wr = _omem00_wr;

  // 1番目の出力用メモリブロックの制御
  reg [5:0] _omem01_bank;
  always @ ( * ) begin
    case ( state )
    24: _omem01_bank = 0;
    25: _omem01_bank = 1;
    26: _omem01_bank = 2;
    27: _omem01_bank = 3;
    28: _omem01_bank = 4;
    29: _omem01_bank = 5;
    30: _omem01_bank = 6;
    31: _omem01_bank = 7;
    32: _omem01_bank = 8;
    33: _omem01_bank = 9;
    34: _omem01_bank = 10;
    35: _omem01_bank = 11;
    36: _omem01_bank = 12;
    37: _omem01_bank = 13;
    38: _omem01_bank = 14;
    39: _omem01_bank = 15;
    40: _omem01_bank = 16;
    41: _omem01_bank = 17;
    42: _omem01_bank = 18;
    43: _omem01_bank = 19;
    44: _omem01_bank = 20;
    45: _omem01_bank = 21;
    46: _omem01_bank = 22;
    47: _omem01_bank = 23;
    48: _omem01_bank = 24;
    49: _omem01_bank = 25;
    50: _omem01_bank = 26;
    51: _omem01_bank = 27;
    52: _omem01_bank = 28;
    53: _omem01_bank = 29;
    54: _omem01_bank = 30;
    55: _omem01_bank = 31;
    56: _omem01_bank = 32;
    57: _omem01_bank = 33;
    58: _omem01_bank = 34;
    59: _omem01_bank = 35;
    60: _omem01_bank = 36;
    61: _omem01_bank = 37;
    62: _omem01_bank = 38;
    63: _omem01_bank = 39;
    64: _omem01_bank = 40;
    65: _omem01_bank = 41;
    66: _omem01_bank = 42;
    67: _omem01_bank = 43;
    68: _omem01_bank = 44;
    69: _omem01_bank = 45;
    70: _omem01_bank = 46;
    71: _omem01_bank = 47;
    72: _omem01_bank = 48;
    73: _omem01_bank = 49;
    74: _omem01_bank = 50;
    75: _omem01_bank = 51;
    76: _omem01_bank = 52;
    77: _omem01_bank = 53;
    78: _omem01_bank = 54;
    79: _omem01_bank = 55;
    80: _omem01_bank = 56;
    81: _omem01_bank = 57;
    82: _omem01_bank = 58;
    83: _omem01_bank = 59;
    default: _omem01_bank = 0;
    endcase
  end // always @ ( * )
  assign omem01_bank = _omem01_bank;
  reg _omem01_wr;
  always @ ( * ) begin
    case ( state )
    24: _omem01_wr = 1;
    25: _omem01_wr = 1;
    26: _omem01_wr = 1;
    27: _omem01_wr = 1;
    28: _omem01_wr = 1;
    29: _omem01_wr = 1;
    30: _omem01_wr = 1;
    31: _omem01_wr = 1;
    32: _omem01_wr = 1;
    33: _omem01_wr = 1;
    34: _omem01_wr = 1;
    35: _omem01_wr = 1;
    36: _omem01_wr = 1;
    37: _omem01_wr = 1;
    38: _omem01_wr = 1;
    39: _omem01_wr = 1;
    40: _omem01_wr = 1;
    41: _omem01_wr = 1;
    42: _omem01_wr = 1;
    43: _omem01_wr = 1;
    44: _omem01_wr = 1;
    45: _omem01_wr = 1;
    46: _omem01_wr = 1;
    47: _omem01_wr = 1;
    48: _omem01_wr = 1;
    49: _omem01_wr = 1;
    50: _omem01_wr = 1;
    51: _omem01_wr = 1;
    52: _omem01_wr = 1;
    53: _omem01_wr = 1;
    54: _omem01_wr = 1;
    55: _omem01_wr = 1;
    56: _omem01_wr = 1;
    57: _omem01_wr = 1;
    58: _omem01_wr = 1;
    59: _omem01_wr = 1;
    60: _omem01_wr = 1;
    61: _omem01_wr = 1;
    62: _omem01_wr = 1;
    63: _omem01_wr = 1;
    64: _omem01_wr = 1;
    65: _omem01_wr = 1;
    66: _omem01_wr = 1;
    67: _omem01_wr = 1;
    68: _omem01_wr = 1;
    69: _omem01_wr = 1;
    70: _omem01_wr = 1;
    71: _omem01_wr = 1;
    72: _omem01_wr = 1;
    73: _omem01_wr = 1;
    74: _omem01_wr = 1;
    75: _omem01_wr = 1;
    76: _omem01_wr = 1;
    77: _omem01_wr = 1;
    78: _omem01_wr = 1;
    79: _omem01_wr = 1;
    80: _omem01_wr = 1;
    81: _omem01_wr = 1;
    82: _omem01_wr = 1;
    83: _omem01_wr = 1;
    default: _omem01_wr = 0;
    endcase
  end // always @ ( * )
  assign omem01_wr = _omem01_wr;

  // 2番目の出力用メモリブロックの制御
  reg [5:0] _omem02_bank;
  always @ ( * ) begin
    case ( state )
    43: _omem02_bank = 0;
    44: _omem02_bank = 1;
    45: _omem02_bank = 2;
    46: _omem02_bank = 3;
    47: _omem02_bank = 4;
    48: _omem02_bank = 5;
    49: _omem02_bank = 6;
    50: _omem02_bank = 7;
    51: _omem02_bank = 8;
    52: _omem02_bank = 9;
    53: _omem02_bank = 10;
    54: _omem02_bank = 11;
    55: _omem02_bank = 12;
    56: _omem02_bank = 13;
    57: _omem02_bank = 14;
    58: _omem02_bank = 15;
    59: _omem02_bank = 16;
    60: _omem02_bank = 17;
    61: _omem02_bank = 18;
    62: _omem02_bank = 19;
    63: _omem02_bank = 20;
    64: _omem02_bank = 21;
    65: _omem02_bank = 22;
    66: _omem02_bank = 23;
    67: _omem02_bank = 24;
    68: _omem02_bank = 25;
    69: _omem02_bank = 26;
    70: _omem02_bank = 27;
    71: _omem02_bank = 28;
    72: _omem02_bank = 29;
    73: _omem02_bank = 30;
    74: _omem02_bank = 31;
    75: _omem02_bank = 32;
    76: _omem02_bank = 33;
    77: _omem02_bank = 34;
    78: _omem02_bank = 35;
    79: _omem02_bank = 36;
    80: _omem02_bank = 37;
    81: _omem02_bank = 38;
    82: _omem02_bank = 39;
    83: _omem02_bank = 40;
    84: _omem02_bank = 41;
    85: _omem02_bank = 42;
    86: _omem02_bank = 43;
    87: _omem02_bank = 44;
    88: _omem02_bank = 45;
    89: _omem02_bank = 46;
    90: _omem02_bank = 47;
    91: _omem02_bank = 48;
    92: _omem02_bank = 49;
    93: _omem02_bank = 50;
    94: _omem02_bank = 51;
    95: _omem02_bank = 52;
    96: _omem02_bank = 53;
    97: _omem02_bank = 54;
    98: _omem02_bank = 55;
    99: _omem02_bank = 56;
    100: _omem02_bank = 57;
    101: _omem02_bank = 58;
    102: _omem02_bank = 59;
    default: _omem02_bank = 0;
    endcase
  end // always @ ( * )
  assign omem02_bank = _omem02_bank;
  reg _omem02_wr;
  always @ ( * ) begin
    case ( state )
    43: _omem02_wr = 1;
    44: _omem02_wr = 1;
    45: _omem02_wr = 1;
    46: _omem02_wr = 1;
    47: _omem02_wr = 1;
    48: _omem02_wr = 1;
    49: _omem02_wr = 1;
    50: _omem02_wr = 1;
    51: _omem02_wr = 1;
    52: _omem02_wr = 1;
    53: _omem02_wr = 1;
    54: _omem02_wr = 1;
    55: _omem02_wr = 1;
    56: _omem02_wr = 1;
    57: _omem02_wr = 1;
    58: _omem02_wr = 1;
    59: _omem02_wr = 1;
    60: _omem02_wr = 1;
    61: _omem02_wr = 1;
    62: _omem02_wr = 1;
    63: _omem02_wr = 1;
    64: _omem02_wr = 1;
    65: _omem02_wr = 1;
    66: _omem02_wr = 1;
    67: _omem02_wr = 1;
    68: _omem02_wr = 1;
    69: _omem02_wr = 1;
    70: _omem02_wr = 1;
    71: _omem02_wr = 1;
    72: _omem02_wr = 1;
    73: _omem02_wr = 1;
    74: _omem02_wr = 1;
    75: _omem02_wr = 1;
    76: _omem02_wr = 1;
    77: _omem02_wr = 1;
    78: _omem02_wr = 1;
    79: _omem02_wr = 1;
    80: _omem02_wr = 1;
    81: _omem02_wr = 1;
    82: _omem02_wr = 1;
    83: _omem02_wr = 1;
    84: _omem02_wr = 1;
    85: _omem02_wr = 1;
    86: _omem02_wr = 1;
    87: _omem02_wr = 1;
    88: _omem02_wr = 1;
    89: _omem02_wr = 1;
    90: _omem02_wr = 1;
    91: _omem02_wr = 1;
    92: _omem02_wr = 1;
    93: _omem02_wr = 1;
    94: _omem02_wr = 1;
    95: _omem02_wr = 1;
    96: _omem02_wr = 1;
    97: _omem02_wr = 1;
    98: _omem02_wr = 1;
    99: _omem02_wr = 1;
    100: _omem02_wr = 1;
    101: _omem02_wr = 1;
    102: _omem02_wr = 1;
    default: _omem02_wr = 0;
    endcase
  end // always @ ( * )
  assign omem02_wr = _omem02_wr;

  // 3番目の出力用メモリブロックの制御
  reg [5:0] _omem03_bank;
  always @ ( * ) begin
    case ( state )
    62: _omem03_bank = 0;
    63: _omem03_bank = 1;
    64: _omem03_bank = 2;
    65: _omem03_bank = 3;
    66: _omem03_bank = 4;
    67: _omem03_bank = 5;
    68: _omem03_bank = 6;
    69: _omem03_bank = 7;
    70: _omem03_bank = 8;
    71: _omem03_bank = 9;
    72: _omem03_bank = 10;
    73: _omem03_bank = 11;
    74: _omem03_bank = 12;
    75: _omem03_bank = 13;
    76: _omem03_bank = 14;
    77: _omem03_bank = 15;
    78: _omem03_bank = 16;
    79: _omem03_bank = 17;
    80: _omem03_bank = 18;
    81: _omem03_bank = 19;
    82: _omem03_bank = 20;
    83: _omem03_bank = 21;
    84: _omem03_bank = 22;
    85: _omem03_bank = 23;
    86: _omem03_bank = 24;
    87: _omem03_bank = 25;
    88: _omem03_bank = 26;
    89: _omem03_bank = 27;
    90: _omem03_bank = 28;
    91: _omem03_bank = 29;
    92: _omem03_bank = 30;
    93: _omem03_bank = 31;
    94: _omem03_bank = 32;
    95: _omem03_bank = 33;
    96: _omem03_bank = 34;
    97: _omem03_bank = 35;
    98: _omem03_bank = 36;
    99: _omem03_bank = 37;
    100: _omem03_bank = 38;
    101: _omem03_bank = 39;
    102: _omem03_bank = 40;
    103: _omem03_bank = 41;
    104: _omem03_bank = 42;
    105: _omem03_bank = 43;
    106: _omem03_bank = 44;
    107: _omem03_bank = 45;
    108: _omem03_bank = 46;
    109: _omem03_bank = 47;
    110: _omem03_bank = 48;
    111: _omem03_bank = 49;
    112: _omem03_bank = 50;
    113: _omem03_bank = 51;
    114: _omem03_bank = 52;
    115: _omem03_bank = 53;
    116: _omem03_bank = 54;
    117: _omem03_bank = 55;
    118: _omem03_bank = 56;
    119: _omem03_bank = 57;
    120: _omem03_bank = 58;
    121: _omem03_bank = 59;
    default: _omem03_bank = 0;
    endcase
  end // always @ ( * )
  assign omem03_bank = _omem03_bank;
  reg _omem03_wr;
  always @ ( * ) begin
    case ( state )
    62: _omem03_wr = 1;
    63: _omem03_wr = 1;
    64: _omem03_wr = 1;
    65: _omem03_wr = 1;
    66: _omem03_wr = 1;
    67: _omem03_wr = 1;
    68: _omem03_wr = 1;
    69: _omem03_wr = 1;
    70: _omem03_wr = 1;
    71: _omem03_wr = 1;
    72: _omem03_wr = 1;
    73: _omem03_wr = 1;
    74: _omem03_wr = 1;
    75: _omem03_wr = 1;
    76: _omem03_wr = 1;
    77: _omem03_wr = 1;
    78: _omem03_wr = 1;
    79: _omem03_wr = 1;
    80: _omem03_wr = 1;
    81: _omem03_wr = 1;
    82: _omem03_wr = 1;
    83: _omem03_wr = 1;
    84: _omem03_wr = 1;
    85: _omem03_wr = 1;
    86: _omem03_wr = 1;
    87: _omem03_wr = 1;
    88: _omem03_wr = 1;
    89: _omem03_wr = 1;
    90: _omem03_wr = 1;
    91: _omem03_wr = 1;
    92: _omem03_wr = 1;
    93: _omem03_wr = 1;
    94: _omem03_wr = 1;
    95: _omem03_wr = 1;
    96: _omem03_wr = 1;
    97: _omem03_wr = 1;
    98: _omem03_wr = 1;
    99: _omem03_wr = 1;
    100: _omem03_wr = 1;
    101: _omem03_wr = 1;
    102: _omem03_wr = 1;
    103: _omem03_wr = 1;
    104: _omem03_wr = 1;
    105: _omem03_wr = 1;
    106: _omem03_wr = 1;
    107: _omem03_wr = 1;
    108: _omem03_wr = 1;
    109: _omem03_wr = 1;
    110: _omem03_wr = 1;
    111: _omem03_wr = 1;
    112: _omem03_wr = 1;
    113: _omem03_wr = 1;
    114: _omem03_wr = 1;
    115: _omem03_wr = 1;
    116: _omem03_wr = 1;
    117: _omem03_wr = 1;
    118: _omem03_wr = 1;
    119: _omem03_wr = 1;
    120: _omem03_wr = 1;
    121: _omem03_wr = 1;
    default: _omem03_wr = 0;
    endcase
  end // always @ ( * )
  assign omem03_wr = _omem03_wr;

  // 4番目の出力用メモリブロックの制御
  reg [5:0] _omem04_bank;
  always @ ( * ) begin
    case ( state )
    81: _omem04_bank = 0;
    82: _omem04_bank = 1;
    83: _omem04_bank = 2;
    84: _omem04_bank = 3;
    85: _omem04_bank = 4;
    86: _omem04_bank = 5;
    87: _omem04_bank = 6;
    88: _omem04_bank = 7;
    89: _omem04_bank = 8;
    90: _omem04_bank = 9;
    91: _omem04_bank = 10;
    92: _omem04_bank = 11;
    93: _omem04_bank = 12;
    94: _omem04_bank = 13;
    95: _omem04_bank = 14;
    96: _omem04_bank = 15;
    97: _omem04_bank = 16;
    98: _omem04_bank = 17;
    99: _omem04_bank = 18;
    100: _omem04_bank = 19;
    101: _omem04_bank = 20;
    102: _omem04_bank = 21;
    103: _omem04_bank = 22;
    104: _omem04_bank = 23;
    105: _omem04_bank = 24;
    106: _omem04_bank = 25;
    107: _omem04_bank = 26;
    108: _omem04_bank = 27;
    109: _omem04_bank = 28;
    110: _omem04_bank = 29;
    111: _omem04_bank = 30;
    112: _omem04_bank = 31;
    113: _omem04_bank = 32;
    114: _omem04_bank = 33;
    115: _omem04_bank = 34;
    116: _omem04_bank = 35;
    117: _omem04_bank = 36;
    118: _omem04_bank = 37;
    119: _omem04_bank = 38;
    120: _omem04_bank = 39;
    121: _omem04_bank = 40;
    122: _omem04_bank = 41;
    123: _omem04_bank = 42;
    124: _omem04_bank = 43;
    125: _omem04_bank = 44;
    126: _omem04_bank = 45;
    127: _omem04_bank = 46;
    128: _omem04_bank = 47;
    129: _omem04_bank = 48;
    130: _omem04_bank = 49;
    131: _omem04_bank = 50;
    132: _omem04_bank = 51;
    133: _omem04_bank = 52;
    134: _omem04_bank = 53;
    135: _omem04_bank = 54;
    136: _omem04_bank = 55;
    137: _omem04_bank = 56;
    138: _omem04_bank = 57;
    default: _omem04_bank = 0;
    endcase
  end // always @ ( * )
  assign omem04_bank = _omem04_bank;
  reg _omem04_wr;
  always @ ( * ) begin
    case ( state )
    81: _omem04_wr = 1;
    82: _omem04_wr = 1;
    83: _omem04_wr = 1;
    84: _omem04_wr = 1;
    85: _omem04_wr = 1;
    86: _omem04_wr = 1;
    87: _omem04_wr = 1;
    88: _omem04_wr = 1;
    89: _omem04_wr = 1;
    90: _omem04_wr = 1;
    91: _omem04_wr = 1;
    92: _omem04_wr = 1;
    93: _omem04_wr = 1;
    94: _omem04_wr = 1;
    95: _omem04_wr = 1;
    96: _omem04_wr = 1;
    97: _omem04_wr = 1;
    98: _omem04_wr = 1;
    99: _omem04_wr = 1;
    100: _omem04_wr = 1;
    101: _omem04_wr = 1;
    102: _omem04_wr = 1;
    103: _omem04_wr = 1;
    104: _omem04_wr = 1;
    105: _omem04_wr = 1;
    106: _omem04_wr = 1;
    107: _omem04_wr = 1;
    108: _omem04_wr = 1;
    109: _omem04_wr = 1;
    110: _omem04_wr = 1;
    111: _omem04_wr = 1;
    112: _omem04_wr = 1;
    113: _omem04_wr = 1;
    114: _omem04_wr = 1;
    115: _omem04_wr = 1;
    116: _omem04_wr = 1;
    117: _omem04_wr = 1;
    118: _omem04_wr = 1;
    119: _omem04_wr = 1;
    120: _omem04_wr = 1;
    121: _omem04_wr = 1;
    122: _omem04_wr = 1;
    123: _omem04_wr = 1;
    124: _omem04_wr = 1;
    125: _omem04_wr = 1;
    126: _omem04_wr = 1;
    127: _omem04_wr = 1;
    128: _omem04_wr = 1;
    129: _omem04_wr = 1;
    130: _omem04_wr = 1;
    131: _omem04_wr = 1;
    132: _omem04_wr = 1;
    133: _omem04_wr = 1;
    134: _omem04_wr = 1;
    135: _omem04_wr = 1;
    136: _omem04_wr = 1;
    137: _omem04_wr = 1;
    138: _omem04_wr = 1;
    default: _omem04_wr = 0;
    endcase
  end // always @ ( * )
  assign omem04_wr = _omem04_wr;
  reg [8:0] _omem00_out;
  always @ ( * ) begin
    case ( state )
    7: _omem00_out = reg_1012;
    8: _omem00_out = reg_1013;
    9: _omem00_out = reg_1014;
    10: _omem00_out = reg_1024;
    11: _omem00_out = reg_1025;
    12: _omem00_out = reg_1026;
    13: _omem00_out = reg_1027;
    14: _omem00_out = reg_1012;
    15: _omem00_out = reg_0796;
    16: _omem00_out = reg_0797;
    17: _omem00_out = reg_0922;
    18: _omem00_out = reg_1013;
    19: _omem00_out = reg_0924;
    20: _omem00_out = reg_1047;
    21: _omem00_out = reg_1048;
    22: _omem00_out = reg_1014;
    23: _omem00_out = reg_1054;
    24: _omem00_out = reg_1024;
    25: _omem00_out = reg_0910;
    26: _omem00_out = reg_0911;
    27: _omem00_out = reg_0789;
    28: _omem00_out = reg_1025;
    29: _omem00_out = reg_0790;
    30: _omem00_out = reg_0890;
    31: _omem00_out = reg_0891;
    32: _omem00_out = reg_1026;
    33: _omem00_out = reg_0893;
    34: _omem00_out = reg_0498;
    35: _omem00_out = reg_0504;
    36: _omem00_out = reg_0505;
    37: _omem00_out = reg_1012;
    38: _omem00_out = reg_0878;
    39: _omem00_out = reg_0879;
    40: _omem00_out = reg_1027;
    41: _omem00_out = reg_0901;
    42: _omem00_out = reg_0796;
    43: _omem00_out = reg_0920;
    44: _omem00_out = reg_0770;
    45: _omem00_out = reg_0791;
    46: _omem00_out = reg_0797;
    47: _omem00_out = reg_0771;
    48: _omem00_out = reg_0794;
    49: _omem00_out = reg_0812;
    50: _omem00_out = reg_0841;
    51: _omem00_out = reg_1013;
    52: _omem00_out = reg_0859;
    53: _omem00_out = reg_0862;
    54: _omem00_out = reg_0742;
    55: _omem00_out = reg_0746;
    56: _omem00_out = reg_0924;
    57: _omem00_out = reg_1047;
    58: _omem00_out = reg_0839;
    59: _omem00_out = reg_0858;
    60: _omem00_out = reg_0861;
    61: _omem00_out = reg_0922;
    62: _omem00_out = reg_1048;
    63: _omem00_out = reg_0881;
    64: _omem00_out = reg_0929;
    65: _omem00_out = reg_0930;
    66: _omem00_out = reg_1014;
    default: _omem00_out = 0;
    endcase
  end // always @ ( * )
  assign omem00_out = _omem00_out[8:0];
  reg [8:0] _omem01_out;
  always @ ( * ) begin
    case ( state )
    24: _omem01_out = reg_0903;
    25: _omem01_out = reg_0527;
    26: _omem01_out = reg_0549;
    27: _omem01_out = reg_0553;
    28: _omem01_out = reg_1024;
    29: _omem01_out = reg_0559;
    30: _omem01_out = reg_0747;
    31: _omem01_out = reg_0903;
    32: _omem01_out = reg_0527;
    33: _omem01_out = reg_0910;
    34: _omem01_out = reg_0788;
    35: _omem01_out = reg_0766;
    36: _omem01_out = reg_0549;
    37: _omem01_out = reg_0911;
    38: _omem01_out = reg_1054;
    39: _omem01_out = reg_0362;
    40: _omem01_out = reg_0379;
    41: _omem01_out = reg_0553;
    42: _omem01_out = reg_1024;
    43: _omem01_out = reg_1025;
    44: _omem01_out = reg_0548;
    45: _omem01_out = reg_0934;
    46: _omem01_out = reg_0559;
    47: _omem01_out = reg_0936;
    48: _omem01_out = reg_0939;
    49: _omem01_out = reg_0600;
    50: _omem01_out = reg_0601;
    51: _omem01_out = reg_0747;
    52: _omem01_out = reg_0801;
    53: _omem01_out = reg_0891;
    54: _omem01_out = reg_0790;
    55: _omem01_out = reg_0527;
    56: _omem01_out = reg_0880;
    57: _omem01_out = reg_1026;
    58: _omem01_out = reg_0887;
    59: _omem01_out = reg_0789;
    60: _omem01_out = reg_0910;
    61: _omem01_out = reg_0800;
    62: _omem01_out = reg_0498;
    63: _omem01_out = reg_0598;
    64: _omem01_out = reg_0788;
    65: _omem01_out = reg_0766;
    66: _omem01_out = reg_0504;
    67: _omem01_out = reg_0561;
    68: _omem01_out = reg_0602;
    69: _omem01_out = reg_0549;
    70: _omem01_out = reg_0505;
    71: _omem01_out = reg_0890;
    72: _omem01_out = reg_0898;
    73: _omem01_out = reg_0911;
    74: _omem01_out = reg_0903;
    75: _omem01_out = reg_1012;
    76: _omem01_out = reg_0878;
    77: _omem01_out = reg_0402;
    78: _omem01_out = reg_0362;
    79: _omem01_out = reg_0606;
    80: _omem01_out = reg_0879;
    81: _omem01_out = reg_0638;
    82: _omem01_out = reg_0379;
    83: _omem01_out = reg_0775;
    default: _omem01_out = 0;
    endcase
  end // always @ ( * )
  assign omem01_out = _omem01_out[8:0];
  reg [8:0] _omem02_out;
  always @ ( * ) begin
    case ( state )
    43: _omem02_out = reg_0901;
    44: _omem02_out = reg_0587;
    45: _omem02_out = reg_0553;
    46: _omem02_out = reg_1024;
    47: _omem02_out = reg_0796;
    48: _omem02_out = reg_0557;
    49: _omem02_out = reg_0618;
    50: _omem02_out = reg_1025;
    51: _omem02_out = reg_0920;
    52: _omem02_out = reg_1027;
    53: _omem02_out = reg_0770;
    54: _omem02_out = reg_0587;
    55: _omem02_out = reg_0582;
    56: _omem02_out = reg_0901;
    57: _omem02_out = reg_0659;
    58: _omem02_out = reg_0553;
    59: _omem02_out = reg_0934;
    60: _omem02_out = reg_0559;
    61: _omem02_out = reg_0548;
    62: _omem02_out = reg_1054;
    63: _omem02_out = reg_1024;
    64: _omem02_out = reg_0796;
    65: _omem02_out = reg_0797;
    66: _omem02_out = reg_0544;
    67: _omem02_out = reg_0546;
    68: _omem02_out = reg_0551;
    69: _omem02_out = reg_0600;
    70: _omem02_out = reg_0791;
    71: _omem02_out = reg_0812;
    72: _omem02_out = reg_0618;
    73: _omem02_out = reg_0601;
    74: _omem02_out = reg_0557;
    75: _omem02_out = reg_0771;
    76: _omem02_out = reg_1013;
    77: _omem02_out = reg_0920;
    78: _omem02_out = reg_0801;
    79: _omem02_out = reg_0794;
    80: _omem02_out = reg_0859;
    81: _omem02_out = reg_0770;
    82: _omem02_out = reg_1025;
    83: _omem02_out = reg_0747;
    84: _omem02_out = reg_0742;
    85: _omem02_out = reg_0587;
    86: _omem02_out = reg_0790;
    87: _omem02_out = reg_0527;
    88: _omem02_out = reg_0891;
    89: _omem02_out = reg_0665;
    90: _omem02_out = reg_0751;
    91: _omem02_out = reg_0880;
    92: _omem02_out = reg_0924;
    93: _omem02_out = reg_1047;
    94: _omem02_out = reg_0659;
    95: _omem02_out = reg_0582;
    96: _omem02_out = reg_0901;
    97: _omem02_out = reg_0839;
    98: _omem02_out = reg_1026;
    99: _omem02_out = reg_0934;
    100: _omem02_out = reg_0746;
    101: _omem02_out = reg_0858;
    102: _omem02_out = reg_0939;
    default: _omem02_out = 0;
    endcase
  end // always @ ( * )
  assign omem02_out = _omem02_out[8:0];
  reg [8:0] _omem03_out;
  always @ ( * ) begin
    case ( state )
    62: _omem03_out = reg_0629;
    63: _omem03_out = reg_0559;
    64: _omem03_out = reg_0922;
    65: _omem03_out = reg_0910;
    66: _omem03_out = reg_0548;
    67: _omem03_out = reg_1027;
    68: _omem03_out = reg_0629;
    69: _omem03_out = reg_1048;
    70: _omem03_out = reg_0553;
    71: _omem03_out = reg_0789;
    72: _omem03_out = reg_0598;
    73: _omem03_out = reg_0881;
    74: _omem03_out = reg_0498;
    75: _omem03_out = reg_0796;
    76: _omem03_out = reg_0388;
    77: _omem03_out = reg_0766;
    78: _omem03_out = reg_0559;
    79: _omem03_out = reg_0797;
    80: _omem03_out = reg_0922;
    81: _omem03_out = reg_0910;
    82: _omem03_out = reg_0548;
    83: _omem03_out = reg_0929;
    84: _omem03_out = reg_0930;
    85: _omem03_out = reg_0561;
    86: _omem03_out = reg_0602;
    87: _omem03_out = reg_0504;
    88: _omem03_out = reg_0936;
    89: _omem03_out = reg_1027;
    90: _omem03_out = reg_0544;
    91: _omem03_out = reg_0549;
    92: _omem03_out = reg_0800;
    93: _omem03_out = reg_0600;
    94: _omem03_out = reg_0791;
    95: _omem03_out = reg_0505;
    96: _omem03_out = reg_0629;
    97: _omem03_out = reg_1048;
    98: _omem03_out = reg_0812;
    99: _omem03_out = reg_1054;
    100: _omem03_out = reg_0618;
    101: _omem03_out = reg_0898;
    102: _omem03_out = reg_0553;
    103: _omem03_out = reg_0890;
    104: _omem03_out = reg_0601;
    105: _omem03_out = reg_0911;
    106: _omem03_out = reg_0498;
    107: _omem03_out = reg_0598;
    108: _omem03_out = reg_0557;
    109: _omem03_out = reg_0771;
    110: _omem03_out = reg_0796;
    111: _omem03_out = reg_0881;
    112: _omem03_out = reg_0861;
    113: _omem03_out = reg_1012;
    114: _omem03_out = reg_0878;
    115: _omem03_out = reg_0388;
    116: _omem03_out = reg_0766;
    117: _omem03_out = reg_1013;
    118: _omem03_out = reg_0920;
    119: _omem03_out = reg_0362;
    120: _omem03_out = reg_0559;
    121: _omem03_out = reg_0801;
    default: _omem03_out = 0;
    endcase
  end // always @ ( * )
  assign omem03_out = _omem03_out[8:0];
  reg [8:0] _omem04_out;
  always @ ( * ) begin
    case ( state )
    81: _omem04_out = reg_0789;
    82: _omem04_out = reg_0606;
    83: _omem04_out = reg_0788;
    84: _omem04_out = reg_0922;
    85: _omem04_out = reg_0649;
    86: _omem04_out = reg_0859;
    87: _omem04_out = reg_0770;
    88: _omem04_out = reg_0910;
    89: _omem04_out = reg_0402;
    90: _omem04_out = reg_0789;
    91: _omem04_out = reg_1025;
    92: _omem04_out = reg_0548;
    93: _omem04_out = reg_0929;
    94: _omem04_out = reg_0794;
    95: _omem04_out = reg_0797;
    96: _omem04_out = reg_0742;
    97: _omem04_out = reg_0930;
    98: _omem04_out = reg_0840;
    99: _omem04_out = reg_0638;
    100: _omem04_out = reg_0649;
    101: _omem04_out = reg_0561;
    102: _omem04_out = reg_0602;
    103: _omem04_out = reg_0835;
    104: _omem04_out = reg_0790;
    105: _omem04_out = reg_0527;
    106: _omem04_out = reg_0504;
    107: _omem04_out = reg_0747;
    108: _omem04_out = reg_0922;
    109: _omem04_out = reg_0546;
    110: _omem04_out = reg_0936;
    111: _omem04_out = reg_0770;
    112: _omem04_out = reg_0910;
    113: _omem04_out = reg_0402;
    114: _omem04_out = reg_1027;
    115: _omem04_out = reg_0751;
    116: _omem04_out = reg_0576;
    117: _omem04_out = reg_0665;
    118: _omem04_out = reg_0841;
    119: _omem04_out = reg_0549;
    120: _omem04_out = reg_0633;
    121: _omem04_out = reg_0189;
    122: _omem04_out = reg_0880;
    123: _omem04_out = reg_0548;
    124: _omem04_out = reg_0862;
    125: _omem04_out = reg_0600;
    126: _omem04_out = reg_0379;
    127: _omem04_out = reg_0800;
    128: _omem04_out = reg_0929;
    129: _omem04_out = reg_0587;
    130: _omem04_out = reg_0879;
    131: _omem04_out = reg_1024;
    132: _omem04_out = reg_0659;
    133: _omem04_out = reg_0551;
    134: _omem04_out = reg_0544;
    135: _omem04_out = reg_0606;
    136: _omem04_out = reg_0582;
    137: _omem04_out = reg_0629;
    138: _omem04_out = reg_0791;
    default: _omem04_out = 0;
    endcase
  end // always @ ( * )
  assign omem04_out = _omem04_out[8:0];

  // OP1#0の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in00 = imem00_in[59:56];
    3: op1_00_in00 = imem07_in[123:120];
    6: op1_00_in00 = imem03_in[95:92];
    4: op1_00_in00 = imem07_in[91:88];
    7: op1_00_in00 = imem00_in[23:20];
    2: op1_00_in00 = imem07_in[115:112];
    8: op1_00_in00 = imem04_in[103:100];
    9: op1_00_in00 = imem06_in[107:104];
    10: op1_00_in00 = imem01_in[107:104];
    11: op1_00_in00 = imem01_in[83:80];
    25: op1_00_in00 = imem01_in[83:80];
    12: op1_00_in00 = imem05_in[99:96];
    13: op1_00_in00 = imem00_in[7:4];
    14: op1_00_in00 = imem05_in[103:100];
    15: op1_00_in00 = imem00_in[27:24];
    30: op1_00_in00 = imem00_in[27:24];
    60: op1_00_in00 = imem00_in[27:24];
    77: op1_00_in00 = imem00_in[27:24];
    16: op1_00_in00 = imem00_in[11:8];
    39: op1_00_in00 = imem00_in[11:8];
    17: op1_00_in00 = imem03_in[91:88];
    18: op1_00_in00 = imem04_in[115:112];
    19: op1_00_in00 = imem04_in[31:28];
    20: op1_00_in00 = imem05_in[35:32];
    21: op1_00_in00 = imem02_in[15:12];
    22: op1_00_in00 = imem06_in[95:92];
    58: op1_00_in00 = imem06_in[95:92];
    23: op1_00_in00 = imem00_in[107:104];
    24: op1_00_in00 = imem04_in[111:108];
    26: op1_00_in00 = imem02_in[119:116];
    27: op1_00_in00 = imem00_in[3:0];
    38: op1_00_in00 = imem00_in[3:0];
    28: op1_00_in00 = imem03_in[127:124];
    29: op1_00_in00 = imem06_in[11:8];
    31: op1_00_in00 = imem03_in[99:96];
    55: op1_00_in00 = imem03_in[99:96];
    32: op1_00_in00 = imem06_in[15:12];
    67: op1_00_in00 = imem06_in[15:12];
    33: op1_00_in00 = imem00_in[35:32];
    47: op1_00_in00 = imem00_in[35:32];
    34: op1_00_in00 = imem00_in[43:40];
    35: op1_00_in00 = imem06_in[111:108];
    36: op1_00_in00 = imem06_in[63:60];
    71: op1_00_in00 = imem06_in[63:60];
    37: op1_00_in00 = imem06_in[103:100];
    40: op1_00_in00 = imem01_in[119:116];
    41: op1_00_in00 = imem01_in[79:76];
    42: op1_00_in00 = imem04_in[59:56];
    43: op1_00_in00 = imem07_in[107:104];
    44: op1_00_in00 = imem00_in[19:16];
    45: op1_00_in00 = imem02_in[63:60];
    72: op1_00_in00 = imem02_in[63:60];
    46: op1_00_in00 = imem04_in[23:20];
    48: op1_00_in00 = imem01_in[71:68];
    49: op1_00_in00 = imem04_in[79:76];
    50: op1_00_in00 = imem05_in[95:92];
    51: op1_00_in00 = imem04_in[95:92];
    52: op1_00_in00 = imem02_in[39:36];
    53: op1_00_in00 = imem01_in[99:96];
    54: op1_00_in00 = imem03_in[55:52];
    56: op1_00_in00 = imem05_in[19:16];
    66: op1_00_in00 = imem05_in[19:16];
    57: op1_00_in00 = imem07_in[111:108];
    59: op1_00_in00 = imem04_in[47:44];
    83: op1_00_in00 = imem04_in[47:44];
    61: op1_00_in00 = imem06_in[35:32];
    89: op1_00_in00 = imem06_in[35:32];
    62: op1_00_in00 = imem00_in[91:88];
    63: op1_00_in00 = imem02_in[7:4];
    64: op1_00_in00 = imem04_in[127:124];
    65: op1_00_in00 = imem05_in[83:80];
    68: op1_00_in00 = imem05_in[47:44];
    69: op1_00_in00 = imem01_in[31:28];
    70: op1_00_in00 = imem03_in[103:100];
    73: op1_00_in00 = imem05_in[59:56];
    74: op1_00_in00 = imem05_in[111:108];
    80: op1_00_in00 = imem05_in[111:108];
    75: op1_00_in00 = imem07_in[43:40];
    76: op1_00_in00 = imem00_in[75:72];
    78: op1_00_in00 = imem03_in[11:8];
    90: op1_00_in00 = imem03_in[11:8];
    79: op1_00_in00 = imem05_in[71:68];
    81: op1_00_in00 = imem07_in[47:44];
    82: op1_00_in00 = imem07_in[35:32];
    84: op1_00_in00 = imem02_in[75:72];
    85: op1_00_in00 = imem02_in[55:52];
    86: op1_00_in00 = imem06_in[75:72];
    87: op1_00_in00 = imem05_in[115:112];
    88: op1_00_in00 = imem03_in[47:44];
    91: op1_00_in00 = imem05_in[123:120];
    92: op1_00_in00 = imem06_in[3:0];
    93: op1_00_in00 = imem01_in[95:92];
    94: op1_00_in00 = imem01_in[27:24];
    95: op1_00_in00 = imem01_in[67:64];
    96: op1_00_in00 = imem00_in[79:76];
    97: op1_00_in00 = imem00_in[15:12];
    default: op1_00_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv00 = 1;
    10: op1_00_inv00 = 1;
    11: op1_00_inv00 = 1;
    14: op1_00_inv00 = 1;
    15: op1_00_inv00 = 1;
    16: op1_00_inv00 = 1;
    17: op1_00_inv00 = 1;
    18: op1_00_inv00 = 1;
    19: op1_00_inv00 = 1;
    20: op1_00_inv00 = 1;
    21: op1_00_inv00 = 1;
    22: op1_00_inv00 = 1;
    25: op1_00_inv00 = 1;
    27: op1_00_inv00 = 1;
    28: op1_00_inv00 = 1;
    29: op1_00_inv00 = 1;
    33: op1_00_inv00 = 1;
    35: op1_00_inv00 = 1;
    40: op1_00_inv00 = 1;
    42: op1_00_inv00 = 1;
    43: op1_00_inv00 = 1;
    44: op1_00_inv00 = 1;
    47: op1_00_inv00 = 1;
    49: op1_00_inv00 = 1;
    50: op1_00_inv00 = 1;
    54: op1_00_inv00 = 1;
    56: op1_00_inv00 = 1;
    57: op1_00_inv00 = 1;
    59: op1_00_inv00 = 1;
    60: op1_00_inv00 = 1;
    61: op1_00_inv00 = 1;
    62: op1_00_inv00 = 1;
    63: op1_00_inv00 = 1;
    64: op1_00_inv00 = 1;
    65: op1_00_inv00 = 1;
    67: op1_00_inv00 = 1;
    69: op1_00_inv00 = 1;
    70: op1_00_inv00 = 1;
    73: op1_00_inv00 = 1;
    74: op1_00_inv00 = 1;
    75: op1_00_inv00 = 1;
    77: op1_00_inv00 = 1;
    78: op1_00_inv00 = 1;
    83: op1_00_inv00 = 1;
    87: op1_00_inv00 = 1;
    88: op1_00_inv00 = 1;
    90: op1_00_inv00 = 1;
    92: op1_00_inv00 = 1;
    94: op1_00_inv00 = 1;
    95: op1_00_inv00 = 1;
    default: op1_00_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in01 = imem00_in[111:108];
    23: op1_00_in01 = imem00_in[111:108];
    33: op1_00_in01 = imem00_in[111:108];
    76: op1_00_in01 = imem00_in[111:108];
    3: op1_00_in01 = reg_0181;
    6: op1_00_in01 = imem04_in[67:64];
    4: op1_00_in01 = reg_0441;
    7: op1_00_in01 = imem00_in[27:24];
    38: op1_00_in01 = imem00_in[27:24];
    8: op1_00_in01 = imem04_in[115:112];
    9: op1_00_in01 = imem07_in[27:24];
    10: op1_00_in01 = imem01_in[111:108];
    53: op1_00_in01 = imem01_in[111:108];
    11: op1_00_in01 = imem01_in[95:92];
    25: op1_00_in01 = imem01_in[95:92];
    95: op1_00_in01 = imem01_in[95:92];
    12: op1_00_in01 = imem05_in[119:116];
    13: op1_00_in01 = imem00_in[39:36];
    15: op1_00_in01 = imem00_in[39:36];
    30: op1_00_in01 = imem00_in[39:36];
    97: op1_00_in01 = imem00_in[39:36];
    14: op1_00_in01 = imem05_in[111:108];
    16: op1_00_in01 = imem00_in[107:104];
    62: op1_00_in01 = imem00_in[107:104];
    17: op1_00_in01 = imem03_in[103:100];
    18: op1_00_in01 = imem05_in[47:44];
    19: op1_00_in01 = imem04_in[51:48];
    59: op1_00_in01 = imem04_in[51:48];
    20: op1_00_in01 = imem05_in[87:84];
    79: op1_00_in01 = imem05_in[87:84];
    21: op1_00_in01 = imem02_in[19:16];
    22: op1_00_in01 = imem06_in[99:96];
    24: op1_00_in01 = reg_0763;
    26: op1_00_in01 = reg_0758;
    27: op1_00_in01 = imem00_in[31:28];
    28: op1_00_in01 = reg_0982;
    29: op1_00_in01 = imem06_in[19:16];
    31: op1_00_in01 = imem03_in[115:112];
    55: op1_00_in01 = imem03_in[115:112];
    32: op1_00_in01 = imem06_in[83:80];
    34: op1_00_in01 = imem00_in[75:72];
    35: op1_00_in01 = reg_0629;
    36: op1_00_in01 = imem06_in[107:104];
    37: op1_00_in01 = imem06_in[111:108];
    39: op1_00_in01 = imem00_in[23:20];
    40: op1_00_in01 = reg_0102;
    41: op1_00_in01 = imem01_in[87:84];
    42: op1_00_in01 = reg_0283;
    43: op1_00_in01 = imem07_in[119:116];
    44: op1_00_in01 = imem00_in[63:60];
    45: op1_00_in01 = imem02_in[79:76];
    46: op1_00_in01 = imem04_in[39:36];
    47: op1_00_in01 = imem00_in[43:40];
    48: op1_00_in01 = imem01_in[75:72];
    49: op1_00_in01 = imem04_in[83:80];
    50: op1_00_in01 = imem05_in[107:104];
    51: op1_00_in01 = reg_0530;
    52: op1_00_in01 = imem02_in[43:40];
    54: op1_00_in01 = imem03_in[59:56];
    90: op1_00_in01 = imem03_in[59:56];
    56: op1_00_in01 = imem05_in[31:28];
    57: op1_00_in01 = imem07_in[115:112];
    58: op1_00_in01 = imem06_in[103:100];
    61: op1_00_in01 = imem06_in[103:100];
    60: op1_00_in01 = imem00_in[51:48];
    77: op1_00_in01 = imem00_in[51:48];
    63: op1_00_in01 = imem02_in[47:44];
    64: op1_00_in01 = reg_0306;
    65: op1_00_in01 = imem05_in[99:96];
    66: op1_00_in01 = imem05_in[43:40];
    67: op1_00_in01 = imem06_in[51:48];
    68: op1_00_in01 = imem05_in[55:52];
    69: op1_00_in01 = imem01_in[43:40];
    70: op1_00_in01 = reg_0987;
    71: op1_00_in01 = imem06_in[95:92];
    72: op1_00_in01 = imem02_in[71:68];
    73: op1_00_in01 = imem05_in[91:88];
    74: op1_00_in01 = imem06_in[43:40];
    75: op1_00_in01 = imem07_in[55:52];
    78: op1_00_in01 = imem03_in[19:16];
    80: op1_00_in01 = reg_0492;
    81: op1_00_in01 = imem07_in[51:48];
    82: op1_00_in01 = imem07_in[59:56];
    83: op1_00_in01 = imem04_in[55:52];
    84: op1_00_in01 = imem02_in[99:96];
    85: op1_00_in01 = imem02_in[91:88];
    86: op1_00_in01 = imem06_in[79:76];
    87: op1_00_in01 = reg_0707;
    88: op1_00_in01 = imem03_in[123:120];
    89: op1_00_in01 = imem06_in[55:52];
    91: op1_00_in01 = reg_0143;
    92: op1_00_in01 = imem06_in[7:4];
    93: op1_00_in01 = imem01_in[115:112];
    94: op1_00_in01 = imem01_in[31:28];
    96: op1_00_in01 = reg_0683;
    default: op1_00_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv01 = 1;
    7: op1_00_inv01 = 1;
    9: op1_00_inv01 = 1;
    10: op1_00_inv01 = 1;
    13: op1_00_inv01 = 1;
    15: op1_00_inv01 = 1;
    18: op1_00_inv01 = 1;
    24: op1_00_inv01 = 1;
    26: op1_00_inv01 = 1;
    27: op1_00_inv01 = 1;
    30: op1_00_inv01 = 1;
    31: op1_00_inv01 = 1;
    32: op1_00_inv01 = 1;
    34: op1_00_inv01 = 1;
    37: op1_00_inv01 = 1;
    38: op1_00_inv01 = 1;
    39: op1_00_inv01 = 1;
    40: op1_00_inv01 = 1;
    41: op1_00_inv01 = 1;
    44: op1_00_inv01 = 1;
    45: op1_00_inv01 = 1;
    46: op1_00_inv01 = 1;
    47: op1_00_inv01 = 1;
    49: op1_00_inv01 = 1;
    50: op1_00_inv01 = 1;
    52: op1_00_inv01 = 1;
    58: op1_00_inv01 = 1;
    59: op1_00_inv01 = 1;
    61: op1_00_inv01 = 1;
    65: op1_00_inv01 = 1;
    67: op1_00_inv01 = 1;
    71: op1_00_inv01 = 1;
    72: op1_00_inv01 = 1;
    73: op1_00_inv01 = 1;
    74: op1_00_inv01 = 1;
    75: op1_00_inv01 = 1;
    76: op1_00_inv01 = 1;
    77: op1_00_inv01 = 1;
    79: op1_00_inv01 = 1;
    80: op1_00_inv01 = 1;
    81: op1_00_inv01 = 1;
    82: op1_00_inv01 = 1;
    83: op1_00_inv01 = 1;
    85: op1_00_inv01 = 1;
    87: op1_00_inv01 = 1;
    88: op1_00_inv01 = 1;
    90: op1_00_inv01 = 1;
    92: op1_00_inv01 = 1;
    93: op1_00_inv01 = 1;
    94: op1_00_inv01 = 1;
    95: op1_00_inv01 = 1;
    96: op1_00_inv01 = 1;
    default: op1_00_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in02 = imem00_in[115:112];
    16: op1_00_in02 = imem00_in[115:112];
    3: op1_00_in02 = reg_0169;
    6: op1_00_in02 = imem04_in[103:100];
    19: op1_00_in02 = imem04_in[103:100];
    4: op1_00_in02 = reg_0428;
    7: op1_00_in02 = imem00_in[63:60];
    8: op1_00_in02 = reg_0545;
    9: op1_00_in02 = imem07_in[95:92];
    10: op1_00_in02 = imem01_in[115:112];
    25: op1_00_in02 = imem01_in[115:112];
    41: op1_00_in02 = imem01_in[115:112];
    11: op1_00_in02 = reg_0905;
    12: op1_00_in02 = reg_0132;
    13: op1_00_in02 = imem00_in[59:56];
    30: op1_00_in02 = imem00_in[59:56];
    14: op1_00_in02 = reg_0973;
    15: op1_00_in02 = imem00_in[47:44];
    97: op1_00_in02 = imem00_in[47:44];
    17: op1_00_in02 = imem03_in[119:116];
    55: op1_00_in02 = imem03_in[119:116];
    18: op1_00_in02 = imem05_in[59:56];
    20: op1_00_in02 = reg_0147;
    21: op1_00_in02 = imem02_in[75:72];
    72: op1_00_in02 = imem02_in[75:72];
    22: op1_00_in02 = imem06_in[103:100];
    23: op1_00_in02 = reg_0684;
    24: op1_00_in02 = reg_0882;
    26: op1_00_in02 = reg_0506;
    27: op1_00_in02 = imem00_in[55:52];
    47: op1_00_in02 = imem00_in[55:52];
    28: op1_00_in02 = reg_0984;
    29: op1_00_in02 = imem06_in[23:20];
    92: op1_00_in02 = imem06_in[23:20];
    31: op1_00_in02 = reg_0377;
    32: op1_00_in02 = imem07_in[3:0];
    33: op1_00_in02 = reg_0689;
    34: op1_00_in02 = imem00_in[79:76];
    35: op1_00_in02 = reg_0630;
    36: op1_00_in02 = reg_0348;
    37: op1_00_in02 = imem06_in[115:112];
    38: op1_00_in02 = imem00_in[31:28];
    39: op1_00_in02 = imem00_in[91:88];
    40: op1_00_in02 = reg_0114;
    42: op1_00_in02 = reg_0736;
    43: op1_00_in02 = reg_0179;
    44: op1_00_in02 = imem00_in[67:64];
    77: op1_00_in02 = imem00_in[67:64];
    45: op1_00_in02 = imem02_in[87:84];
    46: op1_00_in02 = imem04_in[67:64];
    48: op1_00_in02 = imem01_in[95:92];
    49: op1_00_in02 = imem04_in[87:84];
    50: op1_00_in02 = imem05_in[115:112];
    51: op1_00_in02 = reg_0511;
    52: op1_00_in02 = imem02_in[59:56];
    53: op1_00_in02 = imem02_in[35:32];
    54: op1_00_in02 = imem03_in[71:68];
    56: op1_00_in02 = imem05_in[71:68];
    57: op1_00_in02 = reg_0721;
    58: op1_00_in02 = imem06_in[127:124];
    59: op1_00_in02 = imem04_in[55:52];
    60: op1_00_in02 = imem00_in[95:92];
    61: op1_00_in02 = imem07_in[19:16];
    62: op1_00_in02 = imem00_in[119:116];
    63: op1_00_in02 = imem02_in[83:80];
    64: op1_00_in02 = reg_1057;
    65: op1_00_in02 = imem05_in[111:108];
    66: op1_00_in02 = imem05_in[83:80];
    67: op1_00_in02 = imem06_in[55:52];
    68: op1_00_in02 = imem05_in[87:84];
    69: op1_00_in02 = imem01_in[91:88];
    70: op1_00_in02 = reg_1002;
    71: op1_00_in02 = imem06_in[99:96];
    73: op1_00_in02 = imem05_in[107:104];
    74: op1_00_in02 = imem06_in[59:56];
    75: op1_00_in02 = reg_0250;
    76: op1_00_in02 = reg_0683;
    78: op1_00_in02 = imem03_in[23:20];
    79: op1_00_in02 = imem05_in[119:116];
    80: op1_00_in02 = reg_0217;
    81: op1_00_in02 = imem07_in[59:56];
    82: op1_00_in02 = imem07_in[63:60];
    83: op1_00_in02 = imem04_in[123:120];
    84: op1_00_in02 = imem02_in[111:108];
    85: op1_00_in02 = imem03_in[43:40];
    86: op1_00_in02 = reg_0857;
    87: op1_00_in02 = reg_0780;
    88: op1_00_in02 = reg_0672;
    89: op1_00_in02 = imem06_in[79:76];
    90: op1_00_in02 = imem03_in[63:60];
    91: op1_00_in02 = reg_0275;
    93: op1_00_in02 = reg_0832;
    94: op1_00_in02 = imem01_in[55:52];
    95: op1_00_in02 = imem01_in[111:108];
    96: op1_00_in02 = reg_0223;
    default: op1_00_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv02 = 1;
    6: op1_00_inv02 = 1;
    7: op1_00_inv02 = 1;
    9: op1_00_inv02 = 1;
    11: op1_00_inv02 = 1;
    12: op1_00_inv02 = 1;
    13: op1_00_inv02 = 1;
    17: op1_00_inv02 = 1;
    19: op1_00_inv02 = 1;
    20: op1_00_inv02 = 1;
    22: op1_00_inv02 = 1;
    24: op1_00_inv02 = 1;
    25: op1_00_inv02 = 1;
    27: op1_00_inv02 = 1;
    28: op1_00_inv02 = 1;
    29: op1_00_inv02 = 1;
    32: op1_00_inv02 = 1;
    33: op1_00_inv02 = 1;
    35: op1_00_inv02 = 1;
    36: op1_00_inv02 = 1;
    37: op1_00_inv02 = 1;
    39: op1_00_inv02 = 1;
    42: op1_00_inv02 = 1;
    45: op1_00_inv02 = 1;
    46: op1_00_inv02 = 1;
    51: op1_00_inv02 = 1;
    53: op1_00_inv02 = 1;
    54: op1_00_inv02 = 1;
    56: op1_00_inv02 = 1;
    57: op1_00_inv02 = 1;
    58: op1_00_inv02 = 1;
    59: op1_00_inv02 = 1;
    60: op1_00_inv02 = 1;
    63: op1_00_inv02 = 1;
    64: op1_00_inv02 = 1;
    67: op1_00_inv02 = 1;
    68: op1_00_inv02 = 1;
    69: op1_00_inv02 = 1;
    70: op1_00_inv02 = 1;
    71: op1_00_inv02 = 1;
    72: op1_00_inv02 = 1;
    74: op1_00_inv02 = 1;
    75: op1_00_inv02 = 1;
    78: op1_00_inv02 = 1;
    80: op1_00_inv02 = 1;
    83: op1_00_inv02 = 1;
    90: op1_00_inv02 = 1;
    92: op1_00_inv02 = 1;
    96: op1_00_inv02 = 1;
    97: op1_00_inv02 = 1;
    default: op1_00_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in03 = reg_0683;
    3: op1_00_in03 = reg_0160;
    6: op1_00_in03 = imem04_in[107:104];
    19: op1_00_in03 = imem04_in[107:104];
    4: op1_00_in03 = reg_0442;
    7: op1_00_in03 = imem00_in[95:92];
    39: op1_00_in03 = imem00_in[95:92];
    8: op1_00_in03 = reg_0557;
    9: op1_00_in03 = imem07_in[107:104];
    10: op1_00_in03 = imem01_in[119:116];
    11: op1_00_in03 = reg_1040;
    12: op1_00_in03 = reg_0146;
    13: op1_00_in03 = imem00_in[67:64];
    14: op1_00_in03 = reg_0954;
    15: op1_00_in03 = imem00_in[51:48];
    38: op1_00_in03 = imem00_in[51:48];
    16: op1_00_in03 = reg_0694;
    17: op1_00_in03 = reg_0573;
    18: op1_00_in03 = imem05_in[99:96];
    20: op1_00_in03 = reg_0148;
    21: op1_00_in03 = imem02_in[87:84];
    22: op1_00_in03 = imem06_in[111:108];
    23: op1_00_in03 = reg_0670;
    24: op1_00_in03 = reg_0015;
    25: op1_00_in03 = reg_1033;
    26: op1_00_in03 = reg_0016;
    27: op1_00_in03 = imem00_in[91:88];
    28: op1_00_in03 = reg_0993;
    29: op1_00_in03 = imem06_in[55:52];
    30: op1_00_in03 = imem00_in[71:68];
    31: op1_00_in03 = reg_0836;
    32: op1_00_in03 = imem07_in[23:20];
    33: op1_00_in03 = reg_0679;
    34: op1_00_in03 = imem00_in[83:80];
    35: op1_00_in03 = reg_0633;
    36: op1_00_in03 = reg_0381;
    37: op1_00_in03 = imem07_in[3:0];
    71: op1_00_in03 = imem07_in[3:0];
    40: op1_00_in03 = reg_0107;
    41: op1_00_in03 = reg_0123;
    42: op1_00_in03 = reg_0043;
    43: op1_00_in03 = reg_0169;
    44: op1_00_in03 = imem00_in[119:116];
    45: op1_00_in03 = imem02_in[119:116];
    46: op1_00_in03 = imem05_in[3:0];
    47: op1_00_in03 = imem00_in[59:56];
    48: op1_00_in03 = imem01_in[99:96];
    49: op1_00_in03 = imem04_in[111:108];
    50: op1_00_in03 = reg_0145;
    51: op1_00_in03 = reg_0265;
    52: op1_00_in03 = imem02_in[95:92];
    63: op1_00_in03 = imem02_in[95:92];
    53: op1_00_in03 = imem02_in[43:40];
    54: op1_00_in03 = imem03_in[87:84];
    90: op1_00_in03 = imem03_in[87:84];
    55: op1_00_in03 = reg_0847;
    56: op1_00_in03 = imem05_in[91:88];
    57: op1_00_in03 = reg_0713;
    58: op1_00_in03 = reg_1029;
    59: op1_00_in03 = imem04_in[59:56];
    60: op1_00_in03 = imem00_in[123:120];
    61: op1_00_in03 = imem07_in[27:24];
    62: op1_00_in03 = imem00_in[127:124];
    64: op1_00_in03 = reg_0850;
    65: op1_00_in03 = reg_0063;
    66: op1_00_in03 = imem05_in[119:116];
    67: op1_00_in03 = imem06_in[67:64];
    68: op1_00_in03 = imem05_in[95:92];
    69: op1_00_in03 = reg_0607;
    70: op1_00_in03 = reg_0992;
    72: op1_00_in03 = reg_0644;
    73: op1_00_in03 = reg_0020;
    74: op1_00_in03 = imem06_in[63:60];
    75: op1_00_in03 = reg_0433;
    76: op1_00_in03 = reg_0843;
    77: op1_00_in03 = imem00_in[75:72];
    78: op1_00_in03 = imem03_in[67:64];
    79: op1_00_in03 = imem05_in[123:120];
    80: op1_00_in03 = reg_0652;
    81: op1_00_in03 = imem07_in[79:76];
    82: op1_00_in03 = imem07_in[115:112];
    83: op1_00_in03 = reg_0848;
    84: op1_00_in03 = reg_0323;
    85: op1_00_in03 = reg_0322;
    86: op1_00_in03 = reg_0032;
    87: op1_00_in03 = reg_0528;
    88: op1_00_in03 = reg_0581;
    89: op1_00_in03 = imem06_in[83:80];
    91: op1_00_in03 = reg_0269;
    92: op1_00_in03 = reg_0391;
    93: op1_00_in03 = reg_1055;
    94: op1_00_in03 = imem01_in[63:60];
    95: op1_00_in03 = reg_0769;
    96: op1_00_in03 = reg_0118;
    97: op1_00_in03 = imem00_in[99:96];
    default: op1_00_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    3: op1_00_inv03 = 1;
    6: op1_00_inv03 = 1;
    4: op1_00_inv03 = 1;
    7: op1_00_inv03 = 1;
    8: op1_00_inv03 = 1;
    10: op1_00_inv03 = 1;
    11: op1_00_inv03 = 1;
    12: op1_00_inv03 = 1;
    15: op1_00_inv03 = 1;
    18: op1_00_inv03 = 1;
    21: op1_00_inv03 = 1;
    23: op1_00_inv03 = 1;
    25: op1_00_inv03 = 1;
    26: op1_00_inv03 = 1;
    28: op1_00_inv03 = 1;
    34: op1_00_inv03 = 1;
    36: op1_00_inv03 = 1;
    38: op1_00_inv03 = 1;
    40: op1_00_inv03 = 1;
    42: op1_00_inv03 = 1;
    43: op1_00_inv03 = 1;
    46: op1_00_inv03 = 1;
    49: op1_00_inv03 = 1;
    51: op1_00_inv03 = 1;
    53: op1_00_inv03 = 1;
    55: op1_00_inv03 = 1;
    62: op1_00_inv03 = 1;
    64: op1_00_inv03 = 1;
    65: op1_00_inv03 = 1;
    69: op1_00_inv03 = 1;
    70: op1_00_inv03 = 1;
    75: op1_00_inv03 = 1;
    76: op1_00_inv03 = 1;
    77: op1_00_inv03 = 1;
    80: op1_00_inv03 = 1;
    84: op1_00_inv03 = 1;
    89: op1_00_inv03 = 1;
    91: op1_00_inv03 = 1;
    94: op1_00_inv03 = 1;
    95: op1_00_inv03 = 1;
    97: op1_00_inv03 = 1;
    default: op1_00_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in04 = reg_0684;
    6: op1_00_in04 = reg_0545;
    4: op1_00_in04 = reg_0443;
    7: op1_00_in04 = imem00_in[107:104];
    30: op1_00_in04 = imem00_in[107:104];
    8: op1_00_in04 = reg_0530;
    9: op1_00_in04 = imem07_in[115:112];
    10: op1_00_in04 = reg_0123;
    11: op1_00_in04 = reg_1035;
    25: op1_00_in04 = reg_1035;
    12: op1_00_in04 = reg_0155;
    13: op1_00_in04 = imem00_in[87:84];
    47: op1_00_in04 = imem00_in[87:84];
    14: op1_00_in04 = reg_0964;
    15: op1_00_in04 = imem00_in[59:56];
    16: op1_00_in04 = reg_0677;
    17: op1_00_in04 = reg_0596;
    18: op1_00_in04 = imem05_in[123:120];
    19: op1_00_in04 = reg_0058;
    20: op1_00_in04 = reg_0153;
    21: op1_00_in04 = imem03_in[27:24];
    22: op1_00_in04 = imem06_in[123:120];
    23: op1_00_in04 = reg_0680;
    24: op1_00_in04 = reg_0278;
    26: op1_00_in04 = reg_0872;
    27: op1_00_in04 = imem00_in[103:100];
    38: op1_00_in04 = imem00_in[103:100];
    28: op1_00_in04 = reg_0980;
    29: op1_00_in04 = reg_0787;
    31: op1_00_in04 = reg_0312;
    32: op1_00_in04 = imem07_in[39:36];
    33: op1_00_in04 = reg_0678;
    34: op1_00_in04 = imem00_in[127:124];
    35: op1_00_in04 = reg_0632;
    36: op1_00_in04 = reg_0393;
    37: op1_00_in04 = imem07_in[15:12];
    39: op1_00_in04 = reg_0683;
    40: op1_00_in04 = imem02_in[47:44];
    41: op1_00_in04 = reg_0103;
    42: op1_00_in04 = reg_0854;
    43: op1_00_in04 = reg_0185;
    44: op1_00_in04 = reg_0681;
    45: op1_00_in04 = reg_0080;
    46: op1_00_in04 = imem05_in[11:8];
    48: op1_00_in04 = reg_0522;
    49: op1_00_in04 = imem05_in[15:12];
    50: op1_00_in04 = reg_0129;
    51: op1_00_in04 = reg_0937;
    52: op1_00_in04 = imem02_in[107:104];
    53: op1_00_in04 = imem02_in[51:48];
    54: op1_00_in04 = imem03_in[91:88];
    55: op1_00_in04 = reg_0836;
    56: op1_00_in04 = reg_0019;
    57: op1_00_in04 = reg_0707;
    58: op1_00_in04 = reg_0241;
    59: op1_00_in04 = imem05_in[3:0];
    60: op1_00_in04 = reg_0768;
    62: op1_00_in04 = reg_0768;
    61: op1_00_in04 = imem07_in[59:56];
    63: op1_00_in04 = imem02_in[119:116];
    64: op1_00_in04 = reg_0066;
    65: op1_00_in04 = reg_0826;
    66: op1_00_in04 = imem05_in[127:124];
    67: op1_00_in04 = imem06_in[83:80];
    74: op1_00_in04 = imem06_in[83:80];
    68: op1_00_in04 = imem05_in[107:104];
    69: op1_00_in04 = reg_0500;
    70: op1_00_in04 = reg_1001;
    71: op1_00_in04 = imem07_in[11:8];
    72: op1_00_in04 = reg_0089;
    73: op1_00_in04 = reg_0125;
    75: op1_00_in04 = reg_0744;
    76: op1_00_in04 = reg_0738;
    77: op1_00_in04 = imem00_in[115:112];
    78: op1_00_in04 = imem03_in[99:96];
    90: op1_00_in04 = imem03_in[99:96];
    79: op1_00_in04 = reg_0135;
    80: op1_00_in04 = reg_0319;
    81: op1_00_in04 = imem07_in[83:80];
    83: op1_00_in04 = reg_0850;
    84: op1_00_in04 = reg_0441;
    85: op1_00_in04 = reg_0298;
    86: op1_00_in04 = reg_0835;
    87: op1_00_in04 = reg_0816;
    88: op1_00_in04 = reg_0385;
    89: op1_00_in04 = imem07_in[7:4];
    91: op1_00_in04 = reg_0583;
    92: op1_00_in04 = reg_0926;
    93: op1_00_in04 = reg_1033;
    95: op1_00_in04 = reg_1033;
    94: op1_00_in04 = reg_0097;
    96: op1_00_in04 = reg_0867;
    97: op1_00_in04 = imem00_in[123:120];
    default: op1_00_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv04 = 1;
    6: op1_00_inv04 = 1;
    8: op1_00_inv04 = 1;
    9: op1_00_inv04 = 1;
    10: op1_00_inv04 = 1;
    11: op1_00_inv04 = 1;
    13: op1_00_inv04 = 1;
    15: op1_00_inv04 = 1;
    16: op1_00_inv04 = 1;
    17: op1_00_inv04 = 1;
    18: op1_00_inv04 = 1;
    20: op1_00_inv04 = 1;
    22: op1_00_inv04 = 1;
    25: op1_00_inv04 = 1;
    26: op1_00_inv04 = 1;
    30: op1_00_inv04 = 1;
    31: op1_00_inv04 = 1;
    32: op1_00_inv04 = 1;
    34: op1_00_inv04 = 1;
    38: op1_00_inv04 = 1;
    39: op1_00_inv04 = 1;
    40: op1_00_inv04 = 1;
    41: op1_00_inv04 = 1;
    43: op1_00_inv04 = 1;
    44: op1_00_inv04 = 1;
    46: op1_00_inv04 = 1;
    47: op1_00_inv04 = 1;
    49: op1_00_inv04 = 1;
    50: op1_00_inv04 = 1;
    51: op1_00_inv04 = 1;
    52: op1_00_inv04 = 1;
    54: op1_00_inv04 = 1;
    55: op1_00_inv04 = 1;
    58: op1_00_inv04 = 1;
    59: op1_00_inv04 = 1;
    60: op1_00_inv04 = 1;
    61: op1_00_inv04 = 1;
    62: op1_00_inv04 = 1;
    64: op1_00_inv04 = 1;
    68: op1_00_inv04 = 1;
    70: op1_00_inv04 = 1;
    71: op1_00_inv04 = 1;
    72: op1_00_inv04 = 1;
    74: op1_00_inv04 = 1;
    76: op1_00_inv04 = 1;
    77: op1_00_inv04 = 1;
    86: op1_00_inv04 = 1;
    87: op1_00_inv04 = 1;
    88: op1_00_inv04 = 1;
    96: op1_00_inv04 = 1;
    default: op1_00_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in05 = reg_0679;
    6: op1_00_in05 = reg_0551;
    4: op1_00_in05 = reg_0172;
    7: op1_00_in05 = imem00_in[123:120];
    8: op1_00_in05 = reg_0550;
    9: op1_00_in05 = reg_0722;
    10: op1_00_in05 = reg_0124;
    11: op1_00_in05 = reg_0913;
    25: op1_00_in05 = reg_0913;
    12: op1_00_in05 = imem06_in[3:0];
    13: op1_00_in05 = reg_0697;
    14: op1_00_in05 = reg_0942;
    15: op1_00_in05 = imem00_in[63:60];
    16: op1_00_in05 = reg_0678;
    17: op1_00_in05 = reg_0583;
    18: op1_00_in05 = reg_0962;
    19: op1_00_in05 = reg_0044;
    20: op1_00_in05 = reg_0134;
    21: op1_00_in05 = imem03_in[43:40];
    22: op1_00_in05 = reg_0604;
    23: op1_00_in05 = reg_0477;
    24: op1_00_in05 = reg_0047;
    26: op1_00_in05 = imem03_in[35:32];
    27: op1_00_in05 = reg_0684;
    28: op1_00_in05 = reg_0977;
    29: op1_00_in05 = reg_0025;
    30: op1_00_in05 = reg_0685;
    34: op1_00_in05 = reg_0685;
    44: op1_00_in05 = reg_0685;
    60: op1_00_in05 = reg_0685;
    31: op1_00_in05 = reg_0820;
    32: op1_00_in05 = imem07_in[43:40];
    33: op1_00_in05 = reg_0688;
    35: op1_00_in05 = reg_0623;
    36: op1_00_in05 = reg_0741;
    37: op1_00_in05 = imem07_in[59:56];
    38: op1_00_in05 = reg_0682;
    39: op1_00_in05 = reg_0681;
    40: op1_00_in05 = imem02_in[51:48];
    41: op1_00_in05 = reg_0118;
    42: op1_00_in05 = imem05_in[15:12];
    43: op1_00_in05 = reg_0173;
    45: op1_00_in05 = reg_0096;
    46: op1_00_in05 = imem05_in[27:24];
    47: op1_00_in05 = imem00_in[119:116];
    48: op1_00_in05 = reg_0829;
    49: op1_00_in05 = imem05_in[19:16];
    50: op1_00_in05 = imem06_in[59:56];
    51: op1_00_in05 = reg_0282;
    52: op1_00_in05 = imem02_in[115:112];
    53: op1_00_in05 = imem02_in[83:80];
    54: op1_00_in05 = imem03_in[103:100];
    78: op1_00_in05 = imem03_in[103:100];
    55: op1_00_in05 = reg_0376;
    56: op1_00_in05 = reg_0757;
    57: op1_00_in05 = reg_0641;
    58: op1_00_in05 = reg_0605;
    59: op1_00_in05 = imem05_in[91:88];
    61: op1_00_in05 = imem07_in[67:64];
    89: op1_00_in05 = imem07_in[67:64];
    62: op1_00_in05 = reg_0686;
    63: op1_00_in05 = imem02_in[127:124];
    64: op1_00_in05 = reg_0076;
    65: op1_00_in05 = reg_0032;
    66: op1_00_in05 = reg_0147;
    67: op1_00_in05 = imem06_in[87:84];
    68: op1_00_in05 = imem05_in[115:112];
    69: op1_00_in05 = reg_0521;
    70: op1_00_in05 = reg_0993;
    71: op1_00_in05 = imem07_in[91:88];
    72: op1_00_in05 = reg_0484;
    73: op1_00_in05 = reg_0784;
    74: op1_00_in05 = imem06_in[95:92];
    75: op1_00_in05 = reg_0353;
    76: op1_00_in05 = reg_0669;
    77: op1_00_in05 = reg_0768;
    79: op1_00_in05 = reg_0706;
    80: op1_00_in05 = reg_0655;
    83: op1_00_in05 = reg_0058;
    84: op1_00_in05 = reg_0359;
    85: op1_00_in05 = reg_0661;
    86: op1_00_in05 = reg_0915;
    87: op1_00_in05 = reg_0326;
    88: op1_00_in05 = reg_0266;
    90: op1_00_in05 = imem03_in[115:112];
    91: op1_00_in05 = reg_0436;
    92: op1_00_in05 = reg_0533;
    93: op1_00_in05 = reg_0273;
    94: op1_00_in05 = reg_0933;
    95: op1_00_in05 = reg_0555;
    96: op1_00_in05 = reg_0762;
    97: op1_00_in05 = reg_0857;
    default: op1_00_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv05 = 1;
    7: op1_00_inv05 = 1;
    9: op1_00_inv05 = 1;
    11: op1_00_inv05 = 1;
    12: op1_00_inv05 = 1;
    14: op1_00_inv05 = 1;
    15: op1_00_inv05 = 1;
    16: op1_00_inv05 = 1;
    17: op1_00_inv05 = 1;
    18: op1_00_inv05 = 1;
    25: op1_00_inv05 = 1;
    32: op1_00_inv05 = 1;
    33: op1_00_inv05 = 1;
    36: op1_00_inv05 = 1;
    43: op1_00_inv05 = 1;
    47: op1_00_inv05 = 1;
    48: op1_00_inv05 = 1;
    49: op1_00_inv05 = 1;
    52: op1_00_inv05 = 1;
    55: op1_00_inv05 = 1;
    56: op1_00_inv05 = 1;
    57: op1_00_inv05 = 1;
    60: op1_00_inv05 = 1;
    65: op1_00_inv05 = 1;
    67: op1_00_inv05 = 1;
    68: op1_00_inv05 = 1;
    69: op1_00_inv05 = 1;
    70: op1_00_inv05 = 1;
    71: op1_00_inv05 = 1;
    74: op1_00_inv05 = 1;
    75: op1_00_inv05 = 1;
    76: op1_00_inv05 = 1;
    77: op1_00_inv05 = 1;
    80: op1_00_inv05 = 1;
    84: op1_00_inv05 = 1;
    88: op1_00_inv05 = 1;
    89: op1_00_inv05 = 1;
    92: op1_00_inv05 = 1;
    default: op1_00_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in06 = reg_0668;
    6: op1_00_in06 = reg_0281;
    4: op1_00_in06 = reg_0157;
    7: op1_00_in06 = reg_0689;
    8: op1_00_in06 = reg_0548;
    9: op1_00_in06 = reg_0709;
    10: op1_00_in06 = reg_0103;
    11: op1_00_in06 = reg_0871;
    25: op1_00_in06 = reg_0871;
    12: op1_00_in06 = imem06_in[115:112];
    13: op1_00_in06 = reg_0451;
    14: op1_00_in06 = reg_0952;
    15: op1_00_in06 = imem00_in[83:80];
    16: op1_00_in06 = reg_0673;
    17: op1_00_in06 = reg_0572;
    97: op1_00_in06 = reg_0572;
    18: op1_00_in06 = reg_0963;
    19: op1_00_in06 = imem05_in[87:84];
    46: op1_00_in06 = imem05_in[87:84];
    20: op1_00_in06 = imem06_in[7:4];
    21: op1_00_in06 = imem03_in[55:52];
    22: op1_00_in06 = reg_0609;
    23: op1_00_in06 = reg_0481;
    24: op1_00_in06 = reg_0528;
    26: op1_00_in06 = imem03_in[47:44];
    27: op1_00_in06 = reg_0677;
    28: op1_00_in06 = reg_0976;
    29: op1_00_in06 = reg_1010;
    30: op1_00_in06 = reg_0694;
    31: op1_00_in06 = reg_0996;
    32: op1_00_in06 = imem07_in[51:48];
    33: op1_00_in06 = reg_0463;
    34: op1_00_in06 = reg_0674;
    35: op1_00_in06 = reg_0356;
    36: op1_00_in06 = reg_0383;
    37: op1_00_in06 = imem07_in[91:88];
    38: op1_00_in06 = reg_0697;
    39: op1_00_in06 = reg_0685;
    40: op1_00_in06 = imem02_in[95:92];
    41: op1_00_in06 = reg_0116;
    42: op1_00_in06 = imem05_in[39:36];
    44: op1_00_in06 = reg_0684;
    60: op1_00_in06 = reg_0684;
    45: op1_00_in06 = reg_0098;
    47: op1_00_in06 = reg_0672;
    48: op1_00_in06 = reg_0830;
    49: op1_00_in06 = imem05_in[31:28];
    50: op1_00_in06 = reg_0073;
    51: op1_00_in06 = reg_0055;
    52: op1_00_in06 = reg_0083;
    53: op1_00_in06 = imem02_in[115:112];
    54: op1_00_in06 = reg_0923;
    55: op1_00_in06 = reg_0518;
    56: op1_00_in06 = reg_0094;
    57: op1_00_in06 = reg_0427;
    58: op1_00_in06 = imem07_in[11:8];
    59: op1_00_in06 = imem05_in[95:92];
    61: op1_00_in06 = imem07_in[71:68];
    62: op1_00_in06 = reg_0828;
    63: op1_00_in06 = reg_0739;
    64: op1_00_in06 = reg_0056;
    65: op1_00_in06 = reg_0813;
    66: op1_00_in06 = reg_0136;
    67: op1_00_in06 = imem06_in[95:92];
    68: op1_00_in06 = reg_0583;
    69: op1_00_in06 = reg_0354;
    70: op1_00_in06 = reg_0975;
    71: op1_00_in06 = imem07_in[99:96];
    89: op1_00_in06 = imem07_in[99:96];
    72: op1_00_in06 = imem03_in[43:40];
    73: op1_00_in06 = reg_0004;
    74: op1_00_in06 = reg_0080;
    75: op1_00_in06 = reg_0165;
    76: op1_00_in06 = reg_0465;
    77: op1_00_in06 = reg_0825;
    78: op1_00_in06 = imem03_in[111:108];
    79: op1_00_in06 = reg_0146;
    80: op1_00_in06 = reg_0448;
    83: op1_00_in06 = reg_0076;
    84: op1_00_in06 = reg_0372;
    85: op1_00_in06 = reg_0823;
    86: op1_00_in06 = reg_0022;
    87: op1_00_in06 = reg_0965;
    88: op1_00_in06 = reg_0551;
    90: op1_00_in06 = imem04_in[71:68];
    91: op1_00_in06 = reg_0437;
    92: op1_00_in06 = reg_0264;
    93: op1_00_in06 = reg_0860;
    94: op1_00_in06 = reg_1056;
    95: op1_00_in06 = reg_0101;
    96: op1_00_in06 = reg_0310;
    default: op1_00_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_00_inv06 = 1;
    8: op1_00_inv06 = 1;
    11: op1_00_inv06 = 1;
    13: op1_00_inv06 = 1;
    15: op1_00_inv06 = 1;
    18: op1_00_inv06 = 1;
    19: op1_00_inv06 = 1;
    20: op1_00_inv06 = 1;
    21: op1_00_inv06 = 1;
    25: op1_00_inv06 = 1;
    26: op1_00_inv06 = 1;
    28: op1_00_inv06 = 1;
    31: op1_00_inv06 = 1;
    33: op1_00_inv06 = 1;
    34: op1_00_inv06 = 1;
    38: op1_00_inv06 = 1;
    42: op1_00_inv06 = 1;
    47: op1_00_inv06 = 1;
    48: op1_00_inv06 = 1;
    49: op1_00_inv06 = 1;
    50: op1_00_inv06 = 1;
    52: op1_00_inv06 = 1;
    54: op1_00_inv06 = 1;
    56: op1_00_inv06 = 1;
    57: op1_00_inv06 = 1;
    60: op1_00_inv06 = 1;
    61: op1_00_inv06 = 1;
    63: op1_00_inv06 = 1;
    64: op1_00_inv06 = 1;
    66: op1_00_inv06 = 1;
    69: op1_00_inv06 = 1;
    71: op1_00_inv06 = 1;
    72: op1_00_inv06 = 1;
    74: op1_00_inv06 = 1;
    75: op1_00_inv06 = 1;
    76: op1_00_inv06 = 1;
    77: op1_00_inv06 = 1;
    80: op1_00_inv06 = 1;
    85: op1_00_inv06 = 1;
    86: op1_00_inv06 = 1;
    89: op1_00_inv06 = 1;
    93: op1_00_inv06 = 1;
    94: op1_00_inv06 = 1;
    96: op1_00_inv06 = 1;
    default: op1_00_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in07 = reg_0680;
    27: op1_00_in07 = reg_0680;
    6: op1_00_in07 = reg_0305;
    4: op1_00_in07 = reg_0173;
    7: op1_00_in07 = reg_0677;
    8: op1_00_in07 = reg_0549;
    9: op1_00_in07 = reg_0421;
    10: op1_00_in07 = reg_0116;
    11: op1_00_in07 = reg_1017;
    12: op1_00_in07 = imem06_in[119:116];
    13: op1_00_in07 = reg_0462;
    14: op1_00_in07 = reg_0834;
    15: op1_00_in07 = imem00_in[115:112];
    16: op1_00_in07 = reg_0457;
    17: op1_00_in07 = reg_0593;
    18: op1_00_in07 = reg_0955;
    19: op1_00_in07 = imem05_in[107:104];
    20: op1_00_in07 = imem06_in[23:20];
    21: op1_00_in07 = imem03_in[87:84];
    22: op1_00_in07 = reg_0611;
    23: op1_00_in07 = reg_0480;
    24: op1_00_in07 = reg_0774;
    25: op1_00_in07 = reg_0228;
    26: op1_00_in07 = imem03_in[51:48];
    28: op1_00_in07 = imem04_in[7:4];
    29: op1_00_in07 = reg_0805;
    30: op1_00_in07 = reg_0668;
    31: op1_00_in07 = reg_0978;
    32: op1_00_in07 = imem07_in[71:68];
    33: op1_00_in07 = reg_0454;
    34: op1_00_in07 = reg_0463;
    35: op1_00_in07 = reg_0382;
    36: op1_00_in07 = reg_0804;
    37: op1_00_in07 = imem07_in[111:108];
    38: op1_00_in07 = reg_0690;
    39: op1_00_in07 = reg_0684;
    40: op1_00_in07 = imem02_in[127:124];
    41: op1_00_in07 = reg_0120;
    42: op1_00_in07 = imem05_in[47:44];
    44: op1_00_in07 = reg_0674;
    45: op1_00_in07 = reg_0336;
    46: op1_00_in07 = imem05_in[123:120];
    47: op1_00_in07 = reg_0686;
    60: op1_00_in07 = reg_0686;
    77: op1_00_in07 = reg_0686;
    48: op1_00_in07 = reg_0354;
    49: op1_00_in07 = imem05_in[43:40];
    50: op1_00_in07 = reg_0883;
    51: op1_00_in07 = reg_1020;
    52: op1_00_in07 = reg_0007;
    53: op1_00_in07 = reg_0326;
    54: op1_00_in07 = reg_0543;
    55: op1_00_in07 = reg_0822;
    56: op1_00_in07 = reg_0438;
    57: op1_00_in07 = reg_0024;
    58: op1_00_in07 = imem07_in[35:32];
    59: op1_00_in07 = imem05_in[99:96];
    61: op1_00_in07 = imem07_in[91:88];
    62: op1_00_in07 = reg_0455;
    63: op1_00_in07 = reg_0359;
    64: op1_00_in07 = reg_0276;
    65: op1_00_in07 = reg_0145;
    66: op1_00_in07 = reg_0152;
    67: op1_00_in07 = reg_0660;
    68: op1_00_in07 = reg_0941;
    69: op1_00_in07 = reg_0610;
    94: op1_00_in07 = reg_0610;
    70: op1_00_in07 = reg_0988;
    71: op1_00_in07 = reg_0716;
    72: op1_00_in07 = imem03_in[47:44];
    73: op1_00_in07 = reg_1046;
    74: op1_00_in07 = reg_0696;
    75: op1_00_in07 = reg_0159;
    76: op1_00_in07 = reg_0464;
    78: op1_00_in07 = reg_0099;
    79: op1_00_in07 = reg_0950;
    80: op1_00_in07 = reg_0689;
    83: op1_00_in07 = reg_0056;
    84: op1_00_in07 = reg_0608;
    85: op1_00_in07 = reg_0238;
    86: op1_00_in07 = reg_0573;
    87: op1_00_in07 = imem06_in[3:0];
    88: op1_00_in07 = reg_0985;
    89: op1_00_in07 = imem07_in[103:100];
    90: op1_00_in07 = imem04_in[119:116];
    91: op1_00_in07 = reg_0972;
    92: op1_00_in07 = reg_0121;
    93: op1_00_in07 = reg_0827;
    95: op1_00_in07 = reg_0115;
    96: op1_00_in07 = reg_0521;
    97: op1_00_in07 = reg_0386;
    default: op1_00_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv07 = 1;
    4: op1_00_inv07 = 1;
    7: op1_00_inv07 = 1;
    12: op1_00_inv07 = 1;
    13: op1_00_inv07 = 1;
    15: op1_00_inv07 = 1;
    17: op1_00_inv07 = 1;
    19: op1_00_inv07 = 1;
    25: op1_00_inv07 = 1;
    28: op1_00_inv07 = 1;
    29: op1_00_inv07 = 1;
    30: op1_00_inv07 = 1;
    31: op1_00_inv07 = 1;
    32: op1_00_inv07 = 1;
    33: op1_00_inv07 = 1;
    38: op1_00_inv07 = 1;
    41: op1_00_inv07 = 1;
    42: op1_00_inv07 = 1;
    44: op1_00_inv07 = 1;
    45: op1_00_inv07 = 1;
    46: op1_00_inv07 = 1;
    47: op1_00_inv07 = 1;
    48: op1_00_inv07 = 1;
    51: op1_00_inv07 = 1;
    53: op1_00_inv07 = 1;
    55: op1_00_inv07 = 1;
    58: op1_00_inv07 = 1;
    59: op1_00_inv07 = 1;
    60: op1_00_inv07 = 1;
    62: op1_00_inv07 = 1;
    63: op1_00_inv07 = 1;
    65: op1_00_inv07 = 1;
    68: op1_00_inv07 = 1;
    69: op1_00_inv07 = 1;
    71: op1_00_inv07 = 1;
    72: op1_00_inv07 = 1;
    73: op1_00_inv07 = 1;
    74: op1_00_inv07 = 1;
    75: op1_00_inv07 = 1;
    76: op1_00_inv07 = 1;
    79: op1_00_inv07 = 1;
    80: op1_00_inv07 = 1;
    84: op1_00_inv07 = 1;
    87: op1_00_inv07 = 1;
    88: op1_00_inv07 = 1;
    89: op1_00_inv07 = 1;
    90: op1_00_inv07 = 1;
    91: op1_00_inv07 = 1;
    92: op1_00_inv07 = 1;
    94: op1_00_inv07 = 1;
    95: op1_00_inv07 = 1;
    96: op1_00_inv07 = 1;
    97: op1_00_inv07 = 1;
    default: op1_00_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in08 = reg_0688;
    6: op1_00_in08 = reg_0277;
    7: op1_00_in08 = reg_0453;
    8: op1_00_in08 = reg_0554;
    9: op1_00_in08 = reg_0426;
    10: op1_00_in08 = reg_0099;
    11: op1_00_in08 = reg_1038;
    25: op1_00_in08 = reg_1038;
    12: op1_00_in08 = reg_0625;
    13: op1_00_in08 = reg_0467;
    14: op1_00_in08 = reg_0835;
    15: op1_00_in08 = reg_0679;
    16: op1_00_in08 = reg_0479;
    17: op1_00_in08 = reg_0321;
    18: op1_00_in08 = reg_0251;
    19: op1_00_in08 = reg_0970;
    91: op1_00_in08 = reg_0970;
    20: op1_00_in08 = imem06_in[27:24];
    87: op1_00_in08 = imem06_in[27:24];
    21: op1_00_in08 = imem03_in[99:96];
    22: op1_00_in08 = reg_0632;
    23: op1_00_in08 = reg_0452;
    24: op1_00_in08 = imem05_in[11:8];
    26: op1_00_in08 = imem03_in[79:76];
    27: op1_00_in08 = reg_0692;
    39: op1_00_in08 = reg_0692;
    28: op1_00_in08 = imem04_in[15:12];
    29: op1_00_in08 = reg_0005;
    30: op1_00_in08 = reg_0673;
    31: op1_00_in08 = reg_0999;
    32: op1_00_in08 = imem07_in[79:76];
    33: op1_00_in08 = reg_0466;
    76: op1_00_in08 = reg_0466;
    34: op1_00_in08 = reg_0450;
    35: op1_00_in08 = reg_0243;
    36: op1_00_in08 = reg_0390;
    37: op1_00_in08 = reg_0704;
    38: op1_00_in08 = reg_0475;
    40: op1_00_in08 = reg_0650;
    41: op1_00_in08 = reg_0112;
    42: op1_00_in08 = imem05_in[87:84];
    49: op1_00_in08 = imem05_in[87:84];
    44: op1_00_in08 = reg_0675;
    45: op1_00_in08 = reg_0867;
    52: op1_00_in08 = reg_0867;
    46: op1_00_in08 = reg_0962;
    47: op1_00_in08 = reg_0677;
    48: op1_00_in08 = reg_0610;
    50: op1_00_in08 = reg_0895;
    51: op1_00_in08 = reg_0888;
    53: op1_00_in08 = reg_0643;
    54: op1_00_in08 = reg_0836;
    55: op1_00_in08 = reg_0992;
    56: op1_00_in08 = reg_0143;
    57: op1_00_in08 = reg_0640;
    58: op1_00_in08 = imem07_in[51:48];
    59: op1_00_in08 = imem05_in[119:116];
    60: op1_00_in08 = reg_0738;
    61: op1_00_in08 = reg_0728;
    62: op1_00_in08 = reg_0474;
    63: op1_00_in08 = reg_0087;
    64: op1_00_in08 = reg_0296;
    65: op1_00_in08 = reg_0135;
    66: op1_00_in08 = reg_0142;
    67: op1_00_in08 = reg_0010;
    68: op1_00_in08 = reg_0274;
    69: op1_00_in08 = reg_1017;
    70: op1_00_in08 = reg_0990;
    71: op1_00_in08 = reg_0720;
    72: op1_00_in08 = imem03_in[59:56];
    73: op1_00_in08 = reg_0147;
    74: op1_00_in08 = reg_0351;
    75: op1_00_in08 = reg_0177;
    77: op1_00_in08 = reg_0674;
    78: op1_00_in08 = reg_0396;
    79: op1_00_in08 = reg_0949;
    80: op1_00_in08 = reg_0057;
    83: op1_00_in08 = reg_0302;
    84: op1_00_in08 = reg_0347;
    85: op1_00_in08 = reg_0756;
    86: op1_00_in08 = imem07_in[11:8];
    88: op1_00_in08 = reg_0993;
    89: op1_00_in08 = reg_0567;
    90: op1_00_in08 = reg_0577;
    92: op1_00_in08 = reg_0783;
    93: op1_00_in08 = reg_0101;
    94: op1_00_in08 = reg_1055;
    95: op1_00_in08 = reg_0109;
    96: op1_00_in08 = reg_0810;
    97: op1_00_in08 = reg_0345;
    default: op1_00_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv08 = 1;
    6: op1_00_inv08 = 1;
    7: op1_00_inv08 = 1;
    9: op1_00_inv08 = 1;
    11: op1_00_inv08 = 1;
    14: op1_00_inv08 = 1;
    15: op1_00_inv08 = 1;
    16: op1_00_inv08 = 1;
    18: op1_00_inv08 = 1;
    21: op1_00_inv08 = 1;
    22: op1_00_inv08 = 1;
    24: op1_00_inv08 = 1;
    25: op1_00_inv08 = 1;
    26: op1_00_inv08 = 1;
    27: op1_00_inv08 = 1;
    30: op1_00_inv08 = 1;
    31: op1_00_inv08 = 1;
    35: op1_00_inv08 = 1;
    36: op1_00_inv08 = 1;
    37: op1_00_inv08 = 1;
    38: op1_00_inv08 = 1;
    39: op1_00_inv08 = 1;
    42: op1_00_inv08 = 1;
    45: op1_00_inv08 = 1;
    46: op1_00_inv08 = 1;
    47: op1_00_inv08 = 1;
    48: op1_00_inv08 = 1;
    51: op1_00_inv08 = 1;
    54: op1_00_inv08 = 1;
    55: op1_00_inv08 = 1;
    56: op1_00_inv08 = 1;
    57: op1_00_inv08 = 1;
    58: op1_00_inv08 = 1;
    60: op1_00_inv08 = 1;
    61: op1_00_inv08 = 1;
    63: op1_00_inv08 = 1;
    65: op1_00_inv08 = 1;
    66: op1_00_inv08 = 1;
    67: op1_00_inv08 = 1;
    68: op1_00_inv08 = 1;
    70: op1_00_inv08 = 1;
    71: op1_00_inv08 = 1;
    73: op1_00_inv08 = 1;
    75: op1_00_inv08 = 1;
    77: op1_00_inv08 = 1;
    79: op1_00_inv08 = 1;
    80: op1_00_inv08 = 1;
    84: op1_00_inv08 = 1;
    85: op1_00_inv08 = 1;
    86: op1_00_inv08 = 1;
    93: op1_00_inv08 = 1;
    94: op1_00_inv08 = 1;
    96: op1_00_inv08 = 1;
    default: op1_00_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in09 = reg_0673;
    6: op1_00_in09 = reg_0306;
    7: op1_00_in09 = reg_0200;
    8: op1_00_in09 = reg_0546;
    9: op1_00_in09 = reg_0418;
    10: op1_00_in09 = reg_0112;
    11: op1_00_in09 = reg_0122;
    12: op1_00_in09 = reg_0612;
    13: op1_00_in09 = reg_0479;
    14: op1_00_in09 = reg_0900;
    15: op1_00_in09 = reg_0691;
    47: op1_00_in09 = reg_0691;
    16: op1_00_in09 = reg_0478;
    17: op1_00_in09 = reg_0311;
    18: op1_00_in09 = reg_0147;
    19: op1_00_in09 = reg_0956;
    20: op1_00_in09 = imem06_in[91:88];
    21: op1_00_in09 = imem03_in[107:104];
    22: op1_00_in09 = reg_0622;
    23: op1_00_in09 = reg_0214;
    24: op1_00_in09 = imem05_in[19:16];
    25: op1_00_in09 = reg_0904;
    26: op1_00_in09 = imem03_in[103:100];
    27: op1_00_in09 = reg_0457;
    39: op1_00_in09 = reg_0457;
    28: op1_00_in09 = imem04_in[51:48];
    29: op1_00_in09 = imem07_in[23:20];
    30: op1_00_in09 = reg_0477;
    31: op1_00_in09 = reg_0975;
    32: op1_00_in09 = imem07_in[115:112];
    33: op1_00_in09 = reg_0462;
    34: op1_00_in09 = reg_0476;
    35: op1_00_in09 = reg_0399;
    36: op1_00_in09 = reg_0349;
    37: op1_00_in09 = reg_0719;
    61: op1_00_in09 = reg_0719;
    38: op1_00_in09 = reg_0480;
    40: op1_00_in09 = reg_0645;
    41: op1_00_in09 = reg_0108;
    42: op1_00_in09 = imem05_in[107:104];
    44: op1_00_in09 = reg_0687;
    77: op1_00_in09 = reg_0687;
    45: op1_00_in09 = reg_0261;
    46: op1_00_in09 = reg_0955;
    48: op1_00_in09 = reg_0304;
    49: op1_00_in09 = imem05_in[95:92];
    50: op1_00_in09 = reg_0533;
    51: op1_00_in09 = reg_0050;
    52: op1_00_in09 = reg_0086;
    53: op1_00_in09 = reg_0818;
    54: op1_00_in09 = reg_0822;
    55: op1_00_in09 = reg_0993;
    56: op1_00_in09 = imem06_in[27:24];
    57: op1_00_in09 = reg_0175;
    58: op1_00_in09 = imem07_in[59:56];
    59: op1_00_in09 = reg_0255;
    60: op1_00_in09 = reg_0883;
    62: op1_00_in09 = reg_0459;
    63: op1_00_in09 = reg_0335;
    64: op1_00_in09 = reg_0627;
    65: op1_00_in09 = reg_0128;
    66: op1_00_in09 = reg_0156;
    67: op1_00_in09 = reg_0694;
    68: op1_00_in09 = reg_0784;
    69: op1_00_in09 = reg_1051;
    70: op1_00_in09 = reg_0983;
    71: op1_00_in09 = reg_0726;
    89: op1_00_in09 = reg_0726;
    72: op1_00_in09 = imem03_in[75:72];
    73: op1_00_in09 = reg_0148;
    74: op1_00_in09 = reg_0267;
    75: op1_00_in09 = reg_0164;
    76: op1_00_in09 = reg_0475;
    78: op1_00_in09 = reg_0661;
    79: op1_00_in09 = reg_0945;
    91: op1_00_in09 = reg_0945;
    80: op1_00_in09 = reg_0149;
    83: op1_00_in09 = reg_0074;
    84: op1_00_in09 = reg_0007;
    85: op1_00_in09 = reg_1008;
    86: op1_00_in09 = imem07_in[43:40];
    87: op1_00_in09 = imem06_in[83:80];
    88: op1_00_in09 = reg_0986;
    90: op1_00_in09 = reg_0937;
    92: op1_00_in09 = reg_0034;
    93: op1_00_in09 = reg_0110;
    94: op1_00_in09 = reg_0769;
    95: op1_00_in09 = reg_0821;
    96: op1_00_in09 = reg_0160;
    97: op1_00_in09 = reg_0186;
    default: op1_00_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_00_inv09 = 1;
    8: op1_00_inv09 = 1;
    11: op1_00_inv09 = 1;
    13: op1_00_inv09 = 1;
    15: op1_00_inv09 = 1;
    17: op1_00_inv09 = 1;
    18: op1_00_inv09 = 1;
    21: op1_00_inv09 = 1;
    24: op1_00_inv09 = 1;
    27: op1_00_inv09 = 1;
    33: op1_00_inv09 = 1;
    35: op1_00_inv09 = 1;
    37: op1_00_inv09 = 1;
    40: op1_00_inv09 = 1;
    41: op1_00_inv09 = 1;
    45: op1_00_inv09 = 1;
    47: op1_00_inv09 = 1;
    48: op1_00_inv09 = 1;
    50: op1_00_inv09 = 1;
    54: op1_00_inv09 = 1;
    55: op1_00_inv09 = 1;
    57: op1_00_inv09 = 1;
    66: op1_00_inv09 = 1;
    67: op1_00_inv09 = 1;
    73: op1_00_inv09 = 1;
    75: op1_00_inv09 = 1;
    76: op1_00_inv09 = 1;
    80: op1_00_inv09 = 1;
    83: op1_00_inv09 = 1;
    86: op1_00_inv09 = 1;
    88: op1_00_inv09 = 1;
    90: op1_00_inv09 = 1;
    93: op1_00_inv09 = 1;
    default: op1_00_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in10 = reg_0669;
    6: op1_00_in10 = reg_0292;
    7: op1_00_in10 = reg_0189;
    8: op1_00_in10 = reg_0558;
    9: op1_00_in10 = reg_0445;
    10: op1_00_in10 = reg_0108;
    11: op1_00_in10 = reg_0119;
    25: op1_00_in10 = reg_0119;
    48: op1_00_in10 = reg_0119;
    12: op1_00_in10 = reg_0402;
    36: op1_00_in10 = reg_0402;
    13: op1_00_in10 = reg_0459;
    34: op1_00_in10 = reg_0459;
    76: op1_00_in10 = reg_0459;
    14: op1_00_in10 = reg_0256;
    15: op1_00_in10 = reg_0678;
    16: op1_00_in10 = reg_0208;
    17: op1_00_in10 = reg_0385;
    18: op1_00_in10 = reg_0136;
    19: op1_00_in10 = reg_0957;
    20: op1_00_in10 = reg_0620;
    21: op1_00_in10 = reg_0569;
    22: op1_00_in10 = reg_0405;
    23: op1_00_in10 = reg_0193;
    24: op1_00_in10 = imem05_in[31:28];
    26: op1_00_in10 = imem03_in[115:112];
    27: op1_00_in10 = reg_0466;
    28: op1_00_in10 = imem04_in[91:88];
    29: op1_00_in10 = imem07_in[27:24];
    30: op1_00_in10 = reg_0456;
    31: op1_00_in10 = reg_0988;
    32: op1_00_in10 = imem07_in[127:124];
    33: op1_00_in10 = reg_0480;
    35: op1_00_in10 = reg_0332;
    37: op1_00_in10 = reg_0700;
    38: op1_00_in10 = reg_0473;
    39: op1_00_in10 = reg_0461;
    40: op1_00_in10 = reg_0646;
    41: op1_00_in10 = reg_0110;
    42: op1_00_in10 = reg_0962;
    44: op1_00_in10 = reg_0454;
    45: op1_00_in10 = reg_0091;
    46: op1_00_in10 = reg_0964;
    47: op1_00_in10 = reg_0674;
    49: op1_00_in10 = imem05_in[103:100];
    50: op1_00_in10 = reg_0782;
    51: op1_00_in10 = reg_0059;
    52: op1_00_in10 = reg_0506;
    53: op1_00_in10 = reg_0482;
    54: op1_00_in10 = reg_0984;
    55: op1_00_in10 = reg_0986;
    56: op1_00_in10 = imem06_in[35:32];
    57: op1_00_in10 = reg_0164;
    58: op1_00_in10 = imem07_in[71:68];
    59: op1_00_in10 = reg_0492;
    60: op1_00_in10 = reg_0668;
    61: op1_00_in10 = reg_0720;
    62: op1_00_in10 = reg_0191;
    63: op1_00_in10 = reg_0347;
    64: op1_00_in10 = reg_0824;
    65: op1_00_in10 = reg_0152;
    66: op1_00_in10 = reg_0144;
    67: op1_00_in10 = reg_1019;
    68: op1_00_in10 = reg_0004;
    69: op1_00_in10 = reg_0109;
    70: op1_00_in10 = imem04_in[11:8];
    71: op1_00_in10 = reg_0705;
    72: op1_00_in10 = imem03_in[103:100];
    73: op1_00_in10 = reg_0150;
    74: op1_00_in10 = reg_0338;
    77: op1_00_in10 = reg_0453;
    78: op1_00_in10 = reg_0576;
    79: op1_00_in10 = imem06_in[23:20];
    80: op1_00_in10 = reg_0107;
    83: op1_00_in10 = reg_0065;
    84: op1_00_in10 = reg_0876;
    85: op1_00_in10 = reg_0779;
    86: op1_00_in10 = imem07_in[47:44];
    87: op1_00_in10 = imem06_in[95:92];
    88: op1_00_in10 = imem04_in[15:12];
    89: op1_00_in10 = reg_0717;
    90: op1_00_in10 = reg_0912;
    91: op1_00_in10 = imem06_in[71:68];
    92: op1_00_in10 = reg_0036;
    93: op1_00_in10 = imem02_in[23:20];
    94: op1_00_in10 = reg_0116;
    95: op1_00_in10 = imem02_in[31:28];
    96: op1_00_in10 = reg_0333;
    97: op1_00_in10 = reg_0871;
    default: op1_00_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_00_inv10 = 1;
    10: op1_00_inv10 = 1;
    12: op1_00_inv10 = 1;
    13: op1_00_inv10 = 1;
    15: op1_00_inv10 = 1;
    17: op1_00_inv10 = 1;
    18: op1_00_inv10 = 1;
    20: op1_00_inv10 = 1;
    21: op1_00_inv10 = 1;
    22: op1_00_inv10 = 1;
    23: op1_00_inv10 = 1;
    24: op1_00_inv10 = 1;
    26: op1_00_inv10 = 1;
    27: op1_00_inv10 = 1;
    28: op1_00_inv10 = 1;
    29: op1_00_inv10 = 1;
    34: op1_00_inv10 = 1;
    37: op1_00_inv10 = 1;
    41: op1_00_inv10 = 1;
    46: op1_00_inv10 = 1;
    47: op1_00_inv10 = 1;
    51: op1_00_inv10 = 1;
    53: op1_00_inv10 = 1;
    55: op1_00_inv10 = 1;
    59: op1_00_inv10 = 1;
    60: op1_00_inv10 = 1;
    62: op1_00_inv10 = 1;
    67: op1_00_inv10 = 1;
    68: op1_00_inv10 = 1;
    69: op1_00_inv10 = 1;
    70: op1_00_inv10 = 1;
    72: op1_00_inv10 = 1;
    74: op1_00_inv10 = 1;
    76: op1_00_inv10 = 1;
    79: op1_00_inv10 = 1;
    83: op1_00_inv10 = 1;
    85: op1_00_inv10 = 1;
    92: op1_00_inv10 = 1;
    94: op1_00_inv10 = 1;
    95: op1_00_inv10 = 1;
    96: op1_00_inv10 = 1;
    97: op1_00_inv10 = 1;
    default: op1_00_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in11 = reg_0465;
    96: op1_00_in11 = reg_0465;
    6: op1_00_in11 = reg_0275;
    7: op1_00_in11 = reg_0204;
    8: op1_00_in11 = reg_0304;
    9: op1_00_in11 = reg_0446;
    10: op1_00_in11 = reg_0114;
    11: op1_00_in11 = reg_0112;
    12: op1_00_in11 = reg_0405;
    13: op1_00_in11 = reg_0214;
    14: op1_00_in11 = reg_0908;
    15: op1_00_in11 = reg_0668;
    16: op1_00_in11 = reg_0188;
    17: op1_00_in11 = reg_0376;
    18: op1_00_in11 = reg_0142;
    65: op1_00_in11 = reg_0142;
    19: op1_00_in11 = reg_0949;
    20: op1_00_in11 = reg_0621;
    21: op1_00_in11 = reg_0563;
    22: op1_00_in11 = reg_0404;
    23: op1_00_in11 = reg_0201;
    34: op1_00_in11 = reg_0201;
    24: op1_00_in11 = imem05_in[59:56];
    25: op1_00_in11 = reg_0110;
    26: op1_00_in11 = reg_0583;
    27: op1_00_in11 = reg_0467;
    28: op1_00_in11 = imem04_in[103:100];
    29: op1_00_in11 = imem07_in[31:28];
    30: op1_00_in11 = reg_0458;
    31: op1_00_in11 = reg_0994;
    32: op1_00_in11 = reg_0729;
    33: op1_00_in11 = reg_0473;
    35: op1_00_in11 = reg_0780;
    36: op1_00_in11 = reg_0808;
    37: op1_00_in11 = reg_0419;
    38: op1_00_in11 = reg_0468;
    39: op1_00_in11 = reg_0460;
    40: op1_00_in11 = reg_0638;
    41: op1_00_in11 = imem02_in[19:16];
    42: op1_00_in11 = reg_0970;
    44: op1_00_in11 = reg_0466;
    45: op1_00_in11 = reg_0840;
    46: op1_00_in11 = reg_0961;
    47: op1_00_in11 = reg_0671;
    48: op1_00_in11 = reg_0108;
    83: op1_00_in11 = reg_0108;
    49: op1_00_in11 = imem05_in[115:112];
    50: op1_00_in11 = reg_0754;
    51: op1_00_in11 = reg_0078;
    52: op1_00_in11 = reg_0261;
    53: op1_00_in11 = reg_0792;
    54: op1_00_in11 = reg_0978;
    55: op1_00_in11 = reg_0974;
    56: op1_00_in11 = imem06_in[59:56];
    57: op1_00_in11 = reg_0157;
    58: op1_00_in11 = imem07_in[83:80];
    59: op1_00_in11 = reg_0952;
    60: op1_00_in11 = reg_0102;
    61: op1_00_in11 = reg_0730;
    62: op1_00_in11 = reg_0210;
    63: op1_00_in11 = reg_0079;
    64: op1_00_in11 = reg_0295;
    66: op1_00_in11 = imem06_in[3:0];
    67: op1_00_in11 = reg_0691;
    68: op1_00_in11 = reg_0135;
    69: op1_00_in11 = imem02_in[31:28];
    70: op1_00_in11 = imem04_in[59:56];
    71: op1_00_in11 = reg_0361;
    72: op1_00_in11 = reg_0006;
    73: op1_00_in11 = imem06_in[7:4];
    74: op1_00_in11 = reg_0533;
    76: op1_00_in11 = reg_0209;
    77: op1_00_in11 = reg_0457;
    78: op1_00_in11 = reg_0281;
    79: op1_00_in11 = imem06_in[63:60];
    80: op1_00_in11 = reg_0967;
    84: op1_00_in11 = reg_0506;
    85: op1_00_in11 = reg_0597;
    86: op1_00_in11 = imem07_in[51:48];
    87: op1_00_in11 = imem06_in[103:100];
    88: op1_00_in11 = imem04_in[19:16];
    89: op1_00_in11 = reg_0374;
    90: op1_00_in11 = reg_0430;
    91: op1_00_in11 = imem06_in[83:80];
    92: op1_00_in11 = reg_0018;
    93: op1_00_in11 = imem02_in[107:104];
    94: op1_00_in11 = reg_0860;
    95: op1_00_in11 = imem02_in[39:36];
    97: op1_00_in11 = reg_0030;
    default: op1_00_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv11 = 1;
    6: op1_00_inv11 = 1;
    7: op1_00_inv11 = 1;
    8: op1_00_inv11 = 1;
    9: op1_00_inv11 = 1;
    10: op1_00_inv11 = 1;
    11: op1_00_inv11 = 1;
    12: op1_00_inv11 = 1;
    15: op1_00_inv11 = 1;
    16: op1_00_inv11 = 1;
    17: op1_00_inv11 = 1;
    18: op1_00_inv11 = 1;
    19: op1_00_inv11 = 1;
    21: op1_00_inv11 = 1;
    23: op1_00_inv11 = 1;
    24: op1_00_inv11 = 1;
    27: op1_00_inv11 = 1;
    28: op1_00_inv11 = 1;
    29: op1_00_inv11 = 1;
    30: op1_00_inv11 = 1;
    34: op1_00_inv11 = 1;
    35: op1_00_inv11 = 1;
    38: op1_00_inv11 = 1;
    41: op1_00_inv11 = 1;
    44: op1_00_inv11 = 1;
    45: op1_00_inv11 = 1;
    46: op1_00_inv11 = 1;
    51: op1_00_inv11 = 1;
    53: op1_00_inv11 = 1;
    54: op1_00_inv11 = 1;
    55: op1_00_inv11 = 1;
    57: op1_00_inv11 = 1;
    58: op1_00_inv11 = 1;
    59: op1_00_inv11 = 1;
    63: op1_00_inv11 = 1;
    65: op1_00_inv11 = 1;
    66: op1_00_inv11 = 1;
    67: op1_00_inv11 = 1;
    69: op1_00_inv11 = 1;
    72: op1_00_inv11 = 1;
    74: op1_00_inv11 = 1;
    76: op1_00_inv11 = 1;
    78: op1_00_inv11 = 1;
    79: op1_00_inv11 = 1;
    84: op1_00_inv11 = 1;
    85: op1_00_inv11 = 1;
    86: op1_00_inv11 = 1;
    91: op1_00_inv11 = 1;
    93: op1_00_inv11 = 1;
    default: op1_00_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in12 = reg_0451;
    15: op1_00_in12 = reg_0451;
    60: op1_00_in12 = reg_0451;
    6: op1_00_in12 = reg_0041;
    7: op1_00_in12 = reg_0193;
    76: op1_00_in12 = reg_0193;
    8: op1_00_in12 = reg_0292;
    9: op1_00_in12 = reg_0442;
    10: op1_00_in12 = reg_0101;
    11: op1_00_in12 = reg_0115;
    12: op1_00_in12 = reg_0409;
    13: op1_00_in12 = reg_0200;
    14: op1_00_in12 = reg_0822;
    16: op1_00_in12 = reg_0213;
    17: op1_00_in12 = reg_1001;
    18: op1_00_in12 = reg_0146;
    19: op1_00_in12 = reg_0946;
    20: op1_00_in12 = reg_0622;
    21: op1_00_in12 = reg_0391;
    22: op1_00_in12 = reg_0486;
    23: op1_00_in12 = reg_0202;
    24: op1_00_in12 = imem05_in[95:92];
    25: op1_00_in12 = imem02_in[7:4];
    26: op1_00_in12 = reg_0572;
    27: op1_00_in12 = reg_0468;
    28: op1_00_in12 = imem04_in[107:104];
    29: op1_00_in12 = imem07_in[35:32];
    30: op1_00_in12 = reg_0204;
    31: op1_00_in12 = imem04_in[3:0];
    32: op1_00_in12 = reg_0432;
    33: op1_00_in12 = reg_0474;
    34: op1_00_in12 = imem01_in[39:36];
    35: op1_00_in12 = reg_0405;
    36: op1_00_in12 = reg_0032;
    37: op1_00_in12 = reg_0434;
    38: op1_00_in12 = reg_0214;
    39: op1_00_in12 = reg_0473;
    40: op1_00_in12 = reg_0665;
    41: op1_00_in12 = imem02_in[47:44];
    42: op1_00_in12 = reg_0944;
    44: op1_00_in12 = reg_0475;
    45: op1_00_in12 = reg_0310;
    46: op1_00_in12 = reg_0953;
    47: op1_00_in12 = reg_0680;
    48: op1_00_in12 = reg_0114;
    49: op1_00_in12 = reg_0958;
    50: op1_00_in12 = reg_0495;
    51: op1_00_in12 = reg_0529;
    52: op1_00_in12 = reg_0084;
    53: op1_00_in12 = imem03_in[7:4];
    54: op1_00_in12 = reg_0999;
    55: op1_00_in12 = reg_0977;
    56: op1_00_in12 = imem06_in[63:60];
    57: op1_00_in12 = reg_0176;
    58: op1_00_in12 = imem07_in[103:100];
    59: op1_00_in12 = reg_0488;
    61: op1_00_in12 = reg_0726;
    62: op1_00_in12 = reg_0188;
    63: op1_00_in12 = imem03_in[87:84];
    64: op1_00_in12 = reg_0044;
    65: op1_00_in12 = reg_0156;
    66: op1_00_in12 = imem06_in[31:28];
    67: op1_00_in12 = reg_0267;
    68: op1_00_in12 = reg_0136;
    69: op1_00_in12 = imem02_in[59:56];
    70: op1_00_in12 = imem04_in[63:60];
    71: op1_00_in12 = reg_0426;
    72: op1_00_in12 = reg_0620;
    73: op1_00_in12 = imem06_in[11:8];
    74: op1_00_in12 = reg_0008;
    77: op1_00_in12 = reg_0461;
    78: op1_00_in12 = reg_0579;
    79: op1_00_in12 = imem06_in[119:116];
    80: op1_00_in12 = reg_0964;
    83: op1_00_in12 = reg_0856;
    84: op1_00_in12 = imem03_in[39:36];
    85: op1_00_in12 = reg_0975;
    86: op1_00_in12 = imem07_in[67:64];
    87: op1_00_in12 = imem06_in[107:104];
    88: op1_00_in12 = imem04_in[51:48];
    89: op1_00_in12 = reg_0560;
    90: op1_00_in12 = reg_0031;
    91: op1_00_in12 = imem06_in[99:96];
    92: op1_00_in12 = reg_0403;
    93: op1_00_in12 = reg_0916;
    94: op1_00_in12 = reg_0827;
    95: op1_00_in12 = imem02_in[71:68];
    96: op1_00_in12 = reg_0472;
    97: op1_00_in12 = reg_0477;
    default: op1_00_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv12 = 1;
    8: op1_00_inv12 = 1;
    9: op1_00_inv12 = 1;
    10: op1_00_inv12 = 1;
    11: op1_00_inv12 = 1;
    12: op1_00_inv12 = 1;
    13: op1_00_inv12 = 1;
    15: op1_00_inv12 = 1;
    16: op1_00_inv12 = 1;
    17: op1_00_inv12 = 1;
    18: op1_00_inv12 = 1;
    19: op1_00_inv12 = 1;
    20: op1_00_inv12 = 1;
    22: op1_00_inv12 = 1;
    23: op1_00_inv12 = 1;
    24: op1_00_inv12 = 1;
    25: op1_00_inv12 = 1;
    27: op1_00_inv12 = 1;
    28: op1_00_inv12 = 1;
    31: op1_00_inv12 = 1;
    32: op1_00_inv12 = 1;
    34: op1_00_inv12 = 1;
    37: op1_00_inv12 = 1;
    38: op1_00_inv12 = 1;
    40: op1_00_inv12 = 1;
    44: op1_00_inv12 = 1;
    46: op1_00_inv12 = 1;
    49: op1_00_inv12 = 1;
    51: op1_00_inv12 = 1;
    53: op1_00_inv12 = 1;
    55: op1_00_inv12 = 1;
    56: op1_00_inv12 = 1;
    60: op1_00_inv12 = 1;
    61: op1_00_inv12 = 1;
    62: op1_00_inv12 = 1;
    64: op1_00_inv12 = 1;
    67: op1_00_inv12 = 1;
    68: op1_00_inv12 = 1;
    70: op1_00_inv12 = 1;
    71: op1_00_inv12 = 1;
    73: op1_00_inv12 = 1;
    76: op1_00_inv12 = 1;
    78: op1_00_inv12 = 1;
    79: op1_00_inv12 = 1;
    86: op1_00_inv12 = 1;
    87: op1_00_inv12 = 1;
    88: op1_00_inv12 = 1;
    89: op1_00_inv12 = 1;
    90: op1_00_inv12 = 1;
    91: op1_00_inv12 = 1;
    93: op1_00_inv12 = 1;
    94: op1_00_inv12 = 1;
    95: op1_00_inv12 = 1;
    96: op1_00_inv12 = 1;
    97: op1_00_inv12 = 1;
    default: op1_00_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in13 = reg_0455;
    6: op1_00_in13 = reg_0065;
    7: op1_00_in13 = reg_0195;
    8: op1_00_in13 = reg_0295;
    9: op1_00_in13 = reg_0443;
    10: op1_00_in13 = reg_0109;
    11: op1_00_in13 = reg_0110;
    12: op1_00_in13 = reg_0337;
    13: op1_00_in13 = reg_0203;
    14: op1_00_in13 = reg_0865;
    15: op1_00_in13 = reg_0466;
    16: op1_00_in13 = reg_0205;
    17: op1_00_in13 = reg_0974;
    18: op1_00_in13 = reg_0143;
    65: op1_00_in13 = reg_0143;
    19: op1_00_in13 = reg_0903;
    20: op1_00_in13 = reg_0348;
    21: op1_00_in13 = reg_0321;
    22: op1_00_in13 = reg_0781;
    23: op1_00_in13 = reg_0199;
    24: op1_00_in13 = imem05_in[103:100];
    25: op1_00_in13 = imem02_in[23:20];
    26: op1_00_in13 = reg_0576;
    27: op1_00_in13 = reg_0459;
    28: op1_00_in13 = reg_0530;
    29: op1_00_in13 = imem07_in[39:36];
    30: op1_00_in13 = reg_0207;
    31: op1_00_in13 = imem04_in[63:60];
    32: op1_00_in13 = reg_0422;
    33: op1_00_in13 = reg_0456;
    34: op1_00_in13 = imem01_in[87:84];
    35: op1_00_in13 = reg_1010;
    36: op1_00_in13 = reg_0405;
    37: op1_00_in13 = reg_0446;
    38: op1_00_in13 = reg_0210;
    39: op1_00_in13 = reg_0470;
    40: op1_00_in13 = reg_0095;
    41: op1_00_in13 = imem02_in[71:68];
    42: op1_00_in13 = reg_0957;
    49: op1_00_in13 = reg_0957;
    44: op1_00_in13 = reg_0481;
    45: op1_00_in13 = reg_0291;
    46: op1_00_in13 = reg_1021;
    47: op1_00_in13 = reg_0673;
    48: op1_00_in13 = reg_0113;
    50: op1_00_in13 = reg_0293;
    51: op1_00_in13 = reg_0764;
    52: op1_00_in13 = reg_0016;
    53: op1_00_in13 = imem03_in[15:12];
    54: op1_00_in13 = imem04_in[7:4];
    55: op1_00_in13 = imem04_in[27:24];
    56: op1_00_in13 = imem06_in[71:68];
    57: op1_00_in13 = reg_0171;
    58: op1_00_in13 = reg_0728;
    59: op1_00_in13 = reg_0148;
    60: op1_00_in13 = reg_0457;
    61: op1_00_in13 = reg_0717;
    62: op1_00_in13 = reg_0201;
    63: op1_00_in13 = imem03_in[123:120];
    64: op1_00_in13 = imem05_in[19:16];
    66: op1_00_in13 = imem06_in[67:64];
    67: op1_00_in13 = reg_0262;
    68: op1_00_in13 = reg_0141;
    69: op1_00_in13 = imem02_in[75:72];
    70: op1_00_in13 = imem04_in[75:72];
    71: op1_00_in13 = reg_0315;
    72: op1_00_in13 = reg_0245;
    73: op1_00_in13 = imem06_in[19:16];
    74: op1_00_in13 = reg_0699;
    76: op1_00_in13 = reg_0186;
    77: op1_00_in13 = reg_0475;
    78: op1_00_in13 = reg_0239;
    79: op1_00_in13 = reg_0391;
    80: op1_00_in13 = reg_0265;
    83: op1_00_in13 = imem05_in[11:8];
    84: op1_00_in13 = imem03_in[51:48];
    85: op1_00_in13 = reg_0988;
    86: op1_00_in13 = imem07_in[87:84];
    87: op1_00_in13 = imem06_in[127:124];
    88: op1_00_in13 = reg_0147;
    89: op1_00_in13 = reg_0515;
    90: op1_00_in13 = reg_0066;
    91: op1_00_in13 = imem06_in[103:100];
    92: op1_00_in13 = imem07_in[3:0];
    93: op1_00_in13 = reg_0543;
    94: op1_00_in13 = reg_0745;
    95: op1_00_in13 = imem02_in[91:88];
    96: op1_00_in13 = reg_0480;
    97: op1_00_in13 = reg_0476;
    default: op1_00_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv13 = 1;
    6: op1_00_inv13 = 1;
    8: op1_00_inv13 = 1;
    9: op1_00_inv13 = 1;
    15: op1_00_inv13 = 1;
    16: op1_00_inv13 = 1;
    17: op1_00_inv13 = 1;
    18: op1_00_inv13 = 1;
    19: op1_00_inv13 = 1;
    20: op1_00_inv13 = 1;
    23: op1_00_inv13 = 1;
    25: op1_00_inv13 = 1;
    26: op1_00_inv13 = 1;
    28: op1_00_inv13 = 1;
    32: op1_00_inv13 = 1;
    33: op1_00_inv13 = 1;
    35: op1_00_inv13 = 1;
    38: op1_00_inv13 = 1;
    39: op1_00_inv13 = 1;
    44: op1_00_inv13 = 1;
    48: op1_00_inv13 = 1;
    49: op1_00_inv13 = 1;
    50: op1_00_inv13 = 1;
    52: op1_00_inv13 = 1;
    53: op1_00_inv13 = 1;
    55: op1_00_inv13 = 1;
    58: op1_00_inv13 = 1;
    59: op1_00_inv13 = 1;
    60: op1_00_inv13 = 1;
    67: op1_00_inv13 = 1;
    69: op1_00_inv13 = 1;
    71: op1_00_inv13 = 1;
    72: op1_00_inv13 = 1;
    74: op1_00_inv13 = 1;
    80: op1_00_inv13 = 1;
    83: op1_00_inv13 = 1;
    85: op1_00_inv13 = 1;
    86: op1_00_inv13 = 1;
    88: op1_00_inv13 = 1;
    91: op1_00_inv13 = 1;
    95: op1_00_inv13 = 1;
    96: op1_00_inv13 = 1;
    default: op1_00_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in14 = reg_0466;
    6: op1_00_in14 = imem05_in[19:16];
    7: op1_00_in14 = imem01_in[3:0];
    8: op1_00_in14 = reg_0065;
    9: op1_00_in14 = reg_0165;
    10: op1_00_in14 = reg_0117;
    11: op1_00_in14 = imem02_in[47:44];
    94: op1_00_in14 = imem02_in[47:44];
    12: op1_00_in14 = reg_0808;
    13: op1_00_in14 = reg_0194;
    14: op1_00_in14 = reg_0145;
    15: op1_00_in14 = reg_0460;
    16: op1_00_in14 = imem01_in[27:24];
    17: op1_00_in14 = imem04_in[47:44];
    55: op1_00_in14 = imem04_in[47:44];
    18: op1_00_in14 = reg_0138;
    19: op1_00_in14 = reg_0250;
    20: op1_00_in14 = reg_0356;
    50: op1_00_in14 = reg_0356;
    21: op1_00_in14 = reg_0369;
    22: op1_00_in14 = reg_1011;
    23: op1_00_in14 = imem01_in[19:16];
    24: op1_00_in14 = imem05_in[119:116];
    25: op1_00_in14 = imem02_in[59:56];
    26: op1_00_in14 = reg_0385;
    27: op1_00_in14 = reg_0452;
    28: op1_00_in14 = reg_0912;
    29: op1_00_in14 = imem07_in[59:56];
    30: op1_00_in14 = reg_0196;
    31: op1_00_in14 = imem04_in[67:64];
    32: op1_00_in14 = reg_0419;
    33: op1_00_in14 = reg_0200;
    34: op1_00_in14 = imem01_in[91:88];
    35: op1_00_in14 = imem07_in[7:4];
    92: op1_00_in14 = imem07_in[7:4];
    36: op1_00_in14 = reg_0018;
    37: op1_00_in14 = reg_0444;
    38: op1_00_in14 = reg_0209;
    39: op1_00_in14 = reg_0468;
    77: op1_00_in14 = reg_0468;
    40: op1_00_in14 = reg_0886;
    41: op1_00_in14 = imem02_in[79:76];
    42: op1_00_in14 = reg_0942;
    44: op1_00_in14 = reg_0480;
    45: op1_00_in14 = imem03_in[27:24];
    46: op1_00_in14 = reg_0835;
    47: op1_00_in14 = reg_0450;
    48: op1_00_in14 = imem02_in[3:0];
    49: op1_00_in14 = reg_0948;
    51: op1_00_in14 = imem05_in[47:44];
    52: op1_00_in14 = reg_0291;
    53: op1_00_in14 = imem03_in[51:48];
    54: op1_00_in14 = imem04_in[31:28];
    56: op1_00_in14 = imem06_in[83:80];
    66: op1_00_in14 = imem06_in[83:80];
    57: op1_00_in14 = reg_0184;
    58: op1_00_in14 = reg_0575;
    59: op1_00_in14 = reg_0154;
    60: op1_00_in14 = reg_0469;
    61: op1_00_in14 = reg_0705;
    62: op1_00_in14 = reg_0212;
    63: op1_00_in14 = reg_0346;
    64: op1_00_in14 = imem05_in[71:68];
    65: op1_00_in14 = imem06_in[35:32];
    67: op1_00_in14 = reg_0626;
    68: op1_00_in14 = reg_0144;
    69: op1_00_in14 = imem02_in[111:108];
    70: op1_00_in14 = imem04_in[123:120];
    71: op1_00_in14 = reg_0427;
    72: op1_00_in14 = reg_0585;
    73: op1_00_in14 = imem06_in[47:44];
    74: op1_00_in14 = reg_0380;
    76: op1_00_in14 = reg_0198;
    78: op1_00_in14 = reg_0040;
    79: op1_00_in14 = reg_0692;
    80: op1_00_in14 = reg_0970;
    83: op1_00_in14 = imem05_in[43:40];
    84: op1_00_in14 = imem03_in[55:52];
    85: op1_00_in14 = reg_1000;
    86: op1_00_in14 = imem07_in[99:96];
    87: op1_00_in14 = reg_0660;
    88: op1_00_in14 = reg_0511;
    89: op1_00_in14 = reg_0718;
    90: op1_00_in14 = reg_0276;
    91: op1_00_in14 = reg_0010;
    93: op1_00_in14 = reg_0358;
    95: op1_00_in14 = imem02_in[119:116];
    96: op1_00_in14 = imem01_in[39:36];
    97: op1_00_in14 = reg_0475;
    default: op1_00_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv14 = 1;
    8: op1_00_inv14 = 1;
    9: op1_00_inv14 = 1;
    10: op1_00_inv14 = 1;
    11: op1_00_inv14 = 1;
    13: op1_00_inv14 = 1;
    15: op1_00_inv14 = 1;
    18: op1_00_inv14 = 1;
    19: op1_00_inv14 = 1;
    20: op1_00_inv14 = 1;
    22: op1_00_inv14 = 1;
    23: op1_00_inv14 = 1;
    24: op1_00_inv14 = 1;
    27: op1_00_inv14 = 1;
    28: op1_00_inv14 = 1;
    33: op1_00_inv14 = 1;
    34: op1_00_inv14 = 1;
    37: op1_00_inv14 = 1;
    38: op1_00_inv14 = 1;
    39: op1_00_inv14 = 1;
    40: op1_00_inv14 = 1;
    44: op1_00_inv14 = 1;
    45: op1_00_inv14 = 1;
    49: op1_00_inv14 = 1;
    50: op1_00_inv14 = 1;
    54: op1_00_inv14 = 1;
    55: op1_00_inv14 = 1;
    56: op1_00_inv14 = 1;
    58: op1_00_inv14 = 1;
    62: op1_00_inv14 = 1;
    68: op1_00_inv14 = 1;
    70: op1_00_inv14 = 1;
    73: op1_00_inv14 = 1;
    74: op1_00_inv14 = 1;
    78: op1_00_inv14 = 1;
    84: op1_00_inv14 = 1;
    86: op1_00_inv14 = 1;
    88: op1_00_inv14 = 1;
    89: op1_00_inv14 = 1;
    90: op1_00_inv14 = 1;
    93: op1_00_inv14 = 1;
    94: op1_00_inv14 = 1;
    95: op1_00_inv14 = 1;
    96: op1_00_inv14 = 1;
    default: op1_00_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in15 = reg_0473;
    6: op1_00_in15 = imem05_in[35:32];
    7: op1_00_in15 = imem01_in[51:48];
    8: op1_00_in15 = reg_0053;
    10: op1_00_in15 = imem02_in[3:0];
    11: op1_00_in15 = imem02_in[51:48];
    12: op1_00_in15 = reg_1028;
    13: op1_00_in15 = reg_0206;
    14: op1_00_in15 = reg_0133;
    15: op1_00_in15 = reg_0209;
    16: op1_00_in15 = imem01_in[127:124];
    17: op1_00_in15 = imem04_in[99:96];
    18: op1_00_in15 = imem06_in[19:16];
    68: op1_00_in15 = imem06_in[19:16];
    19: op1_00_in15 = reg_0908;
    20: op1_00_in15 = reg_0383;
    21: op1_00_in15 = reg_0995;
    22: op1_00_in15 = imem07_in[15:12];
    23: op1_00_in15 = imem01_in[23:20];
    24: op1_00_in15 = reg_0956;
    25: op1_00_in15 = imem02_in[67:64];
    94: op1_00_in15 = imem02_in[67:64];
    26: op1_00_in15 = reg_0374;
    27: op1_00_in15 = reg_0456;
    28: op1_00_in15 = reg_1020;
    29: op1_00_in15 = imem07_in[63:60];
    30: op1_00_in15 = reg_0202;
    31: op1_00_in15 = reg_1004;
    70: op1_00_in15 = reg_1004;
    32: op1_00_in15 = reg_0431;
    33: op1_00_in15 = reg_0211;
    34: op1_00_in15 = imem01_in[103:100];
    35: op1_00_in15 = imem07_in[59:56];
    36: op1_00_in15 = reg_0597;
    78: op1_00_in15 = reg_0597;
    37: op1_00_in15 = reg_0437;
    38: op1_00_in15 = reg_0188;
    39: op1_00_in15 = reg_0459;
    44: op1_00_in15 = reg_0459;
    40: op1_00_in15 = reg_0338;
    41: op1_00_in15 = reg_0666;
    42: op1_00_in15 = reg_0968;
    45: op1_00_in15 = imem03_in[39:36];
    46: op1_00_in15 = reg_0491;
    47: op1_00_in15 = reg_0469;
    48: op1_00_in15 = imem02_in[15:12];
    49: op1_00_in15 = reg_0951;
    50: op1_00_in15 = reg_0395;
    51: op1_00_in15 = imem05_in[103:100];
    52: op1_00_in15 = imem03_in[7:4];
    53: op1_00_in15 = imem03_in[95:92];
    54: op1_00_in15 = imem04_in[47:44];
    55: op1_00_in15 = imem04_in[59:56];
    56: op1_00_in15 = imem06_in[115:112];
    58: op1_00_in15 = reg_0421;
    59: op1_00_in15 = reg_0139;
    60: op1_00_in15 = reg_0467;
    61: op1_00_in15 = reg_0713;
    62: op1_00_in15 = imem01_in[71:68];
    63: op1_00_in15 = reg_0836;
    64: op1_00_in15 = imem05_in[91:88];
    65: op1_00_in15 = imem06_in[47:44];
    66: op1_00_in15 = imem06_in[91:88];
    67: op1_00_in15 = reg_0679;
    69: op1_00_in15 = reg_0905;
    71: op1_00_in15 = reg_0024;
    72: op1_00_in15 = reg_0434;
    73: op1_00_in15 = reg_0351;
    74: op1_00_in15 = reg_0857;
    76: op1_00_in15 = reg_0196;
    77: op1_00_in15 = reg_0191;
    79: op1_00_in15 = reg_0614;
    80: op1_00_in15 = reg_0965;
    83: op1_00_in15 = imem05_in[55:52];
    84: op1_00_in15 = imem03_in[63:60];
    85: op1_00_in15 = reg_0976;
    86: op1_00_in15 = imem07_in[115:112];
    87: op1_00_in15 = reg_0010;
    88: op1_00_in15 = reg_0008;
    89: op1_00_in15 = reg_0002;
    90: op1_00_in15 = reg_0401;
    91: op1_00_in15 = reg_0694;
    92: op1_00_in15 = imem07_in[55:52];
    93: op1_00_in15 = reg_0052;
    95: op1_00_in15 = reg_0750;
    96: op1_00_in15 = imem01_in[67:64];
    97: op1_00_in15 = reg_0480;
    default: op1_00_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv15 = 1;
    6: op1_00_inv15 = 1;
    12: op1_00_inv15 = 1;
    16: op1_00_inv15 = 1;
    18: op1_00_inv15 = 1;
    19: op1_00_inv15 = 1;
    21: op1_00_inv15 = 1;
    24: op1_00_inv15 = 1;
    27: op1_00_inv15 = 1;
    29: op1_00_inv15 = 1;
    30: op1_00_inv15 = 1;
    31: op1_00_inv15 = 1;
    34: op1_00_inv15 = 1;
    35: op1_00_inv15 = 1;
    41: op1_00_inv15 = 1;
    42: op1_00_inv15 = 1;
    45: op1_00_inv15 = 1;
    46: op1_00_inv15 = 1;
    48: op1_00_inv15 = 1;
    52: op1_00_inv15 = 1;
    54: op1_00_inv15 = 1;
    55: op1_00_inv15 = 1;
    56: op1_00_inv15 = 1;
    58: op1_00_inv15 = 1;
    59: op1_00_inv15 = 1;
    60: op1_00_inv15 = 1;
    61: op1_00_inv15 = 1;
    63: op1_00_inv15 = 1;
    65: op1_00_inv15 = 1;
    66: op1_00_inv15 = 1;
    67: op1_00_inv15 = 1;
    68: op1_00_inv15 = 1;
    69: op1_00_inv15 = 1;
    73: op1_00_inv15 = 1;
    74: op1_00_inv15 = 1;
    77: op1_00_inv15 = 1;
    84: op1_00_inv15 = 1;
    85: op1_00_inv15 = 1;
    86: op1_00_inv15 = 1;
    88: op1_00_inv15 = 1;
    90: op1_00_inv15 = 1;
    92: op1_00_inv15 = 1;
    93: op1_00_inv15 = 1;
    94: op1_00_inv15 = 1;
    95: op1_00_inv15 = 1;
    97: op1_00_inv15 = 1;
    default: op1_00_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in16 = reg_0467;
    6: op1_00_in16 = imem05_in[79:76];
    7: op1_00_in16 = imem01_in[123:120];
    8: op1_00_in16 = reg_0068;
    10: op1_00_in16 = imem02_in[19:16];
    11: op1_00_in16 = imem02_in[91:88];
    12: op1_00_in16 = reg_0801;
    13: op1_00_in16 = imem01_in[39:36];
    14: op1_00_in16 = reg_0139;
    15: op1_00_in16 = reg_0203;
    16: op1_00_in16 = reg_1055;
    17: op1_00_in16 = reg_0544;
    18: op1_00_in16 = imem06_in[27:24];
    19: op1_00_in16 = reg_0865;
    20: op1_00_in16 = reg_0752;
    21: op1_00_in16 = reg_1000;
    22: op1_00_in16 = imem07_in[19:16];
    23: op1_00_in16 = imem01_in[47:44];
    24: op1_00_in16 = reg_0951;
    25: op1_00_in16 = imem02_in[75:72];
    94: op1_00_in16 = imem02_in[75:72];
    26: op1_00_in16 = reg_0389;
    27: op1_00_in16 = reg_0214;
    28: op1_00_in16 = reg_1005;
    29: op1_00_in16 = imem07_in[127:124];
    30: op1_00_in16 = imem01_in[19:16];
    31: op1_00_in16 = reg_1009;
    32: op1_00_in16 = reg_0159;
    33: op1_00_in16 = reg_0198;
    34: op1_00_in16 = reg_0786;
    35: op1_00_in16 = imem07_in[67:64];
    36: op1_00_in16 = imem07_in[11:8];
    37: op1_00_in16 = reg_0420;
    38: op1_00_in16 = imem01_in[59:56];
    39: op1_00_in16 = reg_0478;
    40: op1_00_in16 = reg_0083;
    41: op1_00_in16 = reg_0655;
    42: op1_00_in16 = reg_0965;
    44: op1_00_in16 = reg_0191;
    45: op1_00_in16 = imem03_in[51:48];
    46: op1_00_in16 = reg_0257;
    47: op1_00_in16 = reg_0481;
    48: op1_00_in16 = imem02_in[43:40];
    49: op1_00_in16 = reg_0968;
    50: op1_00_in16 = reg_0391;
    51: op1_00_in16 = reg_0962;
    52: op1_00_in16 = imem03_in[27:24];
    53: op1_00_in16 = imem03_in[99:96];
    54: op1_00_in16 = imem04_in[91:88];
    85: op1_00_in16 = imem04_in[91:88];
    55: op1_00_in16 = imem04_in[63:60];
    56: op1_00_in16 = imem06_in[119:116];
    58: op1_00_in16 = reg_0047;
    59: op1_00_in16 = imem06_in[19:16];
    60: op1_00_in16 = reg_0468;
    61: op1_00_in16 = reg_0715;
    62: op1_00_in16 = reg_0918;
    63: op1_00_in16 = reg_0518;
    64: op1_00_in16 = imem05_in[99:96];
    65: op1_00_in16 = imem06_in[87:84];
    66: op1_00_in16 = imem06_in[107:104];
    67: op1_00_in16 = reg_0817;
    68: op1_00_in16 = imem06_in[31:28];
    69: op1_00_in16 = reg_0654;
    70: op1_00_in16 = reg_0483;
    71: op1_00_in16 = reg_0431;
    72: op1_00_in16 = reg_0240;
    73: op1_00_in16 = reg_0754;
    74: op1_00_in16 = reg_0220;
    76: op1_00_in16 = reg_0202;
    77: op1_00_in16 = reg_0209;
    78: op1_00_in16 = reg_0588;
    79: op1_00_in16 = reg_0028;
    80: op1_00_in16 = reg_0490;
    83: op1_00_in16 = imem05_in[59:56];
    84: op1_00_in16 = imem03_in[75:72];
    86: op1_00_in16 = reg_0720;
    87: op1_00_in16 = reg_0625;
    88: op1_00_in16 = reg_0507;
    89: op1_00_in16 = reg_0315;
    90: op1_00_in16 = reg_0432;
    91: op1_00_in16 = reg_1018;
    92: op1_00_in16 = imem07_in[91:88];
    93: op1_00_in16 = reg_0644;
    95: op1_00_in16 = reg_0666;
    96: op1_00_in16 = imem01_in[71:68];
    97: op1_00_in16 = reg_0479;
    default: op1_00_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv16 = 1;
    8: op1_00_inv16 = 1;
    11: op1_00_inv16 = 1;
    12: op1_00_inv16 = 1;
    15: op1_00_inv16 = 1;
    17: op1_00_inv16 = 1;
    19: op1_00_inv16 = 1;
    21: op1_00_inv16 = 1;
    24: op1_00_inv16 = 1;
    27: op1_00_inv16 = 1;
    29: op1_00_inv16 = 1;
    30: op1_00_inv16 = 1;
    31: op1_00_inv16 = 1;
    32: op1_00_inv16 = 1;
    33: op1_00_inv16 = 1;
    35: op1_00_inv16 = 1;
    39: op1_00_inv16 = 1;
    41: op1_00_inv16 = 1;
    45: op1_00_inv16 = 1;
    50: op1_00_inv16 = 1;
    53: op1_00_inv16 = 1;
    55: op1_00_inv16 = 1;
    56: op1_00_inv16 = 1;
    58: op1_00_inv16 = 1;
    60: op1_00_inv16 = 1;
    63: op1_00_inv16 = 1;
    64: op1_00_inv16 = 1;
    65: op1_00_inv16 = 1;
    66: op1_00_inv16 = 1;
    67: op1_00_inv16 = 1;
    70: op1_00_inv16 = 1;
    71: op1_00_inv16 = 1;
    72: op1_00_inv16 = 1;
    73: op1_00_inv16 = 1;
    74: op1_00_inv16 = 1;
    76: op1_00_inv16 = 1;
    78: op1_00_inv16 = 1;
    84: op1_00_inv16 = 1;
    85: op1_00_inv16 = 1;
    86: op1_00_inv16 = 1;
    87: op1_00_inv16 = 1;
    89: op1_00_inv16 = 1;
    90: op1_00_inv16 = 1;
    91: op1_00_inv16 = 1;
    92: op1_00_inv16 = 1;
    94: op1_00_inv16 = 1;
    97: op1_00_inv16 = 1;
    default: op1_00_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in17 = reg_0474;
    6: op1_00_in17 = imem05_in[115:112];
    7: op1_00_in17 = reg_0501;
    8: op1_00_in17 = reg_0074;
    10: op1_00_in17 = imem02_in[27:24];
    11: op1_00_in17 = reg_0658;
    12: op1_00_in17 = reg_0802;
    13: op1_00_in17 = imem01_in[59:56];
    14: op1_00_in17 = reg_0140;
    15: op1_00_in17 = reg_0193;
    16: op1_00_in17 = reg_0511;
    17: op1_00_in17 = reg_0553;
    18: op1_00_in17 = imem06_in[35:32];
    19: op1_00_in17 = reg_0828;
    20: op1_00_in17 = reg_0486;
    21: op1_00_in17 = reg_0994;
    22: op1_00_in17 = imem07_in[27:24];
    23: op1_00_in17 = imem01_in[63:60];
    24: op1_00_in17 = reg_0949;
    25: op1_00_in17 = reg_0666;
    26: op1_00_in17 = reg_0979;
    27: op1_00_in17 = reg_0194;
    28: op1_00_in17 = reg_0778;
    29: op1_00_in17 = reg_0728;
    92: op1_00_in17 = reg_0728;
    30: op1_00_in17 = imem01_in[31:28];
    31: op1_00_in17 = reg_0277;
    32: op1_00_in17 = reg_0173;
    33: op1_00_in17 = reg_0190;
    34: op1_00_in17 = reg_0224;
    35: op1_00_in17 = imem07_in[87:84];
    36: op1_00_in17 = imem07_in[15:12];
    37: op1_00_in17 = reg_0162;
    38: op1_00_in17 = reg_0218;
    39: op1_00_in17 = reg_0189;
    40: op1_00_in17 = reg_0482;
    41: op1_00_in17 = reg_0653;
    42: op1_00_in17 = reg_0947;
    44: op1_00_in17 = reg_0206;
    45: op1_00_in17 = imem03_in[63:60];
    46: op1_00_in17 = reg_0138;
    47: op1_00_in17 = reg_0468;
    48: op1_00_in17 = imem02_in[51:48];
    49: op1_00_in17 = reg_0827;
    50: op1_00_in17 = reg_0295;
    90: op1_00_in17 = reg_0295;
    51: op1_00_in17 = reg_0973;
    52: op1_00_in17 = imem03_in[59:56];
    53: op1_00_in17 = reg_1050;
    54: op1_00_in17 = reg_0301;
    55: op1_00_in17 = reg_0539;
    56: op1_00_in17 = reg_0613;
    58: op1_00_in17 = reg_0160;
    59: op1_00_in17 = imem06_in[27:24];
    60: op1_00_in17 = reg_0458;
    61: op1_00_in17 = reg_0718;
    62: op1_00_in17 = reg_0510;
    63: op1_00_in17 = reg_0991;
    64: op1_00_in17 = reg_0941;
    65: op1_00_in17 = imem06_in[103:100];
    66: op1_00_in17 = imem06_in[119:116];
    67: op1_00_in17 = reg_0926;
    68: op1_00_in17 = imem06_in[43:40];
    69: op1_00_in17 = reg_0637;
    70: op1_00_in17 = reg_1003;
    71: op1_00_in17 = reg_0164;
    72: op1_00_in17 = reg_0576;
    73: op1_00_in17 = reg_0384;
    74: op1_00_in17 = reg_0369;
    76: op1_00_in17 = reg_0199;
    77: op1_00_in17 = reg_0201;
    78: op1_00_in17 = reg_0987;
    79: op1_00_in17 = reg_0392;
    80: op1_00_in17 = imem06_in[19:16];
    83: op1_00_in17 = imem05_in[71:68];
    84: op1_00_in17 = imem03_in[91:88];
    85: op1_00_in17 = reg_0405;
    86: op1_00_in17 = reg_0710;
    87: op1_00_in17 = reg_0344;
    88: op1_00_in17 = reg_0799;
    89: op1_00_in17 = reg_0641;
    91: op1_00_in17 = reg_0626;
    93: op1_00_in17 = reg_0155;
    94: op1_00_in17 = imem02_in[79:76];
    95: op1_00_in17 = reg_0285;
    96: op1_00_in17 = imem01_in[103:100];
    97: op1_00_in17 = reg_0214;
    default: op1_00_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv17 = 1;
    10: op1_00_inv17 = 1;
    14: op1_00_inv17 = 1;
    17: op1_00_inv17 = 1;
    20: op1_00_inv17 = 1;
    21: op1_00_inv17 = 1;
    28: op1_00_inv17 = 1;
    30: op1_00_inv17 = 1;
    31: op1_00_inv17 = 1;
    32: op1_00_inv17 = 1;
    36: op1_00_inv17 = 1;
    37: op1_00_inv17 = 1;
    39: op1_00_inv17 = 1;
    40: op1_00_inv17 = 1;
    44: op1_00_inv17 = 1;
    49: op1_00_inv17 = 1;
    50: op1_00_inv17 = 1;
    59: op1_00_inv17 = 1;
    60: op1_00_inv17 = 1;
    67: op1_00_inv17 = 1;
    69: op1_00_inv17 = 1;
    70: op1_00_inv17 = 1;
    72: op1_00_inv17 = 1;
    76: op1_00_inv17 = 1;
    77: op1_00_inv17 = 1;
    80: op1_00_inv17 = 1;
    84: op1_00_inv17 = 1;
    85: op1_00_inv17 = 1;
    87: op1_00_inv17 = 1;
    89: op1_00_inv17 = 1;
    90: op1_00_inv17 = 1;
    91: op1_00_inv17 = 1;
    96: op1_00_inv17 = 1;
    97: op1_00_inv17 = 1;
    default: op1_00_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in18 = reg_0452;
    6: op1_00_in18 = imem05_in[127:124];
    7: op1_00_in18 = reg_0522;
    8: op1_00_in18 = reg_0064;
    10: op1_00_in18 = imem02_in[39:36];
    11: op1_00_in18 = reg_0653;
    12: op1_00_in18 = imem07_in[7:4];
    13: op1_00_in18 = imem01_in[75:72];
    14: op1_00_in18 = imem06_in[11:8];
    15: op1_00_in18 = reg_0205;
    16: op1_00_in18 = reg_0735;
    17: op1_00_in18 = reg_0552;
    18: op1_00_in18 = imem06_in[39:36];
    19: op1_00_in18 = reg_0145;
    20: op1_00_in18 = reg_0018;
    21: op1_00_in18 = imem04_in[59:56];
    22: op1_00_in18 = imem07_in[39:36];
    23: op1_00_in18 = imem01_in[79:76];
    24: op1_00_in18 = reg_0968;
    25: op1_00_in18 = reg_0667;
    26: op1_00_in18 = reg_0988;
    63: op1_00_in18 = reg_0988;
    27: op1_00_in18 = reg_0201;
    28: op1_00_in18 = reg_0050;
    29: op1_00_in18 = reg_0731;
    30: op1_00_in18 = imem01_in[35:32];
    31: op1_00_in18 = reg_1020;
    33: op1_00_in18 = imem01_in[51:48];
    34: op1_00_in18 = reg_0555;
    35: op1_00_in18 = reg_0710;
    36: op1_00_in18 = imem07_in[19:16];
    37: op1_00_in18 = reg_0167;
    38: op1_00_in18 = reg_0544;
    39: op1_00_in18 = reg_0193;
    40: op1_00_in18 = reg_0776;
    41: op1_00_in18 = reg_0656;
    42: op1_00_in18 = reg_0972;
    44: op1_00_in18 = reg_0197;
    45: op1_00_in18 = imem03_in[99:96];
    46: op1_00_in18 = reg_0153;
    47: op1_00_in18 = reg_0459;
    48: op1_00_in18 = imem02_in[67:64];
    49: op1_00_in18 = reg_0136;
    50: op1_00_in18 = reg_0804;
    51: op1_00_in18 = reg_0959;
    52: op1_00_in18 = imem03_in[107:104];
    53: op1_00_in18 = reg_1049;
    54: op1_00_in18 = reg_0055;
    55: op1_00_in18 = reg_1057;
    56: op1_00_in18 = reg_0073;
    58: op1_00_in18 = reg_0163;
    59: op1_00_in18 = imem06_in[75:72];
    60: op1_00_in18 = reg_0189;
    61: op1_00_in18 = reg_0701;
    62: op1_00_in18 = reg_1035;
    64: op1_00_in18 = reg_0942;
    65: op1_00_in18 = imem06_in[127:124];
    66: op1_00_in18 = imem06_in[127:124];
    67: op1_00_in18 = reg_0384;
    68: op1_00_in18 = imem06_in[47:44];
    69: op1_00_in18 = reg_0565;
    70: op1_00_in18 = reg_0540;
    71: op1_00_in18 = reg_0170;
    72: op1_00_in18 = reg_0823;
    73: op1_00_in18 = reg_0614;
    74: op1_00_in18 = reg_0573;
    76: op1_00_in18 = imem01_in[23:20];
    77: op1_00_in18 = reg_0190;
    78: op1_00_in18 = reg_0982;
    79: op1_00_in18 = reg_0595;
    80: op1_00_in18 = imem06_in[31:28];
    83: op1_00_in18 = imem05_in[99:96];
    84: op1_00_in18 = imem03_in[103:100];
    85: op1_00_in18 = reg_0390;
    86: op1_00_in18 = reg_0250;
    87: op1_00_in18 = reg_0244;
    88: op1_00_in18 = reg_0076;
    89: op1_00_in18 = reg_0161;
    90: op1_00_in18 = reg_0332;
    91: op1_00_in18 = reg_0926;
    92: op1_00_in18 = reg_0720;
    93: op1_00_in18 = reg_0082;
    94: op1_00_in18 = imem02_in[111:108];
    95: op1_00_in18 = reg_0075;
    96: op1_00_in18 = reg_0869;
    97: op1_00_in18 = reg_0208;
    default: op1_00_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv18 = 1;
    6: op1_00_inv18 = 1;
    8: op1_00_inv18 = 1;
    10: op1_00_inv18 = 1;
    11: op1_00_inv18 = 1;
    12: op1_00_inv18 = 1;
    14: op1_00_inv18 = 1;
    16: op1_00_inv18 = 1;
    22: op1_00_inv18 = 1;
    24: op1_00_inv18 = 1;
    25: op1_00_inv18 = 1;
    28: op1_00_inv18 = 1;
    29: op1_00_inv18 = 1;
    30: op1_00_inv18 = 1;
    31: op1_00_inv18 = 1;
    38: op1_00_inv18 = 1;
    40: op1_00_inv18 = 1;
    41: op1_00_inv18 = 1;
    42: op1_00_inv18 = 1;
    46: op1_00_inv18 = 1;
    47: op1_00_inv18 = 1;
    49: op1_00_inv18 = 1;
    55: op1_00_inv18 = 1;
    56: op1_00_inv18 = 1;
    58: op1_00_inv18 = 1;
    59: op1_00_inv18 = 1;
    61: op1_00_inv18 = 1;
    68: op1_00_inv18 = 1;
    70: op1_00_inv18 = 1;
    72: op1_00_inv18 = 1;
    73: op1_00_inv18 = 1;
    74: op1_00_inv18 = 1;
    76: op1_00_inv18 = 1;
    77: op1_00_inv18 = 1;
    79: op1_00_inv18 = 1;
    83: op1_00_inv18 = 1;
    85: op1_00_inv18 = 1;
    87: op1_00_inv18 = 1;
    88: op1_00_inv18 = 1;
    90: op1_00_inv18 = 1;
    95: op1_00_inv18 = 1;
    default: op1_00_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in19 = reg_0189;
    6: op1_00_in19 = reg_0241;
    7: op1_00_in19 = reg_0520;
    8: op1_00_in19 = imem05_in[15:12];
    10: op1_00_in19 = imem02_in[59:56];
    11: op1_00_in19 = reg_0654;
    12: op1_00_in19 = imem07_in[15:12];
    13: op1_00_in19 = reg_0240;
    14: op1_00_in19 = imem06_in[15:12];
    15: op1_00_in19 = imem01_in[31:28];
    16: op1_00_in19 = reg_0487;
    17: op1_00_in19 = reg_0540;
    18: op1_00_in19 = imem06_in[119:116];
    19: op1_00_in19 = imem06_in[127:124];
    20: op1_00_in19 = reg_0011;
    21: op1_00_in19 = imem04_in[71:68];
    22: op1_00_in19 = imem07_in[43:40];
    23: op1_00_in19 = imem01_in[107:104];
    24: op1_00_in19 = reg_0229;
    25: op1_00_in19 = reg_0352;
    26: op1_00_in19 = imem04_in[23:20];
    27: op1_00_in19 = reg_0206;
    28: op1_00_in19 = reg_0541;
    29: op1_00_in19 = reg_0721;
    35: op1_00_in19 = reg_0721;
    30: op1_00_in19 = imem01_in[83:80];
    31: op1_00_in19 = reg_1005;
    33: op1_00_in19 = imem01_in[63:60];
    34: op1_00_in19 = reg_0274;
    36: op1_00_in19 = imem07_in[67:64];
    37: op1_00_in19 = reg_0163;
    38: op1_00_in19 = reg_1039;
    39: op1_00_in19 = reg_0212;
    40: op1_00_in19 = reg_0091;
    41: op1_00_in19 = reg_0649;
    42: op1_00_in19 = reg_0821;
    44: op1_00_in19 = imem01_in[59:56];
    45: op1_00_in19 = imem03_in[103:100];
    46: op1_00_in19 = imem06_in[39:36];
    80: op1_00_in19 = imem06_in[39:36];
    47: op1_00_in19 = reg_0458;
    48: op1_00_in19 = imem02_in[83:80];
    49: op1_00_in19 = reg_0133;
    50: op1_00_in19 = reg_0349;
    51: op1_00_in19 = reg_0946;
    52: op1_00_in19 = reg_0006;
    53: op1_00_in19 = reg_0327;
    54: op1_00_in19 = reg_1020;
    55: op1_00_in19 = reg_0888;
    56: op1_00_in19 = reg_0759;
    58: op1_00_in19 = reg_0166;
    59: op1_00_in19 = imem06_in[103:100];
    60: op1_00_in19 = reg_0194;
    61: op1_00_in19 = reg_0706;
    62: op1_00_in19 = reg_0285;
    63: op1_00_in19 = reg_0976;
    64: op1_00_in19 = reg_0947;
    65: op1_00_in19 = reg_0660;
    66: op1_00_in19 = reg_0694;
    67: op1_00_in19 = reg_1030;
    68: op1_00_in19 = imem06_in[91:88];
    69: op1_00_in19 = reg_0887;
    70: op1_00_in19 = reg_0931;
    72: op1_00_in19 = reg_0609;
    73: op1_00_in19 = reg_0297;
    74: op1_00_in19 = reg_0566;
    76: op1_00_in19 = imem01_in[35:32];
    77: op1_00_in19 = reg_0199;
    78: op1_00_in19 = reg_0979;
    79: op1_00_in19 = reg_0699;
    83: op1_00_in19 = imem05_in[103:100];
    84: op1_00_in19 = reg_0060;
    85: op1_00_in19 = reg_0031;
    86: op1_00_in19 = reg_0315;
    87: op1_00_in19 = reg_0294;
    88: op1_00_in19 = reg_0815;
    89: op1_00_in19 = reg_0703;
    90: op1_00_in19 = imem05_in[47:44];
    91: op1_00_in19 = reg_0889;
    92: op1_00_in19 = reg_0221;
    93: op1_00_in19 = reg_0624;
    94: op1_00_in19 = imem02_in[119:116];
    95: op1_00_in19 = reg_0543;
    96: op1_00_in19 = reg_0594;
    97: op1_00_in19 = reg_0210;
    default: op1_00_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_00_inv19 = 1;
    11: op1_00_inv19 = 1;
    15: op1_00_inv19 = 1;
    18: op1_00_inv19 = 1;
    19: op1_00_inv19 = 1;
    22: op1_00_inv19 = 1;
    23: op1_00_inv19 = 1;
    26: op1_00_inv19 = 1;
    30: op1_00_inv19 = 1;
    36: op1_00_inv19 = 1;
    41: op1_00_inv19 = 1;
    44: op1_00_inv19 = 1;
    45: op1_00_inv19 = 1;
    46: op1_00_inv19 = 1;
    47: op1_00_inv19 = 1;
    54: op1_00_inv19 = 1;
    56: op1_00_inv19 = 1;
    58: op1_00_inv19 = 1;
    67: op1_00_inv19 = 1;
    72: op1_00_inv19 = 1;
    77: op1_00_inv19 = 1;
    80: op1_00_inv19 = 1;
    85: op1_00_inv19 = 1;
    87: op1_00_inv19 = 1;
    88: op1_00_inv19 = 1;
    89: op1_00_inv19 = 1;
    90: op1_00_inv19 = 1;
    94: op1_00_inv19 = 1;
    95: op1_00_inv19 = 1;
    96: op1_00_inv19 = 1;
    default: op1_00_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in20 = reg_0207;
    6: op1_00_in20 = reg_0264;
    7: op1_00_in20 = reg_0499;
    8: op1_00_in20 = imem05_in[23:20];
    10: op1_00_in20 = imem02_in[103:100];
    48: op1_00_in20 = imem02_in[103:100];
    11: op1_00_in20 = reg_0664;
    12: op1_00_in20 = imem07_in[75:72];
    13: op1_00_in20 = reg_0502;
    14: op1_00_in20 = imem06_in[71:68];
    15: op1_00_in20 = imem01_in[75:72];
    16: op1_00_in20 = reg_0245;
    17: op1_00_in20 = reg_0532;
    18: op1_00_in20 = reg_0368;
    19: op1_00_in20 = reg_0617;
    20: op1_00_in20 = reg_0798;
    21: op1_00_in20 = imem04_in[83:80];
    22: op1_00_in20 = imem07_in[59:56];
    23: op1_00_in20 = reg_1055;
    24: op1_00_in20 = reg_0832;
    25: op1_00_in20 = reg_0357;
    26: op1_00_in20 = imem04_in[59:56];
    27: op1_00_in20 = reg_0192;
    28: op1_00_in20 = reg_0313;
    29: op1_00_in20 = reg_0725;
    30: op1_00_in20 = imem01_in[87:84];
    31: op1_00_in20 = reg_0932;
    33: op1_00_in20 = imem01_in[95:92];
    34: op1_00_in20 = reg_0544;
    35: op1_00_in20 = reg_0715;
    36: op1_00_in20 = imem07_in[79:76];
    37: op1_00_in20 = reg_0164;
    38: op1_00_in20 = reg_0226;
    39: op1_00_in20 = reg_0205;
    40: op1_00_in20 = reg_0484;
    41: op1_00_in20 = reg_0665;
    42: op1_00_in20 = reg_0251;
    44: op1_00_in20 = imem01_in[115:112];
    45: op1_00_in20 = reg_1007;
    46: op1_00_in20 = imem06_in[43:40];
    47: op1_00_in20 = reg_0198;
    49: op1_00_in20 = reg_0154;
    50: op1_00_in20 = reg_0222;
    51: op1_00_in20 = reg_0953;
    52: op1_00_in20 = reg_0317;
    53: op1_00_in20 = reg_0046;
    54: op1_00_in20 = reg_1005;
    55: op1_00_in20 = reg_0931;
    56: op1_00_in20 = reg_0220;
    58: op1_00_in20 = reg_0157;
    59: op1_00_in20 = imem06_in[111:108];
    60: op1_00_in20 = imem01_in[3:0];
    61: op1_00_in20 = reg_0361;
    62: op1_00_in20 = reg_0249;
    63: op1_00_in20 = imem04_in[3:0];
    64: op1_00_in20 = reg_0032;
    65: op1_00_in20 = reg_1019;
    66: op1_00_in20 = reg_0626;
    67: op1_00_in20 = reg_0440;
    68: op1_00_in20 = imem06_in[127:124];
    69: op1_00_in20 = reg_0336;
    70: op1_00_in20 = reg_0076;
    72: op1_00_in20 = reg_0581;
    73: op1_00_in20 = reg_0698;
    74: op1_00_in20 = imem07_in[15:12];
    76: op1_00_in20 = imem01_in[63:60];
    77: op1_00_in20 = imem01_in[43:40];
    78: op1_00_in20 = reg_0993;
    79: op1_00_in20 = reg_0921;
    80: op1_00_in20 = imem06_in[83:80];
    83: op1_00_in20 = imem05_in[123:120];
    84: op1_00_in20 = reg_0012;
    85: op1_00_in20 = reg_0016;
    86: op1_00_in20 = reg_0406;
    87: op1_00_in20 = reg_0391;
    88: op1_00_in20 = reg_0494;
    89: op1_00_in20 = reg_0183;
    90: op1_00_in20 = imem05_in[55:52];
    91: op1_00_in20 = reg_0692;
    92: op1_00_in20 = reg_0710;
    93: op1_00_in20 = imem03_in[3:0];
    94: op1_00_in20 = reg_0916;
    95: op1_00_in20 = reg_0637;
    96: op1_00_in20 = reg_0591;
    97: op1_00_in20 = reg_0209;
    default: op1_00_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv20 = 1;
    6: op1_00_inv20 = 1;
    10: op1_00_inv20 = 1;
    12: op1_00_inv20 = 1;
    16: op1_00_inv20 = 1;
    20: op1_00_inv20 = 1;
    21: op1_00_inv20 = 1;
    24: op1_00_inv20 = 1;
    25: op1_00_inv20 = 1;
    28: op1_00_inv20 = 1;
    30: op1_00_inv20 = 1;
    34: op1_00_inv20 = 1;
    35: op1_00_inv20 = 1;
    36: op1_00_inv20 = 1;
    37: op1_00_inv20 = 1;
    39: op1_00_inv20 = 1;
    42: op1_00_inv20 = 1;
    44: op1_00_inv20 = 1;
    45: op1_00_inv20 = 1;
    46: op1_00_inv20 = 1;
    48: op1_00_inv20 = 1;
    54: op1_00_inv20 = 1;
    58: op1_00_inv20 = 1;
    59: op1_00_inv20 = 1;
    60: op1_00_inv20 = 1;
    65: op1_00_inv20 = 1;
    68: op1_00_inv20 = 1;
    69: op1_00_inv20 = 1;
    70: op1_00_inv20 = 1;
    74: op1_00_inv20 = 1;
    78: op1_00_inv20 = 1;
    83: op1_00_inv20 = 1;
    84: op1_00_inv20 = 1;
    85: op1_00_inv20 = 1;
    87: op1_00_inv20 = 1;
    88: op1_00_inv20 = 1;
    90: op1_00_inv20 = 1;
    91: op1_00_inv20 = 1;
    95: op1_00_inv20 = 1;
    97: op1_00_inv20 = 1;
    default: op1_00_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in21 = reg_0194;
    6: op1_00_in21 = reg_0265;
    7: op1_00_in21 = reg_0498;
    8: op1_00_in21 = imem05_in[27:24];
    10: op1_00_in21 = imem02_in[119:116];
    11: op1_00_in21 = reg_0660;
    12: op1_00_in21 = imem07_in[99:96];
    13: op1_00_in21 = reg_0247;
    14: op1_00_in21 = imem06_in[99:96];
    15: op1_00_in21 = imem01_in[83:80];
    16: op1_00_in21 = reg_1032;
    17: op1_00_in21 = reg_0559;
    18: op1_00_in21 = reg_0787;
    19: op1_00_in21 = reg_0618;
    20: op1_00_in21 = imem07_in[31:28];
    21: op1_00_in21 = imem04_in[87:84];
    22: op1_00_in21 = imem07_in[107:104];
    23: op1_00_in21 = reg_0240;
    24: op1_00_in21 = reg_0819;
    25: op1_00_in21 = reg_0358;
    26: op1_00_in21 = imem04_in[71:68];
    27: op1_00_in21 = imem01_in[63:60];
    28: op1_00_in21 = reg_0763;
    29: op1_00_in21 = reg_0709;
    30: op1_00_in21 = imem01_in[99:96];
    76: op1_00_in21 = imem01_in[99:96];
    31: op1_00_in21 = reg_0078;
    33: op1_00_in21 = reg_0563;
    34: op1_00_in21 = reg_0487;
    35: op1_00_in21 = reg_0700;
    36: op1_00_in21 = reg_0712;
    37: op1_00_in21 = reg_0170;
    38: op1_00_in21 = reg_1042;
    39: op1_00_in21 = reg_0202;
    40: op1_00_in21 = imem03_in[7:4];
    41: op1_00_in21 = reg_0225;
    42: op1_00_in21 = reg_0257;
    44: op1_00_in21 = reg_0786;
    45: op1_00_in21 = reg_0327;
    46: op1_00_in21 = imem06_in[63:60];
    47: op1_00_in21 = reg_0201;
    48: op1_00_in21 = imem02_in[107:104];
    49: op1_00_in21 = reg_0143;
    50: op1_00_in21 = reg_0380;
    51: op1_00_in21 = reg_0215;
    52: op1_00_in21 = reg_1019;
    53: op1_00_in21 = reg_0396;
    54: op1_00_in21 = reg_0540;
    55: op1_00_in21 = reg_0568;
    56: op1_00_in21 = reg_0395;
    58: op1_00_in21 = reg_0176;
    59: op1_00_in21 = reg_0344;
    60: op1_00_in21 = imem01_in[27:24];
    61: op1_00_in21 = reg_0532;
    62: op1_00_in21 = reg_0869;
    63: op1_00_in21 = imem04_in[15:12];
    64: op1_00_in21 = reg_0446;
    65: op1_00_in21 = reg_0691;
    66: op1_00_in21 = reg_0679;
    67: op1_00_in21 = reg_0895;
    68: op1_00_in21 = reg_0080;
    69: op1_00_in21 = reg_0837;
    70: op1_00_in21 = reg_0584;
    72: op1_00_in21 = reg_1001;
    73: op1_00_in21 = reg_0591;
    74: op1_00_in21 = imem07_in[43:40];
    77: op1_00_in21 = imem01_in[75:72];
    78: op1_00_in21 = reg_0980;
    79: op1_00_in21 = reg_0807;
    80: op1_00_in21 = imem06_in[87:84];
    83: op1_00_in21 = imem05_in[127:124];
    84: op1_00_in21 = reg_1007;
    85: op1_00_in21 = reg_0802;
    86: op1_00_in21 = reg_0640;
    87: op1_00_in21 = reg_0817;
    88: op1_00_in21 = imem05_in[3:0];
    89: op1_00_in21 = reg_0724;
    90: op1_00_in21 = imem05_in[63:60];
    91: op1_00_in21 = reg_0792;
    92: op1_00_in21 = reg_0721;
    93: op1_00_in21 = imem03_in[31:28];
    94: op1_00_in21 = reg_0605;
    95: op1_00_in21 = reg_0349;
    96: op1_00_in21 = reg_0769;
    97: op1_00_in21 = reg_0207;
    default: op1_00_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv21 = 1;
    13: op1_00_inv21 = 1;
    16: op1_00_inv21 = 1;
    17: op1_00_inv21 = 1;
    18: op1_00_inv21 = 1;
    22: op1_00_inv21 = 1;
    23: op1_00_inv21 = 1;
    24: op1_00_inv21 = 1;
    26: op1_00_inv21 = 1;
    29: op1_00_inv21 = 1;
    34: op1_00_inv21 = 1;
    35: op1_00_inv21 = 1;
    36: op1_00_inv21 = 1;
    37: op1_00_inv21 = 1;
    38: op1_00_inv21 = 1;
    39: op1_00_inv21 = 1;
    40: op1_00_inv21 = 1;
    41: op1_00_inv21 = 1;
    42: op1_00_inv21 = 1;
    44: op1_00_inv21 = 1;
    45: op1_00_inv21 = 1;
    46: op1_00_inv21 = 1;
    47: op1_00_inv21 = 1;
    48: op1_00_inv21 = 1;
    51: op1_00_inv21 = 1;
    55: op1_00_inv21 = 1;
    56: op1_00_inv21 = 1;
    58: op1_00_inv21 = 1;
    59: op1_00_inv21 = 1;
    60: op1_00_inv21 = 1;
    62: op1_00_inv21 = 1;
    63: op1_00_inv21 = 1;
    65: op1_00_inv21 = 1;
    66: op1_00_inv21 = 1;
    68: op1_00_inv21 = 1;
    69: op1_00_inv21 = 1;
    70: op1_00_inv21 = 1;
    76: op1_00_inv21 = 1;
    78: op1_00_inv21 = 1;
    79: op1_00_inv21 = 1;
    80: op1_00_inv21 = 1;
    84: op1_00_inv21 = 1;
    85: op1_00_inv21 = 1;
    86: op1_00_inv21 = 1;
    87: op1_00_inv21 = 1;
    89: op1_00_inv21 = 1;
    90: op1_00_inv21 = 1;
    93: op1_00_inv21 = 1;
    94: op1_00_inv21 = 1;
    95: op1_00_inv21 = 1;
    default: op1_00_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in22 = reg_0201;
    6: op1_00_in22 = reg_0266;
    7: op1_00_in22 = reg_0218;
    8: op1_00_in22 = imem05_in[63:60];
    10: op1_00_in22 = reg_0666;
    11: op1_00_in22 = reg_0639;
    12: op1_00_in22 = reg_0704;
    22: op1_00_in22 = reg_0704;
    13: op1_00_in22 = reg_0503;
    14: op1_00_in22 = imem06_in[115:112];
    15: op1_00_in22 = imem01_in[103:100];
    16: op1_00_in22 = reg_0216;
    17: op1_00_in22 = reg_0556;
    18: op1_00_in22 = reg_0808;
    19: op1_00_in22 = reg_0627;
    20: op1_00_in22 = imem07_in[39:36];
    21: op1_00_in22 = imem04_in[99:96];
    23: op1_00_in22 = reg_0247;
    24: op1_00_in22 = reg_0128;
    25: op1_00_in22 = reg_0354;
    26: op1_00_in22 = imem04_in[79:76];
    27: op1_00_in22 = imem01_in[71:68];
    28: op1_00_in22 = reg_0760;
    29: op1_00_in22 = reg_0718;
    30: op1_00_in22 = imem01_in[127:124];
    31: op1_00_in22 = reg_0067;
    33: op1_00_in22 = reg_0003;
    34: op1_00_in22 = reg_0087;
    35: op1_00_in22 = reg_0436;
    36: op1_00_in22 = reg_0729;
    38: op1_00_in22 = reg_0496;
    39: op1_00_in22 = imem01_in[7:4];
    40: op1_00_in22 = imem03_in[15:12];
    41: op1_00_in22 = reg_0330;
    42: op1_00_in22 = reg_0132;
    44: op1_00_in22 = reg_0779;
    45: op1_00_in22 = reg_0046;
    46: op1_00_in22 = imem06_in[67:64];
    47: op1_00_in22 = reg_0196;
    48: op1_00_in22 = reg_0363;
    49: op1_00_in22 = imem06_in[51:48];
    50: op1_00_in22 = reg_0332;
    51: op1_00_in22 = reg_0508;
    52: op1_00_in22 = reg_0245;
    53: op1_00_in22 = reg_0795;
    54: op1_00_in22 = reg_0050;
    55: op1_00_in22 = reg_0816;
    56: op1_00_in22 = reg_0741;
    58: op1_00_in22 = reg_0158;
    59: op1_00_in22 = reg_0244;
    60: op1_00_in22 = imem01_in[59:56];
    61: op1_00_in22 = reg_0160;
    62: op1_00_in22 = reg_0514;
    63: op1_00_in22 = imem04_in[71:68];
    64: op1_00_in22 = reg_1046;
    65: op1_00_in22 = reg_0267;
    66: op1_00_in22 = reg_0021;
    67: op1_00_in22 = reg_0439;
    68: op1_00_in22 = reg_0297;
    69: op1_00_in22 = reg_0818;
    70: op1_00_in22 = reg_0732;
    72: op1_00_in22 = reg_0978;
    73: op1_00_in22 = reg_0863;
    74: op1_00_in22 = imem07_in[75:72];
    76: op1_00_in22 = imem01_in[115:112];
    77: op1_00_in22 = imem01_in[115:112];
    78: op1_00_in22 = imem04_in[3:0];
    79: op1_00_in22 = reg_0220;
    80: op1_00_in22 = reg_1019;
    83: op1_00_in22 = reg_1021;
    84: op1_00_in22 = reg_0445;
    85: op1_00_in22 = reg_0568;
    86: op1_00_in22 = reg_0181;
    87: op1_00_in22 = reg_0754;
    88: op1_00_in22 = imem05_in[23:20];
    90: op1_00_in22 = imem05_in[75:72];
    91: op1_00_in22 = reg_0822;
    92: op1_00_in22 = reg_0717;
    93: op1_00_in22 = imem03_in[43:40];
    94: op1_00_in22 = reg_0091;
    95: op1_00_in22 = reg_0739;
    96: op1_00_in22 = reg_0112;
    97: op1_00_in22 = reg_0211;
    default: op1_00_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_00_inv22 = 1;
    8: op1_00_inv22 = 1;
    10: op1_00_inv22 = 1;
    12: op1_00_inv22 = 1;
    13: op1_00_inv22 = 1;
    15: op1_00_inv22 = 1;
    16: op1_00_inv22 = 1;
    17: op1_00_inv22 = 1;
    18: op1_00_inv22 = 1;
    20: op1_00_inv22 = 1;
    22: op1_00_inv22 = 1;
    23: op1_00_inv22 = 1;
    25: op1_00_inv22 = 1;
    28: op1_00_inv22 = 1;
    29: op1_00_inv22 = 1;
    30: op1_00_inv22 = 1;
    33: op1_00_inv22 = 1;
    34: op1_00_inv22 = 1;
    36: op1_00_inv22 = 1;
    38: op1_00_inv22 = 1;
    40: op1_00_inv22 = 1;
    41: op1_00_inv22 = 1;
    49: op1_00_inv22 = 1;
    51: op1_00_inv22 = 1;
    55: op1_00_inv22 = 1;
    56: op1_00_inv22 = 1;
    58: op1_00_inv22 = 1;
    59: op1_00_inv22 = 1;
    60: op1_00_inv22 = 1;
    61: op1_00_inv22 = 1;
    63: op1_00_inv22 = 1;
    64: op1_00_inv22 = 1;
    65: op1_00_inv22 = 1;
    72: op1_00_inv22 = 1;
    73: op1_00_inv22 = 1;
    76: op1_00_inv22 = 1;
    79: op1_00_inv22 = 1;
    80: op1_00_inv22 = 1;
    83: op1_00_inv22 = 1;
    85: op1_00_inv22 = 1;
    86: op1_00_inv22 = 1;
    87: op1_00_inv22 = 1;
    88: op1_00_inv22 = 1;
    90: op1_00_inv22 = 1;
    91: op1_00_inv22 = 1;
    92: op1_00_inv22 = 1;
    93: op1_00_inv22 = 1;
    94: op1_00_inv22 = 1;
    96: op1_00_inv22 = 1;
    97: op1_00_inv22 = 1;
    default: op1_00_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in23 = reg_0190;
    6: op1_00_in23 = reg_0139;
    7: op1_00_in23 = reg_0219;
    8: op1_00_in23 = imem05_in[75:72];
    10: op1_00_in23 = reg_0653;
    11: op1_00_in23 = reg_0640;
    12: op1_00_in23 = reg_0723;
    13: op1_00_in23 = reg_0248;
    14: op1_00_in23 = reg_0628;
    15: op1_00_in23 = imem01_in[107:104];
    16: op1_00_in23 = reg_1036;
    38: op1_00_in23 = reg_1036;
    17: op1_00_in23 = reg_0294;
    18: op1_00_in23 = reg_1028;
    19: op1_00_in23 = reg_0622;
    20: op1_00_in23 = imem07_in[83:80];
    74: op1_00_in23 = imem07_in[83:80];
    21: op1_00_in23 = imem04_in[107:104];
    22: op1_00_in23 = reg_0703;
    23: op1_00_in23 = reg_0503;
    24: op1_00_in23 = reg_0130;
    25: op1_00_in23 = reg_0346;
    45: op1_00_in23 = reg_0346;
    26: op1_00_in23 = reg_0530;
    27: op1_00_in23 = imem01_in[87:84];
    28: op1_00_in23 = reg_0009;
    29: op1_00_in23 = reg_0421;
    30: op1_00_in23 = reg_0013;
    31: op1_00_in23 = reg_0259;
    33: op1_00_in23 = reg_0299;
    34: op1_00_in23 = reg_0496;
    35: op1_00_in23 = reg_0418;
    36: op1_00_in23 = reg_0715;
    39: op1_00_in23 = imem01_in[23:20];
    40: op1_00_in23 = imem03_in[47:44];
    41: op1_00_in23 = reg_0007;
    42: op1_00_in23 = reg_0145;
    44: op1_00_in23 = reg_0274;
    46: op1_00_in23 = reg_0892;
    47: op1_00_in23 = reg_0195;
    48: op1_00_in23 = reg_0082;
    49: op1_00_in23 = imem06_in[63:60];
    50: op1_00_in23 = reg_0629;
    51: op1_00_in23 = reg_0813;
    52: op1_00_in23 = reg_0397;
    53: op1_00_in23 = reg_0509;
    54: op1_00_in23 = reg_0313;
    55: op1_00_in23 = reg_0027;
    56: op1_00_in23 = reg_0382;
    58: op1_00_in23 = reg_0173;
    59: op1_00_in23 = reg_0328;
    66: op1_00_in23 = reg_0328;
    60: op1_00_in23 = imem01_in[75:72];
    61: op1_00_in23 = reg_0166;
    62: op1_00_in23 = reg_0830;
    63: op1_00_in23 = imem04_in[79:76];
    64: op1_00_in23 = reg_0447;
    65: op1_00_in23 = reg_0262;
    67: op1_00_in23 = reg_0804;
    68: op1_00_in23 = reg_0895;
    69: op1_00_in23 = reg_0776;
    70: op1_00_in23 = reg_0284;
    72: op1_00_in23 = reg_0974;
    73: op1_00_in23 = reg_0917;
    76: op1_00_in23 = reg_0106;
    77: op1_00_in23 = imem01_in[119:116];
    78: op1_00_in23 = imem04_in[35:32];
    79: op1_00_in23 = reg_0915;
    80: op1_00_in23 = reg_0021;
    83: op1_00_in23 = reg_0215;
    84: op1_00_in23 = reg_0585;
    85: op1_00_in23 = reg_0296;
    86: op1_00_in23 = reg_0714;
    87: op1_00_in23 = reg_0735;
    88: op1_00_in23 = imem05_in[31:28];
    90: op1_00_in23 = imem05_in[91:88];
    91: op1_00_in23 = reg_0121;
    92: op1_00_in23 = reg_0515;
    93: op1_00_in23 = imem03_in[67:64];
    94: op1_00_in23 = reg_0348;
    95: op1_00_in23 = reg_0664;
    96: op1_00_in23 = reg_0114;
    97: op1_00_in23 = reg_0213;
    default: op1_00_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    13: op1_00_inv23 = 1;
    16: op1_00_inv23 = 1;
    17: op1_00_inv23 = 1;
    20: op1_00_inv23 = 1;
    23: op1_00_inv23 = 1;
    24: op1_00_inv23 = 1;
    25: op1_00_inv23 = 1;
    29: op1_00_inv23 = 1;
    35: op1_00_inv23 = 1;
    36: op1_00_inv23 = 1;
    41: op1_00_inv23 = 1;
    44: op1_00_inv23 = 1;
    49: op1_00_inv23 = 1;
    51: op1_00_inv23 = 1;
    52: op1_00_inv23 = 1;
    53: op1_00_inv23 = 1;
    54: op1_00_inv23 = 1;
    56: op1_00_inv23 = 1;
    58: op1_00_inv23 = 1;
    59: op1_00_inv23 = 1;
    62: op1_00_inv23 = 1;
    63: op1_00_inv23 = 1;
    65: op1_00_inv23 = 1;
    67: op1_00_inv23 = 1;
    68: op1_00_inv23 = 1;
    70: op1_00_inv23 = 1;
    74: op1_00_inv23 = 1;
    76: op1_00_inv23 = 1;
    77: op1_00_inv23 = 1;
    80: op1_00_inv23 = 1;
    83: op1_00_inv23 = 1;
    84: op1_00_inv23 = 1;
    86: op1_00_inv23 = 1;
    91: op1_00_inv23 = 1;
    92: op1_00_inv23 = 1;
    95: op1_00_inv23 = 1;
    96: op1_00_inv23 = 1;
    97: op1_00_inv23 = 1;
    default: op1_00_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in24 = reg_0202;
    6: op1_00_in24 = imem06_in[3:0];
    7: op1_00_in24 = reg_0123;
    8: op1_00_in24 = imem05_in[99:96];
    10: op1_00_in24 = reg_0664;
    11: op1_00_in24 = reg_0662;
    12: op1_00_in24 = reg_0425;
    13: op1_00_in24 = reg_0905;
    14: op1_00_in24 = reg_0625;
    15: op1_00_in24 = reg_1051;
    16: op1_00_in24 = reg_1015;
    17: op1_00_in24 = reg_0297;
    59: op1_00_in24 = reg_0297;
    66: op1_00_in24 = reg_0297;
    18: op1_00_in24 = reg_0005;
    19: op1_00_in24 = reg_0392;
    20: op1_00_in24 = imem07_in[103:100];
    21: op1_00_in24 = imem04_in[115:112];
    22: op1_00_in24 = reg_0712;
    23: op1_00_in24 = reg_0248;
    24: op1_00_in24 = reg_0131;
    25: op1_00_in24 = reg_0347;
    26: op1_00_in24 = reg_0265;
    27: op1_00_in24 = reg_0235;
    28: op1_00_in24 = reg_0738;
    29: op1_00_in24 = reg_0440;
    30: op1_00_in24 = reg_0223;
    31: op1_00_in24 = reg_0276;
    33: op1_00_in24 = reg_0810;
    34: op1_00_in24 = reg_1033;
    35: op1_00_in24 = reg_0419;
    36: op1_00_in24 = reg_0441;
    38: op1_00_in24 = reg_1038;
    39: op1_00_in24 = imem01_in[43:40];
    97: op1_00_in24 = imem01_in[43:40];
    40: op1_00_in24 = imem03_in[127:124];
    41: op1_00_in24 = reg_0506;
    42: op1_00_in24 = reg_0154;
    44: op1_00_in24 = reg_0544;
    45: op1_00_in24 = reg_0833;
    46: op1_00_in24 = reg_0403;
    47: op1_00_in24 = imem01_in[7:4];
    48: op1_00_in24 = reg_0637;
    49: op1_00_in24 = imem06_in[71:68];
    50: op1_00_in24 = reg_0630;
    51: op1_00_in24 = reg_0336;
    52: op1_00_in24 = reg_0874;
    53: op1_00_in24 = reg_0051;
    54: op1_00_in24 = reg_0507;
    55: op1_00_in24 = reg_0777;
    56: op1_00_in24 = reg_0380;
    60: op1_00_in24 = imem01_in[107:104];
    61: op1_00_in24 = reg_0157;
    62: op1_00_in24 = reg_1037;
    63: op1_00_in24 = imem04_in[87:84];
    64: op1_00_in24 = reg_0489;
    65: op1_00_in24 = reg_0229;
    67: op1_00_in24 = reg_0699;
    68: op1_00_in24 = reg_0008;
    69: op1_00_in24 = reg_0867;
    70: op1_00_in24 = reg_0764;
    72: op1_00_in24 = reg_0983;
    73: op1_00_in24 = reg_0857;
    74: op1_00_in24 = reg_0728;
    76: op1_00_in24 = reg_0968;
    77: op1_00_in24 = reg_0969;
    78: op1_00_in24 = imem04_in[103:100];
    79: op1_00_in24 = reg_0755;
    80: op1_00_in24 = reg_0817;
    83: op1_00_in24 = reg_0866;
    84: op1_00_in24 = reg_0434;
    85: op1_00_in24 = reg_0288;
    86: op1_00_in24 = reg_0185;
    87: op1_00_in24 = reg_0692;
    88: op1_00_in24 = imem05_in[55:52];
    90: op1_00_in24 = imem05_in[111:108];
    91: op1_00_in24 = reg_0781;
    92: op1_00_in24 = reg_0653;
    93: op1_00_in24 = imem03_in[75:72];
    94: op1_00_in24 = reg_0077;
    95: op1_00_in24 = reg_0052;
    96: op1_00_in24 = reg_0821;
    default: op1_00_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_00_inv24 = 1;
    10: op1_00_inv24 = 1;
    11: op1_00_inv24 = 1;
    14: op1_00_inv24 = 1;
    15: op1_00_inv24 = 1;
    20: op1_00_inv24 = 1;
    21: op1_00_inv24 = 1;
    22: op1_00_inv24 = 1;
    23: op1_00_inv24 = 1;
    24: op1_00_inv24 = 1;
    25: op1_00_inv24 = 1;
    26: op1_00_inv24 = 1;
    28: op1_00_inv24 = 1;
    30: op1_00_inv24 = 1;
    31: op1_00_inv24 = 1;
    34: op1_00_inv24 = 1;
    35: op1_00_inv24 = 1;
    39: op1_00_inv24 = 1;
    40: op1_00_inv24 = 1;
    41: op1_00_inv24 = 1;
    44: op1_00_inv24 = 1;
    48: op1_00_inv24 = 1;
    49: op1_00_inv24 = 1;
    51: op1_00_inv24 = 1;
    53: op1_00_inv24 = 1;
    54: op1_00_inv24 = 1;
    55: op1_00_inv24 = 1;
    61: op1_00_inv24 = 1;
    62: op1_00_inv24 = 1;
    64: op1_00_inv24 = 1;
    66: op1_00_inv24 = 1;
    67: op1_00_inv24 = 1;
    68: op1_00_inv24 = 1;
    69: op1_00_inv24 = 1;
    72: op1_00_inv24 = 1;
    73: op1_00_inv24 = 1;
    78: op1_00_inv24 = 1;
    80: op1_00_inv24 = 1;
    85: op1_00_inv24 = 1;
    87: op1_00_inv24 = 1;
    88: op1_00_inv24 = 1;
    91: op1_00_inv24 = 1;
    92: op1_00_inv24 = 1;
    97: op1_00_inv24 = 1;
    default: op1_00_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in25 = reg_0195;
    6: op1_00_in25 = imem06_in[7:4];
    7: op1_00_in25 = imem02_in[39:36];
    8: op1_00_in25 = imem05_in[107:104];
    10: op1_00_in25 = reg_0657;
    11: op1_00_in25 = reg_0665;
    12: op1_00_in25 = reg_0441;
    13: op1_00_in25 = reg_0496;
    14: op1_00_in25 = reg_0616;
    15: op1_00_in25 = reg_0735;
    16: op1_00_in25 = reg_0871;
    17: op1_00_in25 = reg_0295;
    18: op1_00_in25 = imem07_in[63:60];
    19: op1_00_in25 = reg_0383;
    20: op1_00_in25 = imem07_in[107:104];
    21: op1_00_in25 = reg_0544;
    22: op1_00_in25 = reg_0706;
    23: op1_00_in25 = reg_1052;
    24: op1_00_in25 = imem06_in[15:12];
    25: op1_00_in25 = reg_0007;
    26: op1_00_in25 = reg_0277;
    27: op1_00_in25 = reg_0223;
    28: op1_00_in25 = reg_0875;
    29: op1_00_in25 = reg_0435;
    30: op1_00_in25 = reg_0510;
    31: op1_00_in25 = reg_0064;
    33: op1_00_in25 = reg_0828;
    34: op1_00_in25 = reg_1037;
    35: op1_00_in25 = reg_0439;
    36: op1_00_in25 = reg_0445;
    38: op1_00_in25 = reg_0904;
    39: op1_00_in25 = imem01_in[47:44];
    40: op1_00_in25 = reg_0535;
    41: op1_00_in25 = reg_0261;
    42: op1_00_in25 = reg_0139;
    44: op1_00_in25 = reg_0087;
    95: op1_00_in25 = reg_0087;
    45: op1_00_in25 = reg_0377;
    46: op1_00_in25 = reg_0495;
    47: op1_00_in25 = imem01_in[31:28];
    48: op1_00_in25 = reg_0621;
    49: op1_00_in25 = imem06_in[111:108];
    50: op1_00_in25 = reg_0241;
    51: op1_00_in25 = reg_0333;
    52: op1_00_in25 = reg_0038;
    53: op1_00_in25 = reg_0820;
    54: op1_00_in25 = reg_0288;
    55: op1_00_in25 = reg_0578;
    56: op1_00_in25 = reg_0780;
    59: op1_00_in25 = reg_0895;
    60: op1_00_in25 = imem01_in[115:112];
    62: op1_00_in25 = reg_0902;
    63: op1_00_in25 = imem04_in[95:92];
    64: op1_00_in25 = reg_0151;
    65: op1_00_in25 = reg_0613;
    66: op1_00_in25 = reg_0624;
    67: op1_00_in25 = reg_0632;
    68: op1_00_in25 = imem07_in[67:64];
    69: op1_00_in25 = reg_0814;
    70: op1_00_in25 = reg_0658;
    72: op1_00_in25 = imem04_in[15:12];
    73: op1_00_in25 = reg_1010;
    74: op1_00_in25 = reg_0720;
    76: op1_00_in25 = reg_0592;
    77: op1_00_in25 = reg_1032;
    78: op1_00_in25 = imem04_in[107:104];
    79: op1_00_in25 = reg_0022;
    80: op1_00_in25 = reg_1011;
    83: op1_00_in25 = reg_0954;
    84: op1_00_in25 = reg_0823;
    85: op1_00_in25 = reg_0065;
    87: op1_00_in25 = reg_0729;
    88: op1_00_in25 = imem05_in[103:100];
    90: op1_00_in25 = imem05_in[115:112];
    91: op1_00_in25 = reg_1020;
    92: op1_00_in25 = reg_0426;
    93: op1_00_in25 = imem03_in[87:84];
    94: op1_00_in25 = reg_0645;
    96: op1_00_in25 = imem02_in[11:8];
    97: op1_00_in25 = imem01_in[55:52];
    default: op1_00_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv25 = 1;
    6: op1_00_inv25 = 1;
    8: op1_00_inv25 = 1;
    16: op1_00_inv25 = 1;
    17: op1_00_inv25 = 1;
    19: op1_00_inv25 = 1;
    21: op1_00_inv25 = 1;
    22: op1_00_inv25 = 1;
    23: op1_00_inv25 = 1;
    24: op1_00_inv25 = 1;
    27: op1_00_inv25 = 1;
    29: op1_00_inv25 = 1;
    30: op1_00_inv25 = 1;
    35: op1_00_inv25 = 1;
    38: op1_00_inv25 = 1;
    39: op1_00_inv25 = 1;
    41: op1_00_inv25 = 1;
    46: op1_00_inv25 = 1;
    47: op1_00_inv25 = 1;
    48: op1_00_inv25 = 1;
    50: op1_00_inv25 = 1;
    51: op1_00_inv25 = 1;
    54: op1_00_inv25 = 1;
    55: op1_00_inv25 = 1;
    56: op1_00_inv25 = 1;
    59: op1_00_inv25 = 1;
    60: op1_00_inv25 = 1;
    62: op1_00_inv25 = 1;
    65: op1_00_inv25 = 1;
    66: op1_00_inv25 = 1;
    67: op1_00_inv25 = 1;
    68: op1_00_inv25 = 1;
    70: op1_00_inv25 = 1;
    74: op1_00_inv25 = 1;
    76: op1_00_inv25 = 1;
    78: op1_00_inv25 = 1;
    79: op1_00_inv25 = 1;
    80: op1_00_inv25 = 1;
    83: op1_00_inv25 = 1;
    85: op1_00_inv25 = 1;
    87: op1_00_inv25 = 1;
    88: op1_00_inv25 = 1;
    90: op1_00_inv25 = 1;
    91: op1_00_inv25 = 1;
    92: op1_00_inv25 = 1;
    95: op1_00_inv25 = 1;
    96: op1_00_inv25 = 1;
    97: op1_00_inv25 = 1;
    default: op1_00_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in26 = imem01_in[47:44];
    6: op1_00_in26 = imem06_in[15:12];
    7: op1_00_in26 = imem02_in[75:72];
    8: op1_00_in26 = reg_0955;
    10: op1_00_in26 = reg_0639;
    11: op1_00_in26 = reg_0659;
    12: op1_00_in26 = reg_0421;
    13: op1_00_in26 = reg_0230;
    14: op1_00_in26 = reg_0626;
    15: op1_00_in26 = reg_0242;
    16: op1_00_in26 = reg_0904;
    17: op1_00_in26 = reg_0298;
    18: op1_00_in26 = imem07_in[71:68];
    19: op1_00_in26 = reg_0406;
    92: op1_00_in26 = reg_0406;
    20: op1_00_in26 = imem07_in[111:108];
    68: op1_00_in26 = imem07_in[111:108];
    21: op1_00_in26 = reg_0560;
    22: op1_00_in26 = reg_0424;
    23: op1_00_in26 = reg_1037;
    24: op1_00_in26 = imem06_in[95:92];
    25: op1_00_in26 = reg_0089;
    26: op1_00_in26 = reg_0541;
    27: op1_00_in26 = reg_0247;
    28: op1_00_in26 = reg_0777;
    29: op1_00_in26 = reg_0175;
    30: op1_00_in26 = reg_0299;
    31: op1_00_in26 = reg_0748;
    33: op1_00_in26 = reg_0248;
    34: op1_00_in26 = reg_1040;
    35: op1_00_in26 = reg_0446;
    36: op1_00_in26 = reg_0428;
    38: op1_00_in26 = reg_0124;
    39: op1_00_in26 = imem01_in[51:48];
    40: op1_00_in26 = reg_0357;
    41: op1_00_in26 = reg_0872;
    42: op1_00_in26 = imem06_in[3:0];
    44: op1_00_in26 = reg_0769;
    45: op1_00_in26 = reg_0807;
    46: op1_00_in26 = reg_0385;
    47: op1_00_in26 = imem01_in[87:84];
    48: op1_00_in26 = reg_0334;
    49: op1_00_in26 = reg_0614;
    50: op1_00_in26 = reg_0609;
    51: op1_00_in26 = reg_0438;
    52: op1_00_in26 = reg_0311;
    53: op1_00_in26 = reg_0518;
    54: op1_00_in26 = reg_0059;
    55: op1_00_in26 = reg_0764;
    56: op1_00_in26 = reg_0241;
    59: op1_00_in26 = reg_0611;
    60: op1_00_in26 = reg_0786;
    62: op1_00_in26 = reg_0610;
    63: op1_00_in26 = reg_0536;
    64: op1_00_in26 = reg_0156;
    65: op1_00_in26 = reg_0533;
    66: op1_00_in26 = reg_0630;
    67: op1_00_in26 = reg_0011;
    69: op1_00_in26 = reg_0091;
    70: op1_00_in26 = reg_0065;
    72: op1_00_in26 = imem04_in[55:52];
    73: op1_00_in26 = imem07_in[3:0];
    74: op1_00_in26 = reg_0723;
    76: op1_00_in26 = reg_0501;
    77: op1_00_in26 = reg_0592;
    78: op1_00_in26 = reg_1004;
    79: op1_00_in26 = reg_0573;
    80: op1_00_in26 = reg_0754;
    83: op1_00_in26 = reg_0647;
    84: op1_00_in26 = reg_0596;
    85: op1_00_in26 = reg_0495;
    87: op1_00_in26 = reg_0510;
    88: op1_00_in26 = imem05_in[127:124];
    90: op1_00_in26 = reg_0866;
    91: op1_00_in26 = reg_0370;
    93: op1_00_in26 = reg_0785;
    94: op1_00_in26 = reg_0359;
    95: op1_00_in26 = reg_0335;
    96: op1_00_in26 = imem02_in[27:24];
    97: op1_00_in26 = imem01_in[71:68];
    default: op1_00_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_00_inv26 = 1;
    10: op1_00_inv26 = 1;
    12: op1_00_inv26 = 1;
    13: op1_00_inv26 = 1;
    14: op1_00_inv26 = 1;
    15: op1_00_inv26 = 1;
    17: op1_00_inv26 = 1;
    18: op1_00_inv26 = 1;
    19: op1_00_inv26 = 1;
    21: op1_00_inv26 = 1;
    26: op1_00_inv26 = 1;
    28: op1_00_inv26 = 1;
    29: op1_00_inv26 = 1;
    31: op1_00_inv26 = 1;
    33: op1_00_inv26 = 1;
    34: op1_00_inv26 = 1;
    36: op1_00_inv26 = 1;
    40: op1_00_inv26 = 1;
    49: op1_00_inv26 = 1;
    53: op1_00_inv26 = 1;
    54: op1_00_inv26 = 1;
    56: op1_00_inv26 = 1;
    60: op1_00_inv26 = 1;
    62: op1_00_inv26 = 1;
    63: op1_00_inv26 = 1;
    66: op1_00_inv26 = 1;
    67: op1_00_inv26 = 1;
    68: op1_00_inv26 = 1;
    72: op1_00_inv26 = 1;
    73: op1_00_inv26 = 1;
    76: op1_00_inv26 = 1;
    79: op1_00_inv26 = 1;
    80: op1_00_inv26 = 1;
    83: op1_00_inv26 = 1;
    87: op1_00_inv26 = 1;
    88: op1_00_inv26 = 1;
    91: op1_00_inv26 = 1;
    94: op1_00_inv26 = 1;
    96: op1_00_inv26 = 1;
    default: op1_00_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in27 = imem01_in[59:56];
    6: op1_00_in27 = imem06_in[71:68];
    7: op1_00_in27 = reg_0658;
    8: op1_00_in27 = reg_0967;
    10: op1_00_in27 = reg_0640;
    11: op1_00_in27 = reg_0667;
    12: op1_00_in27 = reg_0434;
    36: op1_00_in27 = reg_0434;
    13: op1_00_in27 = reg_0500;
    14: op1_00_in27 = reg_0618;
    15: op1_00_in27 = reg_0503;
    16: op1_00_in27 = reg_0103;
    38: op1_00_in27 = reg_0103;
    17: op1_00_in27 = reg_0288;
    18: op1_00_in27 = reg_0724;
    19: op1_00_in27 = reg_0401;
    20: op1_00_in27 = imem07_in[119:116];
    21: op1_00_in27 = reg_0546;
    22: op1_00_in27 = reg_0430;
    23: op1_00_in27 = reg_1040;
    24: op1_00_in27 = imem06_in[103:100];
    25: op1_00_in27 = reg_0776;
    26: op1_00_in27 = reg_0062;
    27: op1_00_in27 = reg_0238;
    28: op1_00_in27 = reg_0044;
    29: op1_00_in27 = reg_0162;
    30: op1_00_in27 = reg_0544;
    33: op1_00_in27 = reg_0544;
    31: op1_00_in27 = reg_0054;
    34: op1_00_in27 = reg_0105;
    35: op1_00_in27 = reg_0440;
    39: op1_00_in27 = imem01_in[95:92];
    40: op1_00_in27 = reg_0343;
    41: op1_00_in27 = imem03_in[3:0];
    42: op1_00_in27 = imem06_in[23:20];
    44: op1_00_in27 = reg_0869;
    45: op1_00_in27 = reg_0376;
    52: op1_00_in27 = reg_0376;
    46: op1_00_in27 = reg_0395;
    47: op1_00_in27 = reg_0786;
    48: op1_00_in27 = reg_0842;
    49: op1_00_in27 = reg_0624;
    80: op1_00_in27 = reg_0624;
    50: op1_00_in27 = reg_0626;
    51: op1_00_in27 = reg_0146;
    53: op1_00_in27 = reg_0513;
    54: op1_00_in27 = reg_0281;
    84: op1_00_in27 = reg_0281;
    55: op1_00_in27 = imem05_in[83:80];
    56: op1_00_in27 = reg_0617;
    59: op1_00_in27 = reg_0781;
    60: op1_00_in27 = reg_0762;
    62: op1_00_in27 = reg_0906;
    63: op1_00_in27 = reg_0282;
    64: op1_00_in27 = reg_0154;
    65: op1_00_in27 = reg_0439;
    87: op1_00_in27 = reg_0439;
    66: op1_00_in27 = reg_0408;
    67: op1_00_in27 = reg_0619;
    68: op1_00_in27 = reg_0728;
    69: op1_00_in27 = reg_0840;
    70: op1_00_in27 = reg_0494;
    72: op1_00_in27 = imem04_in[67:64];
    73: op1_00_in27 = imem07_in[11:8];
    74: op1_00_in27 = reg_0717;
    76: op1_00_in27 = reg_0798;
    77: op1_00_in27 = reg_0234;
    78: op1_00_in27 = reg_0483;
    79: op1_00_in27 = reg_0566;
    83: op1_00_in27 = reg_0143;
    85: op1_00_in27 = imem05_in[47:44];
    88: op1_00_in27 = reg_0944;
    90: op1_00_in27 = reg_0492;
    91: op1_00_in27 = reg_0914;
    92: op1_00_in27 = reg_0868;
    93: op1_00_in27 = reg_0357;
    94: op1_00_in27 = reg_0389;
    95: op1_00_in27 = reg_0516;
    96: op1_00_in27 = imem02_in[63:60];
    97: op1_00_in27 = imem01_in[87:84];
    default: op1_00_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv27 = 1;
    10: op1_00_inv27 = 1;
    11: op1_00_inv27 = 1;
    13: op1_00_inv27 = 1;
    14: op1_00_inv27 = 1;
    17: op1_00_inv27 = 1;
    19: op1_00_inv27 = 1;
    20: op1_00_inv27 = 1;
    21: op1_00_inv27 = 1;
    22: op1_00_inv27 = 1;
    23: op1_00_inv27 = 1;
    24: op1_00_inv27 = 1;
    26: op1_00_inv27 = 1;
    27: op1_00_inv27 = 1;
    29: op1_00_inv27 = 1;
    31: op1_00_inv27 = 1;
    33: op1_00_inv27 = 1;
    42: op1_00_inv27 = 1;
    45: op1_00_inv27 = 1;
    46: op1_00_inv27 = 1;
    48: op1_00_inv27 = 1;
    49: op1_00_inv27 = 1;
    50: op1_00_inv27 = 1;
    52: op1_00_inv27 = 1;
    56: op1_00_inv27 = 1;
    59: op1_00_inv27 = 1;
    60: op1_00_inv27 = 1;
    62: op1_00_inv27 = 1;
    63: op1_00_inv27 = 1;
    66: op1_00_inv27 = 1;
    68: op1_00_inv27 = 1;
    69: op1_00_inv27 = 1;
    74: op1_00_inv27 = 1;
    76: op1_00_inv27 = 1;
    77: op1_00_inv27 = 1;
    78: op1_00_inv27 = 1;
    80: op1_00_inv27 = 1;
    83: op1_00_inv27 = 1;
    84: op1_00_inv27 = 1;
    85: op1_00_inv27 = 1;
    88: op1_00_inv27 = 1;
    90: op1_00_inv27 = 1;
    91: op1_00_inv27 = 1;
    93: op1_00_inv27 = 1;
    95: op1_00_inv27 = 1;
    97: op1_00_inv27 = 1;
    default: op1_00_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in28 = imem01_in[83:80];
    6: op1_00_in28 = imem06_in[75:72];
    7: op1_00_in28 = reg_0654;
    8: op1_00_in28 = reg_0964;
    10: op1_00_in28 = reg_0648;
    11: op1_00_in28 = reg_0341;
    12: op1_00_in28 = reg_0166;
    13: op1_00_in28 = reg_0913;
    14: op1_00_in28 = reg_0348;
    15: op1_00_in28 = reg_0236;
    16: op1_00_in28 = reg_0111;
    17: op1_00_in28 = reg_0061;
    18: op1_00_in28 = reg_0729;
    19: op1_00_in28 = reg_1029;
    20: op1_00_in28 = reg_0716;
    21: op1_00_in28 = reg_0065;
    22: op1_00_in28 = reg_0436;
    23: op1_00_in28 = reg_0122;
    24: op1_00_in28 = imem06_in[119:116];
    25: op1_00_in28 = reg_0792;
    26: op1_00_in28 = reg_0276;
    27: op1_00_in28 = reg_0230;
    28: op1_00_in28 = imem05_in[87:84];
    29: op1_00_in28 = reg_0163;
    30: op1_00_in28 = reg_0219;
    33: op1_00_in28 = reg_0219;
    31: op1_00_in28 = reg_0751;
    34: op1_00_in28 = reg_0118;
    38: op1_00_in28 = reg_0118;
    35: op1_00_in28 = reg_0443;
    36: op1_00_in28 = reg_0444;
    39: op1_00_in28 = reg_0235;
    40: op1_00_in28 = reg_0938;
    41: op1_00_in28 = imem03_in[11:8];
    69: op1_00_in28 = imem03_in[11:8];
    42: op1_00_in28 = imem06_in[71:68];
    44: op1_00_in28 = reg_0829;
    45: op1_00_in28 = reg_0518;
    46: op1_00_in28 = reg_0391;
    47: op1_00_in28 = reg_0003;
    48: op1_00_in28 = reg_0093;
    49: op1_00_in28 = reg_0892;
    50: op1_00_in28 = reg_0633;
    51: op1_00_in28 = reg_0139;
    83: op1_00_in28 = reg_0139;
    52: op1_00_in28 = reg_0234;
    53: op1_00_in28 = reg_0993;
    54: op1_00_in28 = reg_0554;
    55: op1_00_in28 = imem05_in[107:104];
    56: op1_00_in28 = reg_0605;
    59: op1_00_in28 = reg_0699;
    60: op1_00_in28 = reg_0933;
    62: op1_00_in28 = reg_0615;
    63: op1_00_in28 = reg_1005;
    64: op1_00_in28 = reg_0153;
    65: op1_00_in28 = reg_0863;
    66: op1_00_in28 = reg_0405;
    67: op1_00_in28 = reg_0293;
    68: op1_00_in28 = reg_0719;
    70: op1_00_in28 = reg_0495;
    72: op1_00_in28 = imem04_in[123:120];
    73: op1_00_in28 = imem07_in[31:28];
    74: op1_00_in28 = reg_0725;
    76: op1_00_in28 = reg_1043;
    77: op1_00_in28 = reg_1024;
    78: op1_00_in28 = reg_0511;
    79: op1_00_in28 = imem07_in[11:8];
    80: op1_00_in28 = reg_0698;
    87: op1_00_in28 = reg_0698;
    84: op1_00_in28 = reg_0609;
    85: op1_00_in28 = reg_1021;
    88: op1_00_in28 = reg_0128;
    90: op1_00_in28 = reg_0142;
    91: op1_00_in28 = reg_0177;
    92: op1_00_in28 = reg_0181;
    93: op1_00_in28 = reg_0743;
    94: op1_00_in28 = reg_0608;
    95: op1_00_in28 = reg_0155;
    96: op1_00_in28 = imem02_in[87:84];
    97: op1_00_in28 = imem01_in[115:112];
    default: op1_00_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv28 = 1;
    7: op1_00_inv28 = 1;
    8: op1_00_inv28 = 1;
    11: op1_00_inv28 = 1;
    13: op1_00_inv28 = 1;
    17: op1_00_inv28 = 1;
    18: op1_00_inv28 = 1;
    21: op1_00_inv28 = 1;
    23: op1_00_inv28 = 1;
    24: op1_00_inv28 = 1;
    27: op1_00_inv28 = 1;
    29: op1_00_inv28 = 1;
    35: op1_00_inv28 = 1;
    40: op1_00_inv28 = 1;
    44: op1_00_inv28 = 1;
    45: op1_00_inv28 = 1;
    47: op1_00_inv28 = 1;
    48: op1_00_inv28 = 1;
    50: op1_00_inv28 = 1;
    55: op1_00_inv28 = 1;
    56: op1_00_inv28 = 1;
    59: op1_00_inv28 = 1;
    62: op1_00_inv28 = 1;
    64: op1_00_inv28 = 1;
    65: op1_00_inv28 = 1;
    66: op1_00_inv28 = 1;
    68: op1_00_inv28 = 1;
    69: op1_00_inv28 = 1;
    70: op1_00_inv28 = 1;
    72: op1_00_inv28 = 1;
    76: op1_00_inv28 = 1;
    77: op1_00_inv28 = 1;
    78: op1_00_inv28 = 1;
    83: op1_00_inv28 = 1;
    85: op1_00_inv28 = 1;
    88: op1_00_inv28 = 1;
    90: op1_00_inv28 = 1;
    92: op1_00_inv28 = 1;
    94: op1_00_inv28 = 1;
    95: op1_00_inv28 = 1;
    96: op1_00_inv28 = 1;
    default: op1_00_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in29 = imem01_in[91:88];
    6: op1_00_in29 = imem06_in[79:76];
    7: op1_00_in29 = reg_0660;
    8: op1_00_in29 = reg_0968;
    10: op1_00_in29 = reg_0364;
    11: op1_00_in29 = reg_0318;
    12: op1_00_in29 = reg_0168;
    13: op1_00_in29 = reg_1034;
    14: op1_00_in29 = reg_0381;
    15: op1_00_in29 = reg_0487;
    16: op1_00_in29 = reg_0116;
    34: op1_00_in29 = reg_0116;
    17: op1_00_in29 = reg_0078;
    18: op1_00_in29 = reg_0705;
    19: op1_00_in29 = reg_0752;
    20: op1_00_in29 = reg_0731;
    21: op1_00_in29 = reg_0076;
    22: op1_00_in29 = reg_0422;
    23: op1_00_in29 = reg_0124;
    47: op1_00_in29 = reg_0124;
    24: op1_00_in29 = reg_0628;
    25: op1_00_in29 = reg_0086;
    26: op1_00_in29 = reg_0732;
    27: op1_00_in29 = reg_1036;
    28: op1_00_in29 = imem05_in[91:88];
    29: op1_00_in29 = reg_0166;
    30: op1_00_in29 = reg_1042;
    33: op1_00_in29 = reg_1042;
    31: op1_00_in29 = reg_0044;
    35: op1_00_in29 = reg_0183;
    36: op1_00_in29 = reg_0448;
    38: op1_00_in29 = reg_0100;
    39: op1_00_in29 = reg_0223;
    40: op1_00_in29 = reg_0245;
    41: op1_00_in29 = imem03_in[39:36];
    42: op1_00_in29 = imem06_in[99:96];
    44: op1_00_in29 = reg_0740;
    45: op1_00_in29 = reg_0987;
    84: op1_00_in29 = reg_0987;
    46: op1_00_in29 = reg_0386;
    66: op1_00_in29 = reg_0386;
    48: op1_00_in29 = reg_0776;
    49: op1_00_in29 = reg_0781;
    50: op1_00_in29 = imem07_in[23:20];
    79: op1_00_in29 = imem07_in[23:20];
    51: op1_00_in29 = imem06_in[15:12];
    52: op1_00_in29 = reg_1000;
    53: op1_00_in29 = reg_0980;
    54: op1_00_in29 = reg_0027;
    55: op1_00_in29 = reg_0962;
    56: op1_00_in29 = reg_0029;
    59: op1_00_in29 = reg_0605;
    60: op1_00_in29 = reg_0919;
    62: op1_00_in29 = reg_0232;
    63: op1_00_in29 = reg_0292;
    64: op1_00_in29 = reg_0137;
    83: op1_00_in29 = reg_0137;
    65: op1_00_in29 = reg_0699;
    67: op1_00_in29 = reg_0257;
    68: op1_00_in29 = reg_0711;
    69: op1_00_in29 = imem03_in[27:24];
    70: op1_00_in29 = reg_0251;
    72: op1_00_in29 = reg_0301;
    73: op1_00_in29 = imem07_in[51:48];
    74: op1_00_in29 = reg_0729;
    76: op1_00_in29 = reg_0304;
    77: op1_00_in29 = reg_0793;
    78: op1_00_in29 = reg_0912;
    80: op1_00_in29 = reg_0619;
    85: op1_00_in29 = reg_0866;
    87: op1_00_in29 = reg_0264;
    88: op1_00_in29 = reg_0235;
    90: op1_00_in29 = reg_0583;
    91: op1_00_in29 = reg_0611;
    92: op1_00_in29 = reg_0447;
    93: op1_00_in29 = reg_0307;
    94: op1_00_in29 = reg_0734;
    95: op1_00_in29 = reg_0885;
    96: op1_00_in29 = imem02_in[115:112];
    97: op1_00_in29 = imem01_in[119:116];
    default: op1_00_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv29 = 1;
    7: op1_00_inv29 = 1;
    10: op1_00_inv29 = 1;
    12: op1_00_inv29 = 1;
    13: op1_00_inv29 = 1;
    14: op1_00_inv29 = 1;
    17: op1_00_inv29 = 1;
    18: op1_00_inv29 = 1;
    20: op1_00_inv29 = 1;
    23: op1_00_inv29 = 1;
    27: op1_00_inv29 = 1;
    28: op1_00_inv29 = 1;
    29: op1_00_inv29 = 1;
    34: op1_00_inv29 = 1;
    36: op1_00_inv29 = 1;
    38: op1_00_inv29 = 1;
    39: op1_00_inv29 = 1;
    40: op1_00_inv29 = 1;
    41: op1_00_inv29 = 1;
    42: op1_00_inv29 = 1;
    44: op1_00_inv29 = 1;
    45: op1_00_inv29 = 1;
    46: op1_00_inv29 = 1;
    47: op1_00_inv29 = 1;
    48: op1_00_inv29 = 1;
    49: op1_00_inv29 = 1;
    51: op1_00_inv29 = 1;
    53: op1_00_inv29 = 1;
    54: op1_00_inv29 = 1;
    55: op1_00_inv29 = 1;
    56: op1_00_inv29 = 1;
    60: op1_00_inv29 = 1;
    63: op1_00_inv29 = 1;
    65: op1_00_inv29 = 1;
    66: op1_00_inv29 = 1;
    69: op1_00_inv29 = 1;
    72: op1_00_inv29 = 1;
    74: op1_00_inv29 = 1;
    79: op1_00_inv29 = 1;
    83: op1_00_inv29 = 1;
    87: op1_00_inv29 = 1;
    88: op1_00_inv29 = 1;
    90: op1_00_inv29 = 1;
    91: op1_00_inv29 = 1;
    92: op1_00_inv29 = 1;
    93: op1_00_inv29 = 1;
    96: op1_00_inv29 = 1;
    default: op1_00_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_00_in30 = reg_0513;
    6: op1_00_in30 = imem06_in[87:84];
    7: op1_00_in30 = reg_0661;
    8: op1_00_in30 = reg_0953;
    10: op1_00_in30 = reg_0359;
    11: op1_00_in30 = reg_0338;
    13: op1_00_in30 = reg_0111;
    14: op1_00_in30 = reg_0367;
    15: op1_00_in30 = reg_0507;
    16: op1_00_in30 = reg_0117;
    17: op1_00_in30 = reg_0066;
    18: op1_00_in30 = reg_0727;
    19: op1_00_in30 = reg_0801;
    20: op1_00_in30 = reg_0708;
    21: op1_00_in30 = reg_0755;
    22: op1_00_in30 = reg_0433;
    23: op1_00_in30 = reg_0103;
    24: op1_00_in30 = reg_0607;
    25: op1_00_in30 = reg_0084;
    26: op1_00_in30 = reg_0285;
    27: op1_00_in30 = reg_0105;
    28: op1_00_in30 = imem05_in[95:92];
    29: op1_00_in30 = reg_0164;
    35: op1_00_in30 = reg_0164;
    30: op1_00_in30 = reg_0871;
    31: op1_00_in30 = imem05_in[99:96];
    33: op1_00_in30 = reg_0230;
    34: op1_00_in30 = reg_0120;
    36: op1_00_in30 = reg_0162;
    38: op1_00_in30 = imem02_in[7:4];
    39: op1_00_in30 = reg_0563;
    40: op1_00_in30 = reg_0581;
    41: op1_00_in30 = imem03_in[43:40];
    42: op1_00_in30 = reg_0614;
    44: op1_00_in30 = reg_0124;
    45: op1_00_in30 = reg_0998;
    46: op1_00_in30 = reg_0388;
    47: op1_00_in30 = reg_0116;
    48: op1_00_in30 = reg_0086;
    49: op1_00_in30 = reg_0403;
    50: op1_00_in30 = imem07_in[39:36];
    51: op1_00_in30 = imem06_in[103:100];
    52: op1_00_in30 = reg_0997;
    53: op1_00_in30 = reg_0978;
    54: op1_00_in30 = reg_0043;
    55: op1_00_in30 = reg_0963;
    56: op1_00_in30 = reg_0005;
    59: op1_00_in30 = reg_0017;
    60: op1_00_in30 = reg_0503;
    62: op1_00_in30 = reg_0832;
    63: op1_00_in30 = reg_0568;
    64: op1_00_in30 = imem06_in[7:4];
    65: op1_00_in30 = reg_0619;
    66: op1_00_in30 = reg_0264;
    67: op1_00_in30 = reg_0630;
    68: op1_00_in30 = reg_0002;
    69: op1_00_in30 = imem03_in[63:60];
    70: op1_00_in30 = reg_0856;
    72: op1_00_in30 = reg_1009;
    73: op1_00_in30 = imem07_in[63:60];
    74: op1_00_in30 = reg_0744;
    76: op1_00_in30 = reg_0906;
    77: op1_00_in30 = reg_0831;
    78: op1_00_in30 = reg_0888;
    79: op1_00_in30 = imem07_in[47:44];
    80: op1_00_in30 = reg_0857;
    83: op1_00_in30 = reg_0365;
    84: op1_00_in30 = reg_0984;
    85: op1_00_in30 = reg_0954;
    87: op1_00_in30 = reg_0029;
    88: op1_00_in30 = reg_0648;
    90: op1_00_in30 = reg_0178;
    91: op1_00_in30 = reg_0782;
    92: op1_00_in30 = reg_0183;
    93: op1_00_in30 = reg_0007;
    94: op1_00_in30 = reg_0776;
    95: op1_00_in30 = reg_0218;
    96: op1_00_in30 = imem02_in[119:116];
    97: op1_00_in30 = imem01_in[123:120];
    default: op1_00_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv30 = 1;
    6: op1_00_inv30 = 1;
    8: op1_00_inv30 = 1;
    11: op1_00_inv30 = 1;
    19: op1_00_inv30 = 1;
    20: op1_00_inv30 = 1;
    28: op1_00_inv30 = 1;
    34: op1_00_inv30 = 1;
    36: op1_00_inv30 = 1;
    40: op1_00_inv30 = 1;
    41: op1_00_inv30 = 1;
    42: op1_00_inv30 = 1;
    44: op1_00_inv30 = 1;
    45: op1_00_inv30 = 1;
    47: op1_00_inv30 = 1;
    49: op1_00_inv30 = 1;
    50: op1_00_inv30 = 1;
    51: op1_00_inv30 = 1;
    53: op1_00_inv30 = 1;
    55: op1_00_inv30 = 1;
    62: op1_00_inv30 = 1;
    63: op1_00_inv30 = 1;
    67: op1_00_inv30 = 1;
    68: op1_00_inv30 = 1;
    70: op1_00_inv30 = 1;
    74: op1_00_inv30 = 1;
    76: op1_00_inv30 = 1;
    77: op1_00_inv30 = 1;
    79: op1_00_inv30 = 1;
    87: op1_00_inv30 = 1;
    90: op1_00_inv30 = 1;
    94: op1_00_inv30 = 1;
    default: op1_00_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_00_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_00_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in00 = reg_0514;
    6: op1_01_in00 = imem06_in[127:124];
    7: op1_01_in00 = reg_0640;
    8: op1_01_in00 = reg_0960;
    4: op1_01_in00 = imem07_in[47:44];
    9: op1_01_in00 = imem00_in[19:16];
    75: op1_01_in00 = imem00_in[19:16];
    3: op1_01_in00 = imem07_in[103:100];
    73: op1_01_in00 = imem07_in[103:100];
    10: op1_01_in00 = reg_0324;
    11: op1_01_in00 = reg_0335;
    12: op1_01_in00 = imem00_in[43:40];
    13: op1_01_in00 = reg_0099;
    2: op1_01_in00 = imem07_in[15:12];
    14: op1_01_in00 = reg_0380;
    15: op1_01_in00 = reg_0508;
    16: op1_01_in00 = imem02_in[31:28];
    17: op1_01_in00 = reg_0070;
    18: op1_01_in00 = imem00_in[3:0];
    20: op1_01_in00 = imem00_in[3:0];
    58: op1_01_in00 = imem00_in[3:0];
    71: op1_01_in00 = imem00_in[3:0];
    19: op1_01_in00 = reg_0011;
    21: op1_01_in00 = reg_0071;
    22: op1_01_in00 = imem00_in[51:48];
    29: op1_01_in00 = imem00_in[51:48];
    86: op1_01_in00 = imem00_in[51:48];
    23: op1_01_in00 = reg_0104;
    24: op1_01_in00 = reg_0616;
    25: op1_01_in00 = imem03_in[3:0];
    26: op1_01_in00 = reg_0286;
    27: op1_01_in00 = reg_0122;
    28: op1_01_in00 = imem05_in[123:120];
    31: op1_01_in00 = imem05_in[123:120];
    30: op1_01_in00 = reg_0228;
    32: op1_01_in00 = imem00_in[27:24];
    33: op1_01_in00 = reg_0885;
    34: op1_01_in00 = reg_0108;
    35: op1_01_in00 = imem00_in[55:52];
    89: op1_01_in00 = imem00_in[55:52];
    36: op1_01_in00 = reg_0182;
    37: op1_01_in00 = imem00_in[39:36];
    38: op1_01_in00 = imem02_in[19:16];
    39: op1_01_in00 = reg_0274;
    40: op1_01_in00 = reg_0370;
    80: op1_01_in00 = reg_0370;
    41: op1_01_in00 = reg_1050;
    42: op1_01_in00 = reg_0782;
    49: op1_01_in00 = reg_0782;
    43: op1_01_in00 = imem00_in[59:56];
    44: op1_01_in00 = reg_0118;
    45: op1_01_in00 = reg_0982;
    46: op1_01_in00 = reg_0222;
    47: op1_01_in00 = reg_0114;
    48: op1_01_in00 = reg_0506;
    50: op1_01_in00 = imem07_in[63:60];
    51: op1_01_in00 = reg_0073;
    52: op1_01_in00 = reg_0994;
    53: op1_01_in00 = reg_0988;
    54: op1_01_in00 = reg_0429;
    55: op1_01_in00 = reg_0958;
    56: op1_01_in00 = imem07_in[11:8];
    57: op1_01_in00 = imem00_in[15:12];
    82: op1_01_in00 = imem00_in[15:12];
    59: op1_01_in00 = reg_1010;
    60: op1_01_in00 = reg_0249;
    61: op1_01_in00 = imem00_in[7:4];
    62: op1_01_in00 = reg_0111;
    63: op1_01_in00 = reg_0524;
    64: op1_01_in00 = imem06_in[43:40];
    65: op1_01_in00 = reg_0348;
    66: op1_01_in00 = imem07_in[83:80];
    67: op1_01_in00 = reg_0241;
    68: op1_01_in00 = reg_0321;
    69: op1_01_in00 = imem03_in[87:84];
    70: op1_01_in00 = imem05_in[51:48];
    72: op1_01_in00 = reg_1016;
    74: op1_01_in00 = reg_0315;
    76: op1_01_in00 = reg_0512;
    77: op1_01_in00 = reg_0225;
    78: op1_01_in00 = reg_0931;
    79: op1_01_in00 = imem07_in[55:52];
    81: op1_01_in00 = imem00_in[31:28];
    83: op1_01_in00 = reg_0525;
    84: op1_01_in00 = reg_1001;
    85: op1_01_in00 = reg_0655;
    87: op1_01_in00 = reg_0783;
    88: op1_01_in00 = reg_0057;
    90: op1_01_in00 = reg_0436;
    91: op1_01_in00 = reg_0804;
    92: op1_01_in00 = reg_0690;
    93: op1_01_in00 = reg_0033;
    94: op1_01_in00 = reg_0408;
    95: op1_01_in00 = reg_0730;
    96: op1_01_in00 = reg_0069;
    97: op1_01_in00 = reg_0786;
    default: op1_01_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv00 = 1;
    6: op1_01_inv00 = 1;
    7: op1_01_inv00 = 1;
    18: op1_01_inv00 = 1;
    21: op1_01_inv00 = 1;
    22: op1_01_inv00 = 1;
    23: op1_01_inv00 = 1;
    25: op1_01_inv00 = 1;
    26: op1_01_inv00 = 1;
    28: op1_01_inv00 = 1;
    30: op1_01_inv00 = 1;
    31: op1_01_inv00 = 1;
    33: op1_01_inv00 = 1;
    34: op1_01_inv00 = 1;
    35: op1_01_inv00 = 1;
    36: op1_01_inv00 = 1;
    38: op1_01_inv00 = 1;
    41: op1_01_inv00 = 1;
    43: op1_01_inv00 = 1;
    44: op1_01_inv00 = 1;
    46: op1_01_inv00 = 1;
    49: op1_01_inv00 = 1;
    51: op1_01_inv00 = 1;
    52: op1_01_inv00 = 1;
    54: op1_01_inv00 = 1;
    56: op1_01_inv00 = 1;
    58: op1_01_inv00 = 1;
    59: op1_01_inv00 = 1;
    60: op1_01_inv00 = 1;
    62: op1_01_inv00 = 1;
    64: op1_01_inv00 = 1;
    68: op1_01_inv00 = 1;
    69: op1_01_inv00 = 1;
    70: op1_01_inv00 = 1;
    71: op1_01_inv00 = 1;
    72: op1_01_inv00 = 1;
    74: op1_01_inv00 = 1;
    75: op1_01_inv00 = 1;
    80: op1_01_inv00 = 1;
    83: op1_01_inv00 = 1;
    87: op1_01_inv00 = 1;
    88: op1_01_inv00 = 1;
    89: op1_01_inv00 = 1;
    90: op1_01_inv00 = 1;
    default: op1_01_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in01 = reg_0502;
    6: op1_01_in01 = reg_0625;
    46: op1_01_in01 = reg_0625;
    7: op1_01_in01 = reg_0649;
    8: op1_01_in01 = reg_0260;
    4: op1_01_in01 = imem07_in[51:48];
    9: op1_01_in01 = imem00_in[59:56];
    37: op1_01_in01 = imem00_in[59:56];
    89: op1_01_in01 = imem00_in[59:56];
    3: op1_01_in01 = imem07_in[115:112];
    10: op1_01_in01 = reg_0353;
    11: op1_01_in01 = reg_0328;
    12: op1_01_in01 = imem00_in[99:96];
    13: op1_01_in01 = reg_0108;
    2: op1_01_in01 = imem07_in[27:24];
    14: op1_01_in01 = reg_0799;
    15: op1_01_in01 = reg_1032;
    16: op1_01_in01 = imem02_in[79:76];
    17: op1_01_in01 = imem05_in[27:24];
    18: op1_01_in01 = imem00_in[27:24];
    75: op1_01_in01 = imem00_in[27:24];
    19: op1_01_in01 = imem07_in[87:84];
    66: op1_01_in01 = imem07_in[87:84];
    20: op1_01_in01 = imem00_in[55:52];
    21: op1_01_in01 = reg_0732;
    22: op1_01_in01 = imem00_in[127:124];
    23: op1_01_in01 = imem02_in[23:20];
    24: op1_01_in01 = reg_0609;
    25: op1_01_in01 = imem03_in[55:52];
    26: op1_01_in01 = imem05_in[19:16];
    27: op1_01_in01 = reg_0124;
    28: op1_01_in01 = imem05_in[127:124];
    29: op1_01_in01 = imem00_in[83:80];
    43: op1_01_in01 = imem00_in[83:80];
    30: op1_01_in01 = reg_1018;
    31: op1_01_in01 = reg_0962;
    32: op1_01_in01 = imem00_in[39:36];
    58: op1_01_in01 = imem00_in[39:36];
    33: op1_01_in01 = reg_1043;
    34: op1_01_in01 = imem02_in[7:4];
    35: op1_01_in01 = imem00_in[79:76];
    86: op1_01_in01 = imem00_in[79:76];
    36: op1_01_in01 = reg_0160;
    38: op1_01_in01 = imem02_in[51:48];
    39: op1_01_in01 = reg_0238;
    40: op1_01_in01 = reg_0795;
    41: op1_01_in01 = reg_0317;
    42: op1_01_in01 = reg_0783;
    44: op1_01_in01 = reg_0114;
    45: op1_01_in01 = reg_0992;
    47: op1_01_in01 = reg_0106;
    48: op1_01_in01 = reg_0084;
    49: op1_01_in01 = reg_0577;
    50: op1_01_in01 = imem07_in[71:68];
    51: op1_01_in01 = reg_0895;
    52: op1_01_in01 = imem04_in[59:56];
    53: op1_01_in01 = reg_0990;
    54: op1_01_in01 = reg_0882;
    55: op1_01_in01 = reg_0971;
    56: op1_01_in01 = imem07_in[83:80];
    57: op1_01_in01 = imem00_in[51:48];
    59: op1_01_in01 = reg_0545;
    60: op1_01_in01 = reg_0522;
    77: op1_01_in01 = reg_0522;
    61: op1_01_in01 = imem00_in[11:8];
    62: op1_01_in01 = reg_1053;
    76: op1_01_in01 = reg_1053;
    63: op1_01_in01 = reg_0809;
    64: op1_01_in01 = imem06_in[91:88];
    65: op1_01_in01 = reg_0816;
    67: op1_01_in01 = reg_0405;
    68: op1_01_in01 = reg_0406;
    69: op1_01_in01 = reg_0012;
    70: op1_01_in01 = imem05_in[59:56];
    71: op1_01_in01 = imem00_in[15:12];
    72: op1_01_in01 = reg_0850;
    73: op1_01_in01 = imem07_in[123:120];
    74: op1_01_in01 = reg_0419;
    78: op1_01_in01 = reg_0752;
    79: op1_01_in01 = imem07_in[67:64];
    80: op1_01_in01 = reg_0834;
    81: op1_01_in01 = imem00_in[47:44];
    82: op1_01_in01 = imem00_in[23:20];
    83: op1_01_in01 = reg_0314;
    84: op1_01_in01 = reg_0978;
    85: op1_01_in01 = reg_0139;
    87: op1_01_in01 = reg_0719;
    88: op1_01_in01 = reg_0063;
    90: op1_01_in01 = reg_0145;
    91: op1_01_in01 = reg_0632;
    92: op1_01_in01 = reg_0157;
    93: op1_01_in01 = reg_0149;
    94: op1_01_in01 = reg_0365;
    95: op1_01_in01 = reg_0624;
    96: op1_01_in01 = reg_0255;
    97: op1_01_in01 = reg_0246;
    default: op1_01_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv01 = 1;
    7: op1_01_inv01 = 1;
    8: op1_01_inv01 = 1;
    10: op1_01_inv01 = 1;
    11: op1_01_inv01 = 1;
    12: op1_01_inv01 = 1;
    13: op1_01_inv01 = 1;
    2: op1_01_inv01 = 1;
    14: op1_01_inv01 = 1;
    15: op1_01_inv01 = 1;
    19: op1_01_inv01 = 1;
    24: op1_01_inv01 = 1;
    30: op1_01_inv01 = 1;
    32: op1_01_inv01 = 1;
    36: op1_01_inv01 = 1;
    37: op1_01_inv01 = 1;
    38: op1_01_inv01 = 1;
    39: op1_01_inv01 = 1;
    41: op1_01_inv01 = 1;
    42: op1_01_inv01 = 1;
    45: op1_01_inv01 = 1;
    46: op1_01_inv01 = 1;
    48: op1_01_inv01 = 1;
    50: op1_01_inv01 = 1;
    57: op1_01_inv01 = 1;
    58: op1_01_inv01 = 1;
    59: op1_01_inv01 = 1;
    60: op1_01_inv01 = 1;
    64: op1_01_inv01 = 1;
    69: op1_01_inv01 = 1;
    71: op1_01_inv01 = 1;
    74: op1_01_inv01 = 1;
    75: op1_01_inv01 = 1;
    76: op1_01_inv01 = 1;
    78: op1_01_inv01 = 1;
    79: op1_01_inv01 = 1;
    81: op1_01_inv01 = 1;
    82: op1_01_inv01 = 1;
    83: op1_01_inv01 = 1;
    84: op1_01_inv01 = 1;
    87: op1_01_inv01 = 1;
    89: op1_01_inv01 = 1;
    91: op1_01_inv01 = 1;
    93: op1_01_inv01 = 1;
    94: op1_01_inv01 = 1;
    95: op1_01_inv01 = 1;
    97: op1_01_inv01 = 1;
    default: op1_01_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in02 = reg_0503;
    6: op1_01_in02 = reg_0604;
    7: op1_01_in02 = reg_0652;
    8: op1_01_in02 = reg_0253;
    4: op1_01_in02 = imem07_in[75:72];
    50: op1_01_in02 = imem07_in[75:72];
    9: op1_01_in02 = imem00_in[75:72];
    3: op1_01_in02 = reg_0179;
    10: op1_01_in02 = reg_0310;
    11: op1_01_in02 = reg_0347;
    12: op1_01_in02 = reg_0682;
    22: op1_01_in02 = reg_0682;
    43: op1_01_in02 = reg_0682;
    13: op1_01_in02 = reg_0100;
    44: op1_01_in02 = reg_0100;
    2: op1_01_in02 = imem07_in[31:28];
    14: op1_01_in02 = reg_1030;
    15: op1_01_in02 = reg_1044;
    16: op1_01_in02 = imem02_in[87:84];
    17: op1_01_in02 = imem05_in[39:36];
    18: op1_01_in02 = imem00_in[31:28];
    75: op1_01_in02 = imem00_in[31:28];
    19: op1_01_in02 = reg_0716;
    20: op1_01_in02 = imem00_in[87:84];
    29: op1_01_in02 = imem00_in[87:84];
    21: op1_01_in02 = reg_0278;
    23: op1_01_in02 = imem02_in[35:32];
    24: op1_01_in02 = reg_0615;
    60: op1_01_in02 = reg_0615;
    25: op1_01_in02 = imem03_in[63:60];
    26: op1_01_in02 = imem05_in[31:28];
    27: op1_01_in02 = reg_0102;
    28: op1_01_in02 = reg_0971;
    30: op1_01_in02 = reg_0116;
    31: op1_01_in02 = reg_0959;
    55: op1_01_in02 = reg_0959;
    32: op1_01_in02 = imem00_in[103:100];
    86: op1_01_in02 = imem00_in[103:100];
    33: op1_01_in02 = reg_0830;
    34: op1_01_in02 = imem02_in[59:56];
    35: op1_01_in02 = imem00_in[83:80];
    37: op1_01_in02 = imem00_in[67:64];
    38: op1_01_in02 = imem02_in[111:108];
    39: op1_01_in02 = reg_0219;
    40: op1_01_in02 = reg_0311;
    41: op1_01_in02 = reg_0933;
    42: op1_01_in02 = reg_0495;
    45: op1_01_in02 = reg_0984;
    46: op1_01_in02 = reg_0633;
    47: op1_01_in02 = reg_0107;
    48: op1_01_in02 = reg_0872;
    49: op1_01_in02 = reg_0632;
    51: op1_01_in02 = reg_0407;
    52: op1_01_in02 = imem04_in[71:68];
    53: op1_01_in02 = reg_0976;
    54: op1_01_in02 = imem05_in[11:8];
    56: op1_01_in02 = imem07_in[123:120];
    57: op1_01_in02 = imem00_in[79:76];
    89: op1_01_in02 = imem00_in[79:76];
    58: op1_01_in02 = imem00_in[55:52];
    82: op1_01_in02 = imem00_in[55:52];
    59: op1_01_in02 = imem07_in[15:12];
    61: op1_01_in02 = imem00_in[71:68];
    62: op1_01_in02 = reg_0827;
    63: op1_01_in02 = reg_0041;
    64: op1_01_in02 = imem06_in[127:124];
    65: op1_01_in02 = reg_0264;
    66: op1_01_in02 = imem07_in[91:88];
    67: op1_01_in02 = reg_0955;
    68: op1_01_in02 = reg_0428;
    69: op1_01_in02 = reg_1007;
    70: op1_01_in02 = imem05_in[79:76];
    71: op1_01_in02 = imem00_in[27:24];
    72: op1_01_in02 = reg_0288;
    73: op1_01_in02 = reg_0720;
    74: op1_01_in02 = reg_0024;
    76: op1_01_in02 = reg_0112;
    77: op1_01_in02 = reg_0869;
    78: op1_01_in02 = reg_0524;
    79: op1_01_in02 = imem07_in[83:80];
    80: op1_01_in02 = reg_0270;
    81: op1_01_in02 = imem00_in[63:60];
    83: op1_01_in02 = reg_0948;
    84: op1_01_in02 = reg_0990;
    85: op1_01_in02 = reg_0141;
    87: op1_01_in02 = reg_0781;
    88: op1_01_in02 = reg_0259;
    90: op1_01_in02 = reg_0806;
    91: op1_01_in02 = imem07_in[3:0];
    92: op1_01_in02 = reg_0184;
    93: op1_01_in02 = reg_0346;
    94: op1_01_in02 = reg_0643;
    95: op1_01_in02 = reg_0643;
    96: op1_01_in02 = reg_0642;
    97: op1_01_in02 = reg_0520;
    default: op1_01_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_01_inv02 = 1;
    7: op1_01_inv02 = 1;
    8: op1_01_inv02 = 1;
    9: op1_01_inv02 = 1;
    11: op1_01_inv02 = 1;
    13: op1_01_inv02 = 1;
    2: op1_01_inv02 = 1;
    14: op1_01_inv02 = 1;
    15: op1_01_inv02 = 1;
    16: op1_01_inv02 = 1;
    17: op1_01_inv02 = 1;
    21: op1_01_inv02 = 1;
    22: op1_01_inv02 = 1;
    24: op1_01_inv02 = 1;
    25: op1_01_inv02 = 1;
    27: op1_01_inv02 = 1;
    28: op1_01_inv02 = 1;
    30: op1_01_inv02 = 1;
    32: op1_01_inv02 = 1;
    34: op1_01_inv02 = 1;
    37: op1_01_inv02 = 1;
    39: op1_01_inv02 = 1;
    40: op1_01_inv02 = 1;
    41: op1_01_inv02 = 1;
    50: op1_01_inv02 = 1;
    52: op1_01_inv02 = 1;
    53: op1_01_inv02 = 1;
    56: op1_01_inv02 = 1;
    57: op1_01_inv02 = 1;
    58: op1_01_inv02 = 1;
    60: op1_01_inv02 = 1;
    61: op1_01_inv02 = 1;
    62: op1_01_inv02 = 1;
    63: op1_01_inv02 = 1;
    65: op1_01_inv02 = 1;
    68: op1_01_inv02 = 1;
    71: op1_01_inv02 = 1;
    72: op1_01_inv02 = 1;
    75: op1_01_inv02 = 1;
    77: op1_01_inv02 = 1;
    79: op1_01_inv02 = 1;
    81: op1_01_inv02 = 1;
    82: op1_01_inv02 = 1;
    84: op1_01_inv02 = 1;
    85: op1_01_inv02 = 1;
    86: op1_01_inv02 = 1;
    88: op1_01_inv02 = 1;
    90: op1_01_inv02 = 1;
    92: op1_01_inv02 = 1;
    93: op1_01_inv02 = 1;
    97: op1_01_inv02 = 1;
    default: op1_01_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in03 = reg_0515;
    6: op1_01_in03 = reg_0617;
    7: op1_01_in03 = reg_0334;
    8: op1_01_in03 = reg_0132;
    4: op1_01_in03 = imem07_in[79:76];
    9: op1_01_in03 = imem00_in[79:76];
    3: op1_01_in03 = reg_0161;
    10: op1_01_in03 = reg_0342;
    11: op1_01_in03 = reg_0092;
    12: op1_01_in03 = reg_0689;
    13: op1_01_in03 = reg_0115;
    2: op1_01_in03 = imem07_in[39:36];
    14: op1_01_in03 = reg_0027;
    63: op1_01_in03 = reg_0027;
    15: op1_01_in03 = reg_1033;
    16: op1_01_in03 = imem02_in[123:120];
    17: op1_01_in03 = imem05_in[55:52];
    26: op1_01_in03 = imem05_in[55:52];
    18: op1_01_in03 = imem00_in[51:48];
    19: op1_01_in03 = reg_0704;
    20: op1_01_in03 = imem00_in[127:124];
    21: op1_01_in03 = reg_0528;
    22: op1_01_in03 = reg_0693;
    23: op1_01_in03 = imem02_in[127:124];
    24: op1_01_in03 = reg_0344;
    25: op1_01_in03 = imem03_in[91:88];
    27: op1_01_in03 = reg_0117;
    28: op1_01_in03 = reg_0954;
    31: op1_01_in03 = reg_0954;
    29: op1_01_in03 = reg_0671;
    30: op1_01_in03 = reg_0104;
    32: op1_01_in03 = imem00_in[111:108];
    33: op1_01_in03 = reg_0216;
    34: op1_01_in03 = imem02_in[115:112];
    38: op1_01_in03 = imem02_in[115:112];
    35: op1_01_in03 = imem00_in[99:96];
    37: op1_01_in03 = imem00_in[123:120];
    82: op1_01_in03 = imem00_in[123:120];
    39: op1_01_in03 = reg_0249;
    40: op1_01_in03 = reg_1002;
    41: op1_01_in03 = reg_0398;
    42: op1_01_in03 = reg_0387;
    43: op1_01_in03 = reg_0672;
    44: op1_01_in03 = reg_0101;
    45: op1_01_in03 = reg_0993;
    46: op1_01_in03 = reg_0029;
    47: op1_01_in03 = reg_0127;
    48: op1_01_in03 = imem03_in[59:56];
    49: op1_01_in03 = reg_0612;
    50: op1_01_in03 = imem07_in[87:84];
    59: op1_01_in03 = imem07_in[87:84];
    51: op1_01_in03 = reg_0533;
    52: op1_01_in03 = imem04_in[87:84];
    53: op1_01_in03 = imem04_in[3:0];
    54: op1_01_in03 = imem05_in[71:68];
    55: op1_01_in03 = reg_0967;
    56: op1_01_in03 = reg_0710;
    57: op1_01_in03 = imem00_in[83:80];
    89: op1_01_in03 = imem00_in[83:80];
    58: op1_01_in03 = imem00_in[63:60];
    60: op1_01_in03 = reg_0832;
    61: op1_01_in03 = imem00_in[87:84];
    62: op1_01_in03 = reg_0821;
    64: op1_01_in03 = reg_0010;
    65: op1_01_in03 = imem07_in[23:20];
    66: op1_01_in03 = imem07_in[95:92];
    67: op1_01_in03 = imem07_in[51:48];
    68: op1_01_in03 = reg_0420;
    69: op1_01_in03 = reg_0580;
    70: op1_01_in03 = imem05_in[119:116];
    71: op1_01_in03 = imem00_in[67:64];
    72: op1_01_in03 = reg_0764;
    73: op1_01_in03 = reg_0721;
    74: op1_01_in03 = reg_0180;
    75: op1_01_in03 = imem00_in[35:32];
    76: op1_01_in03 = imem02_in[3:0];
    77: op1_01_in03 = reg_0604;
    78: op1_01_in03 = reg_0067;
    79: op1_01_in03 = imem07_in[99:96];
    80: op1_01_in03 = reg_0915;
    81: op1_01_in03 = reg_0825;
    83: op1_01_in03 = reg_0892;
    84: op1_01_in03 = reg_0983;
    85: op1_01_in03 = reg_0958;
    86: op1_01_in03 = reg_0674;
    87: op1_01_in03 = reg_0857;
    88: op1_01_in03 = reg_0675;
    90: op1_01_in03 = reg_0706;
    91: op1_01_in03 = imem07_in[15:12];
    93: op1_01_in03 = reg_0662;
    94: op1_01_in03 = imem03_in[39:36];
    95: op1_01_in03 = reg_0367;
    96: op1_01_in03 = reg_0323;
    97: op1_01_in03 = reg_0064;
    default: op1_01_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_01_inv03 = 1;
    10: op1_01_inv03 = 1;
    13: op1_01_inv03 = 1;
    14: op1_01_inv03 = 1;
    16: op1_01_inv03 = 1;
    20: op1_01_inv03 = 1;
    22: op1_01_inv03 = 1;
    23: op1_01_inv03 = 1;
    24: op1_01_inv03 = 1;
    25: op1_01_inv03 = 1;
    27: op1_01_inv03 = 1;
    28: op1_01_inv03 = 1;
    29: op1_01_inv03 = 1;
    34: op1_01_inv03 = 1;
    38: op1_01_inv03 = 1;
    40: op1_01_inv03 = 1;
    41: op1_01_inv03 = 1;
    42: op1_01_inv03 = 1;
    45: op1_01_inv03 = 1;
    47: op1_01_inv03 = 1;
    51: op1_01_inv03 = 1;
    54: op1_01_inv03 = 1;
    57: op1_01_inv03 = 1;
    61: op1_01_inv03 = 1;
    62: op1_01_inv03 = 1;
    63: op1_01_inv03 = 1;
    64: op1_01_inv03 = 1;
    65: op1_01_inv03 = 1;
    68: op1_01_inv03 = 1;
    71: op1_01_inv03 = 1;
    72: op1_01_inv03 = 1;
    73: op1_01_inv03 = 1;
    74: op1_01_inv03 = 1;
    75: op1_01_inv03 = 1;
    76: op1_01_inv03 = 1;
    77: op1_01_inv03 = 1;
    78: op1_01_inv03 = 1;
    79: op1_01_inv03 = 1;
    82: op1_01_inv03 = 1;
    85: op1_01_inv03 = 1;
    86: op1_01_inv03 = 1;
    88: op1_01_inv03 = 1;
    96: op1_01_inv03 = 1;
    97: op1_01_inv03 = 1;
    default: op1_01_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in04 = reg_0498;
    6: op1_01_in04 = reg_0605;
    7: op1_01_in04 = reg_0357;
    8: op1_01_in04 = reg_0147;
    4: op1_01_in04 = imem07_in[83:80];
    9: op1_01_in04 = imem00_in[111:108];
    3: op1_01_in04 = reg_0169;
    10: op1_01_in04 = reg_0350;
    11: op1_01_in04 = reg_0045;
    12: op1_01_in04 = reg_0684;
    13: op1_01_in04 = reg_0113;
    47: op1_01_in04 = reg_0113;
    2: op1_01_in04 = imem07_in[63:60];
    14: op1_01_in04 = reg_0486;
    15: op1_01_in04 = reg_0830;
    16: op1_01_in04 = imem02_in[127:124];
    17: op1_01_in04 = imem05_in[63:60];
    18: op1_01_in04 = imem00_in[59:56];
    19: op1_01_in04 = reg_0702;
    20: op1_01_in04 = reg_0681;
    21: op1_01_in04 = reg_0286;
    22: op1_01_in04 = reg_0683;
    23: op1_01_in04 = reg_0654;
    24: op1_01_in04 = reg_0372;
    25: op1_01_in04 = reg_0586;
    26: op1_01_in04 = imem05_in[119:116];
    27: op1_01_in04 = reg_0110;
    60: op1_01_in04 = reg_0110;
    28: op1_01_in04 = reg_0969;
    55: op1_01_in04 = reg_0969;
    29: op1_01_in04 = reg_0678;
    30: op1_01_in04 = reg_0115;
    31: op1_01_in04 = reg_0949;
    32: op1_01_in04 = imem00_in[115:112];
    33: op1_01_in04 = reg_1035;
    34: op1_01_in04 = imem02_in[119:116];
    38: op1_01_in04 = imem02_in[119:116];
    35: op1_01_in04 = reg_0697;
    37: op1_01_in04 = reg_0695;
    39: op1_01_in04 = reg_1043;
    40: op1_01_in04 = imem04_in[43:40];
    41: op1_01_in04 = reg_0580;
    42: op1_01_in04 = reg_0381;
    51: op1_01_in04 = reg_0381;
    43: op1_01_in04 = reg_0679;
    44: op1_01_in04 = reg_0117;
    45: op1_01_in04 = reg_0976;
    46: op1_01_in04 = reg_0622;
    48: op1_01_in04 = imem03_in[67:64];
    49: op1_01_in04 = reg_0385;
    50: op1_01_in04 = reg_0717;
    52: op1_01_in04 = imem04_in[91:88];
    53: op1_01_in04 = imem04_in[11:8];
    54: op1_01_in04 = imem05_in[87:84];
    56: op1_01_in04 = reg_0729;
    57: op1_01_in04 = imem00_in[91:88];
    89: op1_01_in04 = imem00_in[91:88];
    58: op1_01_in04 = imem00_in[71:68];
    71: op1_01_in04 = imem00_in[71:68];
    59: op1_01_in04 = reg_0728;
    61: op1_01_in04 = reg_0671;
    62: op1_01_in04 = reg_0745;
    63: op1_01_in04 = reg_0409;
    64: op1_01_in04 = reg_0344;
    65: op1_01_in04 = imem07_in[119:116];
    79: op1_01_in04 = imem07_in[119:116];
    66: op1_01_in04 = imem07_in[107:104];
    67: op1_01_in04 = imem07_in[59:56];
    68: op1_01_in04 = reg_0174;
    69: op1_01_in04 = reg_0445;
    70: op1_01_in04 = reg_0655;
    72: op1_01_in04 = reg_0658;
    73: op1_01_in04 = reg_0723;
    74: op1_01_in04 = reg_0162;
    75: op1_01_in04 = imem00_in[39:36];
    76: op1_01_in04 = imem02_in[23:20];
    77: op1_01_in04 = reg_0860;
    78: op1_01_in04 = reg_0296;
    80: op1_01_in04 = reg_0755;
    81: op1_01_in04 = reg_0900;
    82: op1_01_in04 = reg_0841;
    83: op1_01_in04 = reg_0957;
    84: op1_01_in04 = imem04_in[3:0];
    85: op1_01_in04 = reg_0223;
    86: op1_01_in04 = reg_0668;
    87: op1_01_in04 = reg_0293;
    88: op1_01_in04 = reg_0892;
    90: op1_01_in04 = imem06_in[7:4];
    91: op1_01_in04 = imem07_in[19:16];
    93: op1_01_in04 = reg_0623;
    94: op1_01_in04 = imem03_in[43:40];
    95: op1_01_in04 = imem03_in[11:8];
    96: op1_01_in04 = reg_0039;
    97: op1_01_in04 = reg_0904;
    default: op1_01_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv04 = 1;
    3: op1_01_inv04 = 1;
    12: op1_01_inv04 = 1;
    13: op1_01_inv04 = 1;
    2: op1_01_inv04 = 1;
    14: op1_01_inv04 = 1;
    16: op1_01_inv04 = 1;
    18: op1_01_inv04 = 1;
    19: op1_01_inv04 = 1;
    20: op1_01_inv04 = 1;
    23: op1_01_inv04 = 1;
    26: op1_01_inv04 = 1;
    28: op1_01_inv04 = 1;
    31: op1_01_inv04 = 1;
    35: op1_01_inv04 = 1;
    40: op1_01_inv04 = 1;
    41: op1_01_inv04 = 1;
    43: op1_01_inv04 = 1;
    44: op1_01_inv04 = 1;
    45: op1_01_inv04 = 1;
    48: op1_01_inv04 = 1;
    49: op1_01_inv04 = 1;
    50: op1_01_inv04 = 1;
    51: op1_01_inv04 = 1;
    54: op1_01_inv04 = 1;
    55: op1_01_inv04 = 1;
    58: op1_01_inv04 = 1;
    59: op1_01_inv04 = 1;
    60: op1_01_inv04 = 1;
    64: op1_01_inv04 = 1;
    65: op1_01_inv04 = 1;
    66: op1_01_inv04 = 1;
    67: op1_01_inv04 = 1;
    70: op1_01_inv04 = 1;
    73: op1_01_inv04 = 1;
    75: op1_01_inv04 = 1;
    76: op1_01_inv04 = 1;
    78: op1_01_inv04 = 1;
    79: op1_01_inv04 = 1;
    80: op1_01_inv04 = 1;
    86: op1_01_inv04 = 1;
    90: op1_01_inv04 = 1;
    91: op1_01_inv04 = 1;
    93: op1_01_inv04 = 1;
    95: op1_01_inv04 = 1;
    96: op1_01_inv04 = 1;
    97: op1_01_inv04 = 1;
    default: op1_01_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in05 = reg_0232;
    6: op1_01_in05 = reg_0626;
    7: op1_01_in05 = reg_0346;
    41: op1_01_in05 = reg_0346;
    8: op1_01_in05 = reg_0149;
    4: op1_01_in05 = imem07_in[119:116];
    9: op1_01_in05 = imem00_in[115:112];
    3: op1_01_in05 = reg_0183;
    10: op1_01_in05 = reg_0081;
    11: op1_01_in05 = reg_0087;
    12: op1_01_in05 = reg_0686;
    13: op1_01_in05 = reg_0121;
    44: op1_01_in05 = reg_0121;
    14: op1_01_in05 = reg_0805;
    15: op1_01_in05 = reg_1031;
    16: op1_01_in05 = reg_0658;
    17: op1_01_in05 = imem05_in[83:80];
    18: op1_01_in05 = imem00_in[95:92];
    89: op1_01_in05 = imem00_in[95:92];
    19: op1_01_in05 = reg_0708;
    20: op1_01_in05 = reg_0696;
    21: op1_01_in05 = reg_0044;
    22: op1_01_in05 = reg_0685;
    37: op1_01_in05 = reg_0685;
    23: op1_01_in05 = reg_0640;
    24: op1_01_in05 = reg_0337;
    25: op1_01_in05 = reg_0587;
    26: op1_01_in05 = reg_0973;
    27: op1_01_in05 = imem02_in[15:12];
    28: op1_01_in05 = reg_0964;
    29: op1_01_in05 = reg_0675;
    30: op1_01_in05 = reg_0107;
    31: op1_01_in05 = reg_0965;
    32: op1_01_in05 = reg_0693;
    33: op1_01_in05 = reg_0913;
    34: op1_01_in05 = imem02_in[123:120];
    35: op1_01_in05 = reg_0676;
    38: op1_01_in05 = reg_0645;
    39: op1_01_in05 = reg_0227;
    40: op1_01_in05 = imem04_in[47:44];
    42: op1_01_in05 = reg_0042;
    43: op1_01_in05 = reg_0691;
    45: op1_01_in05 = reg_0997;
    46: op1_01_in05 = imem07_in[23:20];
    47: op1_01_in05 = imem02_in[7:4];
    48: op1_01_in05 = imem03_in[91:88];
    49: op1_01_in05 = reg_0293;
    50: op1_01_in05 = reg_0718;
    51: op1_01_in05 = reg_0395;
    52: op1_01_in05 = imem04_in[123:120];
    53: op1_01_in05 = imem04_in[31:28];
    54: op1_01_in05 = imem05_in[103:100];
    55: op1_01_in05 = reg_0972;
    56: op1_01_in05 = reg_0705;
    57: op1_01_in05 = imem00_in[107:104];
    58: op1_01_in05 = imem00_in[107:104];
    59: op1_01_in05 = reg_0720;
    60: op1_01_in05 = imem02_in[27:24];
    61: op1_01_in05 = reg_0842;
    62: op1_01_in05 = imem02_in[19:16];
    63: op1_01_in05 = reg_0332;
    64: op1_01_in05 = reg_0817;
    65: op1_01_in05 = imem07_in[123:120];
    66: op1_01_in05 = imem07_in[127:124];
    79: op1_01_in05 = imem07_in[127:124];
    67: op1_01_in05 = imem07_in[99:96];
    68: op1_01_in05 = reg_0175;
    69: op1_01_in05 = reg_0327;
    70: op1_01_in05 = reg_0963;
    71: op1_01_in05 = imem00_in[99:96];
    72: op1_01_in05 = reg_0777;
    73: op1_01_in05 = reg_0714;
    74: op1_01_in05 = reg_0167;
    75: op1_01_in05 = imem00_in[71:68];
    76: op1_01_in05 = imem02_in[103:100];
    77: op1_01_in05 = reg_0827;
    78: op1_01_in05 = reg_0432;
    80: op1_01_in05 = reg_0320;
    81: op1_01_in05 = reg_0478;
    82: op1_01_in05 = reg_0738;
    83: op1_01_in05 = reg_0943;
    84: op1_01_in05 = imem04_in[19:16];
    85: op1_01_in05 = reg_0265;
    86: op1_01_in05 = reg_0669;
    87: op1_01_in05 = reg_0026;
    88: op1_01_in05 = reg_0436;
    90: op1_01_in05 = imem06_in[23:20];
    91: op1_01_in05 = imem07_in[27:24];
    93: op1_01_in05 = reg_0596;
    94: op1_01_in05 = imem03_in[47:44];
    95: op1_01_in05 = imem03_in[39:36];
    96: op1_01_in05 = reg_0425;
    97: op1_01_in05 = reg_1022;
    default: op1_01_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_01_inv05 = 1;
    14: op1_01_inv05 = 1;
    16: op1_01_inv05 = 1;
    18: op1_01_inv05 = 1;
    19: op1_01_inv05 = 1;
    21: op1_01_inv05 = 1;
    25: op1_01_inv05 = 1;
    27: op1_01_inv05 = 1;
    28: op1_01_inv05 = 1;
    29: op1_01_inv05 = 1;
    30: op1_01_inv05 = 1;
    31: op1_01_inv05 = 1;
    34: op1_01_inv05 = 1;
    35: op1_01_inv05 = 1;
    37: op1_01_inv05 = 1;
    38: op1_01_inv05 = 1;
    39: op1_01_inv05 = 1;
    40: op1_01_inv05 = 1;
    41: op1_01_inv05 = 1;
    43: op1_01_inv05 = 1;
    45: op1_01_inv05 = 1;
    46: op1_01_inv05 = 1;
    47: op1_01_inv05 = 1;
    48: op1_01_inv05 = 1;
    49: op1_01_inv05 = 1;
    50: op1_01_inv05 = 1;
    56: op1_01_inv05 = 1;
    58: op1_01_inv05 = 1;
    61: op1_01_inv05 = 1;
    67: op1_01_inv05 = 1;
    68: op1_01_inv05 = 1;
    69: op1_01_inv05 = 1;
    70: op1_01_inv05 = 1;
    72: op1_01_inv05 = 1;
    73: op1_01_inv05 = 1;
    75: op1_01_inv05 = 1;
    76: op1_01_inv05 = 1;
    80: op1_01_inv05 = 1;
    82: op1_01_inv05 = 1;
    83: op1_01_inv05 = 1;
    85: op1_01_inv05 = 1;
    87: op1_01_inv05 = 1;
    89: op1_01_inv05 = 1;
    90: op1_01_inv05 = 1;
    91: op1_01_inv05 = 1;
    93: op1_01_inv05 = 1;
    96: op1_01_inv05 = 1;
    97: op1_01_inv05 = 1;
    default: op1_01_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in06 = reg_0226;
    6: op1_01_in06 = reg_0627;
    7: op1_01_in06 = reg_0324;
    8: op1_01_in06 = reg_0153;
    4: op1_01_in06 = imem07_in[123:120];
    9: op1_01_in06 = reg_0682;
    3: op1_01_in06 = reg_0178;
    10: op1_01_in06 = reg_0095;
    11: op1_01_in06 = reg_0093;
    12: op1_01_in06 = reg_0679;
    13: op1_01_in06 = imem02_in[23:20];
    14: op1_01_in06 = imem07_in[3:0];
    15: op1_01_in06 = reg_0913;
    16: op1_01_in06 = reg_0358;
    17: op1_01_in06 = imem05_in[95:92];
    18: op1_01_in06 = imem00_in[127:124];
    71: op1_01_in06 = imem00_in[127:124];
    19: op1_01_in06 = reg_0715;
    20: op1_01_in06 = reg_0688;
    43: op1_01_in06 = reg_0688;
    21: op1_01_in06 = imem05_in[7:4];
    22: op1_01_in06 = reg_0684;
    23: op1_01_in06 = reg_0641;
    24: op1_01_in06 = reg_1029;
    25: op1_01_in06 = reg_0592;
    26: op1_01_in06 = reg_0955;
    27: op1_01_in06 = imem02_in[43:40];
    28: op1_01_in06 = reg_0949;
    29: op1_01_in06 = reg_0692;
    30: op1_01_in06 = reg_0126;
    31: op1_01_in06 = reg_0961;
    32: op1_01_in06 = reg_0697;
    33: op1_01_in06 = reg_1036;
    34: op1_01_in06 = reg_0637;
    35: op1_01_in06 = reg_0698;
    37: op1_01_in06 = reg_0677;
    38: op1_01_in06 = reg_0658;
    39: op1_01_in06 = reg_0216;
    40: op1_01_in06 = imem04_in[55:52];
    41: op1_01_in06 = reg_0823;
    42: op1_01_in06 = reg_0392;
    44: op1_01_in06 = imem02_in[7:4];
    45: op1_01_in06 = imem04_in[35:32];
    46: op1_01_in06 = imem07_in[43:40];
    47: op1_01_in06 = imem02_in[55:52];
    48: op1_01_in06 = imem03_in[127:124];
    49: op1_01_in06 = reg_0356;
    50: op1_01_in06 = reg_0711;
    51: op1_01_in06 = reg_0386;
    52: op1_01_in06 = reg_0536;
    53: op1_01_in06 = imem04_in[47:44];
    54: op1_01_in06 = imem05_in[127:124];
    55: op1_01_in06 = reg_0032;
    56: op1_01_in06 = reg_0713;
    57: op1_01_in06 = imem00_in[115:112];
    58: op1_01_in06 = reg_0900;
    59: op1_01_in06 = reg_0731;
    60: op1_01_in06 = imem02_in[87:84];
    61: op1_01_in06 = reg_0463;
    62: op1_01_in06 = imem02_in[47:44];
    63: op1_01_in06 = imem05_in[27:24];
    64: op1_01_in06 = reg_0439;
    65: op1_01_in06 = reg_0704;
    66: op1_01_in06 = reg_0730;
    67: op1_01_in06 = imem07_in[103:100];
    68: op1_01_in06 = reg_0163;
    69: op1_01_in06 = reg_0662;
    70: op1_01_in06 = reg_0784;
    72: op1_01_in06 = imem05_in[63:60];
    73: op1_01_in06 = reg_0718;
    74: op1_01_in06 = reg_0169;
    75: op1_01_in06 = reg_0841;
    76: op1_01_in06 = imem02_in[107:104];
    77: op1_01_in06 = imem02_in[3:0];
    78: op1_01_in06 = reg_0407;
    79: op1_01_in06 = reg_0426;
    80: op1_01_in06 = imem07_in[39:36];
    81: op1_01_in06 = reg_0214;
    82: op1_01_in06 = reg_0828;
    83: op1_01_in06 = reg_0707;
    84: op1_01_in06 = imem04_in[43:40];
    85: op1_01_in06 = reg_0952;
    86: op1_01_in06 = reg_0455;
    87: op1_01_in06 = reg_0834;
    88: op1_01_in06 = reg_0617;
    89: op1_01_in06 = imem00_in[119:116];
    90: op1_01_in06 = imem06_in[43:40];
    91: op1_01_in06 = imem07_in[59:56];
    93: op1_01_in06 = reg_0239;
    94: op1_01_in06 = imem03_in[67:64];
    95: op1_01_in06 = imem03_in[91:88];
    96: op1_01_in06 = reg_0054;
    97: op1_01_in06 = reg_0104;
    default: op1_01_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv06 = 1;
    7: op1_01_inv06 = 1;
    8: op1_01_inv06 = 1;
    4: op1_01_inv06 = 1;
    9: op1_01_inv06 = 1;
    3: op1_01_inv06 = 1;
    13: op1_01_inv06 = 1;
    14: op1_01_inv06 = 1;
    19: op1_01_inv06 = 1;
    23: op1_01_inv06 = 1;
    26: op1_01_inv06 = 1;
    28: op1_01_inv06 = 1;
    31: op1_01_inv06 = 1;
    32: op1_01_inv06 = 1;
    38: op1_01_inv06 = 1;
    39: op1_01_inv06 = 1;
    41: op1_01_inv06 = 1;
    45: op1_01_inv06 = 1;
    50: op1_01_inv06 = 1;
    51: op1_01_inv06 = 1;
    52: op1_01_inv06 = 1;
    53: op1_01_inv06 = 1;
    54: op1_01_inv06 = 1;
    55: op1_01_inv06 = 1;
    57: op1_01_inv06 = 1;
    61: op1_01_inv06 = 1;
    62: op1_01_inv06 = 1;
    63: op1_01_inv06 = 1;
    64: op1_01_inv06 = 1;
    65: op1_01_inv06 = 1;
    66: op1_01_inv06 = 1;
    68: op1_01_inv06 = 1;
    72: op1_01_inv06 = 1;
    73: op1_01_inv06 = 1;
    75: op1_01_inv06 = 1;
    77: op1_01_inv06 = 1;
    79: op1_01_inv06 = 1;
    81: op1_01_inv06 = 1;
    83: op1_01_inv06 = 1;
    84: op1_01_inv06 = 1;
    86: op1_01_inv06 = 1;
    88: op1_01_inv06 = 1;
    89: op1_01_inv06 = 1;
    93: op1_01_inv06 = 1;
    94: op1_01_inv06 = 1;
    95: op1_01_inv06 = 1;
    default: op1_01_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in07 = reg_0233;
    6: op1_01_in07 = reg_0348;
    7: op1_01_in07 = reg_0342;
    8: op1_01_in07 = reg_0140;
    4: op1_01_in07 = reg_0425;
    9: op1_01_in07 = reg_0693;
    3: op1_01_in07 = reg_0157;
    10: op1_01_in07 = reg_0060;
    11: op1_01_in07 = reg_0073;
    12: op1_01_in07 = reg_0677;
    13: op1_01_in07 = imem02_in[39:36];
    14: op1_01_in07 = imem07_in[15:12];
    15: op1_01_in07 = reg_0871;
    16: op1_01_in07 = reg_0364;
    17: op1_01_in07 = reg_0973;
    18: op1_01_in07 = reg_0698;
    19: op1_01_in07 = reg_0701;
    20: op1_01_in07 = reg_0692;
    21: op1_01_in07 = imem05_in[19:16];
    22: op1_01_in07 = reg_0690;
    23: op1_01_in07 = reg_0320;
    24: op1_01_in07 = reg_0752;
    25: op1_01_in07 = reg_0585;
    26: op1_01_in07 = reg_0964;
    27: op1_01_in07 = imem02_in[107:104];
    28: op1_01_in07 = reg_1021;
    29: op1_01_in07 = reg_0465;
    58: op1_01_in07 = reg_0465;
    30: op1_01_in07 = imem02_in[11:8];
    31: op1_01_in07 = reg_0953;
    32: op1_01_in07 = reg_0674;
    33: op1_01_in07 = reg_1038;
    34: op1_01_in07 = reg_0660;
    35: op1_01_in07 = reg_0679;
    37: op1_01_in07 = reg_0450;
    38: op1_01_in07 = reg_0656;
    39: op1_01_in07 = reg_1045;
    40: op1_01_in07 = imem04_in[71:68];
    41: op1_01_in07 = reg_0370;
    42: op1_01_in07 = reg_0391;
    43: op1_01_in07 = reg_0453;
    61: op1_01_in07 = reg_0453;
    44: op1_01_in07 = imem02_in[23:20];
    45: op1_01_in07 = imem04_in[87:84];
    46: op1_01_in07 = imem07_in[47:44];
    47: op1_01_in07 = imem02_in[99:96];
    48: op1_01_in07 = reg_0006;
    49: op1_01_in07 = reg_0395;
    50: op1_01_in07 = reg_0706;
    51: op1_01_in07 = reg_0741;
    52: op1_01_in07 = reg_0937;
    53: op1_01_in07 = imem04_in[107:104];
    54: op1_01_in07 = reg_0966;
    55: op1_01_in07 = reg_0094;
    56: op1_01_in07 = reg_0303;
    57: op1_01_in07 = reg_0001;
    89: op1_01_in07 = reg_0001;
    59: op1_01_in07 = reg_0721;
    60: op1_01_in07 = imem02_in[119:116];
    62: op1_01_in07 = imem02_in[91:88];
    63: op1_01_in07 = imem05_in[47:44];
    64: op1_01_in07 = reg_0695;
    65: op1_01_in07 = reg_0719;
    66: op1_01_in07 = reg_0723;
    67: op1_01_in07 = imem07_in[115:112];
    68: op1_01_in07 = reg_0176;
    69: op1_01_in07 = reg_0923;
    70: op1_01_in07 = reg_0865;
    71: op1_01_in07 = reg_0683;
    72: op1_01_in07 = imem05_in[67:64];
    73: op1_01_in07 = reg_0727;
    74: op1_01_in07 = reg_0166;
    75: op1_01_in07 = reg_0523;
    76: op1_01_in07 = reg_0916;
    77: op1_01_in07 = imem02_in[15:12];
    78: op1_01_in07 = reg_0243;
    79: op1_01_in07 = reg_0641;
    80: op1_01_in07 = imem07_in[79:76];
    81: op1_01_in07 = reg_0191;
    82: op1_01_in07 = reg_0687;
    83: op1_01_in07 = reg_0816;
    84: op1_01_in07 = imem04_in[51:48];
    85: op1_01_in07 = reg_0943;
    86: op1_01_in07 = reg_0481;
    87: op1_01_in07 = reg_0612;
    88: op1_01_in07 = reg_0707;
    90: op1_01_in07 = imem06_in[71:68];
    91: op1_01_in07 = imem07_in[67:64];
    93: op1_01_in07 = reg_0377;
    94: op1_01_in07 = imem03_in[75:72];
    95: op1_01_in07 = imem03_in[99:96];
    96: op1_01_in07 = reg_0085;
    97: op1_01_in07 = reg_0398;
    default: op1_01_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv07 = 1;
    6: op1_01_inv07 = 1;
    4: op1_01_inv07 = 1;
    10: op1_01_inv07 = 1;
    13: op1_01_inv07 = 1;
    16: op1_01_inv07 = 1;
    17: op1_01_inv07 = 1;
    18: op1_01_inv07 = 1;
    19: op1_01_inv07 = 1;
    24: op1_01_inv07 = 1;
    25: op1_01_inv07 = 1;
    29: op1_01_inv07 = 1;
    32: op1_01_inv07 = 1;
    35: op1_01_inv07 = 1;
    37: op1_01_inv07 = 1;
    38: op1_01_inv07 = 1;
    42: op1_01_inv07 = 1;
    43: op1_01_inv07 = 1;
    44: op1_01_inv07 = 1;
    45: op1_01_inv07 = 1;
    50: op1_01_inv07 = 1;
    51: op1_01_inv07 = 1;
    52: op1_01_inv07 = 1;
    53: op1_01_inv07 = 1;
    54: op1_01_inv07 = 1;
    55: op1_01_inv07 = 1;
    57: op1_01_inv07 = 1;
    59: op1_01_inv07 = 1;
    66: op1_01_inv07 = 1;
    67: op1_01_inv07 = 1;
    69: op1_01_inv07 = 1;
    71: op1_01_inv07 = 1;
    72: op1_01_inv07 = 1;
    73: op1_01_inv07 = 1;
    74: op1_01_inv07 = 1;
    76: op1_01_inv07 = 1;
    78: op1_01_inv07 = 1;
    79: op1_01_inv07 = 1;
    80: op1_01_inv07 = 1;
    81: op1_01_inv07 = 1;
    82: op1_01_inv07 = 1;
    83: op1_01_inv07 = 1;
    85: op1_01_inv07 = 1;
    91: op1_01_inv07 = 1;
    94: op1_01_inv07 = 1;
    97: op1_01_inv07 = 1;
    default: op1_01_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in08 = reg_0218;
    6: op1_01_in08 = reg_0386;
    7: op1_01_in08 = reg_0338;
    8: op1_01_in08 = imem06_in[7:4];
    4: op1_01_in08 = reg_0418;
    9: op1_01_in08 = reg_0697;
    3: op1_01_in08 = reg_0171;
    10: op1_01_in08 = reg_0094;
    11: op1_01_in08 = imem03_in[31:28];
    12: op1_01_in08 = reg_0688;
    13: op1_01_in08 = imem02_in[51:48];
    14: op1_01_in08 = imem07_in[23:20];
    15: op1_01_in08 = reg_1018;
    16: op1_01_in08 = reg_0324;
    17: op1_01_in08 = reg_0966;
    18: op1_01_in08 = reg_0670;
    19: op1_01_in08 = reg_0441;
    20: op1_01_in08 = reg_0669;
    21: op1_01_in08 = imem05_in[31:28];
    22: op1_01_in08 = reg_0677;
    23: op1_01_in08 = reg_0326;
    83: op1_01_in08 = reg_0326;
    24: op1_01_in08 = reg_0780;
    49: op1_01_in08 = reg_0780;
    25: op1_01_in08 = reg_0570;
    26: op1_01_in08 = reg_0947;
    70: op1_01_in08 = reg_0947;
    27: op1_01_in08 = imem02_in[119:116];
    28: op1_01_in08 = reg_0835;
    29: op1_01_in08 = reg_0451;
    30: op1_01_in08 = imem02_in[43:40];
    44: op1_01_in08 = imem02_in[43:40];
    31: op1_01_in08 = reg_1021;
    32: op1_01_in08 = reg_0678;
    33: op1_01_in08 = reg_0108;
    34: op1_01_in08 = reg_0647;
    38: op1_01_in08 = reg_0647;
    35: op1_01_in08 = reg_0680;
    37: op1_01_in08 = reg_0462;
    39: op1_01_in08 = reg_0122;
    40: op1_01_in08 = reg_0530;
    41: op1_01_in08 = reg_0038;
    42: op1_01_in08 = reg_0384;
    43: op1_01_in08 = reg_0454;
    45: op1_01_in08 = imem04_in[95:92];
    46: op1_01_in08 = imem07_in[75:72];
    47: op1_01_in08 = imem02_in[107:104];
    48: op1_01_in08 = reg_0343;
    50: op1_01_in08 = reg_0422;
    51: op1_01_in08 = reg_0349;
    52: op1_01_in08 = reg_1009;
    53: op1_01_in08 = imem04_in[123:120];
    54: op1_01_in08 = reg_0955;
    55: op1_01_in08 = reg_0448;
    56: op1_01_in08 = reg_0250;
    57: op1_01_in08 = reg_0825;
    58: op1_01_in08 = reg_0476;
    59: op1_01_in08 = reg_0714;
    60: op1_01_in08 = imem02_in[123:120];
    61: op1_01_in08 = reg_0457;
    62: op1_01_in08 = imem02_in[115:112];
    63: op1_01_in08 = imem05_in[79:76];
    64: op1_01_in08 = reg_0293;
    65: op1_01_in08 = reg_0730;
    66: op1_01_in08 = reg_0712;
    67: op1_01_in08 = reg_0722;
    68: op1_01_in08 = reg_0158;
    69: op1_01_in08 = reg_0369;
    71: op1_01_in08 = reg_0668;
    72: op1_01_in08 = reg_0693;
    73: op1_01_in08 = reg_0047;
    74: op1_01_in08 = reg_0164;
    75: op1_01_in08 = reg_0842;
    76: op1_01_in08 = reg_0762;
    77: op1_01_in08 = imem02_in[75:72];
    78: op1_01_in08 = reg_0044;
    79: op1_01_in08 = reg_0350;
    80: op1_01_in08 = imem07_in[115:112];
    81: op1_01_in08 = reg_0212;
    82: op1_01_in08 = reg_0663;
    84: op1_01_in08 = imem04_in[67:64];
    85: op1_01_in08 = reg_0819;
    86: op1_01_in08 = reg_0471;
    87: op1_01_in08 = reg_0017;
    88: op1_01_in08 = reg_0019;
    89: op1_01_in08 = reg_0463;
    90: op1_01_in08 = imem06_in[95:92];
    91: op1_01_in08 = imem07_in[83:80];
    93: op1_01_in08 = reg_0767;
    94: op1_01_in08 = imem03_in[83:80];
    95: op1_01_in08 = imem03_in[107:104];
    96: op1_01_in08 = reg_0381;
    97: op1_01_in08 = reg_0120;
    default: op1_01_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv08 = 1;
    10: op1_01_inv08 = 1;
    15: op1_01_inv08 = 1;
    22: op1_01_inv08 = 1;
    25: op1_01_inv08 = 1;
    26: op1_01_inv08 = 1;
    29: op1_01_inv08 = 1;
    32: op1_01_inv08 = 1;
    33: op1_01_inv08 = 1;
    40: op1_01_inv08 = 1;
    41: op1_01_inv08 = 1;
    44: op1_01_inv08 = 1;
    48: op1_01_inv08 = 1;
    49: op1_01_inv08 = 1;
    52: op1_01_inv08 = 1;
    54: op1_01_inv08 = 1;
    56: op1_01_inv08 = 1;
    59: op1_01_inv08 = 1;
    66: op1_01_inv08 = 1;
    68: op1_01_inv08 = 1;
    69: op1_01_inv08 = 1;
    71: op1_01_inv08 = 1;
    75: op1_01_inv08 = 1;
    78: op1_01_inv08 = 1;
    79: op1_01_inv08 = 1;
    80: op1_01_inv08 = 1;
    82: op1_01_inv08 = 1;
    85: op1_01_inv08 = 1;
    89: op1_01_inv08 = 1;
    91: op1_01_inv08 = 1;
    94: op1_01_inv08 = 1;
    97: op1_01_inv08 = 1;
    default: op1_01_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in09 = reg_0234;
    6: op1_01_in09 = reg_0033;
    7: op1_01_in09 = reg_0355;
    8: op1_01_in09 = imem06_in[15:12];
    4: op1_01_in09 = reg_0428;
    73: op1_01_in09 = reg_0428;
    9: op1_01_in09 = reg_0698;
    10: op1_01_in09 = imem03_in[15:12];
    11: op1_01_in09 = imem03_in[59:56];
    12: op1_01_in09 = reg_0463;
    13: op1_01_in09 = imem02_in[107:104];
    14: op1_01_in09 = imem07_in[43:40];
    15: op1_01_in09 = reg_0904;
    16: op1_01_in09 = reg_0338;
    17: op1_01_in09 = reg_0969;
    18: op1_01_in09 = reg_0679;
    19: op1_01_in09 = reg_0446;
    20: op1_01_in09 = reg_0454;
    21: op1_01_in09 = imem05_in[63:60];
    22: op1_01_in09 = reg_0674;
    23: op1_01_in09 = reg_0359;
    24: op1_01_in09 = reg_0798;
    25: op1_01_in09 = reg_0360;
    26: op1_01_in09 = reg_0900;
    28: op1_01_in09 = reg_0900;
    27: op1_01_in09 = reg_0661;
    29: op1_01_in09 = reg_0472;
    30: op1_01_in09 = imem02_in[59:56];
    31: op1_01_in09 = reg_0826;
    32: op1_01_in09 = reg_0688;
    33: op1_01_in09 = imem02_in[23:20];
    34: op1_01_in09 = reg_0659;
    35: op1_01_in09 = reg_0450;
    37: op1_01_in09 = reg_0481;
    38: op1_01_in09 = reg_0640;
    39: op1_01_in09 = reg_0116;
    40: op1_01_in09 = reg_1009;
    41: op1_01_in09 = reg_0040;
    42: op1_01_in09 = reg_0626;
    43: op1_01_in09 = reg_0451;
    44: op1_01_in09 = imem02_in[47:44];
    45: op1_01_in09 = imem04_in[115:112];
    46: op1_01_in09 = imem07_in[115:112];
    47: op1_01_in09 = reg_0363;
    60: op1_01_in09 = reg_0363;
    48: op1_01_in09 = reg_0046;
    49: op1_01_in09 = reg_0605;
    50: op1_01_in09 = reg_0174;
    51: op1_01_in09 = reg_0384;
    52: op1_01_in09 = reg_1020;
    53: op1_01_in09 = reg_0530;
    54: op1_01_in09 = reg_0954;
    55: op1_01_in09 = reg_0333;
    56: op1_01_in09 = reg_0321;
    57: op1_01_in09 = reg_0842;
    58: op1_01_in09 = reg_0462;
    59: op1_01_in09 = reg_0729;
    61: op1_01_in09 = reg_0458;
    62: op1_01_in09 = reg_0655;
    63: op1_01_in09 = imem05_in[107:104];
    64: op1_01_in09 = reg_0630;
    65: op1_01_in09 = reg_0710;
    66: op1_01_in09 = reg_0707;
    67: op1_01_in09 = reg_0719;
    69: op1_01_in09 = reg_1002;
    70: op1_01_in09 = reg_0145;
    85: op1_01_in09 = reg_0145;
    71: op1_01_in09 = reg_0680;
    72: op1_01_in09 = reg_0967;
    74: op1_01_in09 = reg_0157;
    75: op1_01_in09 = reg_0883;
    76: op1_01_in09 = reg_0837;
    77: op1_01_in09 = imem02_in[127:124];
    78: op1_01_in09 = imem05_in[7:4];
    79: op1_01_in09 = reg_0502;
    80: op1_01_in09 = reg_0722;
    81: op1_01_in09 = reg_0199;
    82: op1_01_in09 = reg_0453;
    83: op1_01_in09 = imem06_in[3:0];
    84: op1_01_in09 = imem04_in[79:76];
    86: op1_01_in09 = reg_0468;
    87: op1_01_in09 = reg_1010;
    88: op1_01_in09 = reg_0486;
    89: op1_01_in09 = reg_0475;
    90: op1_01_in09 = reg_0393;
    91: op1_01_in09 = imem07_in[87:84];
    93: op1_01_in09 = reg_0312;
    94: op1_01_in09 = reg_0631;
    95: op1_01_in09 = imem03_in[123:120];
    96: op1_01_in09 = reg_0894;
    97: op1_01_in09 = reg_0594;
    default: op1_01_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv09 = 1;
    6: op1_01_inv09 = 1;
    7: op1_01_inv09 = 1;
    8: op1_01_inv09 = 1;
    4: op1_01_inv09 = 1;
    12: op1_01_inv09 = 1;
    13: op1_01_inv09 = 1;
    15: op1_01_inv09 = 1;
    16: op1_01_inv09 = 1;
    18: op1_01_inv09 = 1;
    19: op1_01_inv09 = 1;
    23: op1_01_inv09 = 1;
    24: op1_01_inv09 = 1;
    28: op1_01_inv09 = 1;
    30: op1_01_inv09 = 1;
    31: op1_01_inv09 = 1;
    37: op1_01_inv09 = 1;
    38: op1_01_inv09 = 1;
    39: op1_01_inv09 = 1;
    40: op1_01_inv09 = 1;
    43: op1_01_inv09 = 1;
    44: op1_01_inv09 = 1;
    45: op1_01_inv09 = 1;
    47: op1_01_inv09 = 1;
    50: op1_01_inv09 = 1;
    52: op1_01_inv09 = 1;
    53: op1_01_inv09 = 1;
    56: op1_01_inv09 = 1;
    57: op1_01_inv09 = 1;
    58: op1_01_inv09 = 1;
    59: op1_01_inv09 = 1;
    60: op1_01_inv09 = 1;
    61: op1_01_inv09 = 1;
    66: op1_01_inv09 = 1;
    70: op1_01_inv09 = 1;
    72: op1_01_inv09 = 1;
    75: op1_01_inv09 = 1;
    76: op1_01_inv09 = 1;
    77: op1_01_inv09 = 1;
    83: op1_01_inv09 = 1;
    84: op1_01_inv09 = 1;
    89: op1_01_inv09 = 1;
    90: op1_01_inv09 = 1;
    default: op1_01_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in10 = reg_0219;
    6: op1_01_in10 = reg_0028;
    7: op1_01_in10 = reg_0335;
    8: op1_01_in10 = imem06_in[19:16];
    4: op1_01_in10 = reg_0444;
    9: op1_01_in10 = reg_0684;
    10: op1_01_in10 = imem03_in[23:20];
    11: op1_01_in10 = imem03_in[111:108];
    12: op1_01_in10 = reg_0453;
    13: op1_01_in10 = reg_0645;
    14: op1_01_in10 = imem07_in[75:72];
    15: op1_01_in10 = reg_0118;
    16: op1_01_in10 = reg_0355;
    17: op1_01_in10 = reg_0949;
    18: op1_01_in10 = reg_0678;
    19: op1_01_in10 = reg_0440;
    20: op1_01_in10 = reg_0455;
    21: op1_01_in10 = imem05_in[67:64];
    22: op1_01_in10 = reg_0450;
    82: op1_01_in10 = reg_0450;
    23: op1_01_in10 = reg_0329;
    24: op1_01_in10 = imem07_in[11:8];
    25: op1_01_in10 = reg_0343;
    26: op1_01_in10 = reg_0757;
    94: op1_01_in10 = reg_0757;
    27: op1_01_in10 = reg_0916;
    28: op1_01_in10 = reg_0489;
    29: op1_01_in10 = reg_0480;
    30: op1_01_in10 = imem02_in[95:92];
    31: op1_01_in10 = reg_0813;
    32: op1_01_in10 = reg_0464;
    35: op1_01_in10 = reg_0464;
    43: op1_01_in10 = reg_0464;
    33: op1_01_in10 = imem02_in[27:24];
    34: op1_01_in10 = reg_0318;
    37: op1_01_in10 = reg_0470;
    38: op1_01_in10 = reg_0641;
    73: op1_01_in10 = reg_0641;
    39: op1_01_in10 = reg_0114;
    40: op1_01_in10 = reg_1005;
    41: op1_01_in10 = reg_0369;
    42: op1_01_in10 = reg_1010;
    44: op1_01_in10 = imem02_in[55:52];
    45: op1_01_in10 = reg_0301;
    46: op1_01_in10 = reg_0720;
    47: op1_01_in10 = reg_0655;
    48: op1_01_in10 = reg_0346;
    49: op1_01_in10 = reg_0609;
    50: op1_01_in10 = reg_0175;
    51: op1_01_in10 = reg_0628;
    52: op1_01_in10 = reg_0050;
    53: op1_01_in10 = reg_0265;
    54: op1_01_in10 = reg_0969;
    55: op1_01_in10 = reg_0819;
    95: op1_01_in10 = reg_0819;
    56: op1_01_in10 = reg_0428;
    57: op1_01_in10 = reg_0828;
    58: op1_01_in10 = reg_0473;
    59: op1_01_in10 = reg_0718;
    60: op1_01_in10 = reg_0656;
    61: op1_01_in10 = reg_0194;
    62: op1_01_in10 = reg_0515;
    63: op1_01_in10 = imem05_in[123:120];
    64: op1_01_in10 = reg_0263;
    65: op1_01_in10 = reg_0703;
    66: op1_01_in10 = reg_0706;
    67: op1_01_in10 = reg_0717;
    69: op1_01_in10 = reg_0982;
    70: op1_01_in10 = reg_0135;
    71: op1_01_in10 = reg_0451;
    72: op1_01_in10 = reg_0528;
    75: op1_01_in10 = reg_0356;
    76: op1_01_in10 = reg_0441;
    77: op1_01_in10 = reg_0649;
    78: op1_01_in10 = imem05_in[31:28];
    79: op1_01_in10 = reg_0174;
    80: op1_01_in10 = reg_0165;
    81: op1_01_in10 = reg_0192;
    83: op1_01_in10 = imem06_in[39:36];
    84: op1_01_in10 = imem04_in[111:108];
    85: op1_01_in10 = imem06_in[87:84];
    86: op1_01_in10 = reg_0210;
    87: op1_01_in10 = reg_0403;
    88: op1_01_in10 = reg_0851;
    89: op1_01_in10 = reg_0460;
    90: op1_01_in10 = reg_0626;
    91: op1_01_in10 = reg_0726;
    93: op1_01_in10 = reg_0581;
    96: op1_01_in10 = reg_0493;
    97: op1_01_in10 = reg_0176;
    default: op1_01_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_01_inv10 = 1;
    7: op1_01_inv10 = 1;
    8: op1_01_inv10 = 1;
    10: op1_01_inv10 = 1;
    11: op1_01_inv10 = 1;
    12: op1_01_inv10 = 1;
    14: op1_01_inv10 = 1;
    15: op1_01_inv10 = 1;
    19: op1_01_inv10 = 1;
    24: op1_01_inv10 = 1;
    25: op1_01_inv10 = 1;
    28: op1_01_inv10 = 1;
    29: op1_01_inv10 = 1;
    30: op1_01_inv10 = 1;
    32: op1_01_inv10 = 1;
    33: op1_01_inv10 = 1;
    34: op1_01_inv10 = 1;
    37: op1_01_inv10 = 1;
    39: op1_01_inv10 = 1;
    41: op1_01_inv10 = 1;
    42: op1_01_inv10 = 1;
    43: op1_01_inv10 = 1;
    44: op1_01_inv10 = 1;
    45: op1_01_inv10 = 1;
    46: op1_01_inv10 = 1;
    49: op1_01_inv10 = 1;
    51: op1_01_inv10 = 1;
    56: op1_01_inv10 = 1;
    57: op1_01_inv10 = 1;
    61: op1_01_inv10 = 1;
    62: op1_01_inv10 = 1;
    63: op1_01_inv10 = 1;
    64: op1_01_inv10 = 1;
    65: op1_01_inv10 = 1;
    66: op1_01_inv10 = 1;
    69: op1_01_inv10 = 1;
    71: op1_01_inv10 = 1;
    75: op1_01_inv10 = 1;
    77: op1_01_inv10 = 1;
    79: op1_01_inv10 = 1;
    81: op1_01_inv10 = 1;
    82: op1_01_inv10 = 1;
    83: op1_01_inv10 = 1;
    84: op1_01_inv10 = 1;
    85: op1_01_inv10 = 1;
    86: op1_01_inv10 = 1;
    89: op1_01_inv10 = 1;
    90: op1_01_inv10 = 1;
    91: op1_01_inv10 = 1;
    93: op1_01_inv10 = 1;
    94: op1_01_inv10 = 1;
    96: op1_01_inv10 = 1;
    97: op1_01_inv10 = 1;
    default: op1_01_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in11 = reg_0118;
    6: op1_01_in11 = reg_0025;
    7: op1_01_in11 = reg_0336;
    8: op1_01_in11 = imem06_in[27:24];
    88: op1_01_in11 = imem06_in[27:24];
    4: op1_01_in11 = reg_0175;
    79: op1_01_in11 = reg_0175;
    9: op1_01_in11 = reg_0671;
    10: op1_01_in11 = imem03_in[39:36];
    11: op1_01_in11 = reg_0602;
    12: op1_01_in11 = reg_0454;
    13: op1_01_in11 = reg_0653;
    14: op1_01_in11 = imem07_in[123:120];
    15: op1_01_in11 = reg_0116;
    16: op1_01_in11 = reg_0052;
    17: op1_01_in11 = reg_0258;
    18: op1_01_in11 = reg_0669;
    19: op1_01_in11 = reg_0427;
    20: op1_01_in11 = reg_0457;
    21: op1_01_in11 = imem05_in[83:80];
    22: op1_01_in11 = reg_0464;
    23: op1_01_in11 = reg_0363;
    24: op1_01_in11 = imem07_in[35:32];
    25: op1_01_in11 = reg_0388;
    26: op1_01_in11 = reg_0229;
    27: op1_01_in11 = reg_0814;
    28: op1_01_in11 = reg_0497;
    29: op1_01_in11 = reg_0467;
    43: op1_01_in11 = reg_0467;
    30: op1_01_in11 = imem02_in[99:96];
    31: op1_01_in11 = reg_0831;
    32: op1_01_in11 = reg_0461;
    33: op1_01_in11 = imem02_in[75:72];
    44: op1_01_in11 = imem02_in[75:72];
    34: op1_01_in11 = reg_0339;
    35: op1_01_in11 = reg_0472;
    37: op1_01_in11 = reg_0468;
    38: op1_01_in11 = reg_0643;
    39: op1_01_in11 = imem02_in[3:0];
    40: op1_01_in11 = reg_0888;
    41: op1_01_in11 = reg_0992;
    42: op1_01_in11 = imem07_in[59:56];
    45: op1_01_in11 = reg_0306;
    46: op1_01_in11 = reg_0724;
    65: op1_01_in11 = reg_0724;
    47: op1_01_in11 = reg_0326;
    48: op1_01_in11 = reg_0847;
    49: op1_01_in11 = reg_0633;
    50: op1_01_in11 = reg_0180;
    51: op1_01_in11 = reg_0332;
    52: op1_01_in11 = reg_0909;
    53: op1_01_in11 = reg_1057;
    54: op1_01_in11 = reg_0964;
    55: op1_01_in11 = reg_0132;
    56: op1_01_in11 = reg_0641;
    57: op1_01_in11 = reg_0465;
    58: op1_01_in11 = reg_0191;
    59: op1_01_in11 = reg_0707;
    60: op1_01_in11 = reg_0651;
    61: op1_01_in11 = reg_0201;
    62: op1_01_in11 = reg_0365;
    63: op1_01_in11 = reg_0935;
    64: op1_01_in11 = imem07_in[11:8];
    66: op1_01_in11 = reg_0406;
    67: op1_01_in11 = reg_0702;
    69: op1_01_in11 = reg_0984;
    70: op1_01_in11 = reg_0133;
    71: op1_01_in11 = reg_0455;
    72: op1_01_in11 = reg_0343;
    73: op1_01_in11 = reg_0166;
    75: op1_01_in11 = reg_0828;
    76: op1_01_in11 = reg_0039;
    77: op1_01_in11 = reg_0763;
    78: op1_01_in11 = imem05_in[35:32];
    80: op1_01_in11 = reg_0159;
    81: op1_01_in11 = imem01_in[11:8];
    82: op1_01_in11 = reg_0462;
    83: op1_01_in11 = imem06_in[67:64];
    84: op1_01_in11 = reg_0446;
    85: op1_01_in11 = imem06_in[107:104];
    86: op1_01_in11 = reg_0195;
    87: op1_01_in11 = reg_0782;
    89: op1_01_in11 = reg_0479;
    90: op1_01_in11 = reg_0754;
    91: op1_01_in11 = reg_0560;
    93: op1_01_in11 = reg_0588;
    94: op1_01_in11 = reg_0049;
    95: op1_01_in11 = reg_1050;
    96: op1_01_in11 = imem03_in[31:28];
    97: op1_01_in11 = reg_0877;
    default: op1_01_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv11 = 1;
    4: op1_01_inv11 = 1;
    10: op1_01_inv11 = 1;
    13: op1_01_inv11 = 1;
    14: op1_01_inv11 = 1;
    16: op1_01_inv11 = 1;
    17: op1_01_inv11 = 1;
    18: op1_01_inv11 = 1;
    19: op1_01_inv11 = 1;
    22: op1_01_inv11 = 1;
    23: op1_01_inv11 = 1;
    26: op1_01_inv11 = 1;
    27: op1_01_inv11 = 1;
    28: op1_01_inv11 = 1;
    29: op1_01_inv11 = 1;
    30: op1_01_inv11 = 1;
    31: op1_01_inv11 = 1;
    32: op1_01_inv11 = 1;
    34: op1_01_inv11 = 1;
    37: op1_01_inv11 = 1;
    39: op1_01_inv11 = 1;
    40: op1_01_inv11 = 1;
    41: op1_01_inv11 = 1;
    44: op1_01_inv11 = 1;
    49: op1_01_inv11 = 1;
    55: op1_01_inv11 = 1;
    58: op1_01_inv11 = 1;
    59: op1_01_inv11 = 1;
    60: op1_01_inv11 = 1;
    61: op1_01_inv11 = 1;
    65: op1_01_inv11 = 1;
    67: op1_01_inv11 = 1;
    69: op1_01_inv11 = 1;
    70: op1_01_inv11 = 1;
    72: op1_01_inv11 = 1;
    75: op1_01_inv11 = 1;
    77: op1_01_inv11 = 1;
    78: op1_01_inv11 = 1;
    79: op1_01_inv11 = 1;
    82: op1_01_inv11 = 1;
    87: op1_01_inv11 = 1;
    91: op1_01_inv11 = 1;
    default: op1_01_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in12 = reg_0104;
    15: op1_01_in12 = reg_0104;
    6: op1_01_in12 = imem07_in[47:44];
    24: op1_01_in12 = imem07_in[47:44];
    7: op1_01_in12 = reg_0089;
    8: op1_01_in12 = imem06_in[91:88];
    4: op1_01_in12 = reg_0180;
    9: op1_01_in12 = reg_0688;
    10: op1_01_in12 = imem03_in[47:44];
    11: op1_01_in12 = reg_0582;
    12: op1_01_in12 = reg_0469;
    22: op1_01_in12 = reg_0469;
    13: op1_01_in12 = reg_0637;
    14: op1_01_in12 = imem07_in[127:124];
    16: op1_01_in12 = reg_0086;
    17: op1_01_in12 = reg_0254;
    18: op1_01_in12 = reg_0481;
    82: op1_01_in12 = reg_0481;
    19: op1_01_in12 = reg_0181;
    50: op1_01_in12 = reg_0181;
    20: op1_01_in12 = reg_0464;
    21: op1_01_in12 = reg_0963;
    23: op1_01_in12 = reg_0338;
    25: op1_01_in12 = reg_0362;
    26: op1_01_in12 = reg_0816;
    27: op1_01_in12 = reg_0091;
    28: op1_01_in12 = reg_0134;
    29: op1_01_in12 = reg_0200;
    30: op1_01_in12 = imem02_in[103:100];
    31: op1_01_in12 = reg_0156;
    32: op1_01_in12 = reg_0466;
    33: op1_01_in12 = reg_0645;
    34: op1_01_in12 = reg_0082;
    35: op1_01_in12 = reg_0479;
    37: op1_01_in12 = reg_0459;
    38: op1_01_in12 = reg_0659;
    39: op1_01_in12 = imem02_in[31:28];
    40: op1_01_in12 = reg_0778;
    41: op1_01_in12 = reg_0984;
    42: op1_01_in12 = imem07_in[83:80];
    43: op1_01_in12 = reg_0214;
    44: op1_01_in12 = imem02_in[91:88];
    45: op1_01_in12 = reg_0539;
    46: op1_01_in12 = reg_0715;
    47: op1_01_in12 = reg_0341;
    48: op1_01_in12 = reg_0874;
    49: op1_01_in12 = imem07_in[11:8];
    51: op1_01_in12 = reg_0625;
    52: op1_01_in12 = reg_0076;
    53: op1_01_in12 = reg_0292;
    54: op1_01_in12 = reg_0952;
    55: op1_01_in12 = reg_0149;
    56: op1_01_in12 = reg_0838;
    57: op1_01_in12 = reg_0476;
    58: op1_01_in12 = reg_0204;
    59: op1_01_in12 = reg_0700;
    60: op1_01_in12 = reg_0052;
    61: op1_01_in12 = reg_0205;
    62: op1_01_in12 = reg_0652;
    63: op1_01_in12 = reg_0956;
    64: op1_01_in12 = imem07_in[31:28];
    65: op1_01_in12 = reg_0729;
    66: op1_01_in12 = reg_0599;
    67: op1_01_in12 = reg_0712;
    69: op1_01_in12 = reg_0974;
    70: op1_01_in12 = reg_0152;
    71: op1_01_in12 = reg_0461;
    72: op1_01_in12 = reg_0940;
    75: op1_01_in12 = reg_0687;
    76: op1_01_in12 = reg_0347;
    77: op1_01_in12 = reg_0643;
    78: op1_01_in12 = imem05_in[47:44];
    79: op1_01_in12 = reg_0172;
    80: op1_01_in12 = reg_0717;
    81: op1_01_in12 = imem01_in[23:20];
    83: op1_01_in12 = imem06_in[75:72];
    84: op1_01_in12 = reg_0395;
    85: op1_01_in12 = imem06_in[119:116];
    86: op1_01_in12 = reg_0206;
    87: op1_01_in12 = reg_0369;
    88: op1_01_in12 = imem06_in[59:56];
    89: op1_01_in12 = reg_0452;
    90: op1_01_in12 = reg_0614;
    91: op1_01_in12 = reg_0563;
    93: op1_01_in12 = reg_0551;
    94: op1_01_in12 = reg_0301;
    95: op1_01_in12 = reg_0357;
    96: op1_01_in12 = imem03_in[91:88];
    97: op1_01_in12 = reg_0740;
    default: op1_01_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv12 = 1;
    7: op1_01_inv12 = 1;
    8: op1_01_inv12 = 1;
    4: op1_01_inv12 = 1;
    10: op1_01_inv12 = 1;
    12: op1_01_inv12 = 1;
    15: op1_01_inv12 = 1;
    17: op1_01_inv12 = 1;
    18: op1_01_inv12 = 1;
    19: op1_01_inv12 = 1;
    21: op1_01_inv12 = 1;
    23: op1_01_inv12 = 1;
    26: op1_01_inv12 = 1;
    27: op1_01_inv12 = 1;
    28: op1_01_inv12 = 1;
    29: op1_01_inv12 = 1;
    30: op1_01_inv12 = 1;
    31: op1_01_inv12 = 1;
    35: op1_01_inv12 = 1;
    40: op1_01_inv12 = 1;
    41: op1_01_inv12 = 1;
    43: op1_01_inv12 = 1;
    46: op1_01_inv12 = 1;
    47: op1_01_inv12 = 1;
    48: op1_01_inv12 = 1;
    50: op1_01_inv12 = 1;
    51: op1_01_inv12 = 1;
    55: op1_01_inv12 = 1;
    56: op1_01_inv12 = 1;
    58: op1_01_inv12 = 1;
    60: op1_01_inv12 = 1;
    61: op1_01_inv12 = 1;
    62: op1_01_inv12 = 1;
    65: op1_01_inv12 = 1;
    66: op1_01_inv12 = 1;
    70: op1_01_inv12 = 1;
    72: op1_01_inv12 = 1;
    75: op1_01_inv12 = 1;
    77: op1_01_inv12 = 1;
    78: op1_01_inv12 = 1;
    83: op1_01_inv12 = 1;
    85: op1_01_inv12 = 1;
    88: op1_01_inv12 = 1;
    93: op1_01_inv12 = 1;
    95: op1_01_inv12 = 1;
    96: op1_01_inv12 = 1;
    97: op1_01_inv12 = 1;
    default: op1_01_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in13 = reg_0100;
    6: op1_01_in13 = imem07_in[123:120];
    7: op1_01_in13 = reg_0096;
    8: op1_01_in13 = imem06_in[95:92];
    4: op1_01_in13 = reg_0162;
    50: op1_01_in13 = reg_0162;
    9: op1_01_in13 = reg_0462;
    10: op1_01_in13 = imem03_in[51:48];
    11: op1_01_in13 = reg_0572;
    12: op1_01_in13 = reg_0472;
    13: op1_01_in13 = reg_0651;
    14: op1_01_in13 = reg_0729;
    15: op1_01_in13 = reg_0119;
    16: op1_01_in13 = reg_0055;
    17: op1_01_in13 = reg_0132;
    18: op1_01_in13 = reg_0473;
    19: op1_01_in13 = reg_0179;
    20: op1_01_in13 = reg_0469;
    21: op1_01_in13 = reg_0959;
    22: op1_01_in13 = reg_0467;
    23: op1_01_in13 = reg_0355;
    24: op1_01_in13 = imem07_in[55:52];
    25: op1_01_in13 = reg_0369;
    26: op1_01_in13 = reg_0275;
    27: op1_01_in13 = reg_0872;
    28: op1_01_in13 = imem06_in[63:60];
    29: op1_01_in13 = reg_0203;
    30: op1_01_in13 = imem02_in[111:108];
    31: op1_01_in13 = reg_0139;
    32: op1_01_in13 = reg_0480;
    82: op1_01_in13 = reg_0480;
    33: op1_01_in13 = reg_0658;
    34: op1_01_in13 = reg_0817;
    35: op1_01_in13 = reg_0452;
    37: op1_01_in13 = reg_0200;
    38: op1_01_in13 = reg_0837;
    62: op1_01_in13 = reg_0837;
    39: op1_01_in13 = imem02_in[39:36];
    40: op1_01_in13 = reg_0050;
    41: op1_01_in13 = reg_0989;
    42: op1_01_in13 = reg_0713;
    65: op1_01_in13 = reg_0713;
    43: op1_01_in13 = reg_0208;
    44: op1_01_in13 = imem02_in[95:92];
    45: op1_01_in13 = reg_0524;
    46: op1_01_in13 = reg_0707;
    47: op1_01_in13 = reg_0515;
    48: op1_01_in13 = reg_0543;
    49: op1_01_in13 = imem07_in[51:48];
    51: op1_01_in13 = reg_0894;
    52: op1_01_in13 = reg_0276;
    53: op1_01_in13 = reg_0540;
    54: op1_01_in13 = reg_0233;
    55: op1_01_in13 = reg_0142;
    56: op1_01_in13 = reg_0180;
    57: op1_01_in13 = reg_0466;
    58: op1_01_in13 = reg_0211;
    59: op1_01_in13 = reg_0361;
    60: op1_01_in13 = reg_0423;
    61: op1_01_in13 = reg_0202;
    63: op1_01_in13 = reg_0491;
    64: op1_01_in13 = imem07_in[47:44];
    66: op1_01_in13 = reg_0502;
    67: op1_01_in13 = reg_0709;
    69: op1_01_in13 = reg_0994;
    70: op1_01_in13 = reg_0153;
    71: op1_01_in13 = reg_0477;
    72: op1_01_in13 = reg_0125;
    75: op1_01_in13 = reg_0749;
    76: op1_01_in13 = reg_0088;
    77: op1_01_in13 = reg_0358;
    78: op1_01_in13 = imem05_in[63:60];
    79: op1_01_in13 = reg_0171;
    80: op1_01_in13 = reg_0374;
    81: op1_01_in13 = imem01_in[51:48];
    83: op1_01_in13 = imem06_in[83:80];
    84: op1_01_in13 = reg_0550;
    85: op1_01_in13 = imem06_in[127:124];
    86: op1_01_in13 = imem01_in[3:0];
    87: op1_01_in13 = reg_0573;
    88: op1_01_in13 = imem06_in[99:96];
    89: op1_01_in13 = reg_0189;
    90: op1_01_in13 = reg_0439;
    91: op1_01_in13 = reg_0653;
    93: op1_01_in13 = reg_0373;
    94: op1_01_in13 = reg_0763;
    95: op1_01_in13 = reg_0558;
    96: op1_01_in13 = reg_0785;
    97: op1_01_in13 = reg_0845;
    default: op1_01_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_01_inv13 = 1;
    11: op1_01_inv13 = 1;
    13: op1_01_inv13 = 1;
    15: op1_01_inv13 = 1;
    16: op1_01_inv13 = 1;
    17: op1_01_inv13 = 1;
    18: op1_01_inv13 = 1;
    20: op1_01_inv13 = 1;
    21: op1_01_inv13 = 1;
    23: op1_01_inv13 = 1;
    24: op1_01_inv13 = 1;
    26: op1_01_inv13 = 1;
    27: op1_01_inv13 = 1;
    28: op1_01_inv13 = 1;
    29: op1_01_inv13 = 1;
    32: op1_01_inv13 = 1;
    33: op1_01_inv13 = 1;
    34: op1_01_inv13 = 1;
    35: op1_01_inv13 = 1;
    37: op1_01_inv13 = 1;
    38: op1_01_inv13 = 1;
    39: op1_01_inv13 = 1;
    40: op1_01_inv13 = 1;
    42: op1_01_inv13 = 1;
    43: op1_01_inv13 = 1;
    44: op1_01_inv13 = 1;
    50: op1_01_inv13 = 1;
    51: op1_01_inv13 = 1;
    53: op1_01_inv13 = 1;
    54: op1_01_inv13 = 1;
    59: op1_01_inv13 = 1;
    60: op1_01_inv13 = 1;
    63: op1_01_inv13 = 1;
    64: op1_01_inv13 = 1;
    65: op1_01_inv13 = 1;
    66: op1_01_inv13 = 1;
    67: op1_01_inv13 = 1;
    72: op1_01_inv13 = 1;
    76: op1_01_inv13 = 1;
    82: op1_01_inv13 = 1;
    84: op1_01_inv13 = 1;
    85: op1_01_inv13 = 1;
    91: op1_01_inv13 = 1;
    93: op1_01_inv13 = 1;
    94: op1_01_inv13 = 1;
    95: op1_01_inv13 = 1;
    96: op1_01_inv13 = 1;
    97: op1_01_inv13 = 1;
    default: op1_01_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in14 = reg_0109;
    6: op1_01_in14 = reg_0717;
    7: op1_01_in14 = reg_0082;
    8: op1_01_in14 = reg_0614;
    4: op1_01_in14 = reg_0169;
    9: op1_01_in14 = reg_0206;
    61: op1_01_in14 = reg_0206;
    10: op1_01_in14 = imem03_in[71:68];
    11: op1_01_in14 = reg_0587;
    12: op1_01_in14 = reg_0473;
    13: op1_01_in14 = reg_0662;
    14: op1_01_in14 = reg_0706;
    46: op1_01_in14 = reg_0706;
    15: op1_01_in14 = reg_0115;
    16: op1_01_in14 = reg_0060;
    17: op1_01_in14 = reg_0148;
    18: op1_01_in14 = reg_0456;
    82: op1_01_in14 = reg_0456;
    19: op1_01_in14 = reg_0167;
    50: op1_01_in14 = reg_0167;
    20: op1_01_in14 = reg_0466;
    21: op1_01_in14 = reg_0957;
    22: op1_01_in14 = reg_0468;
    23: op1_01_in14 = reg_0336;
    24: op1_01_in14 = imem07_in[63:60];
    25: op1_01_in14 = reg_0393;
    26: op1_01_in14 = reg_0832;
    27: op1_01_in14 = imem03_in[43:40];
    28: op1_01_in14 = imem06_in[95:92];
    29: op1_01_in14 = reg_0193;
    43: op1_01_in14 = reg_0193;
    30: op1_01_in14 = imem02_in[123:120];
    31: op1_01_in14 = reg_0138;
    32: op1_01_in14 = reg_0470;
    75: op1_01_in14 = reg_0470;
    33: op1_01_in14 = reg_0653;
    34: op1_01_in14 = reg_0762;
    35: op1_01_in14 = reg_0478;
    37: op1_01_in14 = reg_0187;
    38: op1_01_in14 = reg_0334;
    39: op1_01_in14 = imem02_in[47:44];
    40: op1_01_in14 = reg_0764;
    41: op1_01_in14 = reg_0974;
    42: op1_01_in14 = reg_0436;
    44: op1_01_in14 = reg_0664;
    45: op1_01_in14 = reg_0068;
    47: op1_01_in14 = reg_0026;
    48: op1_01_in14 = reg_0038;
    49: op1_01_in14 = imem07_in[95:92];
    51: op1_01_in14 = reg_0780;
    52: op1_01_in14 = reg_0284;
    53: op1_01_in14 = reg_0537;
    54: op1_01_in14 = reg_0826;
    55: op1_01_in14 = imem06_in[7:4];
    56: op1_01_in14 = reg_0159;
    57: op1_01_in14 = reg_0480;
    58: op1_01_in14 = reg_0205;
    59: op1_01_in14 = reg_0641;
    60: op1_01_in14 = reg_0818;
    62: op1_01_in14 = reg_0358;
    63: op1_01_in14 = reg_0945;
    64: op1_01_in14 = imem07_in[51:48];
    65: op1_01_in14 = reg_0701;
    66: op1_01_in14 = reg_0175;
    67: op1_01_in14 = reg_0705;
    69: op1_01_in14 = imem04_in[7:4];
    70: op1_01_in14 = reg_0137;
    71: op1_01_in14 = reg_0474;
    72: op1_01_in14 = reg_0865;
    76: op1_01_in14 = reg_0867;
    77: op1_01_in14 = reg_0368;
    78: op1_01_in14 = imem05_in[87:84];
    79: op1_01_in14 = reg_0184;
    80: op1_01_in14 = reg_0959;
    81: op1_01_in14 = imem01_in[83:80];
    83: op1_01_in14 = reg_0660;
    84: op1_01_in14 = reg_0937;
    85: op1_01_in14 = reg_0735;
    86: op1_01_in14 = imem01_in[23:20];
    87: op1_01_in14 = imem07_in[3:0];
    88: op1_01_in14 = reg_0696;
    89: op1_01_in14 = reg_0188;
    90: op1_01_in14 = reg_0382;
    91: op1_01_in14 = reg_0727;
    93: op1_01_in14 = reg_0242;
    94: op1_01_in14 = reg_0623;
    95: op1_01_in14 = reg_0596;
    96: op1_01_in14 = reg_0357;
    97: op1_01_in14 = reg_0925;
    default: op1_01_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_01_inv14 = 1;
    4: op1_01_inv14 = 1;
    11: op1_01_inv14 = 1;
    12: op1_01_inv14 = 1;
    16: op1_01_inv14 = 1;
    18: op1_01_inv14 = 1;
    20: op1_01_inv14 = 1;
    21: op1_01_inv14 = 1;
    22: op1_01_inv14 = 1;
    23: op1_01_inv14 = 1;
    27: op1_01_inv14 = 1;
    29: op1_01_inv14 = 1;
    30: op1_01_inv14 = 1;
    32: op1_01_inv14 = 1;
    35: op1_01_inv14 = 1;
    37: op1_01_inv14 = 1;
    45: op1_01_inv14 = 1;
    48: op1_01_inv14 = 1;
    53: op1_01_inv14 = 1;
    54: op1_01_inv14 = 1;
    56: op1_01_inv14 = 1;
    58: op1_01_inv14 = 1;
    63: op1_01_inv14 = 1;
    65: op1_01_inv14 = 1;
    67: op1_01_inv14 = 1;
    71: op1_01_inv14 = 1;
    72: op1_01_inv14 = 1;
    81: op1_01_inv14 = 1;
    84: op1_01_inv14 = 1;
    88: op1_01_inv14 = 1;
    89: op1_01_inv14 = 1;
    94: op1_01_inv14 = 1;
    default: op1_01_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in15 = imem02_in[23:20];
    6: op1_01_in15 = reg_0725;
    7: op1_01_in15 = reg_0091;
    8: op1_01_in15 = reg_0607;
    4: op1_01_in15 = reg_0177;
    9: op1_01_in15 = reg_0199;
    58: op1_01_in15 = reg_0199;
    10: op1_01_in15 = imem03_in[83:80];
    11: op1_01_in15 = reg_0600;
    12: op1_01_in15 = reg_0452;
    13: op1_01_in15 = reg_0644;
    14: op1_01_in15 = reg_0432;
    15: op1_01_in15 = reg_0110;
    16: op1_01_in15 = reg_0094;
    17: op1_01_in15 = reg_0135;
    18: op1_01_in15 = reg_0188;
    82: op1_01_in15 = reg_0188;
    20: op1_01_in15 = reg_0467;
    21: op1_01_in15 = reg_0969;
    22: op1_01_in15 = reg_0459;
    23: op1_01_in15 = reg_0083;
    24: op1_01_in15 = imem07_in[75:72];
    25: op1_01_in15 = reg_0396;
    26: op1_01_in15 = reg_0819;
    27: op1_01_in15 = imem03_in[47:44];
    28: op1_01_in15 = imem06_in[107:104];
    29: op1_01_in15 = reg_0194;
    35: op1_01_in15 = reg_0194;
    30: op1_01_in15 = reg_0666;
    31: op1_01_in15 = reg_0140;
    32: op1_01_in15 = reg_0456;
    33: op1_01_in15 = reg_0639;
    34: op1_01_in15 = reg_0336;
    37: op1_01_in15 = reg_0211;
    38: op1_01_in15 = reg_0916;
    39: op1_01_in15 = imem02_in[59:56];
    40: op1_01_in15 = reg_0760;
    41: op1_01_in15 = reg_0990;
    42: op1_01_in15 = reg_0445;
    43: op1_01_in15 = reg_0207;
    89: op1_01_in15 = reg_0207;
    44: op1_01_in15 = reg_0659;
    45: op1_01_in15 = reg_0732;
    46: op1_01_in15 = reg_0700;
    47: op1_01_in15 = reg_0637;
    48: op1_01_in15 = reg_0377;
    49: op1_01_in15 = reg_0722;
    50: op1_01_in15 = reg_0163;
    51: op1_01_in15 = reg_0609;
    52: op1_01_in15 = reg_0893;
    53: op1_01_in15 = reg_0802;
    54: op1_01_in15 = reg_0259;
    55: op1_01_in15 = imem06_in[15:12];
    56: op1_01_in15 = reg_0183;
    57: op1_01_in15 = reg_0471;
    59: op1_01_in15 = reg_0350;
    60: op1_01_in15 = reg_0037;
    61: op1_01_in15 = imem01_in[7:4];
    62: op1_01_in15 = reg_0664;
    63: op1_01_in15 = reg_0254;
    64: op1_01_in15 = imem07_in[63:60];
    65: op1_01_in15 = reg_0002;
    66: op1_01_in15 = reg_0181;
    67: op1_01_in15 = reg_0325;
    69: op1_01_in15 = imem04_in[15:12];
    70: op1_01_in15 = imem06_in[19:16];
    71: op1_01_in15 = reg_0214;
    72: op1_01_in15 = reg_0947;
    75: op1_01_in15 = reg_0209;
    76: op1_01_in15 = reg_0090;
    77: op1_01_in15 = reg_0372;
    78: op1_01_in15 = imem05_in[111:108];
    80: op1_01_in15 = reg_0903;
    81: op1_01_in15 = imem01_in[107:104];
    83: op1_01_in15 = reg_0694;
    84: op1_01_in15 = reg_1009;
    85: op1_01_in15 = reg_0591;
    86: op1_01_in15 = imem01_in[87:84];
    87: op1_01_in15 = imem07_in[35:32];
    88: op1_01_in15 = reg_0267;
    90: op1_01_in15 = reg_0380;
    91: op1_01_in15 = reg_0744;
    93: op1_01_in15 = reg_0979;
    94: op1_01_in15 = reg_0596;
    95: op1_01_in15 = reg_0281;
    96: op1_01_in15 = reg_0558;
    97: op1_01_in15 = reg_0827;
    default: op1_01_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_01_inv15 = 1;
    4: op1_01_inv15 = 1;
    9: op1_01_inv15 = 1;
    11: op1_01_inv15 = 1;
    13: op1_01_inv15 = 1;
    15: op1_01_inv15 = 1;
    16: op1_01_inv15 = 1;
    17: op1_01_inv15 = 1;
    23: op1_01_inv15 = 1;
    24: op1_01_inv15 = 1;
    25: op1_01_inv15 = 1;
    27: op1_01_inv15 = 1;
    28: op1_01_inv15 = 1;
    30: op1_01_inv15 = 1;
    33: op1_01_inv15 = 1;
    34: op1_01_inv15 = 1;
    35: op1_01_inv15 = 1;
    37: op1_01_inv15 = 1;
    38: op1_01_inv15 = 1;
    39: op1_01_inv15 = 1;
    40: op1_01_inv15 = 1;
    41: op1_01_inv15 = 1;
    43: op1_01_inv15 = 1;
    44: op1_01_inv15 = 1;
    46: op1_01_inv15 = 1;
    53: op1_01_inv15 = 1;
    54: op1_01_inv15 = 1;
    55: op1_01_inv15 = 1;
    57: op1_01_inv15 = 1;
    59: op1_01_inv15 = 1;
    61: op1_01_inv15 = 1;
    62: op1_01_inv15 = 1;
    67: op1_01_inv15 = 1;
    72: op1_01_inv15 = 1;
    76: op1_01_inv15 = 1;
    81: op1_01_inv15 = 1;
    82: op1_01_inv15 = 1;
    83: op1_01_inv15 = 1;
    84: op1_01_inv15 = 1;
    85: op1_01_inv15 = 1;
    86: op1_01_inv15 = 1;
    90: op1_01_inv15 = 1;
    91: op1_01_inv15 = 1;
    93: op1_01_inv15 = 1;
    95: op1_01_inv15 = 1;
    97: op1_01_inv15 = 1;
    default: op1_01_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in16 = imem02_in[43:40];
    6: op1_01_in16 = reg_0701;
    7: op1_01_in16 = reg_0094;
    8: op1_01_in16 = reg_0608;
    4: op1_01_in16 = reg_0170;
    9: op1_01_in16 = imem01_in[23:20];
    61: op1_01_in16 = imem01_in[23:20];
    10: op1_01_in16 = imem03_in[87:84];
    11: op1_01_in16 = reg_0578;
    12: op1_01_in16 = reg_0478;
    22: op1_01_in16 = reg_0478;
    13: op1_01_in16 = reg_0643;
    14: op1_01_in16 = reg_0426;
    15: op1_01_in16 = imem02_in[31:28];
    16: op1_01_in16 = imem03_in[7:4];
    17: op1_01_in16 = reg_0143;
    18: op1_01_in16 = reg_0198;
    20: op1_01_in16 = reg_0471;
    21: op1_01_in16 = reg_0943;
    23: op1_01_in16 = reg_0758;
    34: op1_01_in16 = reg_0758;
    24: op1_01_in16 = imem07_in[91:88];
    25: op1_01_in16 = reg_0374;
    26: op1_01_in16 = reg_0149;
    27: op1_01_in16 = imem03_in[67:64];
    28: op1_01_in16 = imem06_in[123:120];
    29: op1_01_in16 = imem01_in[15:12];
    30: op1_01_in16 = reg_0646;
    31: op1_01_in16 = reg_0155;
    32: op1_01_in16 = reg_0187;
    71: op1_01_in16 = reg_0187;
    33: op1_01_in16 = reg_0662;
    35: op1_01_in16 = reg_0199;
    37: op1_01_in16 = reg_0194;
    38: op1_01_in16 = reg_0330;
    39: op1_01_in16 = imem02_in[83:80];
    40: op1_01_in16 = reg_0066;
    41: op1_01_in16 = reg_0976;
    42: op1_01_in16 = reg_0439;
    43: op1_01_in16 = reg_0211;
    44: op1_01_in16 = reg_0667;
    45: op1_01_in16 = reg_0748;
    46: op1_01_in16 = reg_0805;
    47: op1_01_in16 = reg_0916;
    48: op1_01_in16 = reg_0807;
    49: op1_01_in16 = reg_0728;
    50: op1_01_in16 = reg_0168;
    51: op1_01_in16 = reg_0626;
    52: op1_01_in16 = reg_0059;
    53: op1_01_in16 = reg_0302;
    54: op1_01_in16 = reg_0508;
    55: op1_01_in16 = imem06_in[35:32];
    56: op1_01_in16 = reg_0166;
    57: op1_01_in16 = reg_0479;
    58: op1_01_in16 = imem01_in[3:0];
    59: op1_01_in16 = reg_0589;
    60: op1_01_in16 = reg_0083;
    62: op1_01_in16 = reg_0052;
    63: op1_01_in16 = reg_0972;
    64: op1_01_in16 = imem07_in[67:64];
    65: op1_01_in16 = reg_0321;
    66: op1_01_in16 = reg_0164;
    67: op1_01_in16 = reg_0422;
    69: op1_01_in16 = imem04_in[47:44];
    70: op1_01_in16 = imem06_in[23:20];
    72: op1_01_in16 = reg_0145;
    75: op1_01_in16 = reg_0193;
    76: op1_01_in16 = imem03_in[31:28];
    77: op1_01_in16 = reg_0331;
    78: op1_01_in16 = imem05_in[119:116];
    80: op1_01_in16 = reg_0575;
    81: op1_01_in16 = reg_0106;
    82: op1_01_in16 = reg_0207;
    83: op1_01_in16 = reg_0691;
    84: op1_01_in16 = reg_0870;
    85: op1_01_in16 = reg_0293;
    86: op1_01_in16 = imem01_in[91:88];
    87: op1_01_in16 = imem07_in[39:36];
    88: op1_01_in16 = reg_0262;
    89: op1_01_in16 = imem01_in[39:36];
    90: op1_01_in16 = reg_0918;
    91: op1_01_in16 = reg_0428;
    93: op1_01_in16 = reg_0290;
    94: op1_01_in16 = reg_0773;
    95: op1_01_in16 = reg_1049;
    96: op1_01_in16 = reg_0581;
    97: op1_01_in16 = reg_0117;
    default: op1_01_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv16 = 1;
    6: op1_01_inv16 = 1;
    8: op1_01_inv16 = 1;
    9: op1_01_inv16 = 1;
    11: op1_01_inv16 = 1;
    13: op1_01_inv16 = 1;
    14: op1_01_inv16 = 1;
    16: op1_01_inv16 = 1;
    23: op1_01_inv16 = 1;
    24: op1_01_inv16 = 1;
    26: op1_01_inv16 = 1;
    30: op1_01_inv16 = 1;
    31: op1_01_inv16 = 1;
    33: op1_01_inv16 = 1;
    34: op1_01_inv16 = 1;
    38: op1_01_inv16 = 1;
    39: op1_01_inv16 = 1;
    41: op1_01_inv16 = 1;
    42: op1_01_inv16 = 1;
    43: op1_01_inv16 = 1;
    45: op1_01_inv16 = 1;
    46: op1_01_inv16 = 1;
    47: op1_01_inv16 = 1;
    49: op1_01_inv16 = 1;
    51: op1_01_inv16 = 1;
    52: op1_01_inv16 = 1;
    54: op1_01_inv16 = 1;
    56: op1_01_inv16 = 1;
    57: op1_01_inv16 = 1;
    58: op1_01_inv16 = 1;
    66: op1_01_inv16 = 1;
    67: op1_01_inv16 = 1;
    77: op1_01_inv16 = 1;
    81: op1_01_inv16 = 1;
    83: op1_01_inv16 = 1;
    85: op1_01_inv16 = 1;
    86: op1_01_inv16 = 1;
    88: op1_01_inv16 = 1;
    89: op1_01_inv16 = 1;
    90: op1_01_inv16 = 1;
    91: op1_01_inv16 = 1;
    93: op1_01_inv16 = 1;
    96: op1_01_inv16 = 1;
    default: op1_01_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in17 = imem02_in[71:68];
    6: op1_01_in17 = reg_0436;
    7: op1_01_in17 = reg_0073;
    8: op1_01_in17 = reg_0618;
    9: op1_01_in17 = imem01_in[43:40];
    10: op1_01_in17 = imem03_in[123:120];
    11: op1_01_in17 = reg_0597;
    12: op1_01_in17 = reg_0210;
    13: op1_01_in17 = reg_0665;
    14: op1_01_in17 = reg_0175;
    15: op1_01_in17 = imem02_in[39:36];
    16: op1_01_in17 = imem03_in[79:76];
    17: op1_01_in17 = reg_0130;
    18: op1_01_in17 = reg_0196;
    20: op1_01_in17 = reg_0459;
    21: op1_01_in17 = reg_0826;
    22: op1_01_in17 = imem01_in[31:28];
    23: op1_01_in17 = reg_0761;
    24: op1_01_in17 = imem07_in[99:96];
    25: op1_01_in17 = reg_0982;
    26: op1_01_in17 = reg_0150;
    27: op1_01_in17 = imem03_in[119:116];
    28: op1_01_in17 = imem06_in[127:124];
    29: op1_01_in17 = imem01_in[99:96];
    30: op1_01_in17 = reg_0647;
    31: op1_01_in17 = imem06_in[7:4];
    72: op1_01_in17 = imem06_in[7:4];
    32: op1_01_in17 = reg_0209;
    33: op1_01_in17 = reg_0863;
    34: op1_01_in17 = reg_0506;
    35: op1_01_in17 = imem01_in[15:12];
    58: op1_01_in17 = imem01_in[15:12];
    37: op1_01_in17 = reg_0198;
    38: op1_01_in17 = reg_0817;
    39: op1_01_in17 = reg_0660;
    40: op1_01_in17 = reg_0009;
    41: op1_01_in17 = imem04_in[35:32];
    42: op1_01_in17 = reg_0446;
    43: op1_01_in17 = reg_0213;
    44: op1_01_in17 = reg_0842;
    45: op1_01_in17 = reg_0044;
    46: op1_01_in17 = reg_0422;
    47: op1_01_in17 = reg_0096;
    48: op1_01_in17 = reg_0513;
    49: op1_01_in17 = reg_0704;
    50: op1_01_in17 = reg_0170;
    51: op1_01_in17 = reg_0029;
    52: op1_01_in17 = reg_0281;
    53: op1_01_in17 = reg_0015;
    54: op1_01_in17 = reg_0757;
    55: op1_01_in17 = imem06_in[59:56];
    56: op1_01_in17 = reg_0158;
    57: op1_01_in17 = reg_0214;
    59: op1_01_in17 = reg_0162;
    60: op1_01_in17 = imem03_in[11:8];
    61: op1_01_in17 = imem01_in[87:84];
    62: op1_01_in17 = reg_0425;
    63: op1_01_in17 = reg_0019;
    64: op1_01_in17 = imem07_in[91:88];
    65: op1_01_in17 = reg_0641;
    66: op1_01_in17 = reg_0168;
    67: op1_01_in17 = reg_0502;
    69: op1_01_in17 = imem04_in[51:48];
    70: op1_01_in17 = imem06_in[39:36];
    71: op1_01_in17 = reg_0203;
    75: op1_01_in17 = reg_0190;
    76: op1_01_in17 = imem03_in[103:100];
    77: op1_01_in17 = reg_0083;
    78: op1_01_in17 = imem05_in[123:120];
    80: op1_01_in17 = reg_0303;
    81: op1_01_in17 = reg_0246;
    82: op1_01_in17 = reg_0201;
    83: op1_01_in17 = reg_0262;
    84: op1_01_in17 = reg_0156;
    85: op1_01_in17 = reg_0915;
    86: op1_01_in17 = imem01_in[119:116];
    87: op1_01_in17 = imem07_in[59:56];
    88: op1_01_in17 = reg_0021;
    89: op1_01_in17 = imem01_in[123:120];
    90: op1_01_in17 = reg_0781;
    91: op1_01_in17 = reg_0427;
    93: op1_01_in17 = reg_0318;
    94: op1_01_in17 = reg_0609;
    95: op1_01_in17 = reg_0767;
    96: op1_01_in17 = reg_0233;
    97: op1_01_in17 = reg_0110;
    default: op1_01_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv17 = 1;
    7: op1_01_inv17 = 1;
    15: op1_01_inv17 = 1;
    16: op1_01_inv17 = 1;
    17: op1_01_inv17 = 1;
    18: op1_01_inv17 = 1;
    21: op1_01_inv17 = 1;
    22: op1_01_inv17 = 1;
    23: op1_01_inv17 = 1;
    24: op1_01_inv17 = 1;
    25: op1_01_inv17 = 1;
    27: op1_01_inv17 = 1;
    28: op1_01_inv17 = 1;
    29: op1_01_inv17 = 1;
    32: op1_01_inv17 = 1;
    33: op1_01_inv17 = 1;
    35: op1_01_inv17 = 1;
    39: op1_01_inv17 = 1;
    41: op1_01_inv17 = 1;
    42: op1_01_inv17 = 1;
    46: op1_01_inv17 = 1;
    48: op1_01_inv17 = 1;
    50: op1_01_inv17 = 1;
    51: op1_01_inv17 = 1;
    56: op1_01_inv17 = 1;
    57: op1_01_inv17 = 1;
    58: op1_01_inv17 = 1;
    59: op1_01_inv17 = 1;
    61: op1_01_inv17 = 1;
    66: op1_01_inv17 = 1;
    67: op1_01_inv17 = 1;
    69: op1_01_inv17 = 1;
    76: op1_01_inv17 = 1;
    83: op1_01_inv17 = 1;
    85: op1_01_inv17 = 1;
    86: op1_01_inv17 = 1;
    87: op1_01_inv17 = 1;
    88: op1_01_inv17 = 1;
    90: op1_01_inv17 = 1;
    93: op1_01_inv17 = 1;
    96: op1_01_inv17 = 1;
    default: op1_01_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in18 = imem02_in[75:72];
    6: op1_01_in18 = reg_0434;
    7: op1_01_in18 = imem03_in[3:0];
    8: op1_01_in18 = reg_0405;
    9: op1_01_in18 = imem01_in[63:60];
    10: op1_01_in18 = reg_0598;
    11: op1_01_in18 = reg_0319;
    12: op1_01_in18 = reg_0188;
    13: op1_01_in18 = reg_0329;
    14: op1_01_in18 = reg_0172;
    15: op1_01_in18 = imem02_in[51:48];
    16: op1_01_in18 = reg_0602;
    17: op1_01_in18 = reg_0155;
    18: op1_01_in18 = imem01_in[3:0];
    20: op1_01_in18 = reg_0208;
    21: op1_01_in18 = reg_0256;
    22: op1_01_in18 = imem01_in[39:36];
    23: op1_01_in18 = reg_0086;
    24: op1_01_in18 = reg_0722;
    25: op1_01_in18 = reg_0979;
    26: op1_01_in18 = reg_0154;
    27: op1_01_in18 = reg_0586;
    28: op1_01_in18 = reg_0614;
    29: op1_01_in18 = reg_0223;
    30: op1_01_in18 = reg_0662;
    31: op1_01_in18 = imem06_in[35:32];
    32: op1_01_in18 = reg_0193;
    33: op1_01_in18 = reg_0039;
    34: op1_01_in18 = imem03_in[51:48];
    35: op1_01_in18 = imem01_in[55:52];
    37: op1_01_in18 = reg_0205;
    38: op1_01_in18 = reg_0007;
    77: op1_01_in18 = reg_0007;
    39: op1_01_in18 = reg_0643;
    40: op1_01_in18 = reg_0059;
    41: op1_01_in18 = imem04_in[43:40];
    42: op1_01_in18 = reg_0440;
    43: op1_01_in18 = reg_0199;
    82: op1_01_in18 = reg_0199;
    44: op1_01_in18 = reg_0318;
    45: op1_01_in18 = imem05_in[3:0];
    46: op1_01_in18 = reg_0426;
    47: op1_01_in18 = reg_0865;
    48: op1_01_in18 = reg_0984;
    49: op1_01_in18 = reg_0726;
    50: op1_01_in18 = reg_0157;
    66: op1_01_in18 = reg_0157;
    51: op1_01_in18 = imem07_in[19:16];
    85: op1_01_in18 = imem07_in[19:16];
    52: op1_01_in18 = reg_0834;
    53: op1_01_in18 = reg_0296;
    54: op1_01_in18 = reg_0493;
    55: op1_01_in18 = imem06_in[67:64];
    57: op1_01_in18 = reg_0194;
    58: op1_01_in18 = imem01_in[35:32];
    59: op1_01_in18 = reg_0166;
    60: op1_01_in18 = imem03_in[15:12];
    61: op1_01_in18 = imem01_in[107:104];
    62: op1_01_in18 = reg_0372;
    63: op1_01_in18 = reg_0022;
    64: op1_01_in18 = imem07_in[95:92];
    65: op1_01_in18 = reg_0589;
    67: op1_01_in18 = reg_0640;
    69: op1_01_in18 = imem04_in[67:64];
    70: op1_01_in18 = imem06_in[95:92];
    71: op1_01_in18 = reg_0211;
    72: op1_01_in18 = imem06_in[51:48];
    75: op1_01_in18 = imem01_in[15:12];
    76: op1_01_in18 = imem03_in[111:108];
    78: op1_01_in18 = reg_0636;
    80: op1_01_in18 = reg_0325;
    81: op1_01_in18 = reg_1023;
    83: op1_01_in18 = reg_0817;
    84: op1_01_in18 = reg_0912;
    86: op1_01_in18 = reg_0105;
    87: op1_01_in18 = imem07_in[123:120];
    88: op1_01_in18 = reg_1011;
    89: op1_01_in18 = reg_0904;
    90: op1_01_in18 = reg_0177;
    91: op1_01_in18 = reg_0868;
    93: op1_01_in18 = imem04_in[3:0];
    94: op1_01_in18 = reg_0051;
    95: op1_01_in18 = reg_0982;
    96: op1_01_in18 = reg_0523;
    97: op1_01_in18 = imem02_in[11:8];
    default: op1_01_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv18 = 1;
    6: op1_01_inv18 = 1;
    7: op1_01_inv18 = 1;
    9: op1_01_inv18 = 1;
    10: op1_01_inv18 = 1;
    12: op1_01_inv18 = 1;
    14: op1_01_inv18 = 1;
    15: op1_01_inv18 = 1;
    18: op1_01_inv18 = 1;
    20: op1_01_inv18 = 1;
    23: op1_01_inv18 = 1;
    26: op1_01_inv18 = 1;
    30: op1_01_inv18 = 1;
    31: op1_01_inv18 = 1;
    32: op1_01_inv18 = 1;
    38: op1_01_inv18 = 1;
    40: op1_01_inv18 = 1;
    43: op1_01_inv18 = 1;
    44: op1_01_inv18 = 1;
    49: op1_01_inv18 = 1;
    50: op1_01_inv18 = 1;
    52: op1_01_inv18 = 1;
    53: op1_01_inv18 = 1;
    54: op1_01_inv18 = 1;
    58: op1_01_inv18 = 1;
    60: op1_01_inv18 = 1;
    61: op1_01_inv18 = 1;
    62: op1_01_inv18 = 1;
    64: op1_01_inv18 = 1;
    67: op1_01_inv18 = 1;
    70: op1_01_inv18 = 1;
    71: op1_01_inv18 = 1;
    76: op1_01_inv18 = 1;
    80: op1_01_inv18 = 1;
    83: op1_01_inv18 = 1;
    88: op1_01_inv18 = 1;
    89: op1_01_inv18 = 1;
    90: op1_01_inv18 = 1;
    93: op1_01_inv18 = 1;
    95: op1_01_inv18 = 1;
    97: op1_01_inv18 = 1;
    default: op1_01_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in19 = reg_0658;
    6: op1_01_in19 = reg_0437;
    42: op1_01_in19 = reg_0437;
    7: op1_01_in19 = imem03_in[75:72];
    8: op1_01_in19 = reg_0404;
    9: op1_01_in19 = imem01_in[71:68];
    10: op1_01_in19 = reg_0586;
    11: op1_01_in19 = reg_0398;
    12: op1_01_in19 = reg_0207;
    13: op1_01_in19 = reg_0353;
    14: op1_01_in19 = reg_0181;
    15: op1_01_in19 = imem02_in[111:108];
    16: op1_01_in19 = reg_0579;
    17: op1_01_in19 = imem06_in[31:28];
    18: op1_01_in19 = imem01_in[75:72];
    20: op1_01_in19 = reg_0210;
    21: op1_01_in19 = reg_0816;
    22: op1_01_in19 = imem01_in[63:60];
    23: op1_01_in19 = reg_0084;
    24: op1_01_in19 = reg_0716;
    25: op1_01_in19 = reg_0999;
    26: op1_01_in19 = reg_0139;
    27: op1_01_in19 = reg_0572;
    28: op1_01_in19 = reg_0624;
    29: op1_01_in19 = reg_0236;
    30: op1_01_in19 = reg_0636;
    31: op1_01_in19 = imem06_in[67:64];
    32: op1_01_in19 = reg_0198;
    71: op1_01_in19 = reg_0198;
    33: op1_01_in19 = reg_0096;
    34: op1_01_in19 = reg_1007;
    35: op1_01_in19 = imem01_in[83:80];
    37: op1_01_in19 = imem01_in[11:8];
    38: op1_01_in19 = reg_0758;
    39: op1_01_in19 = reg_0652;
    40: op1_01_in19 = reg_0279;
    41: op1_01_in19 = imem04_in[63:60];
    43: op1_01_in19 = reg_0197;
    44: op1_01_in19 = reg_0817;
    45: op1_01_in19 = imem05_in[51:48];
    46: op1_01_in19 = reg_0428;
    80: op1_01_in19 = reg_0428;
    47: op1_01_in19 = reg_0772;
    48: op1_01_in19 = reg_1001;
    49: op1_01_in19 = reg_0709;
    50: op1_01_in19 = reg_0158;
    51: op1_01_in19 = imem07_in[23:20];
    52: op1_01_in19 = reg_0554;
    53: op1_01_in19 = imem05_in[63:60];
    54: op1_01_in19 = reg_0336;
    55: op1_01_in19 = imem06_in[83:80];
    57: op1_01_in19 = reg_0213;
    58: op1_01_in19 = imem01_in[99:96];
    60: op1_01_in19 = imem03_in[19:16];
    61: op1_01_in19 = reg_0510;
    62: op1_01_in19 = reg_0506;
    63: op1_01_in19 = reg_0259;
    64: op1_01_in19 = reg_0710;
    65: op1_01_in19 = reg_0640;
    66: op1_01_in19 = reg_0173;
    67: op1_01_in19 = reg_0838;
    69: op1_01_in19 = imem04_in[83:80];
    70: op1_01_in19 = reg_0025;
    72: op1_01_in19 = imem06_in[63:60];
    75: op1_01_in19 = imem01_in[31:28];
    76: op1_01_in19 = imem03_in[119:116];
    77: op1_01_in19 = imem03_in[7:4];
    78: op1_01_in19 = reg_0226;
    81: op1_01_in19 = reg_0501;
    82: op1_01_in19 = imem01_in[51:48];
    83: op1_01_in19 = reg_0692;
    84: op1_01_in19 = reg_0540;
    85: op1_01_in19 = imem07_in[79:76];
    86: op1_01_in19 = reg_0968;
    87: op1_01_in19 = imem07_in[127:124];
    88: op1_01_in19 = reg_0297;
    89: op1_01_in19 = reg_0225;
    90: op1_01_in19 = reg_0782;
    91: op1_01_in19 = reg_0431;
    93: op1_01_in19 = imem04_in[15:12];
    94: op1_01_in19 = reg_0779;
    95: op1_01_in19 = reg_0613;
    96: op1_01_in19 = reg_0825;
    97: op1_01_in19 = imem02_in[31:28];
    default: op1_01_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_01_inv19 = 1;
    9: op1_01_inv19 = 1;
    10: op1_01_inv19 = 1;
    11: op1_01_inv19 = 1;
    13: op1_01_inv19 = 1;
    14: op1_01_inv19 = 1;
    15: op1_01_inv19 = 1;
    16: op1_01_inv19 = 1;
    18: op1_01_inv19 = 1;
    20: op1_01_inv19 = 1;
    22: op1_01_inv19 = 1;
    27: op1_01_inv19 = 1;
    28: op1_01_inv19 = 1;
    29: op1_01_inv19 = 1;
    34: op1_01_inv19 = 1;
    37: op1_01_inv19 = 1;
    39: op1_01_inv19 = 1;
    40: op1_01_inv19 = 1;
    41: op1_01_inv19 = 1;
    48: op1_01_inv19 = 1;
    53: op1_01_inv19 = 1;
    54: op1_01_inv19 = 1;
    57: op1_01_inv19 = 1;
    62: op1_01_inv19 = 1;
    64: op1_01_inv19 = 1;
    65: op1_01_inv19 = 1;
    67: op1_01_inv19 = 1;
    70: op1_01_inv19 = 1;
    71: op1_01_inv19 = 1;
    72: op1_01_inv19 = 1;
    80: op1_01_inv19 = 1;
    82: op1_01_inv19 = 1;
    84: op1_01_inv19 = 1;
    85: op1_01_inv19 = 1;
    86: op1_01_inv19 = 1;
    87: op1_01_inv19 = 1;
    88: op1_01_inv19 = 1;
    91: op1_01_inv19 = 1;
    93: op1_01_inv19 = 1;
    97: op1_01_inv19 = 1;
    default: op1_01_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in20 = reg_0646;
    6: op1_01_in20 = reg_0438;
    42: op1_01_in20 = reg_0438;
    7: op1_01_in20 = imem03_in[107:104];
    8: op1_01_in20 = reg_0406;
    9: op1_01_in20 = imem01_in[75:72];
    82: op1_01_in20 = imem01_in[75:72];
    10: op1_01_in20 = reg_0582;
    11: op1_01_in20 = reg_0374;
    12: op1_01_in20 = reg_0201;
    13: op1_01_in20 = reg_0342;
    14: op1_01_in20 = reg_0169;
    15: op1_01_in20 = reg_0650;
    16: op1_01_in20 = reg_0563;
    17: op1_01_in20 = imem06_in[79:76];
    18: op1_01_in20 = imem01_in[115:112];
    20: op1_01_in20 = reg_0189;
    21: op1_01_in20 = reg_0275;
    22: op1_01_in20 = imem01_in[103:100];
    23: op1_01_in20 = reg_0077;
    24: op1_01_in20 = reg_0704;
    25: op1_01_in20 = reg_0997;
    26: op1_01_in20 = reg_0138;
    27: op1_01_in20 = reg_0569;
    28: op1_01_in20 = reg_0617;
    29: op1_01_in20 = reg_0249;
    30: op1_01_in20 = reg_0865;
    31: op1_01_in20 = reg_0605;
    32: op1_01_in20 = imem01_in[3:0];
    33: op1_01_in20 = reg_0762;
    34: op1_01_in20 = reg_0327;
    35: op1_01_in20 = imem01_in[107:104];
    37: op1_01_in20 = imem01_in[39:36];
    75: op1_01_in20 = imem01_in[39:36];
    38: op1_01_in20 = reg_0761;
    47: op1_01_in20 = reg_0761;
    39: op1_01_in20 = reg_0837;
    40: op1_01_in20 = reg_0528;
    41: op1_01_in20 = imem04_in[71:68];
    43: op1_01_in20 = imem01_in[23:20];
    44: op1_01_in20 = reg_0093;
    45: op1_01_in20 = imem05_in[63:60];
    46: op1_01_in20 = reg_0641;
    48: op1_01_in20 = reg_0986;
    49: op1_01_in20 = reg_0433;
    51: op1_01_in20 = imem07_in[39:36];
    52: op1_01_in20 = reg_0517;
    53: op1_01_in20 = imem05_in[103:100];
    54: op1_01_in20 = reg_0094;
    55: op1_01_in20 = imem06_in[103:100];
    57: op1_01_in20 = reg_0199;
    58: op1_01_in20 = imem01_in[119:116];
    60: op1_01_in20 = imem03_in[47:44];
    61: op1_01_in20 = reg_0285;
    62: op1_01_in20 = reg_0840;
    63: op1_01_in20 = reg_0488;
    64: op1_01_in20 = reg_0731;
    65: op1_01_in20 = reg_0838;
    67: op1_01_in20 = reg_0431;
    69: op1_01_in20 = imem04_in[95:92];
    70: op1_01_in20 = reg_0926;
    71: op1_01_in20 = reg_0202;
    72: op1_01_in20 = imem06_in[67:64];
    76: op1_01_in20 = reg_0535;
    77: op1_01_in20 = imem03_in[67:64];
    78: op1_01_in20 = reg_0583;
    80: op1_01_in20 = reg_0599;
    81: op1_01_in20 = reg_1043;
    83: op1_01_in20 = reg_1030;
    84: op1_01_in20 = reg_0882;
    85: op1_01_in20 = imem07_in[107:104];
    86: op1_01_in20 = reg_1035;
    87: op1_01_in20 = reg_0726;
    88: op1_01_in20 = reg_0895;
    89: op1_01_in20 = reg_0607;
    90: op1_01_in20 = imem07_in[19:16];
    91: op1_01_in20 = reg_0182;
    93: op1_01_in20 = imem04_in[35:32];
    94: op1_01_in20 = reg_0588;
    95: op1_01_in20 = reg_0961;
    96: op1_01_in20 = reg_0547;
    97: op1_01_in20 = imem02_in[79:76];
    default: op1_01_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv20 = 1;
    7: op1_01_inv20 = 1;
    8: op1_01_inv20 = 1;
    9: op1_01_inv20 = 1;
    10: op1_01_inv20 = 1;
    15: op1_01_inv20 = 1;
    20: op1_01_inv20 = 1;
    21: op1_01_inv20 = 1;
    22: op1_01_inv20 = 1;
    23: op1_01_inv20 = 1;
    29: op1_01_inv20 = 1;
    32: op1_01_inv20 = 1;
    33: op1_01_inv20 = 1;
    34: op1_01_inv20 = 1;
    35: op1_01_inv20 = 1;
    37: op1_01_inv20 = 1;
    38: op1_01_inv20 = 1;
    40: op1_01_inv20 = 1;
    43: op1_01_inv20 = 1;
    44: op1_01_inv20 = 1;
    45: op1_01_inv20 = 1;
    46: op1_01_inv20 = 1;
    47: op1_01_inv20 = 1;
    48: op1_01_inv20 = 1;
    49: op1_01_inv20 = 1;
    51: op1_01_inv20 = 1;
    53: op1_01_inv20 = 1;
    55: op1_01_inv20 = 1;
    58: op1_01_inv20 = 1;
    61: op1_01_inv20 = 1;
    62: op1_01_inv20 = 1;
    69: op1_01_inv20 = 1;
    70: op1_01_inv20 = 1;
    71: op1_01_inv20 = 1;
    75: op1_01_inv20 = 1;
    76: op1_01_inv20 = 1;
    77: op1_01_inv20 = 1;
    78: op1_01_inv20 = 1;
    82: op1_01_inv20 = 1;
    83: op1_01_inv20 = 1;
    84: op1_01_inv20 = 1;
    86: op1_01_inv20 = 1;
    88: op1_01_inv20 = 1;
    89: op1_01_inv20 = 1;
    90: op1_01_inv20 = 1;
    91: op1_01_inv20 = 1;
    93: op1_01_inv20 = 1;
    94: op1_01_inv20 = 1;
    96: op1_01_inv20 = 1;
    default: op1_01_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in21 = reg_0647;
    6: op1_01_in21 = reg_0162;
    42: op1_01_in21 = reg_0162;
    7: op1_01_in21 = reg_0591;
    8: op1_01_in21 = reg_0028;
    9: op1_01_in21 = imem01_in[95:92];
    10: op1_01_in21 = reg_0596;
    11: op1_01_in21 = reg_0991;
    12: op1_01_in21 = imem01_in[31:28];
    43: op1_01_in21 = imem01_in[31:28];
    13: op1_01_in21 = reg_0082;
    14: op1_01_in21 = reg_0183;
    15: op1_01_in21 = reg_0658;
    16: op1_01_in21 = reg_0576;
    17: op1_01_in21 = imem06_in[83:80];
    18: op1_01_in21 = reg_0013;
    35: op1_01_in21 = reg_0013;
    20: op1_01_in21 = reg_0201;
    21: op1_01_in21 = reg_1046;
    22: op1_01_in21 = imem01_in[107:104];
    23: op1_01_in21 = reg_0079;
    24: op1_01_in21 = reg_0721;
    25: op1_01_in21 = imem04_in[15:12];
    26: op1_01_in21 = imem06_in[23:20];
    27: op1_01_in21 = reg_0594;
    28: op1_01_in21 = reg_0621;
    29: op1_01_in21 = reg_1039;
    30: op1_01_in21 = reg_0098;
    31: op1_01_in21 = reg_0606;
    32: op1_01_in21 = imem01_in[27:24];
    33: op1_01_in21 = reg_0007;
    34: op1_01_in21 = reg_0311;
    37: op1_01_in21 = imem01_in[67:64];
    38: op1_01_in21 = reg_0085;
    39: op1_01_in21 = reg_0330;
    40: op1_01_in21 = reg_0774;
    41: op1_01_in21 = imem04_in[91:88];
    44: op1_01_in21 = reg_0762;
    45: op1_01_in21 = imem05_in[71:68];
    46: op1_01_in21 = reg_0532;
    47: op1_01_in21 = reg_0091;
    48: op1_01_in21 = reg_0990;
    49: op1_01_in21 = reg_0047;
    51: op1_01_in21 = imem07_in[127:124];
    52: op1_01_in21 = reg_0578;
    53: op1_01_in21 = reg_0963;
    54: op1_01_in21 = reg_0819;
    55: op1_01_in21 = imem06_in[107:104];
    57: op1_01_in21 = imem01_in[47:44];
    58: op1_01_in21 = reg_0918;
    60: op1_01_in21 = imem03_in[87:84];
    61: op1_01_in21 = reg_0249;
    62: op1_01_in21 = reg_0484;
    63: op1_01_in21 = reg_0508;
    64: op1_01_in21 = reg_0725;
    65: op1_01_in21 = reg_0431;
    67: op1_01_in21 = reg_0180;
    69: op1_01_in21 = imem04_in[107:104];
    70: op1_01_in21 = reg_0392;
    71: op1_01_in21 = imem01_in[15:12];
    72: op1_01_in21 = imem06_in[95:92];
    75: op1_01_in21 = imem01_in[63:60];
    76: op1_01_in21 = reg_0245;
    77: op1_01_in21 = imem03_in[119:116];
    78: op1_01_in21 = reg_0940;
    80: op1_01_in21 = reg_0181;
    81: op1_01_in21 = reg_0829;
    82: op1_01_in21 = imem01_in[79:76];
    83: op1_01_in21 = reg_0439;
    84: op1_01_in21 = reg_0586;
    85: op1_01_in21 = reg_0159;
    86: op1_01_in21 = reg_0862;
    87: op1_01_in21 = reg_0374;
    88: op1_01_in21 = reg_0792;
    89: op1_01_in21 = reg_0216;
    90: op1_01_in21 = imem07_in[31:28];
    93: op1_01_in21 = imem04_in[51:48];
    94: op1_01_in21 = reg_0979;
    95: op1_01_in21 = reg_0523;
    96: op1_01_in21 = reg_0396;
    97: op1_01_in21 = imem02_in[95:92];
    default: op1_01_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    13: op1_01_inv21 = 1;
    14: op1_01_inv21 = 1;
    15: op1_01_inv21 = 1;
    21: op1_01_inv21 = 1;
    23: op1_01_inv21 = 1;
    25: op1_01_inv21 = 1;
    29: op1_01_inv21 = 1;
    30: op1_01_inv21 = 1;
    33: op1_01_inv21 = 1;
    34: op1_01_inv21 = 1;
    35: op1_01_inv21 = 1;
    37: op1_01_inv21 = 1;
    38: op1_01_inv21 = 1;
    40: op1_01_inv21 = 1;
    41: op1_01_inv21 = 1;
    47: op1_01_inv21 = 1;
    55: op1_01_inv21 = 1;
    57: op1_01_inv21 = 1;
    58: op1_01_inv21 = 1;
    60: op1_01_inv21 = 1;
    63: op1_01_inv21 = 1;
    64: op1_01_inv21 = 1;
    65: op1_01_inv21 = 1;
    67: op1_01_inv21 = 1;
    69: op1_01_inv21 = 1;
    71: op1_01_inv21 = 1;
    77: op1_01_inv21 = 1;
    81: op1_01_inv21 = 1;
    82: op1_01_inv21 = 1;
    85: op1_01_inv21 = 1;
    86: op1_01_inv21 = 1;
    90: op1_01_inv21 = 1;
    96: op1_01_inv21 = 1;
    default: op1_01_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in22 = reg_0648;
    6: op1_01_in22 = reg_0163;
    7: op1_01_in22 = reg_0589;
    8: op1_01_in22 = reg_0037;
    9: op1_01_in22 = reg_0506;
    10: op1_01_in22 = reg_0583;
    11: op1_01_in22 = reg_0995;
    12: op1_01_in22 = imem01_in[39:36];
    13: op1_01_in22 = imem03_in[71:68];
    14: op1_01_in22 = reg_0166;
    15: op1_01_in22 = reg_0653;
    16: op1_01_in22 = reg_0394;
    17: op1_01_in22 = imem06_in[91:88];
    18: op1_01_in22 = reg_1053;
    20: op1_01_in22 = reg_0213;
    21: op1_01_in22 = reg_0896;
    22: op1_01_in22 = reg_0013;
    23: op1_01_in22 = imem03_in[23:20];
    62: op1_01_in22 = imem03_in[23:20];
    24: op1_01_in22 = reg_0713;
    25: op1_01_in22 = imem04_in[19:16];
    26: op1_01_in22 = imem06_in[59:56];
    27: op1_01_in22 = reg_0597;
    28: op1_01_in22 = reg_0611;
    29: op1_01_in22 = reg_1032;
    30: op1_01_in22 = reg_0335;
    31: op1_01_in22 = reg_0609;
    32: op1_01_in22 = imem01_in[107:104];
    33: op1_01_in22 = reg_0088;
    34: op1_01_in22 = reg_0991;
    35: op1_01_in22 = reg_0235;
    37: op1_01_in22 = imem01_in[111:108];
    38: op1_01_in22 = reg_0016;
    39: op1_01_in22 = reg_0098;
    40: op1_01_in22 = reg_0855;
    41: op1_01_in22 = imem04_in[107:104];
    42: op1_01_in22 = reg_0168;
    43: op1_01_in22 = imem01_in[51:48];
    44: op1_01_in22 = reg_0867;
    45: op1_01_in22 = imem05_in[75:72];
    46: op1_01_in22 = reg_0431;
    47: op1_01_in22 = reg_0049;
    48: op1_01_in22 = imem04_in[11:8];
    49: op1_01_in22 = reg_0641;
    51: op1_01_in22 = reg_0728;
    52: op1_01_in22 = reg_0864;
    53: op1_01_in22 = reg_0022;
    54: op1_01_in22 = reg_0130;
    55: op1_01_in22 = imem06_in[123:120];
    57: op1_01_in22 = imem01_in[55:52];
    58: op1_01_in22 = reg_0586;
    60: op1_01_in22 = imem03_in[95:92];
    61: op1_01_in22 = reg_0521;
    63: op1_01_in22 = reg_0404;
    64: op1_01_in22 = reg_0712;
    65: op1_01_in22 = reg_0180;
    67: op1_01_in22 = reg_0164;
    69: op1_01_in22 = imem04_in[115:112];
    70: op1_01_in22 = reg_0698;
    71: op1_01_in22 = imem01_in[31:28];
    72: op1_01_in22 = imem06_in[103:100];
    75: op1_01_in22 = imem01_in[71:68];
    76: op1_01_in22 = reg_0046;
    77: op1_01_in22 = imem03_in[123:120];
    78: op1_01_in22 = reg_0806;
    80: op1_01_in22 = reg_0184;
    81: op1_01_in22 = reg_0500;
    82: op1_01_in22 = imem01_in[99:96];
    83: op1_01_in22 = reg_0863;
    84: op1_01_in22 = reg_0537;
    85: op1_01_in22 = reg_0374;
    86: op1_01_in22 = reg_0225;
    87: op1_01_in22 = reg_0247;
    88: op1_01_in22 = reg_0595;
    89: op1_01_in22 = reg_1031;
    90: op1_01_in22 = imem07_in[43:40];
    93: op1_01_in22 = imem04_in[55:52];
    94: op1_01_in22 = reg_0445;
    95: op1_01_in22 = reg_0986;
    96: op1_01_in22 = imem04_in[7:4];
    97: op1_01_in22 = imem02_in[119:116];
    default: op1_01_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_01_inv22 = 1;
    9: op1_01_inv22 = 1;
    10: op1_01_inv22 = 1;
    11: op1_01_inv22 = 1;
    13: op1_01_inv22 = 1;
    16: op1_01_inv22 = 1;
    17: op1_01_inv22 = 1;
    20: op1_01_inv22 = 1;
    21: op1_01_inv22 = 1;
    22: op1_01_inv22 = 1;
    23: op1_01_inv22 = 1;
    24: op1_01_inv22 = 1;
    25: op1_01_inv22 = 1;
    27: op1_01_inv22 = 1;
    28: op1_01_inv22 = 1;
    32: op1_01_inv22 = 1;
    37: op1_01_inv22 = 1;
    39: op1_01_inv22 = 1;
    41: op1_01_inv22 = 1;
    42: op1_01_inv22 = 1;
    44: op1_01_inv22 = 1;
    48: op1_01_inv22 = 1;
    51: op1_01_inv22 = 1;
    52: op1_01_inv22 = 1;
    60: op1_01_inv22 = 1;
    61: op1_01_inv22 = 1;
    63: op1_01_inv22 = 1;
    65: op1_01_inv22 = 1;
    67: op1_01_inv22 = 1;
    71: op1_01_inv22 = 1;
    75: op1_01_inv22 = 1;
    77: op1_01_inv22 = 1;
    78: op1_01_inv22 = 1;
    81: op1_01_inv22 = 1;
    83: op1_01_inv22 = 1;
    85: op1_01_inv22 = 1;
    86: op1_01_inv22 = 1;
    87: op1_01_inv22 = 1;
    88: op1_01_inv22 = 1;
    89: op1_01_inv22 = 1;
    90: op1_01_inv22 = 1;
    93: op1_01_inv22 = 1;
    94: op1_01_inv22 = 1;
    95: op1_01_inv22 = 1;
    96: op1_01_inv22 = 1;
    default: op1_01_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in23 = reg_0649;
    6: op1_01_in23 = reg_0168;
    7: op1_01_in23 = reg_0593;
    52: op1_01_in23 = reg_0593;
    8: op1_01_in23 = reg_0029;
    9: op1_01_in23 = reg_0510;
    10: op1_01_in23 = reg_0585;
    11: op1_01_in23 = reg_0984;
    12: op1_01_in23 = imem01_in[71:68];
    43: op1_01_in23 = imem01_in[71:68];
    13: op1_01_in23 = reg_0598;
    14: op1_01_in23 = reg_0157;
    42: op1_01_in23 = reg_0157;
    15: op1_01_in23 = reg_0654;
    16: op1_01_in23 = reg_0362;
    17: op1_01_in23 = reg_0613;
    18: op1_01_in23 = reg_1050;
    20: op1_01_in23 = reg_0190;
    21: op1_01_in23 = reg_0831;
    22: op1_01_in23 = reg_1049;
    23: op1_01_in23 = imem03_in[43:40];
    24: op1_01_in23 = reg_0430;
    25: op1_01_in23 = imem04_in[51:48];
    26: op1_01_in23 = imem06_in[119:116];
    27: op1_01_in23 = reg_0570;
    28: op1_01_in23 = reg_0633;
    29: op1_01_in23 = reg_0227;
    30: op1_01_in23 = reg_0876;
    31: op1_01_in23 = reg_0618;
    32: op1_01_in23 = imem01_in[119:116];
    33: op1_01_in23 = reg_0086;
    34: op1_01_in23 = reg_0974;
    35: op1_01_in23 = reg_0779;
    37: op1_01_in23 = imem01_in[115:112];
    38: op1_01_in23 = reg_0077;
    39: op1_01_in23 = reg_0338;
    40: op1_01_in23 = imem05_in[83:80];
    41: op1_01_in23 = imem04_in[111:108];
    44: op1_01_in23 = reg_0085;
    45: op1_01_in23 = reg_0973;
    46: op1_01_in23 = reg_0181;
    47: op1_01_in23 = reg_0084;
    48: op1_01_in23 = imem04_in[55:52];
    49: op1_01_in23 = reg_0158;
    51: op1_01_in23 = reg_0716;
    53: op1_01_in23 = reg_0252;
    54: op1_01_in23 = imem06_in[3:0];
    55: op1_01_in23 = reg_0407;
    57: op1_01_in23 = imem01_in[75:72];
    58: op1_01_in23 = reg_0223;
    60: op1_01_in23 = reg_0006;
    61: op1_01_in23 = reg_0610;
    62: op1_01_in23 = imem03_in[39:36];
    63: op1_01_in23 = reg_0153;
    64: op1_01_in23 = reg_0705;
    65: op1_01_in23 = reg_0160;
    67: op1_01_in23 = reg_0185;
    69: op1_01_in23 = reg_0301;
    70: op1_01_in23 = reg_0699;
    71: op1_01_in23 = imem01_in[63:60];
    72: op1_01_in23 = reg_0294;
    75: op1_01_in23 = imem01_in[87:84];
    76: op1_01_in23 = reg_0396;
    77: op1_01_in23 = reg_0060;
    78: op1_01_in23 = reg_0950;
    81: op1_01_in23 = reg_0615;
    82: op1_01_in23 = imem01_in[107:104];
    83: op1_01_in23 = reg_0804;
    84: op1_01_in23 = reg_0802;
    85: op1_01_in23 = reg_0718;
    86: op1_01_in23 = reg_0607;
    87: op1_01_in23 = reg_0759;
    88: op1_01_in23 = reg_0264;
    89: op1_01_in23 = reg_0925;
    90: op1_01_in23 = imem07_in[67:64];
    93: op1_01_in23 = imem04_in[59:56];
    94: op1_01_in23 = imem04_in[7:4];
    95: op1_01_in23 = reg_0445;
    96: op1_01_in23 = imem04_in[15:12];
    97: op1_01_in23 = reg_0334;
    default: op1_01_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv23 = 1;
    14: op1_01_inv23 = 1;
    16: op1_01_inv23 = 1;
    17: op1_01_inv23 = 1;
    22: op1_01_inv23 = 1;
    23: op1_01_inv23 = 1;
    24: op1_01_inv23 = 1;
    25: op1_01_inv23 = 1;
    28: op1_01_inv23 = 1;
    29: op1_01_inv23 = 1;
    33: op1_01_inv23 = 1;
    35: op1_01_inv23 = 1;
    37: op1_01_inv23 = 1;
    38: op1_01_inv23 = 1;
    39: op1_01_inv23 = 1;
    40: op1_01_inv23 = 1;
    42: op1_01_inv23 = 1;
    48: op1_01_inv23 = 1;
    53: op1_01_inv23 = 1;
    55: op1_01_inv23 = 1;
    57: op1_01_inv23 = 1;
    58: op1_01_inv23 = 1;
    60: op1_01_inv23 = 1;
    64: op1_01_inv23 = 1;
    65: op1_01_inv23 = 1;
    70: op1_01_inv23 = 1;
    71: op1_01_inv23 = 1;
    81: op1_01_inv23 = 1;
    83: op1_01_inv23 = 1;
    84: op1_01_inv23 = 1;
    85: op1_01_inv23 = 1;
    87: op1_01_inv23 = 1;
    88: op1_01_inv23 = 1;
    89: op1_01_inv23 = 1;
    90: op1_01_inv23 = 1;
    93: op1_01_inv23 = 1;
    95: op1_01_inv23 = 1;
    96: op1_01_inv23 = 1;
    97: op1_01_inv23 = 1;
    default: op1_01_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in24 = reg_0659;
    6: op1_01_in24 = reg_0170;
    7: op1_01_in24 = reg_0580;
    10: op1_01_in24 = reg_0580;
    8: op1_01_in24 = reg_0038;
    9: op1_01_in24 = reg_0232;
    11: op1_01_in24 = reg_0999;
    12: op1_01_in24 = imem01_in[95:92];
    13: op1_01_in24 = reg_0602;
    14: op1_01_in24 = reg_0173;
    49: op1_01_in24 = reg_0173;
    15: op1_01_in24 = reg_0656;
    16: op1_01_in24 = reg_0373;
    17: op1_01_in24 = reg_0605;
    18: op1_01_in24 = reg_1039;
    20: op1_01_in24 = imem01_in[51:48];
    21: op1_01_in24 = reg_0497;
    22: op1_01_in24 = reg_0735;
    23: op1_01_in24 = imem03_in[83:80];
    62: op1_01_in24 = imem03_in[83:80];
    24: op1_01_in24 = reg_0419;
    25: op1_01_in24 = imem04_in[67:64];
    93: op1_01_in24 = imem04_in[67:64];
    26: op1_01_in24 = imem06_in[127:124];
    27: op1_01_in24 = reg_0394;
    28: op1_01_in24 = reg_0618;
    29: op1_01_in24 = reg_1040;
    30: op1_01_in24 = reg_0506;
    31: op1_01_in24 = reg_0627;
    32: op1_01_in24 = reg_0239;
    33: op1_01_in24 = reg_0291;
    38: op1_01_in24 = reg_0291;
    34: op1_01_in24 = reg_0977;
    35: op1_01_in24 = reg_0218;
    37: op1_01_in24 = imem01_in[119:116];
    75: op1_01_in24 = imem01_in[119:116];
    39: op1_01_in24 = reg_0516;
    40: op1_01_in24 = reg_0963;
    41: op1_01_in24 = reg_0511;
    43: op1_01_in24 = imem01_in[87:84];
    44: op1_01_in24 = reg_0310;
    45: op1_01_in24 = reg_0966;
    46: op1_01_in24 = reg_0161;
    47: op1_01_in24 = reg_0079;
    48: op1_01_in24 = imem04_in[59:56];
    51: op1_01_in24 = reg_0710;
    52: op1_01_in24 = imem05_in[7:4];
    53: op1_01_in24 = reg_0237;
    54: op1_01_in24 = imem06_in[11:8];
    55: op1_01_in24 = reg_0533;
    57: op1_01_in24 = imem01_in[99:96];
    58: op1_01_in24 = reg_1036;
    60: op1_01_in24 = reg_0535;
    61: op1_01_in24 = reg_1055;
    81: op1_01_in24 = reg_1055;
    63: op1_01_in24 = imem06_in[3:0];
    64: op1_01_in24 = reg_0706;
    65: op1_01_in24 = reg_0185;
    67: op1_01_in24 = reg_0176;
    69: op1_01_in24 = reg_1003;
    70: op1_01_in24 = reg_0380;
    71: op1_01_in24 = imem01_in[79:76];
    72: op1_01_in24 = reg_0338;
    76: op1_01_in24 = reg_0590;
    77: op1_01_in24 = reg_0681;
    78: op1_01_in24 = reg_0326;
    82: op1_01_in24 = reg_0122;
    83: op1_01_in24 = reg_0222;
    84: op1_01_in24 = reg_0848;
    85: op1_01_in24 = reg_0727;
    86: op1_01_in24 = reg_0501;
    87: op1_01_in24 = reg_0653;
    88: op1_01_in24 = reg_0369;
    89: op1_01_in24 = reg_0111;
    90: op1_01_in24 = reg_0726;
    94: op1_01_in24 = imem04_in[19:16];
    95: op1_01_in24 = reg_0825;
    96: op1_01_in24 = imem04_in[27:24];
    97: op1_01_in24 = reg_0536;
    default: op1_01_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv24 = 1;
    6: op1_01_inv24 = 1;
    9: op1_01_inv24 = 1;
    12: op1_01_inv24 = 1;
    15: op1_01_inv24 = 1;
    17: op1_01_inv24 = 1;
    21: op1_01_inv24 = 1;
    22: op1_01_inv24 = 1;
    24: op1_01_inv24 = 1;
    25: op1_01_inv24 = 1;
    26: op1_01_inv24 = 1;
    33: op1_01_inv24 = 1;
    34: op1_01_inv24 = 1;
    37: op1_01_inv24 = 1;
    39: op1_01_inv24 = 1;
    45: op1_01_inv24 = 1;
    49: op1_01_inv24 = 1;
    51: op1_01_inv24 = 1;
    54: op1_01_inv24 = 1;
    55: op1_01_inv24 = 1;
    57: op1_01_inv24 = 1;
    60: op1_01_inv24 = 1;
    62: op1_01_inv24 = 1;
    67: op1_01_inv24 = 1;
    69: op1_01_inv24 = 1;
    78: op1_01_inv24 = 1;
    81: op1_01_inv24 = 1;
    82: op1_01_inv24 = 1;
    83: op1_01_inv24 = 1;
    84: op1_01_inv24 = 1;
    85: op1_01_inv24 = 1;
    87: op1_01_inv24 = 1;
    88: op1_01_inv24 = 1;
    89: op1_01_inv24 = 1;
    93: op1_01_inv24 = 1;
    95: op1_01_inv24 = 1;
    97: op1_01_inv24 = 1;
    default: op1_01_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in25 = reg_0320;
    6: op1_01_in25 = reg_0171;
    7: op1_01_in25 = reg_0576;
    8: op1_01_in25 = imem07_in[39:36];
    9: op1_01_in25 = reg_0249;
    10: op1_01_in25 = reg_0578;
    11: op1_01_in25 = reg_1000;
    12: op1_01_in25 = imem01_in[127:124];
    13: op1_01_in25 = reg_0579;
    15: op1_01_in25 = reg_0665;
    16: op1_01_in25 = reg_0327;
    17: op1_01_in25 = reg_0611;
    18: op1_01_in25 = reg_1031;
    20: op1_01_in25 = imem01_in[71:68];
    21: op1_01_in25 = reg_0147;
    22: op1_01_in25 = reg_0242;
    35: op1_01_in25 = reg_0242;
    23: op1_01_in25 = imem03_in[99:96];
    24: op1_01_in25 = reg_0434;
    25: op1_01_in25 = imem04_in[71:68];
    48: op1_01_in25 = imem04_in[71:68];
    26: op1_01_in25 = reg_0610;
    27: op1_01_in25 = reg_0391;
    28: op1_01_in25 = reg_0632;
    29: op1_01_in25 = reg_0228;
    30: op1_01_in25 = reg_0091;
    31: op1_01_in25 = reg_0623;
    32: op1_01_in25 = reg_0299;
    33: op1_01_in25 = reg_0884;
    34: op1_01_in25 = reg_0988;
    37: op1_01_in25 = reg_0786;
    38: op1_01_in25 = imem03_in[43:40];
    39: op1_01_in25 = reg_0758;
    40: op1_01_in25 = reg_0966;
    41: op1_01_in25 = reg_0937;
    43: op1_01_in25 = imem01_in[103:100];
    44: op1_01_in25 = imem03_in[7:4];
    45: op1_01_in25 = reg_0955;
    46: op1_01_in25 = reg_0169;
    47: op1_01_in25 = imem03_in[3:0];
    51: op1_01_in25 = reg_0714;
    52: op1_01_in25 = imem05_in[11:8];
    53: op1_01_in25 = reg_0269;
    54: op1_01_in25 = imem06_in[23:20];
    55: op1_01_in25 = reg_0892;
    57: op1_01_in25 = imem01_in[111:108];
    58: op1_01_in25 = reg_0871;
    60: op1_01_in25 = reg_0099;
    61: op1_01_in25 = reg_0512;
    62: op1_01_in25 = imem03_in[91:88];
    63: op1_01_in25 = imem06_in[63:60];
    64: op1_01_in25 = reg_0303;
    67: op1_01_in25 = reg_0184;
    69: op1_01_in25 = reg_1009;
    70: op1_01_in25 = reg_1029;
    71: op1_01_in25 = imem01_in[83:80];
    72: op1_01_in25 = reg_0328;
    75: op1_01_in25 = reg_1042;
    76: op1_01_in25 = reg_0756;
    77: op1_01_in25 = reg_0572;
    78: op1_01_in25 = reg_0965;
    81: op1_01_in25 = reg_0769;
    82: op1_01_in25 = reg_1044;
    83: op1_01_in25 = reg_0619;
    84: op1_01_in25 = reg_0568;
    85: op1_01_in25 = reg_0419;
    86: op1_01_in25 = reg_0522;
    87: op1_01_in25 = reg_0325;
    88: op1_01_in25 = imem07_in[3:0];
    89: op1_01_in25 = reg_0114;
    90: op1_01_in25 = reg_0717;
    93: op1_01_in25 = imem04_in[75:72];
    94: op1_01_in25 = imem04_in[43:40];
    95: op1_01_in25 = reg_0975;
    96: op1_01_in25 = imem04_in[35:32];
    97: op1_01_in25 = reg_0348;
    default: op1_01_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_01_inv25 = 1;
    12: op1_01_inv25 = 1;
    13: op1_01_inv25 = 1;
    15: op1_01_inv25 = 1;
    21: op1_01_inv25 = 1;
    22: op1_01_inv25 = 1;
    24: op1_01_inv25 = 1;
    25: op1_01_inv25 = 1;
    26: op1_01_inv25 = 1;
    30: op1_01_inv25 = 1;
    32: op1_01_inv25 = 1;
    33: op1_01_inv25 = 1;
    38: op1_01_inv25 = 1;
    40: op1_01_inv25 = 1;
    44: op1_01_inv25 = 1;
    45: op1_01_inv25 = 1;
    46: op1_01_inv25 = 1;
    47: op1_01_inv25 = 1;
    48: op1_01_inv25 = 1;
    51: op1_01_inv25 = 1;
    52: op1_01_inv25 = 1;
    54: op1_01_inv25 = 1;
    57: op1_01_inv25 = 1;
    58: op1_01_inv25 = 1;
    60: op1_01_inv25 = 1;
    61: op1_01_inv25 = 1;
    69: op1_01_inv25 = 1;
    70: op1_01_inv25 = 1;
    71: op1_01_inv25 = 1;
    75: op1_01_inv25 = 1;
    76: op1_01_inv25 = 1;
    77: op1_01_inv25 = 1;
    78: op1_01_inv25 = 1;
    82: op1_01_inv25 = 1;
    84: op1_01_inv25 = 1;
    85: op1_01_inv25 = 1;
    87: op1_01_inv25 = 1;
    88: op1_01_inv25 = 1;
    93: op1_01_inv25 = 1;
    94: op1_01_inv25 = 1;
    95: op1_01_inv25 = 1;
    default: op1_01_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in26 = reg_0341;
    15: op1_01_in26 = reg_0341;
    7: op1_01_in26 = reg_0321;
    8: op1_01_in26 = imem07_in[43:40];
    9: op1_01_in26 = imem02_in[15:12];
    10: op1_01_in26 = reg_0394;
    11: op1_01_in26 = imem04_in[7:4];
    12: op1_01_in26 = reg_1049;
    13: op1_01_in26 = reg_0568;
    16: op1_01_in26 = reg_0985;
    17: op1_01_in26 = reg_0615;
    18: op1_01_in26 = reg_1041;
    20: op1_01_in26 = imem01_in[75:72];
    21: op1_01_in26 = reg_0133;
    22: op1_01_in26 = reg_1050;
    23: op1_01_in26 = imem03_in[123:120];
    24: op1_01_in26 = reg_0446;
    25: op1_01_in26 = imem04_in[83:80];
    26: op1_01_in26 = reg_0607;
    27: op1_01_in26 = reg_0388;
    28: op1_01_in26 = reg_0408;
    29: op1_01_in26 = reg_1038;
    30: op1_01_in26 = reg_0840;
    31: op1_01_in26 = reg_0612;
    32: op1_01_in26 = reg_0828;
    33: op1_01_in26 = imem03_in[3:0];
    34: op1_01_in26 = reg_0983;
    35: op1_01_in26 = reg_1042;
    37: op1_01_in26 = reg_0221;
    38: op1_01_in26 = imem03_in[71:68];
    39: op1_01_in26 = reg_0776;
    40: op1_01_in26 = reg_0942;
    41: op1_01_in26 = reg_1009;
    43: op1_01_in26 = reg_0544;
    44: op1_01_in26 = imem03_in[27:24];
    45: op1_01_in26 = reg_0957;
    46: op1_01_in26 = reg_0178;
    47: op1_01_in26 = imem03_in[11:8];
    48: op1_01_in26 = imem04_in[99:96];
    51: op1_01_in26 = reg_0729;
    52: op1_01_in26 = imem05_in[71:68];
    53: op1_01_in26 = reg_0147;
    54: op1_01_in26 = imem06_in[67:64];
    55: op1_01_in26 = reg_0754;
    57: op1_01_in26 = reg_0223;
    58: op1_01_in26 = reg_1052;
    60: op1_01_in26 = reg_0760;
    61: op1_01_in26 = reg_0114;
    62: op1_01_in26 = imem03_in[115:112];
    63: op1_01_in26 = imem06_in[75:72];
    64: op1_01_in26 = reg_0250;
    69: op1_01_in26 = reg_0912;
    70: op1_01_in26 = reg_0780;
    71: op1_01_in26 = imem01_in[95:92];
    72: op1_01_in26 = reg_0692;
    75: op1_01_in26 = reg_1032;
    76: op1_01_in26 = reg_0820;
    77: op1_01_in26 = reg_0327;
    78: op1_01_in26 = imem06_in[39:36];
    81: op1_01_in26 = reg_0111;
    82: op1_01_in26 = reg_0488;
    83: op1_01_in26 = reg_0370;
    84: op1_01_in26 = reg_0066;
    85: op1_01_in26 = reg_0532;
    86: op1_01_in26 = reg_0521;
    87: op1_01_in26 = reg_0428;
    88: op1_01_in26 = imem07_in[19:16];
    89: op1_01_in26 = reg_0115;
    90: op1_01_in26 = reg_0718;
    93: op1_01_in26 = imem04_in[91:88];
    94: op1_01_in26 = imem04_in[47:44];
    96: op1_01_in26 = imem04_in[47:44];
    95: op1_01_in26 = imem04_in[3:0];
    97: op1_01_in26 = reg_0765;
    default: op1_01_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv26 = 1;
    7: op1_01_inv26 = 1;
    10: op1_01_inv26 = 1;
    12: op1_01_inv26 = 1;
    13: op1_01_inv26 = 1;
    17: op1_01_inv26 = 1;
    18: op1_01_inv26 = 1;
    22: op1_01_inv26 = 1;
    24: op1_01_inv26 = 1;
    25: op1_01_inv26 = 1;
    29: op1_01_inv26 = 1;
    31: op1_01_inv26 = 1;
    32: op1_01_inv26 = 1;
    34: op1_01_inv26 = 1;
    35: op1_01_inv26 = 1;
    38: op1_01_inv26 = 1;
    40: op1_01_inv26 = 1;
    41: op1_01_inv26 = 1;
    43: op1_01_inv26 = 1;
    47: op1_01_inv26 = 1;
    52: op1_01_inv26 = 1;
    54: op1_01_inv26 = 1;
    55: op1_01_inv26 = 1;
    57: op1_01_inv26 = 1;
    58: op1_01_inv26 = 1;
    60: op1_01_inv26 = 1;
    61: op1_01_inv26 = 1;
    63: op1_01_inv26 = 1;
    64: op1_01_inv26 = 1;
    69: op1_01_inv26 = 1;
    72: op1_01_inv26 = 1;
    77: op1_01_inv26 = 1;
    81: op1_01_inv26 = 1;
    83: op1_01_inv26 = 1;
    85: op1_01_inv26 = 1;
    86: op1_01_inv26 = 1;
    87: op1_01_inv26 = 1;
    88: op1_01_inv26 = 1;
    89: op1_01_inv26 = 1;
    90: op1_01_inv26 = 1;
    93: op1_01_inv26 = 1;
    94: op1_01_inv26 = 1;
    default: op1_01_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in27 = reg_0329;
    7: op1_01_in27 = reg_0369;
    8: op1_01_in27 = imem07_in[59:56];
    9: op1_01_in27 = imem02_in[39:36];
    10: op1_01_in27 = reg_0387;
    11: op1_01_in27 = imem04_in[43:40];
    12: op1_01_in27 = reg_0735;
    13: op1_01_in27 = reg_0592;
    15: op1_01_in27 = reg_0359;
    16: op1_01_in27 = reg_0995;
    17: op1_01_in27 = reg_0356;
    18: op1_01_in27 = reg_0119;
    20: op1_01_in27 = imem01_in[95:92];
    21: op1_01_in27 = reg_0155;
    22: op1_01_in27 = reg_0230;
    23: op1_01_in27 = reg_0598;
    24: op1_01_in27 = reg_0443;
    25: op1_01_in27 = imem04_in[91:88];
    26: op1_01_in27 = reg_0630;
    27: op1_01_in27 = reg_0397;
    28: op1_01_in27 = reg_0407;
    29: op1_01_in27 = reg_0108;
    30: op1_01_in27 = reg_0884;
    31: op1_01_in27 = reg_0348;
    32: op1_01_in27 = reg_0544;
    33: op1_01_in27 = imem03_in[31:28];
    34: op1_01_in27 = reg_0997;
    35: op1_01_in27 = reg_1033;
    37: op1_01_in27 = reg_1032;
    38: op1_01_in27 = reg_1050;
    39: op1_01_in27 = reg_0079;
    40: op1_01_in27 = reg_0961;
    41: op1_01_in27 = reg_0277;
    43: op1_01_in27 = reg_0087;
    44: op1_01_in27 = imem03_in[51:48];
    45: op1_01_in27 = reg_0806;
    46: op1_01_in27 = reg_0157;
    47: op1_01_in27 = imem03_in[23:20];
    48: op1_01_in27 = imem04_in[115:112];
    51: op1_01_in27 = reg_0715;
    52: op1_01_in27 = imem05_in[87:84];
    53: op1_01_in27 = reg_0128;
    54: op1_01_in27 = imem06_in[111:108];
    55: op1_01_in27 = reg_0595;
    57: op1_01_in27 = reg_0762;
    58: op1_01_in27 = reg_0522;
    60: op1_01_in27 = reg_0298;
    61: op1_01_in27 = reg_0860;
    62: op1_01_in27 = reg_0060;
    63: op1_01_in27 = imem06_in[119:116];
    64: op1_01_in27 = reg_0047;
    69: op1_01_in27 = reg_0306;
    70: op1_01_in27 = reg_0241;
    71: op1_01_in27 = imem01_in[115:112];
    72: op1_01_in27 = reg_0534;
    75: op1_01_in27 = reg_0246;
    76: op1_01_in27 = reg_0588;
    77: op1_01_in27 = reg_0585;
    78: op1_01_in27 = imem06_in[79:76];
    81: op1_01_in27 = reg_0512;
    82: op1_01_in27 = reg_0501;
    83: op1_01_in27 = reg_0032;
    84: op1_01_in27 = reg_0815;
    85: op1_01_in27 = reg_0350;
    86: op1_01_in27 = reg_0610;
    87: op1_01_in27 = reg_0589;
    88: op1_01_in27 = imem07_in[31:28];
    89: op1_01_in27 = reg_0109;
    90: op1_01_in27 = reg_0575;
    93: op1_01_in27 = imem04_in[107:104];
    94: op1_01_in27 = imem04_in[123:120];
    95: op1_01_in27 = imem04_in[71:68];
    96: op1_01_in27 = imem04_in[55:52];
    97: op1_01_in27 = reg_0323;
    default: op1_01_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv27 = 1;
    7: op1_01_inv27 = 1;
    8: op1_01_inv27 = 1;
    11: op1_01_inv27 = 1;
    12: op1_01_inv27 = 1;
    13: op1_01_inv27 = 1;
    17: op1_01_inv27 = 1;
    18: op1_01_inv27 = 1;
    20: op1_01_inv27 = 1;
    22: op1_01_inv27 = 1;
    24: op1_01_inv27 = 1;
    28: op1_01_inv27 = 1;
    34: op1_01_inv27 = 1;
    40: op1_01_inv27 = 1;
    45: op1_01_inv27 = 1;
    48: op1_01_inv27 = 1;
    53: op1_01_inv27 = 1;
    54: op1_01_inv27 = 1;
    55: op1_01_inv27 = 1;
    57: op1_01_inv27 = 1;
    60: op1_01_inv27 = 1;
    61: op1_01_inv27 = 1;
    62: op1_01_inv27 = 1;
    69: op1_01_inv27 = 1;
    70: op1_01_inv27 = 1;
    71: op1_01_inv27 = 1;
    72: op1_01_inv27 = 1;
    78: op1_01_inv27 = 1;
    81: op1_01_inv27 = 1;
    84: op1_01_inv27 = 1;
    85: op1_01_inv27 = 1;
    86: op1_01_inv27 = 1;
    88: op1_01_inv27 = 1;
    89: op1_01_inv27 = 1;
    90: op1_01_inv27 = 1;
    95: op1_01_inv27 = 1;
    96: op1_01_inv27 = 1;
    default: op1_01_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in28 = reg_0330;
    7: op1_01_in28 = reg_0361;
    8: op1_01_in28 = imem07_in[75:72];
    9: op1_01_in28 = imem02_in[83:80];
    10: op1_01_in28 = reg_0370;
    11: op1_01_in28 = imem04_in[59:56];
    12: op1_01_in28 = reg_0766;
    13: op1_01_in28 = reg_0589;
    15: op1_01_in28 = reg_0318;
    16: op1_01_in28 = reg_0980;
    17: op1_01_in28 = reg_0406;
    18: op1_01_in28 = reg_0120;
    20: op1_01_in28 = imem01_in[99:96];
    21: op1_01_in28 = reg_0134;
    22: op1_01_in28 = reg_1015;
    23: op1_01_in28 = reg_0573;
    24: op1_01_in28 = reg_0437;
    25: op1_01_in28 = imem04_in[107:104];
    26: op1_01_in28 = reg_0633;
    27: op1_01_in28 = reg_0393;
    28: op1_01_in28 = reg_0405;
    29: op1_01_in28 = reg_0100;
    30: op1_01_in28 = imem03_in[15:12];
    31: op1_01_in28 = reg_0391;
    32: op1_01_in28 = reg_0238;
    33: op1_01_in28 = imem03_in[39:36];
    34: op1_01_in28 = imem04_in[39:36];
    35: op1_01_in28 = reg_0216;
    37: op1_01_in28 = reg_1043;
    38: op1_01_in28 = reg_1008;
    39: op1_01_in28 = imem03_in[31:28];
    40: op1_01_in28 = reg_0757;
    41: op1_01_in28 = reg_0912;
    43: op1_01_in28 = reg_0249;
    44: op1_01_in28 = imem03_in[55:52];
    47: op1_01_in28 = imem03_in[55:52];
    45: op1_01_in28 = reg_0148;
    46: op1_01_in28 = reg_0176;
    48: op1_01_in28 = reg_0530;
    51: op1_01_in28 = reg_0706;
    52: op1_01_in28 = imem05_in[91:88];
    53: op1_01_in28 = reg_0152;
    54: op1_01_in28 = imem06_in[127:124];
    55: op1_01_in28 = reg_0495;
    57: op1_01_in28 = reg_0928;
    58: op1_01_in28 = reg_1041;
    60: op1_01_in28 = reg_0662;
    61: op1_01_in28 = imem02_in[23:20];
    62: op1_01_in28 = reg_0535;
    63: op1_01_in28 = reg_0625;
    64: op1_01_in28 = reg_0744;
    69: op1_01_in28 = reg_0055;
    70: op1_01_in28 = reg_1028;
    71: op1_01_in28 = reg_0105;
    72: op1_01_in28 = reg_0297;
    75: op1_01_in28 = reg_1014;
    76: op1_01_in28 = reg_0551;
    77: op1_01_in28 = reg_0278;
    78: op1_01_in28 = imem06_in[91:88];
    81: op1_01_in28 = reg_1033;
    82: op1_01_in28 = reg_0227;
    83: op1_01_in28 = reg_0755;
    84: op1_01_in28 = reg_0064;
    85: op1_01_in28 = reg_0838;
    86: op1_01_in28 = reg_0232;
    87: op1_01_in28 = reg_0427;
    88: op1_01_in28 = reg_0923;
    89: op1_01_in28 = imem02_in[35:32];
    90: op1_01_in28 = reg_0002;
    93: op1_01_in28 = reg_0577;
    94: op1_01_in28 = reg_0147;
    95: op1_01_in28 = imem04_in[99:96];
    96: op1_01_in28 = imem04_in[63:60];
    97: op1_01_in28 = reg_0739;
    default: op1_01_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv28 = 1;
    7: op1_01_inv28 = 1;
    12: op1_01_inv28 = 1;
    13: op1_01_inv28 = 1;
    15: op1_01_inv28 = 1;
    17: op1_01_inv28 = 1;
    21: op1_01_inv28 = 1;
    22: op1_01_inv28 = 1;
    27: op1_01_inv28 = 1;
    29: op1_01_inv28 = 1;
    32: op1_01_inv28 = 1;
    33: op1_01_inv28 = 1;
    34: op1_01_inv28 = 1;
    35: op1_01_inv28 = 1;
    37: op1_01_inv28 = 1;
    39: op1_01_inv28 = 1;
    40: op1_01_inv28 = 1;
    41: op1_01_inv28 = 1;
    43: op1_01_inv28 = 1;
    47: op1_01_inv28 = 1;
    51: op1_01_inv28 = 1;
    55: op1_01_inv28 = 1;
    60: op1_01_inv28 = 1;
    63: op1_01_inv28 = 1;
    69: op1_01_inv28 = 1;
    70: op1_01_inv28 = 1;
    71: op1_01_inv28 = 1;
    72: op1_01_inv28 = 1;
    76: op1_01_inv28 = 1;
    78: op1_01_inv28 = 1;
    82: op1_01_inv28 = 1;
    83: op1_01_inv28 = 1;
    84: op1_01_inv28 = 1;
    85: op1_01_inv28 = 1;
    86: op1_01_inv28 = 1;
    87: op1_01_inv28 = 1;
    89: op1_01_inv28 = 1;
    90: op1_01_inv28 = 1;
    93: op1_01_inv28 = 1;
    94: op1_01_inv28 = 1;
    96: op1_01_inv28 = 1;
    default: op1_01_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in29 = reg_0342;
    7: op1_01_in29 = reg_0389;
    8: op1_01_in29 = reg_0728;
    9: op1_01_in29 = imem02_in[95:92];
    10: op1_01_in29 = reg_0343;
    11: op1_01_in29 = imem04_in[83:80];
    12: op1_01_in29 = reg_0237;
    13: op1_01_in29 = reg_0594;
    15: op1_01_in29 = reg_0310;
    16: op1_01_in29 = reg_0978;
    17: op1_01_in29 = reg_0367;
    18: op1_01_in29 = reg_0109;
    20: op1_01_in29 = reg_0496;
    21: op1_01_in29 = reg_0144;
    22: op1_01_in29 = reg_1041;
    23: op1_01_in29 = reg_0591;
    24: op1_01_in29 = reg_0162;
    25: op1_01_in29 = reg_0530;
    26: op1_01_in29 = reg_0618;
    27: op1_01_in29 = reg_0993;
    28: op1_01_in29 = reg_0403;
    29: op1_01_in29 = imem02_in[3:0];
    30: op1_01_in29 = imem03_in[27:24];
    31: op1_01_in29 = reg_0243;
    32: op1_01_in29 = reg_0226;
    33: op1_01_in29 = imem03_in[47:44];
    39: op1_01_in29 = imem03_in[47:44];
    34: op1_01_in29 = imem04_in[47:44];
    35: op1_01_in29 = reg_1035;
    37: op1_01_in29 = reg_0500;
    38: op1_01_in29 = reg_1019;
    63: op1_01_in29 = reg_1019;
    40: op1_01_in29 = reg_0152;
    41: op1_01_in29 = reg_0292;
    43: op1_01_in29 = reg_0522;
    44: op1_01_in29 = imem03_in[107:104];
    45: op1_01_in29 = reg_0145;
    47: op1_01_in29 = imem03_in[83:80];
    48: op1_01_in29 = reg_0055;
    51: op1_01_in29 = reg_0727;
    52: op1_01_in29 = imem05_in[99:96];
    53: op1_01_in29 = reg_0143;
    54: op1_01_in29 = reg_0614;
    55: op1_01_in29 = reg_0042;
    57: op1_01_in29 = reg_1045;
    58: op1_01_in29 = reg_0740;
    60: op1_01_in29 = reg_0923;
    61: op1_01_in29 = imem02_in[71:68];
    62: op1_01_in29 = reg_0572;
    64: op1_01_in29 = reg_0353;
    69: op1_01_in29 = reg_0931;
    70: op1_01_in29 = reg_0605;
    71: op1_01_in29 = reg_0122;
    72: op1_01_in29 = reg_0895;
    75: op1_01_in29 = reg_1023;
    76: op1_01_in29 = reg_0979;
    77: op1_01_in29 = reg_0038;
    78: op1_01_in29 = imem06_in[111:108];
    81: op1_01_in29 = reg_0115;
    82: op1_01_in29 = reg_0354;
    83: op1_01_in29 = reg_1010;
    84: op1_01_in29 = reg_0288;
    85: op1_01_in29 = reg_0161;
    86: op1_01_in29 = reg_1051;
    87: op1_01_in29 = reg_0868;
    88: op1_01_in29 = reg_0708;
    89: op1_01_in29 = imem02_in[115:112];
    90: op1_01_in29 = reg_0419;
    93: op1_01_in29 = reg_1009;
    94: op1_01_in29 = reg_0912;
    95: op1_01_in29 = imem04_in[119:116];
    96: op1_01_in29 = imem04_in[71:68];
    97: op1_01_in29 = reg_0441;
    default: op1_01_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_01_inv29 = 1;
    10: op1_01_inv29 = 1;
    13: op1_01_inv29 = 1;
    17: op1_01_inv29 = 1;
    18: op1_01_inv29 = 1;
    23: op1_01_inv29 = 1;
    26: op1_01_inv29 = 1;
    28: op1_01_inv29 = 1;
    31: op1_01_inv29 = 1;
    34: op1_01_inv29 = 1;
    35: op1_01_inv29 = 1;
    37: op1_01_inv29 = 1;
    38: op1_01_inv29 = 1;
    39: op1_01_inv29 = 1;
    41: op1_01_inv29 = 1;
    44: op1_01_inv29 = 1;
    51: op1_01_inv29 = 1;
    52: op1_01_inv29 = 1;
    53: op1_01_inv29 = 1;
    54: op1_01_inv29 = 1;
    55: op1_01_inv29 = 1;
    57: op1_01_inv29 = 1;
    58: op1_01_inv29 = 1;
    60: op1_01_inv29 = 1;
    61: op1_01_inv29 = 1;
    72: op1_01_inv29 = 1;
    75: op1_01_inv29 = 1;
    78: op1_01_inv29 = 1;
    84: op1_01_inv29 = 1;
    86: op1_01_inv29 = 1;
    87: op1_01_inv29 = 1;
    88: op1_01_inv29 = 1;
    90: op1_01_inv29 = 1;
    95: op1_01_inv29 = 1;
    97: op1_01_inv29 = 1;
    default: op1_01_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_01_in30 = reg_0083;
    7: op1_01_in30 = reg_0992;
    8: op1_01_in30 = reg_0719;
    9: op1_01_in30 = imem02_in[111:108];
    10: op1_01_in30 = reg_0385;
    11: op1_01_in30 = imem04_in[91:88];
    34: op1_01_in30 = imem04_in[91:88];
    96: op1_01_in30 = imem04_in[91:88];
    12: op1_01_in30 = reg_0234;
    71: op1_01_in30 = reg_0234;
    13: op1_01_in30 = reg_0581;
    15: op1_01_in30 = reg_0092;
    16: op1_01_in30 = reg_0989;
    76: op1_01_in30 = reg_0989;
    17: op1_01_in30 = reg_0800;
    18: op1_01_in30 = reg_0107;
    20: op1_01_in30 = reg_0119;
    21: op1_01_in30 = imem06_in[123:120];
    22: op1_01_in30 = reg_0124;
    23: op1_01_in30 = reg_0563;
    24: op1_01_in30 = reg_0158;
    25: op1_01_in30 = reg_0511;
    26: op1_01_in30 = reg_0623;
    27: op1_01_in30 = reg_0986;
    28: op1_01_in30 = reg_0406;
    29: op1_01_in30 = imem02_in[43:40];
    30: op1_01_in30 = imem03_in[47:44];
    31: op1_01_in30 = reg_0222;
    32: op1_01_in30 = reg_1032;
    33: op1_01_in30 = imem03_in[51:48];
    35: op1_01_in30 = reg_0904;
    37: op1_01_in30 = reg_1018;
    38: op1_01_in30 = reg_1049;
    39: op1_01_in30 = imem03_in[59:56];
    40: op1_01_in30 = reg_0129;
    41: op1_01_in30 = reg_0065;
    43: op1_01_in30 = reg_1017;
    82: op1_01_in30 = reg_1017;
    44: op1_01_in30 = reg_0327;
    45: op1_01_in30 = reg_0142;
    47: op1_01_in30 = imem03_in[99:96];
    48: op1_01_in30 = reg_0292;
    51: op1_01_in30 = reg_0426;
    52: op1_01_in30 = imem05_in[107:104];
    53: op1_01_in30 = reg_0153;
    54: op1_01_in30 = reg_0020;
    55: op1_01_in30 = reg_0393;
    57: op1_01_in30 = reg_0871;
    58: op1_01_in30 = reg_0925;
    60: op1_01_in30 = reg_0377;
    61: op1_01_in30 = imem02_in[95:92];
    62: op1_01_in30 = reg_1007;
    63: op1_01_in30 = reg_0244;
    64: op1_01_in30 = reg_0599;
    69: op1_01_in30 = reg_0541;
    70: op1_01_in30 = reg_0633;
    72: op1_01_in30 = reg_0595;
    75: op1_01_in30 = reg_1035;
    77: op1_01_in30 = reg_0773;
    78: op1_01_in30 = reg_0625;
    81: op1_01_in30 = imem02_in[51:48];
    83: op1_01_in30 = reg_0403;
    84: op1_01_in30 = reg_0041;
    85: op1_01_in30 = reg_0690;
    86: op1_01_in30 = reg_1033;
    87: op1_01_in30 = reg_0024;
    88: op1_01_in30 = reg_0299;
    89: op1_01_in30 = reg_0069;
    90: op1_01_in30 = reg_0532;
    93: op1_01_in30 = reg_0048;
    94: op1_01_in30 = reg_0306;
    95: op1_01_in30 = imem04_in[123:120];
    97: op1_01_in30 = reg_0039;
    default: op1_01_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_01_inv30 = 1;
    9: op1_01_inv30 = 1;
    10: op1_01_inv30 = 1;
    13: op1_01_inv30 = 1;
    15: op1_01_inv30 = 1;
    16: op1_01_inv30 = 1;
    20: op1_01_inv30 = 1;
    24: op1_01_inv30 = 1;
    26: op1_01_inv30 = 1;
    28: op1_01_inv30 = 1;
    29: op1_01_inv30 = 1;
    30: op1_01_inv30 = 1;
    33: op1_01_inv30 = 1;
    38: op1_01_inv30 = 1;
    43: op1_01_inv30 = 1;
    45: op1_01_inv30 = 1;
    51: op1_01_inv30 = 1;
    53: op1_01_inv30 = 1;
    57: op1_01_inv30 = 1;
    58: op1_01_inv30 = 1;
    61: op1_01_inv30 = 1;
    62: op1_01_inv30 = 1;
    64: op1_01_inv30 = 1;
    69: op1_01_inv30 = 1;
    70: op1_01_inv30 = 1;
    77: op1_01_inv30 = 1;
    81: op1_01_inv30 = 1;
    86: op1_01_inv30 = 1;
    90: op1_01_inv30 = 1;
    97: op1_01_inv30 = 1;
    default: op1_01_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_01_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in00 = reg_0042;
    6: op1_02_in00 = imem00_in[43:40];
    7: op1_02_in00 = reg_0993;
    8: op1_02_in00 = imem00_in[27:24];
    68: op1_02_in00 = imem00_in[27:24];
    9: op1_02_in00 = imem02_in[115:112];
    4: op1_02_in00 = imem07_in[75:72];
    10: op1_02_in00 = reg_0322;
    3: op1_02_in00 = imem07_in[43:40];
    11: op1_02_in00 = imem04_in[107:104];
    12: op1_02_in00 = reg_0487;
    13: op1_02_in00 = reg_0387;
    14: op1_02_in00 = imem00_in[15:12];
    73: op1_02_in00 = imem00_in[15:12];
    91: op1_02_in00 = imem00_in[15:12];
    15: op1_02_in00 = reg_0089;
    2: op1_02_in00 = imem07_in[23:20];
    16: op1_02_in00 = reg_0981;
    17: op1_02_in00 = reg_0486;
    18: op1_02_in00 = imem02_in[27:24];
    19: op1_02_in00 = imem00_in[3:0];
    56: op1_02_in00 = imem00_in[3:0];
    74: op1_02_in00 = imem00_in[3:0];
    90: op1_02_in00 = imem00_in[3:0];
    92: op1_02_in00 = imem00_in[3:0];
    20: op1_02_in00 = reg_0115;
    21: op1_02_in00 = reg_0628;
    22: op1_02_in00 = reg_0108;
    23: op1_02_in00 = reg_0585;
    24: op1_02_in00 = imem00_in[111:108];
    25: op1_02_in00 = reg_1020;
    26: op1_02_in00 = reg_0615;
    82: op1_02_in00 = reg_0615;
    27: op1_02_in00 = imem04_in[15:12];
    28: op1_02_in00 = reg_0787;
    29: op1_02_in00 = reg_0661;
    30: op1_02_in00 = imem03_in[119:116];
    31: op1_02_in00 = reg_1030;
    32: op1_02_in00 = reg_1037;
    33: op1_02_in00 = imem03_in[55:52];
    34: op1_02_in00 = imem04_in[115:112];
    35: op1_02_in00 = reg_0124;
    36: op1_02_in00 = imem00_in[87:84];
    37: op1_02_in00 = reg_0118;
    38: op1_02_in00 = reg_0581;
    39: op1_02_in00 = imem03_in[115:112];
    47: op1_02_in00 = imem03_in[115:112];
    40: op1_02_in00 = reg_0130;
    41: op1_02_in00 = reg_0075;
    42: op1_02_in00 = imem00_in[59:56];
    43: op1_02_in00 = reg_0925;
    44: op1_02_in00 = reg_0580;
    45: op1_02_in00 = reg_0146;
    46: op1_02_in00 = imem00_in[39:36];
    49: op1_02_in00 = imem00_in[39:36];
    48: op1_02_in00 = reg_0050;
    50: op1_02_in00 = imem00_in[7:4];
    66: op1_02_in00 = imem00_in[7:4];
    80: op1_02_in00 = imem00_in[7:4];
    51: op1_02_in00 = reg_0641;
    52: op1_02_in00 = reg_0962;
    53: op1_02_in00 = imem06_in[11:8];
    54: op1_02_in00 = reg_0371;
    55: op1_02_in00 = reg_0917;
    72: op1_02_in00 = reg_0917;
    57: op1_02_in00 = reg_1043;
    58: op1_02_in00 = reg_0832;
    59: op1_02_in00 = imem00_in[35:32];
    79: op1_02_in00 = imem00_in[35:32];
    60: op1_02_in00 = reg_0807;
    61: op1_02_in00 = imem02_in[99:96];
    62: op1_02_in00 = reg_0307;
    63: op1_02_in00 = reg_0021;
    64: op1_02_in00 = reg_0427;
    65: op1_02_in00 = imem00_in[19:16];
    67: op1_02_in00 = imem00_in[75:72];
    69: op1_02_in00 = reg_0752;
    70: op1_02_in00 = reg_0955;
    71: op1_02_in00 = reg_0793;
    75: op1_02_in00 = reg_1031;
    76: op1_02_in00 = reg_0990;
    77: op1_02_in00 = reg_0672;
    78: op1_02_in00 = reg_0694;
    81: op1_02_in00 = imem02_in[59:56];
    83: op1_02_in00 = reg_0369;
    84: op1_02_in00 = reg_0854;
    85: op1_02_in00 = imem00_in[31:28];
    86: op1_02_in00 = reg_0112;
    87: op1_02_in00 = reg_0429;
    88: op1_02_in00 = reg_0903;
    89: op1_02_in00 = reg_0639;
    93: op1_02_in00 = reg_1005;
    94: op1_02_in00 = reg_1005;
    95: op1_02_in00 = reg_0395;
    96: op1_02_in00 = imem04_in[123:120];
    97: op1_02_in00 = reg_0425;
    default: op1_02_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv00 = 1;
    6: op1_02_inv00 = 1;
    7: op1_02_inv00 = 1;
    9: op1_02_inv00 = 1;
    12: op1_02_inv00 = 1;
    14: op1_02_inv00 = 1;
    15: op1_02_inv00 = 1;
    16: op1_02_inv00 = 1;
    20: op1_02_inv00 = 1;
    21: op1_02_inv00 = 1;
    22: op1_02_inv00 = 1;
    23: op1_02_inv00 = 1;
    24: op1_02_inv00 = 1;
    25: op1_02_inv00 = 1;
    26: op1_02_inv00 = 1;
    28: op1_02_inv00 = 1;
    30: op1_02_inv00 = 1;
    33: op1_02_inv00 = 1;
    34: op1_02_inv00 = 1;
    37: op1_02_inv00 = 1;
    38: op1_02_inv00 = 1;
    40: op1_02_inv00 = 1;
    41: op1_02_inv00 = 1;
    44: op1_02_inv00 = 1;
    46: op1_02_inv00 = 1;
    50: op1_02_inv00 = 1;
    53: op1_02_inv00 = 1;
    54: op1_02_inv00 = 1;
    55: op1_02_inv00 = 1;
    57: op1_02_inv00 = 1;
    59: op1_02_inv00 = 1;
    60: op1_02_inv00 = 1;
    63: op1_02_inv00 = 1;
    64: op1_02_inv00 = 1;
    67: op1_02_inv00 = 1;
    69: op1_02_inv00 = 1;
    70: op1_02_inv00 = 1;
    71: op1_02_inv00 = 1;
    74: op1_02_inv00 = 1;
    77: op1_02_inv00 = 1;
    78: op1_02_inv00 = 1;
    79: op1_02_inv00 = 1;
    81: op1_02_inv00 = 1;
    82: op1_02_inv00 = 1;
    86: op1_02_inv00 = 1;
    87: op1_02_inv00 = 1;
    88: op1_02_inv00 = 1;
    90: op1_02_inv00 = 1;
    92: op1_02_inv00 = 1;
    94: op1_02_inv00 = 1;
    96: op1_02_inv00 = 1;
    97: op1_02_inv00 = 1;
    default: op1_02_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in01 = reg_0080;
    15: op1_02_in01 = reg_0080;
    6: op1_02_in01 = imem00_in[127:124];
    7: op1_02_in01 = reg_0980;
    8: op1_02_in01 = imem00_in[51:48];
    14: op1_02_in01 = imem00_in[51:48];
    49: op1_02_in01 = imem00_in[51:48];
    9: op1_02_in01 = imem02_in[119:116];
    4: op1_02_in01 = reg_0425;
    10: op1_02_in01 = reg_0398;
    3: op1_02_in01 = imem07_in[71:68];
    11: op1_02_in01 = imem04_in[119:116];
    12: op1_02_in01 = reg_1050;
    13: op1_02_in01 = reg_0391;
    2: op1_02_in01 = imem07_in[27:24];
    16: op1_02_in01 = imem04_in[7:4];
    17: op1_02_in01 = reg_0805;
    18: op1_02_in01 = imem02_in[87:84];
    81: op1_02_in01 = imem02_in[87:84];
    19: op1_02_in01 = imem00_in[23:20];
    50: op1_02_in01 = imem00_in[23:20];
    20: op1_02_in01 = reg_0127;
    21: op1_02_in01 = reg_0610;
    22: op1_02_in01 = reg_0126;
    23: op1_02_in01 = reg_0597;
    24: op1_02_in01 = imem00_in[119:116];
    25: op1_02_in01 = reg_1005;
    26: op1_02_in01 = reg_0381;
    27: op1_02_in01 = imem04_in[19:16];
    28: op1_02_in01 = reg_0027;
    29: op1_02_in01 = reg_0639;
    30: op1_02_in01 = imem03_in[123:120];
    39: op1_02_in01 = imem03_in[123:120];
    31: op1_02_in01 = reg_0803;
    32: op1_02_in01 = reg_0216;
    33: op1_02_in01 = imem03_in[59:56];
    34: op1_02_in01 = reg_0511;
    35: op1_02_in01 = reg_0107;
    36: op1_02_in01 = imem00_in[99:96];
    37: op1_02_in01 = reg_0112;
    38: op1_02_in01 = reg_0004;
    44: op1_02_in01 = reg_0004;
    40: op1_02_in01 = reg_0140;
    41: op1_02_in01 = reg_0047;
    42: op1_02_in01 = imem00_in[79:76];
    43: op1_02_in01 = reg_0099;
    45: op1_02_in01 = reg_0154;
    46: op1_02_in01 = imem00_in[63:60];
    59: op1_02_in01 = imem00_in[63:60];
    47: op1_02_in01 = reg_0394;
    48: op1_02_in01 = reg_0507;
    51: op1_02_in01 = reg_0420;
    52: op1_02_in01 = reg_0970;
    53: op1_02_in01 = imem06_in[47:44];
    54: op1_02_in01 = reg_0611;
    55: op1_02_in01 = reg_0241;
    56: op1_02_in01 = imem00_in[47:44];
    79: op1_02_in01 = imem00_in[47:44];
    90: op1_02_in01 = imem00_in[47:44];
    91: op1_02_in01 = imem00_in[47:44];
    57: op1_02_in01 = reg_0829;
    58: op1_02_in01 = reg_1055;
    75: op1_02_in01 = reg_1055;
    60: op1_02_in01 = reg_0836;
    61: op1_02_in01 = reg_0341;
    62: op1_02_in01 = reg_0434;
    63: op1_02_in01 = reg_0926;
    64: op1_02_in01 = reg_0024;
    65: op1_02_in01 = imem00_in[31:28];
    74: op1_02_in01 = imem00_in[31:28];
    66: op1_02_in01 = imem00_in[27:24];
    80: op1_02_in01 = imem00_in[27:24];
    67: op1_02_in01 = imem00_in[87:84];
    73: op1_02_in01 = imem00_in[87:84];
    68: op1_02_in01 = imem00_in[67:64];
    69: op1_02_in01 = reg_0014;
    70: op1_02_in01 = reg_0957;
    71: op1_02_in01 = reg_0604;
    72: op1_02_in01 = reg_0619;
    76: op1_02_in01 = reg_1000;
    77: op1_02_in01 = reg_0982;
    78: op1_02_in01 = reg_1019;
    82: op1_02_in01 = reg_1053;
    83: op1_02_in01 = reg_0022;
    84: op1_02_in01 = reg_0332;
    85: op1_02_in01 = imem00_in[59:56];
    86: op1_02_in01 = reg_0745;
    87: op1_02_in01 = reg_0181;
    88: op1_02_in01 = reg_0727;
    89: op1_02_in01 = reg_0091;
    92: op1_02_in01 = imem00_in[35:32];
    93: op1_02_in01 = reg_0888;
    94: op1_02_in01 = reg_0292;
    95: op1_02_in01 = reg_0550;
    96: op1_02_in01 = reg_0430;
    97: op1_02_in01 = reg_0775;
    default: op1_02_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_02_inv01 = 1;
    9: op1_02_inv01 = 1;
    4: op1_02_inv01 = 1;
    3: op1_02_inv01 = 1;
    11: op1_02_inv01 = 1;
    13: op1_02_inv01 = 1;
    19: op1_02_inv01 = 1;
    20: op1_02_inv01 = 1;
    27: op1_02_inv01 = 1;
    31: op1_02_inv01 = 1;
    32: op1_02_inv01 = 1;
    33: op1_02_inv01 = 1;
    35: op1_02_inv01 = 1;
    36: op1_02_inv01 = 1;
    38: op1_02_inv01 = 1;
    39: op1_02_inv01 = 1;
    42: op1_02_inv01 = 1;
    43: op1_02_inv01 = 1;
    44: op1_02_inv01 = 1;
    45: op1_02_inv01 = 1;
    46: op1_02_inv01 = 1;
    49: op1_02_inv01 = 1;
    50: op1_02_inv01 = 1;
    54: op1_02_inv01 = 1;
    56: op1_02_inv01 = 1;
    57: op1_02_inv01 = 1;
    59: op1_02_inv01 = 1;
    61: op1_02_inv01 = 1;
    63: op1_02_inv01 = 1;
    64: op1_02_inv01 = 1;
    66: op1_02_inv01 = 1;
    68: op1_02_inv01 = 1;
    69: op1_02_inv01 = 1;
    71: op1_02_inv01 = 1;
    72: op1_02_inv01 = 1;
    73: op1_02_inv01 = 1;
    74: op1_02_inv01 = 1;
    76: op1_02_inv01 = 1;
    80: op1_02_inv01 = 1;
    81: op1_02_inv01 = 1;
    82: op1_02_inv01 = 1;
    84: op1_02_inv01 = 1;
    89: op1_02_inv01 = 1;
    90: op1_02_inv01 = 1;
    93: op1_02_inv01 = 1;
    95: op1_02_inv01 = 1;
    default: op1_02_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in02 = imem03_in[7:4];
    6: op1_02_in02 = reg_0675;
    7: op1_02_in02 = reg_0978;
    8: op1_02_in02 = imem00_in[71:68];
    46: op1_02_in02 = imem00_in[71:68];
    65: op1_02_in02 = imem00_in[71:68];
    9: op1_02_in02 = reg_0649;
    4: op1_02_in02 = reg_0430;
    10: op1_02_in02 = reg_0312;
    3: op1_02_in02 = imem07_in[115:112];
    11: op1_02_in02 = imem04_in[127:124];
    12: op1_02_in02 = reg_0885;
    13: op1_02_in02 = reg_0370;
    14: op1_02_in02 = imem00_in[91:88];
    68: op1_02_in02 = imem00_in[91:88];
    15: op1_02_in02 = reg_0095;
    2: op1_02_in02 = imem07_in[87:84];
    16: op1_02_in02 = imem04_in[11:8];
    17: op1_02_in02 = reg_0782;
    31: op1_02_in02 = reg_0782;
    18: op1_02_in02 = imem02_in[99:96];
    19: op1_02_in02 = imem00_in[35:32];
    20: op1_02_in02 = imem02_in[43:40];
    35: op1_02_in02 = imem02_in[43:40];
    21: op1_02_in02 = reg_0629;
    22: op1_02_in02 = imem02_in[7:4];
    23: op1_02_in02 = reg_0581;
    24: op1_02_in02 = reg_0698;
    25: op1_02_in02 = reg_0778;
    26: op1_02_in02 = reg_0372;
    27: op1_02_in02 = imem04_in[51:48];
    28: op1_02_in02 = reg_0026;
    29: op1_02_in02 = reg_0647;
    30: op1_02_in02 = reg_0602;
    32: op1_02_in02 = reg_0913;
    33: op1_02_in02 = reg_0006;
    39: op1_02_in02 = reg_0006;
    34: op1_02_in02 = reg_0277;
    36: op1_02_in02 = imem00_in[103:100];
    42: op1_02_in02 = imem00_in[103:100];
    37: op1_02_in02 = reg_0106;
    38: op1_02_in02 = reg_0824;
    44: op1_02_in02 = reg_0824;
    40: op1_02_in02 = reg_0144;
    41: op1_02_in02 = reg_0751;
    43: op1_02_in02 = reg_0120;
    45: op1_02_in02 = reg_0140;
    47: op1_02_in02 = reg_0317;
    48: op1_02_in02 = reg_0524;
    49: op1_02_in02 = imem00_in[75:72];
    91: op1_02_in02 = imem00_in[75:72];
    50: op1_02_in02 = imem00_in[31:28];
    51: op1_02_in02 = reg_0502;
    52: op1_02_in02 = reg_0955;
    53: op1_02_in02 = imem06_in[67:64];
    54: op1_02_in02 = reg_0619;
    55: op1_02_in02 = reg_0605;
    56: op1_02_in02 = imem00_in[55:52];
    92: op1_02_in02 = imem00_in[55:52];
    57: op1_02_in02 = reg_0830;
    58: op1_02_in02 = reg_0111;
    59: op1_02_in02 = imem00_in[95:92];
    73: op1_02_in02 = imem00_in[95:92];
    60: op1_02_in02 = reg_0820;
    61: op1_02_in02 = reg_0565;
    62: op1_02_in02 = reg_0298;
    63: op1_02_in02 = reg_0384;
    64: op1_02_in02 = reg_0169;
    66: op1_02_in02 = imem00_in[39:36];
    67: op1_02_in02 = imem00_in[107:104];
    69: op1_02_in02 = reg_0276;
    70: op1_02_in02 = reg_0897;
    71: op1_02_in02 = reg_0520;
    72: op1_02_in02 = reg_0220;
    74: op1_02_in02 = imem00_in[59:56];
    79: op1_02_in02 = imem00_in[59:56];
    75: op1_02_in02 = reg_0116;
    76: op1_02_in02 = imem04_in[31:28];
    77: op1_02_in02 = reg_1001;
    78: op1_02_in02 = reg_0294;
    80: op1_02_in02 = imem00_in[63:60];
    81: op1_02_in02 = imem02_in[103:100];
    82: op1_02_in02 = reg_0273;
    83: op1_02_in02 = reg_0545;
    84: op1_02_in02 = imem05_in[7:4];
    85: op1_02_in02 = imem00_in[83:80];
    86: op1_02_in02 = imem02_in[31:28];
    87: op1_02_in02 = reg_0731;
    88: op1_02_in02 = reg_0250;
    89: op1_02_in02 = reg_0055;
    90: op1_02_in02 = imem00_in[115:112];
    93: op1_02_in02 = reg_0802;
    94: op1_02_in02 = reg_0540;
    95: op1_02_in02 = reg_0937;
    96: op1_02_in02 = reg_0123;
    97: op1_02_in02 = reg_0700;
    default: op1_02_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv02 = 1;
    6: op1_02_inv02 = 1;
    7: op1_02_inv02 = 1;
    8: op1_02_inv02 = 1;
    10: op1_02_inv02 = 1;
    3: op1_02_inv02 = 1;
    11: op1_02_inv02 = 1;
    14: op1_02_inv02 = 1;
    15: op1_02_inv02 = 1;
    2: op1_02_inv02 = 1;
    16: op1_02_inv02 = 1;
    18: op1_02_inv02 = 1;
    21: op1_02_inv02 = 1;
    27: op1_02_inv02 = 1;
    28: op1_02_inv02 = 1;
    29: op1_02_inv02 = 1;
    31: op1_02_inv02 = 1;
    32: op1_02_inv02 = 1;
    33: op1_02_inv02 = 1;
    34: op1_02_inv02 = 1;
    36: op1_02_inv02 = 1;
    37: op1_02_inv02 = 1;
    38: op1_02_inv02 = 1;
    40: op1_02_inv02 = 1;
    42: op1_02_inv02 = 1;
    43: op1_02_inv02 = 1;
    47: op1_02_inv02 = 1;
    50: op1_02_inv02 = 1;
    52: op1_02_inv02 = 1;
    53: op1_02_inv02 = 1;
    55: op1_02_inv02 = 1;
    56: op1_02_inv02 = 1;
    58: op1_02_inv02 = 1;
    59: op1_02_inv02 = 1;
    62: op1_02_inv02 = 1;
    63: op1_02_inv02 = 1;
    68: op1_02_inv02 = 1;
    72: op1_02_inv02 = 1;
    73: op1_02_inv02 = 1;
    74: op1_02_inv02 = 1;
    76: op1_02_inv02 = 1;
    77: op1_02_inv02 = 1;
    78: op1_02_inv02 = 1;
    79: op1_02_inv02 = 1;
    80: op1_02_inv02 = 1;
    81: op1_02_inv02 = 1;
    83: op1_02_inv02 = 1;
    89: op1_02_inv02 = 1;
    90: op1_02_inv02 = 1;
    91: op1_02_inv02 = 1;
    92: op1_02_inv02 = 1;
    94: op1_02_inv02 = 1;
    95: op1_02_inv02 = 1;
    97: op1_02_inv02 = 1;
    default: op1_02_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in03 = imem03_in[39:36];
    6: op1_02_in03 = reg_0680;
    7: op1_02_in03 = reg_0994;
    8: op1_02_in03 = imem00_in[79:76];
    80: op1_02_in03 = imem00_in[79:76];
    9: op1_02_in03 = reg_0320;
    4: op1_02_in03 = reg_0431;
    10: op1_02_in03 = reg_0361;
    3: op1_02_in03 = imem07_in[119:116];
    11: op1_02_in03 = reg_0545;
    12: op1_02_in03 = reg_0830;
    13: op1_02_in03 = reg_0388;
    14: op1_02_in03 = imem00_in[111:108];
    42: op1_02_in03 = imem00_in[111:108];
    85: op1_02_in03 = imem00_in[111:108];
    15: op1_02_in03 = reg_0090;
    2: op1_02_in03 = imem07_in[91:88];
    16: op1_02_in03 = imem04_in[51:48];
    17: op1_02_in03 = imem07_in[71:68];
    18: op1_02_in03 = imem02_in[103:100];
    19: op1_02_in03 = imem00_in[39:36];
    20: op1_02_in03 = imem02_in[47:44];
    21: op1_02_in03 = reg_0607;
    22: op1_02_in03 = imem02_in[67:64];
    23: op1_02_in03 = reg_0391;
    24: op1_02_in03 = reg_0688;
    25: op1_02_in03 = reg_0050;
    26: op1_02_in03 = reg_0408;
    27: op1_02_in03 = imem04_in[127:124];
    28: op1_02_in03 = reg_0808;
    29: op1_02_in03 = reg_0636;
    30: op1_02_in03 = reg_0586;
    94: op1_02_in03 = reg_0586;
    31: op1_02_in03 = imem07_in[47:44];
    32: op1_02_in03 = reg_1036;
    33: op1_02_in03 = reg_0571;
    34: op1_02_in03 = reg_0541;
    35: op1_02_in03 = imem02_in[55:52];
    36: op1_02_in03 = reg_0681;
    37: op1_02_in03 = reg_0110;
    38: op1_02_in03 = reg_0823;
    39: op1_02_in03 = reg_0938;
    40: op1_02_in03 = imem06_in[63:60];
    41: op1_02_in03 = reg_0774;
    43: op1_02_in03 = imem02_in[7:4];
    44: op1_02_in03 = reg_0923;
    45: op1_02_in03 = imem06_in[43:40];
    46: op1_02_in03 = imem00_in[83:80];
    65: op1_02_in03 = imem00_in[83:80];
    47: op1_02_in03 = reg_0327;
    48: op1_02_in03 = reg_0584;
    49: op1_02_in03 = imem00_in[87:84];
    50: op1_02_in03 = imem00_in[35:32];
    51: op1_02_in03 = reg_0174;
    52: op1_02_in03 = reg_0969;
    53: op1_02_in03 = imem06_in[95:92];
    54: op1_02_in03 = reg_0754;
    55: op1_02_in03 = reg_0025;
    56: op1_02_in03 = imem00_in[91:88];
    57: op1_02_in03 = reg_0216;
    58: op1_02_in03 = reg_0821;
    59: op1_02_in03 = imem00_in[107:104];
    60: op1_02_in03 = reg_0374;
    61: op1_02_in03 = reg_0648;
    62: op1_02_in03 = reg_0346;
    63: op1_02_in03 = reg_0440;
    64: op1_02_in03 = reg_0182;
    66: op1_02_in03 = imem00_in[47:44];
    67: op1_02_in03 = imem00_in[127:124];
    68: op1_02_in03 = imem00_in[103:100];
    69: op1_02_in03 = reg_0072;
    70: op1_02_in03 = imem07_in[7:4];
    71: op1_02_in03 = reg_0829;
    72: op1_02_in03 = reg_0485;
    73: op1_02_in03 = imem00_in[99:96];
    74: op1_02_in03 = imem00_in[75:72];
    75: op1_02_in03 = reg_0101;
    76: op1_02_in03 = reg_0511;
    77: op1_02_in03 = reg_0993;
    78: op1_02_in03 = reg_0351;
    79: op1_02_in03 = imem00_in[63:60];
    81: op1_02_in03 = reg_0810;
    82: op1_02_in03 = reg_0745;
    83: op1_02_in03 = reg_0573;
    84: op1_02_in03 = imem05_in[71:68];
    86: op1_02_in03 = imem02_in[63:60];
    87: op1_02_in03 = reg_0703;
    88: op1_02_in03 = reg_0421;
    89: op1_02_in03 = reg_0621;
    90: op1_02_in03 = reg_0841;
    91: op1_02_in03 = imem00_in[95:92];
    92: op1_02_in03 = imem00_in[59:56];
    93: op1_02_in03 = reg_0058;
    95: op1_02_in03 = reg_0888;
    96: op1_02_in03 = reg_0014;
    97: op1_02_in03 = reg_0778;
    default: op1_02_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_02_inv03 = 1;
    9: op1_02_inv03 = 1;
    10: op1_02_inv03 = 1;
    11: op1_02_inv03 = 1;
    12: op1_02_inv03 = 1;
    13: op1_02_inv03 = 1;
    15: op1_02_inv03 = 1;
    17: op1_02_inv03 = 1;
    19: op1_02_inv03 = 1;
    20: op1_02_inv03 = 1;
    21: op1_02_inv03 = 1;
    22: op1_02_inv03 = 1;
    26: op1_02_inv03 = 1;
    27: op1_02_inv03 = 1;
    28: op1_02_inv03 = 1;
    30: op1_02_inv03 = 1;
    32: op1_02_inv03 = 1;
    36: op1_02_inv03 = 1;
    37: op1_02_inv03 = 1;
    38: op1_02_inv03 = 1;
    40: op1_02_inv03 = 1;
    43: op1_02_inv03 = 1;
    44: op1_02_inv03 = 1;
    48: op1_02_inv03 = 1;
    51: op1_02_inv03 = 1;
    55: op1_02_inv03 = 1;
    59: op1_02_inv03 = 1;
    60: op1_02_inv03 = 1;
    61: op1_02_inv03 = 1;
    63: op1_02_inv03 = 1;
    64: op1_02_inv03 = 1;
    65: op1_02_inv03 = 1;
    66: op1_02_inv03 = 1;
    68: op1_02_inv03 = 1;
    75: op1_02_inv03 = 1;
    76: op1_02_inv03 = 1;
    79: op1_02_inv03 = 1;
    82: op1_02_inv03 = 1;
    84: op1_02_inv03 = 1;
    87: op1_02_inv03 = 1;
    88: op1_02_inv03 = 1;
    91: op1_02_inv03 = 1;
    92: op1_02_inv03 = 1;
    93: op1_02_inv03 = 1;
    96: op1_02_inv03 = 1;
    default: op1_02_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in04 = imem03_in[43:40];
    6: op1_02_in04 = reg_0692;
    7: op1_02_in04 = imem04_in[123:120];
    8: op1_02_in04 = imem00_in[83:80];
    92: op1_02_in04 = imem00_in[83:80];
    9: op1_02_in04 = reg_0318;
    4: op1_02_in04 = reg_0184;
    10: op1_02_in04 = reg_0396;
    3: op1_02_in04 = reg_0175;
    51: op1_02_in04 = reg_0175;
    11: op1_02_in04 = reg_0550;
    12: op1_02_in04 = reg_0216;
    13: op1_02_in04 = reg_0362;
    14: op1_02_in04 = reg_0695;
    15: op1_02_in04 = reg_0087;
    2: op1_02_in04 = imem07_in[103:100];
    16: op1_02_in04 = imem04_in[67:64];
    17: op1_02_in04 = imem07_in[115:112];
    18: op1_02_in04 = imem02_in[119:116];
    19: op1_02_in04 = imem00_in[43:40];
    20: op1_02_in04 = reg_0658;
    21: op1_02_in04 = reg_0605;
    22: op1_02_in04 = imem02_in[83:80];
    23: op1_02_in04 = reg_0321;
    88: op1_02_in04 = reg_0321;
    24: op1_02_in04 = reg_0463;
    25: op1_02_in04 = reg_0061;
    26: op1_02_in04 = reg_0405;
    27: op1_02_in04 = reg_0265;
    28: op1_02_in04 = reg_0018;
    29: op1_02_in04 = reg_0663;
    30: op1_02_in04 = reg_0599;
    31: op1_02_in04 = imem07_in[67:64];
    32: op1_02_in04 = reg_0228;
    33: op1_02_in04 = reg_1019;
    34: op1_02_in04 = reg_0537;
    35: op1_02_in04 = imem02_in[59:56];
    36: op1_02_in04 = reg_0676;
    37: op1_02_in04 = imem02_in[11:8];
    38: op1_02_in04 = reg_0038;
    39: op1_02_in04 = reg_0923;
    40: op1_02_in04 = imem06_in[71:68];
    41: op1_02_in04 = reg_0773;
    42: op1_02_in04 = reg_0682;
    43: op1_02_in04 = imem02_in[23:20];
    44: op1_02_in04 = reg_0807;
    45: op1_02_in04 = imem06_in[47:44];
    46: op1_02_in04 = imem00_in[99:96];
    47: op1_02_in04 = reg_0580;
    48: op1_02_in04 = reg_0401;
    96: op1_02_in04 = reg_0401;
    49: op1_02_in04 = imem00_in[95:92];
    74: op1_02_in04 = imem00_in[95:92];
    50: op1_02_in04 = imem00_in[51:48];
    52: op1_02_in04 = reg_0947;
    53: op1_02_in04 = imem06_in[123:120];
    54: op1_02_in04 = reg_0612;
    55: op1_02_in04 = reg_0626;
    56: op1_02_in04 = reg_0519;
    57: op1_02_in04 = reg_0902;
    58: op1_02_in04 = imem02_in[43:40];
    59: op1_02_in04 = imem00_in[119:116];
    60: op1_02_in04 = reg_0991;
    61: op1_02_in04 = reg_0636;
    62: op1_02_in04 = reg_0661;
    63: op1_02_in04 = reg_0617;
    64: op1_02_in04 = reg_0164;
    65: op1_02_in04 = imem00_in[91:88];
    66: op1_02_in04 = imem00_in[71:68];
    67: op1_02_in04 = reg_0001;
    68: op1_02_in04 = imem00_in[107:104];
    69: op1_02_in04 = reg_0495;
    70: op1_02_in04 = imem07_in[19:16];
    71: op1_02_in04 = reg_1037;
    72: op1_02_in04 = imem07_in[11:8];
    73: op1_02_in04 = reg_0670;
    75: op1_02_in04 = reg_0821;
    76: op1_02_in04 = reg_1005;
    77: op1_02_in04 = reg_0980;
    78: op1_02_in04 = reg_0267;
    79: op1_02_in04 = imem00_in[75:72];
    80: op1_02_in04 = reg_0768;
    81: op1_02_in04 = reg_0637;
    82: op1_02_in04 = imem02_in[63:60];
    83: op1_02_in04 = imem07_in[7:4];
    84: op1_02_in04 = imem05_in[75:72];
    85: op1_02_in04 = imem00_in[115:112];
    86: op1_02_in04 = imem02_in[87:84];
    87: op1_02_in04 = reg_0447;
    89: op1_02_in04 = reg_0077;
    90: op1_02_in04 = reg_0685;
    91: op1_02_in04 = imem00_in[103:100];
    93: op1_02_in04 = reg_0302;
    94: op1_02_in04 = reg_0802;
    95: op1_02_in04 = reg_0864;
    97: op1_02_in04 = reg_0086;
    default: op1_02_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv04 = 1;
    4: op1_02_inv04 = 1;
    11: op1_02_inv04 = 1;
    12: op1_02_inv04 = 1;
    13: op1_02_inv04 = 1;
    2: op1_02_inv04 = 1;
    16: op1_02_inv04 = 1;
    17: op1_02_inv04 = 1;
    21: op1_02_inv04 = 1;
    22: op1_02_inv04 = 1;
    26: op1_02_inv04 = 1;
    28: op1_02_inv04 = 1;
    31: op1_02_inv04 = 1;
    32: op1_02_inv04 = 1;
    33: op1_02_inv04 = 1;
    37: op1_02_inv04 = 1;
    38: op1_02_inv04 = 1;
    40: op1_02_inv04 = 1;
    42: op1_02_inv04 = 1;
    43: op1_02_inv04 = 1;
    45: op1_02_inv04 = 1;
    46: op1_02_inv04 = 1;
    47: op1_02_inv04 = 1;
    48: op1_02_inv04 = 1;
    49: op1_02_inv04 = 1;
    52: op1_02_inv04 = 1;
    53: op1_02_inv04 = 1;
    55: op1_02_inv04 = 1;
    56: op1_02_inv04 = 1;
    60: op1_02_inv04 = 1;
    62: op1_02_inv04 = 1;
    64: op1_02_inv04 = 1;
    65: op1_02_inv04 = 1;
    68: op1_02_inv04 = 1;
    69: op1_02_inv04 = 1;
    72: op1_02_inv04 = 1;
    73: op1_02_inv04 = 1;
    74: op1_02_inv04 = 1;
    75: op1_02_inv04 = 1;
    83: op1_02_inv04 = 1;
    85: op1_02_inv04 = 1;
    86: op1_02_inv04 = 1;
    87: op1_02_inv04 = 1;
    89: op1_02_inv04 = 1;
    92: op1_02_inv04 = 1;
    94: op1_02_inv04 = 1;
    95: op1_02_inv04 = 1;
    96: op1_02_inv04 = 1;
    default: op1_02_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in05 = imem03_in[79:76];
    6: op1_02_in05 = reg_0453;
    24: op1_02_in05 = reg_0453;
    7: op1_02_in05 = reg_0529;
    8: op1_02_in05 = imem00_in[107:104];
    9: op1_02_in05 = reg_0338;
    10: op1_02_in05 = reg_0309;
    3: op1_02_in05 = reg_0183;
    87: op1_02_in05 = reg_0183;
    11: op1_02_in05 = reg_0546;
    12: op1_02_in05 = reg_1041;
    13: op1_02_in05 = reg_0369;
    14: op1_02_in05 = reg_0688;
    15: op1_02_in05 = reg_0093;
    16: op1_02_in05 = reg_0560;
    17: op1_02_in05 = reg_0731;
    18: op1_02_in05 = reg_0661;
    20: op1_02_in05 = reg_0661;
    19: op1_02_in05 = imem00_in[71:68];
    21: op1_02_in05 = reg_0609;
    22: op1_02_in05 = imem02_in[95:92];
    23: op1_02_in05 = reg_0396;
    25: op1_02_in05 = reg_0733;
    26: op1_02_in05 = reg_0371;
    27: op1_02_in05 = reg_1009;
    28: op1_02_in05 = reg_1010;
    29: op1_02_in05 = reg_0334;
    30: op1_02_in05 = reg_0587;
    31: op1_02_in05 = imem07_in[71:68];
    32: op1_02_in05 = reg_1038;
    33: op1_02_in05 = reg_1049;
    34: op1_02_in05 = reg_0313;
    35: op1_02_in05 = imem02_in[99:96];
    36: op1_02_in05 = reg_0698;
    37: op1_02_in05 = imem02_in[23:20];
    38: op1_02_in05 = reg_0051;
    39: op1_02_in05 = reg_0795;
    40: op1_02_in05 = imem06_in[79:76];
    41: op1_02_in05 = reg_0044;
    42: op1_02_in05 = reg_0693;
    46: op1_02_in05 = reg_0693;
    43: op1_02_in05 = imem02_in[31:28];
    44: op1_02_in05 = reg_0767;
    45: op1_02_in05 = imem06_in[67:64];
    47: op1_02_in05 = reg_0397;
    48: op1_02_in05 = reg_0054;
    49: op1_02_in05 = reg_0683;
    50: op1_02_in05 = imem00_in[63:60];
    51: op1_02_in05 = reg_0165;
    52: op1_02_in05 = reg_0063;
    53: op1_02_in05 = reg_0915;
    54: op1_02_in05 = reg_0295;
    55: op1_02_in05 = reg_0263;
    56: op1_02_in05 = reg_0523;
    57: op1_02_in05 = reg_0111;
    58: op1_02_in05 = imem02_in[51:48];
    59: op1_02_in05 = reg_0768;
    60: op1_02_in05 = reg_0996;
    61: op1_02_in05 = reg_0424;
    62: op1_02_in05 = reg_0662;
    63: op1_02_in05 = reg_0595;
    64: op1_02_in05 = reg_0168;
    65: op1_02_in05 = imem00_in[103:100];
    66: op1_02_in05 = imem00_in[119:116];
    67: op1_02_in05 = reg_0671;
    68: op1_02_in05 = imem00_in[115:112];
    69: op1_02_in05 = imem05_in[15:12];
    70: op1_02_in05 = imem07_in[31:28];
    71: op1_02_in05 = reg_1040;
    72: op1_02_in05 = imem07_in[35:32];
    73: op1_02_in05 = reg_0738;
    74: op1_02_in05 = reg_0001;
    75: op1_02_in05 = reg_0110;
    76: op1_02_in05 = reg_0537;
    77: op1_02_in05 = reg_0994;
    78: op1_02_in05 = reg_0262;
    79: op1_02_in05 = reg_0843;
    90: op1_02_in05 = reg_0843;
    80: op1_02_in05 = reg_0825;
    81: op1_02_in05 = reg_0896;
    82: op1_02_in05 = reg_0650;
    83: op1_02_in05 = imem07_in[15:12];
    84: op1_02_in05 = imem05_in[83:80];
    85: op1_02_in05 = reg_0455;
    86: op1_02_in05 = imem02_in[107:104];
    88: op1_02_in05 = reg_0315;
    89: op1_02_in05 = reg_0644;
    91: op1_02_in05 = reg_0463;
    92: op1_02_in05 = imem00_in[99:96];
    93: op1_02_in05 = reg_0251;
    94: op1_02_in05 = reg_0067;
    95: op1_02_in05 = reg_0586;
    96: op1_02_in05 = reg_0815;
    97: op1_02_in05 = reg_0885;
    default: op1_02_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv05 = 1;
    8: op1_02_inv05 = 1;
    9: op1_02_inv05 = 1;
    3: op1_02_inv05 = 1;
    14: op1_02_inv05 = 1;
    16: op1_02_inv05 = 1;
    21: op1_02_inv05 = 1;
    23: op1_02_inv05 = 1;
    25: op1_02_inv05 = 1;
    27: op1_02_inv05 = 1;
    29: op1_02_inv05 = 1;
    32: op1_02_inv05 = 1;
    37: op1_02_inv05 = 1;
    40: op1_02_inv05 = 1;
    42: op1_02_inv05 = 1;
    44: op1_02_inv05 = 1;
    45: op1_02_inv05 = 1;
    51: op1_02_inv05 = 1;
    54: op1_02_inv05 = 1;
    55: op1_02_inv05 = 1;
    56: op1_02_inv05 = 1;
    58: op1_02_inv05 = 1;
    61: op1_02_inv05 = 1;
    62: op1_02_inv05 = 1;
    63: op1_02_inv05 = 1;
    64: op1_02_inv05 = 1;
    65: op1_02_inv05 = 1;
    68: op1_02_inv05 = 1;
    70: op1_02_inv05 = 1;
    71: op1_02_inv05 = 1;
    72: op1_02_inv05 = 1;
    74: op1_02_inv05 = 1;
    75: op1_02_inv05 = 1;
    76: op1_02_inv05 = 1;
    77: op1_02_inv05 = 1;
    79: op1_02_inv05 = 1;
    83: op1_02_inv05 = 1;
    84: op1_02_inv05 = 1;
    85: op1_02_inv05 = 1;
    86: op1_02_inv05 = 1;
    88: op1_02_inv05 = 1;
    92: op1_02_inv05 = 1;
    96: op1_02_inv05 = 1;
    default: op1_02_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in06 = imem03_in[99:96];
    6: op1_02_in06 = reg_0461;
    7: op1_02_in06 = reg_0539;
    8: op1_02_in06 = reg_0672;
    9: op1_02_in06 = reg_0335;
    89: op1_02_in06 = reg_0335;
    10: op1_02_in06 = reg_0985;
    3: op1_02_in06 = reg_0177;
    11: op1_02_in06 = reg_0531;
    12: op1_02_in06 = reg_1038;
    13: op1_02_in06 = reg_0322;
    14: op1_02_in06 = reg_0687;
    15: op1_02_in06 = reg_0073;
    16: op1_02_in06 = reg_0535;
    17: op1_02_in06 = reg_0721;
    18: op1_02_in06 = reg_0638;
    19: op1_02_in06 = imem00_in[83:80];
    20: op1_02_in06 = reg_0663;
    21: op1_02_in06 = reg_0619;
    22: op1_02_in06 = imem02_in[107:104];
    23: op1_02_in06 = reg_1002;
    24: op1_02_in06 = reg_0457;
    25: op1_02_in06 = reg_0276;
    26: op1_02_in06 = reg_0367;
    27: op1_02_in06 = reg_0066;
    28: op1_02_in06 = reg_0805;
    29: op1_02_in06 = reg_0045;
    30: op1_02_in06 = reg_0592;
    31: op1_02_in06 = imem07_in[91:88];
    32: op1_02_in06 = reg_0104;
    33: op1_02_in06 = reg_0581;
    34: op1_02_in06 = reg_0764;
    35: op1_02_in06 = imem02_in[111:108];
    36: op1_02_in06 = reg_0690;
    37: op1_02_in06 = imem02_in[35:32];
    38: op1_02_in06 = reg_0377;
    39: op1_02_in06 = reg_0784;
    40: op1_02_in06 = imem06_in[91:88];
    41: op1_02_in06 = reg_0021;
    42: op1_02_in06 = reg_0683;
    43: op1_02_in06 = imem02_in[43:40];
    44: op1_02_in06 = reg_0844;
    45: op1_02_in06 = imem06_in[71:68];
    46: op1_02_in06 = reg_0676;
    47: op1_02_in06 = reg_0923;
    48: op1_02_in06 = reg_0057;
    49: op1_02_in06 = reg_0681;
    50: op1_02_in06 = imem00_in[71:68];
    51: op1_02_in06 = reg_0162;
    52: op1_02_in06 = reg_0259;
    53: op1_02_in06 = reg_0759;
    54: op1_02_in06 = reg_0917;
    55: op1_02_in06 = imem07_in[11:8];
    56: op1_02_in06 = reg_0670;
    57: op1_02_in06 = reg_1053;
    58: op1_02_in06 = imem02_in[71:68];
    59: op1_02_in06 = reg_0686;
    60: op1_02_in06 = reg_0999;
    61: op1_02_in06 = reg_0052;
    62: op1_02_in06 = reg_0765;
    63: op1_02_in06 = reg_0380;
    65: op1_02_in06 = imem00_in[111:108];
    66: op1_02_in06 = reg_0841;
    74: op1_02_in06 = reg_0841;
    67: op1_02_in06 = reg_0843;
    68: op1_02_in06 = reg_0001;
    69: op1_02_in06 = imem05_in[27:24];
    70: op1_02_in06 = imem07_in[35:32];
    71: op1_02_in06 = reg_1031;
    72: op1_02_in06 = imem07_in[39:36];
    73: op1_02_in06 = reg_0668;
    75: op1_02_in06 = imem02_in[59:56];
    76: op1_02_in06 = reg_0524;
    77: op1_02_in06 = imem04_in[3:0];
    78: op1_02_in06 = reg_0626;
    79: op1_02_in06 = reg_0523;
    80: op1_02_in06 = reg_0523;
    81: op1_02_in06 = reg_0885;
    82: op1_02_in06 = reg_0916;
    83: op1_02_in06 = imem07_in[59:56];
    84: op1_02_in06 = imem05_in[107:104];
    85: op1_02_in06 = reg_0466;
    86: op1_02_in06 = reg_0277;
    87: op1_02_in06 = reg_0157;
    88: op1_02_in06 = reg_0175;
    90: op1_02_in06 = reg_0842;
    91: op1_02_in06 = reg_0465;
    92: op1_02_in06 = imem00_in[103:100];
    93: op1_02_in06 = reg_0070;
    94: op1_02_in06 = reg_0302;
    95: op1_02_in06 = reg_0016;
    96: op1_02_in06 = reg_0074;
    97: op1_02_in06 = reg_0365;
    default: op1_02_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv06 = 1;
    8: op1_02_inv06 = 1;
    9: op1_02_inv06 = 1;
    12: op1_02_inv06 = 1;
    17: op1_02_inv06 = 1;
    18: op1_02_inv06 = 1;
    22: op1_02_inv06 = 1;
    23: op1_02_inv06 = 1;
    25: op1_02_inv06 = 1;
    34: op1_02_inv06 = 1;
    35: op1_02_inv06 = 1;
    36: op1_02_inv06 = 1;
    37: op1_02_inv06 = 1;
    38: op1_02_inv06 = 1;
    39: op1_02_inv06 = 1;
    42: op1_02_inv06 = 1;
    43: op1_02_inv06 = 1;
    44: op1_02_inv06 = 1;
    45: op1_02_inv06 = 1;
    46: op1_02_inv06 = 1;
    49: op1_02_inv06 = 1;
    51: op1_02_inv06 = 1;
    52: op1_02_inv06 = 1;
    53: op1_02_inv06 = 1;
    59: op1_02_inv06 = 1;
    61: op1_02_inv06 = 1;
    62: op1_02_inv06 = 1;
    66: op1_02_inv06 = 1;
    68: op1_02_inv06 = 1;
    69: op1_02_inv06 = 1;
    73: op1_02_inv06 = 1;
    74: op1_02_inv06 = 1;
    75: op1_02_inv06 = 1;
    77: op1_02_inv06 = 1;
    80: op1_02_inv06 = 1;
    81: op1_02_inv06 = 1;
    83: op1_02_inv06 = 1;
    84: op1_02_inv06 = 1;
    86: op1_02_inv06 = 1;
    88: op1_02_inv06 = 1;
    89: op1_02_inv06 = 1;
    91: op1_02_inv06 = 1;
    92: op1_02_inv06 = 1;
    96: op1_02_inv06 = 1;
    default: op1_02_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in07 = reg_0582;
    6: op1_02_in07 = reg_0469;
    7: op1_02_in07 = reg_0537;
    95: op1_02_in07 = reg_0537;
    8: op1_02_in07 = reg_0679;
    9: op1_02_in07 = reg_0314;
    10: op1_02_in07 = reg_0998;
    3: op1_02_in07 = reg_0164;
    11: op1_02_in07 = reg_0556;
    12: op1_02_in07 = reg_0118;
    13: op1_02_in07 = reg_0397;
    14: op1_02_in07 = reg_0669;
    15: op1_02_in07 = imem03_in[11:8];
    16: op1_02_in07 = reg_0532;
    17: op1_02_in07 = reg_0714;
    18: op1_02_in07 = reg_0665;
    19: op1_02_in07 = imem00_in[87:84];
    50: op1_02_in07 = imem00_in[87:84];
    20: op1_02_in07 = reg_0352;
    21: op1_02_in07 = reg_0612;
    22: op1_02_in07 = reg_0334;
    23: op1_02_in07 = reg_1001;
    24: op1_02_in07 = reg_0189;
    25: op1_02_in07 = reg_0069;
    26: op1_02_in07 = reg_1029;
    27: op1_02_in07 = reg_0072;
    94: op1_02_in07 = reg_0072;
    28: op1_02_in07 = reg_0005;
    29: op1_02_in07 = reg_0842;
    66: op1_02_in07 = reg_0842;
    30: op1_02_in07 = reg_0594;
    31: op1_02_in07 = imem07_in[95:92];
    32: op1_02_in07 = reg_0119;
    33: op1_02_in07 = reg_0389;
    34: op1_02_in07 = reg_0740;
    35: op1_02_in07 = reg_0642;
    36: op1_02_in07 = reg_0699;
    37: op1_02_in07 = reg_0653;
    38: op1_02_in07 = reg_0807;
    39: op1_02_in07 = reg_0374;
    40: op1_02_in07 = imem06_in[107:104];
    41: op1_02_in07 = imem05_in[123:120];
    42: op1_02_in07 = reg_0696;
    43: op1_02_in07 = imem02_in[55:52];
    44: op1_02_in07 = reg_0822;
    45: op1_02_in07 = imem06_in[79:76];
    46: op1_02_in07 = reg_0698;
    47: op1_02_in07 = reg_0793;
    48: op1_02_in07 = reg_0286;
    49: op1_02_in07 = reg_0672;
    51: op1_02_in07 = reg_0167;
    52: op1_02_in07 = reg_0774;
    53: op1_02_in07 = reg_0624;
    54: op1_02_in07 = reg_0630;
    55: op1_02_in07 = imem07_in[31:28];
    56: op1_02_in07 = reg_0455;
    57: op1_02_in07 = reg_0110;
    58: op1_02_in07 = imem02_in[79:76];
    59: op1_02_in07 = reg_0668;
    60: op1_02_in07 = reg_0977;
    61: op1_02_in07 = reg_0423;
    62: op1_02_in07 = reg_0373;
    63: op1_02_in07 = reg_0348;
    65: op1_02_in07 = reg_0768;
    67: op1_02_in07 = reg_0686;
    68: op1_02_in07 = reg_0102;
    80: op1_02_in07 = reg_0102;
    69: op1_02_in07 = imem05_in[31:28];
    70: op1_02_in07 = imem07_in[83:80];
    71: op1_02_in07 = reg_1041;
    72: op1_02_in07 = imem07_in[47:44];
    73: op1_02_in07 = reg_0463;
    74: op1_02_in07 = reg_0671;
    75: op1_02_in07 = imem02_in[67:64];
    76: op1_02_in07 = reg_0014;
    77: op1_02_in07 = imem04_in[31:28];
    78: op1_02_in07 = reg_0328;
    79: op1_02_in07 = reg_0748;
    81: op1_02_in07 = reg_0907;
    82: op1_02_in07 = reg_0700;
    83: op1_02_in07 = imem07_in[87:84];
    84: op1_02_in07 = imem05_in[127:124];
    85: op1_02_in07 = reg_0475;
    86: op1_02_in07 = reg_0349;
    87: op1_02_in07 = reg_0371;
    88: op1_02_in07 = reg_0179;
    89: op1_02_in07 = reg_0381;
    90: op1_02_in07 = reg_0674;
    91: op1_02_in07 = reg_0454;
    92: op1_02_in07 = imem00_in[127:124];
    93: op1_02_in07 = reg_0856;
    96: op1_02_in07 = reg_0732;
    97: op1_02_in07 = reg_0894;
    default: op1_02_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv07 = 1;
    13: op1_02_inv07 = 1;
    14: op1_02_inv07 = 1;
    15: op1_02_inv07 = 1;
    17: op1_02_inv07 = 1;
    22: op1_02_inv07 = 1;
    24: op1_02_inv07 = 1;
    25: op1_02_inv07 = 1;
    26: op1_02_inv07 = 1;
    28: op1_02_inv07 = 1;
    30: op1_02_inv07 = 1;
    31: op1_02_inv07 = 1;
    33: op1_02_inv07 = 1;
    34: op1_02_inv07 = 1;
    37: op1_02_inv07 = 1;
    39: op1_02_inv07 = 1;
    41: op1_02_inv07 = 1;
    43: op1_02_inv07 = 1;
    46: op1_02_inv07 = 1;
    47: op1_02_inv07 = 1;
    48: op1_02_inv07 = 1;
    49: op1_02_inv07 = 1;
    52: op1_02_inv07 = 1;
    53: op1_02_inv07 = 1;
    56: op1_02_inv07 = 1;
    57: op1_02_inv07 = 1;
    58: op1_02_inv07 = 1;
    60: op1_02_inv07 = 1;
    62: op1_02_inv07 = 1;
    63: op1_02_inv07 = 1;
    65: op1_02_inv07 = 1;
    75: op1_02_inv07 = 1;
    81: op1_02_inv07 = 1;
    83: op1_02_inv07 = 1;
    84: op1_02_inv07 = 1;
    85: op1_02_inv07 = 1;
    86: op1_02_inv07 = 1;
    87: op1_02_inv07 = 1;
    91: op1_02_inv07 = 1;
    92: op1_02_inv07 = 1;
    94: op1_02_inv07 = 1;
    97: op1_02_inv07 = 1;
    default: op1_02_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in08 = reg_0583;
    6: op1_02_in08 = reg_0462;
    7: op1_02_in08 = reg_0301;
    16: op1_02_in08 = reg_0301;
    8: op1_02_in08 = reg_0673;
    9: op1_02_in08 = reg_0083;
    10: op1_02_in08 = reg_0982;
    3: op1_02_in08 = reg_0157;
    11: op1_02_in08 = reg_0304;
    12: op1_02_in08 = reg_0101;
    13: op1_02_in08 = reg_0393;
    14: op1_02_in08 = reg_0453;
    15: op1_02_in08 = imem03_in[19:16];
    17: op1_02_in08 = reg_0729;
    18: op1_02_in08 = reg_0659;
    19: op1_02_in08 = reg_0693;
    20: op1_02_in08 = reg_0358;
    21: op1_02_in08 = reg_0402;
    22: op1_02_in08 = reg_0339;
    23: op1_02_in08 = reg_1000;
    24: op1_02_in08 = reg_0188;
    25: op1_02_in08 = reg_0059;
    26: op1_02_in08 = reg_0787;
    27: op1_02_in08 = reg_0283;
    28: op1_02_in08 = reg_0011;
    29: op1_02_in08 = reg_0097;
    30: op1_02_in08 = reg_0543;
    47: op1_02_in08 = reg_0543;
    31: op1_02_in08 = reg_0717;
    32: op1_02_in08 = reg_0120;
    33: op1_02_in08 = reg_0795;
    34: op1_02_in08 = reg_0733;
    35: op1_02_in08 = reg_0666;
    36: op1_02_in08 = reg_0463;
    37: op1_02_in08 = reg_0661;
    38: op1_02_in08 = reg_0984;
    39: op1_02_in08 = reg_0998;
    40: op1_02_in08 = reg_0614;
    41: op1_02_in08 = reg_0973;
    42: op1_02_in08 = reg_0698;
    43: op1_02_in08 = imem02_in[59:56];
    44: op1_02_in08 = reg_0995;
    45: op1_02_in08 = imem06_in[87:84];
    46: op1_02_in08 = reg_0684;
    79: op1_02_in08 = reg_0684;
    48: op1_02_in08 = imem05_in[3:0];
    49: op1_02_in08 = reg_0676;
    50: op1_02_in08 = imem00_in[99:96];
    51: op1_02_in08 = reg_0160;
    52: op1_02_in08 = reg_0493;
    53: op1_02_in08 = reg_0556;
    54: op1_02_in08 = reg_0241;
    63: op1_02_in08 = reg_0241;
    55: op1_02_in08 = imem07_in[71:68];
    56: op1_02_in08 = reg_0466;
    57: op1_02_in08 = imem02_in[3:0];
    58: op1_02_in08 = imem02_in[111:108];
    59: op1_02_in08 = reg_0680;
    60: op1_02_in08 = imem04_in[11:8];
    61: op1_02_in08 = reg_0389;
    62: op1_02_in08 = reg_0807;
    65: op1_02_in08 = reg_0843;
    66: op1_02_in08 = reg_0668;
    67: op1_02_in08 = reg_0883;
    68: op1_02_in08 = reg_0460;
    69: op1_02_in08 = imem05_in[75:72];
    70: op1_02_in08 = imem07_in[107:104];
    71: op1_02_in08 = reg_0906;
    72: op1_02_in08 = imem07_in[63:60];
    73: op1_02_in08 = reg_0465;
    74: op1_02_in08 = reg_0748;
    75: op1_02_in08 = imem02_in[87:84];
    76: op1_02_in08 = reg_0302;
    77: op1_02_in08 = imem04_in[47:44];
    78: op1_02_in08 = reg_0028;
    80: op1_02_in08 = reg_0687;
    81: op1_02_in08 = reg_0082;
    82: op1_02_in08 = reg_0833;
    83: op1_02_in08 = imem07_in[95:92];
    84: op1_02_in08 = reg_0215;
    85: op1_02_in08 = reg_0470;
    86: op1_02_in08 = reg_0642;
    88: op1_02_in08 = reg_0703;
    89: op1_02_in08 = reg_0086;
    90: op1_02_in08 = reg_0477;
    91: op1_02_in08 = reg_0450;
    92: op1_02_in08 = reg_0166;
    93: op1_02_in08 = imem05_in[7:4];
    94: op1_02_in08 = reg_0288;
    95: op1_02_in08 = reg_0568;
    96: op1_02_in08 = reg_0284;
    97: op1_02_in08 = imem03_in[27:24];
    default: op1_02_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_02_inv08 = 1;
    8: op1_02_inv08 = 1;
    9: op1_02_inv08 = 1;
    3: op1_02_inv08 = 1;
    11: op1_02_inv08 = 1;
    15: op1_02_inv08 = 1;
    16: op1_02_inv08 = 1;
    17: op1_02_inv08 = 1;
    18: op1_02_inv08 = 1;
    21: op1_02_inv08 = 1;
    22: op1_02_inv08 = 1;
    25: op1_02_inv08 = 1;
    29: op1_02_inv08 = 1;
    30: op1_02_inv08 = 1;
    31: op1_02_inv08 = 1;
    33: op1_02_inv08 = 1;
    36: op1_02_inv08 = 1;
    38: op1_02_inv08 = 1;
    40: op1_02_inv08 = 1;
    41: op1_02_inv08 = 1;
    44: op1_02_inv08 = 1;
    47: op1_02_inv08 = 1;
    48: op1_02_inv08 = 1;
    49: op1_02_inv08 = 1;
    50: op1_02_inv08 = 1;
    52: op1_02_inv08 = 1;
    53: op1_02_inv08 = 1;
    54: op1_02_inv08 = 1;
    55: op1_02_inv08 = 1;
    56: op1_02_inv08 = 1;
    57: op1_02_inv08 = 1;
    58: op1_02_inv08 = 1;
    59: op1_02_inv08 = 1;
    60: op1_02_inv08 = 1;
    62: op1_02_inv08 = 1;
    65: op1_02_inv08 = 1;
    69: op1_02_inv08 = 1;
    70: op1_02_inv08 = 1;
    72: op1_02_inv08 = 1;
    73: op1_02_inv08 = 1;
    74: op1_02_inv08 = 1;
    78: op1_02_inv08 = 1;
    82: op1_02_inv08 = 1;
    88: op1_02_inv08 = 1;
    90: op1_02_inv08 = 1;
    92: op1_02_inv08 = 1;
    93: op1_02_inv08 = 1;
    94: op1_02_inv08 = 1;
    95: op1_02_inv08 = 1;
    96: op1_02_inv08 = 1;
    97: op1_02_inv08 = 1;
    default: op1_02_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in09 = reg_0568;
    6: op1_02_in09 = reg_0467;
    7: op1_02_in09 = reg_0292;
    8: op1_02_in09 = reg_0687;
    9: op1_02_in09 = reg_0090;
    10: op1_02_in09 = reg_0995;
    3: op1_02_in09 = reg_0173;
    11: op1_02_in09 = reg_0281;
    12: op1_02_in09 = imem02_in[3:0];
    13: op1_02_in09 = reg_0389;
    14: op1_02_in09 = reg_0451;
    73: op1_02_in09 = reg_0451;
    15: op1_02_in09 = imem03_in[47:44];
    16: op1_02_in09 = reg_0283;
    17: op1_02_in09 = reg_0425;
    18: op1_02_in09 = reg_0636;
    19: op1_02_in09 = reg_0676;
    20: op1_02_in09 = reg_0330;
    21: op1_02_in09 = reg_0349;
    22: op1_02_in09 = reg_0342;
    23: op1_02_in09 = imem04_in[15:12];
    24: op1_02_in09 = reg_0207;
    25: op1_02_in09 = reg_0875;
    26: op1_02_in09 = reg_0027;
    27: op1_02_in09 = reg_0279;
    28: op1_02_in09 = imem07_in[23:20];
    29: op1_02_in09 = reg_0290;
    30: op1_02_in09 = reg_0038;
    31: op1_02_in09 = reg_0709;
    32: op1_02_in09 = reg_0108;
    33: op1_02_in09 = reg_0836;
    34: op1_02_in09 = reg_0076;
    35: op1_02_in09 = reg_0660;
    36: op1_02_in09 = reg_0457;
    37: op1_02_in09 = reg_0639;
    38: op1_02_in09 = reg_0980;
    39: op1_02_in09 = reg_0982;
    40: op1_02_in09 = reg_0856;
    41: op1_02_in09 = reg_0944;
    42: op1_02_in09 = reg_0686;
    43: op1_02_in09 = imem02_in[79:76];
    44: op1_02_in09 = reg_1001;
    45: op1_02_in09 = imem06_in[127:124];
    46: op1_02_in09 = reg_0668;
    47: op1_02_in09 = reg_0509;
    48: op1_02_in09 = imem05_in[7:4];
    49: op1_02_in09 = reg_0684;
    50: op1_02_in09 = imem00_in[123:120];
    51: op1_02_in09 = reg_0163;
    52: op1_02_in09 = reg_0237;
    53: op1_02_in09 = reg_0632;
    54: op1_02_in09 = reg_0609;
    55: op1_02_in09 = imem07_in[79:76];
    56: op1_02_in09 = reg_0479;
    57: op1_02_in09 = imem02_in[35:32];
    58: op1_02_in09 = reg_0326;
    59: op1_02_in09 = reg_0453;
    60: op1_02_in09 = imem04_in[35:32];
    61: op1_02_in09 = reg_0331;
    62: op1_02_in09 = reg_0376;
    63: op1_02_in09 = reg_0371;
    65: op1_02_in09 = reg_0499;
    66: op1_02_in09 = reg_0680;
    67: op1_02_in09 = reg_0069;
    68: op1_02_in09 = reg_0480;
    69: op1_02_in09 = imem05_in[87:84];
    70: op1_02_in09 = reg_0325;
    71: op1_02_in09 = reg_0832;
    72: op1_02_in09 = imem07_in[99:96];
    74: op1_02_in09 = reg_0900;
    75: op1_02_in09 = reg_0750;
    76: op1_02_in09 = reg_0276;
    77: op1_02_in09 = imem04_in[55:52];
    78: op1_02_in09 = reg_0440;
    79: op1_02_in09 = reg_0356;
    80: op1_02_in09 = reg_0749;
    81: op1_02_in09 = reg_0034;
    82: op1_02_in09 = reg_0887;
    83: op1_02_in09 = imem07_in[103:100];
    84: op1_02_in09 = reg_0136;
    85: op1_02_in09 = reg_0474;
    86: op1_02_in09 = reg_0664;
    88: op1_02_in09 = reg_0714;
    89: op1_02_in09 = reg_0656;
    90: op1_02_in09 = reg_0472;
    91: op1_02_in09 = reg_0455;
    92: op1_02_in09 = reg_0386;
    93: op1_02_in09 = imem05_in[83:80];
    94: op1_02_in09 = reg_0432;
    96: op1_02_in09 = reg_0432;
    95: op1_02_in09 = reg_0015;
    97: op1_02_in09 = imem03_in[39:36];
    default: op1_02_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv09 = 1;
    7: op1_02_inv09 = 1;
    8: op1_02_inv09 = 1;
    11: op1_02_inv09 = 1;
    15: op1_02_inv09 = 1;
    16: op1_02_inv09 = 1;
    17: op1_02_inv09 = 1;
    18: op1_02_inv09 = 1;
    19: op1_02_inv09 = 1;
    21: op1_02_inv09 = 1;
    22: op1_02_inv09 = 1;
    23: op1_02_inv09 = 1;
    24: op1_02_inv09 = 1;
    25: op1_02_inv09 = 1;
    26: op1_02_inv09 = 1;
    27: op1_02_inv09 = 1;
    28: op1_02_inv09 = 1;
    30: op1_02_inv09 = 1;
    35: op1_02_inv09 = 1;
    36: op1_02_inv09 = 1;
    41: op1_02_inv09 = 1;
    43: op1_02_inv09 = 1;
    45: op1_02_inv09 = 1;
    46: op1_02_inv09 = 1;
    47: op1_02_inv09 = 1;
    49: op1_02_inv09 = 1;
    52: op1_02_inv09 = 1;
    61: op1_02_inv09 = 1;
    68: op1_02_inv09 = 1;
    69: op1_02_inv09 = 1;
    70: op1_02_inv09 = 1;
    72: op1_02_inv09 = 1;
    75: op1_02_inv09 = 1;
    76: op1_02_inv09 = 1;
    78: op1_02_inv09 = 1;
    79: op1_02_inv09 = 1;
    81: op1_02_inv09 = 1;
    83: op1_02_inv09 = 1;
    86: op1_02_inv09 = 1;
    92: op1_02_inv09 = 1;
    94: op1_02_inv09 = 1;
    default: op1_02_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in10 = reg_0569;
    6: op1_02_in10 = reg_0470;
    7: op1_02_in10 = reg_0062;
    8: op1_02_in10 = reg_0451;
    9: op1_02_in10 = imem03_in[31:28];
    10: op1_02_in10 = reg_0984;
    3: op1_02_in10 = reg_0171;
    11: op1_02_in10 = reg_0305;
    12: op1_02_in10 = imem02_in[39:36];
    13: op1_02_in10 = reg_0982;
    14: op1_02_in10 = reg_0455;
    73: op1_02_in10 = reg_0455;
    15: op1_02_in10 = imem03_in[51:48];
    16: op1_02_in10 = reg_0289;
    17: op1_02_in10 = reg_0433;
    18: op1_02_in10 = reg_0663;
    19: op1_02_in10 = reg_0689;
    20: op1_02_in10 = reg_0363;
    21: op1_02_in10 = reg_0403;
    22: op1_02_in10 = reg_0338;
    23: op1_02_in10 = imem04_in[43:40];
    24: op1_02_in10 = reg_0201;
    25: op1_02_in10 = reg_0057;
    26: op1_02_in10 = reg_0026;
    27: op1_02_in10 = reg_0751;
    28: op1_02_in10 = imem07_in[95:92];
    29: op1_02_in10 = reg_0817;
    30: op1_02_in10 = reg_0373;
    31: op1_02_in10 = reg_0727;
    32: op1_02_in10 = reg_0110;
    33: op1_02_in10 = reg_0987;
    34: op1_02_in10 = reg_0067;
    35: op1_02_in10 = reg_0651;
    36: op1_02_in10 = reg_0481;
    37: op1_02_in10 = reg_0638;
    38: op1_02_in10 = reg_0977;
    39: op1_02_in10 = reg_0979;
    40: op1_02_in10 = reg_0371;
    41: op1_02_in10 = reg_0969;
    42: op1_02_in10 = reg_0670;
    49: op1_02_in10 = reg_0670;
    43: op1_02_in10 = imem02_in[119:116];
    44: op1_02_in10 = reg_0990;
    45: op1_02_in10 = reg_0856;
    46: op1_02_in10 = reg_0477;
    47: op1_02_in10 = reg_0807;
    48: op1_02_in10 = imem05_in[39:36];
    50: op1_02_in10 = reg_0693;
    51: op1_02_in10 = reg_0183;
    52: op1_02_in10 = reg_1046;
    53: op1_02_in10 = reg_0612;
    54: op1_02_in10 = reg_0626;
    55: op1_02_in10 = reg_0716;
    72: op1_02_in10 = reg_0716;
    56: op1_02_in10 = reg_0478;
    57: op1_02_in10 = imem02_in[55:52];
    58: op1_02_in10 = reg_0515;
    59: op1_02_in10 = reg_0457;
    91: op1_02_in10 = reg_0457;
    60: op1_02_in10 = imem04_in[59:56];
    61: op1_02_in10 = reg_0772;
    62: op1_02_in10 = reg_0991;
    63: op1_02_in10 = imem07_in[3:0];
    65: op1_02_in10 = reg_0069;
    66: op1_02_in10 = reg_0465;
    67: op1_02_in10 = reg_0463;
    68: op1_02_in10 = reg_0459;
    85: op1_02_in10 = reg_0459;
    69: op1_02_in10 = imem05_in[107:104];
    70: op1_02_in10 = reg_0321;
    71: op1_02_in10 = reg_0003;
    74: op1_02_in10 = reg_0475;
    75: op1_02_in10 = reg_0844;
    76: op1_02_in10 = reg_0296;
    77: op1_02_in10 = imem04_in[79:76];
    78: op1_02_in10 = reg_0895;
    79: op1_02_in10 = reg_0466;
    80: op1_02_in10 = reg_0450;
    81: op1_02_in10 = reg_0643;
    82: op1_02_in10 = reg_0643;
    83: op1_02_in10 = reg_0165;
    84: op1_02_in10 = reg_0652;
    86: op1_02_in10 = reg_0423;
    88: op1_02_in10 = reg_0185;
    89: op1_02_in10 = reg_0713;
    90: op1_02_in10 = reg_0480;
    92: op1_02_in10 = reg_0223;
    93: op1_02_in10 = reg_0217;
    94: op1_02_in10 = reg_0065;
    95: op1_02_in10 = reg_0732;
    96: op1_02_in10 = reg_0027;
    97: op1_02_in10 = imem03_in[83:80];
    default: op1_02_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv10 = 1;
    8: op1_02_inv10 = 1;
    9: op1_02_inv10 = 1;
    10: op1_02_inv10 = 1;
    3: op1_02_inv10 = 1;
    11: op1_02_inv10 = 1;
    14: op1_02_inv10 = 1;
    15: op1_02_inv10 = 1;
    16: op1_02_inv10 = 1;
    17: op1_02_inv10 = 1;
    18: op1_02_inv10 = 1;
    23: op1_02_inv10 = 1;
    24: op1_02_inv10 = 1;
    25: op1_02_inv10 = 1;
    33: op1_02_inv10 = 1;
    34: op1_02_inv10 = 1;
    35: op1_02_inv10 = 1;
    36: op1_02_inv10 = 1;
    37: op1_02_inv10 = 1;
    38: op1_02_inv10 = 1;
    39: op1_02_inv10 = 1;
    41: op1_02_inv10 = 1;
    43: op1_02_inv10 = 1;
    45: op1_02_inv10 = 1;
    47: op1_02_inv10 = 1;
    48: op1_02_inv10 = 1;
    51: op1_02_inv10 = 1;
    52: op1_02_inv10 = 1;
    53: op1_02_inv10 = 1;
    55: op1_02_inv10 = 1;
    56: op1_02_inv10 = 1;
    58: op1_02_inv10 = 1;
    59: op1_02_inv10 = 1;
    61: op1_02_inv10 = 1;
    65: op1_02_inv10 = 1;
    67: op1_02_inv10 = 1;
    68: op1_02_inv10 = 1;
    69: op1_02_inv10 = 1;
    70: op1_02_inv10 = 1;
    71: op1_02_inv10 = 1;
    74: op1_02_inv10 = 1;
    76: op1_02_inv10 = 1;
    77: op1_02_inv10 = 1;
    78: op1_02_inv10 = 1;
    81: op1_02_inv10 = 1;
    82: op1_02_inv10 = 1;
    84: op1_02_inv10 = 1;
    86: op1_02_inv10 = 1;
    88: op1_02_inv10 = 1;
    89: op1_02_inv10 = 1;
    92: op1_02_inv10 = 1;
    96: op1_02_inv10 = 1;
    97: op1_02_inv10 = 1;
    default: op1_02_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in11 = reg_0584;
    6: op1_02_in11 = reg_0474;
    7: op1_02_in11 = reg_0058;
    8: op1_02_in11 = reg_0469;
    46: op1_02_in11 = reg_0469;
    9: op1_02_in11 = imem03_in[47:44];
    10: op1_02_in11 = reg_0980;
    3: op1_02_in11 = reg_0184;
    11: op1_02_in11 = reg_0299;
    12: op1_02_in11 = imem02_in[71:68];
    13: op1_02_in11 = reg_0989;
    14: op1_02_in11 = reg_0461;
    15: op1_02_in11 = imem03_in[67:64];
    16: op1_02_in11 = reg_0290;
    17: op1_02_in11 = reg_0419;
    70: op1_02_in11 = reg_0419;
    18: op1_02_in11 = reg_0358;
    19: op1_02_in11 = reg_0684;
    20: op1_02_in11 = reg_0365;
    21: op1_02_in11 = reg_0337;
    22: op1_02_in11 = reg_0083;
    23: op1_02_in11 = imem04_in[99:96];
    24: op1_02_in11 = imem01_in[35:32];
    25: op1_02_in11 = reg_0044;
    26: op1_02_in11 = reg_0486;
    27: op1_02_in11 = reg_0057;
    28: op1_02_in11 = reg_0716;
    29: op1_02_in11 = reg_0007;
    30: op1_02_in11 = reg_0509;
    31: op1_02_in11 = reg_0429;
    32: op1_02_in11 = imem02_in[7:4];
    33: op1_02_in11 = reg_0986;
    34: op1_02_in11 = reg_0259;
    35: op1_02_in11 = reg_0641;
    36: op1_02_in11 = reg_0203;
    37: op1_02_in11 = reg_0636;
    38: op1_02_in11 = reg_0975;
    39: op1_02_in11 = reg_0984;
    40: op1_02_in11 = reg_0783;
    41: op1_02_in11 = reg_0951;
    42: op1_02_in11 = reg_0679;
    43: op1_02_in11 = imem02_in[127:124];
    44: op1_02_in11 = imem04_in[7:4];
    45: op1_02_in11 = reg_0892;
    47: op1_02_in11 = reg_0513;
    48: op1_02_in11 = imem05_in[79:76];
    49: op1_02_in11 = reg_0673;
    50: op1_02_in11 = reg_0672;
    51: op1_02_in11 = reg_0164;
    52: op1_02_in11 = reg_0447;
    53: op1_02_in11 = reg_0387;
    54: op1_02_in11 = reg_0531;
    55: op1_02_in11 = reg_0720;
    56: op1_02_in11 = reg_0189;
    57: op1_02_in11 = imem02_in[59:56];
    58: op1_02_in11 = reg_0651;
    59: op1_02_in11 = reg_0478;
    60: op1_02_in11 = imem04_in[79:76];
    61: op1_02_in11 = reg_0090;
    62: op1_02_in11 = reg_0976;
    63: op1_02_in11 = imem07_in[11:8];
    65: op1_02_in11 = reg_0687;
    66: op1_02_in11 = reg_0475;
    67: op1_02_in11 = reg_0477;
    68: op1_02_in11 = reg_0456;
    69: op1_02_in11 = imem05_in[111:108];
    71: op1_02_in11 = reg_0273;
    72: op1_02_in11 = reg_0719;
    73: op1_02_in11 = reg_0457;
    74: op1_02_in11 = reg_0460;
    75: op1_02_in11 = reg_0916;
    76: op1_02_in11 = reg_0288;
    77: op1_02_in11 = reg_0301;
    78: op1_02_in11 = reg_0863;
    79: op1_02_in11 = reg_0470;
    80: op1_02_in11 = reg_0451;
    81: op1_02_in11 = reg_0279;
    82: op1_02_in11 = reg_0908;
    83: op1_02_in11 = reg_0162;
    84: op1_02_in11 = reg_0128;
    85: op1_02_in11 = reg_0208;
    86: op1_02_in11 = reg_0516;
    88: op1_02_in11 = reg_0697;
    89: op1_02_in11 = imem03_in[75:72];
    90: op1_02_in11 = reg_0204;
    91: op1_02_in11 = reg_0464;
    92: op1_02_in11 = reg_0030;
    93: op1_02_in11 = reg_0652;
    94: op1_02_in11 = reg_0627;
    95: op1_02_in11 = reg_0893;
    96: op1_02_in11 = reg_0295;
    97: op1_02_in11 = reg_0819;
    default: op1_02_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv11 = 1;
    6: op1_02_inv11 = 1;
    8: op1_02_inv11 = 1;
    9: op1_02_inv11 = 1;
    3: op1_02_inv11 = 1;
    11: op1_02_inv11 = 1;
    12: op1_02_inv11 = 1;
    13: op1_02_inv11 = 1;
    14: op1_02_inv11 = 1;
    21: op1_02_inv11 = 1;
    22: op1_02_inv11 = 1;
    24: op1_02_inv11 = 1;
    26: op1_02_inv11 = 1;
    27: op1_02_inv11 = 1;
    31: op1_02_inv11 = 1;
    32: op1_02_inv11 = 1;
    34: op1_02_inv11 = 1;
    35: op1_02_inv11 = 1;
    37: op1_02_inv11 = 1;
    38: op1_02_inv11 = 1;
    39: op1_02_inv11 = 1;
    41: op1_02_inv11 = 1;
    45: op1_02_inv11 = 1;
    46: op1_02_inv11 = 1;
    47: op1_02_inv11 = 1;
    48: op1_02_inv11 = 1;
    51: op1_02_inv11 = 1;
    52: op1_02_inv11 = 1;
    53: op1_02_inv11 = 1;
    55: op1_02_inv11 = 1;
    57: op1_02_inv11 = 1;
    58: op1_02_inv11 = 1;
    59: op1_02_inv11 = 1;
    60: op1_02_inv11 = 1;
    66: op1_02_inv11 = 1;
    67: op1_02_inv11 = 1;
    69: op1_02_inv11 = 1;
    74: op1_02_inv11 = 1;
    75: op1_02_inv11 = 1;
    81: op1_02_inv11 = 1;
    84: op1_02_inv11 = 1;
    85: op1_02_inv11 = 1;
    86: op1_02_inv11 = 1;
    88: op1_02_inv11 = 1;
    89: op1_02_inv11 = 1;
    92: op1_02_inv11 = 1;
    93: op1_02_inv11 = 1;
    94: op1_02_inv11 = 1;
    default: op1_02_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in12 = reg_0585;
    6: op1_02_in12 = reg_0468;
    66: op1_02_in12 = reg_0468;
    7: op1_02_in12 = reg_0064;
    8: op1_02_in12 = reg_0480;
    9: op1_02_in12 = imem03_in[87:84];
    10: op1_02_in12 = reg_0999;
    11: op1_02_in12 = reg_0285;
    12: op1_02_in12 = reg_0653;
    13: op1_02_in12 = reg_0974;
    14: op1_02_in12 = reg_0460;
    15: op1_02_in12 = imem03_in[83:80];
    16: op1_02_in12 = reg_0292;
    17: op1_02_in12 = reg_0446;
    18: op1_02_in12 = reg_0320;
    19: op1_02_in12 = reg_0686;
    20: op1_02_in12 = reg_0097;
    21: op1_02_in12 = reg_0401;
    22: op1_02_in12 = reg_0776;
    23: op1_02_in12 = imem04_in[107:104];
    24: op1_02_in12 = imem01_in[47:44];
    25: op1_02_in12 = reg_0021;
    26: op1_02_in12 = reg_0801;
    27: op1_02_in12 = reg_0286;
    28: op1_02_in12 = reg_0725;
    29: op1_02_in12 = reg_0482;
    30: op1_02_in12 = reg_0836;
    31: op1_02_in12 = reg_0432;
    32: op1_02_in12 = imem02_in[15:12];
    33: op1_02_in12 = reg_0981;
    34: op1_02_in12 = reg_0071;
    35: op1_02_in12 = reg_0318;
    36: op1_02_in12 = imem01_in[31:28];
    37: op1_02_in12 = reg_0007;
    38: op1_02_in12 = reg_1000;
    39: op1_02_in12 = reg_0980;
    40: op1_02_in12 = reg_0612;
    41: op1_02_in12 = reg_0953;
    42: op1_02_in12 = reg_0675;
    43: op1_02_in12 = reg_0646;
    44: op1_02_in12 = reg_0277;
    45: op1_02_in12 = reg_0627;
    46: op1_02_in12 = reg_0459;
    47: op1_02_in12 = reg_0822;
    48: op1_02_in12 = reg_0963;
    49: op1_02_in12 = reg_0465;
    50: op1_02_in12 = reg_0676;
    51: op1_02_in12 = reg_0168;
    52: op1_02_in12 = reg_0269;
    53: op1_02_in12 = reg_0344;
    54: op1_02_in12 = reg_0029;
    55: op1_02_in12 = reg_0723;
    56: op1_02_in12 = reg_0194;
    57: op1_02_in12 = imem02_in[67:64];
    58: op1_02_in12 = reg_0636;
    59: op1_02_in12 = reg_0458;
    60: op1_02_in12 = imem04_in[119:116];
    61: op1_02_in12 = reg_0091;
    62: op1_02_in12 = imem04_in[7:4];
    63: op1_02_in12 = imem07_in[71:68];
    65: op1_02_in12 = reg_0451;
    67: op1_02_in12 = reg_0476;
    68: op1_02_in12 = reg_0186;
    69: op1_02_in12 = reg_0655;
    70: op1_02_in12 = reg_0180;
    71: op1_02_in12 = reg_0101;
    72: op1_02_in12 = reg_0731;
    73: op1_02_in12 = reg_0477;
    74: op1_02_in12 = reg_0191;
    75: op1_02_in12 = reg_0666;
    76: op1_02_in12 = reg_0284;
    77: op1_02_in12 = reg_0537;
    78: op1_02_in12 = reg_0804;
    79: op1_02_in12 = reg_0452;
    80: op1_02_in12 = reg_0457;
    81: op1_02_in12 = reg_0425;
    82: op1_02_in12 = reg_0418;
    83: op1_02_in12 = reg_0726;
    84: op1_02_in12 = reg_0142;
    85: op1_02_in12 = reg_0193;
    86: op1_02_in12 = reg_0355;
    89: op1_02_in12 = imem03_in[79:76];
    90: op1_02_in12 = reg_0203;
    91: op1_02_in12 = reg_0461;
    92: op1_02_in12 = reg_0455;
    93: op1_02_in12 = reg_0954;
    94: op1_02_in12 = reg_0854;
    95: op1_02_in12 = reg_0243;
    96: op1_02_in12 = imem05_in[7:4];
    97: op1_02_in12 = reg_0357;
    default: op1_02_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_02_inv12 = 1;
    8: op1_02_inv12 = 1;
    10: op1_02_inv12 = 1;
    13: op1_02_inv12 = 1;
    14: op1_02_inv12 = 1;
    16: op1_02_inv12 = 1;
    17: op1_02_inv12 = 1;
    20: op1_02_inv12 = 1;
    23: op1_02_inv12 = 1;
    25: op1_02_inv12 = 1;
    26: op1_02_inv12 = 1;
    27: op1_02_inv12 = 1;
    28: op1_02_inv12 = 1;
    30: op1_02_inv12 = 1;
    34: op1_02_inv12 = 1;
    38: op1_02_inv12 = 1;
    39: op1_02_inv12 = 1;
    40: op1_02_inv12 = 1;
    41: op1_02_inv12 = 1;
    42: op1_02_inv12 = 1;
    43: op1_02_inv12 = 1;
    46: op1_02_inv12 = 1;
    47: op1_02_inv12 = 1;
    48: op1_02_inv12 = 1;
    52: op1_02_inv12 = 1;
    53: op1_02_inv12 = 1;
    54: op1_02_inv12 = 1;
    55: op1_02_inv12 = 1;
    57: op1_02_inv12 = 1;
    60: op1_02_inv12 = 1;
    65: op1_02_inv12 = 1;
    69: op1_02_inv12 = 1;
    71: op1_02_inv12 = 1;
    75: op1_02_inv12 = 1;
    77: op1_02_inv12 = 1;
    79: op1_02_inv12 = 1;
    84: op1_02_inv12 = 1;
    85: op1_02_inv12 = 1;
    86: op1_02_inv12 = 1;
    90: op1_02_inv12 = 1;
    92: op1_02_inv12 = 1;
    93: op1_02_inv12 = 1;
    95: op1_02_inv12 = 1;
    96: op1_02_inv12 = 1;
    97: op1_02_inv12 = 1;
    default: op1_02_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in13 = reg_0578;
    6: op1_02_in13 = reg_0459;
    66: op1_02_in13 = reg_0459;
    7: op1_02_in13 = reg_0044;
    8: op1_02_in13 = reg_0468;
    9: op1_02_in13 = imem03_in[103:100];
    10: op1_02_in13 = reg_0989;
    11: op1_02_in13 = reg_0295;
    12: op1_02_in13 = reg_0657;
    13: op1_02_in13 = reg_0983;
    14: op1_02_in13 = reg_0462;
    15: op1_02_in13 = imem03_in[99:96];
    16: op1_02_in13 = reg_0286;
    17: op1_02_in13 = reg_0168;
    18: op1_02_in13 = reg_0363;
    19: op1_02_in13 = reg_0691;
    20: op1_02_in13 = imem03_in[3:0];
    21: op1_02_in13 = reg_0799;
    77: op1_02_in13 = reg_0799;
    22: op1_02_in13 = reg_0761;
    29: op1_02_in13 = reg_0761;
    23: op1_02_in13 = imem04_in[123:120];
    24: op1_02_in13 = imem01_in[123:120];
    25: op1_02_in13 = imem05_in[11:8];
    94: op1_02_in13 = imem05_in[11:8];
    26: op1_02_in13 = reg_0025;
    27: op1_02_in13 = reg_0856;
    28: op1_02_in13 = reg_0724;
    30: op1_02_in13 = reg_0986;
    31: op1_02_in13 = reg_0422;
    32: op1_02_in13 = imem02_in[31:28];
    33: op1_02_in13 = reg_0997;
    34: op1_02_in13 = reg_0075;
    35: op1_02_in13 = reg_0857;
    36: op1_02_in13 = imem01_in[35:32];
    37: op1_02_in13 = reg_0482;
    38: op1_02_in13 = imem04_in[15:12];
    39: op1_02_in13 = reg_0974;
    40: op1_02_in13 = reg_0386;
    41: op1_02_in13 = reg_0972;
    42: op1_02_in13 = reg_0688;
    43: op1_02_in13 = reg_0660;
    44: op1_02_in13 = reg_0539;
    45: op1_02_in13 = reg_0495;
    46: op1_02_in13 = reg_0208;
    47: op1_02_in13 = reg_0985;
    48: op1_02_in13 = reg_0958;
    49: op1_02_in13 = reg_0450;
    50: op1_02_in13 = reg_0686;
    51: op1_02_in13 = reg_0170;
    52: op1_02_in13 = reg_0128;
    53: op1_02_in13 = reg_0399;
    54: op1_02_in13 = reg_0622;
    55: op1_02_in13 = reg_0725;
    56: op1_02_in13 = reg_0197;
    57: op1_02_in13 = imem02_in[75:72];
    58: op1_02_in13 = reg_0739;
    59: op1_02_in13 = reg_0214;
    60: op1_02_in13 = reg_0277;
    61: op1_02_in13 = reg_0840;
    62: op1_02_in13 = imem04_in[23:20];
    63: op1_02_in13 = imem07_in[83:80];
    65: op1_02_in13 = reg_0461;
    67: op1_02_in13 = reg_0481;
    68: op1_02_in13 = reg_0212;
    69: op1_02_in13 = reg_0030;
    70: op1_02_in13 = reg_0162;
    71: op1_02_in13 = reg_0117;
    72: op1_02_in13 = reg_0721;
    73: op1_02_in13 = reg_0470;
    74: op1_02_in13 = reg_0190;
    75: op1_02_in13 = reg_0810;
    76: op1_02_in13 = reg_0893;
    78: op1_02_in13 = reg_0026;
    79: op1_02_in13 = reg_0478;
    80: op1_02_in13 = reg_0475;
    81: op1_02_in13 = reg_0248;
    82: op1_02_in13 = reg_0279;
    83: op1_02_in13 = reg_0717;
    84: op1_02_in13 = reg_0143;
    85: op1_02_in13 = reg_0196;
    86: op1_02_in13 = reg_0086;
    89: op1_02_in13 = imem03_in[95:92];
    90: op1_02_in13 = reg_0211;
    91: op1_02_in13 = reg_0479;
    92: op1_02_in13 = reg_0457;
    93: op1_02_in13 = reg_0655;
    95: op1_02_in13 = reg_0041;
    96: op1_02_in13 = imem05_in[31:28];
    97: op1_02_in13 = reg_0317;
    default: op1_02_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv13 = 1;
    8: op1_02_inv13 = 1;
    9: op1_02_inv13 = 1;
    10: op1_02_inv13 = 1;
    12: op1_02_inv13 = 1;
    13: op1_02_inv13 = 1;
    14: op1_02_inv13 = 1;
    17: op1_02_inv13 = 1;
    18: op1_02_inv13 = 1;
    22: op1_02_inv13 = 1;
    23: op1_02_inv13 = 1;
    25: op1_02_inv13 = 1;
    28: op1_02_inv13 = 1;
    29: op1_02_inv13 = 1;
    30: op1_02_inv13 = 1;
    33: op1_02_inv13 = 1;
    39: op1_02_inv13 = 1;
    43: op1_02_inv13 = 1;
    46: op1_02_inv13 = 1;
    48: op1_02_inv13 = 1;
    49: op1_02_inv13 = 1;
    52: op1_02_inv13 = 1;
    53: op1_02_inv13 = 1;
    54: op1_02_inv13 = 1;
    55: op1_02_inv13 = 1;
    57: op1_02_inv13 = 1;
    58: op1_02_inv13 = 1;
    59: op1_02_inv13 = 1;
    60: op1_02_inv13 = 1;
    65: op1_02_inv13 = 1;
    66: op1_02_inv13 = 1;
    68: op1_02_inv13 = 1;
    71: op1_02_inv13 = 1;
    74: op1_02_inv13 = 1;
    76: op1_02_inv13 = 1;
    77: op1_02_inv13 = 1;
    79: op1_02_inv13 = 1;
    82: op1_02_inv13 = 1;
    90: op1_02_inv13 = 1;
    91: op1_02_inv13 = 1;
    92: op1_02_inv13 = 1;
    93: op1_02_inv13 = 1;
    default: op1_02_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in14 = reg_0570;
    6: op1_02_in14 = reg_0211;
    7: op1_02_in14 = imem05_in[7:4];
    8: op1_02_in14 = reg_0459;
    91: op1_02_in14 = reg_0459;
    9: op1_02_in14 = reg_0598;
    10: op1_02_in14 = reg_0981;
    11: op1_02_in14 = reg_0275;
    12: op1_02_in14 = reg_0661;
    13: op1_02_in14 = reg_0997;
    14: op1_02_in14 = reg_0479;
    15: op1_02_in14 = reg_0573;
    16: op1_02_in14 = reg_0307;
    17: op1_02_in14 = reg_0158;
    18: op1_02_in14 = reg_0088;
    19: op1_02_in14 = reg_0692;
    20: op1_02_in14 = imem03_in[15:12];
    21: op1_02_in14 = reg_0787;
    22: op1_02_in14 = reg_0867;
    29: op1_02_in14 = reg_0867;
    23: op1_02_in14 = reg_0303;
    24: op1_02_in14 = reg_0233;
    25: op1_02_in14 = imem05_in[15:12];
    26: op1_02_in14 = reg_1011;
    27: op1_02_in14 = imem05_in[79:76];
    28: op1_02_in14 = reg_0706;
    30: op1_02_in14 = reg_0977;
    31: op1_02_in14 = reg_0419;
    32: op1_02_in14 = imem02_in[47:44];
    33: op1_02_in14 = imem04_in[7:4];
    34: op1_02_in14 = reg_0283;
    35: op1_02_in14 = reg_0037;
    36: op1_02_in14 = imem01_in[75:72];
    37: op1_02_in14 = reg_0758;
    38: op1_02_in14 = imem04_in[55:52];
    39: op1_02_in14 = reg_0983;
    40: op1_02_in14 = reg_0264;
    41: op1_02_in14 = reg_0821;
    42: op1_02_in14 = reg_0673;
    43: op1_02_in14 = reg_0651;
    44: op1_02_in14 = reg_0888;
    45: op1_02_in14 = reg_0395;
    46: op1_02_in14 = reg_0205;
    47: op1_02_in14 = reg_0998;
    48: op1_02_in14 = reg_0971;
    49: op1_02_in14 = reg_0464;
    50: op1_02_in14 = reg_0670;
    52: op1_02_in14 = reg_0142;
    53: op1_02_in14 = reg_0917;
    54: op1_02_in14 = imem07_in[19:16];
    55: op1_02_in14 = reg_0701;
    56: op1_02_in14 = imem01_in[31:28];
    57: op1_02_in14 = imem02_in[103:100];
    58: op1_02_in14 = reg_0052;
    59: op1_02_in14 = reg_0212;
    60: op1_02_in14 = reg_0055;
    61: op1_02_in14 = reg_0291;
    62: op1_02_in14 = imem04_in[39:36];
    63: op1_02_in14 = imem07_in[95:92];
    65: op1_02_in14 = reg_0481;
    66: op1_02_in14 = reg_0458;
    67: op1_02_in14 = reg_0470;
    68: op1_02_in14 = imem01_in[3:0];
    69: op1_02_in14 = reg_0949;
    70: op1_02_in14 = reg_0169;
    71: op1_02_in14 = reg_0745;
    72: op1_02_in14 = reg_0709;
    73: op1_02_in14 = reg_0452;
    74: op1_02_in14 = reg_0202;
    85: op1_02_in14 = reg_0202;
    75: op1_02_in14 = reg_0896;
    76: op1_02_in14 = imem05_in[55:52];
    77: op1_02_in14 = reg_0802;
    78: op1_02_in14 = reg_0485;
    79: op1_02_in14 = reg_0203;
    80: op1_02_in14 = reg_0199;
    81: op1_02_in14 = reg_0772;
    82: op1_02_in14 = reg_0359;
    83: op1_02_in14 = reg_0569;
    84: op1_02_in14 = reg_0958;
    86: op1_02_in14 = reg_0885;
    89: op1_02_in14 = imem03_in[119:116];
    90: op1_02_in14 = reg_0195;
    92: op1_02_in14 = reg_0476;
    93: op1_02_in14 = reg_0647;
    94: op1_02_in14 = imem05_in[19:16];
    95: op1_02_in14 = reg_0517;
    96: op1_02_in14 = imem05_in[39:36];
    97: op1_02_in14 = reg_0836;
    default: op1_02_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_02_inv14 = 1;
    11: op1_02_inv14 = 1;
    12: op1_02_inv14 = 1;
    13: op1_02_inv14 = 1;
    14: op1_02_inv14 = 1;
    20: op1_02_inv14 = 1;
    21: op1_02_inv14 = 1;
    23: op1_02_inv14 = 1;
    24: op1_02_inv14 = 1;
    26: op1_02_inv14 = 1;
    27: op1_02_inv14 = 1;
    30: op1_02_inv14 = 1;
    31: op1_02_inv14 = 1;
    32: op1_02_inv14 = 1;
    33: op1_02_inv14 = 1;
    34: op1_02_inv14 = 1;
    36: op1_02_inv14 = 1;
    42: op1_02_inv14 = 1;
    43: op1_02_inv14 = 1;
    46: op1_02_inv14 = 1;
    49: op1_02_inv14 = 1;
    50: op1_02_inv14 = 1;
    55: op1_02_inv14 = 1;
    59: op1_02_inv14 = 1;
    60: op1_02_inv14 = 1;
    61: op1_02_inv14 = 1;
    62: op1_02_inv14 = 1;
    63: op1_02_inv14 = 1;
    65: op1_02_inv14 = 1;
    67: op1_02_inv14 = 1;
    70: op1_02_inv14 = 1;
    71: op1_02_inv14 = 1;
    72: op1_02_inv14 = 1;
    75: op1_02_inv14 = 1;
    76: op1_02_inv14 = 1;
    79: op1_02_inv14 = 1;
    81: op1_02_inv14 = 1;
    83: op1_02_inv14 = 1;
    85: op1_02_inv14 = 1;
    90: op1_02_inv14 = 1;
    91: op1_02_inv14 = 1;
    92: op1_02_inv14 = 1;
    94: op1_02_inv14 = 1;
    96: op1_02_inv14 = 1;
    97: op1_02_inv14 = 1;
    default: op1_02_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in15 = reg_0321;
    6: op1_02_in15 = reg_0212;
    7: op1_02_in15 = imem05_in[23:20];
    8: op1_02_in15 = reg_0191;
    9: op1_02_in15 = reg_0586;
    10: op1_02_in15 = reg_0988;
    11: op1_02_in15 = reg_0061;
    12: op1_02_in15 = reg_0643;
    13: op1_02_in15 = imem04_in[103:100];
    14: op1_02_in15 = reg_0478;
    15: op1_02_in15 = reg_0596;
    16: op1_02_in15 = reg_0284;
    18: op1_02_in15 = reg_0081;
    19: op1_02_in15 = reg_0457;
    20: op1_02_in15 = imem03_in[35:32];
    21: op1_02_in15 = reg_1030;
    22: op1_02_in15 = reg_0090;
    37: op1_02_in15 = reg_0090;
    23: op1_02_in15 = reg_0305;
    24: op1_02_in15 = reg_0735;
    25: op1_02_in15 = imem05_in[55:52];
    26: op1_02_in15 = reg_0798;
    27: op1_02_in15 = imem05_in[111:108];
    28: op1_02_in15 = reg_0423;
    31: op1_02_in15 = reg_0423;
    29: op1_02_in15 = reg_0876;
    30: op1_02_in15 = reg_0975;
    32: op1_02_in15 = imem02_in[51:48];
    33: op1_02_in15 = imem04_in[11:8];
    34: op1_02_in15 = imem05_in[11:8];
    35: op1_02_in15 = reg_0085;
    36: op1_02_in15 = reg_0235;
    93: op1_02_in15 = reg_0235;
    38: op1_02_in15 = imem04_in[59:56];
    62: op1_02_in15 = imem04_in[59:56];
    39: op1_02_in15 = imem04_in[23:20];
    40: op1_02_in15 = reg_0804;
    41: op1_02_in15 = reg_0835;
    42: op1_02_in15 = reg_0453;
    43: op1_02_in15 = reg_0647;
    44: op1_02_in15 = reg_0778;
    60: op1_02_in15 = reg_0778;
    45: op1_02_in15 = reg_0351;
    46: op1_02_in15 = reg_0192;
    74: op1_02_in15 = reg_0192;
    47: op1_02_in15 = reg_1001;
    48: op1_02_in15 = reg_0955;
    49: op1_02_in15 = reg_0462;
    50: op1_02_in15 = reg_0677;
    52: op1_02_in15 = reg_0155;
    53: op1_02_in15 = reg_0017;
    54: op1_02_in15 = imem07_in[59:56];
    55: op1_02_in15 = reg_0706;
    56: op1_02_in15 = imem01_in[43:40];
    57: op1_02_in15 = reg_0655;
    58: op1_02_in15 = reg_0248;
    59: op1_02_in15 = imem01_in[15:12];
    61: op1_02_in15 = imem03_in[11:8];
    63: op1_02_in15 = imem07_in[123:120];
    65: op1_02_in15 = reg_0473;
    66: op1_02_in15 = reg_0188;
    67: op1_02_in15 = reg_0452;
    68: op1_02_in15 = imem01_in[47:44];
    69: op1_02_in15 = reg_0945;
    70: op1_02_in15 = reg_0182;
    71: op1_02_in15 = imem02_in[23:20];
    72: op1_02_in15 = reg_0361;
    73: op1_02_in15 = reg_0456;
    75: op1_02_in15 = reg_0082;
    76: op1_02_in15 = imem05_in[59:56];
    77: op1_02_in15 = reg_0850;
    78: op1_02_in15 = reg_0383;
    79: op1_02_in15 = reg_0207;
    80: op1_02_in15 = reg_0197;
    81: op1_02_in15 = reg_0089;
    82: op1_02_in15 = reg_0389;
    83: op1_02_in15 = reg_0708;
    84: op1_02_in15 = reg_0966;
    85: op1_02_in15 = imem01_in[23:20];
    86: op1_02_in15 = reg_0624;
    89: op1_02_in15 = reg_0009;
    90: op1_02_in15 = imem01_in[11:8];
    91: op1_02_in15 = reg_0214;
    92: op1_02_in15 = reg_0475;
    94: op1_02_in15 = imem05_in[35:32];
    95: op1_02_in15 = reg_0108;
    96: op1_02_in15 = imem05_in[47:44];
    97: op1_02_in15 = reg_0301;
    default: op1_02_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv15 = 1;
    7: op1_02_inv15 = 1;
    9: op1_02_inv15 = 1;
    10: op1_02_inv15 = 1;
    12: op1_02_inv15 = 1;
    13: op1_02_inv15 = 1;
    15: op1_02_inv15 = 1;
    16: op1_02_inv15 = 1;
    18: op1_02_inv15 = 1;
    21: op1_02_inv15 = 1;
    23: op1_02_inv15 = 1;
    24: op1_02_inv15 = 1;
    26: op1_02_inv15 = 1;
    27: op1_02_inv15 = 1;
    28: op1_02_inv15 = 1;
    29: op1_02_inv15 = 1;
    30: op1_02_inv15 = 1;
    31: op1_02_inv15 = 1;
    35: op1_02_inv15 = 1;
    36: op1_02_inv15 = 1;
    37: op1_02_inv15 = 1;
    38: op1_02_inv15 = 1;
    40: op1_02_inv15 = 1;
    42: op1_02_inv15 = 1;
    43: op1_02_inv15 = 1;
    45: op1_02_inv15 = 1;
    47: op1_02_inv15 = 1;
    48: op1_02_inv15 = 1;
    50: op1_02_inv15 = 1;
    53: op1_02_inv15 = 1;
    55: op1_02_inv15 = 1;
    56: op1_02_inv15 = 1;
    57: op1_02_inv15 = 1;
    58: op1_02_inv15 = 1;
    62: op1_02_inv15 = 1;
    63: op1_02_inv15 = 1;
    65: op1_02_inv15 = 1;
    68: op1_02_inv15 = 1;
    69: op1_02_inv15 = 1;
    72: op1_02_inv15 = 1;
    75: op1_02_inv15 = 1;
    76: op1_02_inv15 = 1;
    77: op1_02_inv15 = 1;
    79: op1_02_inv15 = 1;
    83: op1_02_inv15 = 1;
    90: op1_02_inv15 = 1;
    94: op1_02_inv15 = 1;
    95: op1_02_inv15 = 1;
    96: op1_02_inv15 = 1;
    97: op1_02_inv15 = 1;
    default: op1_02_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in16 = reg_0343;
    6: op1_02_in16 = imem01_in[27:24];
    85: op1_02_in16 = imem01_in[27:24];
    7: op1_02_in16 = imem05_in[43:40];
    8: op1_02_in16 = imem01_in[19:16];
    9: op1_02_in16 = reg_0571;
    10: op1_02_in16 = reg_0997;
    11: op1_02_in16 = reg_0046;
    12: op1_02_in16 = reg_0665;
    13: op1_02_in16 = imem04_in[115:112];
    14: op1_02_in16 = reg_0204;
    73: op1_02_in16 = reg_0204;
    15: op1_02_in16 = reg_0568;
    16: op1_02_in16 = reg_0054;
    18: op1_02_in16 = reg_0080;
    19: op1_02_in16 = reg_0469;
    42: op1_02_in16 = reg_0469;
    20: op1_02_in16 = imem03_in[47:44];
    61: op1_02_in16 = imem03_in[47:44];
    21: op1_02_in16 = reg_0027;
    22: op1_02_in16 = reg_0484;
    23: op1_02_in16 = reg_0309;
    24: op1_02_in16 = reg_1042;
    25: op1_02_in16 = imem05_in[67:64];
    26: op1_02_in16 = imem07_in[23:20];
    27: op1_02_in16 = imem05_in[115:112];
    28: op1_02_in16 = reg_0442;
    83: op1_02_in16 = reg_0442;
    29: op1_02_in16 = reg_0792;
    30: op1_02_in16 = imem04_in[23:20];
    31: op1_02_in16 = reg_0428;
    32: op1_02_in16 = reg_0653;
    33: op1_02_in16 = imem04_in[31:28];
    34: op1_02_in16 = imem05_in[47:44];
    35: op1_02_in16 = reg_0876;
    36: op1_02_in16 = reg_0779;
    37: op1_02_in16 = reg_0049;
    38: op1_02_in16 = imem04_in[71:68];
    39: op1_02_in16 = imem04_in[71:68];
    40: op1_02_in16 = reg_0390;
    41: op1_02_in16 = reg_0256;
    43: op1_02_in16 = reg_0837;
    44: op1_02_in16 = reg_0058;
    77: op1_02_in16 = reg_0058;
    45: op1_02_in16 = reg_0017;
    46: op1_02_in16 = reg_0197;
    47: op1_02_in16 = reg_0990;
    48: op1_02_in16 = reg_0964;
    49: op1_02_in16 = reg_0481;
    92: op1_02_in16 = reg_0481;
    50: op1_02_in16 = reg_0691;
    52: op1_02_in16 = imem06_in[3:0];
    53: op1_02_in16 = reg_0005;
    54: op1_02_in16 = imem07_in[71:68];
    55: op1_02_in16 = reg_0421;
    72: op1_02_in16 = reg_0421;
    56: op1_02_in16 = imem01_in[59:56];
    57: op1_02_in16 = reg_0654;
    58: op1_02_in16 = reg_0037;
    59: op1_02_in16 = imem01_in[39:36];
    80: op1_02_in16 = imem01_in[39:36];
    60: op1_02_in16 = reg_0931;
    62: op1_02_in16 = imem04_in[67:64];
    63: op1_02_in16 = reg_0726;
    65: op1_02_in16 = reg_0471;
    66: op1_02_in16 = imem01_in[83:80];
    68: op1_02_in16 = imem01_in[83:80];
    67: op1_02_in16 = reg_0200;
    69: op1_02_in16 = reg_0953;
    70: op1_02_in16 = reg_0173;
    71: op1_02_in16 = imem02_in[39:36];
    74: op1_02_in16 = imem01_in[23:20];
    75: op1_02_in16 = reg_0098;
    76: op1_02_in16 = imem05_in[71:68];
    78: op1_02_in16 = reg_0369;
    79: op1_02_in16 = reg_0198;
    81: op1_02_in16 = reg_0776;
    82: op1_02_in16 = reg_0425;
    84: op1_02_in16 = reg_0948;
    86: op1_02_in16 = reg_0493;
    89: op1_02_in16 = reg_0758;
    90: op1_02_in16 = imem01_in[47:44];
    91: op1_02_in16 = reg_0207;
    93: op1_02_in16 = reg_0140;
    94: op1_02_in16 = imem05_in[55:52];
    95: op1_02_in16 = reg_0071;
    96: op1_02_in16 = imem05_in[59:56];
    97: op1_02_in16 = reg_0062;
    default: op1_02_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv16 = 1;
    7: op1_02_inv16 = 1;
    8: op1_02_inv16 = 1;
    10: op1_02_inv16 = 1;
    11: op1_02_inv16 = 1;
    12: op1_02_inv16 = 1;
    13: op1_02_inv16 = 1;
    16: op1_02_inv16 = 1;
    18: op1_02_inv16 = 1;
    19: op1_02_inv16 = 1;
    24: op1_02_inv16 = 1;
    27: op1_02_inv16 = 1;
    28: op1_02_inv16 = 1;
    31: op1_02_inv16 = 1;
    32: op1_02_inv16 = 1;
    35: op1_02_inv16 = 1;
    36: op1_02_inv16 = 1;
    39: op1_02_inv16 = 1;
    41: op1_02_inv16 = 1;
    42: op1_02_inv16 = 1;
    43: op1_02_inv16 = 1;
    47: op1_02_inv16 = 1;
    56: op1_02_inv16 = 1;
    59: op1_02_inv16 = 1;
    60: op1_02_inv16 = 1;
    61: op1_02_inv16 = 1;
    66: op1_02_inv16 = 1;
    69: op1_02_inv16 = 1;
    72: op1_02_inv16 = 1;
    73: op1_02_inv16 = 1;
    76: op1_02_inv16 = 1;
    77: op1_02_inv16 = 1;
    79: op1_02_inv16 = 1;
    80: op1_02_inv16 = 1;
    84: op1_02_inv16 = 1;
    85: op1_02_inv16 = 1;
    86: op1_02_inv16 = 1;
    91: op1_02_inv16 = 1;
    92: op1_02_inv16 = 1;
    93: op1_02_inv16 = 1;
    95: op1_02_inv16 = 1;
    97: op1_02_inv16 = 1;
    default: op1_02_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in17 = reg_0331;
    6: op1_02_in17 = imem01_in[59:56];
    7: op1_02_in17 = imem05_in[47:44];
    8: op1_02_in17 = imem01_in[35:32];
    9: op1_02_in17 = reg_0599;
    10: op1_02_in17 = reg_0994;
    11: op1_02_in17 = reg_0078;
    12: op1_02_in17 = reg_0659;
    13: op1_02_in17 = imem04_in[127:124];
    14: op1_02_in17 = reg_0212;
    15: op1_02_in17 = reg_0591;
    16: op1_02_in17 = reg_0056;
    18: op1_02_in17 = reg_0082;
    19: op1_02_in17 = reg_0462;
    20: op1_02_in17 = imem03_in[71:68];
    21: op1_02_in17 = reg_0781;
    22: op1_02_in17 = reg_0291;
    37: op1_02_in17 = reg_0291;
    23: op1_02_in17 = reg_0060;
    24: op1_02_in17 = reg_1031;
    25: op1_02_in17 = imem05_in[75:72];
    26: op1_02_in17 = imem07_in[79:76];
    27: op1_02_in17 = reg_0963;
    69: op1_02_in17 = reg_0963;
    28: op1_02_in17 = reg_0420;
    29: op1_02_in17 = reg_0814;
    30: op1_02_in17 = imem04_in[63:60];
    31: op1_02_in17 = reg_0172;
    32: op1_02_in17 = reg_0637;
    33: op1_02_in17 = imem04_in[71:68];
    34: op1_02_in17 = imem05_in[67:64];
    35: op1_02_in17 = reg_0091;
    36: op1_02_in17 = reg_0560;
    38: op1_02_in17 = imem04_in[95:92];
    39: op1_02_in17 = imem04_in[75:72];
    40: op1_02_in17 = reg_0332;
    41: op1_02_in17 = reg_0827;
    42: op1_02_in17 = reg_0466;
    43: op1_02_in17 = reg_0097;
    44: op1_02_in17 = reg_0066;
    45: op1_02_in17 = reg_0596;
    46: op1_02_in17 = imem01_in[23:20];
    47: op1_02_in17 = imem04_in[7:4];
    48: op1_02_in17 = reg_0965;
    49: op1_02_in17 = reg_0198;
    50: op1_02_in17 = reg_0674;
    52: op1_02_in17 = imem06_in[47:44];
    53: op1_02_in17 = imem07_in[27:24];
    54: op1_02_in17 = reg_0722;
    55: op1_02_in17 = reg_0175;
    56: op1_02_in17 = imem01_in[75:72];
    57: op1_02_in17 = reg_0300;
    58: op1_02_in17 = reg_0335;
    59: op1_02_in17 = imem01_in[47:44];
    60: op1_02_in17 = reg_0541;
    61: op1_02_in17 = imem03_in[119:116];
    62: op1_02_in17 = imem04_in[99:96];
    63: op1_02_in17 = reg_0729;
    65: op1_02_in17 = reg_0479;
    66: op1_02_in17 = imem01_in[107:104];
    67: op1_02_in17 = reg_0204;
    68: op1_02_in17 = imem01_in[95:92];
    70: op1_02_in17 = reg_0171;
    71: op1_02_in17 = imem02_in[55:52];
    72: op1_02_in17 = reg_0426;
    73: op1_02_in17 = reg_0193;
    74: op1_02_in17 = imem01_in[31:28];
    75: op1_02_in17 = reg_0783;
    76: op1_02_in17 = imem05_in[87:84];
    77: op1_02_in17 = reg_0808;
    78: op1_02_in17 = imem07_in[3:0];
    79: op1_02_in17 = reg_0201;
    80: op1_02_in17 = imem01_in[67:64];
    81: op1_02_in17 = reg_0876;
    82: op1_02_in17 = reg_0248;
    83: op1_02_in17 = reg_0759;
    84: op1_02_in17 = reg_0892;
    85: op1_02_in17 = imem01_in[71:68];
    86: op1_02_in17 = imem03_in[11:8];
    89: op1_02_in17 = reg_0761;
    90: op1_02_in17 = imem01_in[79:76];
    91: op1_02_in17 = imem01_in[103:100];
    92: op1_02_in17 = reg_0191;
    93: op1_02_in17 = reg_0648;
    94: op1_02_in17 = imem05_in[59:56];
    95: op1_02_in17 = reg_0824;
    96: op1_02_in17 = imem05_in[63:60];
    97: op1_02_in17 = reg_0823;
    default: op1_02_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_02_inv17 = 1;
    8: op1_02_inv17 = 1;
    10: op1_02_inv17 = 1;
    11: op1_02_inv17 = 1;
    21: op1_02_inv17 = 1;
    22: op1_02_inv17 = 1;
    25: op1_02_inv17 = 1;
    27: op1_02_inv17 = 1;
    28: op1_02_inv17 = 1;
    30: op1_02_inv17 = 1;
    35: op1_02_inv17 = 1;
    36: op1_02_inv17 = 1;
    38: op1_02_inv17 = 1;
    39: op1_02_inv17 = 1;
    40: op1_02_inv17 = 1;
    41: op1_02_inv17 = 1;
    44: op1_02_inv17 = 1;
    45: op1_02_inv17 = 1;
    46: op1_02_inv17 = 1;
    47: op1_02_inv17 = 1;
    48: op1_02_inv17 = 1;
    49: op1_02_inv17 = 1;
    50: op1_02_inv17 = 1;
    53: op1_02_inv17 = 1;
    58: op1_02_inv17 = 1;
    59: op1_02_inv17 = 1;
    60: op1_02_inv17 = 1;
    62: op1_02_inv17 = 1;
    63: op1_02_inv17 = 1;
    67: op1_02_inv17 = 1;
    69: op1_02_inv17 = 1;
    71: op1_02_inv17 = 1;
    73: op1_02_inv17 = 1;
    76: op1_02_inv17 = 1;
    78: op1_02_inv17 = 1;
    81: op1_02_inv17 = 1;
    82: op1_02_inv17 = 1;
    83: op1_02_inv17 = 1;
    84: op1_02_inv17 = 1;
    89: op1_02_inv17 = 1;
    90: op1_02_inv17 = 1;
    91: op1_02_inv17 = 1;
    93: op1_02_inv17 = 1;
    94: op1_02_inv17 = 1;
    95: op1_02_inv17 = 1;
    97: op1_02_inv17 = 1;
    default: op1_02_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in18 = reg_0000;
    6: op1_02_in18 = imem01_in[103:100];
    7: op1_02_in18 = imem05_in[59:56];
    8: op1_02_in18 = imem01_in[43:40];
    9: op1_02_in18 = reg_0591;
    10: op1_02_in18 = imem04_in[79:76];
    11: op1_02_in18 = reg_0062;
    12: op1_02_in18 = reg_0333;
    13: op1_02_in18 = reg_0545;
    14: op1_02_in18 = reg_0197;
    15: op1_02_in18 = reg_0594;
    16: op1_02_in18 = reg_0053;
    18: op1_02_in18 = imem03_in[23:20];
    86: op1_02_in18 = imem03_in[23:20];
    19: op1_02_in18 = reg_0472;
    42: op1_02_in18 = reg_0472;
    20: op1_02_in18 = imem03_in[79:76];
    21: op1_02_in18 = reg_0805;
    22: op1_02_in18 = imem03_in[31:28];
    23: op1_02_in18 = reg_0764;
    24: op1_02_in18 = reg_1038;
    25: op1_02_in18 = imem05_in[111:108];
    26: op1_02_in18 = reg_0719;
    54: op1_02_in18 = reg_0719;
    27: op1_02_in18 = reg_0973;
    28: op1_02_in18 = reg_0431;
    29: op1_02_in18 = imem03_in[3:0];
    30: op1_02_in18 = imem04_in[107:104];
    31: op1_02_in18 = reg_0157;
    32: op1_02_in18 = reg_0659;
    33: op1_02_in18 = imem04_in[95:92];
    34: op1_02_in18 = imem05_in[71:68];
    35: op1_02_in18 = imem03_in[91:88];
    36: op1_02_in18 = reg_0218;
    37: op1_02_in18 = imem03_in[87:84];
    38: op1_02_in18 = imem04_in[111:108];
    39: op1_02_in18 = imem04_in[99:96];
    40: op1_02_in18 = reg_0780;
    41: op1_02_in18 = reg_0260;
    43: op1_02_in18 = reg_0339;
    44: op1_02_in18 = reg_0056;
    45: op1_02_in18 = reg_0029;
    46: op1_02_in18 = imem01_in[63:60];
    47: op1_02_in18 = imem04_in[11:8];
    48: op1_02_in18 = reg_0947;
    49: op1_02_in18 = reg_0190;
    50: op1_02_in18 = reg_0671;
    52: op1_02_in18 = imem06_in[71:68];
    53: op1_02_in18 = imem07_in[43:40];
    55: op1_02_in18 = reg_0172;
    56: op1_02_in18 = imem01_in[87:84];
    57: op1_02_in18 = reg_0081;
    58: op1_02_in18 = reg_0089;
    59: op1_02_in18 = imem01_in[127:124];
    60: op1_02_in18 = reg_0507;
    61: op1_02_in18 = reg_0099;
    62: op1_02_in18 = imem04_in[119:116];
    63: op1_02_in18 = reg_0002;
    65: op1_02_in18 = reg_0210;
    66: op1_02_in18 = reg_0242;
    67: op1_02_in18 = reg_0188;
    68: op1_02_in18 = reg_0779;
    69: op1_02_in18 = reg_0255;
    71: op1_02_in18 = imem02_in[79:76];
    72: op1_02_in18 = reg_0315;
    73: op1_02_in18 = reg_0194;
    74: op1_02_in18 = imem01_in[83:80];
    75: op1_02_in18 = reg_0423;
    76: op1_02_in18 = reg_0866;
    77: op1_02_in18 = reg_0444;
    78: op1_02_in18 = imem07_in[11:8];
    79: op1_02_in18 = imem01_in[23:20];
    80: op1_02_in18 = imem01_in[95:92];
    81: op1_02_in18 = reg_0884;
    82: op1_02_in18 = reg_0608;
    83: op1_02_in18 = reg_0727;
    84: op1_02_in18 = reg_0336;
    85: op1_02_in18 = imem01_in[79:76];
    89: op1_02_in18 = reg_0578;
    90: op1_02_in18 = imem01_in[99:96];
    91: op1_02_in18 = reg_1042;
    92: op1_02_in18 = reg_0199;
    93: op1_02_in18 = reg_0057;
    94: op1_02_in18 = imem05_in[107:104];
    95: op1_02_in18 = imem05_in[15:12];
    96: op1_02_in18 = imem05_in[67:64];
    97: op1_02_in18 = reg_0278;
    default: op1_02_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv18 = 1;
    6: op1_02_inv18 = 1;
    7: op1_02_inv18 = 1;
    8: op1_02_inv18 = 1;
    9: op1_02_inv18 = 1;
    10: op1_02_inv18 = 1;
    12: op1_02_inv18 = 1;
    13: op1_02_inv18 = 1;
    16: op1_02_inv18 = 1;
    19: op1_02_inv18 = 1;
    21: op1_02_inv18 = 1;
    22: op1_02_inv18 = 1;
    23: op1_02_inv18 = 1;
    26: op1_02_inv18 = 1;
    27: op1_02_inv18 = 1;
    29: op1_02_inv18 = 1;
    30: op1_02_inv18 = 1;
    31: op1_02_inv18 = 1;
    32: op1_02_inv18 = 1;
    33: op1_02_inv18 = 1;
    35: op1_02_inv18 = 1;
    36: op1_02_inv18 = 1;
    37: op1_02_inv18 = 1;
    38: op1_02_inv18 = 1;
    39: op1_02_inv18 = 1;
    40: op1_02_inv18 = 1;
    41: op1_02_inv18 = 1;
    42: op1_02_inv18 = 1;
    43: op1_02_inv18 = 1;
    47: op1_02_inv18 = 1;
    49: op1_02_inv18 = 1;
    54: op1_02_inv18 = 1;
    55: op1_02_inv18 = 1;
    58: op1_02_inv18 = 1;
    60: op1_02_inv18 = 1;
    61: op1_02_inv18 = 1;
    62: op1_02_inv18 = 1;
    66: op1_02_inv18 = 1;
    67: op1_02_inv18 = 1;
    68: op1_02_inv18 = 1;
    69: op1_02_inv18 = 1;
    73: op1_02_inv18 = 1;
    75: op1_02_inv18 = 1;
    77: op1_02_inv18 = 1;
    82: op1_02_inv18 = 1;
    83: op1_02_inv18 = 1;
    84: op1_02_inv18 = 1;
    85: op1_02_inv18 = 1;
    86: op1_02_inv18 = 1;
    89: op1_02_inv18 = 1;
    90: op1_02_inv18 = 1;
    91: op1_02_inv18 = 1;
    92: op1_02_inv18 = 1;
    93: op1_02_inv18 = 1;
    95: op1_02_inv18 = 1;
    default: op1_02_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in19 = reg_0001;
    6: op1_02_in19 = reg_0496;
    7: op1_02_in19 = imem05_in[79:76];
    8: op1_02_in19 = imem01_in[51:48];
    9: op1_02_in19 = reg_0589;
    10: op1_02_in19 = imem04_in[87:84];
    11: op1_02_in19 = reg_0065;
    12: op1_02_in19 = reg_0359;
    57: op1_02_in19 = reg_0359;
    13: op1_02_in19 = reg_0532;
    14: op1_02_in19 = imem01_in[11:8];
    15: op1_02_in19 = reg_0576;
    16: op1_02_in19 = reg_0063;
    18: op1_02_in19 = imem03_in[31:28];
    19: op1_02_in19 = reg_0214;
    20: op1_02_in19 = reg_0598;
    21: op1_02_in19 = reg_0011;
    22: op1_02_in19 = imem03_in[43:40];
    23: op1_02_in19 = reg_0078;
    24: op1_02_in19 = reg_0122;
    25: op1_02_in19 = reg_0962;
    26: op1_02_in19 = reg_0730;
    27: op1_02_in19 = reg_0966;
    28: op1_02_in19 = reg_0172;
    29: op1_02_in19 = imem03_in[51:48];
    30: op1_02_in19 = imem04_in[127:124];
    31: op1_02_in19 = reg_0171;
    32: op1_02_in19 = reg_0663;
    33: op1_02_in19 = imem04_in[107:104];
    34: op1_02_in19 = reg_0958;
    35: op1_02_in19 = imem03_in[103:100];
    36: op1_02_in19 = reg_0240;
    37: op1_02_in19 = imem03_in[111:108];
    38: op1_02_in19 = reg_1004;
    39: op1_02_in19 = imem04_in[103:100];
    40: op1_02_in19 = reg_0025;
    41: op1_02_in19 = reg_0896;
    42: op1_02_in19 = reg_0480;
    43: op1_02_in19 = reg_0865;
    44: op1_02_in19 = reg_0584;
    45: op1_02_in19 = imem07_in[3:0];
    46: op1_02_in19 = reg_0828;
    47: op1_02_in19 = imem04_in[71:68];
    48: op1_02_in19 = reg_0900;
    49: op1_02_in19 = imem01_in[23:20];
    50: op1_02_in19 = reg_0463;
    52: op1_02_in19 = imem06_in[119:116];
    53: op1_02_in19 = imem07_in[47:44];
    54: op1_02_in19 = reg_0744;
    55: op1_02_in19 = reg_0163;
    56: op1_02_in19 = imem01_in[95:92];
    58: op1_02_in19 = reg_0876;
    59: op1_02_in19 = reg_0786;
    60: op1_02_in19 = reg_0276;
    61: op1_02_in19 = reg_0445;
    62: op1_02_in19 = imem04_in[123:120];
    63: op1_02_in19 = reg_0433;
    65: op1_02_in19 = reg_0198;
    66: op1_02_in19 = reg_1056;
    67: op1_02_in19 = reg_0207;
    68: op1_02_in19 = reg_0928;
    69: op1_02_in19 = reg_0274;
    71: op1_02_in19 = imem02_in[119:116];
    72: op1_02_in19 = reg_0167;
    73: op1_02_in19 = reg_0213;
    74: op1_02_in19 = imem01_in[107:104];
    75: op1_02_in19 = reg_0516;
    76: op1_02_in19 = reg_0142;
    77: op1_02_in19 = reg_0295;
    78: op1_02_in19 = imem07_in[15:12];
    79: op1_02_in19 = imem01_in[27:24];
    80: op1_02_in19 = reg_0973;
    81: op1_02_in19 = imem03_in[7:4];
    82: op1_02_in19 = reg_0335;
    83: op1_02_in19 = reg_0361;
    84: op1_02_in19 = reg_0223;
    85: op1_02_in19 = imem01_in[115:112];
    86: op1_02_in19 = imem03_in[63:60];
    89: op1_02_in19 = reg_0596;
    97: op1_02_in19 = reg_0596;
    90: op1_02_in19 = reg_0969;
    91: op1_02_in19 = reg_1044;
    92: op1_02_in19 = imem01_in[19:16];
    93: op1_02_in19 = reg_0268;
    94: op1_02_in19 = reg_0866;
    95: op1_02_in19 = imem05_in[39:36];
    96: op1_02_in19 = imem05_in[103:100];
    default: op1_02_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv19 = 1;
    7: op1_02_inv19 = 1;
    9: op1_02_inv19 = 1;
    10: op1_02_inv19 = 1;
    15: op1_02_inv19 = 1;
    16: op1_02_inv19 = 1;
    21: op1_02_inv19 = 1;
    23: op1_02_inv19 = 1;
    24: op1_02_inv19 = 1;
    26: op1_02_inv19 = 1;
    29: op1_02_inv19 = 1;
    33: op1_02_inv19 = 1;
    34: op1_02_inv19 = 1;
    36: op1_02_inv19 = 1;
    37: op1_02_inv19 = 1;
    40: op1_02_inv19 = 1;
    42: op1_02_inv19 = 1;
    43: op1_02_inv19 = 1;
    46: op1_02_inv19 = 1;
    56: op1_02_inv19 = 1;
    58: op1_02_inv19 = 1;
    59: op1_02_inv19 = 1;
    60: op1_02_inv19 = 1;
    61: op1_02_inv19 = 1;
    63: op1_02_inv19 = 1;
    65: op1_02_inv19 = 1;
    69: op1_02_inv19 = 1;
    73: op1_02_inv19 = 1;
    76: op1_02_inv19 = 1;
    78: op1_02_inv19 = 1;
    79: op1_02_inv19 = 1;
    83: op1_02_inv19 = 1;
    84: op1_02_inv19 = 1;
    85: op1_02_inv19 = 1;
    86: op1_02_inv19 = 1;
    91: op1_02_inv19 = 1;
    93: op1_02_inv19 = 1;
    95: op1_02_inv19 = 1;
    default: op1_02_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in20 = reg_0002;
    6: op1_02_in20 = reg_0513;
    7: op1_02_in20 = imem05_in[115:112];
    8: op1_02_in20 = reg_0504;
    9: op1_02_in20 = reg_0594;
    10: op1_02_in20 = imem04_in[111:108];
    11: op1_02_in20 = reg_0058;
    12: op1_02_in20 = reg_0363;
    13: op1_02_in20 = reg_0301;
    14: op1_02_in20 = imem01_in[15:12];
    15: op1_02_in20 = reg_0384;
    16: op1_02_in20 = reg_0074;
    18: op1_02_in20 = imem03_in[63:60];
    19: op1_02_in20 = reg_0210;
    20: op1_02_in20 = reg_0579;
    21: op1_02_in20 = reg_0798;
    22: op1_02_in20 = imem03_in[47:44];
    23: op1_02_in20 = reg_0014;
    24: op1_02_in20 = reg_0124;
    25: op1_02_in20 = reg_0973;
    26: op1_02_in20 = reg_0721;
    27: op1_02_in20 = reg_0951;
    28: op1_02_in20 = reg_0169;
    29: op1_02_in20 = imem03_in[111:108];
    35: op1_02_in20 = imem03_in[111:108];
    30: op1_02_in20 = reg_0282;
    32: op1_02_in20 = reg_0863;
    33: op1_02_in20 = imem04_in[119:116];
    34: op1_02_in20 = reg_0948;
    36: op1_02_in20 = reg_0122;
    74: op1_02_in20 = reg_0122;
    37: op1_02_in20 = reg_0571;
    38: op1_02_in20 = reg_0536;
    39: op1_02_in20 = imem04_in[123:120];
    40: op1_02_in20 = reg_1010;
    41: op1_02_in20 = reg_0819;
    42: op1_02_in20 = reg_0468;
    43: op1_02_in20 = reg_0335;
    44: op1_02_in20 = reg_0401;
    45: op1_02_in20 = imem07_in[43:40];
    46: op1_02_in20 = reg_0604;
    47: op1_02_in20 = imem04_in[83:80];
    48: op1_02_in20 = reg_0827;
    49: op1_02_in20 = imem01_in[47:44];
    50: op1_02_in20 = reg_0450;
    52: op1_02_in20 = imem06_in[127:124];
    53: op1_02_in20 = imem07_in[87:84];
    54: op1_02_in20 = reg_0428;
    55: op1_02_in20 = reg_0177;
    56: op1_02_in20 = imem01_in[99:96];
    57: op1_02_in20 = reg_0248;
    58: op1_02_in20 = reg_0484;
    59: op1_02_in20 = reg_0904;
    60: op1_02_in20 = reg_0288;
    61: op1_02_in20 = reg_0240;
    62: op1_02_in20 = reg_0483;
    63: op1_02_in20 = reg_0321;
    83: op1_02_in20 = reg_0321;
    65: op1_02_in20 = reg_0196;
    66: op1_02_in20 = reg_0592;
    67: op1_02_in20 = reg_0212;
    73: op1_02_in20 = reg_0212;
    68: op1_02_in20 = reg_0933;
    69: op1_02_in20 = reg_0688;
    71: op1_02_in20 = reg_0845;
    72: op1_02_in20 = reg_0159;
    75: op1_02_in20 = reg_0758;
    76: op1_02_in20 = reg_0143;
    77: op1_02_in20 = reg_0531;
    78: op1_02_in20 = imem07_in[51:48];
    79: op1_02_in20 = imem01_in[31:28];
    80: op1_02_in20 = reg_0337;
    81: op1_02_in20 = imem03_in[55:52];
    82: op1_02_in20 = reg_0516;
    84: op1_02_in20 = reg_0153;
    85: op1_02_in20 = imem01_in[123:120];
    86: op1_02_in20 = imem03_in[71:68];
    89: op1_02_in20 = reg_0239;
    90: op1_02_in20 = reg_0971;
    91: op1_02_in20 = reg_1035;
    92: op1_02_in20 = reg_0106;
    93: op1_02_in20 = reg_0178;
    94: op1_02_in20 = reg_0492;
    95: op1_02_in20 = imem05_in[59:56];
    96: op1_02_in20 = reg_0215;
    97: op1_02_in20 = reg_0597;
    default: op1_02_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_02_inv20 = 1;
    8: op1_02_inv20 = 1;
    9: op1_02_inv20 = 1;
    10: op1_02_inv20 = 1;
    11: op1_02_inv20 = 1;
    12: op1_02_inv20 = 1;
    18: op1_02_inv20 = 1;
    19: op1_02_inv20 = 1;
    20: op1_02_inv20 = 1;
    21: op1_02_inv20 = 1;
    22: op1_02_inv20 = 1;
    23: op1_02_inv20 = 1;
    28: op1_02_inv20 = 1;
    33: op1_02_inv20 = 1;
    34: op1_02_inv20 = 1;
    36: op1_02_inv20 = 1;
    37: op1_02_inv20 = 1;
    38: op1_02_inv20 = 1;
    41: op1_02_inv20 = 1;
    42: op1_02_inv20 = 1;
    43: op1_02_inv20 = 1;
    44: op1_02_inv20 = 1;
    46: op1_02_inv20 = 1;
    50: op1_02_inv20 = 1;
    56: op1_02_inv20 = 1;
    58: op1_02_inv20 = 1;
    60: op1_02_inv20 = 1;
    63: op1_02_inv20 = 1;
    65: op1_02_inv20 = 1;
    72: op1_02_inv20 = 1;
    80: op1_02_inv20 = 1;
    81: op1_02_inv20 = 1;
    82: op1_02_inv20 = 1;
    85: op1_02_inv20 = 1;
    90: op1_02_inv20 = 1;
    91: op1_02_inv20 = 1;
    92: op1_02_inv20 = 1;
    94: op1_02_inv20 = 1;
    95: op1_02_inv20 = 1;
    96: op1_02_inv20 = 1;
    default: op1_02_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in21 = reg_0003;
    6: op1_02_in21 = reg_0499;
    7: op1_02_in21 = imem05_in[119:116];
    8: op1_02_in21 = reg_0501;
    9: op1_02_in21 = reg_0600;
    10: op1_02_in21 = reg_0544;
    11: op1_02_in21 = reg_0074;
    12: op1_02_in21 = reg_0353;
    13: op1_02_in21 = reg_0283;
    14: op1_02_in21 = imem01_in[27:24];
    73: op1_02_in21 = imem01_in[27:24];
    15: op1_02_in21 = reg_0387;
    16: op1_02_in21 = imem05_in[15:12];
    18: op1_02_in21 = imem03_in[99:96];
    19: op1_02_in21 = reg_0209;
    20: op1_02_in21 = reg_0568;
    21: op1_02_in21 = imem07_in[7:4];
    22: op1_02_in21 = imem03_in[51:48];
    23: op1_02_in21 = reg_0075;
    24: op1_02_in21 = reg_0118;
    25: op1_02_in21 = reg_0954;
    26: op1_02_in21 = reg_0726;
    27: op1_02_in21 = reg_0968;
    28: op1_02_in21 = reg_0166;
    29: op1_02_in21 = reg_0579;
    30: op1_02_in21 = reg_1005;
    32: op1_02_in21 = reg_0096;
    33: op1_02_in21 = reg_0511;
    38: op1_02_in21 = reg_0511;
    34: op1_02_in21 = reg_0942;
    35: op1_02_in21 = reg_0394;
    36: op1_02_in21 = reg_0103;
    46: op1_02_in21 = reg_0103;
    37: op1_02_in21 = reg_0046;
    39: op1_02_in21 = imem04_in[127:124];
    40: op1_02_in21 = reg_0008;
    41: op1_02_in21 = reg_0831;
    42: op1_02_in21 = reg_0191;
    43: op1_02_in21 = reg_0083;
    44: op1_02_in21 = reg_0015;
    45: op1_02_in21 = imem07_in[47:44];
    47: op1_02_in21 = imem04_in[99:96];
    48: op1_02_in21 = reg_0491;
    49: op1_02_in21 = imem01_in[111:108];
    50: op1_02_in21 = reg_0457;
    52: op1_02_in21 = reg_0614;
    53: op1_02_in21 = imem07_in[119:116];
    54: op1_02_in21 = reg_0599;
    55: op1_02_in21 = reg_0170;
    56: op1_02_in21 = imem01_in[103:100];
    57: op1_02_in21 = reg_0331;
    58: op1_02_in21 = reg_0291;
    59: op1_02_in21 = reg_1052;
    60: op1_02_in21 = reg_0552;
    61: op1_02_in21 = reg_0784;
    62: op1_02_in21 = reg_0306;
    63: op1_02_in21 = reg_0744;
    65: op1_02_in21 = reg_0205;
    66: op1_02_in21 = reg_0253;
    67: op1_02_in21 = imem01_in[59:56];
    68: op1_02_in21 = reg_0870;
    69: op1_02_in21 = reg_0221;
    71: op1_02_in21 = reg_0036;
    72: op1_02_in21 = reg_0169;
    74: op1_02_in21 = reg_0337;
    75: op1_02_in21 = reg_0089;
    76: op1_02_in21 = reg_0275;
    94: op1_02_in21 = reg_0275;
    77: op1_02_in21 = imem05_in[95:92];
    78: op1_02_in21 = imem07_in[91:88];
    79: op1_02_in21 = imem01_in[47:44];
    80: op1_02_in21 = reg_1035;
    81: op1_02_in21 = imem03_in[103:100];
    82: op1_02_in21 = reg_0347;
    83: op1_02_in21 = reg_0406;
    84: op1_02_in21 = reg_0148;
    85: op1_02_in21 = reg_0105;
    86: op1_02_in21 = imem03_in[107:104];
    89: op1_02_in21 = reg_0230;
    90: op1_02_in21 = reg_1056;
    91: op1_02_in21 = reg_0503;
    92: op1_02_in21 = reg_1032;
    93: op1_02_in21 = reg_0063;
    95: op1_02_in21 = imem05_in[87:84];
    96: op1_02_in21 = reg_0217;
    97: op1_02_in21 = reg_0385;
    default: op1_02_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv21 = 1;
    6: op1_02_inv21 = 1;
    7: op1_02_inv21 = 1;
    8: op1_02_inv21 = 1;
    9: op1_02_inv21 = 1;
    10: op1_02_inv21 = 1;
    12: op1_02_inv21 = 1;
    13: op1_02_inv21 = 1;
    14: op1_02_inv21 = 1;
    16: op1_02_inv21 = 1;
    18: op1_02_inv21 = 1;
    19: op1_02_inv21 = 1;
    20: op1_02_inv21 = 1;
    21: op1_02_inv21 = 1;
    26: op1_02_inv21 = 1;
    29: op1_02_inv21 = 1;
    32: op1_02_inv21 = 1;
    33: op1_02_inv21 = 1;
    36: op1_02_inv21 = 1;
    40: op1_02_inv21 = 1;
    42: op1_02_inv21 = 1;
    48: op1_02_inv21 = 1;
    49: op1_02_inv21 = 1;
    52: op1_02_inv21 = 1;
    54: op1_02_inv21 = 1;
    55: op1_02_inv21 = 1;
    58: op1_02_inv21 = 1;
    61: op1_02_inv21 = 1;
    62: op1_02_inv21 = 1;
    69: op1_02_inv21 = 1;
    71: op1_02_inv21 = 1;
    72: op1_02_inv21 = 1;
    75: op1_02_inv21 = 1;
    78: op1_02_inv21 = 1;
    79: op1_02_inv21 = 1;
    80: op1_02_inv21 = 1;
    84: op1_02_inv21 = 1;
    86: op1_02_inv21 = 1;
    89: op1_02_inv21 = 1;
    91: op1_02_inv21 = 1;
    92: op1_02_inv21 = 1;
    95: op1_02_inv21 = 1;
    97: op1_02_inv21 = 1;
    default: op1_02_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in22 = reg_0004;
    69: op1_02_in22 = reg_0004;
    6: op1_02_in22 = reg_0518;
    91: op1_02_in22 = reg_0518;
    7: op1_02_in22 = reg_0963;
    8: op1_02_in22 = reg_0500;
    9: op1_02_in22 = reg_0595;
    10: op1_02_in22 = reg_0545;
    11: op1_02_in22 = reg_0044;
    12: op1_02_in22 = reg_0355;
    13: op1_02_in22 = reg_0294;
    14: op1_02_in22 = imem01_in[95:92];
    15: op1_02_in22 = reg_0321;
    16: op1_02_in22 = imem05_in[19:16];
    18: op1_02_in22 = reg_0596;
    19: op1_02_in22 = reg_0186;
    20: op1_02_in22 = reg_0569;
    21: op1_02_in22 = imem07_in[19:16];
    22: op1_02_in22 = imem03_in[67:64];
    23: op1_02_in22 = reg_0074;
    24: op1_02_in22 = reg_0125;
    25: op1_02_in22 = reg_0900;
    26: op1_02_in22 = reg_0729;
    27: op1_02_in22 = reg_0945;
    29: op1_02_in22 = reg_0580;
    37: op1_02_in22 = reg_0580;
    30: op1_02_in22 = reg_0292;
    32: op1_02_in22 = reg_0330;
    33: op1_02_in22 = reg_0937;
    34: op1_02_in22 = reg_0835;
    35: op1_02_in22 = reg_0938;
    36: op1_02_in22 = reg_0108;
    38: op1_02_in22 = reg_0048;
    39: op1_02_in22 = reg_1004;
    40: op1_02_in22 = imem07_in[99:96];
    41: op1_02_in22 = reg_0132;
    42: op1_02_in22 = reg_0187;
    43: op1_02_in22 = reg_0088;
    44: op1_02_in22 = reg_0296;
    45: op1_02_in22 = imem07_in[95:92];
    78: op1_02_in22 = imem07_in[95:92];
    46: op1_02_in22 = reg_0111;
    47: op1_02_in22 = imem04_in[123:120];
    48: op1_02_in22 = reg_0832;
    49: op1_02_in22 = reg_0830;
    50: op1_02_in22 = reg_0469;
    52: op1_02_in22 = reg_0624;
    53: op1_02_in22 = reg_0718;
    54: op1_02_in22 = reg_0420;
    63: op1_02_in22 = reg_0420;
    56: op1_02_in22 = imem01_in[111:108];
    57: op1_02_in22 = reg_0347;
    58: op1_02_in22 = imem03_in[31:28];
    59: op1_02_in22 = reg_0249;
    60: op1_02_in22 = reg_0824;
    61: op1_02_in22 = reg_0509;
    62: op1_02_in22 = reg_0537;
    65: op1_02_in22 = reg_0199;
    66: op1_02_in22 = reg_0520;
    67: op1_02_in22 = imem01_in[91:88];
    68: op1_02_in22 = reg_1036;
    71: op1_02_in22 = reg_0224;
    72: op1_02_in22 = reg_0160;
    73: op1_02_in22 = imem01_in[47:44];
    74: op1_02_in22 = reg_0488;
    80: op1_02_in22 = reg_0488;
    90: op1_02_in22 = reg_0488;
    75: op1_02_in22 = reg_0761;
    76: op1_02_in22 = reg_0689;
    94: op1_02_in22 = reg_0689;
    77: op1_02_in22 = imem05_in[111:108];
    79: op1_02_in22 = imem01_in[67:64];
    81: op1_02_in22 = imem03_in[119:116];
    82: op1_02_in22 = reg_0772;
    83: op1_02_in22 = reg_0641;
    84: op1_02_in22 = reg_0404;
    85: op1_02_in22 = reg_1042;
    86: op1_02_in22 = reg_0012;
    89: op1_02_in22 = reg_0820;
    92: op1_02_in22 = reg_1023;
    93: op1_02_in22 = reg_0958;
    95: op1_02_in22 = imem05_in[99:96];
    96: op1_02_in22 = reg_0652;
    97: op1_02_in22 = reg_0060;
    default: op1_02_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv22 = 1;
    6: op1_02_inv22 = 1;
    8: op1_02_inv22 = 1;
    9: op1_02_inv22 = 1;
    11: op1_02_inv22 = 1;
    12: op1_02_inv22 = 1;
    13: op1_02_inv22 = 1;
    16: op1_02_inv22 = 1;
    18: op1_02_inv22 = 1;
    19: op1_02_inv22 = 1;
    20: op1_02_inv22 = 1;
    22: op1_02_inv22 = 1;
    24: op1_02_inv22 = 1;
    29: op1_02_inv22 = 1;
    30: op1_02_inv22 = 1;
    32: op1_02_inv22 = 1;
    34: op1_02_inv22 = 1;
    36: op1_02_inv22 = 1;
    37: op1_02_inv22 = 1;
    40: op1_02_inv22 = 1;
    41: op1_02_inv22 = 1;
    43: op1_02_inv22 = 1;
    44: op1_02_inv22 = 1;
    45: op1_02_inv22 = 1;
    46: op1_02_inv22 = 1;
    50: op1_02_inv22 = 1;
    53: op1_02_inv22 = 1;
    56: op1_02_inv22 = 1;
    58: op1_02_inv22 = 1;
    59: op1_02_inv22 = 1;
    65: op1_02_inv22 = 1;
    68: op1_02_inv22 = 1;
    71: op1_02_inv22 = 1;
    72: op1_02_inv22 = 1;
    74: op1_02_inv22 = 1;
    76: op1_02_inv22 = 1;
    79: op1_02_inv22 = 1;
    80: op1_02_inv22 = 1;
    81: op1_02_inv22 = 1;
    82: op1_02_inv22 = 1;
    84: op1_02_inv22 = 1;
    89: op1_02_inv22 = 1;
    90: op1_02_inv22 = 1;
    95: op1_02_inv22 = 1;
    97: op1_02_inv22 = 1;
    default: op1_02_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in23 = imem04_in[7:4];
    6: op1_02_in23 = reg_0507;
    7: op1_02_in23 = reg_0966;
    8: op1_02_in23 = reg_0521;
    9: op1_02_in23 = reg_0576;
    10: op1_02_in23 = reg_0530;
    11: op1_02_in23 = imem05_in[7:4];
    12: op1_02_in23 = reg_0328;
    13: op1_02_in23 = reg_0293;
    14: op1_02_in23 = reg_0236;
    15: op1_02_in23 = reg_0360;
    16: op1_02_in23 = imem05_in[87:84];
    18: op1_02_in23 = reg_0599;
    19: op1_02_in23 = reg_0195;
    20: op1_02_in23 = reg_0592;
    21: op1_02_in23 = imem07_in[27:24];
    22: op1_02_in23 = imem03_in[127:124];
    23: op1_02_in23 = reg_0059;
    24: op1_02_in23 = reg_0099;
    25: op1_02_in23 = reg_0491;
    26: op1_02_in23 = reg_0715;
    27: op1_02_in23 = reg_0946;
    29: op1_02_in23 = reg_0590;
    30: op1_02_in23 = reg_0932;
    32: op1_02_in23 = reg_0082;
    33: op1_02_in23 = reg_0282;
    34: op1_02_in23 = reg_0256;
    76: op1_02_in23 = reg_0256;
    35: op1_02_in23 = reg_0327;
    36: op1_02_in23 = reg_0114;
    37: op1_02_in23 = reg_0397;
    38: op1_02_in23 = reg_0292;
    39: op1_02_in23 = reg_0483;
    40: op1_02_in23 = imem07_in[119:116];
    41: op1_02_in23 = reg_0128;
    42: op1_02_in23 = imem01_in[19:16];
    65: op1_02_in23 = imem01_in[19:16];
    43: op1_02_in23 = reg_0484;
    44: op1_02_in23 = reg_0736;
    45: op1_02_in23 = imem07_in[111:108];
    46: op1_02_in23 = reg_0118;
    47: op1_02_in23 = reg_0536;
    48: op1_02_in23 = reg_0819;
    49: op1_02_in23 = reg_0123;
    50: op1_02_in23 = reg_0476;
    52: op1_02_in23 = reg_0856;
    53: op1_02_in23 = reg_0711;
    54: op1_02_in23 = reg_0161;
    56: op1_02_in23 = reg_0918;
    57: op1_02_in23 = reg_0482;
    58: op1_02_in23 = imem03_in[35:32];
    59: op1_02_in23 = reg_1034;
    60: op1_02_in23 = reg_0332;
    61: op1_02_in23 = reg_0377;
    62: op1_02_in23 = reg_0066;
    63: op1_02_in23 = reg_0838;
    66: op1_02_in23 = reg_1040;
    67: op1_02_in23 = imem01_in[107:104];
    68: op1_02_in23 = reg_0798;
    69: op1_02_in23 = reg_0142;
    71: op1_02_in23 = reg_0894;
    72: op1_02_in23 = reg_0168;
    73: op1_02_in23 = imem01_in[59:56];
    74: op1_02_in23 = reg_1022;
    75: op1_02_in23 = reg_0086;
    77: op1_02_in23 = reg_0140;
    78: op1_02_in23 = imem07_in[99:96];
    79: op1_02_in23 = imem01_in[75:72];
    80: op1_02_in23 = reg_0793;
    81: op1_02_in23 = reg_0535;
    82: op1_02_in23 = reg_0876;
    83: op1_02_in23 = reg_0532;
    84: op1_02_in23 = reg_0957;
    85: op1_02_in23 = reg_1014;
    86: op1_02_in23 = reg_0345;
    89: op1_02_in23 = reg_0385;
    90: op1_02_in23 = reg_0962;
    91: op1_02_in23 = reg_0234;
    92: op1_02_in23 = reg_0500;
    93: op1_02_in23 = reg_0330;
    94: op1_02_in23 = reg_0648;
    95: op1_02_in23 = imem05_in[103:100];
    96: op1_02_in23 = reg_0647;
    97: op1_02_in23 = reg_0961;
    default: op1_02_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv23 = 1;
    6: op1_02_inv23 = 1;
    8: op1_02_inv23 = 1;
    10: op1_02_inv23 = 1;
    13: op1_02_inv23 = 1;
    15: op1_02_inv23 = 1;
    18: op1_02_inv23 = 1;
    22: op1_02_inv23 = 1;
    23: op1_02_inv23 = 1;
    25: op1_02_inv23 = 1;
    27: op1_02_inv23 = 1;
    32: op1_02_inv23 = 1;
    33: op1_02_inv23 = 1;
    35: op1_02_inv23 = 1;
    37: op1_02_inv23 = 1;
    38: op1_02_inv23 = 1;
    39: op1_02_inv23 = 1;
    41: op1_02_inv23 = 1;
    44: op1_02_inv23 = 1;
    45: op1_02_inv23 = 1;
    46: op1_02_inv23 = 1;
    54: op1_02_inv23 = 1;
    59: op1_02_inv23 = 1;
    60: op1_02_inv23 = 1;
    61: op1_02_inv23 = 1;
    66: op1_02_inv23 = 1;
    67: op1_02_inv23 = 1;
    68: op1_02_inv23 = 1;
    69: op1_02_inv23 = 1;
    72: op1_02_inv23 = 1;
    73: op1_02_inv23 = 1;
    75: op1_02_inv23 = 1;
    76: op1_02_inv23 = 1;
    77: op1_02_inv23 = 1;
    79: op1_02_inv23 = 1;
    84: op1_02_inv23 = 1;
    85: op1_02_inv23 = 1;
    89: op1_02_inv23 = 1;
    93: op1_02_inv23 = 1;
    95: op1_02_inv23 = 1;
    96: op1_02_inv23 = 1;
    97: op1_02_inv23 = 1;
    default: op1_02_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in24 = imem04_in[11:8];
    6: op1_02_in24 = reg_0508;
    7: op1_02_in24 = reg_0967;
    8: op1_02_in24 = reg_0510;
    9: op1_02_in24 = reg_0321;
    10: op1_02_in24 = reg_0534;
    11: op1_02_in24 = imem05_in[75:72];
    12: op1_02_in24 = reg_0089;
    13: op1_02_in24 = reg_0285;
    14: op1_02_in24 = reg_0248;
    15: op1_02_in24 = reg_0385;
    16: op1_02_in24 = imem05_in[107:104];
    18: op1_02_in24 = reg_0572;
    19: op1_02_in24 = reg_0199;
    20: op1_02_in24 = reg_0563;
    21: op1_02_in24 = imem07_in[43:40];
    22: op1_02_in24 = reg_0586;
    23: op1_02_in24 = reg_0748;
    24: op1_02_in24 = reg_0107;
    25: op1_02_in24 = reg_0254;
    26: op1_02_in24 = reg_0706;
    27: op1_02_in24 = reg_0834;
    29: op1_02_in24 = reg_0847;
    30: op1_02_in24 = reg_0760;
    32: op1_02_in24 = reg_0037;
    33: op1_02_in24 = reg_0912;
    34: op1_02_in24 = reg_0757;
    35: op1_02_in24 = reg_0398;
    36: op1_02_in24 = reg_0127;
    37: op1_02_in24 = reg_0396;
    38: op1_02_in24 = reg_0888;
    39: op1_02_in24 = reg_0536;
    40: op1_02_in24 = reg_0719;
    41: op1_02_in24 = reg_0142;
    42: op1_02_in24 = imem01_in[43:40];
    43: op1_02_in24 = reg_0872;
    44: op1_02_in24 = reg_0057;
    45: op1_02_in24 = reg_0720;
    46: op1_02_in24 = reg_0099;
    86: op1_02_in24 = reg_0099;
    47: op1_02_in24 = reg_0507;
    48: op1_02_in24 = reg_0136;
    49: op1_02_in24 = reg_0103;
    50: op1_02_in24 = reg_0470;
    52: op1_02_in24 = reg_0892;
    53: op1_02_in24 = reg_0700;
    54: op1_02_in24 = reg_0162;
    56: op1_02_in24 = reg_0936;
    57: op1_02_in24 = reg_0876;
    58: op1_02_in24 = imem03_in[39:36];
    59: op1_02_in24 = reg_1039;
    90: op1_02_in24 = reg_1039;
    60: op1_02_in24 = reg_0856;
    61: op1_02_in24 = reg_0822;
    62: op1_02_in24 = reg_0302;
    63: op1_02_in24 = reg_0180;
    65: op1_02_in24 = imem01_in[23:20];
    66: op1_02_in24 = reg_0902;
    67: op1_02_in24 = reg_0592;
    68: op1_02_in24 = reg_1017;
    69: op1_02_in24 = reg_0146;
    71: op1_02_in24 = reg_0358;
    73: op1_02_in24 = imem01_in[75:72];
    74: op1_02_in24 = reg_0962;
    75: op1_02_in24 = reg_0090;
    76: op1_02_in24 = reg_0963;
    77: op1_02_in24 = reg_0648;
    78: op1_02_in24 = reg_0919;
    79: op1_02_in24 = imem01_in[79:76];
    80: op1_02_in24 = reg_0501;
    81: op1_02_in24 = reg_0357;
    82: op1_02_in24 = reg_0086;
    83: op1_02_in24 = reg_0350;
    84: op1_02_in24 = reg_0736;
    85: op1_02_in24 = reg_0488;
    89: op1_02_in24 = reg_0551;
    91: op1_02_in24 = reg_0520;
    92: op1_02_in24 = reg_1041;
    93: op1_02_in24 = reg_0960;
    94: op1_02_in24 = reg_0646;
    95: op1_02_in24 = imem05_in[119:116];
    96: op1_02_in24 = reg_0013;
    97: op1_02_in24 = reg_0523;
    default: op1_02_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv24 = 1;
    8: op1_02_inv24 = 1;
    10: op1_02_inv24 = 1;
    11: op1_02_inv24 = 1;
    13: op1_02_inv24 = 1;
    15: op1_02_inv24 = 1;
    18: op1_02_inv24 = 1;
    19: op1_02_inv24 = 1;
    21: op1_02_inv24 = 1;
    22: op1_02_inv24 = 1;
    24: op1_02_inv24 = 1;
    26: op1_02_inv24 = 1;
    27: op1_02_inv24 = 1;
    33: op1_02_inv24 = 1;
    38: op1_02_inv24 = 1;
    41: op1_02_inv24 = 1;
    42: op1_02_inv24 = 1;
    44: op1_02_inv24 = 1;
    46: op1_02_inv24 = 1;
    50: op1_02_inv24 = 1;
    52: op1_02_inv24 = 1;
    53: op1_02_inv24 = 1;
    54: op1_02_inv24 = 1;
    59: op1_02_inv24 = 1;
    65: op1_02_inv24 = 1;
    66: op1_02_inv24 = 1;
    68: op1_02_inv24 = 1;
    71: op1_02_inv24 = 1;
    76: op1_02_inv24 = 1;
    77: op1_02_inv24 = 1;
    78: op1_02_inv24 = 1;
    79: op1_02_inv24 = 1;
    81: op1_02_inv24 = 1;
    85: op1_02_inv24 = 1;
    86: op1_02_inv24 = 1;
    89: op1_02_inv24 = 1;
    90: op1_02_inv24 = 1;
    92: op1_02_inv24 = 1;
    95: op1_02_inv24 = 1;
    default: op1_02_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in25 = imem04_in[23:20];
    6: op1_02_in25 = reg_0232;
    7: op1_02_in25 = reg_0968;
    8: op1_02_in25 = reg_0226;
    9: op1_02_in25 = reg_0373;
    10: op1_02_in25 = reg_0529;
    11: op1_02_in25 = imem05_in[79:76];
    12: op1_02_in25 = reg_0084;
    13: op1_02_in25 = reg_0286;
    14: op1_02_in25 = reg_0245;
    15: op1_02_in25 = reg_0323;
    16: op1_02_in25 = imem05_in[123:120];
    95: op1_02_in25 = imem05_in[123:120];
    18: op1_02_in25 = reg_0576;
    19: op1_02_in25 = imem01_in[67:64];
    20: op1_02_in25 = reg_0597;
    21: op1_02_in25 = imem07_in[47:44];
    22: op1_02_in25 = reg_0582;
    23: op1_02_in25 = reg_0054;
    24: op1_02_in25 = reg_0127;
    25: op1_02_in25 = reg_0832;
    34: op1_02_in25 = reg_0832;
    26: op1_02_in25 = reg_0727;
    27: op1_02_in25 = reg_0257;
    29: op1_02_in25 = reg_0311;
    30: op1_02_in25 = reg_0296;
    32: op1_02_in25 = reg_0762;
    33: op1_02_in25 = reg_0540;
    35: op1_02_in25 = reg_0004;
    36: op1_02_in25 = imem02_in[39:36];
    37: op1_02_in25 = reg_0377;
    38: op1_02_in25 = reg_0778;
    39: op1_02_in25 = reg_1020;
    40: op1_02_in25 = reg_0723;
    41: op1_02_in25 = reg_0153;
    42: op1_02_in25 = imem01_in[55:52];
    43: op1_02_in25 = imem03_in[23:20];
    44: op1_02_in25 = reg_0773;
    45: op1_02_in25 = reg_0721;
    46: op1_02_in25 = reg_0108;
    47: op1_02_in25 = reg_0909;
    48: op1_02_in25 = reg_0128;
    49: op1_02_in25 = reg_0104;
    50: op1_02_in25 = reg_0193;
    52: op1_02_in25 = reg_0782;
    53: op1_02_in25 = reg_0575;
    54: op1_02_in25 = reg_0160;
    56: op1_02_in25 = reg_1056;
    57: op1_02_in25 = reg_0506;
    58: op1_02_in25 = imem03_in[47:44];
    59: op1_02_in25 = reg_0501;
    60: op1_02_in25 = reg_0044;
    61: op1_02_in25 = reg_0991;
    89: op1_02_in25 = reg_0991;
    62: op1_02_in25 = reg_0068;
    63: op1_02_in25 = reg_0177;
    65: op1_02_in25 = imem01_in[39:36];
    66: op1_02_in25 = reg_0354;
    67: op1_02_in25 = reg_0253;
    68: op1_02_in25 = reg_0111;
    69: op1_02_in25 = imem06_in[31:28];
    71: op1_02_in25 = reg_0739;
    73: op1_02_in25 = imem01_in[79:76];
    74: op1_02_in25 = reg_0496;
    75: op1_02_in25 = reg_0261;
    76: op1_02_in25 = reg_0255;
    77: op1_02_in25 = reg_0966;
    78: op1_02_in25 = reg_0784;
    79: op1_02_in25 = imem01_in[87:84];
    80: op1_02_in25 = reg_0216;
    81: op1_02_in25 = reg_0445;
    82: op1_02_in25 = reg_0077;
    83: op1_02_in25 = reg_0589;
    84: op1_02_in25 = reg_0943;
    85: op1_02_in25 = reg_1024;
    86: op1_02_in25 = reg_0434;
    90: op1_02_in25 = reg_0830;
    91: op1_02_in25 = reg_0616;
    92: op1_02_in25 = reg_1033;
    93: op1_02_in25 = reg_0707;
    94: op1_02_in25 = reg_0259;
    96: op1_02_in25 = reg_0648;
    97: op1_02_in25 = reg_0986;
    default: op1_02_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv25 = 1;
    7: op1_02_inv25 = 1;
    8: op1_02_inv25 = 1;
    10: op1_02_inv25 = 1;
    11: op1_02_inv25 = 1;
    12: op1_02_inv25 = 1;
    14: op1_02_inv25 = 1;
    15: op1_02_inv25 = 1;
    16: op1_02_inv25 = 1;
    18: op1_02_inv25 = 1;
    20: op1_02_inv25 = 1;
    21: op1_02_inv25 = 1;
    23: op1_02_inv25 = 1;
    24: op1_02_inv25 = 1;
    25: op1_02_inv25 = 1;
    34: op1_02_inv25 = 1;
    36: op1_02_inv25 = 1;
    39: op1_02_inv25 = 1;
    40: op1_02_inv25 = 1;
    42: op1_02_inv25 = 1;
    44: op1_02_inv25 = 1;
    47: op1_02_inv25 = 1;
    50: op1_02_inv25 = 1;
    53: op1_02_inv25 = 1;
    56: op1_02_inv25 = 1;
    57: op1_02_inv25 = 1;
    58: op1_02_inv25 = 1;
    61: op1_02_inv25 = 1;
    63: op1_02_inv25 = 1;
    65: op1_02_inv25 = 1;
    66: op1_02_inv25 = 1;
    67: op1_02_inv25 = 1;
    69: op1_02_inv25 = 1;
    71: op1_02_inv25 = 1;
    74: op1_02_inv25 = 1;
    78: op1_02_inv25 = 1;
    80: op1_02_inv25 = 1;
    85: op1_02_inv25 = 1;
    86: op1_02_inv25 = 1;
    90: op1_02_inv25 = 1;
    91: op1_02_inv25 = 1;
    92: op1_02_inv25 = 1;
    93: op1_02_inv25 = 1;
    94: op1_02_inv25 = 1;
    96: op1_02_inv25 = 1;
    97: op1_02_inv25 = 1;
    default: op1_02_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in26 = imem04_in[71:68];
    6: op1_02_in26 = reg_0218;
    7: op1_02_in26 = reg_0946;
    8: op1_02_in26 = reg_0239;
    9: op1_02_in26 = reg_0377;
    10: op1_02_in26 = reg_0548;
    11: op1_02_in26 = reg_0962;
    12: op1_02_in26 = reg_0087;
    13: op1_02_in26 = reg_0307;
    14: op1_02_in26 = reg_0507;
    15: op1_02_in26 = reg_0393;
    16: op1_02_in26 = reg_0958;
    18: op1_02_in26 = reg_0322;
    19: op1_02_in26 = imem01_in[79:76];
    20: op1_02_in26 = reg_0319;
    21: op1_02_in26 = imem07_in[79:76];
    22: op1_02_in26 = reg_0573;
    23: op1_02_in26 = reg_0283;
    24: op1_02_in26 = reg_0121;
    25: op1_02_in26 = reg_0819;
    84: op1_02_in26 = reg_0819;
    26: op1_02_in26 = reg_0438;
    27: op1_02_in26 = reg_1046;
    29: op1_02_in26 = reg_0807;
    30: op1_02_in26 = reg_0009;
    32: op1_02_in26 = reg_0336;
    33: op1_02_in26 = reg_0050;
    34: op1_02_in26 = reg_0138;
    35: op1_02_in26 = reg_0389;
    36: op1_02_in26 = imem02_in[95:92];
    37: op1_02_in26 = reg_0836;
    38: op1_02_in26 = reg_0537;
    39: op1_02_in26 = reg_0888;
    40: op1_02_in26 = reg_0708;
    41: op1_02_in26 = reg_0137;
    42: op1_02_in26 = reg_0235;
    43: op1_02_in26 = imem03_in[47:44];
    44: op1_02_in26 = imem05_in[3:0];
    60: op1_02_in26 = imem05_in[3:0];
    45: op1_02_in26 = reg_0713;
    46: op1_02_in26 = reg_0109;
    47: op1_02_in26 = reg_0056;
    48: op1_02_in26 = reg_0152;
    49: op1_02_in26 = reg_0117;
    50: op1_02_in26 = reg_0202;
    52: op1_02_in26 = reg_0627;
    53: op1_02_in26 = reg_0303;
    54: op1_02_in26 = reg_0164;
    56: op1_02_in26 = reg_1045;
    57: op1_02_in26 = reg_0310;
    58: op1_02_in26 = imem03_in[51:48];
    59: op1_02_in26 = reg_0500;
    61: op1_02_in26 = reg_0979;
    62: op1_02_in26 = reg_0074;
    63: op1_02_in26 = reg_0178;
    65: op1_02_in26 = imem01_in[59:56];
    66: op1_02_in26 = reg_0304;
    67: op1_02_in26 = reg_0501;
    68: op1_02_in26 = reg_0116;
    69: op1_02_in26 = imem06_in[71:68];
    71: op1_02_in26 = reg_0664;
    73: op1_02_in26 = imem01_in[87:84];
    74: op1_02_in26 = reg_0798;
    75: op1_02_in26 = reg_0840;
    76: op1_02_in26 = reg_0447;
    77: op1_02_in26 = reg_0935;
    78: op1_02_in26 = reg_0371;
    79: op1_02_in26 = imem01_in[127:124];
    80: op1_02_in26 = reg_0354;
    91: op1_02_in26 = reg_0354;
    81: op1_02_in26 = reg_0577;
    82: op1_02_in26 = reg_0884;
    83: op1_02_in26 = reg_0174;
    85: op1_02_in26 = reg_0522;
    86: op1_02_in26 = reg_0046;
    89: op1_02_in26 = reg_0992;
    90: op1_02_in26 = reg_0740;
    92: op1_02_in26 = reg_0827;
    93: op1_02_in26 = reg_0780;
    94: op1_02_in26 = reg_0892;
    95: op1_02_in26 = imem05_in[127:124];
    96: op1_02_in26 = reg_0063;
    97: op1_02_in26 = reg_0445;
    default: op1_02_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_02_inv26 = 1;
    10: op1_02_inv26 = 1;
    12: op1_02_inv26 = 1;
    14: op1_02_inv26 = 1;
    15: op1_02_inv26 = 1;
    16: op1_02_inv26 = 1;
    20: op1_02_inv26 = 1;
    26: op1_02_inv26 = 1;
    29: op1_02_inv26 = 1;
    32: op1_02_inv26 = 1;
    33: op1_02_inv26 = 1;
    34: op1_02_inv26 = 1;
    35: op1_02_inv26 = 1;
    38: op1_02_inv26 = 1;
    41: op1_02_inv26 = 1;
    45: op1_02_inv26 = 1;
    46: op1_02_inv26 = 1;
    47: op1_02_inv26 = 1;
    48: op1_02_inv26 = 1;
    49: op1_02_inv26 = 1;
    50: op1_02_inv26 = 1;
    52: op1_02_inv26 = 1;
    53: op1_02_inv26 = 1;
    57: op1_02_inv26 = 1;
    58: op1_02_inv26 = 1;
    59: op1_02_inv26 = 1;
    65: op1_02_inv26 = 1;
    66: op1_02_inv26 = 1;
    67: op1_02_inv26 = 1;
    68: op1_02_inv26 = 1;
    71: op1_02_inv26 = 1;
    73: op1_02_inv26 = 1;
    74: op1_02_inv26 = 1;
    75: op1_02_inv26 = 1;
    76: op1_02_inv26 = 1;
    81: op1_02_inv26 = 1;
    82: op1_02_inv26 = 1;
    85: op1_02_inv26 = 1;
    86: op1_02_inv26 = 1;
    94: op1_02_inv26 = 1;
    95: op1_02_inv26 = 1;
    97: op1_02_inv26 = 1;
    default: op1_02_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in27 = reg_0543;
    6: op1_02_in27 = reg_0242;
    7: op1_02_in27 = reg_0961;
    8: op1_02_in27 = reg_0227;
    9: op1_02_in27 = reg_0987;
    10: op1_02_in27 = reg_0555;
    68: op1_02_in27 = reg_0555;
    11: op1_02_in27 = reg_0963;
    12: op1_02_in27 = imem03_in[7:4];
    13: op1_02_in27 = reg_0063;
    14: op1_02_in27 = reg_0905;
    15: op1_02_in27 = reg_0396;
    16: op1_02_in27 = reg_0971;
    18: op1_02_in27 = reg_0374;
    19: op1_02_in27 = imem01_in[111:108];
    20: op1_02_in27 = reg_0998;
    21: op1_02_in27 = imem07_in[91:88];
    22: op1_02_in27 = reg_0587;
    23: op1_02_in27 = reg_0043;
    24: op1_02_in27 = reg_0126;
    25: op1_02_in27 = reg_0135;
    26: op1_02_in27 = reg_0175;
    27: op1_02_in27 = reg_0497;
    29: op1_02_in27 = reg_0513;
    30: op1_02_in27 = reg_0732;
    32: op1_02_in27 = reg_0007;
    33: op1_02_in27 = reg_0541;
    34: op1_02_in27 = reg_0140;
    35: op1_02_in27 = reg_0874;
    36: op1_02_in27 = imem02_in[99:96];
    37: op1_02_in27 = reg_0376;
    38: op1_02_in27 = reg_0760;
    39: op1_02_in27 = reg_0778;
    40: op1_02_in27 = reg_0425;
    41: op1_02_in27 = reg_0134;
    42: op1_02_in27 = reg_0779;
    43: op1_02_in27 = imem03_in[91:88];
    44: op1_02_in27 = imem05_in[39:36];
    45: op1_02_in27 = reg_0701;
    46: op1_02_in27 = imem02_in[19:16];
    47: op1_02_in27 = reg_0815;
    48: op1_02_in27 = reg_0156;
    49: op1_02_in27 = imem02_in[51:48];
    50: op1_02_in27 = imem01_in[3:0];
    52: op1_02_in27 = reg_0754;
    53: op1_02_in27 = reg_0426;
    56: op1_02_in27 = reg_0238;
    57: op1_02_in27 = reg_0016;
    58: op1_02_in27 = imem03_in[103:100];
    59: op1_02_in27 = reg_0610;
    60: op1_02_in27 = imem05_in[19:16];
    61: op1_02_in27 = reg_0984;
    62: op1_02_in27 = reg_0072;
    63: op1_02_in27 = reg_0158;
    65: op1_02_in27 = imem01_in[67:64];
    66: op1_02_in27 = reg_0003;
    67: op1_02_in27 = reg_0830;
    69: op1_02_in27 = reg_0294;
    71: op1_02_in27 = reg_0052;
    73: op1_02_in27 = imem01_in[103:100];
    74: op1_02_in27 = reg_0514;
    75: op1_02_in27 = imem03_in[3:0];
    76: op1_02_in27 = reg_0960;
    77: op1_02_in27 = reg_0948;
    78: op1_02_in27 = reg_0805;
    79: op1_02_in27 = reg_0122;
    80: op1_02_in27 = reg_1055;
    81: op1_02_in27 = reg_0585;
    82: op1_02_in27 = imem03_in[55:52];
    83: op1_02_in27 = reg_0429;
    84: op1_02_in27 = reg_0780;
    85: op1_02_in27 = reg_0520;
    86: op1_02_in27 = reg_0547;
    89: op1_02_in27 = reg_0999;
    90: op1_02_in27 = reg_0304;
    91: op1_02_in27 = reg_1041;
    92: op1_02_in27 = imem02_in[31:28];
    93: op1_02_in27 = reg_0486;
    94: op1_02_in27 = reg_0964;
    95: op1_02_in27 = reg_0492;
    96: op1_02_in27 = reg_0958;
    97: op1_02_in27 = reg_0989;
    default: op1_02_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv27 = 1;
    6: op1_02_inv27 = 1;
    7: op1_02_inv27 = 1;
    8: op1_02_inv27 = 1;
    10: op1_02_inv27 = 1;
    12: op1_02_inv27 = 1;
    13: op1_02_inv27 = 1;
    21: op1_02_inv27 = 1;
    34: op1_02_inv27 = 1;
    36: op1_02_inv27 = 1;
    38: op1_02_inv27 = 1;
    41: op1_02_inv27 = 1;
    45: op1_02_inv27 = 1;
    47: op1_02_inv27 = 1;
    50: op1_02_inv27 = 1;
    53: op1_02_inv27 = 1;
    56: op1_02_inv27 = 1;
    60: op1_02_inv27 = 1;
    65: op1_02_inv27 = 1;
    66: op1_02_inv27 = 1;
    67: op1_02_inv27 = 1;
    68: op1_02_inv27 = 1;
    74: op1_02_inv27 = 1;
    77: op1_02_inv27 = 1;
    78: op1_02_inv27 = 1;
    79: op1_02_inv27 = 1;
    81: op1_02_inv27 = 1;
    82: op1_02_inv27 = 1;
    83: op1_02_inv27 = 1;
    84: op1_02_inv27 = 1;
    85: op1_02_inv27 = 1;
    86: op1_02_inv27 = 1;
    90: op1_02_inv27 = 1;
    91: op1_02_inv27 = 1;
    92: op1_02_inv27 = 1;
    94: op1_02_inv27 = 1;
    default: op1_02_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in28 = reg_0544;
    6: op1_02_in28 = reg_0240;
    7: op1_02_in28 = reg_0251;
    8: op1_02_in28 = reg_0105;
    9: op1_02_in28 = reg_0998;
    10: op1_02_in28 = reg_0531;
    11: op1_02_in28 = reg_0956;
    12: op1_02_in28 = imem03_in[87:84];
    13: op1_02_in28 = reg_0070;
    14: op1_02_in28 = reg_1033;
    15: op1_02_in28 = reg_0309;
    16: op1_02_in28 = reg_0942;
    18: op1_02_in28 = reg_0331;
    19: op1_02_in28 = reg_1051;
    74: op1_02_in28 = reg_1051;
    20: op1_02_in28 = reg_1002;
    21: op1_02_in28 = imem07_in[95:92];
    22: op1_02_in28 = reg_0594;
    23: op1_02_in28 = reg_0774;
    24: op1_02_in28 = imem02_in[55:52];
    25: op1_02_in28 = reg_0142;
    26: op1_02_in28 = reg_0179;
    27: op1_02_in28 = reg_0128;
    29: op1_02_in28 = reg_0374;
    30: op1_02_in28 = reg_0278;
    32: op1_02_in28 = reg_0758;
    33: op1_02_in28 = reg_0537;
    34: op1_02_in28 = imem06_in[27:24];
    35: op1_02_in28 = reg_0234;
    36: op1_02_in28 = imem02_in[103:100];
    37: op1_02_in28 = reg_0820;
    38: op1_02_in28 = reg_0075;
    39: op1_02_in28 = reg_0931;
    40: op1_02_in28 = reg_0423;
    41: op1_02_in28 = reg_0144;
    42: op1_02_in28 = reg_0560;
    43: op1_02_in28 = imem03_in[99:96];
    44: op1_02_in28 = imem05_in[63:60];
    45: op1_02_in28 = reg_0428;
    46: op1_02_in28 = imem02_in[23:20];
    47: op1_02_in28 = reg_0284;
    48: op1_02_in28 = reg_0130;
    49: op1_02_in28 = imem02_in[71:68];
    50: op1_02_in28 = imem01_in[19:16];
    52: op1_02_in28 = reg_0387;
    53: op1_02_in28 = reg_0175;
    56: op1_02_in28 = reg_0285;
    57: op1_02_in28 = reg_0884;
    58: op1_02_in28 = imem03_in[111:108];
    59: op1_02_in28 = reg_1017;
    91: op1_02_in28 = reg_1017;
    60: op1_02_in28 = imem05_in[43:40];
    61: op1_02_in28 = reg_0996;
    62: op1_02_in28 = reg_0041;
    63: op1_02_in28 = reg_0184;
    65: op1_02_in28 = imem01_in[71:68];
    66: op1_02_in28 = reg_0733;
    67: op1_02_in28 = reg_0616;
    68: op1_02_in28 = reg_0877;
    69: op1_02_in28 = reg_0393;
    71: op1_02_in28 = reg_0394;
    73: op1_02_in28 = reg_0122;
    75: op1_02_in28 = imem03_in[39:36];
    76: op1_02_in28 = reg_0528;
    77: op1_02_in28 = reg_0221;
    78: op1_02_in28 = reg_0589;
    79: op1_02_in28 = reg_0973;
    80: op1_02_in28 = reg_0769;
    81: op1_02_in28 = reg_0346;
    82: op1_02_in28 = imem03_in[91:88];
    83: op1_02_in28 = reg_0161;
    84: op1_02_in28 = reg_0135;
    85: op1_02_in28 = reg_1041;
    86: op1_02_in28 = reg_0609;
    89: op1_02_in28 = reg_0990;
    90: op1_02_in28 = reg_0115;
    92: op1_02_in28 = imem02_in[79:76];
    93: op1_02_in28 = reg_0806;
    94: op1_02_in28 = reg_0587;
    95: op1_02_in28 = reg_0139;
    96: op1_02_in28 = reg_0675;
    97: op1_02_in28 = reg_0286;
    default: op1_02_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv28 = 1;
    8: op1_02_inv28 = 1;
    9: op1_02_inv28 = 1;
    10: op1_02_inv28 = 1;
    12: op1_02_inv28 = 1;
    20: op1_02_inv28 = 1;
    27: op1_02_inv28 = 1;
    30: op1_02_inv28 = 1;
    32: op1_02_inv28 = 1;
    33: op1_02_inv28 = 1;
    38: op1_02_inv28 = 1;
    39: op1_02_inv28 = 1;
    40: op1_02_inv28 = 1;
    41: op1_02_inv28 = 1;
    42: op1_02_inv28 = 1;
    48: op1_02_inv28 = 1;
    50: op1_02_inv28 = 1;
    53: op1_02_inv28 = 1;
    57: op1_02_inv28 = 1;
    58: op1_02_inv28 = 1;
    59: op1_02_inv28 = 1;
    60: op1_02_inv28 = 1;
    62: op1_02_inv28 = 1;
    63: op1_02_inv28 = 1;
    66: op1_02_inv28 = 1;
    75: op1_02_inv28 = 1;
    76: op1_02_inv28 = 1;
    82: op1_02_inv28 = 1;
    85: op1_02_inv28 = 1;
    92: op1_02_inv28 = 1;
    97: op1_02_inv28 = 1;
    default: op1_02_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in29 = reg_0545;
    6: op1_02_in29 = reg_0227;
    7: op1_02_in29 = reg_0223;
    8: op1_02_in29 = reg_0124;
    9: op1_02_in29 = imem04_in[7:4];
    10: op1_02_in29 = reg_0556;
    11: op1_02_in29 = reg_0964;
    12: op1_02_in29 = imem03_in[91:88];
    13: op1_02_in29 = imem05_in[15:12];
    14: op1_02_in29 = reg_1036;
    15: op1_02_in29 = reg_0374;
    16: op1_02_in29 = reg_0968;
    18: op1_02_in29 = reg_0991;
    19: op1_02_in29 = reg_0503;
    79: op1_02_in29 = reg_0503;
    20: op1_02_in29 = reg_0992;
    21: op1_02_in29 = imem07_in[107:104];
    22: op1_02_in29 = reg_0387;
    23: op1_02_in29 = reg_0057;
    24: op1_02_in29 = imem02_in[103:100];
    25: op1_02_in29 = reg_0144;
    26: op1_02_in29 = reg_0161;
    27: op1_02_in29 = imem06_in[7:4];
    76: op1_02_in29 = imem06_in[7:4];
    29: op1_02_in29 = reg_0984;
    30: op1_02_in29 = reg_0748;
    32: op1_02_in29 = reg_0876;
    33: op1_02_in29 = reg_0313;
    34: op1_02_in29 = imem06_in[99:96];
    35: op1_02_in29 = reg_0989;
    36: op1_02_in29 = reg_0637;
    37: op1_02_in29 = reg_0844;
    38: op1_02_in29 = reg_0072;
    39: op1_02_in29 = reg_0050;
    40: op1_02_in29 = reg_0445;
    41: op1_02_in29 = imem06_in[3:0];
    42: op1_02_in29 = reg_0242;
    43: op1_02_in29 = imem03_in[107:104];
    44: op1_02_in29 = imem05_in[87:84];
    45: op1_02_in29 = reg_0024;
    46: op1_02_in29 = imem02_in[67:64];
    47: op1_02_in29 = reg_0308;
    48: op1_02_in29 = imem06_in[59:56];
    49: op1_02_in29 = imem02_in[87:84];
    50: op1_02_in29 = imem01_in[51:48];
    52: op1_02_in29 = reg_0294;
    53: op1_02_in29 = reg_0180;
    56: op1_02_in29 = reg_1043;
    57: op1_02_in29 = imem03_in[3:0];
    58: op1_02_in29 = reg_0099;
    59: op1_02_in29 = reg_1055;
    60: op1_02_in29 = imem05_in[63:60];
    61: op1_02_in29 = reg_0978;
    62: op1_02_in29 = reg_0494;
    65: op1_02_in29 = imem01_in[111:108];
    66: op1_02_in29 = reg_0555;
    67: op1_02_in29 = reg_0925;
    68: op1_02_in29 = imem02_in[23:20];
    69: op1_02_in29 = reg_0534;
    71: op1_02_in29 = reg_0054;
    73: op1_02_in29 = reg_1042;
    74: op1_02_in29 = reg_0112;
    75: op1_02_in29 = imem03_in[47:44];
    77: op1_02_in29 = reg_0865;
    78: op1_02_in29 = reg_0175;
    80: op1_02_in29 = reg_0860;
    81: op1_02_in29 = reg_0661;
    82: op1_02_in29 = imem03_in[103:100];
    83: op1_02_in29 = reg_0182;
    84: op1_02_in29 = reg_0508;
    85: op1_02_in29 = reg_0610;
    86: op1_02_in29 = reg_0995;
    89: op1_02_in29 = reg_1000;
    90: op1_02_in29 = reg_0109;
    91: op1_02_in29 = reg_0906;
    92: op1_02_in29 = imem02_in[115:112];
    93: op1_02_in29 = reg_0951;
    94: op1_02_in29 = reg_0617;
    95: op1_02_in29 = reg_0141;
    96: op1_02_in29 = reg_0129;
    97: op1_02_in29 = reg_0975;
    default: op1_02_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv29 = 1;
    7: op1_02_inv29 = 1;
    8: op1_02_inv29 = 1;
    10: op1_02_inv29 = 1;
    12: op1_02_inv29 = 1;
    13: op1_02_inv29 = 1;
    15: op1_02_inv29 = 1;
    16: op1_02_inv29 = 1;
    18: op1_02_inv29 = 1;
    19: op1_02_inv29 = 1;
    20: op1_02_inv29 = 1;
    23: op1_02_inv29 = 1;
    26: op1_02_inv29 = 1;
    27: op1_02_inv29 = 1;
    29: op1_02_inv29 = 1;
    32: op1_02_inv29 = 1;
    33: op1_02_inv29 = 1;
    35: op1_02_inv29 = 1;
    37: op1_02_inv29 = 1;
    39: op1_02_inv29 = 1;
    41: op1_02_inv29 = 1;
    44: op1_02_inv29 = 1;
    50: op1_02_inv29 = 1;
    53: op1_02_inv29 = 1;
    56: op1_02_inv29 = 1;
    58: op1_02_inv29 = 1;
    59: op1_02_inv29 = 1;
    62: op1_02_inv29 = 1;
    65: op1_02_inv29 = 1;
    73: op1_02_inv29 = 1;
    74: op1_02_inv29 = 1;
    75: op1_02_inv29 = 1;
    76: op1_02_inv29 = 1;
    78: op1_02_inv29 = 1;
    85: op1_02_inv29 = 1;
    90: op1_02_inv29 = 1;
    93: op1_02_inv29 = 1;
    94: op1_02_inv29 = 1;
    95: op1_02_inv29 = 1;
    default: op1_02_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_02_in30 = reg_0546;
    6: op1_02_in30 = reg_0219;
    7: op1_02_in30 = reg_0147;
    8: op1_02_in30 = reg_0111;
    9: op1_02_in30 = imem04_in[67:64];
    10: op1_02_in30 = reg_0547;
    97: op1_02_in30 = reg_0547;
    11: op1_02_in30 = reg_0951;
    12: op1_02_in30 = imem03_in[107:104];
    13: op1_02_in30 = imem05_in[39:36];
    14: op1_02_in30 = reg_0871;
    15: op1_02_in30 = reg_0991;
    16: op1_02_in30 = reg_0900;
    18: op1_02_in30 = reg_0993;
    29: op1_02_in30 = reg_0993;
    19: op1_02_in30 = reg_1052;
    20: op1_02_in30 = reg_0995;
    21: op1_02_in30 = reg_0720;
    22: op1_02_in30 = reg_0317;
    23: op1_02_in30 = reg_0044;
    24: op1_02_in30 = reg_0654;
    25: op1_02_in30 = reg_0962;
    26: op1_02_in30 = reg_0169;
    53: op1_02_in30 = reg_0169;
    27: op1_02_in30 = imem06_in[59:56];
    30: op1_02_in30 = reg_0043;
    32: op1_02_in30 = reg_0090;
    33: op1_02_in30 = reg_0764;
    34: op1_02_in30 = reg_0617;
    35: op1_02_in30 = reg_0994;
    89: op1_02_in30 = reg_0994;
    36: op1_02_in30 = reg_0657;
    37: op1_02_in30 = reg_0822;
    38: op1_02_in30 = reg_0278;
    39: op1_02_in30 = reg_0740;
    40: op1_02_in30 = reg_0427;
    41: op1_02_in30 = imem06_in[39:36];
    42: op1_02_in30 = reg_0555;
    43: op1_02_in30 = reg_0357;
    58: op1_02_in30 = reg_0357;
    44: op1_02_in30 = imem05_in[127:124];
    45: op1_02_in30 = reg_0167;
    46: op1_02_in30 = imem02_in[75:72];
    47: op1_02_in30 = reg_0763;
    48: op1_02_in30 = imem06_in[67:64];
    49: op1_02_in30 = imem02_in[107:104];
    50: op1_02_in30 = imem01_in[55:52];
    52: op1_02_in30 = reg_0391;
    56: op1_02_in30 = reg_0829;
    57: op1_02_in30 = imem03_in[63:60];
    59: op1_02_in30 = reg_0116;
    60: op1_02_in30 = imem05_in[71:68];
    61: op1_02_in30 = reg_0990;
    62: op1_02_in30 = imem05_in[23:20];
    65: op1_02_in30 = reg_0223;
    66: op1_02_in30 = reg_0827;
    67: op1_02_in30 = reg_1055;
    68: op1_02_in30 = imem02_in[51:48];
    69: op1_02_in30 = reg_1030;
    71: op1_02_in30 = reg_0083;
    73: op1_02_in30 = reg_1023;
    74: op1_02_in30 = reg_0860;
    75: op1_02_in30 = imem03_in[59:56];
    76: op1_02_in30 = imem06_in[11:8];
    77: op1_02_in30 = reg_0004;
    78: op1_02_in30 = reg_0172;
    79: op1_02_in30 = reg_0518;
    80: op1_02_in30 = reg_0745;
    81: op1_02_in30 = reg_0576;
    82: op1_02_in30 = imem03_in[115:112];
    83: op1_02_in30 = reg_0183;
    84: op1_02_in30 = reg_0706;
    85: op1_02_in30 = reg_0232;
    86: op1_02_in30 = reg_0978;
    90: op1_02_in30 = imem02_in[15:12];
    91: op1_02_in30 = reg_0769;
    92: op1_02_in30 = reg_0554;
    93: op1_02_in30 = reg_0326;
    94: op1_02_in30 = reg_0019;
    95: op1_02_in30 = reg_0226;
    96: op1_02_in30 = reg_0257;
    default: op1_02_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv30 = 1;
    6: op1_02_inv30 = 1;
    8: op1_02_inv30 = 1;
    9: op1_02_inv30 = 1;
    10: op1_02_inv30 = 1;
    11: op1_02_inv30 = 1;
    15: op1_02_inv30 = 1;
    18: op1_02_inv30 = 1;
    19: op1_02_inv30 = 1;
    23: op1_02_inv30 = 1;
    24: op1_02_inv30 = 1;
    27: op1_02_inv30 = 1;
    34: op1_02_inv30 = 1;
    35: op1_02_inv30 = 1;
    37: op1_02_inv30 = 1;
    41: op1_02_inv30 = 1;
    42: op1_02_inv30 = 1;
    48: op1_02_inv30 = 1;
    50: op1_02_inv30 = 1;
    53: op1_02_inv30 = 1;
    60: op1_02_inv30 = 1;
    67: op1_02_inv30 = 1;
    69: op1_02_inv30 = 1;
    71: op1_02_inv30 = 1;
    73: op1_02_inv30 = 1;
    74: op1_02_inv30 = 1;
    75: op1_02_inv30 = 1;
    77: op1_02_inv30 = 1;
    78: op1_02_inv30 = 1;
    79: op1_02_inv30 = 1;
    82: op1_02_inv30 = 1;
    84: op1_02_inv30 = 1;
    90: op1_02_inv30 = 1;
    93: op1_02_inv30 = 1;
    97: op1_02_inv30 = 1;
    default: op1_02_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_02_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_02_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in00 = reg_0547;
    6: op1_03_in00 = reg_0122;
    7: op1_03_in00 = reg_0149;
    8: op1_03_in00 = reg_0125;
    9: op1_03_in00 = imem04_in[91:88];
    10: op1_03_in00 = reg_0281;
    4: op1_03_in00 = imem07_in[27:24];
    3: op1_03_in00 = imem07_in[47:44];
    11: op1_03_in00 = reg_0942;
    44: op1_03_in00 = reg_0942;
    12: op1_03_in00 = imem03_in[127:124];
    13: op1_03_in00 = imem05_in[47:44];
    14: op1_03_in00 = reg_0904;
    15: op1_03_in00 = reg_0979;
    20: op1_03_in00 = reg_0979;
    16: op1_03_in00 = reg_0229;
    17: op1_03_in00 = imem00_in[27:24];
    18: op1_03_in00 = reg_0749;
    19: op1_03_in00 = reg_1039;
    2: op1_03_in00 = imem07_in[91:88];
    21: op1_03_in00 = imem00_in[59:56];
    22: op1_03_in00 = reg_0319;
    23: op1_03_in00 = imem05_in[31:28];
    24: op1_03_in00 = reg_0647;
    25: op1_03_in00 = imem06_in[39:36];
    26: op1_03_in00 = imem00_in[3:0];
    27: op1_03_in00 = imem06_in[71:68];
    28: op1_03_in00 = imem00_in[11:8];
    31: op1_03_in00 = imem00_in[11:8];
    63: op1_03_in00 = imem00_in[11:8];
    29: op1_03_in00 = reg_0990;
    30: op1_03_in00 = reg_0875;
    32: op1_03_in00 = reg_0077;
    33: op1_03_in00 = reg_0733;
    34: op1_03_in00 = reg_0619;
    35: op1_03_in00 = imem04_in[11:8];
    36: op1_03_in00 = reg_0665;
    37: op1_03_in00 = reg_0984;
    38: op1_03_in00 = reg_0059;
    39: op1_03_in00 = reg_0071;
    40: op1_03_in00 = reg_0437;
    41: op1_03_in00 = imem06_in[51:48];
    42: op1_03_in00 = reg_0087;
    43: op1_03_in00 = reg_0933;
    45: op1_03_in00 = imem00_in[55:52];
    46: op1_03_in00 = imem02_in[79:76];
    47: op1_03_in00 = imem05_in[11:8];
    48: op1_03_in00 = imem06_in[87:84];
    49: op1_03_in00 = imem02_in[123:120];
    50: op1_03_in00 = imem01_in[63:60];
    51: op1_03_in00 = imem00_in[83:80];
    52: op1_03_in00 = reg_0399;
    53: op1_03_in00 = reg_0160;
    54: op1_03_in00 = imem00_in[15:12];
    70: op1_03_in00 = imem00_in[15:12];
    55: op1_03_in00 = imem00_in[123:120];
    64: op1_03_in00 = imem00_in[123:120];
    56: op1_03_in00 = reg_1031;
    57: op1_03_in00 = imem03_in[79:76];
    58: op1_03_in00 = reg_0580;
    59: op1_03_in00 = reg_1053;
    60: op1_03_in00 = imem05_in[79:76];
    61: op1_03_in00 = reg_0994;
    62: op1_03_in00 = imem05_in[27:24];
    65: op1_03_in00 = reg_0870;
    66: op1_03_in00 = reg_0109;
    67: op1_03_in00 = reg_0769;
    68: op1_03_in00 = imem02_in[103:100];
    69: op1_03_in00 = reg_0008;
    71: op1_03_in00 = reg_0758;
    72: op1_03_in00 = imem00_in[7:4];
    73: op1_03_in00 = reg_0503;
    74: op1_03_in00 = imem02_in[23:20];
    75: op1_03_in00 = imem03_in[83:80];
    76: op1_03_in00 = imem06_in[43:40];
    77: op1_03_in00 = reg_0333;
    78: op1_03_in00 = reg_0169;
    79: op1_03_in00 = reg_0501;
    80: op1_03_in00 = imem02_in[3:0];
    81: op1_03_in00 = reg_0579;
    82: op1_03_in00 = reg_0620;
    83: op1_03_in00 = reg_0701;
    84: op1_03_in00 = reg_0816;
    85: op1_03_in00 = reg_0114;
    86: op1_03_in00 = imem04_in[15:12];
    87: op1_03_in00 = imem00_in[35:32];
    88: op1_03_in00 = imem00_in[99:96];
    89: op1_03_in00 = imem04_in[39:36];
    90: op1_03_in00 = imem02_in[19:16];
    91: op1_03_in00 = reg_0512;
    92: op1_03_in00 = reg_0348;
    93: op1_03_in00 = reg_0851;
    94: op1_03_in00 = reg_0709;
    95: op1_03_in00 = reg_0256;
    96: op1_03_in00 = reg_0780;
    97: op1_03_in00 = reg_0396;
    default: op1_03_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv00 = 1;
    4: op1_03_inv00 = 1;
    15: op1_03_inv00 = 1;
    16: op1_03_inv00 = 1;
    17: op1_03_inv00 = 1;
    18: op1_03_inv00 = 1;
    19: op1_03_inv00 = 1;
    2: op1_03_inv00 = 1;
    22: op1_03_inv00 = 1;
    31: op1_03_inv00 = 1;
    32: op1_03_inv00 = 1;
    35: op1_03_inv00 = 1;
    41: op1_03_inv00 = 1;
    42: op1_03_inv00 = 1;
    44: op1_03_inv00 = 1;
    47: op1_03_inv00 = 1;
    48: op1_03_inv00 = 1;
    51: op1_03_inv00 = 1;
    57: op1_03_inv00 = 1;
    58: op1_03_inv00 = 1;
    60: op1_03_inv00 = 1;
    61: op1_03_inv00 = 1;
    62: op1_03_inv00 = 1;
    63: op1_03_inv00 = 1;
    64: op1_03_inv00 = 1;
    65: op1_03_inv00 = 1;
    68: op1_03_inv00 = 1;
    69: op1_03_inv00 = 1;
    70: op1_03_inv00 = 1;
    71: op1_03_inv00 = 1;
    73: op1_03_inv00 = 1;
    77: op1_03_inv00 = 1;
    79: op1_03_inv00 = 1;
    80: op1_03_inv00 = 1;
    82: op1_03_inv00 = 1;
    86: op1_03_inv00 = 1;
    88: op1_03_inv00 = 1;
    89: op1_03_inv00 = 1;
    92: op1_03_inv00 = 1;
    93: op1_03_inv00 = 1;
    94: op1_03_inv00 = 1;
    96: op1_03_inv00 = 1;
    default: op1_03_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in01 = reg_0301;
    6: op1_03_in01 = reg_0114;
    7: op1_03_in01 = reg_0134;
    8: op1_03_in01 = reg_0116;
    9: op1_03_in01 = imem04_in[107:104];
    10: op1_03_in01 = reg_0283;
    59: op1_03_in01 = reg_0283;
    4: op1_03_in01 = imem07_in[51:48];
    3: op1_03_in01 = imem07_in[63:60];
    11: op1_03_in01 = reg_0271;
    97: op1_03_in01 = reg_0271;
    12: op1_03_in01 = reg_0596;
    13: op1_03_in01 = imem05_in[71:68];
    14: op1_03_in01 = reg_0127;
    15: op1_03_in01 = reg_0981;
    16: op1_03_in01 = reg_0133;
    17: op1_03_in01 = imem00_in[115:112];
    63: op1_03_in01 = imem00_in[115:112];
    18: op1_03_in01 = reg_0776;
    19: op1_03_in01 = reg_0913;
    20: op1_03_in01 = reg_0993;
    21: op1_03_in01 = imem00_in[119:116];
    22: op1_03_in01 = reg_0377;
    23: op1_03_in01 = imem05_in[35:32];
    62: op1_03_in01 = imem05_in[35:32];
    24: op1_03_in01 = reg_0334;
    25: op1_03_in01 = reg_0625;
    26: op1_03_in01 = imem00_in[19:16];
    70: op1_03_in01 = imem00_in[19:16];
    72: op1_03_in01 = imem00_in[19:16];
    27: op1_03_in01 = imem06_in[75:72];
    41: op1_03_in01 = imem06_in[75:72];
    28: op1_03_in01 = imem00_in[43:40];
    29: op1_03_in01 = reg_0997;
    30: op1_03_in01 = reg_0286;
    31: op1_03_in01 = imem00_in[35:32];
    32: op1_03_in01 = imem03_in[19:16];
    33: op1_03_in01 = reg_0062;
    34: op1_03_in01 = reg_0618;
    35: op1_03_in01 = imem04_in[15:12];
    36: op1_03_in01 = reg_0291;
    37: op1_03_in01 = imem04_in[55:52];
    38: op1_03_in01 = reg_0056;
    39: op1_03_in01 = reg_0069;
    40: op1_03_in01 = reg_0435;
    42: op1_03_in01 = reg_0769;
    43: op1_03_in01 = reg_0397;
    44: op1_03_in01 = reg_0949;
    45: op1_03_in01 = imem00_in[59:56];
    46: op1_03_in01 = imem02_in[107:104];
    68: op1_03_in01 = imem02_in[107:104];
    47: op1_03_in01 = imem05_in[27:24];
    48: op1_03_in01 = imem06_in[115:112];
    49: op1_03_in01 = reg_0341;
    50: op1_03_in01 = imem01_in[75:72];
    51: op1_03_in01 = imem00_in[91:88];
    52: op1_03_in01 = reg_0222;
    53: op1_03_in01 = reg_0166;
    78: op1_03_in01 = reg_0166;
    54: op1_03_in01 = imem00_in[63:60];
    55: op1_03_in01 = reg_0472;
    56: op1_03_in01 = reg_0304;
    57: op1_03_in01 = reg_0445;
    58: op1_03_in01 = reg_0434;
    60: op1_03_in01 = imem05_in[107:104];
    61: op1_03_in01 = imem04_in[19:16];
    64: op1_03_in01 = reg_0523;
    65: op1_03_in01 = reg_1056;
    66: op1_03_in01 = reg_0877;
    67: op1_03_in01 = reg_0111;
    69: op1_03_in01 = reg_1010;
    71: op1_03_in01 = reg_0867;
    73: op1_03_in01 = reg_0487;
    74: op1_03_in01 = imem02_in[47:44];
    75: op1_03_in01 = reg_0357;
    76: op1_03_in01 = imem06_in[83:80];
    77: op1_03_in01 = reg_0709;
    79: op1_03_in01 = reg_1040;
    80: op1_03_in01 = imem02_in[119:116];
    81: op1_03_in01 = reg_0230;
    82: op1_03_in01 = reg_0760;
    83: op1_03_in01 = reg_0157;
    84: op1_03_in01 = reg_0258;
    85: op1_03_in01 = reg_0860;
    86: op1_03_in01 = imem04_in[51:48];
    87: op1_03_in01 = imem00_in[39:36];
    88: op1_03_in01 = reg_0685;
    89: op1_03_in01 = imem04_in[59:56];
    90: op1_03_in01 = imem02_in[91:88];
    91: op1_03_in01 = reg_0003;
    92: op1_03_in01 = reg_0855;
    93: op1_03_in01 = reg_0657;
    94: op1_03_in01 = reg_0795;
    95: op1_03_in01 = reg_0152;
    96: op1_03_in01 = reg_0145;
    default: op1_03_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv01 = 1;
    6: op1_03_inv01 = 1;
    8: op1_03_inv01 = 1;
    10: op1_03_inv01 = 1;
    11: op1_03_inv01 = 1;
    12: op1_03_inv01 = 1;
    13: op1_03_inv01 = 1;
    14: op1_03_inv01 = 1;
    17: op1_03_inv01 = 1;
    19: op1_03_inv01 = 1;
    20: op1_03_inv01 = 1;
    21: op1_03_inv01 = 1;
    23: op1_03_inv01 = 1;
    24: op1_03_inv01 = 1;
    25: op1_03_inv01 = 1;
    26: op1_03_inv01 = 1;
    27: op1_03_inv01 = 1;
    28: op1_03_inv01 = 1;
    32: op1_03_inv01 = 1;
    34: op1_03_inv01 = 1;
    35: op1_03_inv01 = 1;
    39: op1_03_inv01 = 1;
    41: op1_03_inv01 = 1;
    44: op1_03_inv01 = 1;
    46: op1_03_inv01 = 1;
    51: op1_03_inv01 = 1;
    53: op1_03_inv01 = 1;
    55: op1_03_inv01 = 1;
    57: op1_03_inv01 = 1;
    58: op1_03_inv01 = 1;
    59: op1_03_inv01 = 1;
    60: op1_03_inv01 = 1;
    61: op1_03_inv01 = 1;
    65: op1_03_inv01 = 1;
    66: op1_03_inv01 = 1;
    67: op1_03_inv01 = 1;
    69: op1_03_inv01 = 1;
    72: op1_03_inv01 = 1;
    73: op1_03_inv01 = 1;
    74: op1_03_inv01 = 1;
    76: op1_03_inv01 = 1;
    81: op1_03_inv01 = 1;
    84: op1_03_inv01 = 1;
    85: op1_03_inv01 = 1;
    91: op1_03_inv01 = 1;
    93: op1_03_inv01 = 1;
    96: op1_03_inv01 = 1;
    default: op1_03_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in02 = reg_0302;
    6: op1_03_in02 = reg_0113;
    7: op1_03_in02 = imem06_in[27:24];
    8: op1_03_in02 = reg_0117;
    9: op1_03_in02 = imem04_in[111:108];
    10: op1_03_in02 = reg_0282;
    4: op1_03_in02 = imem07_in[79:76];
    3: op1_03_in02 = imem07_in[79:76];
    11: op1_03_in02 = reg_0273;
    59: op1_03_in02 = reg_0273;
    12: op1_03_in02 = reg_0578;
    13: op1_03_in02 = reg_0952;
    14: op1_03_in02 = reg_0110;
    66: op1_03_in02 = reg_0110;
    15: op1_03_in02 = reg_1000;
    16: op1_03_in02 = reg_0151;
    17: op1_03_in02 = reg_0693;
    18: op1_03_in02 = reg_0041;
    19: op1_03_in02 = reg_0871;
    20: op1_03_in02 = reg_0981;
    21: op1_03_in02 = reg_0672;
    22: op1_03_in02 = reg_0397;
    23: op1_03_in02 = imem05_in[51:48];
    24: op1_03_in02 = reg_0333;
    25: op1_03_in02 = reg_0613;
    26: op1_03_in02 = imem00_in[35:32];
    27: op1_03_in02 = imem06_in[95:92];
    41: op1_03_in02 = imem06_in[95:92];
    28: op1_03_in02 = imem00_in[127:124];
    29: op1_03_in02 = imem04_in[55:52];
    30: op1_03_in02 = imem05_in[67:64];
    31: op1_03_in02 = imem00_in[71:68];
    32: op1_03_in02 = imem03_in[43:40];
    36: op1_03_in02 = imem03_in[43:40];
    33: op1_03_in02 = reg_0066;
    34: op1_03_in02 = reg_0632;
    35: op1_03_in02 = imem04_in[19:16];
    37: op1_03_in02 = imem04_in[87:84];
    38: op1_03_in02 = reg_0053;
    39: op1_03_in02 = reg_0738;
    40: op1_03_in02 = reg_0179;
    42: op1_03_in02 = reg_0501;
    43: op1_03_in02 = reg_0874;
    44: op1_03_in02 = reg_0946;
    45: op1_03_in02 = imem00_in[63:60];
    46: op1_03_in02 = reg_0341;
    47: op1_03_in02 = imem05_in[71:68];
    48: op1_03_in02 = reg_0759;
    49: op1_03_in02 = reg_0026;
    50: op1_03_in02 = imem01_in[83:80];
    51: op1_03_in02 = imem00_in[95:92];
    70: op1_03_in02 = imem00_in[95:92];
    52: op1_03_in02 = reg_0628;
    53: op1_03_in02 = reg_0177;
    54: op1_03_in02 = imem00_in[67:64];
    55: op1_03_in02 = imem01_in[19:16];
    56: op1_03_in02 = reg_0283;
    57: op1_03_in02 = reg_0585;
    58: op1_03_in02 = reg_0662;
    60: op1_03_in02 = reg_0944;
    61: op1_03_in02 = imem04_in[35:32];
    62: op1_03_in02 = imem05_in[75:72];
    63: op1_03_in02 = reg_0519;
    64: op1_03_in02 = reg_0463;
    65: op1_03_in02 = reg_0607;
    67: op1_03_in02 = reg_0112;
    68: op1_03_in02 = reg_0914;
    69: op1_03_in02 = imem07_in[63:60];
    71: op1_03_in02 = reg_0792;
    72: op1_03_in02 = imem00_in[75:72];
    73: op1_03_in02 = reg_1024;
    74: op1_03_in02 = imem02_in[51:48];
    75: op1_03_in02 = reg_0445;
    76: op1_03_in02 = imem06_in[99:96];
    77: op1_03_in02 = reg_0806;
    96: op1_03_in02 = reg_0806;
    78: op1_03_in02 = reg_0173;
    79: op1_03_in02 = reg_1041;
    80: op1_03_in02 = reg_0096;
    81: op1_03_in02 = reg_0779;
    82: op1_03_in02 = reg_0580;
    83: op1_03_in02 = reg_0697;
    84: op1_03_in02 = reg_0326;
    94: op1_03_in02 = reg_0326;
    85: op1_03_in02 = reg_0877;
    86: op1_03_in02 = imem04_in[99:96];
    87: op1_03_in02 = imem00_in[47:44];
    88: op1_03_in02 = reg_0686;
    89: op1_03_in02 = imem04_in[127:124];
    90: op1_03_in02 = imem02_in[127:124];
    91: op1_03_in02 = reg_0745;
    92: op1_03_in02 = reg_0095;
    93: op1_03_in02 = imem06_in[59:56];
    95: op1_03_in02 = reg_0129;
    97: op1_03_in02 = imem04_in[23:20];
    default: op1_03_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_03_inv02 = 1;
    9: op1_03_inv02 = 1;
    10: op1_03_inv02 = 1;
    4: op1_03_inv02 = 1;
    12: op1_03_inv02 = 1;
    14: op1_03_inv02 = 1;
    19: op1_03_inv02 = 1;
    20: op1_03_inv02 = 1;
    22: op1_03_inv02 = 1;
    24: op1_03_inv02 = 1;
    25: op1_03_inv02 = 1;
    30: op1_03_inv02 = 1;
    31: op1_03_inv02 = 1;
    34: op1_03_inv02 = 1;
    36: op1_03_inv02 = 1;
    40: op1_03_inv02 = 1;
    44: op1_03_inv02 = 1;
    50: op1_03_inv02 = 1;
    51: op1_03_inv02 = 1;
    52: op1_03_inv02 = 1;
    53: op1_03_inv02 = 1;
    54: op1_03_inv02 = 1;
    55: op1_03_inv02 = 1;
    56: op1_03_inv02 = 1;
    60: op1_03_inv02 = 1;
    62: op1_03_inv02 = 1;
    63: op1_03_inv02 = 1;
    65: op1_03_inv02 = 1;
    67: op1_03_inv02 = 1;
    69: op1_03_inv02 = 1;
    71: op1_03_inv02 = 1;
    72: op1_03_inv02 = 1;
    73: op1_03_inv02 = 1;
    75: op1_03_inv02 = 1;
    77: op1_03_inv02 = 1;
    78: op1_03_inv02 = 1;
    79: op1_03_inv02 = 1;
    80: op1_03_inv02 = 1;
    82: op1_03_inv02 = 1;
    83: op1_03_inv02 = 1;
    84: op1_03_inv02 = 1;
    87: op1_03_inv02 = 1;
    89: op1_03_inv02 = 1;
    92: op1_03_inv02 = 1;
    93: op1_03_inv02 = 1;
    94: op1_03_inv02 = 1;
    96: op1_03_inv02 = 1;
    default: op1_03_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in03 = reg_0276;
    6: op1_03_in03 = imem02_in[7:4];
    66: op1_03_in03 = imem02_in[7:4];
    7: op1_03_in03 = imem06_in[43:40];
    8: op1_03_in03 = imem02_in[27:24];
    9: op1_03_in03 = imem04_in[115:112];
    10: op1_03_in03 = reg_0293;
    4: op1_03_in03 = imem07_in[87:84];
    3: op1_03_in03 = imem07_in[107:104];
    11: op1_03_in03 = reg_0260;
    12: op1_03_in03 = reg_0384;
    13: op1_03_in03 = reg_0215;
    14: op1_03_in03 = imem02_in[11:8];
    15: op1_03_in03 = imem04_in[67:64];
    16: op1_03_in03 = reg_0128;
    17: op1_03_in03 = reg_0683;
    63: op1_03_in03 = reg_0683;
    18: op1_03_in03 = reg_0050;
    19: op1_03_in03 = reg_0111;
    20: op1_03_in03 = reg_1000;
    21: op1_03_in03 = reg_0684;
    22: op1_03_in03 = reg_0361;
    23: op1_03_in03 = imem05_in[55:52];
    24: op1_03_in03 = reg_0345;
    25: op1_03_in03 = reg_0609;
    26: op1_03_in03 = imem00_in[39:36];
    27: op1_03_in03 = reg_0610;
    28: op1_03_in03 = reg_0690;
    29: op1_03_in03 = imem04_in[63:60];
    35: op1_03_in03 = imem04_in[63:60];
    30: op1_03_in03 = imem05_in[91:88];
    31: op1_03_in03 = imem00_in[75:72];
    32: op1_03_in03 = imem03_in[51:48];
    36: op1_03_in03 = imem03_in[51:48];
    33: op1_03_in03 = reg_0076;
    34: op1_03_in03 = reg_0392;
    37: op1_03_in03 = reg_0537;
    38: op1_03_in03 = reg_0285;
    39: op1_03_in03 = reg_0043;
    40: op1_03_in03 = reg_0163;
    41: op1_03_in03 = imem06_in[127:124];
    42: op1_03_in03 = reg_0798;
    43: op1_03_in03 = reg_0833;
    44: op1_03_in03 = reg_0961;
    45: op1_03_in03 = imem00_in[91:88];
    46: op1_03_in03 = reg_0649;
    47: op1_03_in03 = reg_0963;
    48: op1_03_in03 = reg_0407;
    49: op1_03_in03 = reg_0365;
    50: op1_03_in03 = reg_1035;
    51: op1_03_in03 = imem00_in[127:124];
    52: op1_03_in03 = reg_0594;
    53: op1_03_in03 = reg_0168;
    54: op1_03_in03 = imem00_in[111:108];
    55: op1_03_in03 = imem01_in[23:20];
    56: op1_03_in03 = reg_0555;
    57: op1_03_in03 = reg_0346;
    58: op1_03_in03 = reg_0369;
    59: op1_03_in03 = reg_0733;
    67: op1_03_in03 = reg_0733;
    60: op1_03_in03 = reg_0269;
    61: op1_03_in03 = imem04_in[51:48];
    62: op1_03_in03 = imem05_in[111:108];
    64: op1_03_in03 = reg_0465;
    65: op1_03_in03 = reg_0522;
    68: op1_03_in03 = reg_0036;
    69: op1_03_in03 = imem07_in[111:108];
    70: op1_03_in03 = imem00_in[123:120];
    71: op1_03_in03 = reg_0084;
    72: op1_03_in03 = imem00_in[79:76];
    87: op1_03_in03 = imem00_in[79:76];
    73: op1_03_in03 = reg_1039;
    74: op1_03_in03 = imem02_in[79:76];
    75: op1_03_in03 = reg_0046;
    76: op1_03_in03 = imem06_in[123:120];
    77: op1_03_in03 = reg_0706;
    79: op1_03_in03 = reg_1017;
    80: op1_03_in03 = reg_0763;
    81: op1_03_in03 = reg_0998;
    82: op1_03_in03 = reg_0307;
    83: op1_03_in03 = reg_0724;
    84: op1_03_in03 = reg_0965;
    94: op1_03_in03 = reg_0965;
    85: op1_03_in03 = reg_0117;
    86: op1_03_in03 = imem04_in[103:100];
    88: op1_03_in03 = reg_0680;
    89: op1_03_in03 = reg_0405;
    90: op1_03_in03 = reg_0334;
    91: op1_03_in03 = imem02_in[99:96];
    92: op1_03_in03 = reg_0441;
    93: op1_03_in03 = imem06_in[83:80];
    95: op1_03_in03 = reg_0530;
    96: op1_03_in03 = reg_0950;
    97: op1_03_in03 = imem04_in[31:28];
    default: op1_03_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv03 = 1;
    6: op1_03_inv03 = 1;
    10: op1_03_inv03 = 1;
    3: op1_03_inv03 = 1;
    13: op1_03_inv03 = 1;
    15: op1_03_inv03 = 1;
    17: op1_03_inv03 = 1;
    19: op1_03_inv03 = 1;
    20: op1_03_inv03 = 1;
    22: op1_03_inv03 = 1;
    23: op1_03_inv03 = 1;
    27: op1_03_inv03 = 1;
    29: op1_03_inv03 = 1;
    30: op1_03_inv03 = 1;
    31: op1_03_inv03 = 1;
    33: op1_03_inv03 = 1;
    34: op1_03_inv03 = 1;
    35: op1_03_inv03 = 1;
    36: op1_03_inv03 = 1;
    39: op1_03_inv03 = 1;
    40: op1_03_inv03 = 1;
    44: op1_03_inv03 = 1;
    45: op1_03_inv03 = 1;
    46: op1_03_inv03 = 1;
    47: op1_03_inv03 = 1;
    48: op1_03_inv03 = 1;
    50: op1_03_inv03 = 1;
    51: op1_03_inv03 = 1;
    53: op1_03_inv03 = 1;
    54: op1_03_inv03 = 1;
    56: op1_03_inv03 = 1;
    57: op1_03_inv03 = 1;
    59: op1_03_inv03 = 1;
    60: op1_03_inv03 = 1;
    61: op1_03_inv03 = 1;
    62: op1_03_inv03 = 1;
    63: op1_03_inv03 = 1;
    65: op1_03_inv03 = 1;
    67: op1_03_inv03 = 1;
    68: op1_03_inv03 = 1;
    71: op1_03_inv03 = 1;
    72: op1_03_inv03 = 1;
    74: op1_03_inv03 = 1;
    77: op1_03_inv03 = 1;
    79: op1_03_inv03 = 1;
    81: op1_03_inv03 = 1;
    83: op1_03_inv03 = 1;
    84: op1_03_inv03 = 1;
    86: op1_03_inv03 = 1;
    87: op1_03_inv03 = 1;
    90: op1_03_inv03 = 1;
    91: op1_03_inv03 = 1;
    94: op1_03_inv03 = 1;
    97: op1_03_inv03 = 1;
    default: op1_03_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in04 = reg_0288;
    6: op1_03_in04 = reg_0653;
    7: op1_03_in04 = imem06_in[79:76];
    8: op1_03_in04 = imem02_in[51:48];
    9: op1_03_in04 = reg_0550;
    10: op1_03_in04 = reg_0285;
    4: op1_03_in04 = imem07_in[95:92];
    3: op1_03_in04 = imem07_in[111:108];
    11: op1_03_in04 = reg_0272;
    12: op1_03_in04 = reg_0388;
    13: op1_03_in04 = reg_0908;
    14: op1_03_in04 = imem02_in[27:24];
    66: op1_03_in04 = imem02_in[27:24];
    15: op1_03_in04 = imem04_in[83:80];
    16: op1_03_in04 = reg_0129;
    17: op1_03_in04 = reg_0672;
    18: op1_03_in04 = reg_0542;
    19: op1_03_in04 = reg_0119;
    20: op1_03_in04 = reg_0994;
    21: op1_03_in04 = reg_0481;
    22: op1_03_in04 = reg_0331;
    23: op1_03_in04 = imem05_in[67:64];
    24: op1_03_in04 = reg_0355;
    25: op1_03_in04 = reg_0618;
    26: op1_03_in04 = imem00_in[47:44];
    27: op1_03_in04 = reg_0631;
    28: op1_03_in04 = reg_0678;
    29: op1_03_in04 = imem04_in[79:76];
    35: op1_03_in04 = imem04_in[79:76];
    30: op1_03_in04 = imem05_in[95:92];
    31: op1_03_in04 = imem00_in[107:104];
    32: op1_03_in04 = imem03_in[59:56];
    36: op1_03_in04 = imem03_in[59:56];
    33: op1_03_in04 = reg_0063;
    34: op1_03_in04 = reg_0391;
    37: op1_03_in04 = reg_0733;
    38: op1_03_in04 = reg_0044;
    39: op1_03_in04 = imem05_in[15:12];
    40: op1_03_in04 = reg_0166;
    41: op1_03_in04 = reg_0073;
    42: op1_03_in04 = reg_0500;
    43: op1_03_in04 = reg_0040;
    44: op1_03_in04 = reg_0947;
    45: op1_03_in04 = imem00_in[103:100];
    46: op1_03_in04 = reg_0656;
    47: op1_03_in04 = reg_0951;
    48: op1_03_in04 = reg_0020;
    49: op1_03_in04 = reg_0643;
    80: op1_03_in04 = reg_0643;
    50: op1_03_in04 = reg_1045;
    51: op1_03_in04 = reg_0682;
    70: op1_03_in04 = reg_0682;
    52: op1_03_in04 = reg_0241;
    53: op1_03_in04 = reg_0158;
    54: op1_03_in04 = imem00_in[123:120];
    55: op1_03_in04 = imem01_in[59:56];
    56: op1_03_in04 = reg_0827;
    67: op1_03_in04 = reg_0827;
    57: op1_03_in04 = reg_0396;
    58: op1_03_in04 = reg_0234;
    59: op1_03_in04 = reg_0101;
    60: op1_03_in04 = reg_0233;
    61: op1_03_in04 = imem04_in[67:64];
    62: op1_03_in04 = imem05_in[127:124];
    63: op1_03_in04 = reg_0900;
    64: op1_03_in04 = reg_0455;
    65: op1_03_in04 = reg_0604;
    73: op1_03_in04 = reg_0604;
    68: op1_03_in04 = reg_0565;
    69: op1_03_in04 = imem07_in[119:116];
    71: op1_03_in04 = reg_0079;
    72: op1_03_in04 = reg_0683;
    74: op1_03_in04 = imem02_in[87:84];
    75: op1_03_in04 = reg_0571;
    76: op1_03_in04 = reg_0691;
    77: op1_03_in04 = reg_0657;
    79: op1_03_in04 = reg_0769;
    81: op1_03_in04 = reg_0978;
    82: op1_03_in04 = reg_0662;
    83: op1_03_in04 = reg_0184;
    84: op1_03_in04 = imem06_in[15:12];
    85: op1_03_in04 = reg_0352;
    86: op1_03_in04 = reg_0577;
    87: op1_03_in04 = imem00_in[83:80];
    88: op1_03_in04 = reg_0469;
    89: op1_03_in04 = reg_0937;
    90: op1_03_in04 = reg_0666;
    91: op1_03_in04 = reg_0255;
    92: op1_03_in04 = reg_0425;
    93: op1_03_in04 = imem06_in[91:88];
    94: op1_03_in04 = reg_0851;
    95: op1_03_in04 = reg_0019;
    96: op1_03_in04 = imem06_in[11:8];
    97: op1_03_in04 = imem04_in[71:68];
    default: op1_03_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_03_inv04 = 1;
    10: op1_03_inv04 = 1;
    4: op1_03_inv04 = 1;
    3: op1_03_inv04 = 1;
    11: op1_03_inv04 = 1;
    14: op1_03_inv04 = 1;
    16: op1_03_inv04 = 1;
    22: op1_03_inv04 = 1;
    25: op1_03_inv04 = 1;
    26: op1_03_inv04 = 1;
    27: op1_03_inv04 = 1;
    29: op1_03_inv04 = 1;
    31: op1_03_inv04 = 1;
    32: op1_03_inv04 = 1;
    33: op1_03_inv04 = 1;
    34: op1_03_inv04 = 1;
    36: op1_03_inv04 = 1;
    37: op1_03_inv04 = 1;
    39: op1_03_inv04 = 1;
    40: op1_03_inv04 = 1;
    43: op1_03_inv04 = 1;
    45: op1_03_inv04 = 1;
    46: op1_03_inv04 = 1;
    49: op1_03_inv04 = 1;
    51: op1_03_inv04 = 1;
    52: op1_03_inv04 = 1;
    53: op1_03_inv04 = 1;
    56: op1_03_inv04 = 1;
    59: op1_03_inv04 = 1;
    61: op1_03_inv04 = 1;
    62: op1_03_inv04 = 1;
    66: op1_03_inv04 = 1;
    67: op1_03_inv04 = 1;
    70: op1_03_inv04 = 1;
    72: op1_03_inv04 = 1;
    73: op1_03_inv04 = 1;
    77: op1_03_inv04 = 1;
    79: op1_03_inv04 = 1;
    80: op1_03_inv04 = 1;
    86: op1_03_inv04 = 1;
    88: op1_03_inv04 = 1;
    89: op1_03_inv04 = 1;
    90: op1_03_inv04 = 1;
    92: op1_03_inv04 = 1;
    93: op1_03_inv04 = 1;
    96: op1_03_inv04 = 1;
    97: op1_03_inv04 = 1;
    default: op1_03_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in05 = reg_0061;
    6: op1_03_in05 = reg_0638;
    7: op1_03_in05 = imem06_in[103:100];
    8: op1_03_in05 = imem02_in[55:52];
    9: op1_03_in05 = reg_0555;
    10: op1_03_in05 = reg_0292;
    4: op1_03_in05 = imem07_in[103:100];
    3: op1_03_in05 = imem07_in[115:112];
    11: op1_03_in05 = reg_0261;
    12: op1_03_in05 = reg_0393;
    76: op1_03_in05 = reg_0393;
    13: op1_03_in05 = reg_0251;
    14: op1_03_in05 = imem02_in[47:44];
    15: op1_03_in05 = imem04_in[91:88];
    16: op1_03_in05 = reg_0153;
    17: op1_03_in05 = reg_0676;
    18: op1_03_in05 = reg_0534;
    19: op1_03_in05 = reg_0120;
    20: op1_03_in05 = imem04_in[11:8];
    21: op1_03_in05 = reg_0470;
    22: op1_03_in05 = reg_0996;
    23: op1_03_in05 = imem05_in[95:92];
    24: op1_03_in05 = reg_0335;
    25: op1_03_in05 = reg_0402;
    26: op1_03_in05 = imem00_in[75:72];
    27: op1_03_in05 = reg_0577;
    28: op1_03_in05 = reg_0688;
    29: op1_03_in05 = reg_0306;
    30: op1_03_in05 = imem05_in[115:112];
    31: op1_03_in05 = reg_0678;
    32: op1_03_in05 = imem03_in[99:96];
    33: op1_03_in05 = reg_0732;
    34: op1_03_in05 = reg_0390;
    35: op1_03_in05 = reg_0483;
    36: op1_03_in05 = imem03_in[63:60];
    37: op1_03_in05 = reg_0760;
    38: op1_03_in05 = imem05_in[7:4];
    39: op1_03_in05 = imem05_in[31:28];
    40: op1_03_in05 = reg_0164;
    41: op1_03_in05 = reg_0381;
    42: op1_03_in05 = reg_0902;
    43: op1_03_in05 = reg_0784;
    44: op1_03_in05 = reg_0953;
    47: op1_03_in05 = reg_0953;
    45: op1_03_in05 = imem00_in[107:104];
    46: op1_03_in05 = reg_0621;
    48: op1_03_in05 = reg_0611;
    49: op1_03_in05 = reg_0854;
    50: op1_03_in05 = reg_1052;
    51: op1_03_in05 = reg_0693;
    52: op1_03_in05 = reg_0605;
    54: op1_03_in05 = reg_0696;
    55: op1_03_in05 = imem01_in[95:92];
    56: op1_03_in05 = reg_0101;
    79: op1_03_in05 = reg_0101;
    57: op1_03_in05 = reg_0661;
    58: op1_03_in05 = reg_0979;
    59: op1_03_in05 = reg_0117;
    60: op1_03_in05 = reg_0826;
    61: op1_03_in05 = imem04_in[103:100];
    62: op1_03_in05 = reg_0940;
    63: op1_03_in05 = reg_0102;
    64: op1_03_in05 = reg_0466;
    65: op1_03_in05 = reg_1037;
    66: op1_03_in05 = imem02_in[43:40];
    67: op1_03_in05 = reg_0115;
    68: op1_03_in05 = reg_0648;
    69: op1_03_in05 = reg_0720;
    70: op1_03_in05 = reg_0519;
    71: op1_03_in05 = imem03_in[47:44];
    72: op1_03_in05 = reg_0069;
    73: op1_03_in05 = reg_0520;
    74: op1_03_in05 = imem02_in[99:96];
    75: op1_03_in05 = reg_0239;
    82: op1_03_in05 = reg_0239;
    77: op1_03_in05 = imem06_in[11:8];
    80: op1_03_in05 = reg_0323;
    81: op1_03_in05 = reg_0974;
    84: op1_03_in05 = imem06_in[31:28];
    85: op1_03_in05 = reg_0089;
    86: op1_03_in05 = reg_0511;
    87: op1_03_in05 = reg_0841;
    88: op1_03_in05 = reg_0460;
    89: op1_03_in05 = reg_0586;
    90: op1_03_in05 = reg_0536;
    91: op1_03_in05 = reg_0277;
    92: op1_03_in05 = reg_0818;
    93: op1_03_in05 = imem06_in[99:96];
    94: op1_03_in05 = reg_0657;
    95: op1_03_in05 = reg_0741;
    96: op1_03_in05 = imem06_in[51:48];
    97: op1_03_in05 = imem04_in[119:116];
    default: op1_03_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv05 = 1;
    6: op1_03_inv05 = 1;
    8: op1_03_inv05 = 1;
    9: op1_03_inv05 = 1;
    10: op1_03_inv05 = 1;
    11: op1_03_inv05 = 1;
    12: op1_03_inv05 = 1;
    13: op1_03_inv05 = 1;
    15: op1_03_inv05 = 1;
    16: op1_03_inv05 = 1;
    21: op1_03_inv05 = 1;
    25: op1_03_inv05 = 1;
    27: op1_03_inv05 = 1;
    29: op1_03_inv05 = 1;
    31: op1_03_inv05 = 1;
    32: op1_03_inv05 = 1;
    33: op1_03_inv05 = 1;
    35: op1_03_inv05 = 1;
    36: op1_03_inv05 = 1;
    37: op1_03_inv05 = 1;
    38: op1_03_inv05 = 1;
    40: op1_03_inv05 = 1;
    42: op1_03_inv05 = 1;
    45: op1_03_inv05 = 1;
    46: op1_03_inv05 = 1;
    47: op1_03_inv05 = 1;
    49: op1_03_inv05 = 1;
    50: op1_03_inv05 = 1;
    51: op1_03_inv05 = 1;
    52: op1_03_inv05 = 1;
    57: op1_03_inv05 = 1;
    60: op1_03_inv05 = 1;
    61: op1_03_inv05 = 1;
    62: op1_03_inv05 = 1;
    63: op1_03_inv05 = 1;
    64: op1_03_inv05 = 1;
    65: op1_03_inv05 = 1;
    67: op1_03_inv05 = 1;
    68: op1_03_inv05 = 1;
    69: op1_03_inv05 = 1;
    71: op1_03_inv05 = 1;
    72: op1_03_inv05 = 1;
    74: op1_03_inv05 = 1;
    75: op1_03_inv05 = 1;
    77: op1_03_inv05 = 1;
    79: op1_03_inv05 = 1;
    80: op1_03_inv05 = 1;
    81: op1_03_inv05 = 1;
    82: op1_03_inv05 = 1;
    85: op1_03_inv05 = 1;
    86: op1_03_inv05 = 1;
    89: op1_03_inv05 = 1;
    90: op1_03_inv05 = 1;
    91: op1_03_inv05 = 1;
    93: op1_03_inv05 = 1;
    95: op1_03_inv05 = 1;
    96: op1_03_inv05 = 1;
    97: op1_03_inv05 = 1;
    default: op1_03_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in06 = reg_0062;
    6: op1_03_in06 = reg_0643;
    7: op1_03_in06 = reg_0629;
    8: op1_03_in06 = imem02_in[111:108];
    9: op1_03_in06 = reg_0546;
    10: op1_03_in06 = reg_0286;
    4: op1_03_in06 = imem07_in[111:108];
    3: op1_03_in06 = reg_0174;
    11: op1_03_in06 = reg_0263;
    12: op1_03_in06 = reg_1001;
    13: op1_03_in06 = reg_0148;
    14: op1_03_in06 = imem02_in[71:68];
    15: op1_03_in06 = reg_0543;
    16: op1_03_in06 = reg_0140;
    17: op1_03_in06 = reg_0671;
    18: op1_03_in06 = reg_0304;
    19: op1_03_in06 = reg_0101;
    20: op1_03_in06 = imem04_in[23:20];
    21: op1_03_in06 = reg_0474;
    22: op1_03_in06 = reg_0989;
    23: op1_03_in06 = imem05_in[115:112];
    24: op1_03_in06 = reg_0088;
    25: op1_03_in06 = reg_0344;
    26: op1_03_in06 = imem00_in[127:124];
    27: op1_03_in06 = reg_0627;
    28: op1_03_in06 = reg_0699;
    29: op1_03_in06 = reg_0539;
    30: op1_03_in06 = reg_0956;
    31: op1_03_in06 = reg_0463;
    32: op1_03_in06 = imem03_in[119:116];
    33: op1_03_in06 = reg_0773;
    34: op1_03_in06 = reg_0594;
    35: op1_03_in06 = reg_1009;
    36: op1_03_in06 = imem03_in[67:64];
    37: op1_03_in06 = reg_0276;
    38: op1_03_in06 = imem05_in[19:16];
    39: op1_03_in06 = reg_0955;
    40: op1_03_in06 = reg_0176;
    41: op1_03_in06 = reg_0042;
    42: op1_03_in06 = reg_0737;
    65: op1_03_in06 = reg_0737;
    43: op1_03_in06 = reg_0234;
    44: op1_03_in06 = reg_1021;
    47: op1_03_in06 = reg_1021;
    45: op1_03_in06 = reg_0695;
    46: op1_03_in06 = reg_0854;
    48: op1_03_in06 = reg_0395;
    49: op1_03_in06 = reg_0334;
    50: op1_03_in06 = reg_0514;
    51: op1_03_in06 = reg_0676;
    52: op1_03_in06 = reg_0609;
    75: op1_03_in06 = reg_0609;
    54: op1_03_in06 = reg_0691;
    55: op1_03_in06 = imem01_in[99:96];
    56: op1_03_in06 = reg_0113;
    57: op1_03_in06 = reg_0793;
    58: op1_03_in06 = reg_0984;
    59: op1_03_in06 = imem02_in[43:40];
    60: op1_03_in06 = reg_0032;
    61: op1_03_in06 = reg_1006;
    62: op1_03_in06 = reg_0237;
    63: op1_03_in06 = reg_0680;
    64: op1_03_in06 = reg_0456;
    66: op1_03_in06 = imem02_in[87:84];
    67: op1_03_in06 = reg_0821;
    68: op1_03_in06 = reg_0908;
    69: op1_03_in06 = reg_0708;
    70: op1_03_in06 = reg_0843;
    71: op1_03_in06 = imem03_in[51:48];
    72: op1_03_in06 = reg_0102;
    73: op1_03_in06 = reg_1037;
    74: op1_03_in06 = reg_0916;
    76: op1_03_in06 = reg_0021;
    77: op1_03_in06 = imem06_in[67:64];
    79: op1_03_in06 = reg_0109;
    80: op1_03_in06 = reg_0368;
    81: op1_03_in06 = imem04_in[15:12];
    82: op1_03_in06 = reg_1008;
    84: op1_03_in06 = imem06_in[51:48];
    85: op1_03_in06 = reg_0308;
    86: op1_03_in06 = reg_0550;
    87: op1_03_in06 = reg_0519;
    88: op1_03_in06 = reg_0473;
    89: op1_03_in06 = reg_0537;
    90: op1_03_in06 = reg_0077;
    91: op1_03_in06 = reg_0837;
    92: op1_03_in06 = reg_0335;
    93: op1_03_in06 = imem06_in[103:100];
    94: op1_03_in06 = imem06_in[23:20];
    95: op1_03_in06 = imem06_in[75:72];
    96: op1_03_in06 = imem06_in[55:52];
    97: op1_03_in06 = imem04_in[123:120];
    default: op1_03_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv06 = 1;
    9: op1_03_inv06 = 1;
    4: op1_03_inv06 = 1;
    13: op1_03_inv06 = 1;
    14: op1_03_inv06 = 1;
    20: op1_03_inv06 = 1;
    22: op1_03_inv06 = 1;
    24: op1_03_inv06 = 1;
    28: op1_03_inv06 = 1;
    31: op1_03_inv06 = 1;
    37: op1_03_inv06 = 1;
    38: op1_03_inv06 = 1;
    39: op1_03_inv06 = 1;
    41: op1_03_inv06 = 1;
    42: op1_03_inv06 = 1;
    45: op1_03_inv06 = 1;
    50: op1_03_inv06 = 1;
    54: op1_03_inv06 = 1;
    56: op1_03_inv06 = 1;
    57: op1_03_inv06 = 1;
    58: op1_03_inv06 = 1;
    59: op1_03_inv06 = 1;
    60: op1_03_inv06 = 1;
    61: op1_03_inv06 = 1;
    65: op1_03_inv06 = 1;
    66: op1_03_inv06 = 1;
    68: op1_03_inv06 = 1;
    69: op1_03_inv06 = 1;
    70: op1_03_inv06 = 1;
    71: op1_03_inv06 = 1;
    72: op1_03_inv06 = 1;
    75: op1_03_inv06 = 1;
    77: op1_03_inv06 = 1;
    81: op1_03_inv06 = 1;
    82: op1_03_inv06 = 1;
    85: op1_03_inv06 = 1;
    86: op1_03_inv06 = 1;
    90: op1_03_inv06 = 1;
    92: op1_03_inv06 = 1;
    94: op1_03_inv06 = 1;
    95: op1_03_inv06 = 1;
    96: op1_03_inv06 = 1;
    default: op1_03_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in07 = reg_0048;
    29: op1_03_in07 = reg_0048;
    6: op1_03_in07 = reg_0325;
    7: op1_03_in07 = reg_0620;
    8: op1_03_in07 = imem02_in[115:112];
    9: op1_03_in07 = reg_0303;
    10: op1_03_in07 = reg_0062;
    4: op1_03_in07 = imem07_in[115:112];
    3: op1_03_in07 = reg_0158;
    11: op1_03_in07 = reg_0151;
    12: op1_03_in07 = reg_0993;
    13: op1_03_in07 = reg_0156;
    86: op1_03_in07 = reg_0156;
    14: op1_03_in07 = imem02_in[75:72];
    15: op1_03_in07 = reg_0544;
    16: op1_03_in07 = reg_0137;
    17: op1_03_in07 = reg_0688;
    18: op1_03_in07 = imem04_in[31:28];
    19: op1_03_in07 = reg_0126;
    20: op1_03_in07 = imem04_in[27:24];
    21: op1_03_in07 = reg_0191;
    22: op1_03_in07 = reg_0983;
    23: op1_03_in07 = imem05_in[127:124];
    24: op1_03_in07 = reg_0867;
    25: op1_03_in07 = reg_0381;
    26: op1_03_in07 = reg_0697;
    45: op1_03_in07 = reg_0697;
    27: op1_03_in07 = reg_0402;
    28: op1_03_in07 = reg_0463;
    72: op1_03_in07 = reg_0463;
    30: op1_03_in07 = reg_0968;
    31: op1_03_in07 = reg_0464;
    32: op1_03_in07 = reg_0317;
    33: op1_03_in07 = imem05_in[7:4];
    34: op1_03_in07 = reg_0405;
    35: op1_03_in07 = reg_1057;
    36: op1_03_in07 = reg_0394;
    37: op1_03_in07 = reg_0732;
    38: op1_03_in07 = imem05_in[27:24];
    39: op1_03_in07 = reg_0967;
    41: op1_03_in07 = reg_0351;
    42: op1_03_in07 = reg_0610;
    43: op1_03_in07 = reg_0987;
    44: op1_03_in07 = reg_0896;
    46: op1_03_in07 = reg_0558;
    47: op1_03_in07 = reg_0834;
    48: op1_03_in07 = reg_0914;
    49: op1_03_in07 = reg_0863;
    50: op1_03_in07 = reg_1041;
    65: op1_03_in07 = reg_1041;
    51: op1_03_in07 = reg_0686;
    52: op1_03_in07 = reg_0626;
    54: op1_03_in07 = reg_0450;
    55: op1_03_in07 = reg_0586;
    56: op1_03_in07 = imem02_in[19:16];
    57: op1_03_in07 = reg_0765;
    58: op1_03_in07 = reg_0996;
    59: op1_03_in07 = reg_0639;
    60: op1_03_in07 = reg_0446;
    61: op1_03_in07 = reg_0937;
    62: op1_03_in07 = reg_0448;
    63: op1_03_in07 = reg_0753;
    64: op1_03_in07 = reg_0478;
    66: op1_03_in07 = imem02_in[95:92];
    67: op1_03_in07 = reg_0745;
    68: op1_03_in07 = reg_0855;
    90: op1_03_in07 = reg_0855;
    69: op1_03_in07 = reg_0707;
    70: op1_03_in07 = reg_0102;
    71: op1_03_in07 = reg_0535;
    73: op1_03_in07 = reg_0902;
    74: op1_03_in07 = reg_0649;
    75: op1_03_in07 = reg_0588;
    76: op1_03_in07 = reg_0328;
    77: op1_03_in07 = imem06_in[99:96];
    79: op1_03_in07 = reg_0117;
    80: op1_03_in07 = reg_0425;
    81: op1_03_in07 = imem04_in[63:60];
    82: op1_03_in07 = reg_0266;
    84: op1_03_in07 = imem06_in[67:64];
    85: op1_03_in07 = reg_0750;
    87: op1_03_in07 = reg_0674;
    88: op1_03_in07 = reg_0467;
    89: op1_03_in07 = reg_0066;
    91: op1_03_in07 = reg_0645;
    92: op1_03_in07 = reg_0516;
    93: op1_03_in07 = reg_0625;
    94: op1_03_in07 = imem06_in[39:36];
    95: op1_03_in07 = imem06_in[83:80];
    96: op1_03_in07 = imem06_in[59:56];
    97: op1_03_in07 = reg_0942;
    default: op1_03_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv07 = 1;
    7: op1_03_inv07 = 1;
    9: op1_03_inv07 = 1;
    4: op1_03_inv07 = 1;
    12: op1_03_inv07 = 1;
    14: op1_03_inv07 = 1;
    18: op1_03_inv07 = 1;
    20: op1_03_inv07 = 1;
    21: op1_03_inv07 = 1;
    23: op1_03_inv07 = 1;
    29: op1_03_inv07 = 1;
    31: op1_03_inv07 = 1;
    33: op1_03_inv07 = 1;
    35: op1_03_inv07 = 1;
    37: op1_03_inv07 = 1;
    39: op1_03_inv07 = 1;
    42: op1_03_inv07 = 1;
    48: op1_03_inv07 = 1;
    49: op1_03_inv07 = 1;
    51: op1_03_inv07 = 1;
    59: op1_03_inv07 = 1;
    60: op1_03_inv07 = 1;
    61: op1_03_inv07 = 1;
    62: op1_03_inv07 = 1;
    65: op1_03_inv07 = 1;
    69: op1_03_inv07 = 1;
    70: op1_03_inv07 = 1;
    72: op1_03_inv07 = 1;
    73: op1_03_inv07 = 1;
    77: op1_03_inv07 = 1;
    81: op1_03_inv07 = 1;
    82: op1_03_inv07 = 1;
    84: op1_03_inv07 = 1;
    86: op1_03_inv07 = 1;
    87: op1_03_inv07 = 1;
    88: op1_03_inv07 = 1;
    90: op1_03_inv07 = 1;
    91: op1_03_inv07 = 1;
    94: op1_03_inv07 = 1;
    95: op1_03_inv07 = 1;
    97: op1_03_inv07 = 1;
    default: op1_03_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in08 = reg_0063;
    6: op1_03_in08 = reg_0326;
    7: op1_03_in08 = reg_0616;
    8: op1_03_in08 = reg_0660;
    9: op1_03_in08 = reg_0290;
    10: op1_03_in08 = reg_0056;
    4: op1_03_in08 = imem07_in[127:124];
    3: op1_03_in08 = reg_0171;
    11: op1_03_in08 = reg_0153;
    12: op1_03_in08 = reg_0980;
    13: op1_03_in08 = reg_0154;
    14: op1_03_in08 = imem02_in[83:80];
    15: op1_03_in08 = reg_0530;
    16: op1_03_in08 = reg_0134;
    17: op1_03_in08 = reg_0453;
    28: op1_03_in08 = reg_0453;
    18: op1_03_in08 = imem04_in[51:48];
    19: op1_03_in08 = reg_0110;
    65: op1_03_in08 = reg_0110;
    20: op1_03_in08 = imem04_in[67:64];
    21: op1_03_in08 = reg_0203;
    22: op1_03_in08 = imem04_in[39:36];
    23: op1_03_in08 = reg_0963;
    24: op1_03_in08 = reg_0484;
    25: op1_03_in08 = reg_0392;
    26: op1_03_in08 = reg_0685;
    27: op1_03_in08 = reg_0379;
    29: op1_03_in08 = reg_1020;
    30: op1_03_in08 = reg_0900;
    31: op1_03_in08 = reg_0472;
    32: op1_03_in08 = reg_1019;
    33: op1_03_in08 = imem05_in[11:8];
    34: op1_03_in08 = reg_0753;
    35: op1_03_in08 = reg_1016;
    36: op1_03_in08 = reg_0571;
    37: op1_03_in08 = reg_0864;
    38: op1_03_in08 = imem05_in[71:68];
    39: op1_03_in08 = reg_0954;
    41: op1_03_in08 = reg_0349;
    42: op1_03_in08 = reg_0925;
    43: op1_03_in08 = reg_0977;
    44: op1_03_in08 = reg_0128;
    45: op1_03_in08 = reg_0694;
    46: op1_03_in08 = reg_0045;
    47: op1_03_in08 = reg_0215;
    48: op1_03_in08 = reg_0351;
    93: op1_03_in08 = reg_0351;
    49: op1_03_in08 = reg_0080;
    50: op1_03_in08 = reg_0740;
    51: op1_03_in08 = reg_0691;
    52: op1_03_in08 = reg_0008;
    54: op1_03_in08 = reg_0477;
    72: op1_03_in08 = reg_0477;
    55: op1_03_in08 = reg_0274;
    56: op1_03_in08 = imem02_in[35:32];
    57: op1_03_in08 = reg_0509;
    58: op1_03_in08 = reg_1001;
    59: op1_03_in08 = reg_0651;
    60: op1_03_in08 = reg_0094;
    61: op1_03_in08 = reg_0055;
    62: op1_03_in08 = reg_1046;
    63: op1_03_in08 = reg_0465;
    64: op1_03_in08 = reg_0200;
    66: op1_03_in08 = reg_0905;
    67: op1_03_in08 = imem02_in[11:8];
    68: op1_03_in08 = reg_0424;
    69: op1_03_in08 = reg_0250;
    70: op1_03_in08 = reg_0669;
    71: op1_03_in08 = reg_0445;
    73: op1_03_in08 = reg_0737;
    74: op1_03_in08 = reg_0260;
    75: op1_03_in08 = reg_0233;
    76: op1_03_in08 = reg_0229;
    77: op1_03_in08 = reg_0817;
    79: op1_03_in08 = reg_0113;
    80: op1_03_in08 = reg_0248;
    81: op1_03_in08 = imem04_in[79:76];
    82: op1_03_in08 = reg_0551;
    84: op1_03_in08 = imem06_in[71:68];
    85: op1_03_in08 = reg_0844;
    86: op1_03_in08 = reg_0430;
    87: op1_03_in08 = reg_0102;
    88: op1_03_in08 = reg_0471;
    89: op1_03_in08 = reg_0276;
    90: op1_03_in08 = reg_0739;
    91: op1_03_in08 = reg_0664;
    92: op1_03_in08 = reg_0734;
    94: op1_03_in08 = imem06_in[79:76];
    95: op1_03_in08 = imem06_in[91:88];
    96: op1_03_in08 = reg_0696;
    97: op1_03_in08 = reg_0937;
    default: op1_03_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_03_inv08 = 1;
    4: op1_03_inv08 = 1;
    12: op1_03_inv08 = 1;
    13: op1_03_inv08 = 1;
    14: op1_03_inv08 = 1;
    15: op1_03_inv08 = 1;
    17: op1_03_inv08 = 1;
    20: op1_03_inv08 = 1;
    21: op1_03_inv08 = 1;
    24: op1_03_inv08 = 1;
    25: op1_03_inv08 = 1;
    26: op1_03_inv08 = 1;
    28: op1_03_inv08 = 1;
    29: op1_03_inv08 = 1;
    31: op1_03_inv08 = 1;
    33: op1_03_inv08 = 1;
    34: op1_03_inv08 = 1;
    35: op1_03_inv08 = 1;
    36: op1_03_inv08 = 1;
    37: op1_03_inv08 = 1;
    39: op1_03_inv08 = 1;
    41: op1_03_inv08 = 1;
    44: op1_03_inv08 = 1;
    48: op1_03_inv08 = 1;
    50: op1_03_inv08 = 1;
    51: op1_03_inv08 = 1;
    56: op1_03_inv08 = 1;
    57: op1_03_inv08 = 1;
    58: op1_03_inv08 = 1;
    59: op1_03_inv08 = 1;
    60: op1_03_inv08 = 1;
    63: op1_03_inv08 = 1;
    66: op1_03_inv08 = 1;
    67: op1_03_inv08 = 1;
    72: op1_03_inv08 = 1;
    73: op1_03_inv08 = 1;
    74: op1_03_inv08 = 1;
    75: op1_03_inv08 = 1;
    76: op1_03_inv08 = 1;
    77: op1_03_inv08 = 1;
    80: op1_03_inv08 = 1;
    81: op1_03_inv08 = 1;
    82: op1_03_inv08 = 1;
    85: op1_03_inv08 = 1;
    87: op1_03_inv08 = 1;
    89: op1_03_inv08 = 1;
    93: op1_03_inv08 = 1;
    95: op1_03_inv08 = 1;
    default: op1_03_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in09 = reg_0064;
    6: op1_03_in09 = reg_0354;
    7: op1_03_in09 = reg_0631;
    8: op1_03_in09 = reg_0353;
    9: op1_03_in09 = reg_0296;
    10: op1_03_in09 = reg_0043;
    4: op1_03_in09 = reg_0424;
    11: op1_03_in09 = reg_0141;
    13: op1_03_in09 = reg_0141;
    12: op1_03_in09 = reg_0978;
    58: op1_03_in09 = reg_0978;
    14: op1_03_in09 = imem02_in[103:100];
    15: op1_03_in09 = reg_0542;
    16: op1_03_in09 = imem06_in[7:4];
    17: op1_03_in09 = reg_0476;
    54: op1_03_in09 = reg_0476;
    70: op1_03_in09 = reg_0476;
    18: op1_03_in09 = imem04_in[63:60];
    19: op1_03_in09 = imem02_in[7:4];
    20: op1_03_in09 = imem04_in[75:72];
    21: op1_03_in09 = reg_0186;
    22: op1_03_in09 = imem04_in[79:76];
    23: op1_03_in09 = reg_0942;
    24: op1_03_in09 = reg_0291;
    25: op1_03_in09 = reg_0351;
    26: op1_03_in09 = reg_0676;
    27: op1_03_in09 = reg_0381;
    28: op1_03_in09 = reg_0451;
    29: op1_03_in09 = reg_1016;
    30: op1_03_in09 = reg_0244;
    31: op1_03_in09 = reg_0470;
    32: op1_03_in09 = reg_1049;
    36: op1_03_in09 = reg_1049;
    33: op1_03_in09 = imem05_in[27:24];
    34: op1_03_in09 = reg_0011;
    77: op1_03_in09 = reg_0011;
    35: op1_03_in09 = reg_0076;
    37: op1_03_in09 = imem05_in[19:16];
    38: op1_03_in09 = imem05_in[99:96];
    39: op1_03_in09 = reg_0950;
    41: op1_03_in09 = reg_0222;
    42: op1_03_in09 = reg_0120;
    43: op1_03_in09 = reg_0975;
    44: op1_03_in09 = reg_0129;
    45: op1_03_in09 = reg_0691;
    46: op1_03_in09 = reg_0096;
    47: op1_03_in09 = reg_1046;
    48: op1_03_in09 = reg_0243;
    49: op1_03_in09 = reg_0817;
    50: op1_03_in09 = reg_1017;
    51: op1_03_in09 = reg_0674;
    52: op1_03_in09 = reg_0029;
    55: op1_03_in09 = reg_0871;
    56: op1_03_in09 = imem02_in[75:72];
    57: op1_03_in09 = reg_0807;
    59: op1_03_in09 = reg_0652;
    60: op1_03_in09 = reg_0404;
    61: op1_03_in09 = reg_0540;
    62: op1_03_in09 = reg_0148;
    63: op1_03_in09 = reg_0457;
    64: op1_03_in09 = reg_0203;
    65: op1_03_in09 = imem02_in[3:0];
    66: op1_03_in09 = reg_0899;
    67: op1_03_in09 = imem02_in[35:32];
    68: op1_03_in09 = reg_0329;
    69: op1_03_in09 = reg_0047;
    71: op1_03_in09 = reg_0585;
    72: op1_03_in09 = reg_0462;
    73: op1_03_in09 = reg_0232;
    74: op1_03_in09 = reg_0095;
    75: op1_03_in09 = reg_0266;
    76: op1_03_in09 = reg_0889;
    79: op1_03_in09 = imem02_in[11:8];
    80: op1_03_in09 = reg_0087;
    81: op1_03_in09 = imem04_in[95:92];
    82: op1_03_in09 = reg_0991;
    84: op1_03_in09 = imem06_in[79:76];
    85: op1_03_in09 = reg_0554;
    86: op1_03_in09 = reg_0031;
    87: op1_03_in09 = reg_0450;
    88: op1_03_in09 = reg_0208;
    89: op1_03_in09 = reg_0584;
    90: op1_03_in09 = reg_0081;
    91: op1_03_in09 = reg_0372;
    92: op1_03_in09 = reg_0778;
    93: op1_03_in09 = reg_0393;
    94: op1_03_in09 = reg_1019;
    95: op1_03_in09 = imem06_in[107:104];
    96: op1_03_in09 = reg_0391;
    97: op1_03_in09 = reg_0912;
    default: op1_03_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv09 = 1;
    6: op1_03_inv09 = 1;
    11: op1_03_inv09 = 1;
    14: op1_03_inv09 = 1;
    15: op1_03_inv09 = 1;
    18: op1_03_inv09 = 1;
    19: op1_03_inv09 = 1;
    20: op1_03_inv09 = 1;
    21: op1_03_inv09 = 1;
    23: op1_03_inv09 = 1;
    24: op1_03_inv09 = 1;
    25: op1_03_inv09 = 1;
    27: op1_03_inv09 = 1;
    29: op1_03_inv09 = 1;
    30: op1_03_inv09 = 1;
    31: op1_03_inv09 = 1;
    32: op1_03_inv09 = 1;
    34: op1_03_inv09 = 1;
    37: op1_03_inv09 = 1;
    38: op1_03_inv09 = 1;
    39: op1_03_inv09 = 1;
    41: op1_03_inv09 = 1;
    42: op1_03_inv09 = 1;
    45: op1_03_inv09 = 1;
    46: op1_03_inv09 = 1;
    47: op1_03_inv09 = 1;
    52: op1_03_inv09 = 1;
    54: op1_03_inv09 = 1;
    55: op1_03_inv09 = 1;
    56: op1_03_inv09 = 1;
    57: op1_03_inv09 = 1;
    64: op1_03_inv09 = 1;
    65: op1_03_inv09 = 1;
    67: op1_03_inv09 = 1;
    69: op1_03_inv09 = 1;
    72: op1_03_inv09 = 1;
    73: op1_03_inv09 = 1;
    74: op1_03_inv09 = 1;
    75: op1_03_inv09 = 1;
    76: op1_03_inv09 = 1;
    77: op1_03_inv09 = 1;
    80: op1_03_inv09 = 1;
    84: op1_03_inv09 = 1;
    85: op1_03_inv09 = 1;
    86: op1_03_inv09 = 1;
    87: op1_03_inv09 = 1;
    95: op1_03_inv09 = 1;
    96: op1_03_inv09 = 1;
    default: op1_03_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in10 = imem05_in[23:20];
    6: op1_03_in10 = reg_0355;
    7: op1_03_in10 = reg_0632;
    8: op1_03_in10 = reg_0350;
    9: op1_03_in10 = reg_0298;
    10: op1_03_in10 = reg_0053;
    4: op1_03_in10 = reg_0446;
    11: op1_03_in10 = reg_0140;
    12: op1_03_in10 = reg_0975;
    13: op1_03_in10 = reg_0130;
    14: op1_03_in10 = reg_0660;
    95: op1_03_in10 = reg_0660;
    15: op1_03_in10 = reg_0548;
    16: op1_03_in10 = imem06_in[47:44];
    17: op1_03_in10 = reg_0470;
    54: op1_03_in10 = reg_0470;
    18: op1_03_in10 = imem04_in[67:64];
    19: op1_03_in10 = imem02_in[11:8];
    20: op1_03_in10 = imem04_in[91:88];
    21: op1_03_in10 = imem01_in[59:56];
    22: op1_03_in10 = imem04_in[83:80];
    23: op1_03_in10 = reg_0952;
    24: op1_03_in10 = reg_0872;
    25: op1_03_in10 = reg_0375;
    26: op1_03_in10 = reg_0466;
    27: op1_03_in10 = reg_0408;
    28: op1_03_in10 = reg_0455;
    87: op1_03_in10 = reg_0455;
    29: op1_03_in10 = reg_0541;
    30: op1_03_in10 = reg_0142;
    31: op1_03_in10 = reg_0474;
    32: op1_03_in10 = reg_0327;
    33: op1_03_in10 = imem05_in[67:64];
    34: op1_03_in10 = imem07_in[23:20];
    35: op1_03_in10 = reg_0009;
    36: op1_03_in10 = reg_0046;
    37: op1_03_in10 = imem05_in[35:32];
    38: op1_03_in10 = reg_0973;
    39: op1_03_in10 = reg_0968;
    41: op1_03_in10 = reg_0000;
    42: op1_03_in10 = reg_0117;
    43: op1_03_in10 = reg_0983;
    44: op1_03_in10 = reg_0153;
    45: op1_03_in10 = reg_0673;
    46: op1_03_in10 = reg_0225;
    47: op1_03_in10 = reg_0832;
    48: op1_03_in10 = reg_0399;
    49: op1_03_in10 = reg_0758;
    50: op1_03_in10 = reg_0925;
    51: op1_03_in10 = reg_0692;
    52: op1_03_in10 = reg_0926;
    55: op1_03_in10 = reg_1052;
    56: op1_03_in10 = imem02_in[111:108];
    57: op1_03_in10 = reg_0991;
    58: op1_03_in10 = reg_0989;
    59: op1_03_in10 = reg_0418;
    60: op1_03_in10 = reg_0819;
    61: op1_03_in10 = reg_0799;
    86: op1_03_in10 = reg_0799;
    62: op1_03_in10 = reg_0135;
    63: op1_03_in10 = reg_0464;
    64: op1_03_in10 = reg_0213;
    65: op1_03_in10 = imem02_in[55:52];
    66: op1_03_in10 = reg_0845;
    67: op1_03_in10 = reg_0741;
    68: op1_03_in10 = reg_0085;
    69: op1_03_in10 = reg_0406;
    70: op1_03_in10 = reg_0187;
    71: op1_03_in10 = reg_0571;
    72: op1_03_in10 = reg_0472;
    73: op1_03_in10 = reg_0003;
    74: op1_03_in10 = reg_0424;
    75: op1_03_in10 = reg_0996;
    76: op1_03_in10 = reg_0297;
    77: op1_03_in10 = reg_0755;
    79: op1_03_in10 = imem02_in[71:68];
    80: op1_03_in10 = reg_0335;
    81: op1_03_in10 = reg_0536;
    82: op1_03_in10 = reg_0979;
    84: op1_03_in10 = imem06_in[87:84];
    85: op1_03_in10 = reg_0483;
    88: op1_03_in10 = reg_0207;
    89: op1_03_in10 = reg_0288;
    90: op1_03_in10 = reg_0441;
    91: op1_03_in10 = reg_0037;
    92: op1_03_in10 = reg_0730;
    93: op1_03_in10 = reg_0817;
    94: op1_03_in10 = reg_0025;
    96: op1_03_in10 = reg_0025;
    97: op1_03_in10 = reg_0224;
    default: op1_03_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv10 = 1;
    8: op1_03_inv10 = 1;
    9: op1_03_inv10 = 1;
    4: op1_03_inv10 = 1;
    11: op1_03_inv10 = 1;
    13: op1_03_inv10 = 1;
    15: op1_03_inv10 = 1;
    17: op1_03_inv10 = 1;
    18: op1_03_inv10 = 1;
    19: op1_03_inv10 = 1;
    20: op1_03_inv10 = 1;
    21: op1_03_inv10 = 1;
    22: op1_03_inv10 = 1;
    23: op1_03_inv10 = 1;
    25: op1_03_inv10 = 1;
    29: op1_03_inv10 = 1;
    30: op1_03_inv10 = 1;
    32: op1_03_inv10 = 1;
    35: op1_03_inv10 = 1;
    38: op1_03_inv10 = 1;
    39: op1_03_inv10 = 1;
    43: op1_03_inv10 = 1;
    45: op1_03_inv10 = 1;
    47: op1_03_inv10 = 1;
    52: op1_03_inv10 = 1;
    55: op1_03_inv10 = 1;
    57: op1_03_inv10 = 1;
    58: op1_03_inv10 = 1;
    60: op1_03_inv10 = 1;
    61: op1_03_inv10 = 1;
    63: op1_03_inv10 = 1;
    65: op1_03_inv10 = 1;
    66: op1_03_inv10 = 1;
    68: op1_03_inv10 = 1;
    70: op1_03_inv10 = 1;
    71: op1_03_inv10 = 1;
    72: op1_03_inv10 = 1;
    73: op1_03_inv10 = 1;
    74: op1_03_inv10 = 1;
    75: op1_03_inv10 = 1;
    76: op1_03_inv10 = 1;
    86: op1_03_inv10 = 1;
    88: op1_03_inv10 = 1;
    89: op1_03_inv10 = 1;
    95: op1_03_inv10 = 1;
    96: op1_03_inv10 = 1;
    97: op1_03_inv10 = 1;
    default: op1_03_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in11 = reg_0482;
    6: op1_03_in11 = reg_0335;
    7: op1_03_in11 = reg_0351;
    8: op1_03_in11 = reg_0083;
    9: op1_03_in11 = reg_0307;
    10: op1_03_in11 = reg_0063;
    4: op1_03_in11 = reg_0174;
    11: op1_03_in11 = reg_0131;
    12: op1_03_in11 = reg_1000;
    13: op1_03_in11 = reg_0137;
    14: op1_03_in11 = reg_0661;
    15: op1_03_in11 = reg_0558;
    16: op1_03_in11 = imem06_in[115:112];
    17: op1_03_in11 = reg_0456;
    72: op1_03_in11 = reg_0456;
    18: op1_03_in11 = imem04_in[79:76];
    19: op1_03_in11 = imem02_in[91:88];
    65: op1_03_in11 = imem02_in[91:88];
    20: op1_03_in11 = reg_0557;
    21: op1_03_in11 = imem01_in[67:64];
    22: op1_03_in11 = imem04_in[95:92];
    23: op1_03_in11 = reg_0943;
    24: op1_03_in11 = imem03_in[59:56];
    92: op1_03_in11 = imem03_in[59:56];
    25: op1_03_in11 = reg_0390;
    26: op1_03_in11 = reg_0475;
    27: op1_03_in11 = reg_0386;
    28: op1_03_in11 = reg_0476;
    29: op1_03_in11 = reg_0072;
    30: op1_03_in11 = reg_0156;
    31: op1_03_in11 = reg_0459;
    32: op1_03_in11 = reg_0046;
    33: op1_03_in11 = reg_0971;
    38: op1_03_in11 = reg_0971;
    34: op1_03_in11 = imem07_in[27:24];
    35: op1_03_in11 = reg_0525;
    36: op1_03_in11 = reg_0923;
    37: op1_03_in11 = imem05_in[51:48];
    39: op1_03_in11 = reg_0965;
    41: op1_03_in11 = reg_0332;
    42: op1_03_in11 = reg_0126;
    43: op1_03_in11 = imem04_in[47:44];
    44: op1_03_in11 = imem06_in[31:28];
    45: op1_03_in11 = reg_0699;
    46: op1_03_in11 = reg_0338;
    47: op1_03_in11 = reg_0831;
    48: op1_03_in11 = reg_0804;
    49: op1_03_in11 = reg_0089;
    50: op1_03_in11 = reg_0111;
    51: op1_03_in11 = reg_0465;
    52: op1_03_in11 = imem07_in[23:20];
    54: op1_03_in11 = reg_0207;
    55: op1_03_in11 = reg_0238;
    56: op1_03_in11 = imem02_in[123:120];
    57: op1_03_in11 = reg_0984;
    58: op1_03_in11 = reg_0988;
    59: op1_03_in11 = reg_0329;
    60: op1_03_in11 = reg_0136;
    61: op1_03_in11 = reg_0524;
    62: op1_03_in11 = reg_0138;
    63: op1_03_in11 = reg_0477;
    64: op1_03_in11 = reg_0205;
    66: op1_03_in11 = reg_0260;
    67: op1_03_in11 = reg_0666;
    68: op1_03_in11 = reg_0876;
    69: op1_03_in11 = reg_0419;
    70: op1_03_in11 = reg_0193;
    71: op1_03_in11 = reg_0281;
    73: op1_03_in11 = reg_0273;
    74: op1_03_in11 = reg_0052;
    75: op1_03_in11 = reg_0989;
    76: op1_03_in11 = reg_0395;
    77: op1_03_in11 = reg_0018;
    79: op1_03_in11 = imem02_in[75:72];
    80: op1_03_in11 = reg_0007;
    81: op1_03_in11 = reg_0048;
    82: op1_03_in11 = reg_0980;
    84: op1_03_in11 = imem06_in[103:100];
    85: op1_03_in11 = reg_0077;
    86: op1_03_in11 = reg_0848;
    87: op1_03_in11 = reg_0469;
    88: op1_03_in11 = reg_0211;
    89: op1_03_in11 = reg_0041;
    90: op1_03_in11 = reg_0425;
    91: op1_03_in11 = reg_0885;
    93: op1_03_in11 = reg_0889;
    94: op1_03_in11 = reg_0328;
    95: op1_03_in11 = reg_1019;
    96: op1_03_in11 = reg_0626;
    97: op1_03_in11 = reg_0292;
    default: op1_03_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_03_inv11 = 1;
    10: op1_03_inv11 = 1;
    11: op1_03_inv11 = 1;
    12: op1_03_inv11 = 1;
    14: op1_03_inv11 = 1;
    15: op1_03_inv11 = 1;
    17: op1_03_inv11 = 1;
    19: op1_03_inv11 = 1;
    20: op1_03_inv11 = 1;
    24: op1_03_inv11 = 1;
    26: op1_03_inv11 = 1;
    30: op1_03_inv11 = 1;
    31: op1_03_inv11 = 1;
    33: op1_03_inv11 = 1;
    36: op1_03_inv11 = 1;
    37: op1_03_inv11 = 1;
    39: op1_03_inv11 = 1;
    41: op1_03_inv11 = 1;
    43: op1_03_inv11 = 1;
    45: op1_03_inv11 = 1;
    46: op1_03_inv11 = 1;
    47: op1_03_inv11 = 1;
    49: op1_03_inv11 = 1;
    50: op1_03_inv11 = 1;
    51: op1_03_inv11 = 1;
    54: op1_03_inv11 = 1;
    57: op1_03_inv11 = 1;
    59: op1_03_inv11 = 1;
    60: op1_03_inv11 = 1;
    62: op1_03_inv11 = 1;
    63: op1_03_inv11 = 1;
    64: op1_03_inv11 = 1;
    66: op1_03_inv11 = 1;
    68: op1_03_inv11 = 1;
    69: op1_03_inv11 = 1;
    71: op1_03_inv11 = 1;
    72: op1_03_inv11 = 1;
    74: op1_03_inv11 = 1;
    76: op1_03_inv11 = 1;
    79: op1_03_inv11 = 1;
    80: op1_03_inv11 = 1;
    81: op1_03_inv11 = 1;
    82: op1_03_inv11 = 1;
    84: op1_03_inv11 = 1;
    89: op1_03_inv11 = 1;
    90: op1_03_inv11 = 1;
    91: op1_03_inv11 = 1;
    92: op1_03_inv11 = 1;
    default: op1_03_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in12 = reg_0483;
    6: op1_03_in12 = reg_0042;
    8: op1_03_in12 = reg_0042;
    7: op1_03_in12 = reg_0025;
    9: op1_03_in12 = reg_0284;
    10: op1_03_in12 = imem05_in[7:4];
    4: op1_03_in12 = reg_0180;
    11: op1_03_in12 = reg_0134;
    12: op1_03_in12 = reg_0983;
    13: op1_03_in12 = imem06_in[39:36];
    14: op1_03_in12 = reg_0636;
    15: op1_03_in12 = reg_0533;
    16: op1_03_in12 = reg_0628;
    17: op1_03_in12 = reg_0200;
    18: op1_03_in12 = imem05_in[91:88];
    19: op1_03_in12 = reg_0655;
    20: op1_03_in12 = reg_0552;
    21: op1_03_in12 = imem01_in[75:72];
    22: op1_03_in12 = reg_0062;
    23: op1_03_in12 = reg_0953;
    24: op1_03_in12 = imem03_in[123:120];
    25: op1_03_in12 = reg_0787;
    26: op1_03_in12 = reg_0472;
    27: op1_03_in12 = reg_0382;
    28: op1_03_in12 = reg_0471;
    29: op1_03_in12 = reg_0058;
    30: op1_03_in12 = reg_0139;
    31: op1_03_in12 = reg_0214;
    72: op1_03_in12 = reg_0214;
    32: op1_03_in12 = reg_0580;
    33: op1_03_in12 = reg_0969;
    34: op1_03_in12 = imem07_in[35:32];
    35: op1_03_in12 = reg_0517;
    36: op1_03_in12 = reg_0833;
    37: op1_03_in12 = imem05_in[75:72];
    38: op1_03_in12 = reg_0967;
    39: op1_03_in12 = reg_0943;
    41: op1_03_in12 = reg_0617;
    42: op1_03_in12 = reg_0110;
    43: op1_03_in12 = imem04_in[55:52];
    44: op1_03_in12 = reg_0407;
    45: op1_03_in12 = reg_0463;
    46: op1_03_in12 = reg_0762;
    47: op1_03_in12 = reg_0149;
    48: op1_03_in12 = reg_0388;
    49: op1_03_in12 = reg_0086;
    50: op1_03_in12 = reg_0108;
    51: op1_03_in12 = reg_0481;
    52: op1_03_in12 = imem07_in[51:48];
    54: op1_03_in12 = reg_0198;
    70: op1_03_in12 = reg_0198;
    55: op1_03_in12 = reg_1039;
    56: op1_03_in12 = reg_0642;
    57: op1_03_in12 = reg_0977;
    58: op1_03_in12 = reg_0994;
    59: op1_03_in12 = reg_0423;
    60: op1_03_in12 = reg_0144;
    61: op1_03_in12 = reg_0066;
    62: op1_03_in12 = reg_0140;
    63: op1_03_in12 = reg_0475;
    64: op1_03_in12 = imem01_in[27:24];
    65: op1_03_in12 = reg_0290;
    66: op1_03_in12 = reg_0894;
    67: op1_03_in12 = reg_0637;
    68: op1_03_in12 = imem03_in[127:124];
    69: op1_03_in12 = reg_0175;
    71: op1_03_in12 = reg_0051;
    73: op1_03_in12 = reg_0555;
    74: op1_03_in12 = reg_0818;
    75: op1_03_in12 = reg_0997;
    76: op1_03_in12 = reg_0624;
    77: op1_03_in12 = reg_0320;
    79: op1_03_in12 = imem02_in[99:96];
    80: op1_03_in12 = reg_0776;
    81: op1_03_in12 = reg_1005;
    82: op1_03_in12 = reg_0974;
    84: op1_03_in12 = reg_0660;
    85: op1_03_in12 = reg_0418;
    86: op1_03_in12 = reg_0067;
    87: op1_03_in12 = reg_0460;
    88: op1_03_in12 = reg_0213;
    89: op1_03_in12 = reg_0495;
    90: op1_03_in12 = reg_0087;
    91: op1_03_in12 = imem03_in[31:28];
    92: op1_03_in12 = imem03_in[83:80];
    93: op1_03_in12 = reg_0814;
    94: op1_03_in12 = reg_0895;
    95: op1_03_in12 = reg_0393;
    96: op1_03_in12 = reg_0338;
    97: op1_03_in12 = reg_0031;
    default: op1_03_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv12 = 1;
    7: op1_03_inv12 = 1;
    8: op1_03_inv12 = 1;
    9: op1_03_inv12 = 1;
    10: op1_03_inv12 = 1;
    4: op1_03_inv12 = 1;
    13: op1_03_inv12 = 1;
    18: op1_03_inv12 = 1;
    20: op1_03_inv12 = 1;
    27: op1_03_inv12 = 1;
    30: op1_03_inv12 = 1;
    32: op1_03_inv12 = 1;
    33: op1_03_inv12 = 1;
    34: op1_03_inv12 = 1;
    35: op1_03_inv12 = 1;
    37: op1_03_inv12 = 1;
    39: op1_03_inv12 = 1;
    41: op1_03_inv12 = 1;
    46: op1_03_inv12 = 1;
    47: op1_03_inv12 = 1;
    48: op1_03_inv12 = 1;
    49: op1_03_inv12 = 1;
    51: op1_03_inv12 = 1;
    52: op1_03_inv12 = 1;
    54: op1_03_inv12 = 1;
    55: op1_03_inv12 = 1;
    56: op1_03_inv12 = 1;
    58: op1_03_inv12 = 1;
    59: op1_03_inv12 = 1;
    60: op1_03_inv12 = 1;
    62: op1_03_inv12 = 1;
    63: op1_03_inv12 = 1;
    67: op1_03_inv12 = 1;
    68: op1_03_inv12 = 1;
    69: op1_03_inv12 = 1;
    74: op1_03_inv12 = 1;
    75: op1_03_inv12 = 1;
    77: op1_03_inv12 = 1;
    81: op1_03_inv12 = 1;
    82: op1_03_inv12 = 1;
    84: op1_03_inv12 = 1;
    85: op1_03_inv12 = 1;
    86: op1_03_inv12 = 1;
    87: op1_03_inv12 = 1;
    89: op1_03_inv12 = 1;
    91: op1_03_inv12 = 1;
    92: op1_03_inv12 = 1;
    93: op1_03_inv12 = 1;
    95: op1_03_inv12 = 1;
    default: op1_03_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in13 = reg_0484;
    6: op1_03_in13 = reg_0088;
    46: op1_03_in13 = reg_0088;
    7: op1_03_in13 = reg_0030;
    8: op1_03_in13 = reg_0089;
    9: op1_03_in13 = reg_0074;
    10: op1_03_in13 = imem05_in[27:24];
    4: op1_03_in13 = reg_0169;
    11: op1_03_in13 = reg_0144;
    12: op1_03_in13 = imem04_in[27:24];
    13: op1_03_in13 = imem06_in[79:76];
    14: op1_03_in13 = reg_0667;
    15: op1_03_in13 = reg_0541;
    16: op1_03_in13 = reg_0610;
    17: op1_03_in13 = reg_0194;
    18: op1_03_in13 = imem05_in[95:92];
    19: op1_03_in13 = reg_0661;
    20: op1_03_in13 = reg_0539;
    21: op1_03_in13 = imem01_in[79:76];
    22: op1_03_in13 = reg_0071;
    23: op1_03_in13 = reg_0136;
    24: op1_03_in13 = reg_0598;
    25: op1_03_in13 = reg_0027;
    26: op1_03_in13 = reg_0213;
    27: op1_03_in13 = reg_0383;
    28: op1_03_in13 = reg_0209;
    29: op1_03_in13 = reg_0517;
    30: op1_03_in13 = reg_0137;
    31: op1_03_in13 = reg_0210;
    32: op1_03_in13 = reg_0847;
    33: op1_03_in13 = reg_0942;
    34: op1_03_in13 = imem07_in[47:44];
    35: op1_03_in13 = reg_0854;
    36: op1_03_in13 = reg_0373;
    37: op1_03_in13 = reg_0970;
    38: op1_03_in13 = reg_0950;
    39: op1_03_in13 = reg_0826;
    41: op1_03_in13 = reg_0017;
    42: op1_03_in13 = imem02_in[19:16];
    43: op1_03_in13 = imem04_in[59:56];
    44: op1_03_in13 = reg_0556;
    45: op1_03_in13 = reg_0451;
    47: op1_03_in13 = reg_0151;
    48: op1_03_in13 = reg_0000;
    49: op1_03_in13 = reg_0090;
    50: op1_03_in13 = reg_0106;
    51: op1_03_in13 = reg_0470;
    52: op1_03_in13 = imem07_in[63:60];
    54: op1_03_in13 = reg_0201;
    70: op1_03_in13 = reg_0201;
    55: op1_03_in13 = reg_0869;
    56: op1_03_in13 = reg_0650;
    57: op1_03_in13 = reg_0988;
    58: op1_03_in13 = imem04_in[11:8];
    59: op1_03_in13 = reg_0007;
    60: op1_03_in13 = imem06_in[31:28];
    61: op1_03_in13 = reg_0276;
    62: op1_03_in13 = reg_0155;
    63: op1_03_in13 = reg_0460;
    64: op1_03_in13 = imem01_in[35:32];
    65: op1_03_in13 = reg_0225;
    66: op1_03_in13 = reg_0233;
    67: op1_03_in13 = reg_0341;
    68: op1_03_in13 = reg_0445;
    69: op1_03_in13 = reg_0162;
    71: op1_03_in13 = reg_0551;
    72: op1_03_in13 = reg_0208;
    73: op1_03_in13 = reg_0113;
    74: op1_03_in13 = reg_0772;
    75: op1_03_in13 = imem04_in[3:0];
    76: op1_03_in13 = reg_0008;
    77: op1_03_in13 = reg_0573;
    79: op1_03_in13 = reg_0813;
    80: op1_03_in13 = reg_0867;
    81: op1_03_in13 = reg_0778;
    82: op1_03_in13 = reg_0981;
    84: op1_03_in13 = reg_0080;
    85: op1_03_in13 = reg_0425;
    86: op1_03_in13 = reg_0302;
    87: op1_03_in13 = reg_0471;
    88: op1_03_in13 = reg_0190;
    89: op1_03_in13 = reg_0627;
    90: op1_03_in13 = reg_0037;
    91: op1_03_in13 = imem03_in[47:44];
    92: op1_03_in13 = imem03_in[87:84];
    93: op1_03_in13 = reg_1028;
    94: op1_03_in13 = reg_0606;
    95: op1_03_in13 = reg_0754;
    96: op1_03_in13 = reg_0614;
    97: op1_03_in13 = reg_0586;
    default: op1_03_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv13 = 1;
    7: op1_03_inv13 = 1;
    4: op1_03_inv13 = 1;
    14: op1_03_inv13 = 1;
    15: op1_03_inv13 = 1;
    16: op1_03_inv13 = 1;
    17: op1_03_inv13 = 1;
    18: op1_03_inv13 = 1;
    19: op1_03_inv13 = 1;
    20: op1_03_inv13 = 1;
    22: op1_03_inv13 = 1;
    25: op1_03_inv13 = 1;
    26: op1_03_inv13 = 1;
    27: op1_03_inv13 = 1;
    30: op1_03_inv13 = 1;
    33: op1_03_inv13 = 1;
    34: op1_03_inv13 = 1;
    36: op1_03_inv13 = 1;
    42: op1_03_inv13 = 1;
    43: op1_03_inv13 = 1;
    44: op1_03_inv13 = 1;
    46: op1_03_inv13 = 1;
    52: op1_03_inv13 = 1;
    54: op1_03_inv13 = 1;
    57: op1_03_inv13 = 1;
    58: op1_03_inv13 = 1;
    59: op1_03_inv13 = 1;
    62: op1_03_inv13 = 1;
    63: op1_03_inv13 = 1;
    64: op1_03_inv13 = 1;
    68: op1_03_inv13 = 1;
    70: op1_03_inv13 = 1;
    71: op1_03_inv13 = 1;
    75: op1_03_inv13 = 1;
    76: op1_03_inv13 = 1;
    77: op1_03_inv13 = 1;
    82: op1_03_inv13 = 1;
    85: op1_03_inv13 = 1;
    86: op1_03_inv13 = 1;
    89: op1_03_inv13 = 1;
    90: op1_03_inv13 = 1;
    91: op1_03_inv13 = 1;
    92: op1_03_inv13 = 1;
    96: op1_03_inv13 = 1;
    default: op1_03_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in14 = reg_0485;
    6: op1_03_in14 = reg_0084;
    7: op1_03_in14 = imem07_in[11:8];
    8: op1_03_in14 = reg_0097;
    9: op1_03_in14 = reg_0072;
    10: op1_03_in14 = imem05_in[51:48];
    4: op1_03_in14 = reg_0164;
    11: op1_03_in14 = imem06_in[19:16];
    12: op1_03_in14 = imem04_in[51:48];
    13: op1_03_in14 = imem06_in[111:108];
    14: op1_03_in14 = reg_0352;
    15: op1_03_in14 = reg_0547;
    16: op1_03_in14 = reg_0608;
    17: op1_03_in14 = imem01_in[3:0];
    18: op1_03_in14 = imem05_in[103:100];
    19: op1_03_in14 = reg_0648;
    20: op1_03_in14 = reg_0551;
    21: op1_03_in14 = imem01_in[107:104];
    22: op1_03_in14 = reg_0063;
    23: op1_03_in14 = reg_0154;
    24: op1_03_in14 = reg_0569;
    25: op1_03_in14 = reg_0781;
    26: op1_03_in14 = reg_0196;
    27: op1_03_in14 = reg_0403;
    28: op1_03_in14 = reg_0211;
    29: op1_03_in14 = reg_0875;
    30: op1_03_in14 = imem06_in[7:4];
    31: op1_03_in14 = reg_0190;
    32: op1_03_in14 = reg_0874;
    33: op1_03_in14 = reg_0961;
    34: op1_03_in14 = reg_0720;
    35: op1_03_in14 = reg_0855;
    36: op1_03_in14 = reg_0509;
    37: op1_03_in14 = reg_0948;
    38: op1_03_in14 = reg_0949;
    39: op1_03_in14 = reg_0244;
    41: op1_03_in14 = reg_0596;
    42: op1_03_in14 = imem02_in[71:68];
    43: op1_03_in14 = imem04_in[63:60];
    44: op1_03_in14 = reg_0783;
    45: op1_03_in14 = reg_0473;
    46: op1_03_in14 = reg_0089;
    59: op1_03_in14 = reg_0089;
    47: op1_03_in14 = reg_0153;
    48: op1_03_in14 = reg_1029;
    49: op1_03_in14 = reg_0091;
    50: op1_03_in14 = reg_0115;
    51: op1_03_in14 = reg_0478;
    52: op1_03_in14 = imem07_in[75:72];
    54: op1_03_in14 = reg_0195;
    70: op1_03_in14 = reg_0195;
    55: op1_03_in14 = reg_0604;
    56: op1_03_in14 = reg_0657;
    57: op1_03_in14 = imem04_in[71:68];
    58: op1_03_in14 = imem04_in[31:28];
    60: op1_03_in14 = imem06_in[75:72];
    61: op1_03_in14 = reg_0732;
    62: op1_03_in14 = imem06_in[11:8];
    63: op1_03_in14 = reg_0462;
    64: op1_03_in14 = imem01_in[71:68];
    65: op1_03_in14 = reg_0873;
    66: op1_03_in14 = reg_0039;
    67: op1_03_in14 = reg_0225;
    68: op1_03_in14 = reg_0577;
    69: op1_03_in14 = reg_0169;
    71: op1_03_in14 = reg_0995;
    72: op1_03_in14 = reg_0193;
    73: op1_03_in14 = reg_0821;
    74: op1_03_in14 = reg_0482;
    75: op1_03_in14 = imem04_in[19:16];
    76: op1_03_in14 = reg_0632;
    77: op1_03_in14 = reg_0566;
    79: op1_03_in14 = reg_0763;
    80: op1_03_in14 = reg_0079;
    81: op1_03_in14 = reg_0537;
    97: op1_03_in14 = reg_0537;
    82: op1_03_in14 = reg_0975;
    84: op1_03_in14 = reg_0625;
    85: op1_03_in14 = reg_0087;
    86: op1_03_in14 = reg_0584;
    87: op1_03_in14 = reg_0214;
    88: op1_03_in14 = reg_0197;
    89: op1_03_in14 = reg_0824;
    90: op1_03_in14 = reg_0083;
    91: op1_03_in14 = imem03_in[71:68];
    92: op1_03_in14 = reg_0631;
    93: op1_03_in14 = reg_0382;
    94: op1_03_in14 = reg_0822;
    95: op1_03_in14 = reg_1028;
    96: op1_03_in14 = reg_0510;
    default: op1_03_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv14 = 1;
    7: op1_03_inv14 = 1;
    8: op1_03_inv14 = 1;
    9: op1_03_inv14 = 1;
    4: op1_03_inv14 = 1;
    13: op1_03_inv14 = 1;
    14: op1_03_inv14 = 1;
    15: op1_03_inv14 = 1;
    16: op1_03_inv14 = 1;
    17: op1_03_inv14 = 1;
    18: op1_03_inv14 = 1;
    21: op1_03_inv14 = 1;
    23: op1_03_inv14 = 1;
    27: op1_03_inv14 = 1;
    29: op1_03_inv14 = 1;
    31: op1_03_inv14 = 1;
    32: op1_03_inv14 = 1;
    35: op1_03_inv14 = 1;
    36: op1_03_inv14 = 1;
    38: op1_03_inv14 = 1;
    39: op1_03_inv14 = 1;
    42: op1_03_inv14 = 1;
    44: op1_03_inv14 = 1;
    47: op1_03_inv14 = 1;
    48: op1_03_inv14 = 1;
    50: op1_03_inv14 = 1;
    51: op1_03_inv14 = 1;
    52: op1_03_inv14 = 1;
    59: op1_03_inv14 = 1;
    64: op1_03_inv14 = 1;
    65: op1_03_inv14 = 1;
    67: op1_03_inv14 = 1;
    68: op1_03_inv14 = 1;
    70: op1_03_inv14 = 1;
    72: op1_03_inv14 = 1;
    75: op1_03_inv14 = 1;
    79: op1_03_inv14 = 1;
    80: op1_03_inv14 = 1;
    82: op1_03_inv14 = 1;
    86: op1_03_inv14 = 1;
    92: op1_03_inv14 = 1;
    96: op1_03_inv14 = 1;
    default: op1_03_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in15 = reg_0486;
    6: op1_03_in15 = reg_0093;
    7: op1_03_in15 = imem07_in[23:20];
    77: op1_03_in15 = imem07_in[23:20];
    8: op1_03_in15 = reg_0073;
    9: op1_03_in15 = imem05_in[19:16];
    10: op1_03_in15 = imem05_in[55:52];
    11: op1_03_in15 = imem06_in[43:40];
    12: op1_03_in15 = imem04_in[107:104];
    13: op1_03_in15 = reg_0606;
    14: op1_03_in15 = reg_0334;
    15: op1_03_in15 = reg_0281;
    16: op1_03_in15 = reg_0618;
    17: op1_03_in15 = imem01_in[11:8];
    18: op1_03_in15 = imem05_in[107:104];
    19: op1_03_in15 = reg_0638;
    20: op1_03_in15 = reg_0733;
    21: op1_03_in15 = reg_0013;
    22: op1_03_in15 = reg_0296;
    23: op1_03_in15 = reg_0139;
    24: op1_03_in15 = reg_0592;
    25: op1_03_in15 = reg_1010;
    26: op1_03_in15 = imem01_in[31:28];
    27: op1_03_in15 = reg_0390;
    28: op1_03_in15 = reg_0194;
    29: op1_03_in15 = reg_0856;
    30: op1_03_in15 = imem06_in[11:8];
    31: op1_03_in15 = reg_0199;
    32: op1_03_in15 = reg_0038;
    33: op1_03_in15 = reg_0835;
    34: op1_03_in15 = reg_0708;
    35: op1_03_in15 = reg_0773;
    36: op1_03_in15 = reg_0820;
    37: op1_03_in15 = reg_0942;
    38: op1_03_in15 = reg_0946;
    39: op1_03_in15 = reg_0831;
    41: op1_03_in15 = reg_0025;
    48: op1_03_in15 = reg_0025;
    42: op1_03_in15 = reg_0657;
    43: op1_03_in15 = imem04_in[95:92];
    44: op1_03_in15 = reg_0754;
    45: op1_03_in15 = reg_0471;
    46: op1_03_in15 = reg_0867;
    47: op1_03_in15 = imem06_in[7:4];
    49: op1_03_in15 = imem03_in[15:12];
    50: op1_03_in15 = reg_0107;
    51: op1_03_in15 = reg_0214;
    52: op1_03_in15 = imem07_in[83:80];
    54: op1_03_in15 = reg_0192;
    55: op1_03_in15 = reg_0616;
    56: op1_03_in15 = reg_0326;
    57: op1_03_in15 = imem04_in[119:116];
    58: op1_03_in15 = imem04_in[43:40];
    59: op1_03_in15 = reg_0840;
    60: op1_03_in15 = imem06_in[83:80];
    61: op1_03_in15 = reg_0495;
    62: op1_03_in15 = imem06_in[15:12];
    63: op1_03_in15 = reg_0456;
    64: op1_03_in15 = imem01_in[107:104];
    65: op1_03_in15 = reg_0052;
    66: op1_03_in15 = reg_0389;
    67: op1_03_in15 = reg_0873;
    68: op1_03_in15 = reg_0590;
    69: op1_03_in15 = reg_0182;
    70: op1_03_in15 = imem01_in[63:60];
    71: op1_03_in15 = reg_0977;
    72: op1_03_in15 = reg_0198;
    73: op1_03_in15 = imem02_in[19:16];
    74: op1_03_in15 = reg_0085;
    75: op1_03_in15 = imem04_in[59:56];
    76: op1_03_in15 = reg_0026;
    79: op1_03_in15 = reg_0765;
    80: op1_03_in15 = imem03_in[11:8];
    81: op1_03_in15 = reg_0802;
    82: op1_03_in15 = reg_0988;
    84: op1_03_in15 = reg_1019;
    85: op1_03_in15 = imem02_in[35:32];
    86: op1_03_in15 = reg_0732;
    87: op1_03_in15 = reg_0200;
    88: op1_03_in15 = imem01_in[75:72];
    89: op1_03_in15 = imem05_in[3:0];
    90: op1_03_in15 = reg_0734;
    91: op1_03_in15 = imem03_in[87:84];
    92: op1_03_in15 = reg_0785;
    93: op1_03_in15 = reg_0029;
    94: op1_03_in15 = reg_0121;
    95: op1_03_in15 = reg_0822;
    96: op1_03_in15 = reg_0781;
    97: op1_03_in15 = reg_0568;
    default: op1_03_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_03_inv15 = 1;
    11: op1_03_inv15 = 1;
    13: op1_03_inv15 = 1;
    14: op1_03_inv15 = 1;
    18: op1_03_inv15 = 1;
    19: op1_03_inv15 = 1;
    21: op1_03_inv15 = 1;
    23: op1_03_inv15 = 1;
    24: op1_03_inv15 = 1;
    25: op1_03_inv15 = 1;
    27: op1_03_inv15 = 1;
    28: op1_03_inv15 = 1;
    29: op1_03_inv15 = 1;
    30: op1_03_inv15 = 1;
    31: op1_03_inv15 = 1;
    35: op1_03_inv15 = 1;
    37: op1_03_inv15 = 1;
    38: op1_03_inv15 = 1;
    41: op1_03_inv15 = 1;
    43: op1_03_inv15 = 1;
    44: op1_03_inv15 = 1;
    47: op1_03_inv15 = 1;
    48: op1_03_inv15 = 1;
    55: op1_03_inv15 = 1;
    56: op1_03_inv15 = 1;
    58: op1_03_inv15 = 1;
    64: op1_03_inv15 = 1;
    65: op1_03_inv15 = 1;
    66: op1_03_inv15 = 1;
    68: op1_03_inv15 = 1;
    71: op1_03_inv15 = 1;
    72: op1_03_inv15 = 1;
    73: op1_03_inv15 = 1;
    74: op1_03_inv15 = 1;
    75: op1_03_inv15 = 1;
    76: op1_03_inv15 = 1;
    77: op1_03_inv15 = 1;
    79: op1_03_inv15 = 1;
    80: op1_03_inv15 = 1;
    85: op1_03_inv15 = 1;
    89: op1_03_inv15 = 1;
    93: op1_03_inv15 = 1;
    97: op1_03_inv15 = 1;
    default: op1_03_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in16 = reg_0259;
    6: op1_03_in16 = reg_0825;
    7: op1_03_in16 = imem07_in[47:44];
    8: op1_03_in16 = imem03_in[115:112];
    9: op1_03_in16 = imem05_in[63:60];
    10: op1_03_in16 = imem05_in[63:60];
    11: op1_03_in16 = imem06_in[87:84];
    12: op1_03_in16 = reg_0545;
    13: op1_03_in16 = reg_0619;
    14: op1_03_in16 = reg_0341;
    15: op1_03_in16 = reg_0285;
    16: op1_03_in16 = reg_0622;
    17: op1_03_in16 = imem01_in[47:44];
    54: op1_03_in16 = imem01_in[47:44];
    18: op1_03_in16 = imem05_in[111:108];
    19: op1_03_in16 = reg_0644;
    42: op1_03_in16 = reg_0644;
    20: op1_03_in16 = reg_0072;
    21: op1_03_in16 = reg_0235;
    22: op1_03_in16 = reg_0525;
    23: op1_03_in16 = reg_0138;
    24: op1_03_in16 = reg_0585;
    25: op1_03_in16 = reg_0805;
    26: op1_03_in16 = imem01_in[63:60];
    27: op1_03_in16 = reg_0380;
    94: op1_03_in16 = reg_0380;
    95: op1_03_in16 = reg_0380;
    28: op1_03_in16 = reg_0206;
    29: op1_03_in16 = imem05_in[39:36];
    30: op1_03_in16 = imem06_in[35:32];
    31: op1_03_in16 = imem01_in[7:4];
    32: op1_03_in16 = reg_0051;
    33: op1_03_in16 = reg_0900;
    34: op1_03_in16 = reg_0709;
    35: op1_03_in16 = imem05_in[15:12];
    36: op1_03_in16 = reg_0513;
    37: op1_03_in16 = reg_0953;
    38: op1_03_in16 = reg_0952;
    39: op1_03_in16 = reg_0145;
    41: op1_03_in16 = imem07_in[23:20];
    43: op1_03_in16 = reg_0536;
    44: op1_03_in16 = reg_0495;
    45: op1_03_in16 = reg_0479;
    46: op1_03_in16 = reg_0506;
    47: op1_03_in16 = reg_0614;
    48: op1_03_in16 = imem07_in[11:8];
    76: op1_03_in16 = imem07_in[11:8];
    49: op1_03_in16 = imem03_in[39:36];
    50: op1_03_in16 = reg_0126;
    51: op1_03_in16 = reg_0209;
    87: op1_03_in16 = reg_0209;
    52: op1_03_in16 = imem07_in[91:88];
    55: op1_03_in16 = reg_0354;
    56: op1_03_in16 = reg_0637;
    57: op1_03_in16 = imem04_in[127:124];
    58: op1_03_in16 = imem04_in[83:80];
    59: op1_03_in16 = imem03_in[3:0];
    60: op1_03_in16 = reg_0344;
    61: op1_03_in16 = reg_0777;
    62: op1_03_in16 = imem06_in[71:68];
    63: op1_03_in16 = reg_0210;
    64: op1_03_in16 = reg_0786;
    65: op1_03_in16 = reg_0372;
    66: op1_03_in16 = reg_0372;
    67: op1_03_in16 = reg_0647;
    68: op1_03_in16 = reg_0833;
    69: op1_03_in16 = reg_0185;
    70: op1_03_in16 = imem01_in[83:80];
    71: op1_03_in16 = reg_0990;
    72: op1_03_in16 = imem01_in[51:48];
    73: op1_03_in16 = imem02_in[55:52];
    74: op1_03_in16 = reg_0090;
    75: op1_03_in16 = imem04_in[99:96];
    77: op1_03_in16 = imem07_in[95:92];
    79: op1_03_in16 = reg_0358;
    80: op1_03_in16 = imem03_in[35:32];
    81: op1_03_in16 = reg_0752;
    82: op1_03_in16 = imem04_in[35:32];
    84: op1_03_in16 = reg_0267;
    85: op1_03_in16 = imem02_in[51:48];
    86: op1_03_in16 = reg_0552;
    88: op1_03_in16 = imem01_in[79:76];
    89: op1_03_in16 = imem05_in[79:76];
    90: op1_03_in16 = reg_0155;
    91: op1_03_in16 = imem03_in[91:88];
    92: op1_03_in16 = reg_0743;
    93: op1_03_in16 = reg_0918;
    96: op1_03_in16 = reg_1020;
    97: op1_03_in16 = reg_0584;
    default: op1_03_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv16 = 1;
    6: op1_03_inv16 = 1;
    11: op1_03_inv16 = 1;
    12: op1_03_inv16 = 1;
    15: op1_03_inv16 = 1;
    20: op1_03_inv16 = 1;
    23: op1_03_inv16 = 1;
    24: op1_03_inv16 = 1;
    25: op1_03_inv16 = 1;
    27: op1_03_inv16 = 1;
    29: op1_03_inv16 = 1;
    32: op1_03_inv16 = 1;
    33: op1_03_inv16 = 1;
    35: op1_03_inv16 = 1;
    39: op1_03_inv16 = 1;
    41: op1_03_inv16 = 1;
    43: op1_03_inv16 = 1;
    44: op1_03_inv16 = 1;
    45: op1_03_inv16 = 1;
    48: op1_03_inv16 = 1;
    49: op1_03_inv16 = 1;
    54: op1_03_inv16 = 1;
    55: op1_03_inv16 = 1;
    56: op1_03_inv16 = 1;
    58: op1_03_inv16 = 1;
    61: op1_03_inv16 = 1;
    65: op1_03_inv16 = 1;
    67: op1_03_inv16 = 1;
    68: op1_03_inv16 = 1;
    69: op1_03_inv16 = 1;
    76: op1_03_inv16 = 1;
    77: op1_03_inv16 = 1;
    81: op1_03_inv16 = 1;
    86: op1_03_inv16 = 1;
    87: op1_03_inv16 = 1;
    88: op1_03_inv16 = 1;
    89: op1_03_inv16 = 1;
    92: op1_03_inv16 = 1;
    96: op1_03_inv16 = 1;
    97: op1_03_inv16 = 1;
    default: op1_03_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in17 = reg_0260;
    6: op1_03_in17 = reg_0568;
    7: op1_03_in17 = imem07_in[51:48];
    8: op1_03_in17 = reg_0573;
    9: op1_03_in17 = imem05_in[67:64];
    10: op1_03_in17 = imem05_in[75:72];
    11: op1_03_in17 = imem06_in[103:100];
    12: op1_03_in17 = reg_0550;
    13: op1_03_in17 = reg_0615;
    14: op1_03_in17 = reg_0330;
    15: op1_03_in17 = reg_0286;
    16: op1_03_in17 = reg_0407;
    17: op1_03_in17 = imem01_in[51:48];
    18: op1_03_in17 = imem05_in[119:116];
    19: op1_03_in17 = reg_0643;
    20: op1_03_in17 = reg_0882;
    21: op1_03_in17 = reg_1049;
    22: op1_03_in17 = reg_0054;
    66: op1_03_in17 = reg_0054;
    23: op1_03_in17 = reg_0153;
    39: op1_03_in17 = reg_0153;
    24: op1_03_in17 = reg_0600;
    25: op1_03_in17 = reg_1011;
    26: op1_03_in17 = imem01_in[95:92];
    88: op1_03_in17 = imem01_in[95:92];
    27: op1_03_in17 = reg_0799;
    28: op1_03_in17 = reg_0197;
    29: op1_03_in17 = imem05_in[63:60];
    30: op1_03_in17 = imem06_in[95:92];
    31: op1_03_in17 = imem01_in[39:36];
    32: op1_03_in17 = reg_0376;
    33: op1_03_in17 = reg_0757;
    34: op1_03_in17 = reg_0718;
    35: op1_03_in17 = imem05_in[59:56];
    36: op1_03_in17 = reg_0979;
    37: op1_03_in17 = reg_0972;
    38: op1_03_in17 = reg_0953;
    41: op1_03_in17 = imem07_in[27:24];
    42: op1_03_in17 = reg_0652;
    43: op1_03_in17 = reg_1003;
    44: op1_03_in17 = reg_0309;
    45: op1_03_in17 = reg_0456;
    46: op1_03_in17 = reg_0884;
    47: op1_03_in17 = reg_0895;
    48: op1_03_in17 = imem07_in[59:56];
    49: op1_03_in17 = imem03_in[47:44];
    50: op1_03_in17 = imem02_in[51:48];
    51: op1_03_in17 = reg_0207;
    52: op1_03_in17 = imem07_in[95:92];
    54: op1_03_in17 = imem01_in[79:76];
    55: op1_03_in17 = reg_1041;
    56: op1_03_in17 = reg_0565;
    57: op1_03_in17 = reg_1004;
    58: op1_03_in17 = reg_1009;
    59: op1_03_in17 = imem03_in[19:16];
    60: op1_03_in17 = reg_0696;
    61: op1_03_in17 = reg_0332;
    62: op1_03_in17 = imem06_in[91:88];
    63: op1_03_in17 = reg_0189;
    64: op1_03_in17 = reg_0592;
    65: op1_03_in17 = reg_0083;
    67: op1_03_in17 = reg_0036;
    68: op1_03_in17 = reg_0992;
    70: op1_03_in17 = imem01_in[87:84];
    72: op1_03_in17 = imem01_in[87:84];
    71: op1_03_in17 = imem04_in[43:40];
    73: op1_03_in17 = imem02_in[59:56];
    74: op1_03_in17 = reg_0840;
    75: op1_03_in17 = reg_0539;
    76: op1_03_in17 = imem07_in[19:16];
    77: op1_03_in17 = imem07_in[123:120];
    79: op1_03_in17 = reg_0081;
    80: op1_03_in17 = imem03_in[83:80];
    81: op1_03_in17 = reg_0056;
    82: op1_03_in17 = imem04_in[51:48];
    84: op1_03_in17 = reg_0021;
    85: op1_03_in17 = imem02_in[75:72];
    86: op1_03_in17 = reg_0409;
    87: op1_03_in17 = reg_0193;
    89: op1_03_in17 = imem05_in[115:112];
    90: op1_03_in17 = reg_0085;
    91: op1_03_in17 = imem03_in[103:100];
    92: op1_03_in17 = reg_0623;
    93: op1_03_in17 = reg_1029;
    94: op1_03_in17 = reg_0804;
    95: op1_03_in17 = reg_0811;
    96: op1_03_in17 = reg_0914;
    97: op1_03_in17 = reg_0296;
    default: op1_03_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv17 = 1;
    7: op1_03_inv17 = 1;
    8: op1_03_inv17 = 1;
    9: op1_03_inv17 = 1;
    11: op1_03_inv17 = 1;
    12: op1_03_inv17 = 1;
    13: op1_03_inv17 = 1;
    14: op1_03_inv17 = 1;
    16: op1_03_inv17 = 1;
    17: op1_03_inv17 = 1;
    19: op1_03_inv17 = 1;
    24: op1_03_inv17 = 1;
    25: op1_03_inv17 = 1;
    26: op1_03_inv17 = 1;
    27: op1_03_inv17 = 1;
    29: op1_03_inv17 = 1;
    30: op1_03_inv17 = 1;
    32: op1_03_inv17 = 1;
    33: op1_03_inv17 = 1;
    36: op1_03_inv17 = 1;
    37: op1_03_inv17 = 1;
    38: op1_03_inv17 = 1;
    41: op1_03_inv17 = 1;
    42: op1_03_inv17 = 1;
    47: op1_03_inv17 = 1;
    51: op1_03_inv17 = 1;
    52: op1_03_inv17 = 1;
    54: op1_03_inv17 = 1;
    55: op1_03_inv17 = 1;
    56: op1_03_inv17 = 1;
    58: op1_03_inv17 = 1;
    59: op1_03_inv17 = 1;
    60: op1_03_inv17 = 1;
    63: op1_03_inv17 = 1;
    70: op1_03_inv17 = 1;
    72: op1_03_inv17 = 1;
    73: op1_03_inv17 = 1;
    74: op1_03_inv17 = 1;
    76: op1_03_inv17 = 1;
    77: op1_03_inv17 = 1;
    80: op1_03_inv17 = 1;
    81: op1_03_inv17 = 1;
    85: op1_03_inv17 = 1;
    87: op1_03_inv17 = 1;
    88: op1_03_inv17 = 1;
    89: op1_03_inv17 = 1;
    90: op1_03_inv17 = 1;
    92: op1_03_inv17 = 1;
    93: op1_03_inv17 = 1;
    94: op1_03_inv17 = 1;
    95: op1_03_inv17 = 1;
    default: op1_03_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in18 = reg_0132;
    6: op1_03_in18 = reg_0589;
    7: op1_03_in18 = imem07_in[67:64];
    8: op1_03_in18 = reg_0579;
    9: op1_03_in18 = imem05_in[75:72];
    35: op1_03_in18 = imem05_in[75:72];
    10: op1_03_in18 = imem05_in[83:80];
    11: op1_03_in18 = reg_0614;
    12: op1_03_in18 = reg_0529;
    13: op1_03_in18 = reg_0379;
    14: op1_03_in18 = reg_0324;
    15: op1_03_in18 = reg_0307;
    16: op1_03_in18 = reg_0371;
    17: op1_03_in18 = imem01_in[67:64];
    18: op1_03_in18 = reg_0956;
    19: op1_03_in18 = reg_0652;
    20: op1_03_in18 = reg_0015;
    21: op1_03_in18 = reg_0248;
    22: op1_03_in18 = reg_0279;
    23: op1_03_in18 = reg_0144;
    24: op1_03_in18 = reg_0597;
    25: op1_03_in18 = imem07_in[23:20];
    76: op1_03_in18 = imem07_in[23:20];
    26: op1_03_in18 = imem01_in[103:100];
    27: op1_03_in18 = reg_1028;
    28: op1_03_in18 = imem01_in[15:12];
    29: op1_03_in18 = imem05_in[91:88];
    30: op1_03_in18 = reg_0628;
    31: op1_03_in18 = imem01_in[55:52];
    32: op1_03_in18 = reg_0312;
    33: op1_03_in18 = reg_0147;
    34: op1_03_in18 = reg_0422;
    36: op1_03_in18 = reg_0974;
    37: op1_03_in18 = reg_0821;
    38: op1_03_in18 = reg_0960;
    39: op1_03_in18 = reg_0140;
    41: op1_03_in18 = imem07_in[55:52];
    42: op1_03_in18 = reg_0334;
    43: op1_03_in18 = reg_0306;
    44: op1_03_in18 = reg_0241;
    45: op1_03_in18 = reg_0214;
    46: op1_03_in18 = imem03_in[3:0];
    47: op1_03_in18 = reg_0624;
    48: op1_03_in18 = imem07_in[87:84];
    49: op1_03_in18 = imem03_in[59:56];
    50: op1_03_in18 = imem02_in[67:64];
    51: op1_03_in18 = reg_0211;
    52: op1_03_in18 = imem07_in[111:108];
    54: op1_03_in18 = reg_0779;
    55: op1_03_in18 = reg_0512;
    56: op1_03_in18 = reg_0636;
    57: op1_03_in18 = reg_0536;
    58: op1_03_in18 = reg_1020;
    59: op1_03_in18 = imem03_in[43:40];
    60: op1_03_in18 = reg_0754;
    61: op1_03_in18 = imem05_in[7:4];
    62: op1_03_in18 = imem06_in[107:104];
    63: op1_03_in18 = reg_0201;
    64: op1_03_in18 = reg_0253;
    65: op1_03_in18 = reg_0007;
    66: op1_03_in18 = reg_0792;
    67: op1_03_in18 = reg_0565;
    68: op1_03_in18 = reg_0979;
    70: op1_03_in18 = reg_0337;
    71: op1_03_in18 = imem04_in[103:100];
    72: op1_03_in18 = imem01_in[95:92];
    73: op1_03_in18 = imem02_in[107:104];
    74: op1_03_in18 = imem03_in[67:64];
    75: op1_03_in18 = reg_1005;
    77: op1_03_in18 = imem07_in[127:124];
    79: op1_03_in18 = reg_0052;
    80: op1_03_in18 = imem03_in[99:96];
    81: op1_03_in18 = reg_0584;
    82: op1_03_in18 = imem04_in[83:80];
    84: op1_03_in18 = reg_0926;
    85: op1_03_in18 = imem02_in[111:108];
    86: op1_03_in18 = reg_0495;
    87: op1_03_in18 = reg_0192;
    88: op1_03_in18 = imem01_in[119:116];
    89: op1_03_in18 = reg_0866;
    90: op1_03_in18 = reg_0656;
    91: op1_03_in18 = reg_0342;
    92: op1_03_in18 = reg_0331;
    93: op1_03_in18 = reg_0289;
    94: op1_03_in18 = imem07_in[39:36];
    95: op1_03_in18 = reg_0914;
    96: op1_03_in18 = reg_0040;
    97: op1_03_in18 = reg_0072;
    default: op1_03_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv18 = 1;
    6: op1_03_inv18 = 1;
    7: op1_03_inv18 = 1;
    8: op1_03_inv18 = 1;
    11: op1_03_inv18 = 1;
    12: op1_03_inv18 = 1;
    14: op1_03_inv18 = 1;
    15: op1_03_inv18 = 1;
    18: op1_03_inv18 = 1;
    20: op1_03_inv18 = 1;
    21: op1_03_inv18 = 1;
    22: op1_03_inv18 = 1;
    24: op1_03_inv18 = 1;
    28: op1_03_inv18 = 1;
    29: op1_03_inv18 = 1;
    30: op1_03_inv18 = 1;
    31: op1_03_inv18 = 1;
    33: op1_03_inv18 = 1;
    34: op1_03_inv18 = 1;
    35: op1_03_inv18 = 1;
    36: op1_03_inv18 = 1;
    37: op1_03_inv18 = 1;
    39: op1_03_inv18 = 1;
    43: op1_03_inv18 = 1;
    47: op1_03_inv18 = 1;
    49: op1_03_inv18 = 1;
    54: op1_03_inv18 = 1;
    56: op1_03_inv18 = 1;
    57: op1_03_inv18 = 1;
    58: op1_03_inv18 = 1;
    59: op1_03_inv18 = 1;
    61: op1_03_inv18 = 1;
    65: op1_03_inv18 = 1;
    68: op1_03_inv18 = 1;
    70: op1_03_inv18 = 1;
    73: op1_03_inv18 = 1;
    74: op1_03_inv18 = 1;
    76: op1_03_inv18 = 1;
    79: op1_03_inv18 = 1;
    81: op1_03_inv18 = 1;
    82: op1_03_inv18 = 1;
    84: op1_03_inv18 = 1;
    85: op1_03_inv18 = 1;
    88: op1_03_inv18 = 1;
    90: op1_03_inv18 = 1;
    91: op1_03_inv18 = 1;
    92: op1_03_inv18 = 1;
    93: op1_03_inv18 = 1;
    94: op1_03_inv18 = 1;
    default: op1_03_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in19 = reg_0136;
    6: op1_03_in19 = reg_0580;
    7: op1_03_in19 = imem07_in[71:68];
    8: op1_03_in19 = reg_0597;
    9: op1_03_in19 = imem05_in[91:88];
    10: op1_03_in19 = imem05_in[119:116];
    11: op1_03_in19 = reg_0604;
    12: op1_03_in19 = reg_0556;
    13: op1_03_in19 = reg_0390;
    14: op1_03_in19 = reg_0365;
    15: op1_03_in19 = reg_0061;
    16: op1_03_in19 = reg_0382;
    17: op1_03_in19 = imem01_in[119:116];
    18: op1_03_in19 = reg_0942;
    19: op1_03_in19 = reg_0357;
    20: op1_03_in19 = reg_0525;
    21: op1_03_in19 = reg_0234;
    22: op1_03_in19 = reg_0854;
    86: op1_03_in19 = reg_0854;
    23: op1_03_in19 = imem06_in[15:12];
    24: op1_03_in19 = reg_0391;
    25: op1_03_in19 = imem07_in[31:28];
    26: op1_03_in19 = reg_0238;
    27: op1_03_in19 = reg_0798;
    28: op1_03_in19 = imem01_in[31:28];
    29: op1_03_in19 = reg_0954;
    30: op1_03_in19 = reg_0621;
    31: op1_03_in19 = imem01_in[87:84];
    32: op1_03_in19 = reg_0374;
    33: op1_03_in19 = reg_0139;
    34: op1_03_in19 = reg_0421;
    35: op1_03_in19 = imem05_in[99:96];
    36: op1_03_in19 = imem04_in[11:8];
    37: op1_03_in19 = reg_0826;
    38: op1_03_in19 = reg_0834;
    39: op1_03_in19 = reg_0155;
    41: op1_03_in19 = imem07_in[59:56];
    94: op1_03_in19 = imem07_in[59:56];
    42: op1_03_in19 = reg_0097;
    43: op1_03_in19 = reg_1057;
    44: op1_03_in19 = reg_1010;
    45: op1_03_in19 = reg_0189;
    46: op1_03_in19 = imem03_in[71:68];
    47: op1_03_in19 = reg_0220;
    48: op1_03_in19 = imem07_in[115:112];
    49: op1_03_in19 = imem03_in[127:124];
    50: op1_03_in19 = imem02_in[119:116];
    51: op1_03_in19 = reg_0192;
    52: op1_03_in19 = reg_0722;
    54: op1_03_in19 = reg_0904;
    55: op1_03_in19 = reg_0827;
    56: op1_03_in19 = reg_0279;
    57: op1_03_in19 = reg_0511;
    58: op1_03_in19 = reg_0909;
    59: op1_03_in19 = imem03_in[95:92];
    60: op1_03_in19 = reg_0692;
    61: op1_03_in19 = imem05_in[23:20];
    62: op1_03_in19 = reg_0694;
    63: op1_03_in19 = reg_0213;
    64: op1_03_in19 = reg_1034;
    65: op1_03_in19 = reg_0506;
    66: op1_03_in19 = reg_0090;
    67: op1_03_in19 = reg_0323;
    68: op1_03_in19 = reg_0993;
    70: op1_03_in19 = reg_0592;
    71: op1_03_in19 = imem04_in[111:108];
    72: op1_03_in19 = imem01_in[99:96];
    73: op1_03_in19 = reg_0700;
    74: op1_03_in19 = imem03_in[91:88];
    75: op1_03_in19 = reg_0067;
    76: op1_03_in19 = imem07_in[39:36];
    77: op1_03_in19 = reg_0919;
    79: op1_03_in19 = reg_0394;
    80: op1_03_in19 = imem03_in[111:108];
    81: op1_03_in19 = reg_0288;
    82: op1_03_in19 = imem04_in[103:100];
    84: op1_03_in19 = reg_0328;
    85: op1_03_in19 = imem03_in[7:4];
    87: op1_03_in19 = imem01_in[35:32];
    88: op1_03_in19 = imem01_in[127:124];
    89: op1_03_in19 = reg_0492;
    90: op1_03_in19 = reg_0788;
    91: op1_03_in19 = reg_0579;
    92: op1_03_in19 = reg_0571;
    93: op1_03_in19 = reg_0133;
    95: op1_03_in19 = reg_0392;
    96: op1_03_in19 = reg_0018;
    97: op1_03_in19 = reg_0658;
    default: op1_03_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_03_inv19 = 1;
    9: op1_03_inv19 = 1;
    14: op1_03_inv19 = 1;
    16: op1_03_inv19 = 1;
    18: op1_03_inv19 = 1;
    19: op1_03_inv19 = 1;
    20: op1_03_inv19 = 1;
    21: op1_03_inv19 = 1;
    24: op1_03_inv19 = 1;
    26: op1_03_inv19 = 1;
    31: op1_03_inv19 = 1;
    33: op1_03_inv19 = 1;
    35: op1_03_inv19 = 1;
    37: op1_03_inv19 = 1;
    41: op1_03_inv19 = 1;
    42: op1_03_inv19 = 1;
    44: op1_03_inv19 = 1;
    45: op1_03_inv19 = 1;
    46: op1_03_inv19 = 1;
    47: op1_03_inv19 = 1;
    51: op1_03_inv19 = 1;
    52: op1_03_inv19 = 1;
    55: op1_03_inv19 = 1;
    57: op1_03_inv19 = 1;
    60: op1_03_inv19 = 1;
    64: op1_03_inv19 = 1;
    65: op1_03_inv19 = 1;
    75: op1_03_inv19 = 1;
    81: op1_03_inv19 = 1;
    82: op1_03_inv19 = 1;
    84: op1_03_inv19 = 1;
    85: op1_03_inv19 = 1;
    89: op1_03_inv19 = 1;
    90: op1_03_inv19 = 1;
    91: op1_03_inv19 = 1;
    93: op1_03_inv19 = 1;
    95: op1_03_inv19 = 1;
    96: op1_03_inv19 = 1;
    97: op1_03_inv19 = 1;
    default: op1_03_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in20 = reg_0137;
    6: op1_03_in20 = reg_0590;
    8: op1_03_in20 = reg_0590;
    7: op1_03_in20 = imem07_in[79:76];
    9: op1_03_in20 = reg_0973;
    10: op1_03_in20 = reg_0973;
    11: op1_03_in20 = reg_0607;
    12: op1_03_in20 = reg_0308;
    13: op1_03_in20 = reg_0486;
    14: op1_03_in20 = reg_0336;
    42: op1_03_in20 = reg_0336;
    15: op1_03_in20 = reg_0062;
    16: op1_03_in20 = reg_0368;
    56: op1_03_in20 = reg_0368;
    17: op1_03_in20 = imem01_in[127:124];
    18: op1_03_in20 = reg_0946;
    19: op1_03_in20 = reg_0341;
    20: op1_03_in20 = reg_0047;
    21: op1_03_in20 = reg_0245;
    22: op1_03_in20 = reg_0286;
    23: op1_03_in20 = imem06_in[91:88];
    24: op1_03_in20 = reg_0360;
    25: op1_03_in20 = imem07_in[39:36];
    26: op1_03_in20 = reg_1033;
    27: op1_03_in20 = imem07_in[35:32];
    28: op1_03_in20 = imem01_in[39:36];
    87: op1_03_in20 = imem01_in[39:36];
    29: op1_03_in20 = reg_0957;
    30: op1_03_in20 = reg_0626;
    31: op1_03_in20 = imem01_in[111:108];
    32: op1_03_in20 = reg_0991;
    33: op1_03_in20 = reg_0131;
    34: op1_03_in20 = reg_0426;
    35: op1_03_in20 = imem05_in[119:116];
    36: op1_03_in20 = imem04_in[39:36];
    37: op1_03_in20 = reg_0835;
    38: op1_03_in20 = reg_0835;
    39: op1_03_in20 = imem06_in[79:76];
    41: op1_03_in20 = reg_0703;
    43: op1_03_in20 = reg_0888;
    44: op1_03_in20 = reg_0005;
    45: op1_03_in20 = reg_0203;
    46: op1_03_in20 = imem03_in[99:96];
    47: op1_03_in20 = reg_0782;
    48: op1_03_in20 = reg_0726;
    49: op1_03_in20 = reg_1049;
    91: op1_03_in20 = reg_1049;
    50: op1_03_in20 = reg_0650;
    51: op1_03_in20 = imem01_in[47:44];
    52: op1_03_in20 = reg_0731;
    54: op1_03_in20 = reg_0870;
    55: op1_03_in20 = reg_0115;
    57: op1_03_in20 = reg_0912;
    58: op1_03_in20 = reg_0066;
    59: op1_03_in20 = imem03_in[103:100];
    60: op1_03_in20 = reg_0440;
    61: op1_03_in20 = imem05_in[31:28];
    62: op1_03_in20 = reg_0294;
    63: op1_03_in20 = reg_0206;
    64: op1_03_in20 = reg_0798;
    65: op1_03_in20 = imem03_in[11:8];
    66: op1_03_in20 = reg_0049;
    67: op1_03_in20 = reg_0441;
    68: op1_03_in20 = reg_0999;
    70: op1_03_in20 = reg_0518;
    71: op1_03_in20 = reg_0483;
    72: op1_03_in20 = imem01_in[119:116];
    73: op1_03_in20 = reg_0886;
    74: op1_03_in20 = imem03_in[95:92];
    75: op1_03_in20 = reg_0815;
    76: op1_03_in20 = imem07_in[47:44];
    77: op1_03_in20 = reg_0713;
    79: op1_03_in20 = reg_0389;
    80: op1_03_in20 = imem03_in[119:116];
    81: op1_03_in20 = reg_0027;
    82: op1_03_in20 = imem04_in[119:116];
    84: op1_03_in20 = reg_0692;
    85: op1_03_in20 = imem03_in[19:16];
    86: op1_03_in20 = reg_0071;
    88: op1_03_in20 = reg_1032;
    89: op1_03_in20 = reg_0217;
    90: op1_03_in20 = reg_0984;
    92: op1_03_in20 = reg_0397;
    93: op1_03_in20 = reg_0914;
    94: op1_03_in20 = imem07_in[83:80];
    95: op1_03_in20 = reg_0036;
    96: op1_03_in20 = reg_0611;
    97: op1_03_in20 = reg_0065;
    default: op1_03_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv20 = 1;
    6: op1_03_inv20 = 1;
    7: op1_03_inv20 = 1;
    8: op1_03_inv20 = 1;
    10: op1_03_inv20 = 1;
    13: op1_03_inv20 = 1;
    14: op1_03_inv20 = 1;
    15: op1_03_inv20 = 1;
    17: op1_03_inv20 = 1;
    19: op1_03_inv20 = 1;
    21: op1_03_inv20 = 1;
    23: op1_03_inv20 = 1;
    24: op1_03_inv20 = 1;
    25: op1_03_inv20 = 1;
    26: op1_03_inv20 = 1;
    30: op1_03_inv20 = 1;
    36: op1_03_inv20 = 1;
    37: op1_03_inv20 = 1;
    41: op1_03_inv20 = 1;
    42: op1_03_inv20 = 1;
    43: op1_03_inv20 = 1;
    45: op1_03_inv20 = 1;
    47: op1_03_inv20 = 1;
    48: op1_03_inv20 = 1;
    51: op1_03_inv20 = 1;
    55: op1_03_inv20 = 1;
    56: op1_03_inv20 = 1;
    57: op1_03_inv20 = 1;
    58: op1_03_inv20 = 1;
    59: op1_03_inv20 = 1;
    63: op1_03_inv20 = 1;
    64: op1_03_inv20 = 1;
    65: op1_03_inv20 = 1;
    66: op1_03_inv20 = 1;
    71: op1_03_inv20 = 1;
    75: op1_03_inv20 = 1;
    80: op1_03_inv20 = 1;
    81: op1_03_inv20 = 1;
    85: op1_03_inv20 = 1;
    90: op1_03_inv20 = 1;
    92: op1_03_inv20 = 1;
    93: op1_03_inv20 = 1;
    96: op1_03_inv20 = 1;
    default: op1_03_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in21 = reg_0144;
    6: op1_03_in21 = reg_0387;
    7: op1_03_in21 = reg_0719;
    8: op1_03_in21 = reg_0360;
    9: op1_03_in21 = reg_0944;
    10: op1_03_in21 = reg_0970;
    11: op1_03_in21 = reg_0624;
    12: op1_03_in21 = reg_0301;
    13: op1_03_in21 = reg_0801;
    14: op1_03_in21 = reg_0081;
    15: op1_03_in21 = reg_0065;
    16: op1_03_in21 = reg_1029;
    17: op1_03_in21 = reg_1055;
    18: op1_03_in21 = reg_0960;
    19: op1_03_in21 = reg_0359;
    20: op1_03_in21 = reg_0286;
    21: op1_03_in21 = reg_1052;
    22: op1_03_in21 = imem05_in[3:0];
    23: op1_03_in21 = reg_0625;
    24: op1_03_in21 = reg_0369;
    25: op1_03_in21 = imem07_in[87:84];
    27: op1_03_in21 = imem07_in[87:84];
    94: op1_03_in21 = imem07_in[87:84];
    26: op1_03_in21 = reg_1041;
    28: op1_03_in21 = imem01_in[67:64];
    29: op1_03_in21 = reg_0965;
    30: op1_03_in21 = reg_0601;
    31: op1_03_in21 = reg_0779;
    91: op1_03_in21 = reg_0779;
    32: op1_03_in21 = reg_0979;
    33: op1_03_in21 = imem06_in[39:36];
    34: op1_03_in21 = reg_0434;
    35: op1_03_in21 = reg_0942;
    36: op1_03_in21 = imem04_in[51:48];
    37: op1_03_in21 = reg_0256;
    38: op1_03_in21 = reg_0229;
    39: op1_03_in21 = imem06_in[119:116];
    41: op1_03_in21 = reg_0712;
    42: op1_03_in21 = reg_0007;
    43: op1_03_in21 = reg_0313;
    44: op1_03_in21 = imem07_in[3:0];
    45: op1_03_in21 = reg_0186;
    46: op1_03_in21 = reg_0357;
    47: op1_03_in21 = reg_0632;
    48: op1_03_in21 = reg_0714;
    49: op1_03_in21 = reg_0765;
    73: op1_03_in21 = reg_0765;
    50: op1_03_in21 = reg_0654;
    51: op1_03_in21 = imem01_in[99:96];
    52: op1_03_in21 = reg_0726;
    54: op1_03_in21 = reg_1036;
    55: op1_03_in21 = reg_0113;
    56: op1_03_in21 = reg_0608;
    57: op1_03_in21 = reg_0292;
    58: op1_03_in21 = reg_0288;
    59: op1_03_in21 = imem03_in[107:104];
    74: op1_03_in21 = imem03_in[107:104];
    60: op1_03_in21 = reg_0297;
    61: op1_03_in21 = imem05_in[55:52];
    62: op1_03_in21 = reg_1011;
    63: op1_03_in21 = imem01_in[31:28];
    64: op1_03_in21 = reg_0869;
    65: op1_03_in21 = imem03_in[43:40];
    66: op1_03_in21 = reg_0291;
    67: op1_03_in21 = reg_0424;
    68: op1_03_in21 = imem04_in[23:20];
    70: op1_03_in21 = reg_0831;
    71: op1_03_in21 = reg_0539;
    72: op1_03_in21 = reg_1014;
    75: op1_03_in21 = reg_0494;
    76: op1_03_in21 = reg_0892;
    77: op1_03_in21 = reg_0515;
    79: op1_03_in21 = reg_0331;
    80: op1_03_in21 = reg_0099;
    81: op1_03_in21 = reg_0517;
    82: op1_03_in21 = imem04_in[127:124];
    84: op1_03_in21 = reg_0028;
    85: op1_03_in21 = imem03_in[39:36];
    86: op1_03_in21 = reg_0070;
    87: op1_03_in21 = imem01_in[51:48];
    88: op1_03_in21 = reg_0968;
    89: op1_03_in21 = reg_0954;
    90: op1_03_in21 = reg_0327;
    92: op1_03_in21 = reg_0579;
    93: op1_03_in21 = reg_0919;
    95: op1_03_in21 = reg_0611;
    96: op1_03_in21 = reg_0403;
    97: op1_03_in21 = reg_0332;
    default: op1_03_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv21 = 1;
    10: op1_03_inv21 = 1;
    13: op1_03_inv21 = 1;
    15: op1_03_inv21 = 1;
    19: op1_03_inv21 = 1;
    21: op1_03_inv21 = 1;
    22: op1_03_inv21 = 1;
    23: op1_03_inv21 = 1;
    24: op1_03_inv21 = 1;
    26: op1_03_inv21 = 1;
    30: op1_03_inv21 = 1;
    33: op1_03_inv21 = 1;
    37: op1_03_inv21 = 1;
    38: op1_03_inv21 = 1;
    41: op1_03_inv21 = 1;
    43: op1_03_inv21 = 1;
    44: op1_03_inv21 = 1;
    48: op1_03_inv21 = 1;
    49: op1_03_inv21 = 1;
    50: op1_03_inv21 = 1;
    51: op1_03_inv21 = 1;
    52: op1_03_inv21 = 1;
    56: op1_03_inv21 = 1;
    57: op1_03_inv21 = 1;
    59: op1_03_inv21 = 1;
    60: op1_03_inv21 = 1;
    61: op1_03_inv21 = 1;
    62: op1_03_inv21 = 1;
    64: op1_03_inv21 = 1;
    65: op1_03_inv21 = 1;
    66: op1_03_inv21 = 1;
    70: op1_03_inv21 = 1;
    71: op1_03_inv21 = 1;
    74: op1_03_inv21 = 1;
    76: op1_03_inv21 = 1;
    80: op1_03_inv21 = 1;
    81: op1_03_inv21 = 1;
    82: op1_03_inv21 = 1;
    84: op1_03_inv21 = 1;
    88: op1_03_inv21 = 1;
    91: op1_03_inv21 = 1;
    93: op1_03_inv21 = 1;
    95: op1_03_inv21 = 1;
    96: op1_03_inv21 = 1;
    default: op1_03_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in22 = imem06_in[35:32];
    6: op1_03_in22 = reg_0388;
    7: op1_03_in22 = reg_0712;
    8: op1_03_in22 = reg_0311;
    9: op1_03_in22 = reg_0955;
    10: op1_03_in22 = reg_0966;
    11: op1_03_in22 = reg_0631;
    12: op1_03_in22 = reg_0289;
    13: op1_03_in22 = reg_0805;
    14: op1_03_in22 = reg_0095;
    15: op1_03_in22 = reg_0070;
    16: op1_03_in22 = reg_0787;
    17: op1_03_in22 = reg_0503;
    18: op1_03_in22 = reg_0834;
    58: op1_03_in22 = reg_0834;
    19: op1_03_in22 = reg_0353;
    20: op1_03_in22 = reg_0512;
    21: op1_03_in22 = reg_0249;
    22: op1_03_in22 = imem05_in[7:4];
    23: op1_03_in22 = reg_0604;
    24: op1_03_in22 = reg_0385;
    25: op1_03_in22 = imem07_in[107:104];
    26: op1_03_in22 = reg_1017;
    27: op1_03_in22 = imem07_in[95:92];
    28: op1_03_in22 = imem01_in[99:96];
    29: op1_03_in22 = reg_0813;
    30: op1_03_in22 = reg_0386;
    31: op1_03_in22 = reg_0223;
    32: op1_03_in22 = reg_0980;
    33: op1_03_in22 = imem06_in[63:60];
    34: op1_03_in22 = reg_0449;
    35: op1_03_in22 = reg_0946;
    36: op1_03_in22 = imem04_in[87:84];
    37: op1_03_in22 = reg_0827;
    38: op1_03_in22 = reg_1046;
    39: op1_03_in22 = imem06_in[127:124];
    41: op1_03_in22 = reg_0701;
    42: op1_03_in22 = reg_0867;
    43: op1_03_in22 = reg_0568;
    44: op1_03_in22 = imem07_in[19:16];
    45: op1_03_in22 = reg_0194;
    46: op1_03_in22 = reg_0343;
    47: op1_03_in22 = reg_0627;
    48: op1_03_in22 = reg_0709;
    49: op1_03_in22 = reg_0807;
    50: op1_03_in22 = reg_0656;
    51: op1_03_in22 = imem01_in[127:124];
    52: op1_03_in22 = reg_0702;
    54: op1_03_in22 = reg_0274;
    55: op1_03_in22 = imem02_in[3:0];
    56: op1_03_in22 = reg_0772;
    57: op1_03_in22 = reg_0050;
    59: op1_03_in22 = reg_0099;
    60: op1_03_in22 = reg_0617;
    61: op1_03_in22 = imem05_in[63:60];
    97: op1_03_in22 = imem05_in[63:60];
    62: op1_03_in22 = reg_0735;
    63: op1_03_in22 = imem01_in[39:36];
    64: op1_03_in22 = reg_0514;
    65: op1_03_in22 = imem03_in[75:72];
    66: op1_03_in22 = imem03_in[23:20];
    67: op1_03_in22 = reg_0664;
    68: op1_03_in22 = imem04_in[91:88];
    70: op1_03_in22 = reg_0520;
    71: op1_03_in22 = reg_1057;
    72: op1_03_in22 = reg_0968;
    73: op1_03_in22 = reg_0837;
    74: op1_03_in22 = imem03_in[123:120];
    75: op1_03_in22 = imem05_in[27:24];
    76: op1_03_in22 = reg_0405;
    77: op1_03_in22 = reg_0446;
    79: op1_03_in22 = reg_0083;
    80: op1_03_in22 = reg_0357;
    81: op1_03_in22 = reg_0409;
    82: op1_03_in22 = reg_0536;
    84: op1_03_in22 = reg_0011;
    85: op1_03_in22 = imem03_in[55:52];
    86: op1_03_in22 = reg_0332;
    87: op1_03_in22 = imem01_in[71:68];
    88: op1_03_in22 = reg_0546;
    89: op1_03_in22 = reg_0448;
    90: op1_03_in22 = reg_0585;
    91: op1_03_in22 = reg_0672;
    92: op1_03_in22 = reg_0312;
    93: op1_03_in22 = reg_0628;
    94: op1_03_in22 = imem07_in[119:116];
    95: op1_03_in22 = imem07_in[27:24];
    96: op1_03_in22 = reg_0084;
    default: op1_03_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv22 = 1;
    6: op1_03_inv22 = 1;
    7: op1_03_inv22 = 1;
    9: op1_03_inv22 = 1;
    11: op1_03_inv22 = 1;
    12: op1_03_inv22 = 1;
    13: op1_03_inv22 = 1;
    14: op1_03_inv22 = 1;
    16: op1_03_inv22 = 1;
    17: op1_03_inv22 = 1;
    19: op1_03_inv22 = 1;
    20: op1_03_inv22 = 1;
    22: op1_03_inv22 = 1;
    24: op1_03_inv22 = 1;
    25: op1_03_inv22 = 1;
    26: op1_03_inv22 = 1;
    28: op1_03_inv22 = 1;
    29: op1_03_inv22 = 1;
    31: op1_03_inv22 = 1;
    32: op1_03_inv22 = 1;
    33: op1_03_inv22 = 1;
    34: op1_03_inv22 = 1;
    36: op1_03_inv22 = 1;
    38: op1_03_inv22 = 1;
    41: op1_03_inv22 = 1;
    42: op1_03_inv22 = 1;
    43: op1_03_inv22 = 1;
    44: op1_03_inv22 = 1;
    45: op1_03_inv22 = 1;
    46: op1_03_inv22 = 1;
    52: op1_03_inv22 = 1;
    55: op1_03_inv22 = 1;
    57: op1_03_inv22 = 1;
    58: op1_03_inv22 = 1;
    59: op1_03_inv22 = 1;
    60: op1_03_inv22 = 1;
    64: op1_03_inv22 = 1;
    66: op1_03_inv22 = 1;
    67: op1_03_inv22 = 1;
    68: op1_03_inv22 = 1;
    71: op1_03_inv22 = 1;
    72: op1_03_inv22 = 1;
    74: op1_03_inv22 = 1;
    76: op1_03_inv22 = 1;
    80: op1_03_inv22 = 1;
    82: op1_03_inv22 = 1;
    89: op1_03_inv22 = 1;
    90: op1_03_inv22 = 1;
    91: op1_03_inv22 = 1;
    93: op1_03_inv22 = 1;
    94: op1_03_inv22 = 1;
    95: op1_03_inv22 = 1;
    96: op1_03_inv22 = 1;
    default: op1_03_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in23 = imem06_in[63:60];
    6: op1_03_in23 = reg_0323;
    7: op1_03_in23 = reg_0708;
    8: op1_03_in23 = reg_0369;
    9: op1_03_in23 = reg_0957;
    10: op1_03_in23 = reg_0944;
    11: op1_03_in23 = reg_0622;
    12: op1_03_in23 = reg_0306;
    13: op1_03_in23 = reg_1011;
    14: op1_03_in23 = reg_0086;
    15: op1_03_in23 = imem05_in[27:24];
    86: op1_03_in23 = imem05_in[27:24];
    16: op1_03_in23 = reg_0800;
    17: op1_03_in23 = reg_0234;
    18: op1_03_in23 = reg_0252;
    19: op1_03_in23 = reg_0347;
    20: op1_03_in23 = reg_0529;
    21: op1_03_in23 = reg_1039;
    22: op1_03_in23 = imem05_in[83:80];
    23: op1_03_in23 = reg_0611;
    24: op1_03_in23 = reg_0376;
    91: op1_03_in23 = reg_0376;
    25: op1_03_in23 = imem07_in[115:112];
    26: op1_03_in23 = reg_1038;
    27: op1_03_in23 = imem07_in[119:116];
    28: op1_03_in23 = imem01_in[115:112];
    29: op1_03_in23 = reg_0816;
    30: op1_03_in23 = reg_0243;
    31: op1_03_in23 = reg_0560;
    32: op1_03_in23 = reg_0983;
    33: op1_03_in23 = imem06_in[67:64];
    34: op1_03_in23 = reg_0444;
    35: op1_03_in23 = reg_0952;
    36: op1_03_in23 = imem04_in[107:104];
    37: op1_03_in23 = reg_0491;
    38: op1_03_in23 = reg_0831;
    39: op1_03_in23 = reg_0385;
    41: op1_03_in23 = reg_0430;
    42: op1_03_in23 = reg_0876;
    43: op1_03_in23 = reg_0066;
    44: op1_03_in23 = imem07_in[127:124];
    45: op1_03_in23 = reg_0206;
    46: op1_03_in23 = reg_1019;
    47: op1_03_in23 = reg_0754;
    48: op1_03_in23 = reg_0711;
    49: op1_03_in23 = reg_0836;
    50: op1_03_in23 = reg_0082;
    51: op1_03_in23 = reg_0786;
    52: op1_03_in23 = reg_0805;
    54: op1_03_in23 = reg_1045;
    55: op1_03_in23 = imem02_in[27:24];
    56: op1_03_in23 = reg_0482;
    79: op1_03_in23 = reg_0482;
    57: op1_03_in23 = reg_0507;
    58: op1_03_in23 = reg_0078;
    59: op1_03_in23 = reg_0245;
    60: op1_03_in23 = reg_0863;
    61: op1_03_in23 = imem05_in[79:76];
    62: op1_03_in23 = reg_0028;
    63: op1_03_in23 = imem01_in[55:52];
    64: op1_03_in23 = reg_0227;
    65: op1_03_in23 = imem03_in[83:80];
    66: op1_03_in23 = imem03_in[27:24];
    67: op1_03_in23 = reg_0394;
    68: op1_03_in23 = reg_0048;
    70: op1_03_in23 = reg_1040;
    71: op1_03_in23 = reg_0540;
    72: op1_03_in23 = reg_0337;
    73: op1_03_in23 = reg_0645;
    74: op1_03_in23 = reg_0012;
    75: op1_03_in23 = imem05_in[31:28];
    76: op1_03_in23 = reg_0264;
    77: op1_03_in23 = reg_0250;
    80: op1_03_in23 = reg_0228;
    81: op1_03_in23 = reg_0251;
    82: op1_03_in23 = reg_0301;
    84: op1_03_in23 = reg_0834;
    85: op1_03_in23 = imem03_in[59:56];
    87: op1_03_in23 = imem01_in[95:92];
    88: op1_03_in23 = reg_1023;
    89: op1_03_in23 = reg_0057;
    90: op1_03_in23 = reg_0352;
    92: op1_03_in23 = reg_0938;
    93: op1_03_in23 = imem07_in[43:40];
    94: op1_03_in23 = imem07_in[123:120];
    95: op1_03_in23 = imem07_in[31:28];
    96: op1_03_in23 = imem07_in[39:36];
    97: op1_03_in23 = imem05_in[71:68];
    default: op1_03_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv23 = 1;
    6: op1_03_inv23 = 1;
    7: op1_03_inv23 = 1;
    8: op1_03_inv23 = 1;
    9: op1_03_inv23 = 1;
    12: op1_03_inv23 = 1;
    14: op1_03_inv23 = 1;
    18: op1_03_inv23 = 1;
    19: op1_03_inv23 = 1;
    24: op1_03_inv23 = 1;
    26: op1_03_inv23 = 1;
    29: op1_03_inv23 = 1;
    32: op1_03_inv23 = 1;
    36: op1_03_inv23 = 1;
    38: op1_03_inv23 = 1;
    39: op1_03_inv23 = 1;
    41: op1_03_inv23 = 1;
    42: op1_03_inv23 = 1;
    44: op1_03_inv23 = 1;
    47: op1_03_inv23 = 1;
    51: op1_03_inv23 = 1;
    54: op1_03_inv23 = 1;
    55: op1_03_inv23 = 1;
    59: op1_03_inv23 = 1;
    60: op1_03_inv23 = 1;
    64: op1_03_inv23 = 1;
    65: op1_03_inv23 = 1;
    67: op1_03_inv23 = 1;
    68: op1_03_inv23 = 1;
    70: op1_03_inv23 = 1;
    71: op1_03_inv23 = 1;
    74: op1_03_inv23 = 1;
    75: op1_03_inv23 = 1;
    77: op1_03_inv23 = 1;
    79: op1_03_inv23 = 1;
    84: op1_03_inv23 = 1;
    85: op1_03_inv23 = 1;
    87: op1_03_inv23 = 1;
    88: op1_03_inv23 = 1;
    90: op1_03_inv23 = 1;
    91: op1_03_inv23 = 1;
    93: op1_03_inv23 = 1;
    94: op1_03_inv23 = 1;
    96: op1_03_inv23 = 1;
    97: op1_03_inv23 = 1;
    default: op1_03_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in24 = imem06_in[111:108];
    6: op1_03_in24 = reg_0389;
    67: op1_03_in24 = reg_0389;
    7: op1_03_in24 = reg_0445;
    8: op1_03_in24 = reg_0323;
    9: op1_03_in24 = reg_0950;
    10: op1_03_in24 = reg_0959;
    11: op1_03_in24 = reg_0381;
    12: op1_03_in24 = reg_0292;
    13: op1_03_in24 = reg_0005;
    14: op1_03_in24 = reg_0094;
    15: op1_03_in24 = imem05_in[47:44];
    16: op1_03_in24 = reg_0802;
    57: op1_03_in24 = reg_0802;
    17: op1_03_in24 = reg_1042;
    18: op1_03_in24 = reg_0832;
    19: op1_03_in24 = reg_0086;
    42: op1_03_in24 = reg_0086;
    20: op1_03_in24 = reg_0962;
    21: op1_03_in24 = reg_1043;
    22: op1_03_in24 = imem05_in[103:100];
    23: op1_03_in24 = reg_0332;
    81: op1_03_in24 = reg_0332;
    24: op1_03_in24 = reg_0331;
    25: op1_03_in24 = reg_0730;
    26: op1_03_in24 = reg_0122;
    27: op1_03_in24 = imem07_in[123:120];
    28: op1_03_in24 = reg_0013;
    29: op1_03_in24 = reg_0275;
    30: op1_03_in24 = reg_0000;
    31: op1_03_in24 = reg_0510;
    32: op1_03_in24 = imem04_in[11:8];
    33: op1_03_in24 = imem06_in[95:92];
    34: op1_03_in24 = reg_0443;
    35: op1_03_in24 = reg_0960;
    36: op1_03_in24 = reg_0536;
    37: op1_03_in24 = reg_0260;
    38: op1_03_in24 = reg_0148;
    39: op1_03_in24 = reg_0295;
    41: op1_03_in24 = reg_0432;
    43: op1_03_in24 = reg_0068;
    44: op1_03_in24 = reg_0703;
    45: op1_03_in24 = imem01_in[39:36];
    46: op1_03_in24 = reg_0046;
    47: op1_03_in24 = reg_0294;
    48: op1_03_in24 = reg_0421;
    49: op1_03_in24 = reg_0999;
    50: op1_03_in24 = reg_0565;
    51: op1_03_in24 = reg_0779;
    52: op1_03_in24 = reg_0422;
    54: op1_03_in24 = reg_0238;
    55: op1_03_in24 = imem02_in[115:112];
    56: op1_03_in24 = reg_0758;
    58: op1_03_in24 = reg_0053;
    59: op1_03_in24 = reg_0585;
    60: op1_03_in24 = reg_0632;
    61: op1_03_in24 = reg_0215;
    62: op1_03_in24 = reg_1030;
    63: op1_03_in24 = imem01_in[79:76];
    64: op1_03_in24 = reg_0740;
    65: op1_03_in24 = reg_0006;
    66: op1_03_in24 = imem03_in[39:36];
    68: op1_03_in24 = reg_1005;
    70: op1_03_in24 = reg_0354;
    71: op1_03_in24 = reg_0909;
    72: op1_03_in24 = reg_0546;
    73: op1_03_in24 = reg_0423;
    74: op1_03_in24 = reg_0345;
    75: op1_03_in24 = imem05_in[75:72];
    76: op1_03_in24 = reg_0715;
    77: op1_03_in24 = reg_0325;
    79: op1_03_in24 = reg_0506;
    80: op1_03_in24 = reg_0756;
    82: op1_03_in24 = reg_0277;
    84: op1_03_in24 = reg_0403;
    85: op1_03_in24 = reg_0760;
    86: op1_03_in24 = imem05_in[43:40];
    87: op1_03_in24 = imem01_in[107:104];
    88: op1_03_in24 = reg_0234;
    89: op1_03_in24 = reg_0646;
    90: op1_03_in24 = reg_0983;
    91: op1_03_in24 = reg_0597;
    92: op1_03_in24 = reg_0989;
    93: op1_03_in24 = imem07_in[79:76];
    94: op1_03_in24 = reg_0728;
    95: op1_03_in24 = imem07_in[63:60];
    96: op1_03_in24 = imem07_in[43:40];
    97: op1_03_in24 = imem05_in[79:76];
    default: op1_03_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_03_inv24 = 1;
    9: op1_03_inv24 = 1;
    10: op1_03_inv24 = 1;
    12: op1_03_inv24 = 1;
    14: op1_03_inv24 = 1;
    15: op1_03_inv24 = 1;
    18: op1_03_inv24 = 1;
    24: op1_03_inv24 = 1;
    25: op1_03_inv24 = 1;
    28: op1_03_inv24 = 1;
    30: op1_03_inv24 = 1;
    31: op1_03_inv24 = 1;
    32: op1_03_inv24 = 1;
    35: op1_03_inv24 = 1;
    36: op1_03_inv24 = 1;
    39: op1_03_inv24 = 1;
    41: op1_03_inv24 = 1;
    43: op1_03_inv24 = 1;
    44: op1_03_inv24 = 1;
    46: op1_03_inv24 = 1;
    47: op1_03_inv24 = 1;
    49: op1_03_inv24 = 1;
    51: op1_03_inv24 = 1;
    54: op1_03_inv24 = 1;
    60: op1_03_inv24 = 1;
    61: op1_03_inv24 = 1;
    62: op1_03_inv24 = 1;
    63: op1_03_inv24 = 1;
    64: op1_03_inv24 = 1;
    65: op1_03_inv24 = 1;
    66: op1_03_inv24 = 1;
    73: op1_03_inv24 = 1;
    74: op1_03_inv24 = 1;
    76: op1_03_inv24 = 1;
    79: op1_03_inv24 = 1;
    84: op1_03_inv24 = 1;
    87: op1_03_inv24 = 1;
    88: op1_03_inv24 = 1;
    90: op1_03_inv24 = 1;
    91: op1_03_inv24 = 1;
    96: op1_03_inv24 = 1;
    97: op1_03_inv24 = 1;
    default: op1_03_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in25 = reg_0620;
    6: op1_03_in25 = imem03_in[3:0];
    7: op1_03_in25 = reg_0435;
    8: op1_03_in25 = reg_0397;
    9: op1_03_in25 = reg_0945;
    10: op1_03_in25 = reg_0955;
    11: op1_03_in25 = reg_0372;
    12: op1_03_in25 = reg_0286;
    13: op1_03_in25 = reg_0754;
    14: op1_03_in25 = reg_0093;
    15: op1_03_in25 = imem05_in[95:92];
    16: op1_03_in25 = imem07_in[3:0];
    17: op1_03_in25 = reg_0500;
    18: op1_03_in25 = reg_0150;
    19: op1_03_in25 = reg_0090;
    42: op1_03_in25 = reg_0090;
    20: op1_03_in25 = reg_0973;
    21: op1_03_in25 = reg_1044;
    51: op1_03_in25 = reg_1044;
    22: op1_03_in25 = imem05_in[111:108];
    23: op1_03_in25 = reg_0356;
    24: op1_03_in25 = reg_0992;
    25: op1_03_in25 = reg_0709;
    26: op1_03_in25 = reg_0113;
    27: op1_03_in25 = reg_0716;
    28: op1_03_in25 = reg_0786;
    29: op1_03_in25 = reg_1046;
    30: op1_03_in25 = reg_0027;
    31: op1_03_in25 = reg_0860;
    32: op1_03_in25 = imem04_in[35:32];
    33: op1_03_in25 = imem06_in[103:100];
    34: op1_03_in25 = reg_0420;
    35: op1_03_in25 = reg_0491;
    36: op1_03_in25 = reg_0511;
    37: op1_03_in25 = reg_0254;
    38: op1_03_in25 = reg_0146;
    39: op1_03_in25 = reg_0399;
    41: op1_03_in25 = reg_0426;
    43: op1_03_in25 = reg_0748;
    44: op1_03_in25 = reg_0729;
    45: op1_03_in25 = imem01_in[71:68];
    46: op1_03_in25 = reg_0824;
    47: op1_03_in25 = reg_0741;
    48: op1_03_in25 = reg_0406;
    77: op1_03_in25 = reg_0406;
    49: op1_03_in25 = reg_0977;
    50: op1_03_in25 = reg_0300;
    52: op1_03_in25 = reg_0315;
    54: op1_03_in25 = reg_0496;
    55: op1_03_in25 = imem02_in[119:116];
    56: op1_03_in25 = reg_0085;
    57: op1_03_in25 = reg_0568;
    58: op1_03_in25 = reg_0578;
    59: op1_03_in25 = reg_0298;
    60: op1_03_in25 = reg_0011;
    61: op1_03_in25 = reg_0757;
    62: op1_03_in25 = reg_0595;
    63: op1_03_in25 = imem01_in[87:84];
    64: op1_03_in25 = reg_0232;
    65: op1_03_in25 = reg_0535;
    66: op1_03_in25 = imem03_in[67:64];
    67: op1_03_in25 = reg_0867;
    68: op1_03_in25 = reg_1016;
    70: op1_03_in25 = reg_1017;
    71: op1_03_in25 = reg_0850;
    72: op1_03_in25 = reg_0962;
    73: op1_03_in25 = reg_0368;
    74: op1_03_in25 = reg_0580;
    75: op1_03_in25 = imem05_in[87:84];
    76: op1_03_in25 = reg_0250;
    79: op1_03_in25 = reg_0310;
    80: op1_03_in25 = reg_0038;
    81: op1_03_in25 = imem05_in[63:60];
    82: op1_03_in25 = reg_1057;
    84: op1_03_in25 = reg_0782;
    85: op1_03_in25 = reg_0445;
    86: op1_03_in25 = imem05_in[103:100];
    87: op1_03_in25 = reg_0122;
    88: op1_03_in25 = reg_0487;
    89: op1_03_in25 = reg_0964;
    90: op1_03_in25 = reg_0240;
    91: op1_03_in25 = reg_0588;
    92: op1_03_in25 = reg_0981;
    93: op1_03_in25 = imem07_in[111:108];
    94: op1_03_in25 = reg_0159;
    95: op1_03_in25 = reg_0567;
    96: op1_03_in25 = imem07_in[115:112];
    97: op1_03_in25 = imem05_in[123:120];
    default: op1_03_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv25 = 1;
    6: op1_03_inv25 = 1;
    7: op1_03_inv25 = 1;
    9: op1_03_inv25 = 1;
    15: op1_03_inv25 = 1;
    21: op1_03_inv25 = 1;
    23: op1_03_inv25 = 1;
    24: op1_03_inv25 = 1;
    30: op1_03_inv25 = 1;
    31: op1_03_inv25 = 1;
    37: op1_03_inv25 = 1;
    38: op1_03_inv25 = 1;
    41: op1_03_inv25 = 1;
    43: op1_03_inv25 = 1;
    44: op1_03_inv25 = 1;
    45: op1_03_inv25 = 1;
    49: op1_03_inv25 = 1;
    54: op1_03_inv25 = 1;
    55: op1_03_inv25 = 1;
    58: op1_03_inv25 = 1;
    60: op1_03_inv25 = 1;
    62: op1_03_inv25 = 1;
    63: op1_03_inv25 = 1;
    64: op1_03_inv25 = 1;
    65: op1_03_inv25 = 1;
    68: op1_03_inv25 = 1;
    70: op1_03_inv25 = 1;
    71: op1_03_inv25 = 1;
    72: op1_03_inv25 = 1;
    75: op1_03_inv25 = 1;
    77: op1_03_inv25 = 1;
    79: op1_03_inv25 = 1;
    82: op1_03_inv25 = 1;
    84: op1_03_inv25 = 1;
    85: op1_03_inv25 = 1;
    88: op1_03_inv25 = 1;
    89: op1_03_inv25 = 1;
    90: op1_03_inv25 = 1;
    94: op1_03_inv25 = 1;
    95: op1_03_inv25 = 1;
    default: op1_03_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in26 = reg_0621;
    6: op1_03_in26 = imem03_in[75:72];
    7: op1_03_in26 = reg_0175;
    8: op1_03_in26 = reg_0393;
    9: op1_03_in26 = reg_0946;
    10: op1_03_in26 = reg_0969;
    11: op1_03_in26 = reg_0405;
    12: op1_03_in26 = reg_0275;
    13: op1_03_in26 = imem07_in[31:28];
    14: op1_03_in26 = imem03_in[3:0];
    15: op1_03_in26 = imem05_in[127:124];
    16: op1_03_in26 = imem07_in[39:36];
    17: op1_03_in26 = reg_1017;
    18: op1_03_in26 = reg_0151;
    19: op1_03_in26 = reg_0087;
    20: op1_03_in26 = reg_0964;
    21: op1_03_in26 = reg_0500;
    22: op1_03_in26 = reg_0973;
    23: op1_03_in26 = reg_0372;
    24: op1_03_in26 = reg_0993;
    25: op1_03_in26 = reg_0718;
    26: op1_03_in26 = reg_0743;
    27: op1_03_in26 = reg_0704;
    28: op1_03_in26 = reg_0218;
    29: op1_03_in26 = reg_0832;
    64: op1_03_in26 = reg_0832;
    30: op1_03_in26 = reg_0026;
    31: op1_03_in26 = reg_0811;
    32: op1_03_in26 = imem04_in[43:40];
    33: op1_03_in26 = imem06_in[115:112];
    34: op1_03_in26 = reg_0180;
    35: op1_03_in26 = reg_0813;
    36: op1_03_in26 = reg_0265;
    37: op1_03_in26 = reg_0896;
    38: op1_03_in26 = reg_0130;
    39: op1_03_in26 = reg_0617;
    41: op1_03_in26 = reg_0428;
    42: op1_03_in26 = reg_0016;
    79: op1_03_in26 = reg_0016;
    43: op1_03_in26 = reg_0777;
    44: op1_03_in26 = reg_0711;
    45: op1_03_in26 = imem01_in[83:80];
    46: op1_03_in26 = reg_0389;
    73: op1_03_in26 = reg_0389;
    47: op1_03_in26 = reg_0264;
    48: op1_03_in26 = reg_0353;
    49: op1_03_in26 = reg_0990;
    50: op1_03_in26 = reg_0648;
    51: op1_03_in26 = reg_0904;
    52: op1_03_in26 = reg_0589;
    54: op1_03_in26 = reg_1043;
    55: op1_03_in26 = reg_0642;
    56: op1_03_in26 = reg_0310;
    57: op1_03_in26 = reg_0058;
    58: op1_03_in26 = reg_0593;
    59: op1_03_in26 = reg_0576;
    60: op1_03_in26 = reg_0628;
    61: op1_03_in26 = reg_0435;
    62: op1_03_in26 = reg_0556;
    63: op1_03_in26 = reg_0918;
    65: op1_03_in26 = reg_0046;
    74: op1_03_in26 = reg_0046;
    66: op1_03_in26 = reg_1007;
    67: op1_03_in26 = reg_0814;
    68: op1_03_in26 = reg_0932;
    70: op1_03_in26 = reg_0906;
    71: op1_03_in26 = reg_0014;
    72: op1_03_in26 = reg_0604;
    88: op1_03_in26 = reg_0604;
    75: op1_03_in26 = reg_0215;
    76: op1_03_in26 = reg_0426;
    77: op1_03_in26 = reg_0532;
    80: op1_03_in26 = reg_0672;
    81: op1_03_in26 = imem05_in[67:64];
    82: op1_03_in26 = reg_1020;
    84: op1_03_in26 = reg_0573;
    85: op1_03_in26 = reg_0547;
    86: op1_03_in26 = reg_1021;
    87: op1_03_in26 = reg_0337;
    89: op1_03_in26 = reg_0530;
    90: op1_03_in26 = reg_0859;
    91: op1_03_in26 = reg_0975;
    92: op1_03_in26 = reg_0825;
    93: op1_03_in26 = reg_0165;
    94: op1_03_in26 = reg_0717;
    95: op1_03_in26 = reg_0717;
    96: op1_03_in26 = reg_0722;
    97: op1_03_in26 = reg_0652;
    default: op1_03_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv26 = 1;
    7: op1_03_inv26 = 1;
    10: op1_03_inv26 = 1;
    11: op1_03_inv26 = 1;
    12: op1_03_inv26 = 1;
    18: op1_03_inv26 = 1;
    19: op1_03_inv26 = 1;
    20: op1_03_inv26 = 1;
    21: op1_03_inv26 = 1;
    22: op1_03_inv26 = 1;
    25: op1_03_inv26 = 1;
    27: op1_03_inv26 = 1;
    28: op1_03_inv26 = 1;
    29: op1_03_inv26 = 1;
    31: op1_03_inv26 = 1;
    32: op1_03_inv26 = 1;
    33: op1_03_inv26 = 1;
    35: op1_03_inv26 = 1;
    37: op1_03_inv26 = 1;
    39: op1_03_inv26 = 1;
    42: op1_03_inv26 = 1;
    44: op1_03_inv26 = 1;
    47: op1_03_inv26 = 1;
    54: op1_03_inv26 = 1;
    56: op1_03_inv26 = 1;
    62: op1_03_inv26 = 1;
    66: op1_03_inv26 = 1;
    67: op1_03_inv26 = 1;
    71: op1_03_inv26 = 1;
    72: op1_03_inv26 = 1;
    75: op1_03_inv26 = 1;
    76: op1_03_inv26 = 1;
    80: op1_03_inv26 = 1;
    82: op1_03_inv26 = 1;
    84: op1_03_inv26 = 1;
    86: op1_03_inv26 = 1;
    87: op1_03_inv26 = 1;
    88: op1_03_inv26 = 1;
    90: op1_03_inv26 = 1;
    91: op1_03_inv26 = 1;
    93: op1_03_inv26 = 1;
    94: op1_03_inv26 = 1;
    95: op1_03_inv26 = 1;
    96: op1_03_inv26 = 1;
    97: op1_03_inv26 = 1;
    default: op1_03_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in27 = reg_0622;
    60: op1_03_in27 = reg_0622;
    6: op1_03_in27 = imem04_in[3:0];
    91: op1_03_in27 = imem04_in[3:0];
    7: op1_03_in27 = reg_0172;
    48: op1_03_in27 = reg_0172;
    8: op1_03_in27 = reg_0985;
    9: op1_03_in27 = reg_0943;
    10: op1_03_in27 = reg_0964;
    11: op1_03_in27 = reg_0375;
    12: op1_03_in27 = reg_0288;
    13: op1_03_in27 = imem07_in[75:72];
    14: op1_03_in27 = imem03_in[11:8];
    15: op1_03_in27 = reg_0958;
    16: op1_03_in27 = imem07_in[43:40];
    17: op1_03_in27 = reg_1038;
    18: op1_03_in27 = reg_0146;
    19: op1_03_in27 = reg_0094;
    20: op1_03_in27 = reg_0965;
    21: op1_03_in27 = reg_1041;
    22: op1_03_in27 = reg_0971;
    23: op1_03_in27 = reg_0407;
    24: op1_03_in27 = reg_0877;
    25: op1_03_in27 = reg_0706;
    26: op1_03_in27 = reg_0833;
    27: op1_03_in27 = reg_0726;
    28: op1_03_in27 = reg_0860;
    29: op1_03_in27 = reg_0831;
    30: op1_03_in27 = reg_0808;
    31: op1_03_in27 = reg_0238;
    32: op1_03_in27 = imem04_in[59:56];
    33: op1_03_in27 = reg_0609;
    39: op1_03_in27 = reg_0609;
    34: op1_03_in27 = reg_0161;
    35: op1_03_in27 = reg_0229;
    36: op1_03_in27 = reg_0912;
    37: op1_03_in27 = reg_0156;
    38: op1_03_in27 = reg_0144;
    41: op1_03_in27 = reg_0443;
    42: op1_03_in27 = reg_0872;
    79: op1_03_in27 = reg_0872;
    43: op1_03_in27 = reg_0057;
    44: op1_03_in27 = reg_0700;
    45: op1_03_in27 = imem01_in[99:96];
    46: op1_03_in27 = reg_0377;
    47: op1_03_in27 = reg_0399;
    49: op1_03_in27 = reg_1000;
    50: op1_03_in27 = reg_0837;
    51: op1_03_in27 = reg_0933;
    52: op1_03_in27 = reg_0175;
    54: op1_03_in27 = reg_0829;
    55: op1_03_in27 = reg_0650;
    56: op1_03_in27 = reg_0016;
    57: op1_03_in27 = reg_0056;
    58: op1_03_in27 = reg_0031;
    59: op1_03_in27 = reg_0784;
    61: op1_03_in27 = reg_0336;
    62: op1_03_in27 = reg_0632;
    63: op1_03_in27 = reg_0586;
    64: op1_03_in27 = reg_0745;
    65: op1_03_in27 = reg_0576;
    66: op1_03_in27 = reg_0240;
    85: op1_03_in27 = reg_0240;
    67: op1_03_in27 = reg_0484;
    68: op1_03_in27 = reg_0061;
    70: op1_03_in27 = reg_0615;
    71: op1_03_in27 = reg_0296;
    72: op1_03_in27 = reg_0520;
    88: op1_03_in27 = reg_0520;
    73: op1_03_in27 = reg_0792;
    74: op1_03_in27 = reg_0396;
    75: op1_03_in27 = reg_0866;
    76: op1_03_in27 = reg_0047;
    77: op1_03_in27 = reg_0599;
    80: op1_03_in27 = reg_0312;
    81: op1_03_in27 = imem05_in[119:116];
    82: op1_03_in27 = reg_0778;
    84: op1_03_in27 = imem07_in[19:16];
    86: op1_03_in27 = reg_0141;
    87: op1_03_in27 = reg_0120;
    89: op1_03_in27 = reg_0795;
    90: op1_03_in27 = reg_0301;
    92: op1_03_in27 = reg_0318;
    93: op1_03_in27 = reg_0720;
    96: op1_03_in27 = reg_0720;
    94: op1_03_in27 = reg_0923;
    95: op1_03_in27 = reg_0560;
    97: op1_03_in27 = reg_0954;
    default: op1_03_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv27 = 1;
    6: op1_03_inv27 = 1;
    10: op1_03_inv27 = 1;
    11: op1_03_inv27 = 1;
    12: op1_03_inv27 = 1;
    14: op1_03_inv27 = 1;
    16: op1_03_inv27 = 1;
    17: op1_03_inv27 = 1;
    25: op1_03_inv27 = 1;
    27: op1_03_inv27 = 1;
    29: op1_03_inv27 = 1;
    34: op1_03_inv27 = 1;
    35: op1_03_inv27 = 1;
    36: op1_03_inv27 = 1;
    37: op1_03_inv27 = 1;
    38: op1_03_inv27 = 1;
    39: op1_03_inv27 = 1;
    41: op1_03_inv27 = 1;
    42: op1_03_inv27 = 1;
    43: op1_03_inv27 = 1;
    44: op1_03_inv27 = 1;
    47: op1_03_inv27 = 1;
    51: op1_03_inv27 = 1;
    55: op1_03_inv27 = 1;
    56: op1_03_inv27 = 1;
    58: op1_03_inv27 = 1;
    60: op1_03_inv27 = 1;
    62: op1_03_inv27 = 1;
    63: op1_03_inv27 = 1;
    65: op1_03_inv27 = 1;
    68: op1_03_inv27 = 1;
    73: op1_03_inv27 = 1;
    76: op1_03_inv27 = 1;
    77: op1_03_inv27 = 1;
    85: op1_03_inv27 = 1;
    90: op1_03_inv27 = 1;
    92: op1_03_inv27 = 1;
    default: op1_03_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in28 = reg_0623;
    6: op1_03_in28 = imem04_in[23:20];
    7: op1_03_in28 = reg_0181;
    8: op1_03_in28 = reg_0994;
    9: op1_03_in28 = reg_0267;
    10: op1_03_in28 = reg_0951;
    11: op1_03_in28 = reg_0404;
    12: op1_03_in28 = reg_0307;
    13: op1_03_in28 = imem07_in[83:80];
    14: op1_03_in28 = imem03_in[15:12];
    15: op1_03_in28 = reg_0955;
    16: op1_03_in28 = imem07_in[47:44];
    17: op1_03_in28 = reg_0105;
    18: op1_03_in28 = reg_0138;
    19: op1_03_in28 = imem03_in[11:8];
    42: op1_03_in28 = imem03_in[11:8];
    56: op1_03_in28 = imem03_in[11:8];
    20: op1_03_in28 = reg_0946;
    21: op1_03_in28 = reg_0871;
    22: op1_03_in28 = reg_0956;
    23: op1_03_in28 = reg_0337;
    24: op1_03_in28 = reg_0554;
    25: op1_03_in28 = reg_0425;
    26: op1_03_in28 = reg_0737;
    27: op1_03_in28 = reg_0725;
    28: op1_03_in28 = reg_0487;
    29: op1_03_in28 = reg_0147;
    30: op1_03_in28 = reg_0486;
    31: op1_03_in28 = reg_0249;
    32: op1_03_in28 = imem04_in[71:68];
    33: op1_03_in28 = reg_0622;
    34: op1_03_in28 = reg_0182;
    35: op1_03_in28 = reg_0254;
    36: op1_03_in28 = reg_0306;
    37: op1_03_in28 = reg_0752;
    82: op1_03_in28 = reg_0752;
    38: op1_03_in28 = imem06_in[23:20];
    39: op1_03_in28 = reg_1010;
    41: op1_03_in28 = reg_0175;
    43: op1_03_in28 = reg_0855;
    44: op1_03_in28 = reg_0361;
    45: op1_03_in28 = reg_0013;
    46: op1_03_in28 = reg_0312;
    47: op1_03_in28 = reg_1029;
    48: op1_03_in28 = reg_0167;
    49: op1_03_in28 = reg_0983;
    50: op1_03_in28 = reg_0334;
    51: op1_03_in28 = reg_0919;
    52: op1_03_in28 = reg_0180;
    54: op1_03_in28 = reg_0227;
    55: op1_03_in28 = reg_0363;
    57: op1_03_in28 = reg_0015;
    58: op1_03_in28 = imem05_in[27:24];
    59: op1_03_in28 = reg_0509;
    60: op1_03_in28 = imem07_in[3:0];
    61: op1_03_in28 = reg_0094;
    62: op1_03_in28 = reg_0386;
    63: op1_03_in28 = reg_0510;
    64: op1_03_in28 = imem02_in[47:44];
    65: op1_03_in28 = reg_0847;
    66: op1_03_in28 = reg_0370;
    67: op1_03_in28 = imem03_in[23:20];
    68: op1_03_in28 = reg_0432;
    70: op1_03_in28 = reg_1055;
    71: op1_03_in28 = reg_0809;
    72: op1_03_in28 = reg_0615;
    73: op1_03_in28 = reg_0484;
    74: op1_03_in28 = reg_0662;
    75: op1_03_in28 = reg_0954;
    76: op1_03_in28 = reg_0321;
    77: op1_03_in28 = reg_0868;
    79: op1_03_in28 = imem03_in[19:16];
    80: op1_03_in28 = reg_0820;
    81: op1_03_in28 = imem05_in[123:120];
    84: op1_03_in28 = imem07_in[59:56];
    85: op1_03_in28 = reg_0278;
    86: op1_03_in28 = reg_0963;
    87: op1_03_in28 = reg_0862;
    88: op1_03_in28 = reg_0514;
    89: op1_03_in28 = reg_0528;
    90: op1_03_in28 = reg_0062;
    91: op1_03_in28 = imem04_in[19:16];
    92: op1_03_in28 = imem04_in[59:56];
    93: op1_03_in28 = reg_0221;
    94: op1_03_in28 = reg_0959;
    95: op1_03_in28 = reg_0903;
    96: op1_03_in28 = reg_0560;
    97: op1_03_in28 = reg_0448;
    default: op1_03_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv28 = 1;
    10: op1_03_inv28 = 1;
    12: op1_03_inv28 = 1;
    13: op1_03_inv28 = 1;
    14: op1_03_inv28 = 1;
    16: op1_03_inv28 = 1;
    17: op1_03_inv28 = 1;
    18: op1_03_inv28 = 1;
    19: op1_03_inv28 = 1;
    20: op1_03_inv28 = 1;
    26: op1_03_inv28 = 1;
    28: op1_03_inv28 = 1;
    29: op1_03_inv28 = 1;
    32: op1_03_inv28 = 1;
    33: op1_03_inv28 = 1;
    37: op1_03_inv28 = 1;
    41: op1_03_inv28 = 1;
    45: op1_03_inv28 = 1;
    47: op1_03_inv28 = 1;
    50: op1_03_inv28 = 1;
    57: op1_03_inv28 = 1;
    58: op1_03_inv28 = 1;
    59: op1_03_inv28 = 1;
    60: op1_03_inv28 = 1;
    61: op1_03_inv28 = 1;
    62: op1_03_inv28 = 1;
    63: op1_03_inv28 = 1;
    66: op1_03_inv28 = 1;
    68: op1_03_inv28 = 1;
    70: op1_03_inv28 = 1;
    73: op1_03_inv28 = 1;
    74: op1_03_inv28 = 1;
    75: op1_03_inv28 = 1;
    77: op1_03_inv28 = 1;
    79: op1_03_inv28 = 1;
    80: op1_03_inv28 = 1;
    82: op1_03_inv28 = 1;
    86: op1_03_inv28 = 1;
    87: op1_03_inv28 = 1;
    89: op1_03_inv28 = 1;
    92: op1_03_inv28 = 1;
    93: op1_03_inv28 = 1;
    94: op1_03_inv28 = 1;
    95: op1_03_inv28 = 1;
    97: op1_03_inv28 = 1;
    default: op1_03_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in29 = reg_0332;
    6: op1_03_in29 = imem04_in[71:68];
    7: op1_03_in29 = reg_0169;
    8: op1_03_in29 = imem04_in[3:0];
    9: op1_03_in29 = reg_0268;
    10: op1_03_in29 = reg_0949;
    11: op1_03_in29 = reg_0315;
    12: op1_03_in29 = reg_0062;
    13: op1_03_in29 = imem07_in[107:104];
    14: op1_03_in29 = imem03_in[55:52];
    15: op1_03_in29 = reg_0954;
    16: op1_03_in29 = imem07_in[63:60];
    17: op1_03_in29 = reg_0122;
    18: op1_03_in29 = reg_0129;
    19: op1_03_in29 = imem03_in[15:12];
    20: op1_03_in29 = imem05_in[59:56];
    21: op1_03_in29 = reg_1018;
    22: op1_03_in29 = reg_0957;
    23: op1_03_in29 = reg_0027;
    24: op1_03_in29 = reg_0559;
    25: op1_03_in29 = reg_0436;
    26: op1_03_in29 = reg_0545;
    27: op1_03_in29 = reg_0712;
    28: op1_03_in29 = reg_0249;
    29: op1_03_in29 = reg_0136;
    30: op1_03_in29 = reg_0783;
    31: op1_03_in29 = reg_0226;
    32: op1_03_in29 = imem04_in[99:96];
    33: op1_03_in29 = reg_0381;
    34: op1_03_in29 = reg_0170;
    35: op1_03_in29 = reg_0896;
    36: op1_03_in29 = reg_1057;
    37: op1_03_in29 = reg_0521;
    38: op1_03_in29 = imem06_in[91:88];
    39: op1_03_in29 = imem07_in[15:12];
    41: op1_03_in29 = reg_0167;
    42: op1_03_in29 = imem03_in[23:20];
    43: op1_03_in29 = imem05_in[11:8];
    44: op1_03_in29 = reg_0433;
    45: op1_03_in29 = reg_0563;
    46: op1_03_in29 = reg_0844;
    47: op1_03_in29 = reg_0894;
    48: op1_03_in29 = reg_0160;
    52: op1_03_in29 = reg_0160;
    49: op1_03_in29 = reg_0337;
    50: op1_03_in29 = reg_0842;
    51: op1_03_in29 = reg_1056;
    54: op1_03_in29 = reg_0216;
    55: op1_03_in29 = reg_0649;
    56: op1_03_in29 = imem03_in[43:40];
    57: op1_03_in29 = reg_0064;
    58: op1_03_in29 = imem05_in[51:48];
    59: op1_03_in29 = reg_0513;
    60: op1_03_in29 = imem07_in[47:44];
    61: op1_03_in29 = reg_0697;
    62: op1_03_in29 = reg_0449;
    63: op1_03_in29 = reg_1036;
    64: op1_03_in29 = imem02_in[55:52];
    65: op1_03_in29 = reg_0793;
    66: op1_03_in29 = reg_0038;
    67: op1_03_in29 = imem03_in[27:24];
    79: op1_03_in29 = imem03_in[27:24];
    68: op1_03_in29 = reg_0407;
    71: op1_03_in29 = reg_0407;
    70: op1_03_in29 = reg_0003;
    72: op1_03_in29 = reg_0832;
    73: op1_03_in29 = reg_0291;
    74: op1_03_in29 = reg_0756;
    75: op1_03_in29 = reg_0655;
    76: op1_03_in29 = reg_0419;
    77: op1_03_in29 = reg_0838;
    80: op1_03_in29 = reg_0996;
    81: op1_03_in29 = imem05_in[127:124];
    82: op1_03_in29 = reg_0568;
    84: op1_03_in29 = imem07_in[71:68];
    85: op1_03_in29 = reg_0239;
    86: op1_03_in29 = reg_0150;
    87: op1_03_in29 = reg_1039;
    88: op1_03_in29 = reg_0500;
    89: op1_03_in29 = reg_0490;
    90: op1_03_in29 = reg_0662;
    91: op1_03_in29 = imem04_in[23:20];
    92: op1_03_in29 = imem04_in[119:116];
    93: op1_03_in29 = reg_0560;
    94: op1_03_in29 = reg_0303;
    95: op1_03_in29 = reg_0350;
    96: op1_03_in29 = reg_0718;
    97: op1_03_in29 = reg_0057;
    default: op1_03_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv29 = 1;
    7: op1_03_inv29 = 1;
    8: op1_03_inv29 = 1;
    10: op1_03_inv29 = 1;
    14: op1_03_inv29 = 1;
    15: op1_03_inv29 = 1;
    17: op1_03_inv29 = 1;
    18: op1_03_inv29 = 1;
    19: op1_03_inv29 = 1;
    23: op1_03_inv29 = 1;
    24: op1_03_inv29 = 1;
    27: op1_03_inv29 = 1;
    28: op1_03_inv29 = 1;
    29: op1_03_inv29 = 1;
    30: op1_03_inv29 = 1;
    31: op1_03_inv29 = 1;
    32: op1_03_inv29 = 1;
    34: op1_03_inv29 = 1;
    37: op1_03_inv29 = 1;
    38: op1_03_inv29 = 1;
    41: op1_03_inv29 = 1;
    46: op1_03_inv29 = 1;
    50: op1_03_inv29 = 1;
    55: op1_03_inv29 = 1;
    57: op1_03_inv29 = 1;
    58: op1_03_inv29 = 1;
    63: op1_03_inv29 = 1;
    68: op1_03_inv29 = 1;
    70: op1_03_inv29 = 1;
    71: op1_03_inv29 = 1;
    73: op1_03_inv29 = 1;
    74: op1_03_inv29 = 1;
    75: op1_03_inv29 = 1;
    80: op1_03_inv29 = 1;
    81: op1_03_inv29 = 1;
    82: op1_03_inv29 = 1;
    84: op1_03_inv29 = 1;
    86: op1_03_inv29 = 1;
    90: op1_03_inv29 = 1;
    94: op1_03_inv29 = 1;
    95: op1_03_inv29 = 1;
    97: op1_03_inv29 = 1;
    default: op1_03_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_03_in30 = reg_0344;
    6: op1_03_in30 = reg_0543;
    7: op1_03_in30 = reg_0176;
    8: op1_03_in30 = imem04_in[7:4];
    9: op1_03_in30 = reg_0259;
    97: op1_03_in30 = reg_0259;
    10: op1_03_in30 = reg_0968;
    11: op1_03_in30 = reg_0406;
    12: op1_03_in30 = reg_0065;
    13: op1_03_in30 = reg_0722;
    14: op1_03_in30 = imem03_in[107:104];
    15: op1_03_in30 = reg_0948;
    16: op1_03_in30 = imem07_in[91:88];
    17: op1_03_in30 = reg_0116;
    72: op1_03_in30 = reg_0116;
    18: op1_03_in30 = reg_0153;
    19: op1_03_in30 = imem03_in[31:28];
    79: op1_03_in30 = imem03_in[31:28];
    20: op1_03_in30 = imem05_in[67:64];
    21: op1_03_in30 = reg_0123;
    22: op1_03_in30 = reg_0951;
    23: op1_03_in30 = reg_0801;
    24: op1_03_in30 = imem04_in[39:36];
    25: op1_03_in30 = reg_0423;
    26: op1_03_in30 = reg_0547;
    27: op1_03_in30 = reg_0709;
    28: op1_03_in30 = reg_0905;
    29: op1_03_in30 = reg_0133;
    30: op1_03_in30 = reg_0011;
    31: op1_03_in30 = reg_0230;
    32: op1_03_in30 = reg_0530;
    33: op1_03_in30 = reg_0395;
    92: op1_03_in30 = reg_0395;
    34: op1_03_in30 = reg_0157;
    35: op1_03_in30 = reg_0135;
    36: op1_03_in30 = reg_1020;
    37: op1_03_in30 = reg_0782;
    38: op1_03_in30 = reg_0799;
    39: op1_03_in30 = imem07_in[51:48];
    41: op1_03_in30 = reg_0177;
    42: op1_03_in30 = imem03_in[99:96];
    43: op1_03_in30 = imem05_in[23:20];
    44: op1_03_in30 = reg_0421;
    45: op1_03_in30 = reg_0860;
    46: op1_03_in30 = reg_0374;
    47: op1_03_in30 = reg_0241;
    48: op1_03_in30 = reg_0183;
    49: op1_03_in30 = reg_0733;
    50: op1_03_in30 = reg_0318;
    51: op1_03_in30 = reg_0592;
    52: op1_03_in30 = imem07_in[75:72];
    54: op1_03_in30 = reg_0902;
    55: op1_03_in30 = reg_0656;
    56: op1_03_in30 = imem03_in[59:56];
    57: op1_03_in30 = reg_0809;
    58: op1_03_in30 = reg_0255;
    59: op1_03_in30 = reg_0985;
    60: op1_03_in30 = imem07_in[59:56];
    61: op1_03_in30 = reg_0759;
    62: op1_03_in30 = reg_1010;
    63: op1_03_in30 = reg_1052;
    64: op1_03_in30 = imem02_in[87:84];
    65: op1_03_in30 = reg_0833;
    66: op1_03_in30 = reg_0312;
    67: op1_03_in30 = imem03_in[39:36];
    68: op1_03_in30 = reg_0044;
    70: op1_03_in30 = reg_1053;
    71: op1_03_in30 = reg_0658;
    73: op1_03_in30 = imem03_in[27:24];
    74: op1_03_in30 = reg_0239;
    75: op1_03_in30 = reg_0139;
    76: op1_03_in30 = reg_0428;
    77: op1_03_in30 = reg_0431;
    80: op1_03_in30 = reg_0986;
    81: op1_03_in30 = reg_0136;
    82: op1_03_in30 = reg_0524;
    84: op1_03_in30 = reg_0712;
    85: op1_03_in30 = reg_0767;
    86: op1_03_in30 = reg_0953;
    87: op1_03_in30 = reg_0501;
    88: op1_03_in30 = reg_0227;
    89: op1_03_in30 = reg_0042;
    90: op1_03_in30 = reg_0623;
    91: op1_03_in30 = imem04_in[47:44];
    93: op1_03_in30 = reg_0164;
    94: op1_03_in30 = reg_0325;
    95: op1_03_in30 = reg_0427;
    96: op1_03_in30 = reg_0303;
    default: op1_03_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv30 = 1;
    8: op1_03_inv30 = 1;
    9: op1_03_inv30 = 1;
    13: op1_03_inv30 = 1;
    14: op1_03_inv30 = 1;
    17: op1_03_inv30 = 1;
    18: op1_03_inv30 = 1;
    19: op1_03_inv30 = 1;
    20: op1_03_inv30 = 1;
    21: op1_03_inv30 = 1;
    23: op1_03_inv30 = 1;
    26: op1_03_inv30 = 1;
    27: op1_03_inv30 = 1;
    29: op1_03_inv30 = 1;
    30: op1_03_inv30 = 1;
    31: op1_03_inv30 = 1;
    33: op1_03_inv30 = 1;
    35: op1_03_inv30 = 1;
    38: op1_03_inv30 = 1;
    39: op1_03_inv30 = 1;
    41: op1_03_inv30 = 1;
    43: op1_03_inv30 = 1;
    44: op1_03_inv30 = 1;
    45: op1_03_inv30 = 1;
    48: op1_03_inv30 = 1;
    51: op1_03_inv30 = 1;
    52: op1_03_inv30 = 1;
    55: op1_03_inv30 = 1;
    56: op1_03_inv30 = 1;
    59: op1_03_inv30 = 1;
    60: op1_03_inv30 = 1;
    61: op1_03_inv30 = 1;
    62: op1_03_inv30 = 1;
    64: op1_03_inv30 = 1;
    66: op1_03_inv30 = 1;
    68: op1_03_inv30 = 1;
    70: op1_03_inv30 = 1;
    71: op1_03_inv30 = 1;
    74: op1_03_inv30 = 1;
    75: op1_03_inv30 = 1;
    84: op1_03_inv30 = 1;
    85: op1_03_inv30 = 1;
    89: op1_03_inv30 = 1;
    90: op1_03_inv30 = 1;
    93: op1_03_inv30 = 1;
    95: op1_03_inv30 = 1;
    96: op1_03_inv30 = 1;
    97: op1_03_inv30 = 1;
    default: op1_03_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_03_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_03_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in00 = reg_0401;
    6: op1_04_in00 = reg_0552;
    7: op1_04_in00 = imem00_in[11:8];
    8: op1_04_in00 = imem04_in[15:12];
    9: op1_04_in00 = reg_0256;
    10: op1_04_in00 = reg_0952;
    11: op1_04_in00 = reg_0367;
    4: op1_04_in00 = imem07_in[39:36];
    3: op1_04_in00 = imem07_in[39:36];
    12: op1_04_in00 = reg_0043;
    13: op1_04_in00 = imem00_in[3:0];
    53: op1_04_in00 = imem00_in[3:0];
    14: op1_04_in00 = reg_0598;
    15: op1_04_in00 = reg_0950;
    16: op1_04_in00 = imem00_in[7:4];
    69: op1_04_in00 = imem00_in[7:4];
    17: op1_04_in00 = reg_0119;
    18: op1_04_in00 = imem06_in[27:24];
    19: op1_04_in00 = imem03_in[43:40];
    20: op1_04_in00 = imem05_in[95:92];
    21: op1_04_in00 = reg_0127;
    22: op1_04_in00 = reg_0949;
    23: op1_04_in00 = reg_0017;
    2: op1_04_in00 = imem07_in[35:32];
    24: op1_04_in00 = imem04_in[67:64];
    25: op1_04_in00 = imem00_in[67:64];
    26: op1_04_in00 = reg_0658;
    27: op1_04_in00 = reg_0697;
    28: op1_04_in00 = reg_0226;
    29: op1_04_in00 = reg_0152;
    97: op1_04_in00 = reg_0152;
    30: op1_04_in00 = imem07_in[27:24];
    31: op1_04_in00 = reg_1043;
    32: op1_04_in00 = reg_0778;
    33: op1_04_in00 = reg_0392;
    34: op1_04_in00 = imem00_in[19:16];
    78: op1_04_in00 = imem00_in[19:16];
    35: op1_04_in00 = reg_0133;
    36: op1_04_in00 = reg_0292;
    37: op1_04_in00 = reg_0577;
    38: op1_04_in00 = reg_0372;
    39: op1_04_in00 = imem07_in[75:72];
    40: op1_04_in00 = imem00_in[27:24];
    41: op1_04_in00 = reg_0171;
    42: op1_04_in00 = reg_0394;
    43: op1_04_in00 = imem05_in[39:36];
    44: op1_04_in00 = reg_0047;
    94: op1_04_in00 = reg_0047;
    45: op1_04_in00 = reg_0544;
    46: op1_04_in00 = reg_0979;
    47: op1_04_in00 = reg_0633;
    48: op1_04_in00 = imem00_in[15:12];
    83: op1_04_in00 = imem00_in[15:12];
    49: op1_04_in00 = reg_0065;
    50: op1_04_in00 = reg_0865;
    89: op1_04_in00 = reg_0865;
    51: op1_04_in00 = reg_0503;
    52: op1_04_in00 = reg_0183;
    54: op1_04_in00 = reg_0737;
    55: op1_04_in00 = reg_0082;
    56: op1_04_in00 = imem03_in[71:68];
    57: op1_04_in00 = reg_0288;
    58: op1_04_in00 = reg_0957;
    59: op1_04_in00 = reg_0987;
    60: op1_04_in00 = imem07_in[71:68];
    61: op1_04_in00 = reg_0734;
    62: op1_04_in00 = reg_0399;
    63: op1_04_in00 = reg_0249;
    64: op1_04_in00 = reg_0355;
    65: op1_04_in00 = reg_0376;
    66: op1_04_in00 = reg_0844;
    67: op1_04_in00 = imem03_in[51:48];
    68: op1_04_in00 = reg_0531;
    70: op1_04_in00 = reg_0821;
    71: op1_04_in00 = reg_0495;
    72: op1_04_in00 = reg_0733;
    73: op1_04_in00 = imem03_in[39:36];
    74: op1_04_in00 = reg_1008;
    75: op1_04_in00 = reg_0137;
    76: op1_04_in00 = reg_0532;
    77: op1_04_in00 = reg_0165;
    79: op1_04_in00 = imem03_in[47:44];
    80: op1_04_in00 = reg_0989;
    81: op1_04_in00 = reg_0944;
    82: op1_04_in00 = reg_0076;
    84: op1_04_in00 = reg_0221;
    85: op1_04_in00 = reg_0581;
    86: op1_04_in00 = reg_0314;
    87: op1_04_in00 = reg_0830;
    88: op1_04_in00 = reg_0521;
    90: op1_04_in00 = reg_0238;
    91: op1_04_in00 = imem04_in[51:48];
    92: op1_04_in00 = reg_0048;
    93: op1_04_in00 = reg_0575;
    95: op1_04_in00 = reg_0174;
    96: op1_04_in00 = reg_0250;
    default: op1_04_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv00 = 1;
    6: op1_04_inv00 = 1;
    7: op1_04_inv00 = 1;
    13: op1_04_inv00 = 1;
    15: op1_04_inv00 = 1;
    16: op1_04_inv00 = 1;
    3: op1_04_inv00 = 1;
    18: op1_04_inv00 = 1;
    20: op1_04_inv00 = 1;
    21: op1_04_inv00 = 1;
    23: op1_04_inv00 = 1;
    24: op1_04_inv00 = 1;
    27: op1_04_inv00 = 1;
    32: op1_04_inv00 = 1;
    35: op1_04_inv00 = 1;
    36: op1_04_inv00 = 1;
    37: op1_04_inv00 = 1;
    38: op1_04_inv00 = 1;
    39: op1_04_inv00 = 1;
    40: op1_04_inv00 = 1;
    42: op1_04_inv00 = 1;
    44: op1_04_inv00 = 1;
    49: op1_04_inv00 = 1;
    52: op1_04_inv00 = 1;
    55: op1_04_inv00 = 1;
    56: op1_04_inv00 = 1;
    57: op1_04_inv00 = 1;
    58: op1_04_inv00 = 1;
    62: op1_04_inv00 = 1;
    63: op1_04_inv00 = 1;
    64: op1_04_inv00 = 1;
    67: op1_04_inv00 = 1;
    68: op1_04_inv00 = 1;
    73: op1_04_inv00 = 1;
    74: op1_04_inv00 = 1;
    75: op1_04_inv00 = 1;
    76: op1_04_inv00 = 1;
    77: op1_04_inv00 = 1;
    80: op1_04_inv00 = 1;
    83: op1_04_inv00 = 1;
    85: op1_04_inv00 = 1;
    87: op1_04_inv00 = 1;
    89: op1_04_inv00 = 1;
    93: op1_04_inv00 = 1;
    94: op1_04_inv00 = 1;
    95: op1_04_inv00 = 1;
    96: op1_04_inv00 = 1;
    default: op1_04_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in01 = reg_0028;
    6: op1_04_in01 = reg_0532;
    7: op1_04_in01 = imem00_in[39:36];
    8: op1_04_in01 = imem04_in[19:16];
    9: op1_04_in01 = reg_0243;
    10: op1_04_in01 = reg_0961;
    11: op1_04_in01 = reg_0799;
    4: op1_04_in01 = imem07_in[51:48];
    2: op1_04_in01 = imem07_in[51:48];
    12: op1_04_in01 = reg_0044;
    13: op1_04_in01 = imem00_in[27:24];
    83: op1_04_in01 = imem00_in[27:24];
    14: op1_04_in01 = reg_0572;
    73: op1_04_in01 = reg_0572;
    15: op1_04_in01 = reg_0835;
    16: op1_04_in01 = imem00_in[23:20];
    17: op1_04_in01 = reg_0108;
    3: op1_04_in01 = imem07_in[63:60];
    18: op1_04_in01 = imem06_in[35:32];
    19: op1_04_in01 = imem03_in[51:48];
    20: op1_04_in01 = imem05_in[103:100];
    21: op1_04_in01 = reg_0121;
    22: op1_04_in01 = reg_0960;
    23: op1_04_in01 = reg_0753;
    24: op1_04_in01 = imem04_in[83:80];
    25: op1_04_in01 = imem00_in[83:80];
    26: op1_04_in01 = reg_0666;
    27: op1_04_in01 = reg_0683;
    28: op1_04_in01 = reg_1031;
    29: op1_04_in01 = reg_0146;
    30: op1_04_in01 = imem07_in[75:72];
    31: op1_04_in01 = reg_0104;
    32: op1_04_in01 = reg_1016;
    33: op1_04_in01 = reg_0391;
    34: op1_04_in01 = imem00_in[47:44];
    35: op1_04_in01 = reg_0151;
    36: op1_04_in01 = reg_0540;
    92: op1_04_in01 = reg_0540;
    37: op1_04_in01 = reg_0735;
    38: op1_04_in01 = reg_0034;
    39: op1_04_in01 = reg_0720;
    40: op1_04_in01 = imem00_in[43:40];
    42: op1_04_in01 = reg_0327;
    43: op1_04_in01 = imem05_in[47:44];
    44: op1_04_in01 = reg_0321;
    45: op1_04_in01 = reg_0811;
    46: op1_04_in01 = reg_0974;
    47: op1_04_in01 = reg_0005;
    48: op1_04_in01 = imem00_in[19:16];
    53: op1_04_in01 = imem00_in[19:16];
    69: op1_04_in01 = imem00_in[19:16];
    49: op1_04_in01 = reg_0877;
    50: op1_04_in01 = reg_0857;
    51: op1_04_in01 = reg_0253;
    52: op1_04_in01 = reg_0177;
    54: op1_04_in01 = reg_0354;
    55: op1_04_in01 = reg_0323;
    56: op1_04_in01 = imem03_in[119:116];
    57: op1_04_in01 = reg_0061;
    58: op1_04_in01 = reg_0221;
    59: op1_04_in01 = reg_1002;
    60: op1_04_in01 = reg_0708;
    61: op1_04_in01 = reg_0864;
    62: op1_04_in01 = imem07_in[11:8];
    63: op1_04_in01 = reg_0829;
    64: op1_04_in01 = reg_0341;
    65: op1_04_in01 = reg_0820;
    66: op1_04_in01 = reg_0995;
    67: op1_04_in01 = imem03_in[75:72];
    79: op1_04_in01 = imem03_in[75:72];
    68: op1_04_in01 = reg_0215;
    70: op1_04_in01 = imem02_in[55:52];
    71: op1_04_in01 = reg_0824;
    72: op1_04_in01 = reg_0115;
    74: op1_04_in01 = reg_0376;
    75: op1_04_in01 = reg_0057;
    76: op1_04_in01 = reg_0420;
    77: op1_04_in01 = reg_0167;
    78: op1_04_in01 = imem00_in[99:96];
    80: op1_04_in01 = reg_0977;
    81: op1_04_in01 = reg_0217;
    82: op1_04_in01 = reg_0302;
    84: op1_04_in01 = reg_0710;
    85: op1_04_in01 = reg_0385;
    86: op1_04_in01 = reg_0154;
    87: op1_04_in01 = reg_0500;
    88: op1_04_in01 = reg_0610;
    89: op1_04_in01 = reg_0622;
    90: op1_04_in01 = reg_0278;
    91: op1_04_in01 = imem04_in[67:64];
    93: op1_04_in01 = reg_0641;
    94: op1_04_in01 = reg_0428;
    95: op1_04_in01 = reg_0175;
    96: op1_04_in01 = reg_0325;
    97: op1_04_in01 = reg_0023;
    default: op1_04_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv01 = 1;
    8: op1_04_inv01 = 1;
    11: op1_04_inv01 = 1;
    12: op1_04_inv01 = 1;
    13: op1_04_inv01 = 1;
    14: op1_04_inv01 = 1;
    18: op1_04_inv01 = 1;
    22: op1_04_inv01 = 1;
    2: op1_04_inv01 = 1;
    25: op1_04_inv01 = 1;
    26: op1_04_inv01 = 1;
    27: op1_04_inv01 = 1;
    28: op1_04_inv01 = 1;
    29: op1_04_inv01 = 1;
    30: op1_04_inv01 = 1;
    34: op1_04_inv01 = 1;
    35: op1_04_inv01 = 1;
    36: op1_04_inv01 = 1;
    37: op1_04_inv01 = 1;
    38: op1_04_inv01 = 1;
    42: op1_04_inv01 = 1;
    45: op1_04_inv01 = 1;
    46: op1_04_inv01 = 1;
    47: op1_04_inv01 = 1;
    49: op1_04_inv01 = 1;
    53: op1_04_inv01 = 1;
    54: op1_04_inv01 = 1;
    55: op1_04_inv01 = 1;
    57: op1_04_inv01 = 1;
    58: op1_04_inv01 = 1;
    60: op1_04_inv01 = 1;
    61: op1_04_inv01 = 1;
    62: op1_04_inv01 = 1;
    63: op1_04_inv01 = 1;
    64: op1_04_inv01 = 1;
    67: op1_04_inv01 = 1;
    70: op1_04_inv01 = 1;
    71: op1_04_inv01 = 1;
    73: op1_04_inv01 = 1;
    76: op1_04_inv01 = 1;
    77: op1_04_inv01 = 1;
    78: op1_04_inv01 = 1;
    81: op1_04_inv01 = 1;
    82: op1_04_inv01 = 1;
    84: op1_04_inv01 = 1;
    85: op1_04_inv01 = 1;
    86: op1_04_inv01 = 1;
    90: op1_04_inv01 = 1;
    91: op1_04_inv01 = 1;
    92: op1_04_inv01 = 1;
    93: op1_04_inv01 = 1;
    default: op1_04_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in02 = reg_0025;
    6: op1_04_in02 = reg_0301;
    7: op1_04_in02 = imem00_in[55:52];
    16: op1_04_in02 = imem00_in[55:52];
    53: op1_04_in02 = imem00_in[55:52];
    8: op1_04_in02 = imem04_in[59:56];
    9: op1_04_in02 = reg_0253;
    10: op1_04_in02 = reg_0943;
    11: op1_04_in02 = reg_0787;
    4: op1_04_in02 = imem07_in[75:72];
    12: op1_04_in02 = reg_1020;
    13: op1_04_in02 = imem00_in[75:72];
    14: op1_04_in02 = reg_0587;
    15: op1_04_in02 = reg_0024;
    17: op1_04_in02 = imem02_in[3:0];
    3: op1_04_in02 = imem07_in[95:92];
    18: op1_04_in02 = reg_0610;
    19: op1_04_in02 = imem03_in[59:56];
    20: op1_04_in02 = imem05_in[115:112];
    21: op1_04_in02 = reg_0768;
    22: op1_04_in02 = reg_0215;
    23: op1_04_in02 = reg_1010;
    2: op1_04_in02 = imem07_in[59:56];
    24: op1_04_in02 = imem04_in[103:100];
    25: op1_04_in02 = imem00_in[87:84];
    26: op1_04_in02 = reg_0655;
    27: op1_04_in02 = reg_0698;
    28: op1_04_in02 = reg_1045;
    29: op1_04_in02 = reg_0156;
    30: op1_04_in02 = imem07_in[99:96];
    31: op1_04_in02 = reg_0119;
    32: op1_04_in02 = reg_0760;
    33: op1_04_in02 = reg_0804;
    34: op1_04_in02 = imem00_in[91:88];
    35: op1_04_in02 = reg_0128;
    81: op1_04_in02 = reg_0128;
    36: op1_04_in02 = reg_0888;
    37: op1_04_in02 = reg_0534;
    38: op1_04_in02 = reg_0593;
    39: op1_04_in02 = reg_0730;
    40: op1_04_in02 = imem00_in[59:56];
    48: op1_04_in02 = imem00_in[59:56];
    42: op1_04_in02 = reg_0346;
    43: op1_04_in02 = imem05_in[55:52];
    44: op1_04_in02 = reg_0599;
    94: op1_04_in02 = reg_0599;
    45: op1_04_in02 = reg_0227;
    63: op1_04_in02 = reg_0227;
    46: op1_04_in02 = reg_0975;
    47: op1_04_in02 = imem07_in[7:4];
    49: op1_04_in02 = reg_0364;
    50: op1_04_in02 = reg_0335;
    51: op1_04_in02 = reg_0869;
    52: op1_04_in02 = reg_0168;
    54: op1_04_in02 = reg_0740;
    55: op1_04_in02 = reg_0358;
    56: op1_04_in02 = imem03_in[123:120];
    57: op1_04_in02 = reg_0078;
    58: op1_04_in02 = reg_0235;
    59: op1_04_in02 = reg_0979;
    66: op1_04_in02 = reg_0979;
    60: op1_04_in02 = reg_0709;
    61: op1_04_in02 = reg_0691;
    62: op1_04_in02 = imem07_in[67:64];
    64: op1_04_in02 = reg_0290;
    65: op1_04_in02 = reg_0246;
    67: op1_04_in02 = imem03_in[83:80];
    68: op1_04_in02 = reg_0581;
    69: op1_04_in02 = imem00_in[31:28];
    70: op1_04_in02 = imem02_in[99:96];
    71: op1_04_in02 = imem05_in[11:8];
    72: op1_04_in02 = reg_0110;
    73: op1_04_in02 = reg_0580;
    74: op1_04_in02 = reg_0820;
    75: op1_04_in02 = reg_0963;
    76: op1_04_in02 = reg_0427;
    77: op1_04_in02 = reg_0163;
    78: op1_04_in02 = imem00_in[127:124];
    79: op1_04_in02 = imem03_in[103:100];
    80: op1_04_in02 = reg_0990;
    82: op1_04_in02 = reg_0584;
    83: op1_04_in02 = imem00_in[47:44];
    84: op1_04_in02 = reg_0721;
    85: op1_04_in02 = reg_0551;
    86: op1_04_in02 = reg_1046;
    87: op1_04_in02 = reg_0216;
    88: op1_04_in02 = reg_0925;
    89: op1_04_in02 = reg_0660;
    90: op1_04_in02 = reg_0230;
    91: op1_04_in02 = imem04_in[91:88];
    92: op1_04_in02 = reg_0058;
    93: op1_04_in02 = reg_0353;
    95: op1_04_in02 = reg_0429;
    96: op1_04_in02 = reg_0315;
    97: op1_04_in02 = reg_0892;
    default: op1_04_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_04_inv02 = 1;
    4: op1_04_inv02 = 1;
    17: op1_04_inv02 = 1;
    3: op1_04_inv02 = 1;
    18: op1_04_inv02 = 1;
    21: op1_04_inv02 = 1;
    22: op1_04_inv02 = 1;
    23: op1_04_inv02 = 1;
    24: op1_04_inv02 = 1;
    28: op1_04_inv02 = 1;
    29: op1_04_inv02 = 1;
    33: op1_04_inv02 = 1;
    36: op1_04_inv02 = 1;
    43: op1_04_inv02 = 1;
    44: op1_04_inv02 = 1;
    46: op1_04_inv02 = 1;
    47: op1_04_inv02 = 1;
    48: op1_04_inv02 = 1;
    51: op1_04_inv02 = 1;
    52: op1_04_inv02 = 1;
    56: op1_04_inv02 = 1;
    59: op1_04_inv02 = 1;
    60: op1_04_inv02 = 1;
    61: op1_04_inv02 = 1;
    62: op1_04_inv02 = 1;
    65: op1_04_inv02 = 1;
    66: op1_04_inv02 = 1;
    67: op1_04_inv02 = 1;
    69: op1_04_inv02 = 1;
    70: op1_04_inv02 = 1;
    71: op1_04_inv02 = 1;
    73: op1_04_inv02 = 1;
    79: op1_04_inv02 = 1;
    80: op1_04_inv02 = 1;
    81: op1_04_inv02 = 1;
    84: op1_04_inv02 = 1;
    86: op1_04_inv02 = 1;
    87: op1_04_inv02 = 1;
    89: op1_04_inv02 = 1;
    91: op1_04_inv02 = 1;
    93: op1_04_inv02 = 1;
    94: op1_04_inv02 = 1;
    97: op1_04_inv02 = 1;
    default: op1_04_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in03 = reg_0029;
    6: op1_04_in03 = reg_0291;
    7: op1_04_in03 = imem00_in[71:68];
    8: op1_04_in03 = imem04_in[79:76];
    9: op1_04_in03 = reg_0147;
    10: op1_04_in03 = reg_0953;
    11: op1_04_in03 = reg_0026;
    4: op1_04_in03 = imem07_in[127:124];
    12: op1_04_in03 = reg_0491;
    13: op1_04_in03 = imem00_in[79:76];
    14: op1_04_in03 = reg_0319;
    81: op1_04_in03 = reg_0319;
    15: op1_04_in03 = reg_0255;
    16: op1_04_in03 = imem00_in[63:60];
    53: op1_04_in03 = imem00_in[63:60];
    17: op1_04_in03 = imem02_in[47:44];
    3: op1_04_in03 = imem07_in[123:120];
    18: op1_04_in03 = reg_0626;
    19: op1_04_in03 = imem03_in[63:60];
    20: op1_04_in03 = imem05_in[123:120];
    43: op1_04_in03 = imem05_in[123:120];
    21: op1_04_in03 = reg_0743;
    22: op1_04_in03 = reg_0826;
    58: op1_04_in03 = reg_0826;
    23: op1_04_in03 = imem07_in[3:0];
    24: op1_04_in03 = imem04_in[111:108];
    25: op1_04_in03 = reg_0693;
    48: op1_04_in03 = reg_0693;
    26: op1_04_in03 = reg_0653;
    27: op1_04_in03 = reg_0686;
    28: op1_04_in03 = reg_1034;
    29: op1_04_in03 = reg_0372;
    30: op1_04_in03 = reg_0720;
    31: op1_04_in03 = reg_0120;
    32: op1_04_in03 = reg_0069;
    33: op1_04_in03 = reg_0388;
    34: op1_04_in03 = reg_0677;
    35: op1_04_in03 = reg_0138;
    36: op1_04_in03 = reg_0931;
    37: op1_04_in03 = reg_0542;
    38: op1_04_in03 = reg_0897;
    39: op1_04_in03 = reg_0702;
    40: op1_04_in03 = imem00_in[87:84];
    42: op1_04_in03 = reg_0793;
    44: op1_04_in03 = reg_0502;
    76: op1_04_in03 = reg_0502;
    45: op1_04_in03 = reg_0616;
    46: op1_04_in03 = reg_0988;
    47: op1_04_in03 = imem07_in[19:16];
    49: op1_04_in03 = reg_0547;
    50: op1_04_in03 = reg_0772;
    51: op1_04_in03 = reg_0500;
    52: op1_04_in03 = reg_0173;
    54: op1_04_in03 = reg_0925;
    55: op1_04_in03 = reg_0664;
    56: op1_04_in03 = reg_0099;
    57: op1_04_in03 = reg_0899;
    59: op1_04_in03 = reg_0993;
    60: op1_04_in03 = reg_0705;
    61: op1_04_in03 = reg_0351;
    62: op1_04_in03 = reg_0703;
    63: op1_04_in03 = reg_0737;
    64: op1_04_in03 = reg_0894;
    65: op1_04_in03 = reg_0234;
    66: op1_04_in03 = reg_1001;
    67: op1_04_in03 = imem03_in[99:96];
    68: op1_04_in03 = reg_0128;
    69: op1_04_in03 = imem00_in[59:56];
    70: op1_04_in03 = reg_0810;
    71: op1_04_in03 = imem05_in[51:48];
    72: op1_04_in03 = reg_0063;
    73: op1_04_in03 = reg_0445;
    74: op1_04_in03 = reg_0581;
    75: op1_04_in03 = reg_0941;
    77: op1_04_in03 = reg_0185;
    78: op1_04_in03 = reg_0001;
    79: op1_04_in03 = reg_0060;
    80: op1_04_in03 = reg_0997;
    82: op1_04_in03 = reg_0072;
    83: op1_04_in03 = imem00_in[83:80];
    84: op1_04_in03 = reg_0718;
    85: op1_04_in03 = reg_0987;
    86: op1_04_in03 = reg_0952;
    87: op1_04_in03 = reg_0902;
    88: op1_04_in03 = reg_0116;
    89: op1_04_in03 = reg_0625;
    90: op1_04_in03 = reg_0820;
    91: op1_04_in03 = reg_0913;
    92: op1_04_in03 = reg_0066;
    93: op1_04_in03 = reg_0599;
    94: op1_04_in03 = reg_0350;
    95: op1_04_in03 = reg_0161;
    96: op1_04_in03 = reg_0419;
    97: op1_04_in03 = reg_0330;
    default: op1_04_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv03 = 1;
    6: op1_04_inv03 = 1;
    9: op1_04_inv03 = 1;
    10: op1_04_inv03 = 1;
    11: op1_04_inv03 = 1;
    12: op1_04_inv03 = 1;
    15: op1_04_inv03 = 1;
    17: op1_04_inv03 = 1;
    3: op1_04_inv03 = 1;
    21: op1_04_inv03 = 1;
    23: op1_04_inv03 = 1;
    25: op1_04_inv03 = 1;
    26: op1_04_inv03 = 1;
    27: op1_04_inv03 = 1;
    28: op1_04_inv03 = 1;
    29: op1_04_inv03 = 1;
    30: op1_04_inv03 = 1;
    33: op1_04_inv03 = 1;
    34: op1_04_inv03 = 1;
    38: op1_04_inv03 = 1;
    39: op1_04_inv03 = 1;
    40: op1_04_inv03 = 1;
    45: op1_04_inv03 = 1;
    48: op1_04_inv03 = 1;
    49: op1_04_inv03 = 1;
    50: op1_04_inv03 = 1;
    51: op1_04_inv03 = 1;
    54: op1_04_inv03 = 1;
    57: op1_04_inv03 = 1;
    58: op1_04_inv03 = 1;
    60: op1_04_inv03 = 1;
    62: op1_04_inv03 = 1;
    63: op1_04_inv03 = 1;
    64: op1_04_inv03 = 1;
    65: op1_04_inv03 = 1;
    66: op1_04_inv03 = 1;
    67: op1_04_inv03 = 1;
    74: op1_04_inv03 = 1;
    75: op1_04_inv03 = 1;
    78: op1_04_inv03 = 1;
    79: op1_04_inv03 = 1;
    81: op1_04_inv03 = 1;
    82: op1_04_inv03 = 1;
    84: op1_04_inv03 = 1;
    85: op1_04_inv03 = 1;
    87: op1_04_inv03 = 1;
    88: op1_04_inv03 = 1;
    91: op1_04_inv03 = 1;
    93: op1_04_inv03 = 1;
    94: op1_04_inv03 = 1;
    95: op1_04_inv03 = 1;
    96: op1_04_inv03 = 1;
    97: op1_04_inv03 = 1;
    default: op1_04_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in04 = reg_0005;
    6: op1_04_in04 = reg_0053;
    7: op1_04_in04 = imem00_in[83:80];
    8: op1_04_in04 = imem04_in[127:124];
    9: op1_04_in04 = reg_0136;
    10: op1_04_in04 = reg_0268;
    11: op1_04_in04 = reg_1010;
    4: op1_04_in04 = reg_0430;
    12: op1_04_in04 = reg_0489;
    13: op1_04_in04 = imem00_in[123:120];
    14: op1_04_in04 = reg_0982;
    15: op1_04_in04 = reg_0819;
    86: op1_04_in04 = reg_0819;
    16: op1_04_in04 = imem00_in[71:68];
    17: op1_04_in04 = imem02_in[95:92];
    3: op1_04_in04 = reg_0172;
    18: op1_04_in04 = reg_0632;
    19: op1_04_in04 = imem03_in[79:76];
    20: op1_04_in04 = reg_0133;
    21: op1_04_in04 = reg_0917;
    22: op1_04_in04 = reg_0229;
    23: op1_04_in04 = imem07_in[7:4];
    24: op1_04_in04 = imem04_in[119:116];
    25: op1_04_in04 = reg_0697;
    48: op1_04_in04 = reg_0697;
    26: op1_04_in04 = reg_0640;
    27: op1_04_in04 = reg_0680;
    28: op1_04_in04 = reg_0120;
    29: op1_04_in04 = reg_0317;
    30: op1_04_in04 = reg_0726;
    31: op1_04_in04 = reg_0112;
    32: op1_04_in04 = reg_0074;
    33: op1_04_in04 = reg_0222;
    34: op1_04_in04 = reg_0191;
    35: op1_04_in04 = reg_0153;
    36: op1_04_in04 = reg_0061;
    37: op1_04_in04 = reg_0407;
    38: op1_04_in04 = reg_0566;
    39: op1_04_in04 = reg_0708;
    40: op1_04_in04 = imem00_in[119:116];
    42: op1_04_in04 = reg_0038;
    43: op1_04_in04 = reg_0963;
    44: op1_04_in04 = reg_0868;
    45: op1_04_in04 = reg_0906;
    46: op1_04_in04 = reg_0976;
    47: op1_04_in04 = imem07_in[75:72];
    49: op1_04_in04 = reg_1003;
    50: op1_04_in04 = reg_0761;
    51: op1_04_in04 = reg_0216;
    53: op1_04_in04 = imem00_in[107:104];
    54: op1_04_in04 = reg_0769;
    55: op1_04_in04 = reg_0818;
    56: op1_04_in04 = reg_0580;
    57: op1_04_in04 = reg_0027;
    58: op1_04_in04 = reg_0022;
    59: op1_04_in04 = reg_0999;
    60: op1_04_in04 = reg_0707;
    61: op1_04_in04 = reg_0025;
    62: op1_04_in04 = reg_0805;
    63: op1_04_in04 = reg_0615;
    64: op1_04_in04 = reg_0643;
    65: op1_04_in04 = reg_0987;
    66: op1_04_in04 = reg_0990;
    67: op1_04_in04 = imem03_in[123:120];
    68: op1_04_in04 = reg_0813;
    69: op1_04_in04 = reg_0001;
    70: op1_04_in04 = reg_0666;
    71: op1_04_in04 = imem05_in[75:72];
    72: op1_04_in04 = reg_0365;
    73: op1_04_in04 = reg_0307;
    74: op1_04_in04 = reg_0266;
    75: op1_04_in04 = reg_0940;
    76: op1_04_in04 = reg_0175;
    77: op1_04_in04 = reg_0173;
    78: op1_04_in04 = reg_0519;
    79: op1_04_in04 = reg_0535;
    80: op1_04_in04 = imem04_in[3:0];
    81: op1_04_in04 = reg_0138;
    82: op1_04_in04 = reg_0288;
    83: op1_04_in04 = imem00_in[91:88];
    84: op1_04_in04 = reg_0563;
    85: op1_04_in04 = reg_1002;
    87: op1_04_in04 = reg_0610;
    88: op1_04_in04 = reg_0273;
    89: op1_04_in04 = reg_0344;
    90: op1_04_in04 = reg_0581;
    91: op1_04_in04 = reg_0540;
    92: op1_04_in04 = reg_0056;
    93: op1_04_in04 = reg_0427;
    94: op1_04_in04 = reg_0429;
    95: op1_04_in04 = reg_0447;
    96: op1_04_in04 = reg_0339;
    97: op1_04_in04 = reg_0530;
    default: op1_04_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv04 = 1;
    6: op1_04_inv04 = 1;
    11: op1_04_inv04 = 1;
    15: op1_04_inv04 = 1;
    16: op1_04_inv04 = 1;
    3: op1_04_inv04 = 1;
    22: op1_04_inv04 = 1;
    27: op1_04_inv04 = 1;
    29: op1_04_inv04 = 1;
    31: op1_04_inv04 = 1;
    33: op1_04_inv04 = 1;
    34: op1_04_inv04 = 1;
    35: op1_04_inv04 = 1;
    36: op1_04_inv04 = 1;
    37: op1_04_inv04 = 1;
    40: op1_04_inv04 = 1;
    43: op1_04_inv04 = 1;
    45: op1_04_inv04 = 1;
    55: op1_04_inv04 = 1;
    59: op1_04_inv04 = 1;
    61: op1_04_inv04 = 1;
    63: op1_04_inv04 = 1;
    64: op1_04_inv04 = 1;
    65: op1_04_inv04 = 1;
    66: op1_04_inv04 = 1;
    68: op1_04_inv04 = 1;
    72: op1_04_inv04 = 1;
    73: op1_04_inv04 = 1;
    74: op1_04_inv04 = 1;
    75: op1_04_inv04 = 1;
    79: op1_04_inv04 = 1;
    80: op1_04_inv04 = 1;
    81: op1_04_inv04 = 1;
    82: op1_04_inv04 = 1;
    84: op1_04_inv04 = 1;
    86: op1_04_inv04 = 1;
    87: op1_04_inv04 = 1;
    93: op1_04_inv04 = 1;
    default: op1_04_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in05 = imem07_in[7:4];
    6: op1_04_in05 = reg_0071;
    7: op1_04_in05 = imem00_in[107:104];
    8: op1_04_in05 = reg_0530;
    9: op1_04_in05 = reg_0133;
    10: op1_04_in05 = reg_0259;
    24: op1_04_in05 = reg_0259;
    11: op1_04_in05 = reg_0803;
    4: op1_04_in05 = reg_0436;
    12: op1_04_in05 = reg_0959;
    13: op1_04_in05 = reg_0681;
    67: op1_04_in05 = reg_0681;
    14: op1_04_in05 = reg_0992;
    15: op1_04_in05 = reg_0150;
    16: op1_04_in05 = imem00_in[79:76];
    17: op1_04_in05 = imem02_in[111:108];
    3: op1_04_in05 = reg_0169;
    18: op1_04_in05 = reg_0622;
    19: op1_04_in05 = reg_0583;
    20: op1_04_in05 = reg_0142;
    21: op1_04_in05 = reg_0887;
    22: op1_04_in05 = reg_0785;
    23: op1_04_in05 = imem07_in[35:32];
    25: op1_04_in05 = reg_0696;
    26: op1_04_in05 = reg_0636;
    64: op1_04_in05 = reg_0636;
    27: op1_04_in05 = reg_0687;
    28: op1_04_in05 = reg_0108;
    29: op1_04_in05 = reg_0036;
    30: op1_04_in05 = reg_0705;
    31: op1_04_in05 = imem02_in[7:4];
    32: op1_04_in05 = reg_0525;
    33: op1_04_in05 = reg_0380;
    34: op1_04_in05 = reg_0188;
    35: op1_04_in05 = imem06_in[15:12];
    36: op1_04_in05 = reg_0078;
    37: op1_04_in05 = reg_0558;
    38: op1_04_in05 = reg_0381;
    39: op1_04_in05 = reg_0709;
    40: op1_04_in05 = imem00_in[123:120];
    42: op1_04_in05 = reg_0795;
    43: op1_04_in05 = reg_0951;
    44: op1_04_in05 = reg_0175;
    93: op1_04_in05 = reg_0175;
    45: op1_04_in05 = reg_0123;
    46: op1_04_in05 = reg_0065;
    47: op1_04_in05 = imem07_in[119:116];
    48: op1_04_in05 = reg_0689;
    53: op1_04_in05 = reg_0689;
    49: op1_04_in05 = reg_1005;
    50: op1_04_in05 = reg_0049;
    51: op1_04_in05 = reg_0616;
    54: op1_04_in05 = reg_0733;
    55: op1_04_in05 = reg_0087;
    56: op1_04_in05 = reg_0046;
    57: op1_04_in05 = imem05_in[19:16];
    58: op1_04_in05 = reg_0094;
    59: op1_04_in05 = reg_0997;
    60: op1_04_in05 = reg_0047;
    61: op1_04_in05 = reg_0021;
    62: op1_04_in05 = reg_0421;
    63: op1_04_in05 = reg_1053;
    65: op1_04_in05 = reg_1002;
    66: op1_04_in05 = reg_1000;
    68: op1_04_in05 = reg_0510;
    69: op1_04_in05 = reg_0682;
    70: op1_04_in05 = reg_0647;
    71: op1_04_in05 = imem05_in[91:88];
    72: op1_04_in05 = reg_0642;
    73: op1_04_in05 = reg_0577;
    74: op1_04_in05 = reg_0994;
    75: op1_04_in05 = reg_0935;
    76: op1_04_in05 = reg_0172;
    78: op1_04_in05 = reg_0825;
    79: op1_04_in05 = reg_0760;
    80: op1_04_in05 = imem04_in[27:24];
    81: op1_04_in05 = reg_0448;
    82: op1_04_in05 = reg_0494;
    83: op1_04_in05 = imem00_in[119:116];
    84: op1_04_in05 = reg_0299;
    85: op1_04_in05 = reg_0991;
    86: op1_04_in05 = reg_0970;
    87: op1_04_in05 = reg_1017;
    88: op1_04_in05 = reg_0114;
    89: op1_04_in05 = reg_0294;
    90: op1_04_in05 = reg_0233;
    91: op1_04_in05 = reg_0008;
    92: op1_04_in05 = reg_0302;
    94: op1_04_in05 = reg_0703;
    95: op1_04_in05 = reg_0339;
    96: op1_04_in05 = reg_0529;
    97: op1_04_in05 = reg_0806;
    default: op1_04_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv05 = 1;
    8: op1_04_inv05 = 1;
    15: op1_04_inv05 = 1;
    16: op1_04_inv05 = 1;
    17: op1_04_inv05 = 1;
    3: op1_04_inv05 = 1;
    18: op1_04_inv05 = 1;
    20: op1_04_inv05 = 1;
    21: op1_04_inv05 = 1;
    23: op1_04_inv05 = 1;
    26: op1_04_inv05 = 1;
    27: op1_04_inv05 = 1;
    28: op1_04_inv05 = 1;
    33: op1_04_inv05 = 1;
    34: op1_04_inv05 = 1;
    35: op1_04_inv05 = 1;
    45: op1_04_inv05 = 1;
    47: op1_04_inv05 = 1;
    48: op1_04_inv05 = 1;
    50: op1_04_inv05 = 1;
    51: op1_04_inv05 = 1;
    53: op1_04_inv05 = 1;
    54: op1_04_inv05 = 1;
    55: op1_04_inv05 = 1;
    57: op1_04_inv05 = 1;
    59: op1_04_inv05 = 1;
    60: op1_04_inv05 = 1;
    61: op1_04_inv05 = 1;
    62: op1_04_inv05 = 1;
    63: op1_04_inv05 = 1;
    64: op1_04_inv05 = 1;
    65: op1_04_inv05 = 1;
    68: op1_04_inv05 = 1;
    69: op1_04_inv05 = 1;
    71: op1_04_inv05 = 1;
    72: op1_04_inv05 = 1;
    73: op1_04_inv05 = 1;
    75: op1_04_inv05 = 1;
    79: op1_04_inv05 = 1;
    80: op1_04_inv05 = 1;
    83: op1_04_inv05 = 1;
    84: op1_04_inv05 = 1;
    85: op1_04_inv05 = 1;
    86: op1_04_inv05 = 1;
    88: op1_04_inv05 = 1;
    96: op1_04_inv05 = 1;
    default: op1_04_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in06 = imem07_in[31:28];
    6: op1_04_in06 = reg_0070;
    7: op1_04_in06 = reg_0695;
    8: op1_04_in06 = reg_0553;
    9: op1_04_in06 = reg_0139;
    10: op1_04_in06 = reg_0273;
    11: op1_04_in06 = reg_0782;
    4: op1_04_in06 = reg_0442;
    12: op1_04_in06 = reg_0967;
    13: op1_04_in06 = reg_0685;
    14: op1_04_in06 = reg_0984;
    15: op1_04_in06 = reg_0142;
    16: op1_04_in06 = imem00_in[91:88];
    17: op1_04_in06 = imem02_in[115:112];
    3: op1_04_in06 = reg_0157;
    18: op1_04_in06 = reg_0348;
    19: op1_04_in06 = reg_0587;
    20: op1_04_in06 = reg_0156;
    21: op1_04_in06 = reg_0650;
    22: op1_04_in06 = reg_0244;
    23: op1_04_in06 = imem07_in[59:56];
    24: op1_04_in06 = reg_0014;
    25: op1_04_in06 = reg_0689;
    26: op1_04_in06 = reg_0667;
    27: op1_04_in06 = reg_0453;
    28: op1_04_in06 = reg_0101;
    29: op1_04_in06 = reg_0557;
    30: op1_04_in06 = reg_0707;
    31: op1_04_in06 = imem02_in[35:32];
    32: op1_04_in06 = reg_0279;
    33: op1_04_in06 = reg_0486;
    86: op1_04_in06 = reg_0486;
    34: op1_04_in06 = reg_0203;
    35: op1_04_in06 = imem06_in[51:48];
    36: op1_04_in06 = reg_0074;
    37: op1_04_in06 = reg_0556;
    38: op1_04_in06 = reg_0294;
    39: op1_04_in06 = reg_0705;
    40: op1_04_in06 = reg_0679;
    42: op1_04_in06 = reg_0784;
    43: op1_04_in06 = reg_0821;
    44: op1_04_in06 = reg_0180;
    45: op1_04_in06 = reg_0118;
    46: op1_04_in06 = reg_0542;
    82: op1_04_in06 = reg_0542;
    47: op1_04_in06 = reg_0722;
    48: op1_04_in06 = reg_0684;
    53: op1_04_in06 = reg_0684;
    49: op1_04_in06 = reg_0584;
    92: op1_04_in06 = reg_0584;
    50: op1_04_in06 = imem03_in[3:0];
    51: op1_04_in06 = reg_0610;
    54: op1_04_in06 = reg_0827;
    88: op1_04_in06 = reg_0827;
    55: op1_04_in06 = reg_0347;
    56: op1_04_in06 = reg_0547;
    57: op1_04_in06 = imem05_in[67:64];
    58: op1_04_in06 = reg_0489;
    59: op1_04_in06 = reg_0126;
    60: op1_04_in06 = reg_0321;
    61: op1_04_in06 = reg_0926;
    62: op1_04_in06 = reg_0350;
    63: op1_04_in06 = reg_0860;
    64: op1_04_in06 = reg_0855;
    65: op1_04_in06 = imem04_in[11:8];
    66: op1_04_in06 = imem04_in[7:4];
    67: op1_04_in06 = reg_1007;
    68: op1_04_in06 = reg_0579;
    69: op1_04_in06 = reg_0519;
    70: op1_04_in06 = reg_0643;
    71: op1_04_in06 = imem05_in[95:92];
    72: op1_04_in06 = reg_0558;
    73: op1_04_in06 = reg_0434;
    74: op1_04_in06 = imem04_in[99:96];
    75: op1_04_in06 = reg_0819;
    76: op1_04_in06 = reg_0161;
    78: op1_04_in06 = reg_0883;
    79: op1_04_in06 = reg_0322;
    80: op1_04_in06 = imem04_in[43:40];
    81: op1_04_in06 = reg_0013;
    83: op1_04_in06 = reg_0768;
    84: op1_04_in06 = reg_0250;
    85: op1_04_in06 = reg_0979;
    87: op1_04_in06 = reg_0769;
    89: op1_04_in06 = reg_0267;
    90: op1_04_in06 = reg_0551;
    91: op1_04_in06 = reg_0123;
    93: op1_04_in06 = reg_0179;
    94: op1_04_in06 = reg_0185;
    97: op1_04_in06 = reg_0951;
    default: op1_04_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv06 = 1;
    7: op1_04_inv06 = 1;
    10: op1_04_inv06 = 1;
    4: op1_04_inv06 = 1;
    12: op1_04_inv06 = 1;
    13: op1_04_inv06 = 1;
    14: op1_04_inv06 = 1;
    15: op1_04_inv06 = 1;
    17: op1_04_inv06 = 1;
    3: op1_04_inv06 = 1;
    19: op1_04_inv06 = 1;
    21: op1_04_inv06 = 1;
    22: op1_04_inv06 = 1;
    23: op1_04_inv06 = 1;
    24: op1_04_inv06 = 1;
    26: op1_04_inv06 = 1;
    27: op1_04_inv06 = 1;
    30: op1_04_inv06 = 1;
    31: op1_04_inv06 = 1;
    32: op1_04_inv06 = 1;
    35: op1_04_inv06 = 1;
    36: op1_04_inv06 = 1;
    37: op1_04_inv06 = 1;
    38: op1_04_inv06 = 1;
    39: op1_04_inv06 = 1;
    42: op1_04_inv06 = 1;
    48: op1_04_inv06 = 1;
    49: op1_04_inv06 = 1;
    56: op1_04_inv06 = 1;
    57: op1_04_inv06 = 1;
    58: op1_04_inv06 = 1;
    59: op1_04_inv06 = 1;
    61: op1_04_inv06 = 1;
    62: op1_04_inv06 = 1;
    66: op1_04_inv06 = 1;
    67: op1_04_inv06 = 1;
    68: op1_04_inv06 = 1;
    70: op1_04_inv06 = 1;
    71: op1_04_inv06 = 1;
    72: op1_04_inv06 = 1;
    73: op1_04_inv06 = 1;
    74: op1_04_inv06 = 1;
    75: op1_04_inv06 = 1;
    79: op1_04_inv06 = 1;
    89: op1_04_inv06 = 1;
    91: op1_04_inv06 = 1;
    92: op1_04_inv06 = 1;
    93: op1_04_inv06 = 1;
    94: op1_04_inv06 = 1;
    97: op1_04_inv06 = 1;
    default: op1_04_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in07 = imem07_in[99:96];
    6: op1_04_in07 = reg_0826;
    7: op1_04_in07 = reg_0696;
    8: op1_04_in07 = reg_0554;
    9: op1_04_in07 = reg_0141;
    10: op1_04_in07 = reg_0256;
    11: op1_04_in07 = reg_1011;
    89: op1_04_in07 = reg_1011;
    4: op1_04_in07 = reg_0427;
    12: op1_04_in07 = reg_0969;
    13: op1_04_in07 = reg_0698;
    14: op1_04_in07 = reg_0980;
    15: op1_04_in07 = reg_0140;
    16: op1_04_in07 = imem00_in[115:112];
    17: op1_04_in07 = imem02_in[123:120];
    18: op1_04_in07 = reg_0372;
    19: op1_04_in07 = reg_0589;
    20: op1_04_in07 = reg_0155;
    21: op1_04_in07 = reg_0665;
    22: op1_04_in07 = reg_0497;
    58: op1_04_in07 = reg_0497;
    23: op1_04_in07 = imem07_in[95:92];
    24: op1_04_in07 = reg_0075;
    25: op1_04_in07 = reg_0679;
    26: op1_04_in07 = imem02_in[11:8];
    27: op1_04_in07 = reg_0450;
    28: op1_04_in07 = reg_0121;
    29: op1_04_in07 = reg_0556;
    30: op1_04_in07 = reg_0430;
    31: op1_04_in07 = imem02_in[67:64];
    32: op1_04_in07 = reg_0738;
    33: op1_04_in07 = reg_0753;
    34: op1_04_in07 = reg_0199;
    35: op1_04_in07 = imem06_in[67:64];
    36: op1_04_in07 = reg_0528;
    37: op1_04_in07 = reg_0585;
    79: op1_04_in07 = reg_0585;
    38: op1_04_in07 = reg_0351;
    39: op1_04_in07 = reg_0701;
    40: op1_04_in07 = reg_0680;
    42: op1_04_in07 = reg_0312;
    43: op1_04_in07 = reg_0813;
    44: op1_04_in07 = reg_0183;
    93: op1_04_in07 = reg_0183;
    45: op1_04_in07 = reg_0125;
    46: op1_04_in07 = reg_0259;
    47: op1_04_in07 = reg_0720;
    48: op1_04_in07 = reg_0686;
    49: op1_04_in07 = reg_0074;
    50: op1_04_in07 = imem03_in[27:24];
    51: op1_04_in07 = reg_0740;
    53: op1_04_in07 = reg_0687;
    54: op1_04_in07 = reg_0110;
    55: op1_04_in07 = reg_0776;
    56: op1_04_in07 = reg_0765;
    57: op1_04_in07 = imem05_in[75:72];
    59: op1_04_in07 = reg_0491;
    60: op1_04_in07 = reg_0744;
    61: op1_04_in07 = reg_0889;
    62: op1_04_in07 = reg_0502;
    63: op1_04_in07 = reg_0485;
    64: op1_04_in07 = reg_0336;
    65: op1_04_in07 = imem04_in[15:12];
    66: op1_04_in07 = imem04_in[79:76];
    67: op1_04_in07 = reg_0307;
    68: op1_04_in07 = reg_0349;
    69: op1_04_in07 = reg_0683;
    70: op1_04_in07 = reg_0323;
    71: op1_04_in07 = imem05_in[127:124];
    72: op1_04_in07 = imem02_in[35:32];
    73: op1_04_in07 = reg_0396;
    74: op1_04_in07 = reg_0483;
    75: op1_04_in07 = reg_0438;
    76: op1_04_in07 = reg_0164;
    78: op1_04_in07 = reg_0356;
    80: op1_04_in07 = imem04_in[71:68];
    81: op1_04_in07 = reg_0226;
    82: op1_04_in07 = reg_0295;
    83: op1_04_in07 = reg_0684;
    84: op1_04_in07 = reg_0422;
    85: op1_04_in07 = reg_1001;
    86: op1_04_in07 = reg_0806;
    87: op1_04_in07 = reg_0003;
    88: op1_04_in07 = imem02_in[75:72];
    90: op1_04_in07 = imem03_in[31:28];
    91: op1_04_in07 = reg_0799;
    92: op1_04_in07 = reg_0815;
    94: op1_04_in07 = reg_0157;
    97: op1_04_in07 = reg_0851;
    default: op1_04_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv07 = 1;
    8: op1_04_inv07 = 1;
    9: op1_04_inv07 = 1;
    11: op1_04_inv07 = 1;
    13: op1_04_inv07 = 1;
    16: op1_04_inv07 = 1;
    19: op1_04_inv07 = 1;
    23: op1_04_inv07 = 1;
    24: op1_04_inv07 = 1;
    26: op1_04_inv07 = 1;
    27: op1_04_inv07 = 1;
    34: op1_04_inv07 = 1;
    36: op1_04_inv07 = 1;
    39: op1_04_inv07 = 1;
    40: op1_04_inv07 = 1;
    43: op1_04_inv07 = 1;
    44: op1_04_inv07 = 1;
    45: op1_04_inv07 = 1;
    48: op1_04_inv07 = 1;
    50: op1_04_inv07 = 1;
    54: op1_04_inv07 = 1;
    55: op1_04_inv07 = 1;
    56: op1_04_inv07 = 1;
    58: op1_04_inv07 = 1;
    60: op1_04_inv07 = 1;
    65: op1_04_inv07 = 1;
    66: op1_04_inv07 = 1;
    67: op1_04_inv07 = 1;
    68: op1_04_inv07 = 1;
    69: op1_04_inv07 = 1;
    70: op1_04_inv07 = 1;
    71: op1_04_inv07 = 1;
    73: op1_04_inv07 = 1;
    75: op1_04_inv07 = 1;
    80: op1_04_inv07 = 1;
    81: op1_04_inv07 = 1;
    82: op1_04_inv07 = 1;
    87: op1_04_inv07 = 1;
    88: op1_04_inv07 = 1;
    89: op1_04_inv07 = 1;
    90: op1_04_inv07 = 1;
    92: op1_04_inv07 = 1;
    93: op1_04_inv07 = 1;
    94: op1_04_inv07 = 1;
    default: op1_04_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in08 = imem07_in[103:100];
    6: op1_04_in08 = reg_0827;
    7: op1_04_in08 = reg_0463;
    78: op1_04_in08 = reg_0463;
    8: op1_04_in08 = reg_0532;
    9: op1_04_in08 = reg_0859;
    10: op1_04_in08 = reg_0274;
    11: op1_04_in08 = imem07_in[3:0];
    4: op1_04_in08 = reg_0437;
    12: op1_04_in08 = reg_0942;
    13: op1_04_in08 = reg_0467;
    14: op1_04_in08 = reg_0975;
    15: op1_04_in08 = reg_0155;
    16: op1_04_in08 = imem00_in[127:124];
    17: op1_04_in08 = reg_0654;
    18: op1_04_in08 = reg_0392;
    19: op1_04_in08 = reg_0600;
    20: op1_04_in08 = reg_0134;
    21: op1_04_in08 = reg_0341;
    22: op1_04_in08 = reg_0132;
    23: op1_04_in08 = imem07_in[107:104];
    24: op1_04_in08 = reg_0072;
    49: op1_04_in08 = reg_0072;
    25: op1_04_in08 = reg_0677;
    26: op1_04_in08 = imem02_in[27:24];
    27: op1_04_in08 = reg_0468;
    28: op1_04_in08 = imem02_in[51:48];
    29: op1_04_in08 = reg_0735;
    30: op1_04_in08 = reg_0432;
    31: op1_04_in08 = imem02_in[71:68];
    32: op1_04_in08 = reg_0058;
    91: op1_04_in08 = reg_0058;
    33: op1_04_in08 = reg_0025;
    34: op1_04_in08 = imem01_in[11:8];
    35: op1_04_in08 = imem06_in[75:72];
    36: op1_04_in08 = reg_0044;
    37: op1_04_in08 = reg_0293;
    38: op1_04_in08 = reg_0264;
    39: op1_04_in08 = reg_0706;
    40: op1_04_in08 = reg_0692;
    42: op1_04_in08 = reg_0844;
    43: op1_04_in08 = reg_0896;
    44: op1_04_in08 = reg_0158;
    45: op1_04_in08 = reg_0104;
    46: op1_04_in08 = reg_0071;
    47: op1_04_in08 = reg_0714;
    48: op1_04_in08 = reg_0679;
    50: op1_04_in08 = imem03_in[39:36];
    51: op1_04_in08 = reg_1017;
    53: op1_04_in08 = reg_0453;
    54: op1_04_in08 = imem02_in[11:8];
    55: op1_04_in08 = reg_0867;
    56: op1_04_in08 = reg_0833;
    57: op1_04_in08 = imem05_in[79:76];
    58: op1_04_in08 = reg_0142;
    59: op1_04_in08 = reg_0750;
    60: op1_04_in08 = reg_0599;
    84: op1_04_in08 = reg_0599;
    61: op1_04_in08 = reg_0384;
    62: op1_04_in08 = reg_0182;
    63: op1_04_in08 = reg_0857;
    64: op1_04_in08 = reg_0052;
    65: op1_04_in08 = imem04_in[31:28];
    66: op1_04_in08 = reg_0277;
    67: op1_04_in08 = reg_0434;
    68: op1_04_in08 = reg_0943;
    69: op1_04_in08 = reg_0685;
    70: op1_04_in08 = reg_0664;
    71: op1_04_in08 = reg_0944;
    72: op1_04_in08 = imem02_in[95:92];
    73: op1_04_in08 = reg_0662;
    74: op1_04_in08 = reg_0301;
    75: op1_04_in08 = reg_0707;
    79: op1_04_in08 = reg_0346;
    80: op1_04_in08 = imem04_in[99:96];
    81: op1_04_in08 = reg_0057;
    82: op1_04_in08 = imem05_in[39:36];
    83: op1_04_in08 = reg_0670;
    85: op1_04_in08 = reg_0974;
    86: op1_04_in08 = reg_0865;
    87: op1_04_in08 = reg_0116;
    88: op1_04_in08 = reg_0334;
    89: op1_04_in08 = reg_0614;
    90: op1_04_in08 = imem03_in[47:44];
    92: op1_04_in08 = reg_0732;
    93: op1_04_in08 = reg_0701;
    97: op1_04_in08 = imem06_in[3:0];
    default: op1_04_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv08 = 1;
    8: op1_04_inv08 = 1;
    4: op1_04_inv08 = 1;
    15: op1_04_inv08 = 1;
    16: op1_04_inv08 = 1;
    17: op1_04_inv08 = 1;
    18: op1_04_inv08 = 1;
    19: op1_04_inv08 = 1;
    20: op1_04_inv08 = 1;
    22: op1_04_inv08 = 1;
    23: op1_04_inv08 = 1;
    24: op1_04_inv08 = 1;
    27: op1_04_inv08 = 1;
    30: op1_04_inv08 = 1;
    31: op1_04_inv08 = 1;
    35: op1_04_inv08 = 1;
    39: op1_04_inv08 = 1;
    40: op1_04_inv08 = 1;
    42: op1_04_inv08 = 1;
    44: op1_04_inv08 = 1;
    47: op1_04_inv08 = 1;
    51: op1_04_inv08 = 1;
    53: op1_04_inv08 = 1;
    55: op1_04_inv08 = 1;
    61: op1_04_inv08 = 1;
    65: op1_04_inv08 = 1;
    68: op1_04_inv08 = 1;
    75: op1_04_inv08 = 1;
    79: op1_04_inv08 = 1;
    83: op1_04_inv08 = 1;
    85: op1_04_inv08 = 1;
    86: op1_04_inv08 = 1;
    87: op1_04_inv08 = 1;
    88: op1_04_inv08 = 1;
    89: op1_04_inv08 = 1;
    91: op1_04_inv08 = 1;
    92: op1_04_inv08 = 1;
    93: op1_04_inv08 = 1;
    default: op1_04_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in09 = imem07_in[115:112];
    6: op1_04_in09 = reg_0828;
    7: op1_04_in09 = reg_0465;
    8: op1_04_in09 = reg_0559;
    9: op1_04_in09 = reg_1019;
    10: op1_04_in09 = reg_0264;
    11: op1_04_in09 = imem07_in[7:4];
    4: op1_04_in09 = reg_0180;
    12: op1_04_in09 = imem05_in[23:20];
    13: op1_04_in09 = reg_0195;
    14: op1_04_in09 = reg_0988;
    15: op1_04_in09 = imem06_in[7:4];
    16: op1_04_in09 = reg_0682;
    17: op1_04_in09 = reg_0333;
    18: op1_04_in09 = reg_0407;
    19: op1_04_in09 = reg_0360;
    20: op1_04_in09 = imem06_in[11:8];
    21: op1_04_in09 = reg_0353;
    22: op1_04_in09 = reg_0142;
    23: op1_04_in09 = imem07_in[123:120];
    24: op1_04_in09 = reg_0882;
    25: op1_04_in09 = reg_0678;
    26: op1_04_in09 = imem02_in[111:108];
    27: op1_04_in09 = reg_0189;
    28: op1_04_in09 = imem02_in[55:52];
    29: op1_04_in09 = reg_0612;
    30: op1_04_in09 = reg_0426;
    31: op1_04_in09 = imem02_in[79:76];
    32: op1_04_in09 = reg_0773;
    33: op1_04_in09 = reg_0404;
    34: op1_04_in09 = imem01_in[31:28];
    35: op1_04_in09 = imem06_in[119:116];
    36: op1_04_in09 = imem05_in[63:60];
    37: op1_04_in09 = reg_0392;
    38: op1_04_in09 = reg_0383;
    39: op1_04_in09 = reg_0727;
    40: op1_04_in09 = reg_0451;
    42: op1_04_in09 = reg_0998;
    43: op1_04_in09 = reg_0832;
    45: op1_04_in09 = reg_0106;
    46: op1_04_in09 = reg_0546;
    47: op1_04_in09 = reg_0713;
    48: op1_04_in09 = reg_0680;
    49: op1_04_in09 = reg_0284;
    50: op1_04_in09 = imem03_in[71:68];
    51: op1_04_in09 = reg_0615;
    53: op1_04_in09 = reg_0455;
    54: op1_04_in09 = imem02_in[35:32];
    55: op1_04_in09 = reg_0484;
    56: op1_04_in09 = reg_0509;
    57: op1_04_in09 = imem05_in[87:84];
    58: op1_04_in09 = reg_0146;
    59: op1_04_in09 = reg_0855;
    60: op1_04_in09 = reg_0640;
    61: op1_04_in09 = reg_0781;
    62: op1_04_in09 = reg_0160;
    63: op1_04_in09 = reg_0642;
    64: op1_04_in09 = reg_0329;
    65: op1_04_in09 = imem04_in[63:60];
    66: op1_04_in09 = reg_0539;
    67: op1_04_in09 = reg_0370;
    68: op1_04_in09 = imem05_in[19:16];
    69: op1_04_in09 = reg_0684;
    70: op1_04_in09 = reg_0007;
    71: op1_04_in09 = reg_0652;
    72: op1_04_in09 = imem02_in[99:96];
    73: op1_04_in09 = reg_0576;
    74: op1_04_in09 = reg_0511;
    75: op1_04_in09 = reg_0970;
    78: op1_04_in09 = reg_0453;
    79: op1_04_in09 = reg_0281;
    80: op1_04_in09 = imem04_in[111:108];
    81: op1_04_in09 = reg_0365;
    82: op1_04_in09 = imem05_in[59:56];
    83: op1_04_in09 = reg_0842;
    84: op1_04_in09 = reg_0350;
    85: op1_04_in09 = reg_0981;
    86: op1_04_in09 = reg_0704;
    87: op1_04_in09 = reg_1033;
    88: op1_04_in09 = reg_0536;
    89: op1_04_in09 = reg_0121;
    90: op1_04_in09 = imem03_in[75:72];
    91: op1_04_in09 = reg_0014;
    92: op1_04_in09 = reg_0893;
    93: op1_04_in09 = reg_0157;
    97: op1_04_in09 = imem06_in[19:16];
    default: op1_04_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_04_inv09 = 1;
    9: op1_04_inv09 = 1;
    11: op1_04_inv09 = 1;
    13: op1_04_inv09 = 1;
    14: op1_04_inv09 = 1;
    15: op1_04_inv09 = 1;
    16: op1_04_inv09 = 1;
    21: op1_04_inv09 = 1;
    23: op1_04_inv09 = 1;
    29: op1_04_inv09 = 1;
    32: op1_04_inv09 = 1;
    33: op1_04_inv09 = 1;
    34: op1_04_inv09 = 1;
    36: op1_04_inv09 = 1;
    37: op1_04_inv09 = 1;
    48: op1_04_inv09 = 1;
    50: op1_04_inv09 = 1;
    51: op1_04_inv09 = 1;
    54: op1_04_inv09 = 1;
    58: op1_04_inv09 = 1;
    59: op1_04_inv09 = 1;
    60: op1_04_inv09 = 1;
    61: op1_04_inv09 = 1;
    66: op1_04_inv09 = 1;
    68: op1_04_inv09 = 1;
    72: op1_04_inv09 = 1;
    78: op1_04_inv09 = 1;
    80: op1_04_inv09 = 1;
    81: op1_04_inv09 = 1;
    82: op1_04_inv09 = 1;
    84: op1_04_inv09 = 1;
    86: op1_04_inv09 = 1;
    91: op1_04_inv09 = 1;
    93: op1_04_inv09 = 1;
    97: op1_04_inv09 = 1;
    default: op1_04_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in10 = reg_0704;
    23: op1_04_in10 = reg_0704;
    6: op1_04_in10 = reg_0829;
    7: op1_04_in10 = reg_0457;
    8: op1_04_in10 = reg_0308;
    9: op1_04_in10 = reg_1021;
    10: op1_04_in10 = reg_0251;
    11: op1_04_in10 = imem07_in[75:72];
    4: op1_04_in10 = reg_0162;
    12: op1_04_in10 = imem05_in[115:112];
    57: op1_04_in10 = imem05_in[115:112];
    13: op1_04_in10 = imem01_in[11:8];
    14: op1_04_in10 = imem04_in[99:96];
    15: op1_04_in10 = imem06_in[31:28];
    16: op1_04_in10 = reg_0672;
    17: op1_04_in10 = reg_0358;
    18: op1_04_in10 = reg_0390;
    19: op1_04_in10 = reg_0370;
    20: op1_04_in10 = imem06_in[39:36];
    97: op1_04_in10 = imem06_in[39:36];
    21: op1_04_in10 = imem02_in[3:0];
    22: op1_04_in10 = reg_0146;
    24: op1_04_in10 = reg_0058;
    25: op1_04_in10 = reg_0688;
    26: op1_04_in10 = imem02_in[119:116];
    27: op1_04_in10 = reg_0190;
    28: op1_04_in10 = imem02_in[59:56];
    29: op1_04_in10 = imem06_in[15:12];
    30: op1_04_in10 = reg_0419;
    31: op1_04_in10 = imem02_in[87:84];
    32: op1_04_in10 = imem05_in[95:92];
    33: op1_04_in10 = reg_0018;
    34: op1_04_in10 = imem01_in[59:56];
    35: op1_04_in10 = reg_0628;
    36: op1_04_in10 = imem05_in[103:100];
    37: op1_04_in10 = reg_0741;
    38: op1_04_in10 = reg_0243;
    39: op1_04_in10 = reg_0436;
    40: op1_04_in10 = reg_0469;
    42: op1_04_in10 = reg_1002;
    43: op1_04_in10 = reg_0831;
    45: op1_04_in10 = reg_0036;
    46: op1_04_in10 = reg_0551;
    47: op1_04_in10 = reg_0701;
    48: op1_04_in10 = reg_0699;
    49: op1_04_in10 = imem04_in[23:20];
    50: op1_04_in10 = imem03_in[83:80];
    51: op1_04_in10 = reg_0124;
    53: op1_04_in10 = reg_0460;
    54: op1_04_in10 = imem02_in[75:72];
    55: op1_04_in10 = reg_0405;
    56: op1_04_in10 = reg_0376;
    58: op1_04_in10 = reg_0143;
    59: op1_04_in10 = reg_0588;
    60: op1_04_in10 = reg_0168;
    61: op1_04_in10 = reg_0382;
    62: op1_04_in10 = reg_0184;
    63: op1_04_in10 = reg_0281;
    64: op1_04_in10 = reg_0818;
    65: op1_04_in10 = imem04_in[87:84];
    66: op1_04_in10 = reg_0541;
    67: op1_04_in10 = reg_0795;
    68: op1_04_in10 = imem05_in[23:20];
    69: op1_04_in10 = reg_0069;
    70: op1_04_in10 = reg_0482;
    71: op1_04_in10 = reg_0655;
    72: op1_04_in10 = reg_0279;
    73: op1_04_in10 = reg_0397;
    74: op1_04_in10 = reg_0306;
    75: op1_04_in10 = reg_0145;
    78: op1_04_in10 = reg_0462;
    79: op1_04_in10 = reg_0040;
    80: op1_04_in10 = reg_0483;
    81: op1_04_in10 = reg_0958;
    82: op1_04_in10 = imem05_in[119:116];
    83: op1_04_in10 = reg_0499;
    84: op1_04_in10 = reg_0589;
    85: op1_04_in10 = reg_0988;
    86: op1_04_in10 = reg_0093;
    87: op1_04_in10 = reg_0101;
    88: op1_04_in10 = reg_0073;
    89: op1_04_in10 = reg_0320;
    90: op1_04_in10 = reg_0147;
    91: op1_04_in10 = reg_0296;
    92: op1_04_in10 = reg_0764;
    default: op1_04_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv10 = 1;
    11: op1_04_inv10 = 1;
    15: op1_04_inv10 = 1;
    16: op1_04_inv10 = 1;
    17: op1_04_inv10 = 1;
    18: op1_04_inv10 = 1;
    19: op1_04_inv10 = 1;
    21: op1_04_inv10 = 1;
    22: op1_04_inv10 = 1;
    24: op1_04_inv10 = 1;
    25: op1_04_inv10 = 1;
    26: op1_04_inv10 = 1;
    27: op1_04_inv10 = 1;
    28: op1_04_inv10 = 1;
    31: op1_04_inv10 = 1;
    33: op1_04_inv10 = 1;
    35: op1_04_inv10 = 1;
    36: op1_04_inv10 = 1;
    38: op1_04_inv10 = 1;
    39: op1_04_inv10 = 1;
    42: op1_04_inv10 = 1;
    43: op1_04_inv10 = 1;
    47: op1_04_inv10 = 1;
    50: op1_04_inv10 = 1;
    51: op1_04_inv10 = 1;
    53: op1_04_inv10 = 1;
    54: op1_04_inv10 = 1;
    57: op1_04_inv10 = 1;
    60: op1_04_inv10 = 1;
    61: op1_04_inv10 = 1;
    62: op1_04_inv10 = 1;
    63: op1_04_inv10 = 1;
    64: op1_04_inv10 = 1;
    69: op1_04_inv10 = 1;
    70: op1_04_inv10 = 1;
    71: op1_04_inv10 = 1;
    72: op1_04_inv10 = 1;
    74: op1_04_inv10 = 1;
    80: op1_04_inv10 = 1;
    84: op1_04_inv10 = 1;
    89: op1_04_inv10 = 1;
    90: op1_04_inv10 = 1;
    97: op1_04_inv10 = 1;
    default: op1_04_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in11 = reg_0717;
    6: op1_04_in11 = imem05_in[59:56];
    7: op1_04_in11 = reg_0477;
    8: op1_04_in11 = reg_0283;
    9: op1_04_in11 = reg_0613;
    10: op1_04_in11 = reg_0257;
    11: op1_04_in11 = imem07_in[87:84];
    4: op1_04_in11 = reg_0169;
    12: op1_04_in11 = reg_0132;
    13: op1_04_in11 = imem01_in[19:16];
    14: op1_04_in11 = imem04_in[111:108];
    15: op1_04_in11 = imem06_in[95:92];
    16: op1_04_in11 = reg_0461;
    17: op1_04_in11 = reg_0341;
    18: op1_04_in11 = reg_0005;
    19: op1_04_in11 = reg_0319;
    20: op1_04_in11 = imem06_in[71:68];
    97: op1_04_in11 = imem06_in[71:68];
    21: op1_04_in11 = imem02_in[19:16];
    22: op1_04_in11 = reg_0138;
    23: op1_04_in11 = reg_0719;
    24: op1_04_in11 = reg_0774;
    25: op1_04_in11 = reg_0673;
    71: op1_04_in11 = reg_0673;
    26: op1_04_in11 = imem02_in[127:124];
    27: op1_04_in11 = imem01_in[79:76];
    28: op1_04_in11 = imem02_in[91:88];
    29: op1_04_in11 = imem06_in[39:36];
    30: op1_04_in11 = reg_0440;
    31: op1_04_in11 = imem02_in[95:92];
    54: op1_04_in11 = imem02_in[95:92];
    32: op1_04_in11 = imem05_in[111:108];
    36: op1_04_in11 = imem05_in[111:108];
    33: op1_04_in11 = reg_0597;
    34: op1_04_in11 = imem01_in[87:84];
    35: op1_04_in11 = reg_0621;
    37: op1_04_in11 = reg_0382;
    38: op1_04_in11 = reg_0349;
    39: op1_04_in11 = reg_0439;
    40: op1_04_in11 = reg_0475;
    42: op1_04_in11 = reg_0991;
    43: op1_04_in11 = reg_0136;
    45: op1_04_in11 = reg_0314;
    46: op1_04_in11 = reg_0547;
    47: op1_04_in11 = reg_0706;
    48: op1_04_in11 = reg_0450;
    49: op1_04_in11 = imem04_in[47:44];
    50: op1_04_in11 = imem03_in[91:88];
    51: op1_04_in11 = reg_0111;
    53: op1_04_in11 = reg_0456;
    55: op1_04_in11 = reg_0743;
    56: op1_04_in11 = reg_0822;
    57: op1_04_in11 = imem05_in[123:120];
    58: op1_04_in11 = reg_0139;
    59: op1_04_in11 = reg_0579;
    61: op1_04_in11 = reg_0699;
    63: op1_04_in11 = reg_0381;
    64: op1_04_in11 = reg_0037;
    65: op1_04_in11 = imem04_in[95:92];
    66: op1_04_in11 = reg_0802;
    67: op1_04_in11 = reg_0311;
    68: op1_04_in11 = imem05_in[43:40];
    69: op1_04_in11 = reg_0669;
    70: op1_04_in11 = reg_0088;
    72: op1_04_in11 = reg_0359;
    73: op1_04_in11 = reg_1008;
    79: op1_04_in11 = reg_1008;
    74: op1_04_in11 = reg_0055;
    75: op1_04_in11 = reg_0651;
    78: op1_04_in11 = reg_0458;
    80: op1_04_in11 = reg_0778;
    81: op1_04_in11 = reg_0150;
    82: op1_04_in11 = reg_0492;
    83: op1_04_in11 = reg_0457;
    84: op1_04_in11 = reg_0420;
    85: op1_04_in11 = reg_1000;
    86: op1_04_in11 = reg_0482;
    87: op1_04_in11 = reg_0877;
    88: op1_04_in11 = reg_0323;
    89: op1_04_in11 = reg_0011;
    90: op1_04_in11 = reg_0540;
    91: op1_04_in11 = reg_0074;
    92: op1_04_in11 = reg_0552;
    default: op1_04_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv11 = 1;
    6: op1_04_inv11 = 1;
    9: op1_04_inv11 = 1;
    4: op1_04_inv11 = 1;
    17: op1_04_inv11 = 1;
    19: op1_04_inv11 = 1;
    21: op1_04_inv11 = 1;
    23: op1_04_inv11 = 1;
    24: op1_04_inv11 = 1;
    25: op1_04_inv11 = 1;
    27: op1_04_inv11 = 1;
    30: op1_04_inv11 = 1;
    35: op1_04_inv11 = 1;
    38: op1_04_inv11 = 1;
    46: op1_04_inv11 = 1;
    50: op1_04_inv11 = 1;
    54: op1_04_inv11 = 1;
    57: op1_04_inv11 = 1;
    64: op1_04_inv11 = 1;
    67: op1_04_inv11 = 1;
    72: op1_04_inv11 = 1;
    74: op1_04_inv11 = 1;
    75: op1_04_inv11 = 1;
    79: op1_04_inv11 = 1;
    82: op1_04_inv11 = 1;
    85: op1_04_inv11 = 1;
    86: op1_04_inv11 = 1;
    88: op1_04_inv11 = 1;
    89: op1_04_inv11 = 1;
    90: op1_04_inv11 = 1;
    91: op1_04_inv11 = 1;
    default: op1_04_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in12 = reg_0718;
    6: op1_04_in12 = imem05_in[99:96];
    7: op1_04_in12 = reg_0466;
    8: op1_04_in12 = reg_0293;
    9: op1_04_in12 = reg_0617;
    10: op1_04_in12 = reg_0272;
    45: op1_04_in12 = reg_0272;
    11: op1_04_in12 = imem07_in[103:100];
    4: op1_04_in12 = reg_0166;
    12: op1_04_in12 = reg_0152;
    13: op1_04_in12 = imem01_in[99:96];
    14: op1_04_in12 = reg_0552;
    15: op1_04_in12 = imem06_in[115:112];
    20: op1_04_in12 = imem06_in[115:112];
    16: op1_04_in12 = reg_0469;
    17: op1_04_in12 = reg_0330;
    18: op1_04_in12 = reg_0754;
    19: op1_04_in12 = reg_0322;
    21: op1_04_in12 = imem02_in[87:84];
    22: op1_04_in12 = reg_0140;
    23: op1_04_in12 = reg_0720;
    24: op1_04_in12 = reg_0057;
    25: op1_04_in12 = reg_0461;
    26: op1_04_in12 = reg_0758;
    27: op1_04_in12 = imem01_in[107:104];
    28: op1_04_in12 = imem02_in[103:100];
    29: op1_04_in12 = imem06_in[103:100];
    30: op1_04_in12 = reg_0442;
    31: op1_04_in12 = reg_0642;
    32: op1_04_in12 = reg_0963;
    33: op1_04_in12 = imem07_in[3:0];
    34: op1_04_in12 = reg_0013;
    71: op1_04_in12 = reg_0013;
    35: op1_04_in12 = reg_0631;
    36: op1_04_in12 = imem05_in[119:116];
    37: op1_04_in12 = reg_0804;
    38: op1_04_in12 = reg_0384;
    39: op1_04_in12 = reg_0167;
    40: op1_04_in12 = reg_0470;
    42: op1_04_in12 = reg_0992;
    43: op1_04_in12 = reg_0150;
    46: op1_04_in12 = reg_1003;
    47: op1_04_in12 = reg_0744;
    48: op1_04_in12 = reg_0451;
    49: op1_04_in12 = imem04_in[63:60];
    50: op1_04_in12 = imem03_in[127:124];
    51: op1_04_in12 = reg_0116;
    53: op1_04_in12 = reg_0186;
    54: op1_04_in12 = reg_0363;
    55: op1_04_in12 = reg_0318;
    56: op1_04_in12 = reg_0987;
    57: op1_04_in12 = imem05_in[127:124];
    58: op1_04_in12 = reg_0131;
    59: op1_04_in12 = reg_1006;
    61: op1_04_in12 = reg_0222;
    63: op1_04_in12 = imem02_in[35:32];
    64: op1_04_in12 = reg_0335;
    65: op1_04_in12 = imem04_in[99:96];
    66: op1_04_in12 = reg_0752;
    67: op1_04_in12 = reg_0991;
    68: op1_04_in12 = imem05_in[47:44];
    69: op1_04_in12 = reg_0477;
    70: op1_04_in12 = reg_0084;
    72: op1_04_in12 = reg_0329;
    73: op1_04_in12 = reg_0376;
    74: op1_04_in12 = reg_0048;
    75: op1_04_in12 = reg_0528;
    78: op1_04_in12 = reg_0200;
    79: op1_04_in12 = reg_0773;
    80: op1_04_in12 = reg_0537;
    81: op1_04_in12 = reg_1015;
    82: op1_04_in12 = reg_0128;
    83: op1_04_in12 = reg_0476;
    84: op1_04_in12 = reg_0640;
    85: op1_04_in12 = imem04_in[15:12];
    86: op1_04_in12 = reg_0263;
    87: op1_04_in12 = reg_0110;
    88: op1_04_in12 = reg_0424;
    89: op1_04_in12 = reg_0781;
    90: op1_04_in12 = reg_0888;
    91: op1_04_in12 = reg_0854;
    92: op1_04_in12 = reg_0494;
    97: op1_04_in12 = imem06_in[91:88];
    default: op1_04_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv12 = 1;
    7: op1_04_inv12 = 1;
    8: op1_04_inv12 = 1;
    9: op1_04_inv12 = 1;
    10: op1_04_inv12 = 1;
    4: op1_04_inv12 = 1;
    12: op1_04_inv12 = 1;
    15: op1_04_inv12 = 1;
    17: op1_04_inv12 = 1;
    18: op1_04_inv12 = 1;
    19: op1_04_inv12 = 1;
    21: op1_04_inv12 = 1;
    22: op1_04_inv12 = 1;
    26: op1_04_inv12 = 1;
    29: op1_04_inv12 = 1;
    35: op1_04_inv12 = 1;
    36: op1_04_inv12 = 1;
    38: op1_04_inv12 = 1;
    42: op1_04_inv12 = 1;
    43: op1_04_inv12 = 1;
    45: op1_04_inv12 = 1;
    46: op1_04_inv12 = 1;
    48: op1_04_inv12 = 1;
    50: op1_04_inv12 = 1;
    54: op1_04_inv12 = 1;
    55: op1_04_inv12 = 1;
    56: op1_04_inv12 = 1;
    58: op1_04_inv12 = 1;
    61: op1_04_inv12 = 1;
    63: op1_04_inv12 = 1;
    65: op1_04_inv12 = 1;
    66: op1_04_inv12 = 1;
    71: op1_04_inv12 = 1;
    72: op1_04_inv12 = 1;
    73: op1_04_inv12 = 1;
    74: op1_04_inv12 = 1;
    79: op1_04_inv12 = 1;
    80: op1_04_inv12 = 1;
    82: op1_04_inv12 = 1;
    83: op1_04_inv12 = 1;
    88: op1_04_inv12 = 1;
    89: op1_04_inv12 = 1;
    90: op1_04_inv12 = 1;
    92: op1_04_inv12 = 1;
    default: op1_04_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in13 = reg_0706;
    6: op1_04_in13 = reg_0267;
    7: op1_04_in13 = reg_0474;
    8: op1_04_in13 = reg_0046;
    9: op1_04_in13 = reg_0606;
    10: op1_04_in13 = reg_0261;
    11: op1_04_in13 = reg_0704;
    4: op1_04_in13 = reg_0185;
    12: op1_04_in13 = reg_0153;
    13: op1_04_in13 = imem01_in[115:112];
    14: op1_04_in13 = reg_0555;
    15: op1_04_in13 = reg_0630;
    16: op1_04_in13 = reg_0472;
    17: op1_04_in13 = reg_0363;
    18: op1_04_in13 = imem07_in[75:72];
    19: op1_04_in13 = reg_0396;
    20: op1_04_in13 = imem06_in[119:116];
    21: op1_04_in13 = imem03_in[7:4];
    22: op1_04_in13 = imem06_in[35:32];
    23: op1_04_in13 = reg_0730;
    24: op1_04_in13 = imem05_in[39:36];
    25: op1_04_in13 = reg_0462;
    83: op1_04_in13 = reg_0462;
    26: op1_04_in13 = reg_0089;
    27: op1_04_in13 = reg_0786;
    28: op1_04_in13 = reg_0650;
    31: op1_04_in13 = reg_0650;
    29: op1_04_in13 = imem06_in[107:104];
    30: op1_04_in13 = reg_0180;
    32: op1_04_in13 = reg_0970;
    33: op1_04_in13 = imem07_in[23:20];
    34: op1_04_in13 = reg_0242;
    35: op1_04_in13 = reg_0626;
    36: op1_04_in13 = reg_0954;
    82: op1_04_in13 = reg_0954;
    37: op1_04_in13 = reg_0388;
    38: op1_04_in13 = reg_0628;
    40: op1_04_in13 = reg_0468;
    42: op1_04_in13 = reg_0989;
    43: op1_04_in13 = reg_0152;
    45: op1_04_in13 = imem02_in[63:60];
    46: op1_04_in13 = reg_0265;
    47: op1_04_in13 = reg_0589;
    48: op1_04_in13 = reg_0455;
    49: op1_04_in13 = imem04_in[75:72];
    50: op1_04_in13 = reg_0492;
    51: op1_04_in13 = reg_0115;
    53: op1_04_in13 = reg_0199;
    54: op1_04_in13 = reg_0656;
    55: op1_04_in13 = reg_0676;
    56: op1_04_in13 = reg_1001;
    57: op1_04_in13 = reg_0581;
    58: op1_04_in13 = reg_0144;
    59: op1_04_in13 = reg_1009;
    61: op1_04_in13 = reg_0619;
    63: op1_04_in13 = imem02_in[47:44];
    64: op1_04_in13 = reg_0516;
    65: op1_04_in13 = reg_0313;
    66: op1_04_in13 = reg_0808;
    67: op1_04_in13 = reg_0980;
    68: op1_04_in13 = imem05_in[51:48];
    69: op1_04_in13 = reg_0459;
    70: op1_04_in13 = reg_0872;
    71: op1_04_in13 = reg_0689;
    72: op1_04_in13 = reg_0644;
    73: op1_04_in13 = reg_0820;
    74: op1_04_in13 = reg_0014;
    75: op1_04_in13 = reg_0490;
    78: op1_04_in13 = reg_0193;
    79: op1_04_in13 = reg_1049;
    80: op1_04_in13 = reg_0276;
    81: op1_04_in13 = reg_0154;
    84: op1_04_in13 = reg_0431;
    85: op1_04_in13 = imem04_in[19:16];
    86: op1_04_in13 = reg_0344;
    87: op1_04_in13 = imem02_in[3:0];
    88: op1_04_in13 = reg_0054;
    89: op1_04_in13 = imem06_in[63:60];
    90: op1_04_in13 = reg_0031;
    91: op1_04_in13 = reg_0071;
    92: op1_04_in13 = reg_0824;
    97: op1_04_in13 = imem06_in[111:108];
    default: op1_04_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv13 = 1;
    6: op1_04_inv13 = 1;
    7: op1_04_inv13 = 1;
    8: op1_04_inv13 = 1;
    9: op1_04_inv13 = 1;
    11: op1_04_inv13 = 1;
    13: op1_04_inv13 = 1;
    15: op1_04_inv13 = 1;
    18: op1_04_inv13 = 1;
    19: op1_04_inv13 = 1;
    20: op1_04_inv13 = 1;
    21: op1_04_inv13 = 1;
    22: op1_04_inv13 = 1;
    23: op1_04_inv13 = 1;
    24: op1_04_inv13 = 1;
    25: op1_04_inv13 = 1;
    26: op1_04_inv13 = 1;
    28: op1_04_inv13 = 1;
    30: op1_04_inv13 = 1;
    31: op1_04_inv13 = 1;
    32: op1_04_inv13 = 1;
    33: op1_04_inv13 = 1;
    42: op1_04_inv13 = 1;
    43: op1_04_inv13 = 1;
    46: op1_04_inv13 = 1;
    48: op1_04_inv13 = 1;
    54: op1_04_inv13 = 1;
    57: op1_04_inv13 = 1;
    64: op1_04_inv13 = 1;
    66: op1_04_inv13 = 1;
    67: op1_04_inv13 = 1;
    69: op1_04_inv13 = 1;
    72: op1_04_inv13 = 1;
    73: op1_04_inv13 = 1;
    74: op1_04_inv13 = 1;
    75: op1_04_inv13 = 1;
    78: op1_04_inv13 = 1;
    83: op1_04_inv13 = 1;
    84: op1_04_inv13 = 1;
    85: op1_04_inv13 = 1;
    86: op1_04_inv13 = 1;
    87: op1_04_inv13 = 1;
    97: op1_04_inv13 = 1;
    default: op1_04_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in14 = reg_0423;
    6: op1_04_in14 = reg_0268;
    7: op1_04_in14 = reg_0471;
    16: op1_04_in14 = reg_0471;
    8: op1_04_in14 = reg_0054;
    9: op1_04_in14 = reg_0577;
    10: op1_04_in14 = reg_0253;
    11: op1_04_in14 = reg_0719;
    4: op1_04_in14 = reg_0173;
    12: op1_04_in14 = reg_0130;
    13: op1_04_in14 = reg_0013;
    14: op1_04_in14 = reg_0547;
    15: op1_04_in14 = reg_0626;
    17: op1_04_in14 = reg_0092;
    18: op1_04_in14 = imem07_in[115:112];
    19: op1_04_in14 = reg_0984;
    20: op1_04_in14 = reg_0614;
    21: op1_04_in14 = imem03_in[27:24];
    22: op1_04_in14 = imem06_in[47:44];
    23: op1_04_in14 = reg_0723;
    24: op1_04_in14 = imem05_in[75:72];
    25: op1_04_in14 = reg_0480;
    26: op1_04_in14 = reg_0084;
    64: op1_04_in14 = reg_0084;
    27: op1_04_in14 = reg_0223;
    28: op1_04_in14 = reg_0645;
    29: op1_04_in14 = imem06_in[111:108];
    30: op1_04_in14 = reg_0163;
    31: op1_04_in14 = reg_0666;
    32: op1_04_in14 = reg_0959;
    33: op1_04_in14 = imem07_in[51:48];
    34: op1_04_in14 = reg_0240;
    35: op1_04_in14 = reg_0622;
    36: op1_04_in14 = reg_0956;
    37: op1_04_in14 = reg_0390;
    38: op1_04_in14 = reg_0625;
    40: op1_04_in14 = reg_0213;
    42: op1_04_in14 = reg_0990;
    43: op1_04_in14 = reg_0153;
    45: op1_04_in14 = imem02_in[99:96];
    46: op1_04_in14 = reg_1009;
    47: op1_04_in14 = reg_0175;
    48: op1_04_in14 = reg_0472;
    49: op1_04_in14 = imem04_in[115:112];
    50: op1_04_in14 = reg_1007;
    51: op1_04_in14 = reg_0110;
    53: op1_04_in14 = reg_0105;
    54: op1_04_in14 = reg_0300;
    55: op1_04_in14 = reg_0567;
    56: op1_04_in14 = reg_0980;
    57: op1_04_in14 = reg_0955;
    58: op1_04_in14 = reg_0387;
    59: op1_04_in14 = reg_0932;
    61: op1_04_in14 = imem06_in[11:8];
    63: op1_04_in14 = imem02_in[95:92];
    65: op1_04_in14 = reg_0799;
    66: op1_04_in14 = reg_0815;
    67: op1_04_in14 = reg_0999;
    68: op1_04_in14 = reg_0675;
    69: op1_04_in14 = reg_0214;
    70: op1_04_in14 = reg_0079;
    71: op1_04_in14 = reg_0784;
    72: op1_04_in14 = reg_0335;
    73: op1_04_in14 = reg_0985;
    74: op1_04_in14 = reg_0276;
    75: op1_04_in14 = reg_0144;
    78: op1_04_in14 = reg_0186;
    79: op1_04_in14 = reg_0779;
    80: op1_04_in14 = reg_0401;
    81: op1_04_in14 = reg_0892;
    82: op1_04_in14 = reg_0235;
    83: op1_04_in14 = reg_0474;
    84: op1_04_in14 = reg_0429;
    85: op1_04_in14 = imem04_in[23:20];
    86: op1_04_in14 = reg_0262;
    87: op1_04_in14 = imem02_in[11:8];
    88: op1_04_in14 = reg_0083;
    89: op1_04_in14 = imem06_in[75:72];
    90: op1_04_in14 = reg_0016;
    91: op1_04_in14 = reg_0542;
    92: op1_04_in14 = reg_0332;
    97: op1_04_in14 = reg_0351;
    default: op1_04_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv14 = 1;
    10: op1_04_inv14 = 1;
    11: op1_04_inv14 = 1;
    4: op1_04_inv14 = 1;
    12: op1_04_inv14 = 1;
    13: op1_04_inv14 = 1;
    14: op1_04_inv14 = 1;
    16: op1_04_inv14 = 1;
    18: op1_04_inv14 = 1;
    21: op1_04_inv14 = 1;
    22: op1_04_inv14 = 1;
    25: op1_04_inv14 = 1;
    26: op1_04_inv14 = 1;
    33: op1_04_inv14 = 1;
    34: op1_04_inv14 = 1;
    36: op1_04_inv14 = 1;
    37: op1_04_inv14 = 1;
    38: op1_04_inv14 = 1;
    42: op1_04_inv14 = 1;
    46: op1_04_inv14 = 1;
    47: op1_04_inv14 = 1;
    49: op1_04_inv14 = 1;
    50: op1_04_inv14 = 1;
    51: op1_04_inv14 = 1;
    54: op1_04_inv14 = 1;
    56: op1_04_inv14 = 1;
    58: op1_04_inv14 = 1;
    59: op1_04_inv14 = 1;
    63: op1_04_inv14 = 1;
    65: op1_04_inv14 = 1;
    68: op1_04_inv14 = 1;
    70: op1_04_inv14 = 1;
    74: op1_04_inv14 = 1;
    75: op1_04_inv14 = 1;
    78: op1_04_inv14 = 1;
    79: op1_04_inv14 = 1;
    81: op1_04_inv14 = 1;
    83: op1_04_inv14 = 1;
    85: op1_04_inv14 = 1;
    86: op1_04_inv14 = 1;
    87: op1_04_inv14 = 1;
    88: op1_04_inv14 = 1;
    90: op1_04_inv14 = 1;
    97: op1_04_inv14 = 1;
    default: op1_04_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in15 = reg_0180;
    6: op1_04_in15 = reg_0252;
    7: op1_04_in15 = reg_0478;
    8: op1_04_in15 = reg_0067;
    9: op1_04_in15 = reg_0402;
    10: op1_04_in15 = reg_0132;
    11: op1_04_in15 = reg_0726;
    4: op1_04_in15 = reg_0184;
    12: op1_04_in15 = reg_0155;
    13: op1_04_in15 = reg_0766;
    14: op1_04_in15 = reg_0308;
    15: op1_04_in15 = reg_0349;
    16: op1_04_in15 = reg_0458;
    17: op1_04_in15 = reg_0084;
    18: op1_04_in15 = reg_0714;
    19: op1_04_in15 = reg_0997;
    20: op1_04_in15 = reg_0617;
    21: op1_04_in15 = imem03_in[107:104];
    22: op1_04_in15 = imem06_in[119:116];
    23: op1_04_in15 = reg_0700;
    24: op1_04_in15 = imem05_in[103:100];
    25: op1_04_in15 = reg_0471;
    26: op1_04_in15 = reg_0310;
    27: op1_04_in15 = reg_0299;
    28: op1_04_in15 = reg_0655;
    29: op1_04_in15 = reg_0787;
    30: op1_04_in15 = reg_0185;
    31: op1_04_in15 = reg_0639;
    32: op1_04_in15 = reg_0956;
    33: op1_04_in15 = imem07_in[63:60];
    34: op1_04_in15 = reg_0828;
    35: op1_04_in15 = reg_0392;
    36: op1_04_in15 = reg_0948;
    37: op1_04_in15 = reg_0222;
    38: op1_04_in15 = reg_1010;
    40: op1_04_in15 = reg_0196;
    42: op1_04_in15 = reg_1000;
    43: op1_04_in15 = imem06_in[67:64];
    45: op1_04_in15 = reg_0334;
    46: op1_04_in15 = reg_0277;
    47: op1_04_in15 = reg_0172;
    48: op1_04_in15 = reg_0480;
    49: op1_04_in15 = imem05_in[15:12];
    50: op1_04_in15 = reg_0358;
    51: op1_04_in15 = imem02_in[51:48];
    53: op1_04_in15 = reg_1042;
    54: op1_04_in15 = reg_0739;
    55: op1_04_in15 = reg_0552;
    56: op1_04_in15 = reg_0999;
    57: op1_04_in15 = reg_0225;
    58: op1_04_in15 = reg_0631;
    59: op1_04_in15 = reg_0050;
    61: op1_04_in15 = imem06_in[27:24];
    63: op1_04_in15 = imem02_in[103:100];
    64: op1_04_in15 = reg_0884;
    65: op1_04_in15 = reg_0076;
    66: op1_04_in15 = reg_0809;
    67: op1_04_in15 = reg_0975;
    68: op1_04_in15 = reg_0125;
    69: op1_04_in15 = reg_0208;
    70: op1_04_in15 = reg_0019;
    71: op1_04_in15 = reg_0438;
    72: op1_04_in15 = reg_0088;
    73: op1_04_in15 = reg_0987;
    74: op1_04_in15 = reg_0808;
    75: op1_04_in15 = imem06_in[23:20];
    78: op1_04_in15 = reg_0194;
    79: op1_04_in15 = reg_0597;
    80: op1_04_in15 = reg_0064;
    81: op1_04_in15 = reg_0336;
    82: op1_04_in15 = reg_0140;
    83: op1_04_in15 = reg_0209;
    84: op1_04_in15 = reg_0181;
    85: op1_04_in15 = imem04_in[35:32];
    86: op1_04_in15 = reg_0679;
    87: op1_04_in15 = imem02_in[47:44];
    88: op1_04_in15 = reg_0381;
    89: op1_04_in15 = imem06_in[115:112];
    90: op1_04_in15 = reg_0909;
    91: op1_04_in15 = reg_0044;
    92: op1_04_in15 = imem05_in[43:40];
    97: op1_04_in15 = reg_0626;
    default: op1_04_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_04_inv15 = 1;
    9: op1_04_inv15 = 1;
    10: op1_04_inv15 = 1;
    11: op1_04_inv15 = 1;
    13: op1_04_inv15 = 1;
    14: op1_04_inv15 = 1;
    20: op1_04_inv15 = 1;
    21: op1_04_inv15 = 1;
    25: op1_04_inv15 = 1;
    26: op1_04_inv15 = 1;
    28: op1_04_inv15 = 1;
    29: op1_04_inv15 = 1;
    31: op1_04_inv15 = 1;
    32: op1_04_inv15 = 1;
    33: op1_04_inv15 = 1;
    34: op1_04_inv15 = 1;
    35: op1_04_inv15 = 1;
    47: op1_04_inv15 = 1;
    48: op1_04_inv15 = 1;
    49: op1_04_inv15 = 1;
    50: op1_04_inv15 = 1;
    51: op1_04_inv15 = 1;
    53: op1_04_inv15 = 1;
    54: op1_04_inv15 = 1;
    55: op1_04_inv15 = 1;
    59: op1_04_inv15 = 1;
    61: op1_04_inv15 = 1;
    63: op1_04_inv15 = 1;
    64: op1_04_inv15 = 1;
    65: op1_04_inv15 = 1;
    67: op1_04_inv15 = 1;
    68: op1_04_inv15 = 1;
    70: op1_04_inv15 = 1;
    71: op1_04_inv15 = 1;
    72: op1_04_inv15 = 1;
    73: op1_04_inv15 = 1;
    74: op1_04_inv15 = 1;
    75: op1_04_inv15 = 1;
    78: op1_04_inv15 = 1;
    79: op1_04_inv15 = 1;
    81: op1_04_inv15 = 1;
    82: op1_04_inv15 = 1;
    84: op1_04_inv15 = 1;
    85: op1_04_inv15 = 1;
    87: op1_04_inv15 = 1;
    88: op1_04_inv15 = 1;
    90: op1_04_inv15 = 1;
    91: op1_04_inv15 = 1;
    92: op1_04_inv15 = 1;
    default: op1_04_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in16 = reg_0166;
    6: op1_04_in16 = reg_0243;
    7: op1_04_in16 = reg_0210;
    16: op1_04_in16 = reg_0210;
    8: op1_04_in16 = reg_0043;
    9: op1_04_in16 = reg_0372;
    10: op1_04_in16 = reg_0147;
    11: op1_04_in16 = reg_0713;
    12: op1_04_in16 = reg_0144;
    13: op1_04_in16 = reg_1042;
    14: op1_04_in16 = reg_0301;
    15: op1_04_in16 = reg_0407;
    17: op1_04_in16 = reg_0073;
    18: op1_04_in16 = reg_0709;
    19: op1_04_in16 = reg_0912;
    20: op1_04_in16 = reg_0615;
    21: op1_04_in16 = reg_0598;
    22: op1_04_in16 = reg_0610;
    23: op1_04_in16 = reg_0727;
    24: op1_04_in16 = reg_0966;
    25: op1_04_in16 = reg_0458;
    26: op1_04_in16 = imem03_in[15:12];
    27: op1_04_in16 = reg_0769;
    28: op1_04_in16 = reg_0661;
    29: op1_04_in16 = reg_0801;
    30: op1_04_in16 = reg_0168;
    31: op1_04_in16 = reg_0652;
    32: op1_04_in16 = reg_0969;
    33: op1_04_in16 = imem07_in[71:68];
    34: op1_04_in16 = reg_0236;
    35: op1_04_in16 = reg_0382;
    36: op1_04_in16 = reg_0961;
    37: op1_04_in16 = reg_0917;
    38: op1_04_in16 = reg_0008;
    40: op1_04_in16 = reg_0271;
    42: op1_04_in16 = reg_0557;
    43: op1_04_in16 = reg_0614;
    45: op1_04_in16 = reg_0081;
    46: op1_04_in16 = reg_1020;
    47: op1_04_in16 = reg_0159;
    48: op1_04_in16 = reg_0468;
    49: op1_04_in16 = imem05_in[23:20];
    50: op1_04_in16 = reg_0581;
    51: op1_04_in16 = reg_0639;
    53: op1_04_in16 = reg_0108;
    54: op1_04_in16 = reg_0664;
    55: op1_04_in16 = imem03_in[51:48];
    56: op1_04_in16 = reg_0988;
    57: op1_04_in16 = reg_0908;
    58: op1_04_in16 = reg_0390;
    59: op1_04_in16 = reg_0507;
    61: op1_04_in16 = imem06_in[63:60];
    63: op1_04_in16 = imem02_in[111:108];
    64: op1_04_in16 = reg_0079;
    65: op1_04_in16 = reg_0056;
    66: op1_04_in16 = reg_0732;
    67: op1_04_in16 = reg_0976;
    68: op1_04_in16 = reg_0149;
    69: op1_04_in16 = reg_0211;
    70: op1_04_in16 = reg_0676;
    71: op1_04_in16 = reg_0960;
    72: op1_04_in16 = reg_0867;
    73: op1_04_in16 = reg_0990;
    74: op1_04_in16 = reg_0893;
    75: op1_04_in16 = imem06_in[59:56];
    78: op1_04_in16 = reg_0190;
    79: op1_04_in16 = reg_0233;
    80: op1_04_in16 = reg_0809;
    81: op1_04_in16 = reg_0952;
    82: op1_04_in16 = reg_0137;
    83: op1_04_in16 = reg_0213;
    84: op1_04_in16 = reg_0731;
    85: op1_04_in16 = imem04_in[43:40];
    86: op1_04_in16 = reg_0328;
    87: op1_04_in16 = imem02_in[59:56];
    88: op1_04_in16 = reg_0656;
    89: op1_04_in16 = imem07_in[31:28];
    90: op1_04_in16 = reg_0752;
    91: op1_04_in16 = imem05_in[7:4];
    92: op1_04_in16 = imem05_in[51:48];
    97: op1_04_in16 = reg_1011;
    default: op1_04_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv16 = 1;
    8: op1_04_inv16 = 1;
    9: op1_04_inv16 = 1;
    10: op1_04_inv16 = 1;
    11: op1_04_inv16 = 1;
    12: op1_04_inv16 = 1;
    13: op1_04_inv16 = 1;
    15: op1_04_inv16 = 1;
    16: op1_04_inv16 = 1;
    17: op1_04_inv16 = 1;
    19: op1_04_inv16 = 1;
    21: op1_04_inv16 = 1;
    23: op1_04_inv16 = 1;
    26: op1_04_inv16 = 1;
    28: op1_04_inv16 = 1;
    29: op1_04_inv16 = 1;
    30: op1_04_inv16 = 1;
    31: op1_04_inv16 = 1;
    34: op1_04_inv16 = 1;
    35: op1_04_inv16 = 1;
    36: op1_04_inv16 = 1;
    37: op1_04_inv16 = 1;
    38: op1_04_inv16 = 1;
    43: op1_04_inv16 = 1;
    46: op1_04_inv16 = 1;
    47: op1_04_inv16 = 1;
    51: op1_04_inv16 = 1;
    57: op1_04_inv16 = 1;
    58: op1_04_inv16 = 1;
    59: op1_04_inv16 = 1;
    63: op1_04_inv16 = 1;
    64: op1_04_inv16 = 1;
    66: op1_04_inv16 = 1;
    68: op1_04_inv16 = 1;
    71: op1_04_inv16 = 1;
    72: op1_04_inv16 = 1;
    73: op1_04_inv16 = 1;
    75: op1_04_inv16 = 1;
    79: op1_04_inv16 = 1;
    83: op1_04_inv16 = 1;
    84: op1_04_inv16 = 1;
    86: op1_04_inv16 = 1;
    89: op1_04_inv16 = 1;
    91: op1_04_inv16 = 1;
    92: op1_04_inv16 = 1;
    default: op1_04_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in17 = reg_0168;
    6: op1_04_in17 = reg_0269;
    7: op1_04_in17 = reg_0203;
    8: op1_04_in17 = reg_0068;
    9: op1_04_in17 = reg_0408;
    10: op1_04_in17 = reg_0148;
    11: op1_04_in17 = reg_0711;
    12: op1_04_in17 = imem06_in[3:0];
    13: op1_04_in17 = reg_0869;
    14: op1_04_in17 = reg_0283;
    15: op1_04_in17 = reg_0405;
    16: op1_04_in17 = reg_0187;
    48: op1_04_in17 = reg_0187;
    17: op1_04_in17 = imem03_in[3:0];
    18: op1_04_in17 = reg_0715;
    19: op1_04_in17 = reg_0776;
    20: op1_04_in17 = reg_0349;
    21: op1_04_in17 = reg_0573;
    22: op1_04_in17 = reg_0617;
    23: op1_04_in17 = reg_0424;
    24: op1_04_in17 = reg_0955;
    25: op1_04_in17 = reg_0200;
    26: op1_04_in17 = imem03_in[23:20];
    27: op1_04_in17 = reg_1039;
    28: op1_04_in17 = reg_0656;
    29: op1_04_in17 = reg_0802;
    59: op1_04_in17 = reg_0802;
    30: op1_04_in17 = reg_0158;
    31: op1_04_in17 = reg_0663;
    32: op1_04_in17 = reg_0964;
    33: op1_04_in17 = imem07_in[123:120];
    34: op1_04_in17 = reg_0274;
    35: op1_04_in17 = reg_0383;
    36: op1_04_in17 = reg_0947;
    37: op1_04_in17 = imem06_in[15:12];
    86: op1_04_in17 = imem06_in[15:12];
    38: op1_04_in17 = reg_0029;
    40: op1_04_in17 = reg_0228;
    42: op1_04_in17 = reg_0063;
    43: op1_04_in17 = reg_0407;
    74: op1_04_in17 = reg_0407;
    45: op1_04_in17 = reg_0097;
    46: op1_04_in17 = reg_0932;
    47: op1_04_in17 = reg_0169;
    49: op1_04_in17 = imem05_in[27:24];
    50: op1_04_in17 = reg_0576;
    51: op1_04_in17 = reg_0651;
    53: op1_04_in17 = reg_0828;
    54: op1_04_in17 = reg_0389;
    55: op1_04_in17 = imem03_in[59:56];
    56: op1_04_in17 = imem04_in[23:20];
    57: op1_04_in17 = reg_0688;
    58: op1_04_in17 = reg_0691;
    61: op1_04_in17 = imem06_in[71:68];
    63: op1_04_in17 = reg_0739;
    64: op1_04_in17 = imem03_in[79:76];
    65: op1_04_in17 = reg_0584;
    66: op1_04_in17 = reg_0494;
    67: op1_04_in17 = imem04_in[7:4];
    68: op1_04_in17 = reg_0142;
    69: op1_04_in17 = reg_0206;
    70: op1_04_in17 = reg_0099;
    71: op1_04_in17 = reg_0143;
    72: op1_04_in17 = reg_0085;
    73: op1_04_in17 = reg_0983;
    75: op1_04_in17 = imem06_in[87:84];
    78: op1_04_in17 = imem01_in[39:36];
    79: op1_04_in17 = reg_0979;
    80: op1_04_in17 = reg_0065;
    81: op1_04_in17 = reg_0508;
    82: op1_04_in17 = reg_0107;
    83: op1_04_in17 = imem01_in[43:40];
    84: op1_04_in17 = reg_0703;
    85: op1_04_in17 = imem04_in[91:88];
    87: op1_04_in17 = reg_0666;
    88: op1_04_in17 = reg_0082;
    89: op1_04_in17 = imem07_in[51:48];
    90: op1_04_in17 = reg_0276;
    91: op1_04_in17 = imem05_in[59:56];
    92: op1_04_in17 = imem05_in[103:100];
    97: op1_04_in17 = reg_0229;
    default: op1_04_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv17 = 1;
    8: op1_04_inv17 = 1;
    9: op1_04_inv17 = 1;
    11: op1_04_inv17 = 1;
    14: op1_04_inv17 = 1;
    16: op1_04_inv17 = 1;
    17: op1_04_inv17 = 1;
    19: op1_04_inv17 = 1;
    22: op1_04_inv17 = 1;
    24: op1_04_inv17 = 1;
    25: op1_04_inv17 = 1;
    27: op1_04_inv17 = 1;
    28: op1_04_inv17 = 1;
    31: op1_04_inv17 = 1;
    34: op1_04_inv17 = 1;
    35: op1_04_inv17 = 1;
    40: op1_04_inv17 = 1;
    45: op1_04_inv17 = 1;
    47: op1_04_inv17 = 1;
    48: op1_04_inv17 = 1;
    49: op1_04_inv17 = 1;
    51: op1_04_inv17 = 1;
    54: op1_04_inv17 = 1;
    55: op1_04_inv17 = 1;
    56: op1_04_inv17 = 1;
    57: op1_04_inv17 = 1;
    58: op1_04_inv17 = 1;
    63: op1_04_inv17 = 1;
    64: op1_04_inv17 = 1;
    66: op1_04_inv17 = 1;
    69: op1_04_inv17 = 1;
    75: op1_04_inv17 = 1;
    79: op1_04_inv17 = 1;
    82: op1_04_inv17 = 1;
    83: op1_04_inv17 = 1;
    86: op1_04_inv17 = 1;
    89: op1_04_inv17 = 1;
    90: op1_04_inv17 = 1;
    92: op1_04_inv17 = 1;
    97: op1_04_inv17 = 1;
    default: op1_04_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の18番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in18 = reg_0244;
    7: op1_04_in18 = reg_0186;
    8: op1_04_in18 = reg_0075;
    9: op1_04_in18 = reg_0392;
    10: op1_04_in18 = reg_0145;
    11: op1_04_in18 = reg_0424;
    12: op1_04_in18 = imem06_in[7:4];
    13: op1_04_in18 = reg_0228;
    64: op1_04_in18 = reg_0228;
    70: op1_04_in18 = reg_0228;
    14: op1_04_in18 = reg_0279;
    15: op1_04_in18 = reg_0375;
    20: op1_04_in18 = reg_0375;
    16: op1_04_in18 = reg_0193;
    17: op1_04_in18 = imem03_in[19:16];
    18: op1_04_in18 = reg_0707;
    19: op1_04_in18 = reg_0048;
    21: op1_04_in18 = reg_0568;
    22: op1_04_in18 = reg_0605;
    23: op1_04_in18 = reg_0430;
    24: op1_04_in18 = reg_0826;
    25: op1_04_in18 = reg_0204;
    48: op1_04_in18 = reg_0204;
    26: op1_04_in18 = imem03_in[47:44];
    27: op1_04_in18 = reg_1032;
    34: op1_04_in18 = reg_1032;
    28: op1_04_in18 = reg_0651;
    29: op1_04_in18 = imem07_in[23:20];
    38: op1_04_in18 = imem07_in[23:20];
    31: op1_04_in18 = reg_0086;
    72: op1_04_in18 = reg_0086;
    32: op1_04_in18 = reg_0900;
    33: op1_04_in18 = reg_0719;
    35: op1_04_in18 = reg_0222;
    36: op1_04_in18 = reg_0960;
    37: op1_04_in18 = imem06_in[63:60];
    40: op1_04_in18 = reg_1018;
    42: op1_04_in18 = reg_0579;
    43: op1_04_in18 = reg_0020;
    45: op1_04_in18 = reg_0318;
    46: op1_04_in18 = reg_0752;
    47: op1_04_in18 = reg_0163;
    49: op1_04_in18 = imem05_in[43:40];
    50: op1_04_in18 = reg_0923;
    55: op1_04_in18 = reg_0923;
    89: op1_04_in18 = reg_0923;
    51: op1_04_in18 = reg_0026;
    53: op1_04_in18 = reg_0913;
    54: op1_04_in18 = reg_0425;
    56: op1_04_in18 = imem04_in[35:32];
    57: op1_04_in18 = reg_0689;
    58: op1_04_in18 = reg_0351;
    59: op1_04_in18 = reg_0067;
    61: op1_04_in18 = imem07_in[19:16];
    63: op1_04_in18 = reg_0389;
    65: op1_04_in18 = reg_0015;
    66: op1_04_in18 = reg_0027;
    67: op1_04_in18 = imem04_in[51:48];
    68: op1_04_in18 = reg_0146;
    81: op1_04_in18 = reg_0146;
    69: op1_04_in18 = reg_0199;
    71: op1_04_in18 = reg_0139;
    73: op1_04_in18 = imem04_in[7:4];
    74: op1_04_in18 = reg_0658;
    75: op1_04_in18 = reg_0626;
    78: op1_04_in18 = imem01_in[55:52];
    83: op1_04_in18 = imem01_in[55:52];
    79: op1_04_in18 = reg_0996;
    80: op1_04_in18 = reg_0071;
    82: op1_04_in18 = reg_0967;
    84: op1_04_in18 = reg_0447;
    85: op1_04_in18 = imem04_in[95:92];
    86: op1_04_in18 = imem06_in[23:20];
    87: op1_04_in18 = reg_0285;
    88: op1_04_in18 = reg_0874;
    90: op1_04_in18 = reg_0284;
    91: op1_04_in18 = imem05_in[63:60];
    92: op1_04_in18 = reg_0944;
    97: op1_04_in18 = reg_0814;
    default: op1_04_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv18 = 1;
    9: op1_04_inv18 = 1;
    10: op1_04_inv18 = 1;
    13: op1_04_inv18 = 1;
    17: op1_04_inv18 = 1;
    19: op1_04_inv18 = 1;
    22: op1_04_inv18 = 1;
    27: op1_04_inv18 = 1;
    35: op1_04_inv18 = 1;
    38: op1_04_inv18 = 1;
    43: op1_04_inv18 = 1;
    46: op1_04_inv18 = 1;
    49: op1_04_inv18 = 1;
    50: op1_04_inv18 = 1;
    54: op1_04_inv18 = 1;
    57: op1_04_inv18 = 1;
    58: op1_04_inv18 = 1;
    59: op1_04_inv18 = 1;
    61: op1_04_inv18 = 1;
    63: op1_04_inv18 = 1;
    64: op1_04_inv18 = 1;
    66: op1_04_inv18 = 1;
    71: op1_04_inv18 = 1;
    72: op1_04_inv18 = 1;
    73: op1_04_inv18 = 1;
    75: op1_04_inv18 = 1;
    78: op1_04_inv18 = 1;
    81: op1_04_inv18 = 1;
    82: op1_04_inv18 = 1;
    83: op1_04_inv18 = 1;
    87: op1_04_inv18 = 1;
    92: op1_04_inv18 = 1;
    97: op1_04_inv18 = 1;
    default: op1_04_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の19番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in19 = reg_0263;
    7: op1_04_in19 = reg_0212;
    16: op1_04_in19 = reg_0212;
    8: op1_04_in19 = reg_0044;
    9: op1_04_in19 = reg_0409;
    10: op1_04_in19 = reg_0136;
    11: op1_04_in19 = reg_0429;
    23: op1_04_in19 = reg_0429;
    12: op1_04_in19 = imem06_in[43:40];
    13: op1_04_in19 = reg_0124;
    14: op1_04_in19 = reg_0300;
    51: op1_04_in19 = reg_0300;
    15: op1_04_in19 = reg_0383;
    17: op1_04_in19 = imem03_in[35:32];
    18: op1_04_in19 = reg_0436;
    19: op1_04_in19 = reg_0892;
    20: op1_04_in19 = reg_0406;
    21: op1_04_in19 = reg_0592;
    22: op1_04_in19 = reg_0632;
    24: op1_04_in19 = reg_0806;
    25: op1_04_in19 = reg_0207;
    26: op1_04_in19 = imem03_in[71:68];
    27: op1_04_in19 = reg_0869;
    28: op1_04_in19 = reg_0649;
    29: op1_04_in19 = imem07_in[71:68];
    31: op1_04_in19 = reg_0310;
    32: op1_04_in19 = reg_0757;
    33: op1_04_in19 = reg_0717;
    34: op1_04_in19 = reg_0830;
    35: op1_04_in19 = reg_0594;
    36: op1_04_in19 = reg_0022;
    37: op1_04_in19 = imem06_in[75:72];
    38: op1_04_in19 = imem07_in[75:72];
    40: op1_04_in19 = reg_1034;
    42: op1_04_in19 = reg_0347;
    54: op1_04_in19 = reg_0347;
    43: op1_04_in19 = reg_0371;
    45: op1_04_in19 = reg_0886;
    46: op1_04_in19 = reg_0524;
    47: op1_04_in19 = reg_0178;
    48: op1_04_in19 = reg_0188;
    49: op1_04_in19 = imem05_in[51:48];
    50: op1_04_in19 = reg_0051;
    53: op1_04_in19 = reg_0240;
    55: op1_04_in19 = reg_0793;
    56: op1_04_in19 = imem04_in[91:88];
    57: op1_04_in19 = reg_0057;
    58: op1_04_in19 = reg_0025;
    59: op1_04_in19 = reg_0068;
    61: op1_04_in19 = imem07_in[27:24];
    63: op1_04_in19 = reg_0425;
    64: op1_04_in19 = reg_0585;
    65: op1_04_in19 = reg_0407;
    66: op1_04_in19 = reg_0108;
    67: op1_04_in19 = imem04_in[55:52];
    68: op1_04_in19 = reg_0129;
    69: op1_04_in19 = reg_0192;
    70: op1_04_in19 = reg_0580;
    71: op1_04_in19 = reg_0153;
    72: op1_04_in19 = reg_0084;
    73: op1_04_in19 = imem04_in[19:16];
    74: op1_04_in19 = reg_0494;
    90: op1_04_in19 = reg_0494;
    75: op1_04_in19 = reg_0754;
    78: op1_04_in19 = imem01_in[115:112];
    79: op1_04_in19 = reg_0994;
    80: op1_04_in19 = reg_0824;
    81: op1_04_in19 = reg_0816;
    82: op1_04_in19 = reg_1015;
    83: op1_04_in19 = imem01_in[63:60];
    84: op1_04_in19 = reg_0339;
    85: op1_04_in19 = imem04_in[119:116];
    86: op1_04_in19 = imem06_in[63:60];
    87: op1_04_in19 = reg_0605;
    88: op1_04_in19 = reg_0613;
    89: op1_04_in19 = reg_0959;
    91: op1_04_in19 = imem05_in[99:96];
    92: op1_04_in19 = reg_0954;
    97: op1_04_in19 = reg_0698;
    default: op1_04_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_04_inv19 = 1;
    10: op1_04_inv19 = 1;
    11: op1_04_inv19 = 1;
    13: op1_04_inv19 = 1;
    15: op1_04_inv19 = 1;
    16: op1_04_inv19 = 1;
    17: op1_04_inv19 = 1;
    20: op1_04_inv19 = 1;
    21: op1_04_inv19 = 1;
    22: op1_04_inv19 = 1;
    23: op1_04_inv19 = 1;
    25: op1_04_inv19 = 1;
    26: op1_04_inv19 = 1;
    35: op1_04_inv19 = 1;
    36: op1_04_inv19 = 1;
    37: op1_04_inv19 = 1;
    43: op1_04_inv19 = 1;
    46: op1_04_inv19 = 1;
    47: op1_04_inv19 = 1;
    49: op1_04_inv19 = 1;
    51: op1_04_inv19 = 1;
    58: op1_04_inv19 = 1;
    59: op1_04_inv19 = 1;
    63: op1_04_inv19 = 1;
    64: op1_04_inv19 = 1;
    67: op1_04_inv19 = 1;
    68: op1_04_inv19 = 1;
    70: op1_04_inv19 = 1;
    71: op1_04_inv19 = 1;
    73: op1_04_inv19 = 1;
    75: op1_04_inv19 = 1;
    80: op1_04_inv19 = 1;
    85: op1_04_inv19 = 1;
    87: op1_04_inv19 = 1;
    88: op1_04_inv19 = 1;
    89: op1_04_inv19 = 1;
    90: op1_04_inv19 = 1;
    91: op1_04_inv19 = 1;
    92: op1_04_inv19 = 1;
    97: op1_04_inv19 = 1;
    default: op1_04_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の20番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in20 = reg_0145;
    7: op1_04_in20 = reg_0197;
    69: op1_04_in20 = reg_0197;
    8: op1_04_in20 = imem05_in[3:0];
    9: op1_04_in20 = reg_0371;
    10: op1_04_in20 = reg_0128;
    11: op1_04_in20 = reg_0423;
    12: op1_04_in20 = imem06_in[47:44];
    13: op1_04_in20 = reg_0125;
    14: op1_04_in20 = reg_0295;
    15: op1_04_in20 = reg_0404;
    16: op1_04_in20 = reg_0202;
    17: op1_04_in20 = imem03_in[55:52];
    18: op1_04_in20 = reg_0419;
    19: op1_04_in20 = reg_0484;
    20: op1_04_in20 = reg_0787;
    21: op1_04_in20 = reg_0591;
    22: op1_04_in20 = reg_0386;
    23: op1_04_in20 = reg_0443;
    24: op1_04_in20 = reg_0251;
    25: op1_04_in20 = reg_0918;
    26: op1_04_in20 = imem03_in[87:84];
    27: op1_04_in20 = reg_0885;
    28: op1_04_in20 = reg_0095;
    29: op1_04_in20 = imem07_in[111:108];
    31: op1_04_in20 = reg_0502;
    32: op1_04_in20 = reg_0813;
    33: op1_04_in20 = reg_0706;
    34: op1_04_in20 = reg_1037;
    35: op1_04_in20 = reg_0405;
    36: op1_04_in20 = reg_0491;
    37: op1_04_in20 = imem06_in[83:80];
    38: op1_04_in20 = imem07_in[95:92];
    40: op1_04_in20 = reg_0013;
    42: op1_04_in20 = reg_0307;
    43: op1_04_in20 = reg_0781;
    45: op1_04_in20 = reg_0865;
    46: op1_04_in20 = imem04_in[39:36];
    47: op1_04_in20 = reg_0173;
    48: op1_04_in20 = reg_0193;
    49: op1_04_in20 = imem05_in[95:92];
    50: op1_04_in20 = reg_0312;
    51: op1_04_in20 = reg_0636;
    53: op1_04_in20 = reg_0905;
    54: op1_04_in20 = reg_0007;
    55: op1_04_in20 = reg_0833;
    56: op1_04_in20 = imem04_in[107:104];
    57: op1_04_in20 = reg_0233;
    58: op1_04_in20 = reg_0626;
    59: op1_04_in20 = reg_0815;
    61: op1_04_in20 = imem07_in[55:52];
    63: op1_04_in20 = reg_0085;
    64: op1_04_in20 = reg_0547;
    70: op1_04_in20 = reg_0547;
    65: op1_04_in20 = reg_0444;
    66: op1_04_in20 = reg_0332;
    67: op1_04_in20 = imem04_in[59:56];
    68: op1_04_in20 = reg_0130;
    71: op1_04_in20 = reg_0141;
    72: op1_04_in20 = imem03_in[15:12];
    73: op1_04_in20 = imem04_in[67:64];
    74: op1_04_in20 = reg_0854;
    75: op1_04_in20 = reg_0384;
    78: op1_04_in20 = reg_0122;
    79: op1_04_in20 = imem04_in[51:48];
    80: op1_04_in20 = reg_0542;
    81: op1_04_in20 = imem06_in[71:68];
    82: op1_04_in20 = reg_0223;
    83: op1_04_in20 = imem01_in[71:68];
    84: op1_04_in20 = reg_0184;
    85: op1_04_in20 = reg_0126;
    86: op1_04_in20 = imem06_in[111:108];
    87: op1_04_in20 = reg_0069;
    88: op1_04_in20 = reg_0961;
    89: op1_04_in20 = reg_0718;
    90: op1_04_in20 = imem05_in[55:52];
    91: op1_04_in20 = reg_0140;
    92: op1_04_in20 = reg_0275;
    97: op1_04_in20 = reg_0783;
    default: op1_04_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv20 = 1;
    13: op1_04_inv20 = 1;
    14: op1_04_inv20 = 1;
    15: op1_04_inv20 = 1;
    16: op1_04_inv20 = 1;
    17: op1_04_inv20 = 1;
    18: op1_04_inv20 = 1;
    20: op1_04_inv20 = 1;
    22: op1_04_inv20 = 1;
    25: op1_04_inv20 = 1;
    27: op1_04_inv20 = 1;
    32: op1_04_inv20 = 1;
    34: op1_04_inv20 = 1;
    36: op1_04_inv20 = 1;
    37: op1_04_inv20 = 1;
    42: op1_04_inv20 = 1;
    49: op1_04_inv20 = 1;
    53: op1_04_inv20 = 1;
    54: op1_04_inv20 = 1;
    55: op1_04_inv20 = 1;
    59: op1_04_inv20 = 1;
    61: op1_04_inv20 = 1;
    63: op1_04_inv20 = 1;
    65: op1_04_inv20 = 1;
    71: op1_04_inv20 = 1;
    73: op1_04_inv20 = 1;
    74: op1_04_inv20 = 1;
    75: op1_04_inv20 = 1;
    79: op1_04_inv20 = 1;
    80: op1_04_inv20 = 1;
    81: op1_04_inv20 = 1;
    82: op1_04_inv20 = 1;
    83: op1_04_inv20 = 1;
    89: op1_04_inv20 = 1;
    90: op1_04_inv20 = 1;
    91: op1_04_inv20 = 1;
    92: op1_04_inv20 = 1;
    default: op1_04_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の21番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in21 = reg_0140;
    71: op1_04_in21 = reg_0140;
    7: op1_04_in21 = imem01_in[107:104];
    8: op1_04_in21 = imem05_in[15:12];
    9: op1_04_in21 = reg_0382;
    10: op1_04_in21 = reg_0142;
    11: op1_04_in21 = reg_0439;
    12: op1_04_in21 = imem06_in[71:68];
    13: op1_04_in21 = reg_0102;
    14: op1_04_in21 = reg_0065;
    15: op1_04_in21 = reg_0315;
    16: op1_04_in21 = imem01_in[11:8];
    17: op1_04_in21 = imem03_in[83:80];
    18: op1_04_in21 = reg_0431;
    19: op1_04_in21 = reg_0876;
    20: op1_04_in21 = reg_0783;
    21: op1_04_in21 = reg_0580;
    22: op1_04_in21 = reg_0399;
    23: op1_04_in21 = reg_0175;
    24: op1_04_in21 = reg_0275;
    25: op1_04_in21 = reg_0532;
    26: op1_04_in21 = imem03_in[91:88];
    27: op1_04_in21 = reg_0830;
    28: op1_04_in21 = reg_0330;
    29: op1_04_in21 = imem07_in[119:116];
    31: op1_04_in21 = reg_0321;
    32: op1_04_in21 = reg_0832;
    33: op1_04_in21 = reg_0700;
    34: op1_04_in21 = reg_1031;
    35: op1_04_in21 = reg_0596;
    36: op1_04_in21 = reg_0260;
    37: op1_04_in21 = imem06_in[95:92];
    38: op1_04_in21 = imem07_in[99:96];
    40: op1_04_in21 = reg_0786;
    42: op1_04_in21 = reg_0301;
    43: op1_04_in21 = reg_0356;
    45: op1_04_in21 = reg_0817;
    46: op1_04_in21 = imem04_in[91:88];
    48: op1_04_in21 = reg_0199;
    49: op1_04_in21 = imem05_in[99:96];
    50: op1_04_in21 = reg_0998;
    51: op1_04_in21 = reg_0097;
    53: op1_04_in21 = reg_0779;
    54: op1_04_in21 = reg_0085;
    55: op1_04_in21 = reg_0795;
    56: op1_04_in21 = imem04_in[119:116];
    57: op1_04_in21 = reg_0032;
    58: op1_04_in21 = reg_0926;
    59: op1_04_in21 = reg_0072;
    61: op1_04_in21 = imem07_in[75:72];
    63: op1_04_in21 = reg_0261;
    64: op1_04_in21 = reg_0298;
    65: op1_04_in21 = reg_0041;
    66: op1_04_in21 = reg_0652;
    67: op1_04_in21 = imem04_in[107:104];
    68: op1_04_in21 = reg_0131;
    69: op1_04_in21 = reg_0918;
    70: op1_04_in21 = reg_0576;
    72: op1_04_in21 = imem03_in[43:40];
    73: op1_04_in21 = imem04_in[75:72];
    74: op1_04_in21 = reg_0824;
    75: op1_04_in21 = reg_0534;
    78: op1_04_in21 = reg_0488;
    79: op1_04_in21 = imem04_in[59:56];
    80: op1_04_in21 = reg_0332;
    81: op1_04_in21 = imem06_in[75:72];
    82: op1_04_in21 = reg_0952;
    83: op1_04_in21 = reg_1023;
    85: op1_04_in21 = reg_0430;
    86: op1_04_in21 = imem06_in[123:120];
    87: op1_04_in21 = reg_0348;
    88: op1_04_in21 = imem03_in[7:4];
    89: op1_04_in21 = reg_0563;
    90: op1_04_in21 = imem05_in[75:72];
    91: op1_04_in21 = reg_0689;
    92: op1_04_in21 = reg_0013;
    97: op1_04_in21 = reg_0011;
    default: op1_04_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv21 = 1;
    9: op1_04_inv21 = 1;
    10: op1_04_inv21 = 1;
    11: op1_04_inv21 = 1;
    13: op1_04_inv21 = 1;
    14: op1_04_inv21 = 1;
    15: op1_04_inv21 = 1;
    16: op1_04_inv21 = 1;
    17: op1_04_inv21 = 1;
    18: op1_04_inv21 = 1;
    19: op1_04_inv21 = 1;
    21: op1_04_inv21 = 1;
    24: op1_04_inv21 = 1;
    25: op1_04_inv21 = 1;
    26: op1_04_inv21 = 1;
    28: op1_04_inv21 = 1;
    31: op1_04_inv21 = 1;
    33: op1_04_inv21 = 1;
    35: op1_04_inv21 = 1;
    38: op1_04_inv21 = 1;
    40: op1_04_inv21 = 1;
    45: op1_04_inv21 = 1;
    46: op1_04_inv21 = 1;
    50: op1_04_inv21 = 1;
    54: op1_04_inv21 = 1;
    56: op1_04_inv21 = 1;
    57: op1_04_inv21 = 1;
    59: op1_04_inv21 = 1;
    61: op1_04_inv21 = 1;
    64: op1_04_inv21 = 1;
    65: op1_04_inv21 = 1;
    69: op1_04_inv21 = 1;
    72: op1_04_inv21 = 1;
    75: op1_04_inv21 = 1;
    78: op1_04_inv21 = 1;
    79: op1_04_inv21 = 1;
    81: op1_04_inv21 = 1;
    83: op1_04_inv21 = 1;
    85: op1_04_inv21 = 1;
    88: op1_04_inv21 = 1;
    89: op1_04_inv21 = 1;
    90: op1_04_inv21 = 1;
    92: op1_04_inv21 = 1;
    default: op1_04_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の22番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in22 = imem06_in[47:44];
    7: op1_04_in22 = imem01_in[111:108];
    8: op1_04_in22 = imem05_in[75:72];
    9: op1_04_in22 = reg_0380;
    10: op1_04_in22 = reg_0146;
    11: op1_04_in22 = reg_0435;
    12: op1_04_in22 = imem06_in[79:76];
    13: op1_04_in22 = reg_0114;
    14: op1_04_in22 = reg_0056;
    15: op1_04_in22 = reg_0390;
    16: op1_04_in22 = imem01_in[23:20];
    17: op1_04_in22 = reg_0582;
    18: op1_04_in22 = reg_0172;
    19: op1_04_in22 = reg_0543;
    20: op1_04_in22 = imem07_in[11:8];
    21: op1_04_in22 = reg_0595;
    22: op1_04_in22 = reg_0027;
    23: op1_04_in22 = reg_0167;
    24: op1_04_in22 = reg_0260;
    25: op1_04_in22 = reg_0775;
    26: op1_04_in22 = imem03_in[95:92];
    27: op1_04_in22 = reg_0216;
    28: op1_04_in22 = reg_0886;
    29: op1_04_in22 = reg_0719;
    31: op1_04_in22 = reg_0568;
    32: op1_04_in22 = reg_0819;
    33: op1_04_in22 = reg_0432;
    34: op1_04_in22 = reg_0913;
    35: op1_04_in22 = reg_0029;
    36: op1_04_in22 = reg_0832;
    37: op1_04_in22 = imem06_in[99:96];
    38: op1_04_in22 = reg_0728;
    40: op1_04_in22 = reg_0779;
    42: op1_04_in22 = reg_0530;
    43: op1_04_in22 = reg_0914;
    45: op1_04_in22 = reg_0083;
    46: op1_04_in22 = imem04_in[103:100];
    48: op1_04_in22 = reg_0597;
    49: op1_04_in22 = reg_0944;
    50: op1_04_in22 = reg_0986;
    51: op1_04_in22 = reg_0318;
    53: op1_04_in22 = reg_1034;
    54: op1_04_in22 = reg_0009;
    55: op1_04_in22 = reg_0784;
    56: op1_04_in22 = imem04_in[127:124];
    57: op1_04_in22 = reg_0488;
    58: op1_04_in22 = reg_0229;
    59: op1_04_in22 = imem04_in[87:84];
    61: op1_04_in22 = imem07_in[91:88];
    63: op1_04_in22 = reg_0077;
    64: op1_04_in22 = reg_0346;
    65: op1_04_in22 = reg_0071;
    66: op1_04_in22 = reg_0314;
    67: op1_04_in22 = reg_0265;
    68: op1_04_in22 = imem06_in[55:52];
    69: op1_04_in22 = reg_0490;
    70: op1_04_in22 = imem03_in[23:20];
    71: op1_04_in22 = reg_0137;
    72: op1_04_in22 = imem03_in[107:104];
    73: op1_04_in22 = imem04_in[79:76];
    74: op1_04_in22 = reg_0332;
    75: op1_04_in22 = reg_0297;
    78: op1_04_in22 = reg_1022;
    79: op1_04_in22 = imem04_in[63:60];
    80: op1_04_in22 = reg_0531;
    81: op1_04_in22 = imem06_in[83:80];
    82: op1_04_in22 = reg_0957;
    83: op1_04_in22 = reg_1035;
    85: op1_04_in22 = reg_1005;
    86: op1_04_in22 = imem06_in[127:124];
    87: op1_04_in22 = reg_0483;
    88: op1_04_in22 = imem03_in[19:16];
    89: op1_04_in22 = reg_0759;
    90: op1_04_in22 = imem05_in[83:80];
    91: op1_04_in22 = reg_0057;
    92: op1_04_in22 = reg_0269;
    97: op1_04_in22 = reg_1029;
    default: op1_04_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_04_inv22 = 1;
    13: op1_04_inv22 = 1;
    14: op1_04_inv22 = 1;
    16: op1_04_inv22 = 1;
    19: op1_04_inv22 = 1;
    21: op1_04_inv22 = 1;
    22: op1_04_inv22 = 1;
    25: op1_04_inv22 = 1;
    29: op1_04_inv22 = 1;
    34: op1_04_inv22 = 1;
    35: op1_04_inv22 = 1;
    36: op1_04_inv22 = 1;
    37: op1_04_inv22 = 1;
    40: op1_04_inv22 = 1;
    46: op1_04_inv22 = 1;
    48: op1_04_inv22 = 1;
    50: op1_04_inv22 = 1;
    51: op1_04_inv22 = 1;
    53: op1_04_inv22 = 1;
    55: op1_04_inv22 = 1;
    56: op1_04_inv22 = 1;
    58: op1_04_inv22 = 1;
    59: op1_04_inv22 = 1;
    61: op1_04_inv22 = 1;
    63: op1_04_inv22 = 1;
    67: op1_04_inv22 = 1;
    68: op1_04_inv22 = 1;
    69: op1_04_inv22 = 1;
    70: op1_04_inv22 = 1;
    73: op1_04_inv22 = 1;
    78: op1_04_inv22 = 1;
    81: op1_04_inv22 = 1;
    82: op1_04_inv22 = 1;
    83: op1_04_inv22 = 1;
    85: op1_04_inv22 = 1;
    87: op1_04_inv22 = 1;
    89: op1_04_inv22 = 1;
    90: op1_04_inv22 = 1;
    97: op1_04_inv22 = 1;
    default: op1_04_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の23番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in23 = imem06_in[67:64];
    7: op1_04_in23 = reg_0499;
    8: op1_04_in23 = imem05_in[83:80];
    9: op1_04_in23 = imem06_in[71:68];
    10: op1_04_in23 = reg_0139;
    11: op1_04_in23 = reg_0175;
    12: op1_04_in23 = imem06_in[83:80];
    13: op1_04_in23 = reg_0107;
    14: op1_04_in23 = reg_0064;
    15: op1_04_in23 = reg_0799;
    16: op1_04_in23 = imem01_in[83:80];
    17: op1_04_in23 = reg_0573;
    19: op1_04_in23 = reg_0536;
    20: op1_04_in23 = imem07_in[31:28];
    21: op1_04_in23 = reg_0576;
    22: op1_04_in23 = imem07_in[55:52];
    23: op1_04_in23 = reg_0160;
    24: op1_04_in23 = reg_0896;
    25: op1_04_in23 = reg_0925;
    26: op1_04_in23 = reg_0583;
    91: op1_04_in23 = reg_0583;
    27: op1_04_in23 = reg_1040;
    28: op1_04_in23 = reg_0516;
    29: op1_04_in23 = reg_0731;
    31: op1_04_in23 = reg_0569;
    32: op1_04_in23 = reg_0831;
    78: op1_04_in23 = reg_0831;
    33: op1_04_in23 = reg_0439;
    34: op1_04_in23 = reg_1036;
    35: op1_04_in23 = reg_0595;
    36: op1_04_in23 = reg_0819;
    37: op1_04_in23 = imem06_in[103:100];
    38: op1_04_in23 = reg_0719;
    40: op1_04_in23 = reg_0563;
    42: op1_04_in23 = reg_0265;
    43: op1_04_in23 = reg_0382;
    75: op1_04_in23 = reg_0382;
    45: op1_04_in23 = reg_0776;
    46: op1_04_in23 = imem05_in[7:4];
    80: op1_04_in23 = imem05_in[7:4];
    48: op1_04_in23 = reg_0849;
    69: op1_04_in23 = reg_0849;
    49: op1_04_in23 = reg_0969;
    50: op1_04_in23 = reg_0980;
    51: op1_04_in23 = reg_0330;
    53: op1_04_in23 = reg_1043;
    54: op1_04_in23 = reg_0743;
    55: op1_04_in23 = reg_0513;
    56: op1_04_in23 = reg_0483;
    57: op1_04_in23 = reg_0252;
    58: op1_04_in23 = imem06_in[59:56];
    59: op1_04_in23 = imem04_in[95:92];
    73: op1_04_in23 = imem04_in[95:92];
    61: op1_04_in23 = imem07_in[127:124];
    63: op1_04_in23 = reg_0291;
    64: op1_04_in23 = reg_0823;
    65: op1_04_in23 = reg_0332;
    66: op1_04_in23 = reg_0782;
    67: op1_04_in23 = reg_0055;
    68: op1_04_in23 = imem06_in[99:96];
    81: op1_04_in23 = imem06_in[99:96];
    70: op1_04_in23 = imem03_in[31:28];
    71: op1_04_in23 = reg_0118;
    72: op1_04_in23 = reg_0012;
    74: op1_04_in23 = reg_0044;
    79: op1_04_in23 = imem04_in[67:64];
    82: op1_04_in23 = reg_0943;
    83: op1_04_in23 = reg_1024;
    85: op1_04_in23 = reg_0296;
    86: op1_04_in23 = reg_0032;
    87: op1_04_in23 = reg_0765;
    88: op1_04_in23 = imem03_in[35:32];
    89: op1_04_in23 = reg_0002;
    90: op1_04_in23 = imem05_in[87:84];
    92: op1_04_in23 = reg_0256;
    97: op1_04_in23 = reg_0133;
    default: op1_04_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv23 = 1;
    8: op1_04_inv23 = 1;
    9: op1_04_inv23 = 1;
    10: op1_04_inv23 = 1;
    12: op1_04_inv23 = 1;
    13: op1_04_inv23 = 1;
    14: op1_04_inv23 = 1;
    22: op1_04_inv23 = 1;
    25: op1_04_inv23 = 1;
    26: op1_04_inv23 = 1;
    27: op1_04_inv23 = 1;
    28: op1_04_inv23 = 1;
    31: op1_04_inv23 = 1;
    34: op1_04_inv23 = 1;
    36: op1_04_inv23 = 1;
    40: op1_04_inv23 = 1;
    42: op1_04_inv23 = 1;
    48: op1_04_inv23 = 1;
    50: op1_04_inv23 = 1;
    54: op1_04_inv23 = 1;
    57: op1_04_inv23 = 1;
    58: op1_04_inv23 = 1;
    59: op1_04_inv23 = 1;
    65: op1_04_inv23 = 1;
    69: op1_04_inv23 = 1;
    71: op1_04_inv23 = 1;
    78: op1_04_inv23 = 1;
    80: op1_04_inv23 = 1;
    83: op1_04_inv23 = 1;
    85: op1_04_inv23 = 1;
    86: op1_04_inv23 = 1;
    87: op1_04_inv23 = 1;
    89: op1_04_inv23 = 1;
    90: op1_04_inv23 = 1;
    91: op1_04_inv23 = 1;
    92: op1_04_inv23 = 1;
    default: op1_04_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の24番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in24 = imem06_in[95:92];
    7: op1_04_in24 = reg_0518;
    8: op1_04_in24 = imem05_in[107:104];
    9: op1_04_in24 = imem06_in[99:96];
    12: op1_04_in24 = imem06_in[99:96];
    10: op1_04_in24 = reg_0137;
    11: op1_04_in24 = reg_0161;
    13: op1_04_in24 = reg_0127;
    14: op1_04_in24 = imem05_in[15:12];
    46: op1_04_in24 = imem05_in[15:12];
    80: op1_04_in24 = imem05_in[15:12];
    15: op1_04_in24 = reg_0787;
    16: op1_04_in24 = imem01_in[103:100];
    17: op1_04_in24 = reg_0583;
    19: op1_04_in24 = reg_0548;
    20: op1_04_in24 = imem07_in[63:60];
    21: op1_04_in24 = reg_0321;
    22: op1_04_in24 = reg_0722;
    23: op1_04_in24 = reg_0183;
    24: op1_04_in24 = reg_0128;
    25: op1_04_in24 = imem01_in[15:12];
    26: op1_04_in24 = reg_0592;
    27: op1_04_in24 = reg_1015;
    28: op1_04_in24 = reg_0336;
    29: op1_04_in24 = reg_0724;
    31: op1_04_in24 = reg_0319;
    32: op1_04_in24 = reg_0135;
    33: op1_04_in24 = reg_0427;
    34: op1_04_in24 = reg_1017;
    35: op1_04_in24 = imem07_in[19:16];
    36: op1_04_in24 = reg_0489;
    37: op1_04_in24 = imem07_in[27:24];
    38: op1_04_in24 = reg_0710;
    40: op1_04_in24 = reg_0248;
    42: op1_04_in24 = reg_1057;
    43: op1_04_in24 = reg_0383;
    45: op1_04_in24 = reg_0091;
    48: op1_04_in24 = reg_0738;
    49: op1_04_in24 = reg_0942;
    50: op1_04_in24 = reg_0975;
    51: op1_04_in24 = reg_0339;
    53: op1_04_in24 = reg_0906;
    54: op1_04_in24 = reg_0343;
    55: op1_04_in24 = reg_0374;
    56: op1_04_in24 = reg_0511;
    57: op1_04_in24 = reg_0813;
    58: op1_04_in24 = imem06_in[67:64];
    59: op1_04_in24 = imem05_in[39:36];
    61: op1_04_in24 = reg_0731;
    63: op1_04_in24 = reg_0079;
    64: op1_04_in24 = reg_0847;
    65: op1_04_in24 = reg_0892;
    66: op1_04_in24 = reg_0968;
    67: op1_04_in24 = reg_1005;
    68: op1_04_in24 = imem06_in[107:104];
    69: op1_04_in24 = reg_0226;
    70: op1_04_in24 = imem03_in[43:40];
    71: op1_04_in24 = reg_0218;
    72: op1_04_in24 = reg_0577;
    73: op1_04_in24 = reg_1004;
    74: op1_04_in24 = reg_0736;
    75: op1_04_in24 = reg_0591;
    78: op1_04_in24 = reg_0522;
    79: op1_04_in24 = imem04_in[87:84];
    81: op1_04_in24 = imem06_in[127:124];
    82: op1_04_in24 = reg_0819;
    83: op1_04_in24 = reg_0501;
    85: op1_04_in24 = reg_0815;
    86: op1_04_in24 = reg_0270;
    87: op1_04_in24 = reg_0095;
    88: op1_04_in24 = imem03_in[75:72];
    89: op1_04_in24 = reg_0422;
    90: op1_04_in24 = imem05_in[91:88];
    91: op1_04_in24 = reg_0178;
    92: op1_04_in24 = reg_0063;
    97: op1_04_in24 = reg_0919;
    default: op1_04_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_04_inv24 = 1;
    10: op1_04_inv24 = 1;
    11: op1_04_inv24 = 1;
    12: op1_04_inv24 = 1;
    14: op1_04_inv24 = 1;
    15: op1_04_inv24 = 1;
    22: op1_04_inv24 = 1;
    24: op1_04_inv24 = 1;
    25: op1_04_inv24 = 1;
    26: op1_04_inv24 = 1;
    27: op1_04_inv24 = 1;
    28: op1_04_inv24 = 1;
    29: op1_04_inv24 = 1;
    37: op1_04_inv24 = 1;
    38: op1_04_inv24 = 1;
    42: op1_04_inv24 = 1;
    43: op1_04_inv24 = 1;
    45: op1_04_inv24 = 1;
    49: op1_04_inv24 = 1;
    50: op1_04_inv24 = 1;
    54: op1_04_inv24 = 1;
    55: op1_04_inv24 = 1;
    64: op1_04_inv24 = 1;
    65: op1_04_inv24 = 1;
    67: op1_04_inv24 = 1;
    69: op1_04_inv24 = 1;
    70: op1_04_inv24 = 1;
    71: op1_04_inv24 = 1;
    72: op1_04_inv24 = 1;
    79: op1_04_inv24 = 1;
    80: op1_04_inv24 = 1;
    85: op1_04_inv24 = 1;
    86: op1_04_inv24 = 1;
    87: op1_04_inv24 = 1;
    88: op1_04_inv24 = 1;
    90: op1_04_inv24 = 1;
    92: op1_04_inv24 = 1;
    97: op1_04_inv24 = 1;
    default: op1_04_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の25番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in25 = reg_0628;
    7: op1_04_in25 = reg_0515;
    8: op1_04_in25 = imem05_in[115:112];
    9: op1_04_in25 = imem06_in[115:112];
    10: op1_04_in25 = imem06_in[15:12];
    11: op1_04_in25 = reg_0163;
    12: op1_04_in25 = imem06_in[119:116];
    13: op1_04_in25 = imem02_in[3:0];
    14: op1_04_in25 = imem05_in[39:36];
    15: op1_04_in25 = reg_0486;
    16: op1_04_in25 = imem01_in[107:104];
    17: op1_04_in25 = reg_0592;
    19: op1_04_in25 = reg_0555;
    20: op1_04_in25 = imem07_in[107:104];
    21: op1_04_in25 = reg_0397;
    22: op1_04_in25 = reg_0716;
    23: op1_04_in25 = reg_0177;
    24: op1_04_in25 = reg_0152;
    25: op1_04_in25 = imem01_in[39:36];
    26: op1_04_in25 = reg_0585;
    72: op1_04_in25 = reg_0585;
    27: op1_04_in25 = reg_1045;
    28: op1_04_in25 = reg_0482;
    29: op1_04_in25 = reg_0715;
    31: op1_04_in25 = imem03_in[7:4];
    45: op1_04_in25 = imem03_in[7:4];
    32: op1_04_in25 = reg_0143;
    33: op1_04_in25 = reg_0448;
    34: op1_04_in25 = reg_0122;
    35: op1_04_in25 = imem07_in[59:56];
    36: op1_04_in25 = reg_0145;
    37: op1_04_in25 = imem07_in[31:28];
    38: op1_04_in25 = reg_0729;
    40: op1_04_in25 = reg_0544;
    42: op1_04_in25 = reg_1020;
    43: op1_04_in25 = reg_0243;
    46: op1_04_in25 = imem05_in[19:16];
    48: op1_04_in25 = imem01_in[47:44];
    49: op1_04_in25 = reg_0961;
    50: op1_04_in25 = reg_0976;
    51: op1_04_in25 = reg_0007;
    53: op1_04_in25 = imem01_in[15:12];
    54: op1_04_in25 = imem03_in[3:0];
    63: op1_04_in25 = imem03_in[3:0];
    55: op1_04_in25 = reg_0974;
    56: op1_04_in25 = reg_1005;
    57: op1_04_in25 = reg_0094;
    58: op1_04_in25 = imem06_in[75:72];
    59: op1_04_in25 = imem05_in[43:40];
    61: op1_04_in25 = reg_0705;
    64: op1_04_in25 = reg_0793;
    65: op1_04_in25 = reg_0235;
    66: op1_04_in25 = reg_0945;
    67: op1_04_in25 = reg_0888;
    68: op1_04_in25 = imem06_in[111:108];
    69: op1_04_in25 = reg_0045;
    70: op1_04_in25 = imem03_in[59:56];
    71: op1_04_in25 = reg_0390;
    73: op1_04_in25 = reg_0483;
    74: op1_04_in25 = reg_0130;
    75: op1_04_in25 = reg_0008;
    78: op1_04_in25 = reg_0798;
    79: op1_04_in25 = imem04_in[119:116];
    80: op1_04_in25 = reg_0826;
    81: op1_04_in25 = reg_0080;
    82: op1_04_in25 = reg_0780;
    83: op1_04_in25 = reg_0869;
    85: op1_04_in25 = reg_0072;
    86: op1_04_in25 = imem07_in[23:20];
    87: op1_04_in25 = reg_0441;
    88: op1_04_in25 = reg_0756;
    89: op1_04_in25 = reg_0589;
    90: op1_04_in25 = imem05_in[95:92];
    91: op1_04_in25 = reg_0063;
    92: op1_04_in25 = reg_0947;
    97: op1_04_in25 = reg_0124;
    default: op1_04_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv25 = 1;
    7: op1_04_inv25 = 1;
    8: op1_04_inv25 = 1;
    10: op1_04_inv25 = 1;
    12: op1_04_inv25 = 1;
    14: op1_04_inv25 = 1;
    19: op1_04_inv25 = 1;
    20: op1_04_inv25 = 1;
    21: op1_04_inv25 = 1;
    22: op1_04_inv25 = 1;
    23: op1_04_inv25 = 1;
    24: op1_04_inv25 = 1;
    26: op1_04_inv25 = 1;
    27: op1_04_inv25 = 1;
    28: op1_04_inv25 = 1;
    29: op1_04_inv25 = 1;
    34: op1_04_inv25 = 1;
    35: op1_04_inv25 = 1;
    36: op1_04_inv25 = 1;
    37: op1_04_inv25 = 1;
    38: op1_04_inv25 = 1;
    40: op1_04_inv25 = 1;
    42: op1_04_inv25 = 1;
    43: op1_04_inv25 = 1;
    48: op1_04_inv25 = 1;
    51: op1_04_inv25 = 1;
    53: op1_04_inv25 = 1;
    54: op1_04_inv25 = 1;
    55: op1_04_inv25 = 1;
    56: op1_04_inv25 = 1;
    57: op1_04_inv25 = 1;
    59: op1_04_inv25 = 1;
    61: op1_04_inv25 = 1;
    63: op1_04_inv25 = 1;
    65: op1_04_inv25 = 1;
    69: op1_04_inv25 = 1;
    71: op1_04_inv25 = 1;
    72: op1_04_inv25 = 1;
    73: op1_04_inv25 = 1;
    74: op1_04_inv25 = 1;
    75: op1_04_inv25 = 1;
    82: op1_04_inv25 = 1;
    87: op1_04_inv25 = 1;
    89: op1_04_inv25 = 1;
    92: op1_04_inv25 = 1;
    97: op1_04_inv25 = 1;
    default: op1_04_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の26番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in26 = reg_0613;
    7: op1_04_in26 = reg_0233;
    8: op1_04_in26 = reg_0955;
    9: op1_04_in26 = imem07_in[39:36];
    86: op1_04_in26 = imem07_in[39:36];
    10: op1_04_in26 = imem06_in[39:36];
    11: op1_04_in26 = reg_0183;
    12: op1_04_in26 = reg_0628;
    13: op1_04_in26 = reg_0645;
    14: op1_04_in26 = imem05_in[43:40];
    15: op1_04_in26 = reg_0801;
    16: op1_04_in26 = reg_0766;
    17: op1_04_in26 = reg_0578;
    19: op1_04_in26 = reg_0549;
    20: op1_04_in26 = reg_0721;
    21: op1_04_in26 = reg_0389;
    22: op1_04_in26 = reg_0712;
    23: op1_04_in26 = reg_0168;
    24: op1_04_in26 = reg_0146;
    25: op1_04_in26 = imem01_in[51:48];
    26: op1_04_in26 = reg_0593;
    27: op1_04_in26 = reg_1018;
    28: op1_04_in26 = reg_0089;
    29: op1_04_in26 = reg_0701;
    31: op1_04_in26 = imem03_in[15:12];
    32: op1_04_in26 = reg_0139;
    33: op1_04_in26 = reg_0435;
    34: op1_04_in26 = reg_0116;
    35: op1_04_in26 = imem07_in[103:100];
    36: op1_04_in26 = reg_0133;
    37: op1_04_in26 = imem07_in[47:44];
    38: op1_04_in26 = reg_0705;
    40: op1_04_in26 = reg_0811;
    42: op1_04_in26 = reg_0537;
    43: op1_04_in26 = reg_1029;
    45: op1_04_in26 = imem03_in[43:40];
    46: op1_04_in26 = imem05_in[27:24];
    48: op1_04_in26 = imem01_in[59:56];
    49: op1_04_in26 = reg_0972;
    50: op1_04_in26 = imem04_in[27:24];
    51: op1_04_in26 = reg_0085;
    53: op1_04_in26 = imem01_in[27:24];
    69: op1_04_in26 = imem01_in[27:24];
    54: op1_04_in26 = imem03_in[19:16];
    55: op1_04_in26 = reg_0977;
    56: op1_04_in26 = reg_0888;
    57: op1_04_in26 = reg_0404;
    58: op1_04_in26 = reg_0780;
    59: op1_04_in26 = imem05_in[47:44];
    61: op1_04_in26 = reg_0707;
    63: op1_04_in26 = imem03_in[7:4];
    64: op1_04_in26 = reg_0784;
    65: op1_04_in26 = reg_0269;
    66: op1_04_in26 = reg_0437;
    67: op1_04_in26 = reg_0313;
    68: op1_04_in26 = imem06_in[119:116];
    70: op1_04_in26 = imem03_in[63:60];
    71: op1_04_in26 = reg_0005;
    72: op1_04_in26 = reg_0434;
    73: op1_04_in26 = reg_0778;
    74: op1_04_in26 = reg_0131;
    75: op1_04_in26 = reg_0804;
    78: op1_04_in26 = reg_0500;
    79: op1_04_in26 = imem04_in[123:120];
    80: op1_04_in26 = reg_0217;
    81: op1_04_in26 = reg_0889;
    82: op1_04_in26 = reg_0806;
    83: op1_04_in26 = reg_0830;
    85: op1_04_in26 = reg_0284;
    87: op1_04_in26 = reg_0664;
    88: op1_04_in26 = reg_0230;
    89: op1_04_in26 = reg_0502;
    90: op1_04_in26 = imem05_in[103:100];
    91: op1_04_in26 = reg_0947;
    92: op1_04_in26 = reg_0023;
    97: op1_04_in26 = reg_0177;
    default: op1_04_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv26 = 1;
    9: op1_04_inv26 = 1;
    10: op1_04_inv26 = 1;
    11: op1_04_inv26 = 1;
    12: op1_04_inv26 = 1;
    13: op1_04_inv26 = 1;
    17: op1_04_inv26 = 1;
    19: op1_04_inv26 = 1;
    21: op1_04_inv26 = 1;
    24: op1_04_inv26 = 1;
    25: op1_04_inv26 = 1;
    26: op1_04_inv26 = 1;
    27: op1_04_inv26 = 1;
    29: op1_04_inv26 = 1;
    32: op1_04_inv26 = 1;
    33: op1_04_inv26 = 1;
    34: op1_04_inv26 = 1;
    36: op1_04_inv26 = 1;
    38: op1_04_inv26 = 1;
    46: op1_04_inv26 = 1;
    49: op1_04_inv26 = 1;
    51: op1_04_inv26 = 1;
    53: op1_04_inv26 = 1;
    55: op1_04_inv26 = 1;
    56: op1_04_inv26 = 1;
    59: op1_04_inv26 = 1;
    64: op1_04_inv26 = 1;
    66: op1_04_inv26 = 1;
    68: op1_04_inv26 = 1;
    71: op1_04_inv26 = 1;
    72: op1_04_inv26 = 1;
    74: op1_04_inv26 = 1;
    75: op1_04_inv26 = 1;
    80: op1_04_inv26 = 1;
    83: op1_04_inv26 = 1;
    85: op1_04_inv26 = 1;
    86: op1_04_inv26 = 1;
    87: op1_04_inv26 = 1;
    90: op1_04_inv26 = 1;
    92: op1_04_inv26 = 1;
    default: op1_04_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の27番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in27 = reg_0612;
    7: op1_04_in27 = reg_0246;
    8: op1_04_in27 = reg_0956;
    9: op1_04_in27 = imem07_in[47:44];
    86: op1_04_in27 = imem07_in[47:44];
    10: op1_04_in27 = imem06_in[67:64];
    12: op1_04_in27 = reg_0351;
    13: op1_04_in27 = reg_0666;
    14: op1_04_in27 = imem05_in[67:64];
    15: op1_04_in27 = reg_0781;
    16: op1_04_in27 = reg_0220;
    17: op1_04_in27 = reg_0360;
    19: op1_04_in27 = reg_0546;
    20: op1_04_in27 = reg_0729;
    21: op1_04_in27 = reg_0985;
    22: op1_04_in27 = reg_0709;
    23: op1_04_in27 = reg_0173;
    24: op1_04_in27 = reg_0138;
    25: op1_04_in27 = imem01_in[79:76];
    26: op1_04_in27 = reg_0597;
    27: op1_04_in27 = reg_0108;
    28: op1_04_in27 = reg_0776;
    29: op1_04_in27 = reg_0429;
    31: op1_04_in27 = imem03_in[35:32];
    32: op1_04_in27 = reg_0153;
    33: op1_04_in27 = reg_0180;
    34: op1_04_in27 = imem02_in[3:0];
    35: op1_04_in27 = reg_0728;
    36: op1_04_in27 = reg_0142;
    80: op1_04_in27 = reg_0142;
    37: op1_04_in27 = reg_0717;
    38: op1_04_in27 = reg_0707;
    40: op1_04_in27 = reg_0219;
    42: op1_04_in27 = imem04_in[39:36];
    43: op1_04_in27 = reg_0605;
    45: op1_04_in27 = imem03_in[55:52];
    46: op1_04_in27 = imem05_in[87:84];
    48: op1_04_in27 = imem01_in[75:72];
    49: op1_04_in27 = reg_0275;
    50: op1_04_in27 = imem04_in[35:32];
    51: op1_04_in27 = reg_0086;
    53: op1_04_in27 = imem01_in[35:32];
    54: op1_04_in27 = imem03_in[39:36];
    55: op1_04_in27 = reg_0988;
    56: op1_04_in27 = reg_0932;
    57: op1_04_in27 = reg_0438;
    58: op1_04_in27 = reg_0241;
    59: op1_04_in27 = imem05_in[107:104];
    61: op1_04_in27 = reg_0706;
    63: op1_04_in27 = imem03_in[15:12];
    64: op1_04_in27 = reg_0509;
    65: op1_04_in27 = reg_0953;
    66: op1_04_in27 = reg_0896;
    67: op1_04_in27 = reg_0802;
    68: op1_04_in27 = imem06_in[123:120];
    69: op1_04_in27 = imem01_in[71:68];
    70: op1_04_in27 = imem03_in[83:80];
    71: op1_04_in27 = reg_0625;
    72: op1_04_in27 = reg_0240;
    73: op1_04_in27 = reg_1016;
    74: op1_04_in27 = reg_0492;
    75: op1_04_in27 = reg_0222;
    78: op1_04_in27 = reg_0227;
    79: op1_04_in27 = imem04_in[127:124];
    81: op1_04_in27 = reg_0028;
    82: op1_04_in27 = reg_0816;
    83: op1_04_in27 = reg_0232;
    85: op1_04_in27 = reg_0658;
    87: op1_04_in27 = reg_0329;
    88: op1_04_in27 = reg_0377;
    89: op1_04_in27 = reg_0640;
    90: op1_04_in27 = imem05_in[111:108];
    91: op1_04_in27 = reg_0023;
    92: op1_04_in27 = reg_0964;
    97: op1_04_in27 = reg_0018;
    default: op1_04_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv27 = 1;
    8: op1_04_inv27 = 1;
    9: op1_04_inv27 = 1;
    13: op1_04_inv27 = 1;
    15: op1_04_inv27 = 1;
    16: op1_04_inv27 = 1;
    21: op1_04_inv27 = 1;
    23: op1_04_inv27 = 1;
    27: op1_04_inv27 = 1;
    31: op1_04_inv27 = 1;
    35: op1_04_inv27 = 1;
    37: op1_04_inv27 = 1;
    45: op1_04_inv27 = 1;
    50: op1_04_inv27 = 1;
    51: op1_04_inv27 = 1;
    53: op1_04_inv27 = 1;
    54: op1_04_inv27 = 1;
    56: op1_04_inv27 = 1;
    57: op1_04_inv27 = 1;
    58: op1_04_inv27 = 1;
    59: op1_04_inv27 = 1;
    61: op1_04_inv27 = 1;
    65: op1_04_inv27 = 1;
    66: op1_04_inv27 = 1;
    67: op1_04_inv27 = 1;
    70: op1_04_inv27 = 1;
    71: op1_04_inv27 = 1;
    74: op1_04_inv27 = 1;
    75: op1_04_inv27 = 1;
    78: op1_04_inv27 = 1;
    86: op1_04_inv27 = 1;
    87: op1_04_inv27 = 1;
    88: op1_04_inv27 = 1;
    89: op1_04_inv27 = 1;
    90: op1_04_inv27 = 1;
    91: op1_04_inv27 = 1;
    97: op1_04_inv27 = 1;
    default: op1_04_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の28番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in28 = reg_0348;
    7: op1_04_in28 = reg_0245;
    8: op1_04_in28 = reg_0964;
    9: op1_04_in28 = imem07_in[83:80];
    10: op1_04_in28 = imem06_in[71:68];
    12: op1_04_in28 = reg_0018;
    13: op1_04_in28 = reg_0639;
    14: op1_04_in28 = imem05_in[79:76];
    15: op1_04_in28 = reg_1010;
    16: op1_04_in28 = reg_0247;
    17: op1_04_in28 = reg_0370;
    19: op1_04_in28 = reg_0540;
    20: op1_04_in28 = reg_0709;
    21: op1_04_in28 = reg_0998;
    22: op1_04_in28 = reg_0718;
    23: op1_04_in28 = reg_0171;
    24: op1_04_in28 = reg_0144;
    25: op1_04_in28 = imem01_in[103:100];
    26: op1_04_in28 = reg_0570;
    27: op1_04_in28 = reg_0114;
    28: op1_04_in28 = reg_0086;
    29: op1_04_in28 = reg_0174;
    31: op1_04_in28 = imem03_in[43:40];
    54: op1_04_in28 = imem03_in[43:40];
    32: op1_04_in28 = reg_0799;
    56: op1_04_in28 = reg_0799;
    33: op1_04_in28 = reg_0165;
    34: op1_04_in28 = imem02_in[11:8];
    35: op1_04_in28 = reg_0720;
    36: op1_04_in28 = reg_0138;
    74: op1_04_in28 = reg_0138;
    37: op1_04_in28 = reg_0729;
    38: op1_04_in28 = reg_0428;
    40: op1_04_in28 = imem01_in[47:44];
    42: op1_04_in28 = imem04_in[55:52];
    43: op1_04_in28 = reg_0626;
    45: op1_04_in28 = imem03_in[111:108];
    46: op1_04_in28 = imem05_in[99:96];
    48: op1_04_in28 = imem01_in[83:80];
    49: op1_04_in28 = reg_0896;
    50: op1_04_in28 = imem04_in[39:36];
    51: op1_04_in28 = imem03_in[15:12];
    53: op1_04_in28 = imem01_in[67:64];
    55: op1_04_in28 = imem04_in[7:4];
    57: op1_04_in28 = reg_0148;
    58: op1_04_in28 = reg_0605;
    59: op1_04_in28 = imem05_in[123:120];
    90: op1_04_in28 = imem05_in[123:120];
    61: op1_04_in28 = reg_0727;
    63: op1_04_in28 = imem03_in[27:24];
    64: op1_04_in28 = reg_0992;
    70: op1_04_in28 = reg_0992;
    65: op1_04_in28 = imem05_in[7:4];
    66: op1_04_in28 = reg_0657;
    67: op1_04_in28 = reg_0066;
    68: op1_04_in28 = reg_0926;
    69: op1_04_in28 = imem01_in[107:104];
    71: op1_04_in28 = reg_0244;
    72: op1_04_in28 = reg_0662;
    73: op1_04_in28 = reg_0058;
    75: op1_04_in28 = reg_0293;
    78: op1_04_in28 = reg_0737;
    79: op1_04_in28 = reg_1004;
    80: op1_04_in28 = reg_0275;
    81: op1_04_in28 = reg_0895;
    82: op1_04_in28 = reg_0951;
    83: op1_04_in28 = reg_1055;
    85: op1_04_in28 = reg_0444;
    86: op1_04_in28 = imem07_in[55:52];
    87: op1_04_in28 = reg_0394;
    88: op1_04_in28 = reg_0376;
    89: op1_04_in28 = reg_0157;
    91: op1_04_in28 = reg_0130;
    92: op1_04_in28 = reg_0330;
    97: op1_04_in28 = reg_0611;
    default: op1_04_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_04_inv28 = 1;
    10: op1_04_inv28 = 1;
    12: op1_04_inv28 = 1;
    16: op1_04_inv28 = 1;
    21: op1_04_inv28 = 1;
    23: op1_04_inv28 = 1;
    25: op1_04_inv28 = 1;
    26: op1_04_inv28 = 1;
    29: op1_04_inv28 = 1;
    31: op1_04_inv28 = 1;
    36: op1_04_inv28 = 1;
    38: op1_04_inv28 = 1;
    46: op1_04_inv28 = 1;
    48: op1_04_inv28 = 1;
    49: op1_04_inv28 = 1;
    50: op1_04_inv28 = 1;
    53: op1_04_inv28 = 1;
    54: op1_04_inv28 = 1;
    58: op1_04_inv28 = 1;
    59: op1_04_inv28 = 1;
    61: op1_04_inv28 = 1;
    63: op1_04_inv28 = 1;
    64: op1_04_inv28 = 1;
    65: op1_04_inv28 = 1;
    66: op1_04_inv28 = 1;
    68: op1_04_inv28 = 1;
    70: op1_04_inv28 = 1;
    72: op1_04_inv28 = 1;
    78: op1_04_inv28 = 1;
    83: op1_04_inv28 = 1;
    87: op1_04_inv28 = 1;
    88: op1_04_inv28 = 1;
    89: op1_04_inv28 = 1;
    90: op1_04_inv28 = 1;
    91: op1_04_inv28 = 1;
    97: op1_04_inv28 = 1;
    default: op1_04_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の29番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in29 = reg_0356;
    7: op1_04_in29 = reg_0221;
    8: op1_04_in29 = reg_0951;
    9: op1_04_in29 = reg_0730;
    10: op1_04_in29 = imem06_in[87:84];
    12: op1_04_in29 = reg_0754;
    68: op1_04_in29 = reg_0754;
    13: op1_04_in29 = reg_0648;
    14: op1_04_in29 = imem05_in[95:92];
    15: op1_04_in29 = reg_1011;
    16: op1_04_in29 = reg_1018;
    17: op1_04_in29 = reg_0319;
    19: op1_04_in29 = imem04_in[15:12];
    20: op1_04_in29 = reg_0425;
    21: op1_04_in29 = reg_1002;
    22: op1_04_in29 = reg_0707;
    24: op1_04_in29 = imem06_in[7:4];
    25: op1_04_in29 = imem01_in[123:120];
    26: op1_04_in29 = reg_0373;
    27: op1_04_in29 = reg_0113;
    28: op1_04_in29 = reg_0506;
    29: op1_04_in29 = reg_0165;
    31: op1_04_in29 = imem03_in[55:52];
    32: op1_04_in29 = reg_0372;
    33: op1_04_in29 = reg_0183;
    34: op1_04_in29 = imem02_in[67:64];
    35: op1_04_in29 = reg_0721;
    36: op1_04_in29 = reg_0153;
    37: op1_04_in29 = reg_0713;
    38: op1_04_in29 = reg_0438;
    40: op1_04_in29 = imem01_in[55:52];
    42: op1_04_in29 = reg_0525;
    43: op1_04_in29 = reg_0531;
    45: op1_04_in29 = reg_0573;
    46: op1_04_in29 = reg_0962;
    48: op1_04_in29 = imem01_in[115:112];
    49: op1_04_in29 = reg_0832;
    50: op1_04_in29 = imem04_in[55:52];
    51: op1_04_in29 = imem03_in[79:76];
    54: op1_04_in29 = imem03_in[79:76];
    53: op1_04_in29 = imem01_in[75:72];
    55: op1_04_in29 = imem04_in[95:92];
    56: op1_04_in29 = reg_0076;
    57: op1_04_in29 = reg_0136;
    90: op1_04_in29 = reg_0136;
    58: op1_04_in29 = reg_0017;
    59: op1_04_in29 = reg_0835;
    61: op1_04_in29 = reg_0002;
    63: op1_04_in29 = imem03_in[103:100];
    64: op1_04_in29 = reg_0984;
    65: op1_04_in29 = imem05_in[99:96];
    66: op1_04_in29 = imem05_in[23:20];
    67: op1_04_in29 = reg_0068;
    69: op1_04_in29 = reg_0520;
    70: op1_04_in29 = reg_1001;
    71: op1_04_in29 = reg_0021;
    72: op1_04_in29 = reg_0238;
    73: op1_04_in29 = reg_0066;
    74: op1_04_in29 = reg_0255;
    75: op1_04_in29 = reg_0403;
    78: op1_04_in29 = reg_0521;
    79: op1_04_in29 = reg_0536;
    80: op1_04_in29 = reg_0952;
    81: op1_04_in29 = reg_0392;
    82: op1_04_in29 = reg_0851;
    83: op1_04_in29 = reg_0283;
    85: op1_04_in29 = reg_0065;
    86: op1_04_in29 = imem07_in[111:108];
    87: op1_04_in29 = reg_0368;
    88: op1_04_in29 = reg_0987;
    91: op1_04_in29 = reg_0437;
    92: op1_04_in29 = reg_0130;
    97: op1_04_in29 = reg_0782;
    default: op1_04_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv29 = 1;
    9: op1_04_inv29 = 1;
    10: op1_04_inv29 = 1;
    12: op1_04_inv29 = 1;
    13: op1_04_inv29 = 1;
    14: op1_04_inv29 = 1;
    17: op1_04_inv29 = 1;
    19: op1_04_inv29 = 1;
    20: op1_04_inv29 = 1;
    22: op1_04_inv29 = 1;
    26: op1_04_inv29 = 1;
    27: op1_04_inv29 = 1;
    29: op1_04_inv29 = 1;
    31: op1_04_inv29 = 1;
    34: op1_04_inv29 = 1;
    35: op1_04_inv29 = 1;
    37: op1_04_inv29 = 1;
    40: op1_04_inv29 = 1;
    43: op1_04_inv29 = 1;
    49: op1_04_inv29 = 1;
    50: op1_04_inv29 = 1;
    54: op1_04_inv29 = 1;
    55: op1_04_inv29 = 1;
    56: op1_04_inv29 = 1;
    59: op1_04_inv29 = 1;
    61: op1_04_inv29 = 1;
    63: op1_04_inv29 = 1;
    64: op1_04_inv29 = 1;
    65: op1_04_inv29 = 1;
    66: op1_04_inv29 = 1;
    67: op1_04_inv29 = 1;
    68: op1_04_inv29 = 1;
    70: op1_04_inv29 = 1;
    72: op1_04_inv29 = 1;
    73: op1_04_inv29 = 1;
    78: op1_04_inv29 = 1;
    79: op1_04_inv29 = 1;
    85: op1_04_inv29 = 1;
    87: op1_04_inv29 = 1;
    90: op1_04_inv29 = 1;
    91: op1_04_inv29 = 1;
    97: op1_04_inv29 = 1;
    default: op1_04_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の30番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_04_in30 = reg_0382;
    7: op1_04_in30 = reg_0123;
    8: op1_04_in30 = reg_0942;
    9: op1_04_in30 = reg_0731;
    10: op1_04_in30 = imem06_in[99:96];
    12: op1_04_in30 = imem07_in[31:28];
    13: op1_04_in30 = reg_0643;
    14: op1_04_in30 = imem05_in[107:104];
    15: op1_04_in30 = reg_0754;
    16: op1_04_in30 = reg_0904;
    17: op1_04_in30 = reg_0385;
    19: op1_04_in30 = imem04_in[35:32];
    20: op1_04_in30 = reg_0436;
    21: op1_04_in30 = reg_0979;
    22: op1_04_in30 = reg_0426;
    24: op1_04_in30 = imem06_in[95:92];
    25: op1_04_in30 = reg_0905;
    26: op1_04_in30 = reg_0986;
    27: op1_04_in30 = reg_0110;
    28: op1_04_in30 = reg_0484;
    29: op1_04_in30 = reg_0162;
    31: op1_04_in30 = imem03_in[75:72];
    32: op1_04_in30 = reg_0556;
    33: op1_04_in30 = reg_0185;
    34: op1_04_in30 = imem02_in[83:80];
    35: op1_04_in30 = reg_0714;
    36: op1_04_in30 = reg_0614;
    37: op1_04_in30 = reg_0718;
    38: op1_04_in30 = reg_0448;
    40: op1_04_in30 = imem01_in[111:108];
    42: op1_04_in30 = reg_0279;
    43: op1_04_in30 = reg_0621;
    45: op1_04_in30 = reg_1007;
    46: op1_04_in30 = reg_0973;
    48: op1_04_in30 = imem01_in[119:116];
    49: op1_04_in30 = reg_0831;
    50: op1_04_in30 = imem04_in[119:116];
    51: op1_04_in30 = imem03_in[111:108];
    53: op1_04_in30 = imem01_in[87:84];
    54: op1_04_in30 = imem03_in[87:84];
    55: op1_04_in30 = imem04_in[103:100];
    56: op1_04_in30 = reg_0056;
    57: op1_04_in30 = reg_0133;
    58: op1_04_in30 = reg_0029;
    59: op1_04_in30 = reg_0955;
    61: op1_04_in30 = reg_0315;
    63: op1_04_in30 = reg_0572;
    64: op1_04_in30 = reg_1001;
    65: op1_04_in30 = imem05_in[123:120];
    66: op1_04_in30 = imem05_in[71:68];
    67: op1_04_in30 = reg_0732;
    68: op1_04_in30 = reg_0028;
    69: op1_04_in30 = reg_0925;
    70: op1_04_in30 = reg_0980;
    71: op1_04_in30 = reg_0817;
    72: op1_04_in30 = reg_0230;
    73: op1_04_in30 = reg_0014;
    74: op1_04_in30 = reg_0960;
    75: op1_04_in30 = reg_0782;
    78: op1_04_in30 = reg_0610;
    79: op1_04_in30 = reg_0301;
    80: op1_04_in30 = reg_0819;
    81: op1_04_in30 = reg_0611;
    82: op1_04_in30 = reg_0490;
    83: op1_04_in30 = imem02_in[7:4];
    85: op1_04_in30 = reg_0027;
    86: op1_04_in30 = reg_0567;
    87: op1_04_in30 = reg_0425;
    88: op1_04_in30 = reg_0989;
    90: op1_04_in30 = reg_0954;
    91: op1_04_in30 = reg_0587;
    92: op1_04_in30 = reg_0272;
    97: op1_04_in30 = reg_0804;
    default: op1_04_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv30 = 1;
    8: op1_04_inv30 = 1;
    10: op1_04_inv30 = 1;
    14: op1_04_inv30 = 1;
    16: op1_04_inv30 = 1;
    17: op1_04_inv30 = 1;
    19: op1_04_inv30 = 1;
    20: op1_04_inv30 = 1;
    24: op1_04_inv30 = 1;
    26: op1_04_inv30 = 1;
    28: op1_04_inv30 = 1;
    29: op1_04_inv30 = 1;
    31: op1_04_inv30 = 1;
    32: op1_04_inv30 = 1;
    35: op1_04_inv30 = 1;
    37: op1_04_inv30 = 1;
    38: op1_04_inv30 = 1;
    40: op1_04_inv30 = 1;
    42: op1_04_inv30 = 1;
    43: op1_04_inv30 = 1;
    48: op1_04_inv30 = 1;
    50: op1_04_inv30 = 1;
    51: op1_04_inv30 = 1;
    53: op1_04_inv30 = 1;
    54: op1_04_inv30 = 1;
    55: op1_04_inv30 = 1;
    57: op1_04_inv30 = 1;
    58: op1_04_inv30 = 1;
    63: op1_04_inv30 = 1;
    65: op1_04_inv30 = 1;
    68: op1_04_inv30 = 1;
    69: op1_04_inv30 = 1;
    70: op1_04_inv30 = 1;
    72: op1_04_inv30 = 1;
    73: op1_04_inv30 = 1;
    75: op1_04_inv30 = 1;
    78: op1_04_inv30 = 1;
    79: op1_04_inv30 = 1;
    82: op1_04_inv30 = 1;
    83: op1_04_inv30 = 1;
    86: op1_04_inv30 = 1;
    87: op1_04_inv30 = 1;
    88: op1_04_inv30 = 1;
    97: op1_04_inv30 = 1;
    default: op1_04_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_04_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_04_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in00 = imem00_in[31:28];
    11: op1_05_in00 = imem00_in[31:28];
    95: op1_05_in00 = imem00_in[31:28];
    6: op1_05_in00 = reg_0315;
    7: op1_05_in00 = reg_0122;
    8: op1_05_in00 = reg_0968;
    9: op1_05_in00 = imem00_in[55:52];
    77: op1_05_in00 = imem00_in[55:52];
    10: op1_05_in00 = reg_0630;
    12: op1_05_in00 = imem07_in[75:72];
    4: op1_05_in00 = imem07_in[47:44];
    13: op1_05_in00 = reg_0667;
    14: op1_05_in00 = imem05_in[127:124];
    15: op1_05_in00 = imem07_in[7:4];
    3: op1_05_in00 = imem07_in[7:4];
    97: op1_05_in00 = imem07_in[7:4];
    16: op1_05_in00 = reg_0124;
    17: op1_05_in00 = reg_0377;
    18: op1_05_in00 = imem00_in[7:4];
    23: op1_05_in00 = imem00_in[7:4];
    30: op1_05_in00 = imem00_in[7:4];
    62: op1_05_in00 = imem00_in[7:4];
    19: op1_05_in00 = imem04_in[51:48];
    20: op1_05_in00 = imem00_in[27:24];
    22: op1_05_in00 = imem00_in[27:24];
    21: op1_05_in00 = reg_0994;
    24: op1_05_in00 = imem06_in[127:124];
    2: op1_05_in00 = imem07_in[63:60];
    25: op1_05_in00 = reg_0869;
    26: op1_05_in00 = reg_0981;
    27: op1_05_in00 = imem02_in[7:4];
    28: op1_05_in00 = reg_0321;
    29: op1_05_in00 = imem00_in[67:64];
    31: op1_05_in00 = reg_0793;
    32: op1_05_in00 = reg_0614;
    33: op1_05_in00 = imem00_in[3:0];
    93: op1_05_in00 = imem00_in[3:0];
    34: op1_05_in00 = imem02_in[99:96];
    35: op1_05_in00 = reg_0711;
    37: op1_05_in00 = reg_0711;
    36: op1_05_in00 = reg_0613;
    38: op1_05_in00 = reg_0172;
    39: op1_05_in00 = imem00_in[95:92];
    40: op1_05_in00 = reg_0116;
    41: op1_05_in00 = imem00_in[35:32];
    47: op1_05_in00 = imem00_in[35:32];
    89: op1_05_in00 = imem00_in[35:32];
    42: op1_05_in00 = reg_0528;
    43: op1_05_in00 = reg_0027;
    44: op1_05_in00 = imem00_in[47:44];
    45: op1_05_in00 = reg_0933;
    46: op1_05_in00 = reg_0966;
    48: op1_05_in00 = reg_0604;
    49: op1_05_in00 = reg_0152;
    50: op1_05_in00 = imem04_in[127:124];
    51: op1_05_in00 = imem03_in[127:124];
    52: op1_05_in00 = imem00_in[15:12];
    76: op1_05_in00 = imem00_in[15:12];
    84: op1_05_in00 = imem00_in[15:12];
    53: op1_05_in00 = imem01_in[95:92];
    54: op1_05_in00 = imem03_in[99:96];
    55: op1_05_in00 = imem04_in[111:108];
    56: op1_05_in00 = reg_0014;
    57: op1_05_in00 = reg_0142;
    58: op1_05_in00 = reg_0545;
    59: op1_05_in00 = reg_0492;
    60: op1_05_in00 = imem00_in[39:36];
    61: op1_05_in00 = reg_0641;
    63: op1_05_in00 = reg_0327;
    64: op1_05_in00 = reg_0975;
    65: op1_05_in00 = reg_0757;
    66: op1_05_in00 = imem05_in[83:80];
    67: op1_05_in00 = reg_0284;
    68: op1_05_in00 = reg_0297;
    69: op1_05_in00 = reg_0769;
    70: op1_05_in00 = reg_0977;
    71: op1_05_in00 = reg_0735;
    72: op1_05_in00 = reg_0984;
    73: op1_05_in00 = reg_0302;
    74: op1_05_in00 = imem05_in[51:48];
    75: op1_05_in00 = reg_0369;
    78: op1_05_in00 = reg_0111;
    79: op1_05_in00 = reg_0511;
    80: op1_05_in00 = reg_0780;
    81: op1_05_in00 = reg_0781;
    82: op1_05_in00 = reg_0144;
    83: op1_05_in00 = imem02_in[35:32];
    85: op1_05_in00 = reg_0495;
    86: op1_05_in00 = reg_0100;
    87: op1_05_in00 = reg_0608;
    88: op1_05_in00 = reg_0988;
    90: op1_05_in00 = reg_0139;
    91: op1_05_in00 = reg_0736;
    92: op1_05_in00 = reg_0530;
    94: op1_05_in00 = imem00_in[43:40];
    96: op1_05_in00 = imem00_in[103:100];
    default: op1_05_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv00 = 1;
    6: op1_05_inv00 = 1;
    7: op1_05_inv00 = 1;
    8: op1_05_inv00 = 1;
    9: op1_05_inv00 = 1;
    12: op1_05_inv00 = 1;
    15: op1_05_inv00 = 1;
    20: op1_05_inv00 = 1;
    21: op1_05_inv00 = 1;
    25: op1_05_inv00 = 1;
    26: op1_05_inv00 = 1;
    28: op1_05_inv00 = 1;
    29: op1_05_inv00 = 1;
    30: op1_05_inv00 = 1;
    31: op1_05_inv00 = 1;
    32: op1_05_inv00 = 1;
    35: op1_05_inv00 = 1;
    41: op1_05_inv00 = 1;
    43: op1_05_inv00 = 1;
    44: op1_05_inv00 = 1;
    46: op1_05_inv00 = 1;
    48: op1_05_inv00 = 1;
    50: op1_05_inv00 = 1;
    51: op1_05_inv00 = 1;
    52: op1_05_inv00 = 1;
    53: op1_05_inv00 = 1;
    55: op1_05_inv00 = 1;
    57: op1_05_inv00 = 1;
    58: op1_05_inv00 = 1;
    59: op1_05_inv00 = 1;
    60: op1_05_inv00 = 1;
    62: op1_05_inv00 = 1;
    64: op1_05_inv00 = 1;
    66: op1_05_inv00 = 1;
    68: op1_05_inv00 = 1;
    70: op1_05_inv00 = 1;
    71: op1_05_inv00 = 1;
    74: op1_05_inv00 = 1;
    77: op1_05_inv00 = 1;
    78: op1_05_inv00 = 1;
    80: op1_05_inv00 = 1;
    81: op1_05_inv00 = 1;
    84: op1_05_inv00 = 1;
    85: op1_05_inv00 = 1;
    86: op1_05_inv00 = 1;
    90: op1_05_inv00 = 1;
    91: op1_05_inv00 = 1;
    92: op1_05_inv00 = 1;
    97: op1_05_inv00 = 1;
    default: op1_05_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in01 = imem00_in[35:32];
    23: op1_05_in01 = imem00_in[35:32];
    6: op1_05_in01 = reg_0390;
    7: op1_05_in01 = imem02_in[3:0];
    8: op1_05_in01 = reg_0965;
    9: op1_05_in01 = imem00_in[79:76];
    10: op1_05_in01 = reg_0613;
    11: op1_05_in01 = imem00_in[47:44];
    47: op1_05_in01 = imem00_in[47:44];
    12: op1_05_in01 = imem07_in[123:120];
    4: op1_05_in01 = imem07_in[59:56];
    58: op1_05_in01 = imem07_in[59:56];
    13: op1_05_in01 = reg_0339;
    14: op1_05_in01 = reg_0958;
    15: op1_05_in01 = imem07_in[23:20];
    16: op1_05_in01 = reg_0125;
    17: op1_05_in01 = reg_0361;
    18: op1_05_in01 = reg_0682;
    19: op1_05_in01 = imem04_in[59:56];
    3: op1_05_in01 = imem07_in[19:16];
    20: op1_05_in01 = imem00_in[99:96];
    39: op1_05_in01 = imem00_in[99:96];
    21: op1_05_in01 = imem04_in[35:32];
    22: op1_05_in01 = imem00_in[51:48];
    44: op1_05_in01 = imem00_in[51:48];
    89: op1_05_in01 = imem00_in[51:48];
    24: op1_05_in01 = reg_0607;
    2: op1_05_in01 = imem07_in[83:80];
    25: op1_05_in01 = reg_0885;
    26: op1_05_in01 = reg_0997;
    27: op1_05_in01 = imem02_in[11:8];
    28: op1_05_in01 = reg_0561;
    29: op1_05_in01 = imem00_in[75:72];
    30: op1_05_in01 = imem00_in[27:24];
    76: op1_05_in01 = imem00_in[27:24];
    31: op1_05_in01 = reg_0370;
    32: op1_05_in01 = reg_0628;
    33: op1_05_in01 = imem00_in[19:16];
    52: op1_05_in01 = imem00_in[19:16];
    84: op1_05_in01 = imem00_in[19:16];
    34: op1_05_in01 = imem02_in[123:120];
    35: op1_05_in01 = reg_0426;
    36: op1_05_in01 = reg_0611;
    37: op1_05_in01 = reg_0424;
    38: op1_05_in01 = reg_0162;
    40: op1_05_in01 = reg_0100;
    41: op1_05_in01 = imem00_in[39:36];
    42: op1_05_in01 = imem05_in[79:76];
    43: op1_05_in01 = reg_0735;
    45: op1_05_in01 = reg_0046;
    46: op1_05_in01 = reg_0959;
    48: op1_05_in01 = reg_0520;
    49: op1_05_in01 = reg_0138;
    50: op1_05_in01 = reg_0301;
    55: op1_05_in01 = reg_0301;
    51: op1_05_in01 = reg_0006;
    53: op1_05_in01 = imem02_in[35:32];
    54: op1_05_in01 = imem03_in[107:104];
    56: op1_05_in01 = reg_0584;
    57: op1_05_in01 = reg_0139;
    59: op1_05_in01 = reg_0689;
    60: op1_05_in01 = imem00_in[43:40];
    61: op1_05_in01 = reg_0532;
    62: op1_05_in01 = reg_0841;
    63: op1_05_in01 = reg_0322;
    64: op1_05_in01 = imem04_in[55:52];
    65: op1_05_in01 = reg_0435;
    66: op1_05_in01 = imem05_in[127:124];
    67: op1_05_in01 = reg_0893;
    68: op1_05_in01 = reg_0392;
    69: op1_05_in01 = reg_0273;
    70: op1_05_in01 = reg_0988;
    71: op1_05_in01 = reg_0028;
    72: op1_05_in01 = reg_0993;
    73: op1_05_in01 = reg_0401;
    74: op1_05_in01 = imem05_in[95:92];
    75: op1_05_in01 = reg_0567;
    77: op1_05_in01 = imem00_in[59:56];
    95: op1_05_in01 = imem00_in[59:56];
    78: op1_05_in01 = reg_0003;
    79: op1_05_in01 = reg_1020;
    80: op1_05_in01 = reg_0145;
    81: op1_05_in01 = reg_0556;
    82: op1_05_in01 = imem06_in[7:4];
    83: op1_05_in01 = imem02_in[63:60];
    85: op1_05_in01 = reg_0108;
    86: op1_05_in01 = reg_0560;
    87: op1_05_in01 = reg_0347;
    88: op1_05_in01 = imem04_in[71:68];
    90: op1_05_in01 = reg_0235;
    91: op1_05_in01 = reg_0530;
    92: op1_05_in01 = reg_0806;
    93: op1_05_in01 = imem00_in[11:8];
    94: op1_05_in01 = imem00_in[87:84];
    96: op1_05_in01 = reg_0223;
    97: op1_05_in01 = imem07_in[39:36];
    default: op1_05_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv01 = 1;
    10: op1_05_inv01 = 1;
    12: op1_05_inv01 = 1;
    13: op1_05_inv01 = 1;
    14: op1_05_inv01 = 1;
    15: op1_05_inv01 = 1;
    16: op1_05_inv01 = 1;
    17: op1_05_inv01 = 1;
    19: op1_05_inv01 = 1;
    22: op1_05_inv01 = 1;
    24: op1_05_inv01 = 1;
    2: op1_05_inv01 = 1;
    25: op1_05_inv01 = 1;
    26: op1_05_inv01 = 1;
    28: op1_05_inv01 = 1;
    29: op1_05_inv01 = 1;
    30: op1_05_inv01 = 1;
    31: op1_05_inv01 = 1;
    32: op1_05_inv01 = 1;
    36: op1_05_inv01 = 1;
    40: op1_05_inv01 = 1;
    42: op1_05_inv01 = 1;
    43: op1_05_inv01 = 1;
    46: op1_05_inv01 = 1;
    47: op1_05_inv01 = 1;
    48: op1_05_inv01 = 1;
    49: op1_05_inv01 = 1;
    54: op1_05_inv01 = 1;
    58: op1_05_inv01 = 1;
    59: op1_05_inv01 = 1;
    60: op1_05_inv01 = 1;
    62: op1_05_inv01 = 1;
    63: op1_05_inv01 = 1;
    64: op1_05_inv01 = 1;
    65: op1_05_inv01 = 1;
    66: op1_05_inv01 = 1;
    68: op1_05_inv01 = 1;
    71: op1_05_inv01 = 1;
    72: op1_05_inv01 = 1;
    73: op1_05_inv01 = 1;
    75: op1_05_inv01 = 1;
    77: op1_05_inv01 = 1;
    80: op1_05_inv01 = 1;
    84: op1_05_inv01 = 1;
    86: op1_05_inv01 = 1;
    87: op1_05_inv01 = 1;
    89: op1_05_inv01 = 1;
    90: op1_05_inv01 = 1;
    91: op1_05_inv01 = 1;
    94: op1_05_inv01 = 1;
    95: op1_05_inv01 = 1;
    97: op1_05_inv01 = 1;
    default: op1_05_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in02 = imem00_in[51:48];
    6: op1_05_in02 = reg_0034;
    7: op1_05_in02 = imem02_in[11:8];
    8: op1_05_in02 = reg_0267;
    9: op1_05_in02 = imem00_in[123:120];
    10: op1_05_in02 = reg_0620;
    11: op1_05_in02 = imem00_in[59:56];
    12: op1_05_in02 = reg_0729;
    4: op1_05_in02 = imem07_in[95:92];
    13: op1_05_in02 = reg_0324;
    14: op1_05_in02 = reg_0967;
    15: op1_05_in02 = imem07_in[31:28];
    16: op1_05_in02 = reg_0115;
    17: op1_05_in02 = reg_0396;
    18: op1_05_in02 = reg_0696;
    19: op1_05_in02 = imem04_in[63:60];
    3: op1_05_in02 = imem07_in[35:32];
    20: op1_05_in02 = reg_0684;
    21: op1_05_in02 = imem04_in[47:44];
    22: op1_05_in02 = imem00_in[55:52];
    44: op1_05_in02 = imem00_in[55:52];
    23: op1_05_in02 = imem00_in[39:36];
    24: op1_05_in02 = reg_0624;
    32: op1_05_in02 = reg_0624;
    25: op1_05_in02 = reg_1040;
    26: op1_05_in02 = imem04_in[15:12];
    27: op1_05_in02 = imem02_in[15:12];
    28: op1_05_in02 = reg_0749;
    29: op1_05_in02 = imem00_in[95:92];
    30: op1_05_in02 = imem00_in[87:84];
    31: op1_05_in02 = reg_0833;
    33: op1_05_in02 = imem00_in[43:40];
    34: op1_05_in02 = reg_0642;
    35: op1_05_in02 = reg_0443;
    36: op1_05_in02 = imem06_in[27:24];
    37: op1_05_in02 = reg_0429;
    38: op1_05_in02 = reg_0167;
    39: op1_05_in02 = reg_0693;
    40: op1_05_in02 = imem02_in[87:84];
    41: op1_05_in02 = imem00_in[115:112];
    42: op1_05_in02 = imem05_in[115:112];
    74: op1_05_in02 = imem05_in[115:112];
    43: op1_05_in02 = reg_0623;
    45: op1_05_in02 = reg_0346;
    46: op1_05_in02 = reg_0957;
    47: op1_05_in02 = imem00_in[67:64];
    95: op1_05_in02 = imem00_in[67:64];
    48: op1_05_in02 = reg_1041;
    49: op1_05_in02 = reg_0153;
    50: op1_05_in02 = reg_0511;
    51: op1_05_in02 = reg_1050;
    52: op1_05_in02 = imem00_in[91:88];
    53: op1_05_in02 = imem02_in[91:88];
    54: op1_05_in02 = reg_0793;
    55: op1_05_in02 = reg_0277;
    56: op1_05_in02 = reg_0809;
    57: op1_05_in02 = reg_0131;
    58: op1_05_in02 = reg_0361;
    59: op1_05_in02 = reg_0943;
    60: op1_05_in02 = imem00_in[83:80];
    61: op1_05_in02 = reg_0502;
    62: op1_05_in02 = reg_0683;
    63: op1_05_in02 = reg_0576;
    64: op1_05_in02 = imem04_in[67:64];
    65: op1_05_in02 = reg_0094;
    66: op1_05_in02 = reg_0152;
    67: op1_05_in02 = reg_0061;
    68: op1_05_in02 = reg_0698;
    69: op1_05_in02 = reg_0555;
    70: op1_05_in02 = imem04_in[3:0];
    71: op1_05_in02 = imem06_in[3:0];
    72: op1_05_in02 = reg_0989;
    73: op1_05_in02 = reg_0296;
    75: op1_05_in02 = reg_0704;
    76: op1_05_in02 = imem00_in[63:60];
    77: op1_05_in02 = reg_0768;
    78: op1_05_in02 = reg_0116;
    79: op1_05_in02 = reg_0932;
    80: op1_05_in02 = reg_0135;
    81: op1_05_in02 = reg_0591;
    82: op1_05_in02 = imem06_in[11:8];
    83: op1_05_in02 = imem02_in[67:64];
    84: op1_05_in02 = imem00_in[27:24];
    85: op1_05_in02 = imem05_in[3:0];
    86: op1_05_in02 = reg_0442;
    87: op1_05_in02 = reg_0772;
    88: op1_05_in02 = imem04_in[91:88];
    89: op1_05_in02 = imem00_in[75:72];
    90: op1_05_in02 = reg_0140;
    91: op1_05_in02 = reg_0960;
    92: op1_05_in02 = reg_0965;
    93: op1_05_in02 = imem00_in[19:16];
    94: op1_05_in02 = reg_0762;
    96: op1_05_in02 = reg_0186;
    97: op1_05_in02 = imem07_in[103:100];
    default: op1_05_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv02 = 1;
    11: op1_05_inv02 = 1;
    13: op1_05_inv02 = 1;
    16: op1_05_inv02 = 1;
    17: op1_05_inv02 = 1;
    18: op1_05_inv02 = 1;
    19: op1_05_inv02 = 1;
    20: op1_05_inv02 = 1;
    22: op1_05_inv02 = 1;
    23: op1_05_inv02 = 1;
    24: op1_05_inv02 = 1;
    26: op1_05_inv02 = 1;
    27: op1_05_inv02 = 1;
    28: op1_05_inv02 = 1;
    29: op1_05_inv02 = 1;
    30: op1_05_inv02 = 1;
    31: op1_05_inv02 = 1;
    35: op1_05_inv02 = 1;
    38: op1_05_inv02 = 1;
    40: op1_05_inv02 = 1;
    41: op1_05_inv02 = 1;
    43: op1_05_inv02 = 1;
    44: op1_05_inv02 = 1;
    45: op1_05_inv02 = 1;
    46: op1_05_inv02 = 1;
    49: op1_05_inv02 = 1;
    50: op1_05_inv02 = 1;
    52: op1_05_inv02 = 1;
    53: op1_05_inv02 = 1;
    54: op1_05_inv02 = 1;
    55: op1_05_inv02 = 1;
    56: op1_05_inv02 = 1;
    59: op1_05_inv02 = 1;
    60: op1_05_inv02 = 1;
    63: op1_05_inv02 = 1;
    64: op1_05_inv02 = 1;
    66: op1_05_inv02 = 1;
    68: op1_05_inv02 = 1;
    70: op1_05_inv02 = 1;
    71: op1_05_inv02 = 1;
    72: op1_05_inv02 = 1;
    74: op1_05_inv02 = 1;
    75: op1_05_inv02 = 1;
    77: op1_05_inv02 = 1;
    78: op1_05_inv02 = 1;
    79: op1_05_inv02 = 1;
    82: op1_05_inv02 = 1;
    83: op1_05_inv02 = 1;
    86: op1_05_inv02 = 1;
    89: op1_05_inv02 = 1;
    91: op1_05_inv02 = 1;
    92: op1_05_inv02 = 1;
    93: op1_05_inv02 = 1;
    95: op1_05_inv02 = 1;
    97: op1_05_inv02 = 1;
    default: op1_05_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in03 = imem00_in[55:52];
    84: op1_05_in03 = imem00_in[55:52];
    6: op1_05_in03 = reg_0035;
    7: op1_05_in03 = imem02_in[19:16];
    8: op1_05_in03 = reg_0271;
    9: op1_05_in03 = reg_0681;
    10: op1_05_in03 = reg_0617;
    11: op1_05_in03 = imem00_in[99:96];
    12: op1_05_in03 = reg_0713;
    4: op1_05_in03 = reg_0424;
    13: op1_05_in03 = reg_0083;
    14: op1_05_in03 = reg_0954;
    15: op1_05_in03 = imem07_in[39:36];
    16: op1_05_in03 = reg_0113;
    17: op1_05_in03 = reg_0374;
    18: op1_05_in03 = reg_0672;
    19: op1_05_in03 = imem04_in[95:92];
    88: op1_05_in03 = imem04_in[95:92];
    3: op1_05_in03 = imem07_in[59:56];
    20: op1_05_in03 = reg_0690;
    21: op1_05_in03 = imem04_in[67:64];
    22: op1_05_in03 = imem00_in[91:88];
    23: op1_05_in03 = imem00_in[43:40];
    24: op1_05_in03 = reg_0620;
    25: op1_05_in03 = reg_0116;
    26: op1_05_in03 = imem04_in[19:16];
    27: op1_05_in03 = imem02_in[51:48];
    28: op1_05_in03 = reg_0323;
    29: op1_05_in03 = imem00_in[103:100];
    30: op1_05_in03 = imem00_in[127:124];
    31: op1_05_in03 = reg_0373;
    32: op1_05_in03 = reg_0613;
    33: op1_05_in03 = imem00_in[47:44];
    34: op1_05_in03 = reg_0656;
    35: op1_05_in03 = reg_0181;
    36: op1_05_in03 = imem06_in[55:52];
    37: op1_05_in03 = reg_0432;
    38: op1_05_in03 = reg_0163;
    39: op1_05_in03 = reg_0697;
    40: op1_05_in03 = imem02_in[111:108];
    41: op1_05_in03 = reg_0696;
    42: op1_05_in03 = imem05_in[123:120];
    43: op1_05_in03 = reg_0717;
    44: op1_05_in03 = imem00_in[67:64];
    45: op1_05_in03 = reg_0847;
    46: op1_05_in03 = reg_0948;
    47: op1_05_in03 = imem00_in[83:80];
    48: op1_05_in03 = reg_0103;
    49: op1_05_in03 = reg_0141;
    50: op1_05_in03 = reg_0937;
    51: op1_05_in03 = reg_0317;
    52: op1_05_in03 = reg_0682;
    53: op1_05_in03 = imem02_in[103:100];
    54: op1_05_in03 = reg_0836;
    55: op1_05_in03 = reg_0539;
    56: op1_05_in03 = reg_0732;
    57: op1_05_in03 = imem06_in[47:44];
    58: op1_05_in03 = reg_0303;
    59: op1_05_in03 = reg_0057;
    60: op1_05_in03 = imem00_in[107:104];
    61: op1_05_in03 = reg_0868;
    62: op1_05_in03 = reg_0825;
    63: op1_05_in03 = reg_0923;
    64: op1_05_in03 = imem04_in[111:108];
    65: op1_05_in03 = reg_0448;
    66: op1_05_in03 = reg_0156;
    67: op1_05_in03 = reg_0027;
    68: op1_05_in03 = reg_0804;
    81: op1_05_in03 = reg_0804;
    69: op1_05_in03 = reg_0117;
    70: op1_05_in03 = imem04_in[31:28];
    71: op1_05_in03 = imem06_in[31:28];
    72: op1_05_in03 = reg_0974;
    73: op1_05_in03 = reg_0658;
    74: op1_05_in03 = imem06_in[7:4];
    75: op1_05_in03 = reg_0678;
    76: op1_05_in03 = reg_0685;
    77: op1_05_in03 = reg_0686;
    78: op1_05_in03 = reg_0733;
    79: op1_05_in03 = reg_0537;
    80: op1_05_in03 = reg_0508;
    82: op1_05_in03 = imem06_in[23:20];
    83: op1_05_in03 = imem02_in[115:112];
    85: op1_05_in03 = imem05_in[11:8];
    86: op1_05_in03 = reg_0805;
    87: op1_05_in03 = reg_0650;
    89: op1_05_in03 = reg_0738;
    96: op1_05_in03 = reg_0738;
    90: op1_05_in03 = reg_0947;
    91: op1_05_in03 = reg_0970;
    92: op1_05_in03 = reg_0657;
    93: op1_05_in03 = imem00_in[31:28];
    94: op1_05_in03 = reg_0521;
    95: op1_05_in03 = imem00_in[79:76];
    97: op1_05_in03 = imem07_in[107:104];
    default: op1_05_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv03 = 1;
    7: op1_05_inv03 = 1;
    8: op1_05_inv03 = 1;
    9: op1_05_inv03 = 1;
    10: op1_05_inv03 = 1;
    11: op1_05_inv03 = 1;
    12: op1_05_inv03 = 1;
    14: op1_05_inv03 = 1;
    16: op1_05_inv03 = 1;
    18: op1_05_inv03 = 1;
    21: op1_05_inv03 = 1;
    23: op1_05_inv03 = 1;
    26: op1_05_inv03 = 1;
    27: op1_05_inv03 = 1;
    31: op1_05_inv03 = 1;
    33: op1_05_inv03 = 1;
    38: op1_05_inv03 = 1;
    41: op1_05_inv03 = 1;
    48: op1_05_inv03 = 1;
    49: op1_05_inv03 = 1;
    51: op1_05_inv03 = 1;
    52: op1_05_inv03 = 1;
    53: op1_05_inv03 = 1;
    55: op1_05_inv03 = 1;
    58: op1_05_inv03 = 1;
    60: op1_05_inv03 = 1;
    61: op1_05_inv03 = 1;
    63: op1_05_inv03 = 1;
    64: op1_05_inv03 = 1;
    65: op1_05_inv03 = 1;
    67: op1_05_inv03 = 1;
    69: op1_05_inv03 = 1;
    70: op1_05_inv03 = 1;
    72: op1_05_inv03 = 1;
    73: op1_05_inv03 = 1;
    74: op1_05_inv03 = 1;
    75: op1_05_inv03 = 1;
    79: op1_05_inv03 = 1;
    83: op1_05_inv03 = 1;
    84: op1_05_inv03 = 1;
    86: op1_05_inv03 = 1;
    88: op1_05_inv03 = 1;
    89: op1_05_inv03 = 1;
    90: op1_05_inv03 = 1;
    91: op1_05_inv03 = 1;
    93: op1_05_inv03 = 1;
    94: op1_05_inv03 = 1;
    97: op1_05_inv03 = 1;
    default: op1_05_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in04 = imem00_in[107:104];
    6: op1_05_in04 = reg_0036;
    7: op1_05_in04 = imem02_in[111:108];
    8: op1_05_in04 = reg_0264;
    9: op1_05_in04 = reg_0696;
    10: op1_05_in04 = reg_0621;
    11: op1_05_in04 = imem00_in[123:120];
    12: op1_05_in04 = reg_0433;
    4: op1_05_in04 = reg_0429;
    13: op1_05_in04 = reg_0096;
    14: op1_05_in04 = reg_0956;
    15: op1_05_in04 = imem07_in[79:76];
    16: op1_05_in04 = imem02_in[7:4];
    17: op1_05_in04 = reg_0389;
    18: op1_05_in04 = reg_0687;
    19: op1_05_in04 = imem04_in[119:116];
    3: op1_05_in04 = imem07_in[75:72];
    20: op1_05_in04 = reg_0691;
    21: op1_05_in04 = imem04_in[71:68];
    22: op1_05_in04 = imem00_in[111:108];
    23: op1_05_in04 = imem00_in[47:44];
    24: op1_05_in04 = reg_0606;
    25: op1_05_in04 = imem02_in[51:48];
    26: op1_05_in04 = imem04_in[83:80];
    27: op1_05_in04 = imem02_in[71:68];
    28: op1_05_in04 = reg_0558;
    29: op1_05_in04 = reg_0695;
    30: op1_05_in04 = reg_0690;
    31: op1_05_in04 = reg_0807;
    32: op1_05_in04 = reg_0617;
    33: op1_05_in04 = imem00_in[51:48];
    34: op1_05_in04 = reg_0647;
    35: op1_05_in04 = reg_0161;
    36: op1_05_in04 = imem06_in[91:88];
    37: op1_05_in04 = reg_0436;
    38: op1_05_in04 = reg_0168;
    39: op1_05_in04 = reg_0676;
    40: op1_05_in04 = imem02_in[127:124];
    41: op1_05_in04 = reg_0672;
    42: op1_05_in04 = imem05_in[127:124];
    43: op1_05_in04 = reg_0708;
    44: op1_05_in04 = imem00_in[71:68];
    45: op1_05_in04 = reg_0923;
    46: op1_05_in04 = reg_0942;
    47: op1_05_in04 = imem00_in[119:116];
    60: op1_05_in04 = imem00_in[119:116];
    48: op1_05_in04 = reg_0116;
    49: op1_05_in04 = reg_0131;
    50: op1_05_in04 = reg_1057;
    51: op1_05_in04 = reg_0397;
    52: op1_05_in04 = reg_0683;
    53: op1_05_in04 = reg_0655;
    54: op1_05_in04 = reg_0312;
    55: op1_05_in04 = reg_0068;
    56: op1_05_in04 = reg_0281;
    57: op1_05_in04 = imem06_in[59:56];
    58: op1_05_in04 = reg_0421;
    59: op1_05_in04 = reg_0488;
    61: op1_05_in04 = reg_0640;
    62: op1_05_in04 = reg_0748;
    63: op1_05_in04 = reg_0038;
    64: op1_05_in04 = reg_1004;
    65: op1_05_in04 = reg_0489;
    66: op1_05_in04 = reg_0154;
    67: op1_05_in04 = reg_0777;
    68: op1_05_in04 = reg_0011;
    81: op1_05_in04 = reg_0011;
    69: op1_05_in04 = reg_0821;
    70: op1_05_in04 = imem04_in[55:52];
    71: op1_05_in04 = imem06_in[55:52];
    72: op1_05_in04 = reg_0997;
    73: op1_05_in04 = reg_0444;
    74: op1_05_in04 = imem06_in[11:8];
    75: op1_05_in04 = reg_0822;
    76: op1_05_in04 = reg_0825;
    77: op1_05_in04 = reg_0842;
    78: op1_05_in04 = reg_0115;
    79: op1_05_in04 = reg_0313;
    80: op1_05_in04 = reg_0706;
    82: op1_05_in04 = imem06_in[31:28];
    83: op1_05_in04 = reg_0908;
    84: op1_05_in04 = reg_0001;
    85: op1_05_in04 = imem05_in[27:24];
    86: op1_05_in04 = reg_0575;
    87: op1_05_in04 = reg_0775;
    88: op1_05_in04 = reg_0577;
    89: op1_05_in04 = reg_0883;
    90: op1_05_in04 = reg_0813;
    91: op1_05_in04 = reg_0949;
    92: op1_05_in04 = reg_0144;
    93: op1_05_in04 = imem00_in[43:40];
    94: op1_05_in04 = reg_0030;
    95: op1_05_in04 = imem00_in[83:80];
    96: op1_05_in04 = reg_0699;
    97: op1_05_in04 = reg_0717;
    default: op1_05_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv04 = 1;
    8: op1_05_inv04 = 1;
    9: op1_05_inv04 = 1;
    10: op1_05_inv04 = 1;
    13: op1_05_inv04 = 1;
    15: op1_05_inv04 = 1;
    18: op1_05_inv04 = 1;
    19: op1_05_inv04 = 1;
    20: op1_05_inv04 = 1;
    21: op1_05_inv04 = 1;
    25: op1_05_inv04 = 1;
    26: op1_05_inv04 = 1;
    27: op1_05_inv04 = 1;
    31: op1_05_inv04 = 1;
    32: op1_05_inv04 = 1;
    34: op1_05_inv04 = 1;
    38: op1_05_inv04 = 1;
    39: op1_05_inv04 = 1;
    41: op1_05_inv04 = 1;
    42: op1_05_inv04 = 1;
    43: op1_05_inv04 = 1;
    44: op1_05_inv04 = 1;
    47: op1_05_inv04 = 1;
    48: op1_05_inv04 = 1;
    52: op1_05_inv04 = 1;
    53: op1_05_inv04 = 1;
    55: op1_05_inv04 = 1;
    59: op1_05_inv04 = 1;
    61: op1_05_inv04 = 1;
    62: op1_05_inv04 = 1;
    63: op1_05_inv04 = 1;
    64: op1_05_inv04 = 1;
    65: op1_05_inv04 = 1;
    68: op1_05_inv04 = 1;
    70: op1_05_inv04 = 1;
    78: op1_05_inv04 = 1;
    79: op1_05_inv04 = 1;
    82: op1_05_inv04 = 1;
    85: op1_05_inv04 = 1;
    88: op1_05_inv04 = 1;
    89: op1_05_inv04 = 1;
    92: op1_05_inv04 = 1;
    93: op1_05_inv04 = 1;
    95: op1_05_inv04 = 1;
    96: op1_05_inv04 = 1;
    97: op1_05_inv04 = 1;
    default: op1_05_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in05 = imem00_in[115:112];
    22: op1_05_in05 = imem00_in[115:112];
    95: op1_05_in05 = imem00_in[115:112];
    6: op1_05_in05 = reg_0021;
    7: op1_05_in05 = imem02_in[115:112];
    8: op1_05_in05 = reg_0229;
    9: op1_05_in05 = reg_0689;
    10: op1_05_in05 = reg_0616;
    32: op1_05_in05 = reg_0616;
    11: op1_05_in05 = reg_0675;
    12: op1_05_in05 = reg_0426;
    4: op1_05_in05 = reg_0436;
    13: op1_05_in05 = reg_0090;
    14: op1_05_in05 = reg_0957;
    15: op1_05_in05 = imem07_in[87:84];
    16: op1_05_in05 = imem02_in[35:32];
    17: op1_05_in05 = reg_0985;
    18: op1_05_in05 = reg_0699;
    19: op1_05_in05 = reg_0283;
    3: op1_05_in05 = imem07_in[127:124];
    20: op1_05_in05 = reg_0688;
    21: op1_05_in05 = imem04_in[127:124];
    23: op1_05_in05 = imem00_in[55:52];
    24: op1_05_in05 = reg_0609;
    25: op1_05_in05 = imem02_in[55:52];
    26: op1_05_in05 = imem04_in[99:96];
    27: op1_05_in05 = imem02_in[103:100];
    28: op1_05_in05 = reg_0551;
    29: op1_05_in05 = reg_0682;
    30: op1_05_in05 = reg_0454;
    31: op1_05_in05 = reg_0376;
    33: op1_05_in05 = imem00_in[83:80];
    34: op1_05_in05 = reg_0636;
    35: op1_05_in05 = reg_0183;
    36: op1_05_in05 = imem06_in[95:92];
    37: op1_05_in05 = reg_0422;
    38: op1_05_in05 = reg_0157;
    39: op1_05_in05 = reg_0686;
    40: op1_05_in05 = reg_0653;
    41: op1_05_in05 = reg_0694;
    42: op1_05_in05 = reg_0973;
    43: op1_05_in05 = reg_0715;
    44: op1_05_in05 = imem00_in[99:96];
    45: op1_05_in05 = reg_0038;
    46: op1_05_in05 = reg_0949;
    47: op1_05_in05 = reg_0693;
    48: op1_05_in05 = reg_0117;
    49: op1_05_in05 = imem06_in[11:8];
    50: op1_05_in05 = reg_1020;
    51: op1_05_in05 = reg_0823;
    52: op1_05_in05 = reg_0469;
    53: op1_05_in05 = reg_0649;
    54: op1_05_in05 = reg_0844;
    55: op1_05_in05 = reg_0015;
    56: op1_05_in05 = reg_0578;
    57: op1_05_in05 = imem06_in[71:68];
    58: op1_05_in05 = reg_0532;
    59: op1_05_in05 = reg_0446;
    60: op1_05_in05 = reg_0523;
    61: op1_05_in05 = reg_0838;
    62: op1_05_in05 = reg_0900;
    63: op1_05_in05 = reg_0807;
    64: op1_05_in05 = reg_0282;
    65: op1_05_in05 = reg_0150;
    66: op1_05_in05 = reg_0155;
    67: op1_05_in05 = reg_0856;
    68: op1_05_in05 = reg_0222;
    69: op1_05_in05 = imem02_in[75:72];
    70: op1_05_in05 = imem04_in[119:116];
    71: op1_05_in05 = imem06_in[83:80];
    72: op1_05_in05 = reg_0994;
    73: op1_05_in05 = reg_0824;
    74: op1_05_in05 = imem06_in[43:40];
    75: op1_05_in05 = reg_0705;
    76: op1_05_in05 = reg_0738;
    77: op1_05_in05 = reg_0102;
    78: op1_05_in05 = reg_0113;
    79: op1_05_in05 = reg_0276;
    80: op1_05_in05 = reg_0326;
    81: op1_05_in05 = reg_0220;
    82: op1_05_in05 = imem06_in[103:100];
    83: op1_05_in05 = reg_0739;
    84: op1_05_in05 = reg_0825;
    85: op1_05_in05 = imem05_in[35:32];
    86: op1_05_in05 = reg_0421;
    87: op1_05_in05 = reg_0656;
    88: op1_05_in05 = reg_0511;
    89: op1_05_in05 = reg_0356;
    90: op1_05_in05 = reg_0831;
    91: op1_05_in05 = reg_0741;
    92: op1_05_in05 = imem06_in[3:0];
    93: op1_05_in05 = imem00_in[71:68];
    94: op1_05_in05 = reg_0455;
    96: op1_05_in05 = reg_0465;
    97: op1_05_in05 = reg_0374;
    default: op1_05_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv05 = 1;
    10: op1_05_inv05 = 1;
    12: op1_05_inv05 = 1;
    4: op1_05_inv05 = 1;
    13: op1_05_inv05 = 1;
    14: op1_05_inv05 = 1;
    15: op1_05_inv05 = 1;
    16: op1_05_inv05 = 1;
    17: op1_05_inv05 = 1;
    3: op1_05_inv05 = 1;
    20: op1_05_inv05 = 1;
    24: op1_05_inv05 = 1;
    25: op1_05_inv05 = 1;
    28: op1_05_inv05 = 1;
    30: op1_05_inv05 = 1;
    34: op1_05_inv05 = 1;
    35: op1_05_inv05 = 1;
    36: op1_05_inv05 = 1;
    41: op1_05_inv05 = 1;
    43: op1_05_inv05 = 1;
    44: op1_05_inv05 = 1;
    50: op1_05_inv05 = 1;
    51: op1_05_inv05 = 1;
    53: op1_05_inv05 = 1;
    56: op1_05_inv05 = 1;
    59: op1_05_inv05 = 1;
    64: op1_05_inv05 = 1;
    65: op1_05_inv05 = 1;
    70: op1_05_inv05 = 1;
    72: op1_05_inv05 = 1;
    73: op1_05_inv05 = 1;
    75: op1_05_inv05 = 1;
    80: op1_05_inv05 = 1;
    81: op1_05_inv05 = 1;
    82: op1_05_inv05 = 1;
    88: op1_05_inv05 = 1;
    89: op1_05_inv05 = 1;
    90: op1_05_inv05 = 1;
    95: op1_05_inv05 = 1;
    default: op1_05_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in06 = reg_0674;
    6: op1_05_in06 = reg_0029;
    7: op1_05_in06 = imem02_in[119:116];
    8: op1_05_in06 = reg_0260;
    9: op1_05_in06 = reg_0671;
    10: op1_05_in06 = reg_0626;
    11: op1_05_in06 = reg_0687;
    77: op1_05_in06 = reg_0687;
    12: op1_05_in06 = reg_0447;
    4: op1_05_in06 = reg_0447;
    13: op1_05_in06 = reg_0051;
    14: op1_05_in06 = reg_0949;
    42: op1_05_in06 = reg_0949;
    15: op1_05_in06 = imem07_in[95:92];
    16: op1_05_in06 = imem02_in[43:40];
    17: op1_05_in06 = reg_0991;
    18: op1_05_in06 = reg_0463;
    19: op1_05_in06 = reg_0517;
    3: op1_05_in06 = reg_0180;
    20: op1_05_in06 = reg_0673;
    21: op1_05_in06 = reg_0545;
    81: op1_05_in06 = reg_0545;
    22: op1_05_in06 = reg_0682;
    23: op1_05_in06 = imem00_in[63:60];
    24: op1_05_in06 = reg_0632;
    25: op1_05_in06 = imem02_in[67:64];
    26: op1_05_in06 = imem04_in[103:100];
    27: op1_05_in06 = reg_0658;
    28: op1_05_in06 = reg_0582;
    29: op1_05_in06 = reg_0698;
    30: op1_05_in06 = reg_0450;
    31: op1_05_in06 = reg_0844;
    32: op1_05_in06 = reg_0631;
    33: op1_05_in06 = imem00_in[87:84];
    34: op1_05_in06 = reg_0667;
    35: op1_05_in06 = reg_0171;
    36: op1_05_in06 = imem06_in[99:96];
    37: op1_05_in06 = reg_0433;
    39: op1_05_in06 = reg_0670;
    40: op1_05_in06 = reg_0654;
    41: op1_05_in06 = reg_0668;
    62: op1_05_in06 = reg_0668;
    43: op1_05_in06 = reg_0701;
    44: op1_05_in06 = imem00_in[119:116];
    45: op1_05_in06 = reg_0311;
    46: op1_05_in06 = reg_0952;
    47: op1_05_in06 = reg_0681;
    48: op1_05_in06 = reg_0126;
    49: op1_05_in06 = imem06_in[55:52];
    74: op1_05_in06 = imem06_in[55:52];
    50: op1_05_in06 = reg_0537;
    51: op1_05_in06 = reg_0543;
    52: op1_05_in06 = reg_0473;
    53: op1_05_in06 = reg_0647;
    54: op1_05_in06 = reg_0374;
    55: op1_05_in06 = reg_0444;
    56: op1_05_in06 = reg_0270;
    57: op1_05_in06 = imem06_in[87:84];
    58: op1_05_in06 = reg_0599;
    59: op1_05_in06 = reg_0023;
    60: op1_05_in06 = reg_0748;
    61: op1_05_in06 = reg_0174;
    63: op1_05_in06 = reg_0518;
    64: op1_05_in06 = reg_1057;
    65: op1_05_in06 = reg_0146;
    66: op1_05_in06 = reg_0144;
    67: op1_05_in06 = imem05_in[19:16];
    68: op1_05_in06 = reg_0946;
    69: op1_05_in06 = imem02_in[107:104];
    70: op1_05_in06 = reg_0483;
    71: op1_05_in06 = imem06_in[103:100];
    72: op1_05_in06 = imem04_in[7:4];
    73: op1_05_in06 = reg_0958;
    75: op1_05_in06 = reg_0437;
    76: op1_05_in06 = reg_0356;
    78: op1_05_in06 = reg_0821;
    79: op1_05_in06 = reg_0584;
    80: op1_05_in06 = imem06_in[19:16];
    82: op1_05_in06 = imem06_in[107:104];
    83: op1_05_in06 = reg_0394;
    84: op1_05_in06 = reg_0843;
    85: op1_05_in06 = imem05_in[79:76];
    86: op1_05_in06 = reg_0428;
    87: op1_05_in06 = reg_0643;
    88: op1_05_in06 = reg_0156;
    89: op1_05_in06 = reg_0480;
    90: op1_05_in06 = reg_0709;
    91: op1_05_in06 = reg_0657;
    92: op1_05_in06 = imem06_in[71:68];
    93: op1_05_in06 = imem00_in[83:80];
    94: op1_05_in06 = reg_0464;
    95: op1_05_in06 = imem00_in[127:124];
    96: op1_05_in06 = reg_0469;
    97: op1_05_in06 = reg_0560;
    default: op1_05_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv06 = 1;
    6: op1_05_inv06 = 1;
    7: op1_05_inv06 = 1;
    9: op1_05_inv06 = 1;
    11: op1_05_inv06 = 1;
    4: op1_05_inv06 = 1;
    13: op1_05_inv06 = 1;
    16: op1_05_inv06 = 1;
    18: op1_05_inv06 = 1;
    20: op1_05_inv06 = 1;
    21: op1_05_inv06 = 1;
    25: op1_05_inv06 = 1;
    27: op1_05_inv06 = 1;
    31: op1_05_inv06 = 1;
    32: op1_05_inv06 = 1;
    33: op1_05_inv06 = 1;
    34: op1_05_inv06 = 1;
    35: op1_05_inv06 = 1;
    39: op1_05_inv06 = 1;
    43: op1_05_inv06 = 1;
    45: op1_05_inv06 = 1;
    47: op1_05_inv06 = 1;
    51: op1_05_inv06 = 1;
    54: op1_05_inv06 = 1;
    56: op1_05_inv06 = 1;
    58: op1_05_inv06 = 1;
    60: op1_05_inv06 = 1;
    62: op1_05_inv06 = 1;
    63: op1_05_inv06 = 1;
    64: op1_05_inv06 = 1;
    66: op1_05_inv06 = 1;
    69: op1_05_inv06 = 1;
    71: op1_05_inv06 = 1;
    75: op1_05_inv06 = 1;
    77: op1_05_inv06 = 1;
    81: op1_05_inv06 = 1;
    88: op1_05_inv06 = 1;
    90: op1_05_inv06 = 1;
    92: op1_05_inv06 = 1;
    93: op1_05_inv06 = 1;
    95: op1_05_inv06 = 1;
    96: op1_05_inv06 = 1;
    default: op1_05_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in07 = reg_0475;
    6: op1_05_in07 = reg_0022;
    7: op1_05_in07 = reg_0357;
    8: op1_05_in07 = reg_0265;
    9: op1_05_in07 = reg_0680;
    76: op1_05_in07 = reg_0680;
    10: op1_05_in07 = reg_0615;
    11: op1_05_in07 = reg_0692;
    12: op1_05_in07 = reg_0419;
    4: op1_05_in07 = reg_0418;
    13: op1_05_in07 = reg_0094;
    14: op1_05_in07 = reg_0945;
    15: op1_05_in07 = imem07_in[107:104];
    16: op1_05_in07 = imem02_in[51:48];
    17: op1_05_in07 = reg_0992;
    18: op1_05_in07 = reg_0464;
    19: op1_05_in07 = reg_0056;
    3: op1_05_in07 = reg_0172;
    20: op1_05_in07 = reg_0687;
    21: op1_05_in07 = reg_0557;
    22: op1_05_in07 = reg_0683;
    23: op1_05_in07 = imem00_in[67:64];
    24: op1_05_in07 = reg_0402;
    25: op1_05_in07 = imem02_in[87:84];
    26: op1_05_in07 = imem04_in[111:108];
    27: op1_05_in07 = reg_0660;
    28: op1_05_in07 = reg_0593;
    29: op1_05_in07 = reg_0679;
    30: op1_05_in07 = reg_0455;
    31: op1_05_in07 = reg_0991;
    32: op1_05_in07 = reg_0381;
    33: op1_05_in07 = imem00_in[91:88];
    34: op1_05_in07 = reg_0663;
    36: op1_05_in07 = imem06_in[115:112];
    37: op1_05_in07 = reg_0421;
    39: op1_05_in07 = reg_0690;
    40: op1_05_in07 = reg_0639;
    41: op1_05_in07 = reg_0465;
    42: op1_05_in07 = reg_0965;
    43: op1_05_in07 = imem07_in[3:0];
    71: op1_05_in07 = imem07_in[3:0];
    75: op1_05_in07 = imem07_in[3:0];
    44: op1_05_in07 = imem00_in[123:120];
    45: op1_05_in07 = reg_0836;
    46: op1_05_in07 = reg_0821;
    47: op1_05_in07 = reg_0672;
    48: op1_05_in07 = imem02_in[55:52];
    49: op1_05_in07 = imem06_in[87:84];
    50: op1_05_in07 = reg_0799;
    51: op1_05_in07 = reg_0312;
    52: op1_05_in07 = reg_0474;
    53: op1_05_in07 = reg_0854;
    54: op1_05_in07 = reg_0234;
    55: op1_05_in07 = reg_0429;
    56: op1_05_in07 = reg_0319;
    57: op1_05_in07 = reg_0914;
    58: op1_05_in07 = reg_0180;
    59: op1_05_in07 = reg_0435;
    60: op1_05_in07 = reg_0900;
    61: op1_05_in07 = reg_0175;
    62: op1_05_in07 = reg_0102;
    63: op1_05_in07 = reg_0513;
    64: op1_05_in07 = reg_1020;
    65: op1_05_in07 = reg_0139;
    66: op1_05_in07 = imem06_in[15:12];
    67: op1_05_in07 = imem05_in[59:56];
    68: op1_05_in07 = reg_0780;
    69: op1_05_in07 = reg_0653;
    70: op1_05_in07 = reg_0937;
    72: op1_05_in07 = imem04_in[63:60];
    73: op1_05_in07 = reg_0133;
    74: op1_05_in07 = imem06_in[103:100];
    77: op1_05_in07 = reg_0749;
    78: op1_05_in07 = reg_0110;
    79: op1_05_in07 = reg_0658;
    80: op1_05_in07 = imem06_in[23:20];
    81: op1_05_in07 = reg_0566;
    82: op1_05_in07 = imem06_in[111:108];
    83: op1_05_in07 = reg_0389;
    84: op1_05_in07 = reg_0523;
    85: op1_05_in07 = imem05_in[91:88];
    86: op1_05_in07 = reg_0532;
    87: op1_05_in07 = reg_0493;
    88: op1_05_in07 = reg_0912;
    89: op1_05_in07 = reg_0467;
    90: op1_05_in07 = reg_0508;
    91: op1_05_in07 = imem06_in[31:28];
    92: op1_05_in07 = reg_0244;
    93: op1_05_in07 = imem00_in[115:112];
    94: op1_05_in07 = reg_0462;
    95: op1_05_in07 = reg_0857;
    96: op1_05_in07 = reg_0466;
    97: op1_05_in07 = reg_0708;
    default: op1_05_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv07 = 1;
    7: op1_05_inv07 = 1;
    9: op1_05_inv07 = 1;
    11: op1_05_inv07 = 1;
    12: op1_05_inv07 = 1;
    14: op1_05_inv07 = 1;
    18: op1_05_inv07 = 1;
    19: op1_05_inv07 = 1;
    21: op1_05_inv07 = 1;
    24: op1_05_inv07 = 1;
    28: op1_05_inv07 = 1;
    29: op1_05_inv07 = 1;
    32: op1_05_inv07 = 1;
    37: op1_05_inv07 = 1;
    40: op1_05_inv07 = 1;
    41: op1_05_inv07 = 1;
    44: op1_05_inv07 = 1;
    45: op1_05_inv07 = 1;
    48: op1_05_inv07 = 1;
    51: op1_05_inv07 = 1;
    52: op1_05_inv07 = 1;
    54: op1_05_inv07 = 1;
    56: op1_05_inv07 = 1;
    57: op1_05_inv07 = 1;
    59: op1_05_inv07 = 1;
    60: op1_05_inv07 = 1;
    65: op1_05_inv07 = 1;
    67: op1_05_inv07 = 1;
    68: op1_05_inv07 = 1;
    71: op1_05_inv07 = 1;
    72: op1_05_inv07 = 1;
    74: op1_05_inv07 = 1;
    81: op1_05_inv07 = 1;
    82: op1_05_inv07 = 1;
    84: op1_05_inv07 = 1;
    85: op1_05_inv07 = 1;
    87: op1_05_inv07 = 1;
    88: op1_05_inv07 = 1;
    94: op1_05_inv07 = 1;
    95: op1_05_inv07 = 1;
    default: op1_05_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in08 = reg_0452;
    6: op1_05_in08 = imem07_in[11:8];
    7: op1_05_in08 = reg_0330;
    8: op1_05_in08 = reg_0255;
    9: op1_05_in08 = reg_0669;
    20: op1_05_in08 = reg_0669;
    10: op1_05_in08 = reg_0332;
    11: op1_05_in08 = reg_0463;
    12: op1_05_in08 = reg_0444;
    4: op1_05_in08 = reg_0437;
    13: op1_05_in08 = imem03_in[27:24];
    14: op1_05_in08 = reg_0943;
    15: op1_05_in08 = reg_0728;
    16: op1_05_in08 = reg_0650;
    17: op1_05_in08 = reg_0979;
    18: op1_05_in08 = reg_0466;
    19: op1_05_in08 = reg_0043;
    3: op1_05_in08 = reg_0165;
    61: op1_05_in08 = reg_0165;
    21: op1_05_in08 = reg_0548;
    22: op1_05_in08 = reg_0676;
    44: op1_05_in08 = reg_0676;
    47: op1_05_in08 = reg_0676;
    23: op1_05_in08 = imem00_in[87:84];
    24: op1_05_in08 = reg_0372;
    25: op1_05_in08 = reg_0665;
    26: op1_05_in08 = reg_0483;
    27: op1_05_in08 = reg_0639;
    28: op1_05_in08 = reg_0576;
    29: op1_05_in08 = reg_0691;
    30: op1_05_in08 = reg_0461;
    41: op1_05_in08 = reg_0461;
    31: op1_05_in08 = reg_0992;
    32: op1_05_in08 = reg_0383;
    33: op1_05_in08 = imem00_in[111:108];
    34: op1_05_in08 = reg_0334;
    36: op1_05_in08 = reg_0386;
    57: op1_05_in08 = reg_0386;
    37: op1_05_in08 = reg_0419;
    39: op1_05_in08 = reg_0677;
    40: op1_05_in08 = reg_0648;
    42: op1_05_in08 = reg_0952;
    43: op1_05_in08 = imem07_in[51:48];
    45: op1_05_in08 = reg_0844;
    46: op1_05_in08 = reg_0813;
    48: op1_05_in08 = imem02_in[71:68];
    49: op1_05_in08 = imem06_in[103:100];
    50: op1_05_in08 = reg_0848;
    51: op1_05_in08 = reg_0513;
    52: op1_05_in08 = reg_0187;
    53: op1_05_in08 = reg_0837;
    54: op1_05_in08 = reg_0822;
    55: op1_05_in08 = reg_0882;
    56: op1_05_in08 = reg_0949;
    58: op1_05_in08 = reg_0185;
    59: op1_05_in08 = reg_1046;
    60: op1_05_in08 = reg_0356;
    62: op1_05_in08 = reg_0663;
    63: op1_05_in08 = reg_0234;
    64: op1_05_in08 = reg_0050;
    65: op1_05_in08 = reg_0137;
    66: op1_05_in08 = imem06_in[31:28];
    80: op1_05_in08 = imem06_in[31:28];
    67: op1_05_in08 = imem05_in[87:84];
    68: op1_05_in08 = reg_0264;
    69: op1_05_in08 = reg_0290;
    70: op1_05_in08 = reg_1005;
    71: op1_05_in08 = imem07_in[15:12];
    72: op1_05_in08 = imem04_in[75:72];
    73: op1_05_in08 = reg_0959;
    74: op1_05_in08 = imem06_in[127:124];
    75: op1_05_in08 = imem07_in[63:60];
    76: op1_05_in08 = reg_0828;
    77: op1_05_in08 = reg_0453;
    78: op1_05_in08 = imem02_in[15:12];
    79: op1_05_in08 = reg_0070;
    81: op1_05_in08 = reg_0678;
    82: op1_05_in08 = imem06_in[119:116];
    83: op1_05_in08 = reg_0335;
    84: op1_05_in08 = reg_0686;
    85: op1_05_in08 = reg_0215;
    86: op1_05_in08 = reg_0024;
    87: op1_05_in08 = imem03_in[15:12];
    88: op1_05_in08 = reg_0540;
    89: op1_05_in08 = reg_0456;
    90: op1_05_in08 = reg_0951;
    91: op1_05_in08 = imem06_in[35:32];
    92: op1_05_in08 = reg_0393;
    93: op1_05_in08 = reg_0684;
    94: op1_05_in08 = reg_0474;
    95: op1_05_in08 = reg_0009;
    96: op1_05_in08 = reg_0473;
    97: op1_05_in08 = reg_0718;
    default: op1_05_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv08 = 1;
    7: op1_05_inv08 = 1;
    9: op1_05_inv08 = 1;
    10: op1_05_inv08 = 1;
    11: op1_05_inv08 = 1;
    12: op1_05_inv08 = 1;
    4: op1_05_inv08 = 1;
    13: op1_05_inv08 = 1;
    21: op1_05_inv08 = 1;
    23: op1_05_inv08 = 1;
    25: op1_05_inv08 = 1;
    29: op1_05_inv08 = 1;
    39: op1_05_inv08 = 1;
    40: op1_05_inv08 = 1;
    47: op1_05_inv08 = 1;
    50: op1_05_inv08 = 1;
    55: op1_05_inv08 = 1;
    56: op1_05_inv08 = 1;
    57: op1_05_inv08 = 1;
    58: op1_05_inv08 = 1;
    59: op1_05_inv08 = 1;
    60: op1_05_inv08 = 1;
    63: op1_05_inv08 = 1;
    67: op1_05_inv08 = 1;
    68: op1_05_inv08 = 1;
    72: op1_05_inv08 = 1;
    73: op1_05_inv08 = 1;
    74: op1_05_inv08 = 1;
    77: op1_05_inv08 = 1;
    85: op1_05_inv08 = 1;
    86: op1_05_inv08 = 1;
    87: op1_05_inv08 = 1;
    90: op1_05_inv08 = 1;
    92: op1_05_inv08 = 1;
    94: op1_05_inv08 = 1;
    97: op1_05_inv08 = 1;
    default: op1_05_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in09 = reg_0208;
    6: op1_05_in09 = imem07_in[15:12];
    7: op1_05_in09 = reg_0310;
    8: op1_05_in09 = reg_0145;
    9: op1_05_in09 = reg_0454;
    10: op1_05_in09 = reg_0381;
    11: op1_05_in09 = reg_0460;
    30: op1_05_in09 = reg_0460;
    12: op1_05_in09 = reg_0437;
    4: op1_05_in09 = reg_0175;
    13: op1_05_in09 = imem03_in[51:48];
    14: op1_05_in09 = reg_0863;
    15: op1_05_in09 = reg_0719;
    16: op1_05_in09 = reg_0656;
    17: op1_05_in09 = reg_0980;
    18: op1_05_in09 = reg_0473;
    19: op1_05_in09 = reg_0854;
    3: op1_05_in09 = reg_0162;
    20: op1_05_in09 = reg_0475;
    21: op1_05_in09 = reg_0554;
    22: op1_05_in09 = reg_0687;
    23: op1_05_in09 = imem00_in[91:88];
    24: op1_05_in09 = reg_1029;
    25: op1_05_in09 = reg_0663;
    26: op1_05_in09 = reg_0301;
    27: op1_05_in09 = reg_0638;
    28: op1_05_in09 = imem03_in[19:16];
    29: op1_05_in09 = reg_0674;
    31: op1_05_in09 = reg_0993;
    32: op1_05_in09 = reg_0399;
    33: op1_05_in09 = imem00_in[123:120];
    34: op1_05_in09 = reg_0916;
    36: op1_05_in09 = reg_0741;
    37: op1_05_in09 = reg_0439;
    39: op1_05_in09 = reg_0691;
    40: op1_05_in09 = reg_0641;
    41: op1_05_in09 = reg_0477;
    42: op1_05_in09 = reg_0953;
    43: op1_05_in09 = imem07_in[75:72];
    44: op1_05_in09 = reg_0684;
    45: op1_05_in09 = reg_0234;
    46: op1_05_in09 = reg_0257;
    47: op1_05_in09 = reg_0686;
    48: op1_05_in09 = imem02_in[95:92];
    49: op1_05_in09 = imem06_in[115:112];
    91: op1_05_in09 = imem06_in[115:112];
    50: op1_05_in09 = reg_0850;
    51: op1_05_in09 = reg_0844;
    52: op1_05_in09 = reg_0209;
    53: op1_05_in09 = reg_0664;
    54: op1_05_in09 = reg_0998;
    55: op1_05_in09 = imem05_in[23:20];
    56: op1_05_in09 = reg_0945;
    57: op1_05_in09 = reg_0295;
    58: op1_05_in09 = reg_0170;
    59: op1_05_in09 = reg_0489;
    60: op1_05_in09 = reg_0668;
    61: op1_05_in09 = reg_0161;
    62: op1_05_in09 = reg_0464;
    63: op1_05_in09 = reg_1002;
    64: op1_05_in09 = reg_0752;
    65: op1_05_in09 = imem06_in[11:8];
    66: op1_05_in09 = imem06_in[35:32];
    80: op1_05_in09 = imem06_in[35:32];
    67: op1_05_in09 = imem05_in[111:108];
    68: op1_05_in09 = reg_0633;
    69: op1_05_in09 = reg_0565;
    70: op1_05_in09 = reg_0931;
    71: op1_05_in09 = imem07_in[39:36];
    72: op1_05_in09 = imem04_in[103:100];
    73: op1_05_in09 = reg_0946;
    74: op1_05_in09 = reg_0010;
    75: op1_05_in09 = imem07_in[91:88];
    76: op1_05_in09 = reg_0457;
    77: op1_05_in09 = reg_0469;
    78: op1_05_in09 = imem02_in[35:32];
    79: op1_05_in09 = reg_0586;
    81: op1_05_in09 = reg_0713;
    82: op1_05_in09 = reg_0660;
    83: op1_05_in09 = reg_0054;
    84: op1_05_in09 = reg_0499;
    85: op1_05_in09 = reg_0142;
    86: op1_05_in09 = reg_0701;
    87: op1_05_in09 = imem03_in[59:56];
    88: op1_05_in09 = reg_0882;
    89: op1_05_in09 = reg_0214;
    90: op1_05_in09 = reg_0965;
    92: op1_05_in09 = reg_0754;
    93: op1_05_in09 = reg_0160;
    94: op1_05_in09 = reg_0479;
    95: op1_05_in09 = reg_0871;
    96: op1_05_in09 = reg_0467;
    97: op1_05_in09 = reg_0903;
    default: op1_05_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv09 = 1;
    11: op1_05_inv09 = 1;
    4: op1_05_inv09 = 1;
    14: op1_05_inv09 = 1;
    17: op1_05_inv09 = 1;
    18: op1_05_inv09 = 1;
    3: op1_05_inv09 = 1;
    21: op1_05_inv09 = 1;
    22: op1_05_inv09 = 1;
    23: op1_05_inv09 = 1;
    24: op1_05_inv09 = 1;
    25: op1_05_inv09 = 1;
    26: op1_05_inv09 = 1;
    27: op1_05_inv09 = 1;
    28: op1_05_inv09 = 1;
    33: op1_05_inv09 = 1;
    36: op1_05_inv09 = 1;
    41: op1_05_inv09 = 1;
    46: op1_05_inv09 = 1;
    48: op1_05_inv09 = 1;
    49: op1_05_inv09 = 1;
    53: op1_05_inv09 = 1;
    56: op1_05_inv09 = 1;
    58: op1_05_inv09 = 1;
    59: op1_05_inv09 = 1;
    60: op1_05_inv09 = 1;
    61: op1_05_inv09 = 1;
    62: op1_05_inv09 = 1;
    64: op1_05_inv09 = 1;
    67: op1_05_inv09 = 1;
    68: op1_05_inv09 = 1;
    70: op1_05_inv09 = 1;
    72: op1_05_inv09 = 1;
    74: op1_05_inv09 = 1;
    75: op1_05_inv09 = 1;
    78: op1_05_inv09 = 1;
    79: op1_05_inv09 = 1;
    81: op1_05_inv09 = 1;
    82: op1_05_inv09 = 1;
    83: op1_05_inv09 = 1;
    85: op1_05_inv09 = 1;
    86: op1_05_inv09 = 1;
    90: op1_05_inv09 = 1;
    92: op1_05_inv09 = 1;
    94: op1_05_inv09 = 1;
    97: op1_05_inv09 = 1;
    default: op1_05_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in10 = reg_0191;
    6: op1_05_in10 = imem07_in[71:68];
    7: op1_05_in10 = reg_0083;
    8: op1_05_in10 = reg_0136;
    9: op1_05_in10 = reg_0466;
    10: op1_05_in10 = reg_0392;
    11: op1_05_in10 = reg_0480;
    12: op1_05_in10 = reg_0448;
    4: op1_05_in10 = reg_0162;
    13: op1_05_in10 = imem03_in[63:60];
    14: op1_05_in10 = reg_0217;
    15: op1_05_in10 = reg_0726;
    16: op1_05_in10 = reg_0649;
    17: op1_05_in10 = imem04_in[7:4];
    18: op1_05_in10 = reg_0470;
    19: op1_05_in10 = imem05_in[15:12];
    3: op1_05_in10 = reg_0167;
    20: op1_05_in10 = reg_0468;
    21: op1_05_in10 = reg_0546;
    22: op1_05_in10 = reg_0669;
    23: op1_05_in10 = reg_0672;
    24: op1_05_in10 = reg_0801;
    25: op1_05_in10 = reg_0364;
    26: op1_05_in10 = reg_0511;
    27: op1_05_in10 = reg_0659;
    28: op1_05_in10 = imem03_in[39:36];
    29: op1_05_in10 = reg_0678;
    30: op1_05_in10 = reg_0462;
    84: op1_05_in10 = reg_0462;
    31: op1_05_in10 = reg_0986;
    32: op1_05_in10 = reg_0804;
    33: op1_05_in10 = reg_0694;
    74: op1_05_in10 = reg_0694;
    34: op1_05_in10 = reg_0863;
    36: op1_05_in10 = reg_0295;
    37: op1_05_in10 = reg_0446;
    39: op1_05_in10 = reg_0671;
    40: op1_05_in10 = reg_0665;
    41: op1_05_in10 = reg_0469;
    42: op1_05_in10 = reg_0821;
    43: op1_05_in10 = imem07_in[119:116];
    44: op1_05_in10 = reg_0670;
    47: op1_05_in10 = reg_0670;
    45: op1_05_in10 = reg_0982;
    46: op1_05_in10 = reg_0497;
    48: op1_05_in10 = reg_0651;
    49: op1_05_in10 = imem06_in[127:124];
    50: op1_05_in10 = reg_0074;
    51: op1_05_in10 = reg_0246;
    52: op1_05_in10 = reg_0186;
    53: op1_05_in10 = reg_0052;
    54: op1_05_in10 = reg_1002;
    55: op1_05_in10 = imem05_in[51:48];
    56: op1_05_in10 = reg_0831;
    57: op1_05_in10 = reg_0243;
    59: op1_05_in10 = reg_0146;
    60: op1_05_in10 = reg_0102;
    61: op1_05_in10 = reg_0183;
    62: op1_05_in10 = reg_0477;
    63: op1_05_in10 = reg_0984;
    64: op1_05_in10 = reg_0276;
    65: op1_05_in10 = imem06_in[23:20];
    66: op1_05_in10 = imem06_in[71:68];
    67: op1_05_in10 = reg_0958;
    68: op1_05_in10 = reg_0263;
    69: op1_05_in10 = reg_0224;
    70: op1_05_in10 = reg_0850;
    71: op1_05_in10 = imem07_in[59:56];
    72: op1_05_in10 = imem04_in[119:116];
    73: op1_05_in10 = imem05_in[23:20];
    75: op1_05_in10 = imem07_in[115:112];
    76: op1_05_in10 = reg_0464;
    77: op1_05_in10 = reg_0452;
    78: op1_05_in10 = imem02_in[51:48];
    79: op1_05_in10 = reg_0334;
    80: op1_05_in10 = imem06_in[43:40];
    81: op1_05_in10 = reg_0160;
    82: op1_05_in10 = reg_0691;
    83: op1_05_in10 = reg_0347;
    85: op1_05_in10 = reg_0139;
    87: op1_05_in10 = imem03_in[75:72];
    88: op1_05_in10 = reg_0752;
    89: op1_05_in10 = reg_0189;
    90: op1_05_in10 = imem06_in[39:36];
    91: op1_05_in10 = imem06_in[123:120];
    92: op1_05_in10 = reg_0297;
    93: op1_05_in10 = reg_0461;
    94: op1_05_in10 = reg_0201;
    95: op1_05_in10 = reg_0463;
    96: op1_05_in10 = reg_0474;
    97: op1_05_in10 = reg_0805;
    default: op1_05_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv10 = 1;
    8: op1_05_inv10 = 1;
    10: op1_05_inv10 = 1;
    14: op1_05_inv10 = 1;
    18: op1_05_inv10 = 1;
    19: op1_05_inv10 = 1;
    21: op1_05_inv10 = 1;
    22: op1_05_inv10 = 1;
    23: op1_05_inv10 = 1;
    24: op1_05_inv10 = 1;
    25: op1_05_inv10 = 1;
    27: op1_05_inv10 = 1;
    30: op1_05_inv10 = 1;
    31: op1_05_inv10 = 1;
    36: op1_05_inv10 = 1;
    37: op1_05_inv10 = 1;
    40: op1_05_inv10 = 1;
    43: op1_05_inv10 = 1;
    46: op1_05_inv10 = 1;
    47: op1_05_inv10 = 1;
    49: op1_05_inv10 = 1;
    54: op1_05_inv10 = 1;
    55: op1_05_inv10 = 1;
    59: op1_05_inv10 = 1;
    60: op1_05_inv10 = 1;
    61: op1_05_inv10 = 1;
    62: op1_05_inv10 = 1;
    65: op1_05_inv10 = 1;
    66: op1_05_inv10 = 1;
    68: op1_05_inv10 = 1;
    69: op1_05_inv10 = 1;
    70: op1_05_inv10 = 1;
    71: op1_05_inv10 = 1;
    74: op1_05_inv10 = 1;
    77: op1_05_inv10 = 1;
    84: op1_05_inv10 = 1;
    87: op1_05_inv10 = 1;
    88: op1_05_inv10 = 1;
    89: op1_05_inv10 = 1;
    92: op1_05_inv10 = 1;
    93: op1_05_inv10 = 1;
    94: op1_05_inv10 = 1;
    95: op1_05_inv10 = 1;
    96: op1_05_inv10 = 1;
    default: op1_05_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in11 = reg_0209;
    6: op1_05_in11 = reg_0722;
    7: op1_05_in11 = reg_0042;
    8: op1_05_in11 = reg_0151;
    9: op1_05_in11 = reg_0471;
    10: op1_05_in11 = reg_0351;
    11: op1_05_in11 = reg_0473;
    12: op1_05_in11 = reg_0174;
    4: op1_05_in11 = reg_0167;
    13: op1_05_in11 = imem03_in[95:92];
    14: op1_05_in11 = reg_0897;
    15: op1_05_in11 = reg_0425;
    16: op1_05_in11 = reg_0644;
    17: op1_05_in11 = imem04_in[39:36];
    18: op1_05_in11 = reg_0479;
    19: op1_05_in11 = imem05_in[47:44];
    73: op1_05_in11 = imem05_in[47:44];
    3: op1_05_in11 = reg_0182;
    20: op1_05_in11 = reg_0478;
    21: op1_05_in11 = reg_0558;
    48: op1_05_in11 = reg_0558;
    22: op1_05_in11 = reg_0477;
    23: op1_05_in11 = reg_0699;
    24: op1_05_in11 = reg_0018;
    25: op1_05_in11 = reg_0359;
    26: op1_05_in11 = reg_0265;
    27: op1_05_in11 = reg_0334;
    28: op1_05_in11 = imem03_in[47:44];
    29: op1_05_in11 = reg_0673;
    30: op1_05_in11 = reg_0474;
    31: op1_05_in11 = reg_0974;
    32: op1_05_in11 = reg_0349;
    33: op1_05_in11 = reg_0676;
    79: op1_05_in11 = reg_0676;
    34: op1_05_in11 = reg_0318;
    36: op1_05_in11 = reg_0402;
    37: op1_05_in11 = reg_0440;
    39: op1_05_in11 = reg_0675;
    40: op1_05_in11 = reg_0097;
    41: op1_05_in11 = reg_0476;
    42: op1_05_in11 = reg_0835;
    44: op1_05_in11 = reg_0679;
    45: op1_05_in11 = reg_0991;
    46: op1_05_in11 = reg_0155;
    47: op1_05_in11 = reg_0668;
    49: op1_05_in11 = reg_0220;
    50: op1_05_in11 = reg_0072;
    51: op1_05_in11 = reg_0234;
    52: op1_05_in11 = reg_0194;
    53: op1_05_in11 = reg_0608;
    54: op1_05_in11 = reg_0990;
    55: op1_05_in11 = imem05_in[79:76];
    56: op1_05_in11 = imem05_in[31:28];
    57: op1_05_in11 = reg_0399;
    59: op1_05_in11 = reg_0129;
    60: op1_05_in11 = reg_0828;
    61: op1_05_in11 = reg_0168;
    62: op1_05_in11 = reg_0469;
    63: op1_05_in11 = reg_0996;
    64: op1_05_in11 = reg_0815;
    65: op1_05_in11 = imem06_in[55:52];
    66: op1_05_in11 = imem06_in[75:72];
    67: op1_05_in11 = reg_0782;
    68: op1_05_in11 = imem07_in[31:28];
    69: op1_05_in11 = reg_0279;
    70: op1_05_in11 = reg_0732;
    71: op1_05_in11 = imem07_in[107:104];
    72: op1_05_in11 = imem04_in[127:124];
    74: op1_05_in11 = reg_1019;
    75: op1_05_in11 = reg_0361;
    76: op1_05_in11 = reg_0460;
    77: op1_05_in11 = reg_0200;
    78: op1_05_in11 = imem02_in[59:56];
    80: op1_05_in11 = imem06_in[71:68];
    81: op1_05_in11 = reg_0127;
    82: op1_05_in11 = reg_0267;
    83: op1_05_in11 = reg_0776;
    84: op1_05_in11 = reg_0480;
    85: op1_05_in11 = reg_0138;
    87: op1_05_in11 = imem03_in[83:80];
    88: op1_05_in11 = reg_0568;
    89: op1_05_in11 = reg_0206;
    90: op1_05_in11 = imem06_in[63:60];
    91: op1_05_in11 = reg_0691;
    92: op1_05_in11 = reg_0533;
    93: op1_05_in11 = reg_0475;
    94: op1_05_in11 = reg_0195;
    95: op1_05_in11 = reg_0466;
    96: op1_05_in11 = reg_0468;
    97: op1_05_in11 = reg_0325;
    default: op1_05_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv11 = 1;
    7: op1_05_inv11 = 1;
    8: op1_05_inv11 = 1;
    9: op1_05_inv11 = 1;
    11: op1_05_inv11 = 1;
    12: op1_05_inv11 = 1;
    4: op1_05_inv11 = 1;
    13: op1_05_inv11 = 1;
    15: op1_05_inv11 = 1;
    17: op1_05_inv11 = 1;
    19: op1_05_inv11 = 1;
    3: op1_05_inv11 = 1;
    22: op1_05_inv11 = 1;
    24: op1_05_inv11 = 1;
    27: op1_05_inv11 = 1;
    28: op1_05_inv11 = 1;
    30: op1_05_inv11 = 1;
    31: op1_05_inv11 = 1;
    33: op1_05_inv11 = 1;
    39: op1_05_inv11 = 1;
    40: op1_05_inv11 = 1;
    41: op1_05_inv11 = 1;
    42: op1_05_inv11 = 1;
    47: op1_05_inv11 = 1;
    49: op1_05_inv11 = 1;
    51: op1_05_inv11 = 1;
    52: op1_05_inv11 = 1;
    53: op1_05_inv11 = 1;
    56: op1_05_inv11 = 1;
    57: op1_05_inv11 = 1;
    60: op1_05_inv11 = 1;
    61: op1_05_inv11 = 1;
    63: op1_05_inv11 = 1;
    66: op1_05_inv11 = 1;
    69: op1_05_inv11 = 1;
    73: op1_05_inv11 = 1;
    74: op1_05_inv11 = 1;
    80: op1_05_inv11 = 1;
    81: op1_05_inv11 = 1;
    84: op1_05_inv11 = 1;
    85: op1_05_inv11 = 1;
    87: op1_05_inv11 = 1;
    90: op1_05_inv11 = 1;
    91: op1_05_inv11 = 1;
    default: op1_05_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in12 = reg_0203;
    77: op1_05_in12 = reg_0203;
    96: op1_05_in12 = reg_0203;
    6: op1_05_in12 = reg_0726;
    7: op1_05_in12 = reg_0095;
    8: op1_05_in12 = reg_0142;
    9: op1_05_in12 = reg_0468;
    39: op1_05_in12 = reg_0468;
    10: op1_05_in12 = reg_0409;
    11: op1_05_in12 = reg_0467;
    12: op1_05_in12 = reg_0165;
    4: op1_05_in12 = reg_0177;
    13: op1_05_in12 = reg_0582;
    14: op1_05_in12 = reg_0254;
    15: op1_05_in12 = reg_0430;
    16: op1_05_in12 = reg_0358;
    17: op1_05_in12 = imem04_in[43:40];
    18: op1_05_in12 = reg_0478;
    19: op1_05_in12 = imem05_in[59:56];
    3: op1_05_in12 = reg_0160;
    20: op1_05_in12 = imem01_in[19:16];
    21: op1_05_in12 = reg_0551;
    22: op1_05_in12 = reg_0462;
    23: op1_05_in12 = reg_0461;
    24: op1_05_in12 = imem07_in[47:44];
    25: op1_05_in12 = reg_0345;
    26: op1_05_in12 = reg_0937;
    27: op1_05_in12 = reg_0225;
    28: op1_05_in12 = imem03_in[59:56];
    29: op1_05_in12 = reg_0463;
    30: op1_05_in12 = reg_0194;
    31: op1_05_in12 = reg_0976;
    32: op1_05_in12 = reg_0222;
    33: op1_05_in12 = reg_0670;
    34: op1_05_in12 = reg_0886;
    36: op1_05_in12 = reg_0011;
    37: op1_05_in12 = reg_0437;
    40: op1_05_in12 = reg_0330;
    41: op1_05_in12 = reg_0480;
    42: op1_05_in12 = reg_0900;
    44: op1_05_in12 = reg_0690;
    45: op1_05_in12 = reg_0984;
    46: op1_05_in12 = imem06_in[31:28];
    47: op1_05_in12 = reg_0477;
    48: op1_05_in12 = reg_0418;
    49: op1_05_in12 = reg_0533;
    50: op1_05_in12 = reg_0517;
    51: op1_05_in12 = reg_1001;
    52: op1_05_in12 = reg_0195;
    53: op1_05_in12 = reg_0335;
    54: op1_05_in12 = imem04_in[7:4];
    55: op1_05_in12 = imem05_in[87:84];
    56: op1_05_in12 = imem05_in[35:32];
    57: op1_05_in12 = reg_0332;
    59: op1_05_in12 = reg_0131;
    60: op1_05_in12 = reg_0687;
    61: op1_05_in12 = reg_0171;
    62: op1_05_in12 = reg_0466;
    63: op1_05_in12 = reg_0986;
    64: op1_05_in12 = reg_0072;
    65: op1_05_in12 = imem06_in[115:112];
    66: op1_05_in12 = imem06_in[119:116];
    67: op1_05_in12 = reg_0941;
    68: op1_05_in12 = imem07_in[39:36];
    69: op1_05_in12 = reg_0329;
    70: op1_05_in12 = reg_0432;
    71: op1_05_in12 = reg_0704;
    72: op1_05_in12 = reg_0530;
    73: op1_05_in12 = imem05_in[55:52];
    74: op1_05_in12 = reg_0617;
    75: op1_05_in12 = reg_0315;
    76: op1_05_in12 = reg_0187;
    78: op1_05_in12 = imem02_in[75:72];
    79: op1_05_in12 = reg_0094;
    80: op1_05_in12 = imem06_in[75:72];
    81: op1_05_in12 = reg_0031;
    82: op1_05_in12 = reg_0025;
    83: op1_05_in12 = reg_0876;
    84: op1_05_in12 = reg_0474;
    85: op1_05_in12 = reg_0141;
    87: op1_05_in12 = imem03_in[107:104];
    88: op1_05_in12 = reg_0288;
    89: op1_05_in12 = imem01_in[71:68];
    90: op1_05_in12 = imem06_in[67:64];
    91: op1_05_in12 = reg_0391;
    92: op1_05_in12 = reg_0380;
    93: op1_05_in12 = reg_0459;
    94: op1_05_in12 = reg_0199;
    95: op1_05_in12 = reg_0475;
    97: op1_05_in12 = reg_0422;
    default: op1_05_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv12 = 1;
    8: op1_05_inv12 = 1;
    9: op1_05_inv12 = 1;
    11: op1_05_inv12 = 1;
    15: op1_05_inv12 = 1;
    17: op1_05_inv12 = 1;
    18: op1_05_inv12 = 1;
    19: op1_05_inv12 = 1;
    3: op1_05_inv12 = 1;
    20: op1_05_inv12 = 1;
    21: op1_05_inv12 = 1;
    24: op1_05_inv12 = 1;
    25: op1_05_inv12 = 1;
    26: op1_05_inv12 = 1;
    28: op1_05_inv12 = 1;
    30: op1_05_inv12 = 1;
    31: op1_05_inv12 = 1;
    33: op1_05_inv12 = 1;
    40: op1_05_inv12 = 1;
    41: op1_05_inv12 = 1;
    44: op1_05_inv12 = 1;
    46: op1_05_inv12 = 1;
    48: op1_05_inv12 = 1;
    49: op1_05_inv12 = 1;
    51: op1_05_inv12 = 1;
    53: op1_05_inv12 = 1;
    54: op1_05_inv12 = 1;
    57: op1_05_inv12 = 1;
    61: op1_05_inv12 = 1;
    63: op1_05_inv12 = 1;
    64: op1_05_inv12 = 1;
    65: op1_05_inv12 = 1;
    66: op1_05_inv12 = 1;
    68: op1_05_inv12 = 1;
    69: op1_05_inv12 = 1;
    73: op1_05_inv12 = 1;
    75: op1_05_inv12 = 1;
    80: op1_05_inv12 = 1;
    83: op1_05_inv12 = 1;
    85: op1_05_inv12 = 1;
    89: op1_05_inv12 = 1;
    92: op1_05_inv12 = 1;
    93: op1_05_inv12 = 1;
    96: op1_05_inv12 = 1;
    default: op1_05_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in13 = reg_0190;
    6: op1_05_in13 = reg_0711;
    7: op1_05_in13 = reg_0096;
    48: op1_05_in13 = reg_0096;
    8: op1_05_in13 = reg_0146;
    9: op1_05_in13 = reg_0479;
    11: op1_05_in13 = reg_0479;
    10: op1_05_in13 = reg_0371;
    4: op1_05_in13 = reg_0157;
    13: op1_05_in13 = reg_0572;
    14: op1_05_in13 = reg_0832;
    15: op1_05_in13 = reg_0447;
    79: op1_05_in13 = reg_0447;
    16: op1_05_in13 = reg_0320;
    17: op1_05_in13 = imem04_in[119:116];
    18: op1_05_in13 = reg_0212;
    30: op1_05_in13 = reg_0212;
    19: op1_05_in13 = imem05_in[71:68];
    3: op1_05_in13 = reg_0176;
    20: op1_05_in13 = imem01_in[23:20];
    21: op1_05_in13 = reg_0559;
    22: op1_05_in13 = reg_0472;
    23: op1_05_in13 = reg_0476;
    24: op1_05_in13 = imem07_in[55:52];
    25: op1_05_in13 = reg_0353;
    26: op1_05_in13 = reg_1009;
    27: op1_05_in13 = reg_0318;
    28: op1_05_in13 = imem03_in[63:60];
    29: op1_05_in13 = reg_0454;
    31: op1_05_in13 = imem04_in[7:4];
    32: op1_05_in13 = reg_0380;
    33: op1_05_in13 = reg_0677;
    34: op1_05_in13 = reg_0338;
    36: op1_05_in13 = reg_0367;
    37: op1_05_in13 = reg_0173;
    39: op1_05_in13 = reg_0187;
    40: op1_05_in13 = reg_0049;
    41: op1_05_in13 = reg_0468;
    42: op1_05_in13 = reg_0252;
    44: op1_05_in13 = reg_0455;
    45: op1_05_in13 = reg_0986;
    51: op1_05_in13 = reg_0986;
    46: op1_05_in13 = imem06_in[87:84];
    47: op1_05_in13 = reg_0469;
    49: op1_05_in13 = reg_0392;
    50: op1_05_in13 = reg_0429;
    52: op1_05_in13 = reg_0199;
    53: op1_05_in13 = reg_0758;
    54: op1_05_in13 = imem04_in[51:48];
    55: op1_05_in13 = reg_0973;
    56: op1_05_in13 = imem05_in[51:48];
    57: op1_05_in13 = reg_0596;
    59: op1_05_in13 = reg_0144;
    60: op1_05_in13 = reg_0749;
    62: op1_05_in13 = reg_0480;
    63: op1_05_in13 = imem04_in[23:20];
    64: op1_05_in13 = reg_0809;
    65: op1_05_in13 = imem06_in[127:124];
    66: op1_05_in13 = reg_0691;
    67: op1_05_in13 = reg_0940;
    68: op1_05_in13 = imem07_in[51:48];
    69: op1_05_in13 = reg_0423;
    70: op1_05_in13 = reg_0552;
    71: op1_05_in13 = reg_0719;
    72: op1_05_in13 = reg_1003;
    73: op1_05_in13 = reg_0004;
    74: op1_05_in13 = reg_0595;
    75: op1_05_in13 = reg_0024;
    76: op1_05_in13 = reg_0193;
    77: op1_05_in13 = reg_0201;
    78: op1_05_in13 = imem02_in[95:92];
    80: op1_05_in13 = reg_0660;
    81: op1_05_in13 = reg_0515;
    82: op1_05_in13 = reg_0626;
    91: op1_05_in13 = reg_0626;
    83: op1_05_in13 = reg_0872;
    84: op1_05_in13 = reg_0478;
    85: op1_05_in13 = reg_0448;
    87: op1_05_in13 = imem03_in[119:116];
    88: op1_05_in13 = reg_0284;
    89: op1_05_in13 = imem01_in[123:120];
    90: op1_05_in13 = imem06_in[75:72];
    92: op1_05_in13 = reg_0811;
    93: op1_05_in13 = reg_0452;
    94: op1_05_in13 = reg_0270;
    95: op1_05_in13 = reg_0462;
    96: op1_05_in13 = reg_0211;
    97: op1_05_in13 = reg_0641;
    default: op1_05_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv13 = 1;
    7: op1_05_inv13 = 1;
    8: op1_05_inv13 = 1;
    9: op1_05_inv13 = 1;
    11: op1_05_inv13 = 1;
    13: op1_05_inv13 = 1;
    14: op1_05_inv13 = 1;
    15: op1_05_inv13 = 1;
    17: op1_05_inv13 = 1;
    19: op1_05_inv13 = 1;
    23: op1_05_inv13 = 1;
    26: op1_05_inv13 = 1;
    27: op1_05_inv13 = 1;
    36: op1_05_inv13 = 1;
    41: op1_05_inv13 = 1;
    42: op1_05_inv13 = 1;
    44: op1_05_inv13 = 1;
    47: op1_05_inv13 = 1;
    53: op1_05_inv13 = 1;
    54: op1_05_inv13 = 1;
    56: op1_05_inv13 = 1;
    59: op1_05_inv13 = 1;
    60: op1_05_inv13 = 1;
    62: op1_05_inv13 = 1;
    63: op1_05_inv13 = 1;
    65: op1_05_inv13 = 1;
    69: op1_05_inv13 = 1;
    72: op1_05_inv13 = 1;
    78: op1_05_inv13 = 1;
    79: op1_05_inv13 = 1;
    80: op1_05_inv13 = 1;
    82: op1_05_inv13 = 1;
    85: op1_05_inv13 = 1;
    87: op1_05_inv13 = 1;
    88: op1_05_inv13 = 1;
    94: op1_05_inv13 = 1;
    95: op1_05_inv13 = 1;
    default: op1_05_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in14 = reg_0202;
    6: op1_05_in14 = reg_0727;
    7: op1_05_in14 = reg_0086;
    8: op1_05_in14 = reg_0139;
    9: op1_05_in14 = reg_0187;
    10: op1_05_in14 = reg_0375;
    11: op1_05_in14 = reg_0208;
    4: op1_05_in14 = reg_0173;
    13: op1_05_in14 = reg_0588;
    14: op1_05_in14 = reg_0149;
    15: op1_05_in14 = reg_0419;
    16: op1_05_in14 = reg_0341;
    17: op1_05_in14 = reg_0552;
    18: op1_05_in14 = reg_0205;
    19: op1_05_in14 = imem05_in[119:116];
    20: op1_05_in14 = imem01_in[39:36];
    21: op1_05_in14 = reg_0547;
    22: op1_05_in14 = reg_0473;
    23: op1_05_in14 = reg_0475;
    24: op1_05_in14 = imem07_in[59:56];
    25: op1_05_in14 = reg_0350;
    97: op1_05_in14 = reg_0350;
    26: op1_05_in14 = reg_0912;
    27: op1_05_in14 = reg_0886;
    28: op1_05_in14 = imem03_in[71:68];
    29: op1_05_in14 = reg_0481;
    30: op1_05_in14 = reg_0197;
    31: op1_05_in14 = imem04_in[11:8];
    32: op1_05_in14 = reg_0917;
    33: op1_05_in14 = reg_0678;
    34: op1_05_in14 = reg_0037;
    36: op1_05_in14 = imem07_in[43:40];
    39: op1_05_in14 = reg_0204;
    40: op1_05_in14 = reg_0077;
    41: op1_05_in14 = reg_0478;
    42: op1_05_in14 = reg_0816;
    44: op1_05_in14 = reg_0472;
    95: op1_05_in14 = reg_0472;
    45: op1_05_in14 = imem04_in[31:28];
    46: op1_05_in14 = reg_0534;
    47: op1_05_in14 = reg_0462;
    48: op1_05_in14 = reg_0290;
    49: op1_05_in14 = reg_0351;
    50: op1_05_in14 = reg_0075;
    51: op1_05_in14 = reg_0980;
    52: op1_05_in14 = reg_0192;
    53: op1_05_in14 = reg_0090;
    54: op1_05_in14 = imem04_in[59:56];
    55: op1_05_in14 = reg_0966;
    56: op1_05_in14 = imem05_in[63:60];
    57: op1_05_in14 = reg_0545;
    59: op1_05_in14 = imem06_in[51:48];
    60: op1_05_in14 = reg_0453;
    62: op1_05_in14 = reg_0474;
    63: op1_05_in14 = imem04_in[51:48];
    64: op1_05_in14 = reg_0432;
    65: op1_05_in14 = reg_0817;
    66: op1_05_in14 = reg_0244;
    67: op1_05_in14 = reg_0259;
    68: op1_05_in14 = imem07_in[95:92];
    69: op1_05_in14 = reg_0331;
    70: op1_05_in14 = reg_0070;
    71: op1_05_in14 = reg_0717;
    72: op1_05_in14 = reg_0937;
    73: op1_05_in14 = reg_0786;
    74: op1_05_in14 = reg_0781;
    75: op1_05_in14 = reg_0431;
    76: op1_05_in14 = reg_0186;
    77: op1_05_in14 = imem01_in[19:16];
    78: op1_05_in14 = imem02_in[107:104];
    79: op1_05_in14 = reg_0263;
    80: op1_05_in14 = reg_0010;
    81: op1_05_in14 = reg_0442;
    82: op1_05_in14 = reg_0328;
    83: op1_05_in14 = imem03_in[43:40];
    84: op1_05_in14 = reg_0210;
    85: op1_05_in14 = reg_0137;
    87: op1_05_in14 = imem03_in[123:120];
    88: op1_05_in14 = reg_0065;
    89: op1_05_in14 = reg_0106;
    90: op1_05_in14 = imem06_in[83:80];
    91: op1_05_in14 = reg_0021;
    92: op1_05_in14 = reg_0918;
    93: op1_05_in14 = reg_0456;
    94: op1_05_in14 = reg_0236;
    96: op1_05_in14 = reg_0201;
    default: op1_05_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv14 = 1;
    7: op1_05_inv14 = 1;
    9: op1_05_inv14 = 1;
    10: op1_05_inv14 = 1;
    11: op1_05_inv14 = 1;
    17: op1_05_inv14 = 1;
    22: op1_05_inv14 = 1;
    24: op1_05_inv14 = 1;
    25: op1_05_inv14 = 1;
    26: op1_05_inv14 = 1;
    27: op1_05_inv14 = 1;
    29: op1_05_inv14 = 1;
    32: op1_05_inv14 = 1;
    33: op1_05_inv14 = 1;
    36: op1_05_inv14 = 1;
    39: op1_05_inv14 = 1;
    40: op1_05_inv14 = 1;
    41: op1_05_inv14 = 1;
    45: op1_05_inv14 = 1;
    46: op1_05_inv14 = 1;
    47: op1_05_inv14 = 1;
    48: op1_05_inv14 = 1;
    49: op1_05_inv14 = 1;
    54: op1_05_inv14 = 1;
    59: op1_05_inv14 = 1;
    62: op1_05_inv14 = 1;
    63: op1_05_inv14 = 1;
    65: op1_05_inv14 = 1;
    66: op1_05_inv14 = 1;
    67: op1_05_inv14 = 1;
    69: op1_05_inv14 = 1;
    70: op1_05_inv14 = 1;
    71: op1_05_inv14 = 1;
    73: op1_05_inv14 = 1;
    78: op1_05_inv14 = 1;
    79: op1_05_inv14 = 1;
    80: op1_05_inv14 = 1;
    81: op1_05_inv14 = 1;
    83: op1_05_inv14 = 1;
    88: op1_05_inv14 = 1;
    90: op1_05_inv14 = 1;
    92: op1_05_inv14 = 1;
    95: op1_05_inv14 = 1;
    96: op1_05_inv14 = 1;
    97: op1_05_inv14 = 1;
    default: op1_05_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in15 = imem01_in[19:16];
    6: op1_05_in15 = reg_0424;
    7: op1_05_in15 = imem03_in[31:28];
    8: op1_05_in15 = reg_0141;
    9: op1_05_in15 = reg_0188;
    10: op1_05_in15 = reg_0382;
    11: op1_05_in15 = reg_0191;
    13: op1_05_in15 = reg_0384;
    82: op1_05_in15 = reg_0384;
    91: op1_05_in15 = reg_0384;
    14: op1_05_in15 = reg_0128;
    15: op1_05_in15 = reg_0442;
    16: op1_05_in15 = reg_0359;
    17: op1_05_in15 = reg_0542;
    18: op1_05_in15 = reg_0190;
    19: op1_05_in15 = imem05_in[123:120];
    20: op1_05_in15 = reg_0235;
    21: op1_05_in15 = reg_0047;
    22: op1_05_in15 = reg_0470;
    23: op1_05_in15 = reg_0474;
    24: op1_05_in15 = imem07_in[67:64];
    25: op1_05_in15 = reg_0347;
    26: op1_05_in15 = reg_1057;
    27: op1_05_in15 = reg_0093;
    28: op1_05_in15 = imem03_in[75:72];
    29: op1_05_in15 = reg_0471;
    62: op1_05_in15 = reg_0471;
    30: op1_05_in15 = imem01_in[3:0];
    31: op1_05_in15 = imem04_in[83:80];
    32: op1_05_in15 = imem06_in[11:8];
    33: op1_05_in15 = reg_0675;
    34: op1_05_in15 = reg_0335;
    36: op1_05_in15 = imem07_in[47:44];
    39: op1_05_in15 = reg_0211;
    40: op1_05_in15 = imem03_in[35:32];
    41: op1_05_in15 = reg_0204;
    42: op1_05_in15 = reg_0257;
    44: op1_05_in15 = reg_0452;
    45: op1_05_in15 = imem04_in[55:52];
    46: op1_05_in15 = reg_0073;
    47: op1_05_in15 = reg_0481;
    48: op1_05_in15 = reg_0865;
    49: op1_05_in15 = reg_0390;
    50: op1_05_in15 = reg_0739;
    51: op1_05_in15 = reg_0997;
    52: op1_05_in15 = imem01_in[39:36];
    53: op1_05_in15 = reg_0506;
    54: op1_05_in15 = imem04_in[75:72];
    55: op1_05_in15 = reg_0964;
    56: op1_05_in15 = imem05_in[75:72];
    57: op1_05_in15 = reg_0263;
    59: op1_05_in15 = reg_0660;
    60: op1_05_in15 = reg_0469;
    63: op1_05_in15 = imem04_in[67:64];
    64: op1_05_in15 = reg_0658;
    65: op1_05_in15 = reg_0328;
    66: op1_05_in15 = reg_0351;
    67: op1_05_in15 = reg_0935;
    68: op1_05_in15 = imem07_in[115:112];
    69: op1_05_in15 = reg_0644;
    70: op1_05_in15 = imem05_in[35:32];
    71: op1_05_in15 = reg_0713;
    72: op1_05_in15 = reg_0888;
    73: op1_05_in15 = reg_0149;
    74: op1_05_in15 = reg_0556;
    75: op1_05_in15 = reg_0175;
    76: op1_05_in15 = reg_0205;
    77: op1_05_in15 = imem01_in[23:20];
    78: op1_05_in15 = imem02_in[111:108];
    79: op1_05_in15 = reg_0647;
    80: op1_05_in15 = reg_0344;
    81: op1_05_in15 = reg_0563;
    83: op1_05_in15 = imem03_in[71:68];
    84: op1_05_in15 = reg_0209;
    93: op1_05_in15 = reg_0209;
    85: op1_05_in15 = reg_0963;
    87: op1_05_in15 = reg_0535;
    88: op1_05_in15 = reg_0071;
    89: op1_05_in15 = reg_0488;
    90: op1_05_in15 = imem06_in[95:92];
    92: op1_05_in15 = reg_0914;
    94: op1_05_in15 = reg_0368;
    95: op1_05_in15 = reg_0459;
    96: op1_05_in15 = reg_0206;
    97: op1_05_in15 = reg_0420;
    default: op1_05_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv15 = 1;
    10: op1_05_inv15 = 1;
    14: op1_05_inv15 = 1;
    18: op1_05_inv15 = 1;
    21: op1_05_inv15 = 1;
    23: op1_05_inv15 = 1;
    24: op1_05_inv15 = 1;
    28: op1_05_inv15 = 1;
    29: op1_05_inv15 = 1;
    31: op1_05_inv15 = 1;
    33: op1_05_inv15 = 1;
    34: op1_05_inv15 = 1;
    42: op1_05_inv15 = 1;
    44: op1_05_inv15 = 1;
    46: op1_05_inv15 = 1;
    47: op1_05_inv15 = 1;
    48: op1_05_inv15 = 1;
    49: op1_05_inv15 = 1;
    51: op1_05_inv15 = 1;
    52: op1_05_inv15 = 1;
    53: op1_05_inv15 = 1;
    54: op1_05_inv15 = 1;
    55: op1_05_inv15 = 1;
    56: op1_05_inv15 = 1;
    57: op1_05_inv15 = 1;
    62: op1_05_inv15 = 1;
    63: op1_05_inv15 = 1;
    64: op1_05_inv15 = 1;
    66: op1_05_inv15 = 1;
    69: op1_05_inv15 = 1;
    70: op1_05_inv15 = 1;
    71: op1_05_inv15 = 1;
    73: op1_05_inv15 = 1;
    75: op1_05_inv15 = 1;
    76: op1_05_inv15 = 1;
    81: op1_05_inv15 = 1;
    82: op1_05_inv15 = 1;
    84: op1_05_inv15 = 1;
    85: op1_05_inv15 = 1;
    88: op1_05_inv15 = 1;
    90: op1_05_inv15 = 1;
    91: op1_05_inv15 = 1;
    93: op1_05_inv15 = 1;
    95: op1_05_inv15 = 1;
    96: op1_05_inv15 = 1;
    default: op1_05_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in16 = imem01_in[63:60];
    6: op1_05_in16 = reg_0419;
    7: op1_05_in16 = imem03_in[35:32];
    8: op1_05_in16 = reg_0137;
    9: op1_05_in16 = reg_0203;
    10: op1_05_in16 = reg_0406;
    11: op1_05_in16 = reg_0188;
    44: op1_05_in16 = reg_0188;
    13: op1_05_in16 = reg_0388;
    14: op1_05_in16 = reg_0154;
    15: op1_05_in16 = reg_0427;
    16: op1_05_in16 = reg_0318;
    17: op1_05_in16 = reg_0549;
    18: op1_05_in16 = reg_0197;
    19: op1_05_in16 = reg_0973;
    20: op1_05_in16 = reg_1055;
    21: op1_05_in16 = reg_0279;
    22: op1_05_in16 = reg_0452;
    23: op1_05_in16 = reg_0471;
    24: op1_05_in16 = imem07_in[87:84];
    25: op1_05_in16 = reg_0089;
    26: op1_05_in16 = reg_0078;
    27: op1_05_in16 = reg_0085;
    28: op1_05_in16 = imem03_in[83:80];
    29: op1_05_in16 = reg_0479;
    30: op1_05_in16 = imem01_in[15:12];
    31: op1_05_in16 = imem04_in[87:84];
    32: op1_05_in16 = imem06_in[23:20];
    33: op1_05_in16 = reg_0669;
    34: op1_05_in16 = reg_0772;
    36: op1_05_in16 = imem07_in[59:56];
    39: op1_05_in16 = reg_0198;
    40: op1_05_in16 = imem03_in[43:40];
    41: op1_05_in16 = reg_0503;
    42: op1_05_in16 = reg_0260;
    45: op1_05_in16 = imem04_in[63:60];
    46: op1_05_in16 = reg_0883;
    47: op1_05_in16 = reg_0472;
    48: op1_05_in16 = reg_0336;
    49: op1_05_in16 = reg_0222;
    50: op1_05_in16 = reg_0258;
    51: op1_05_in16 = reg_0994;
    52: op1_05_in16 = imem01_in[59:56];
    53: op1_05_in16 = imem03_in[51:48];
    54: op1_05_in16 = imem04_in[91:88];
    55: op1_05_in16 = reg_0965;
    56: op1_05_in16 = imem05_in[87:84];
    57: op1_05_in16 = imem07_in[15:12];
    59: op1_05_in16 = reg_0080;
    60: op1_05_in16 = reg_0470;
    62: op1_05_in16 = reg_0189;
    63: op1_05_in16 = imem04_in[99:96];
    64: op1_05_in16 = reg_0027;
    65: op1_05_in16 = reg_0229;
    66: op1_05_in16 = reg_0391;
    67: op1_05_in16 = reg_0020;
    68: op1_05_in16 = reg_0725;
    69: op1_05_in16 = reg_0037;
    70: op1_05_in16 = imem05_in[51:48];
    71: op1_05_in16 = reg_0715;
    72: op1_05_in16 = reg_0076;
    73: op1_05_in16 = reg_0155;
    74: op1_05_in16 = reg_0632;
    75: op1_05_in16 = reg_0161;
    76: op1_05_in16 = reg_0206;
    77: op1_05_in16 = imem01_in[27:24];
    78: op1_05_in16 = reg_0813;
    79: op1_05_in16 = reg_0139;
    80: op1_05_in16 = reg_0691;
    81: op1_05_in16 = reg_0653;
    82: op1_05_in16 = reg_1030;
    83: op1_05_in16 = imem03_in[91:88];
    84: op1_05_in16 = imem01_in[55:52];
    85: op1_05_in16 = reg_0150;
    87: op1_05_in16 = reg_0760;
    88: op1_05_in16 = reg_0777;
    89: op1_05_in16 = reg_1039;
    90: op1_05_in16 = imem06_in[107:104];
    91: op1_05_in16 = reg_0614;
    92: op1_05_in16 = reg_0034;
    93: op1_05_in16 = reg_0211;
    94: op1_05_in16 = reg_0304;
    95: op1_05_in16 = reg_0208;
    96: op1_05_in16 = reg_0270;
    97: op1_05_in16 = reg_0172;
    default: op1_05_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv16 = 1;
    10: op1_05_inv16 = 1;
    16: op1_05_inv16 = 1;
    17: op1_05_inv16 = 1;
    18: op1_05_inv16 = 1;
    20: op1_05_inv16 = 1;
    21: op1_05_inv16 = 1;
    22: op1_05_inv16 = 1;
    25: op1_05_inv16 = 1;
    27: op1_05_inv16 = 1;
    28: op1_05_inv16 = 1;
    30: op1_05_inv16 = 1;
    34: op1_05_inv16 = 1;
    40: op1_05_inv16 = 1;
    41: op1_05_inv16 = 1;
    44: op1_05_inv16 = 1;
    47: op1_05_inv16 = 1;
    49: op1_05_inv16 = 1;
    50: op1_05_inv16 = 1;
    52: op1_05_inv16 = 1;
    54: op1_05_inv16 = 1;
    55: op1_05_inv16 = 1;
    59: op1_05_inv16 = 1;
    64: op1_05_inv16 = 1;
    66: op1_05_inv16 = 1;
    71: op1_05_inv16 = 1;
    74: op1_05_inv16 = 1;
    77: op1_05_inv16 = 1;
    78: op1_05_inv16 = 1;
    79: op1_05_inv16 = 1;
    82: op1_05_inv16 = 1;
    84: op1_05_inv16 = 1;
    85: op1_05_inv16 = 1;
    89: op1_05_inv16 = 1;
    91: op1_05_inv16 = 1;
    93: op1_05_inv16 = 1;
    95: op1_05_inv16 = 1;
    96: op1_05_inv16 = 1;
    default: op1_05_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in17 = imem01_in[91:88];
    6: op1_05_in17 = reg_0439;
    7: op1_05_in17 = imem03_in[63:60];
    8: op1_05_in17 = imem06_in[19:16];
    9: op1_05_in17 = reg_0207;
    62: op1_05_in17 = reg_0207;
    10: op1_05_in17 = reg_0799;
    11: op1_05_in17 = reg_0203;
    13: op1_05_in17 = reg_0373;
    14: op1_05_in17 = reg_0153;
    15: op1_05_in17 = reg_0172;
    16: op1_05_in17 = reg_0092;
    17: op1_05_in17 = reg_0546;
    18: op1_05_in17 = imem01_in[67:64];
    19: op1_05_in17 = reg_0955;
    20: op1_05_in17 = reg_0239;
    21: op1_05_in17 = reg_0058;
    22: op1_05_in17 = reg_0458;
    23: op1_05_in17 = reg_0186;
    24: op1_05_in17 = imem07_in[95:92];
    25: op1_05_in17 = reg_0761;
    26: op1_05_in17 = reg_0760;
    27: op1_05_in17 = reg_0814;
    91: op1_05_in17 = reg_0814;
    28: op1_05_in17 = imem03_in[87:84];
    29: op1_05_in17 = reg_0478;
    30: op1_05_in17 = imem01_in[35:32];
    31: op1_05_in17 = imem04_in[107:104];
    32: op1_05_in17 = imem06_in[67:64];
    33: op1_05_in17 = reg_0461;
    34: op1_05_in17 = reg_0007;
    36: op1_05_in17 = imem07_in[127:124];
    39: op1_05_in17 = reg_0195;
    40: op1_05_in17 = imem03_in[103:100];
    41: op1_05_in17 = reg_0228;
    42: op1_05_in17 = reg_0832;
    44: op1_05_in17 = imem01_in[51:48];
    76: op1_05_in17 = imem01_in[51:48];
    45: op1_05_in17 = imem04_in[67:64];
    46: op1_05_in17 = reg_0895;
    65: op1_05_in17 = reg_0895;
    47: op1_05_in17 = reg_0208;
    48: op1_05_in17 = reg_0083;
    49: op1_05_in17 = reg_0384;
    50: op1_05_in17 = reg_0494;
    51: op1_05_in17 = imem04_in[3:0];
    52: op1_05_in17 = imem01_in[83:80];
    84: op1_05_in17 = imem01_in[83:80];
    53: op1_05_in17 = imem03_in[59:56];
    54: op1_05_in17 = imem04_in[95:92];
    55: op1_05_in17 = reg_0019;
    56: op1_05_in17 = imem05_in[103:100];
    57: op1_05_in17 = imem07_in[23:20];
    59: op1_05_in17 = reg_0351;
    60: op1_05_in17 = reg_0479;
    63: op1_05_in17 = imem04_in[115:112];
    64: op1_05_in17 = reg_0856;
    66: op1_05_in17 = reg_0262;
    67: op1_05_in17 = reg_0948;
    68: op1_05_in17 = reg_0729;
    69: op1_05_in17 = reg_0608;
    70: op1_05_in17 = imem05_in[91:88];
    71: op1_05_in17 = reg_0727;
    81: op1_05_in17 = reg_0727;
    72: op1_05_in17 = reg_0815;
    73: op1_05_in17 = imem06_in[39:36];
    74: op1_05_in17 = reg_0917;
    75: op1_05_in17 = reg_0167;
    77: op1_05_in17 = imem01_in[55:52];
    78: op1_05_in17 = reg_0637;
    79: op1_05_in17 = reg_0689;
    80: op1_05_in17 = reg_0391;
    82: op1_05_in17 = reg_0556;
    83: op1_05_in17 = reg_0535;
    85: op1_05_in17 = reg_0943;
    87: op1_05_in17 = reg_0572;
    88: op1_05_in17 = reg_0542;
    89: op1_05_in17 = reg_0869;
    90: op1_05_in17 = imem06_in[115:112];
    92: op1_05_in17 = reg_0628;
    93: op1_05_in17 = reg_0198;
    94: op1_05_in17 = imem01_in[7:4];
    95: op1_05_in17 = reg_0210;
    96: op1_05_in17 = reg_0519;
    97: op1_05_in17 = reg_0181;
    default: op1_05_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv17 = 1;
    8: op1_05_inv17 = 1;
    9: op1_05_inv17 = 1;
    14: op1_05_inv17 = 1;
    18: op1_05_inv17 = 1;
    19: op1_05_inv17 = 1;
    20: op1_05_inv17 = 1;
    21: op1_05_inv17 = 1;
    26: op1_05_inv17 = 1;
    29: op1_05_inv17 = 1;
    30: op1_05_inv17 = 1;
    31: op1_05_inv17 = 1;
    33: op1_05_inv17 = 1;
    36: op1_05_inv17 = 1;
    40: op1_05_inv17 = 1;
    44: op1_05_inv17 = 1;
    45: op1_05_inv17 = 1;
    49: op1_05_inv17 = 1;
    50: op1_05_inv17 = 1;
    51: op1_05_inv17 = 1;
    52: op1_05_inv17 = 1;
    54: op1_05_inv17 = 1;
    57: op1_05_inv17 = 1;
    60: op1_05_inv17 = 1;
    66: op1_05_inv17 = 1;
    67: op1_05_inv17 = 1;
    68: op1_05_inv17 = 1;
    69: op1_05_inv17 = 1;
    70: op1_05_inv17 = 1;
    71: op1_05_inv17 = 1;
    72: op1_05_inv17 = 1;
    73: op1_05_inv17 = 1;
    75: op1_05_inv17 = 1;
    76: op1_05_inv17 = 1;
    77: op1_05_inv17 = 1;
    78: op1_05_inv17 = 1;
    79: op1_05_inv17 = 1;
    80: op1_05_inv17 = 1;
    81: op1_05_inv17 = 1;
    82: op1_05_inv17 = 1;
    84: op1_05_inv17 = 1;
    88: op1_05_inv17 = 1;
    89: op1_05_inv17 = 1;
    90: op1_05_inv17 = 1;
    91: op1_05_inv17 = 1;
    93: op1_05_inv17 = 1;
    95: op1_05_inv17 = 1;
    97: op1_05_inv17 = 1;
    default: op1_05_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in18 = reg_0504;
    6: op1_05_in18 = reg_0440;
    7: op1_05_in18 = imem03_in[91:88];
    8: op1_05_in18 = imem06_in[23:20];
    9: op1_05_in18 = reg_0186;
    10: op1_05_in18 = reg_0808;
    11: op1_05_in18 = reg_0207;
    13: op1_05_in18 = reg_0398;
    14: op1_05_in18 = reg_0130;
    15: op1_05_in18 = reg_0167;
    16: op1_05_in18 = reg_0091;
    17: op1_05_in18 = reg_0308;
    18: op1_05_in18 = imem01_in[83:80];
    19: op1_05_in18 = reg_0954;
    20: op1_05_in18 = reg_0242;
    21: op1_05_in18 = reg_0057;
    22: op1_05_in18 = reg_0191;
    23: op1_05_in18 = reg_0199;
    39: op1_05_in18 = reg_0199;
    24: op1_05_in18 = reg_0728;
    25: op1_05_in18 = reg_0085;
    26: op1_05_in18 = reg_0063;
    27: op1_05_in18 = reg_0840;
    28: op1_05_in18 = imem03_in[99:96];
    53: op1_05_in18 = imem03_in[99:96];
    29: op1_05_in18 = reg_0200;
    60: op1_05_in18 = reg_0200;
    30: op1_05_in18 = imem01_in[63:60];
    31: op1_05_in18 = imem04_in[111:108];
    32: op1_05_in18 = imem06_in[71:68];
    33: op1_05_in18 = reg_0462;
    34: op1_05_in18 = reg_0089;
    36: op1_05_in18 = reg_0704;
    40: op1_05_in18 = reg_0535;
    41: op1_05_in18 = reg_1018;
    42: op1_05_in18 = reg_0137;
    44: op1_05_in18 = imem01_in[111:108];
    45: op1_05_in18 = imem04_in[79:76];
    46: op1_05_in18 = reg_0220;
    47: op1_05_in18 = reg_0190;
    62: op1_05_in18 = reg_0190;
    48: op1_05_in18 = imem03_in[31:28];
    49: op1_05_in18 = reg_0609;
    50: op1_05_in18 = reg_0828;
    51: op1_05_in18 = imem04_in[11:8];
    52: op1_05_in18 = reg_0936;
    54: op1_05_in18 = imem04_in[107:104];
    55: op1_05_in18 = reg_0032;
    74: op1_05_in18 = reg_0032;
    56: op1_05_in18 = imem05_in[119:116];
    57: op1_05_in18 = imem07_in[39:36];
    59: op1_05_in18 = reg_0626;
    66: op1_05_in18 = reg_0626;
    63: op1_05_in18 = reg_0530;
    64: op1_05_in18 = reg_0044;
    65: op1_05_in18 = reg_0392;
    67: op1_05_in18 = reg_0132;
    68: op1_05_in18 = reg_0713;
    69: op1_05_in18 = reg_0347;
    70: op1_05_in18 = imem05_in[115:112];
    71: op1_05_in18 = reg_0361;
    72: op1_05_in18 = reg_0064;
    73: op1_05_in18 = imem06_in[47:44];
    75: op1_05_in18 = reg_0163;
    76: op1_05_in18 = imem01_in[67:64];
    77: op1_05_in18 = imem01_in[67:64];
    78: op1_05_in18 = reg_0649;
    79: op1_05_in18 = reg_0269;
    80: op1_05_in18 = reg_0267;
    81: op1_05_in18 = reg_0321;
    82: op1_05_in18 = reg_0591;
    83: op1_05_in18 = reg_0661;
    84: op1_05_in18 = imem01_in[91:88];
    85: op1_05_in18 = reg_0486;
    87: op1_05_in18 = reg_0445;
    88: op1_05_in18 = reg_0332;
    89: op1_05_in18 = reg_0520;
    90: op1_05_in18 = reg_0025;
    91: op1_05_in18 = reg_0439;
    92: op1_05_in18 = reg_0611;
    93: op1_05_in18 = reg_0196;
    94: op1_05_in18 = imem01_in[47:44];
    95: op1_05_in18 = reg_0541;
    96: op1_05_in18 = reg_0245;
    97: op1_05_in18 = reg_0447;
    default: op1_05_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv18 = 1;
    6: op1_05_inv18 = 1;
    7: op1_05_inv18 = 1;
    9: op1_05_inv18 = 1;
    10: op1_05_inv18 = 1;
    11: op1_05_inv18 = 1;
    13: op1_05_inv18 = 1;
    14: op1_05_inv18 = 1;
    15: op1_05_inv18 = 1;
    16: op1_05_inv18 = 1;
    18: op1_05_inv18 = 1;
    24: op1_05_inv18 = 1;
    25: op1_05_inv18 = 1;
    28: op1_05_inv18 = 1;
    29: op1_05_inv18 = 1;
    30: op1_05_inv18 = 1;
    31: op1_05_inv18 = 1;
    34: op1_05_inv18 = 1;
    39: op1_05_inv18 = 1;
    40: op1_05_inv18 = 1;
    44: op1_05_inv18 = 1;
    45: op1_05_inv18 = 1;
    46: op1_05_inv18 = 1;
    49: op1_05_inv18 = 1;
    50: op1_05_inv18 = 1;
    52: op1_05_inv18 = 1;
    54: op1_05_inv18 = 1;
    55: op1_05_inv18 = 1;
    56: op1_05_inv18 = 1;
    59: op1_05_inv18 = 1;
    60: op1_05_inv18 = 1;
    62: op1_05_inv18 = 1;
    64: op1_05_inv18 = 1;
    66: op1_05_inv18 = 1;
    68: op1_05_inv18 = 1;
    69: op1_05_inv18 = 1;
    72: op1_05_inv18 = 1;
    75: op1_05_inv18 = 1;
    76: op1_05_inv18 = 1;
    77: op1_05_inv18 = 1;
    78: op1_05_inv18 = 1;
    79: op1_05_inv18 = 1;
    80: op1_05_inv18 = 1;
    81: op1_05_inv18 = 1;
    84: op1_05_inv18 = 1;
    85: op1_05_inv18 = 1;
    90: op1_05_inv18 = 1;
    96: op1_05_inv18 = 1;
    default: op1_05_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in19 = reg_0515;
    6: op1_05_in19 = reg_0427;
    7: op1_05_in19 = imem03_in[115:112];
    8: op1_05_in19 = imem06_in[35:32];
    9: op1_05_in19 = reg_0192;
    39: op1_05_in19 = reg_0192;
    10: op1_05_in19 = reg_0801;
    11: op1_05_in19 = reg_0212;
    13: op1_05_in19 = reg_0982;
    28: op1_05_in19 = reg_0982;
    14: op1_05_in19 = reg_0131;
    15: op1_05_in19 = reg_0169;
    16: op1_05_in19 = reg_0084;
    17: op1_05_in19 = reg_0305;
    18: op1_05_in19 = imem01_in[127:124];
    19: op1_05_in19 = reg_0951;
    20: op1_05_in19 = reg_0766;
    21: op1_05_in19 = reg_0864;
    22: op1_05_in19 = reg_0210;
    23: op1_05_in19 = imem01_in[3:0];
    24: op1_05_in19 = reg_0704;
    25: op1_05_in19 = reg_0091;
    26: op1_05_in19 = reg_0882;
    27: op1_05_in19 = reg_0872;
    29: op1_05_in19 = reg_0189;
    30: op1_05_in19 = imem01_in[67:64];
    31: op1_05_in19 = reg_1004;
    32: op1_05_in19 = imem06_in[75:72];
    33: op1_05_in19 = reg_0472;
    34: op1_05_in19 = reg_0792;
    36: op1_05_in19 = reg_0723;
    40: op1_05_in19 = reg_1050;
    41: op1_05_in19 = reg_0013;
    42: op1_05_in19 = reg_0134;
    44: op1_05_in19 = reg_0235;
    45: op1_05_in19 = reg_0536;
    46: op1_05_in19 = reg_0782;
    47: op1_05_in19 = reg_0197;
    48: op1_05_in19 = imem03_in[35:32];
    49: op1_05_in19 = imem07_in[39:36];
    50: op1_05_in19 = reg_0750;
    51: op1_05_in19 = imem04_in[59:56];
    52: op1_05_in19 = reg_0242;
    53: op1_05_in19 = imem03_in[127:124];
    54: op1_05_in19 = imem04_in[115:112];
    55: op1_05_in19 = reg_0023;
    56: op1_05_in19 = reg_0448;
    57: op1_05_in19 = imem07_in[91:88];
    59: op1_05_in19 = reg_0754;
    60: op1_05_in19 = reg_0208;
    62: op1_05_in19 = reg_0206;
    63: op1_05_in19 = reg_1003;
    64: op1_05_in19 = imem05_in[27:24];
    65: op1_05_in19 = reg_0439;
    66: op1_05_in19 = reg_0021;
    67: op1_05_in19 = reg_0154;
    68: op1_05_in19 = reg_0361;
    69: op1_05_in19 = reg_0482;
    70: op1_05_in19 = imem05_in[127:124];
    71: op1_05_in19 = reg_0002;
    72: op1_05_in19 = reg_0764;
    73: op1_05_in19 = imem06_in[51:48];
    74: op1_05_in19 = reg_0834;
    75: op1_05_in19 = reg_0183;
    97: op1_05_in19 = reg_0183;
    76: op1_05_in19 = imem01_in[71:68];
    77: op1_05_in19 = imem01_in[91:88];
    78: op1_05_in19 = reg_0846;
    79: op1_05_in19 = imem05_in[15:12];
    80: op1_05_in19 = reg_0328;
    81: op1_05_in19 = reg_0419;
    82: op1_05_in19 = reg_0220;
    83: op1_05_in19 = reg_0662;
    84: op1_05_in19 = imem01_in[99:96];
    85: op1_05_in19 = reg_0651;
    87: op1_05_in19 = reg_0590;
    88: op1_05_in19 = imem05_in[43:40];
    89: op1_05_in19 = reg_0227;
    90: op1_05_in19 = reg_0679;
    91: op1_05_in19 = reg_0343;
    92: op1_05_in19 = reg_0632;
    93: op1_05_in19 = reg_0202;
    94: op1_05_in19 = imem01_in[51:48];
    95: op1_05_in19 = reg_0240;
    96: op1_05_in19 = reg_0368;
    default: op1_05_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv19 = 1;
    9: op1_05_inv19 = 1;
    11: op1_05_inv19 = 1;
    14: op1_05_inv19 = 1;
    15: op1_05_inv19 = 1;
    16: op1_05_inv19 = 1;
    17: op1_05_inv19 = 1;
    19: op1_05_inv19 = 1;
    22: op1_05_inv19 = 1;
    24: op1_05_inv19 = 1;
    31: op1_05_inv19 = 1;
    32: op1_05_inv19 = 1;
    34: op1_05_inv19 = 1;
    40: op1_05_inv19 = 1;
    48: op1_05_inv19 = 1;
    49: op1_05_inv19 = 1;
    51: op1_05_inv19 = 1;
    53: op1_05_inv19 = 1;
    54: op1_05_inv19 = 1;
    55: op1_05_inv19 = 1;
    56: op1_05_inv19 = 1;
    57: op1_05_inv19 = 1;
    64: op1_05_inv19 = 1;
    67: op1_05_inv19 = 1;
    69: op1_05_inv19 = 1;
    72: op1_05_inv19 = 1;
    76: op1_05_inv19 = 1;
    77: op1_05_inv19 = 1;
    79: op1_05_inv19 = 1;
    80: op1_05_inv19 = 1;
    82: op1_05_inv19 = 1;
    85: op1_05_inv19 = 1;
    89: op1_05_inv19 = 1;
    93: op1_05_inv19 = 1;
    94: op1_05_inv19 = 1;
    95: op1_05_inv19 = 1;
    97: op1_05_inv19 = 1;
    default: op1_05_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in20 = reg_0487;
    6: op1_05_in20 = reg_0167;
    7: op1_05_in20 = reg_0571;
    8: op1_05_in20 = imem06_in[63:60];
    9: op1_05_in20 = imem01_in[91:88];
    10: op1_05_in20 = reg_0017;
    82: op1_05_in20 = reg_0017;
    11: op1_05_in20 = reg_0222;
    13: op1_05_in20 = reg_0999;
    14: op1_05_in20 = imem06_in[39:36];
    15: op1_05_in20 = reg_0177;
    16: op1_05_in20 = reg_0098;
    17: op1_05_in20 = reg_0293;
    18: op1_05_in20 = reg_0235;
    19: op1_05_in20 = reg_0942;
    20: op1_05_in20 = reg_1056;
    21: op1_05_in20 = imem05_in[19:16];
    22: op1_05_in20 = reg_0187;
    23: op1_05_in20 = imem01_in[39:36];
    47: op1_05_in20 = imem01_in[39:36];
    24: op1_05_in20 = reg_0723;
    25: op1_05_in20 = reg_0016;
    26: op1_05_in20 = reg_0056;
    27: op1_05_in20 = imem03_in[23:20];
    28: op1_05_in20 = reg_0995;
    29: op1_05_in20 = reg_0211;
    30: op1_05_in20 = imem01_in[99:96];
    31: op1_05_in20 = reg_1006;
    32: op1_05_in20 = imem06_in[95:92];
    33: op1_05_in20 = reg_0474;
    34: op1_05_in20 = reg_0090;
    36: op1_05_in20 = reg_0717;
    39: op1_05_in20 = imem01_in[7:4];
    40: op1_05_in20 = reg_0245;
    53: op1_05_in20 = reg_0245;
    41: op1_05_in20 = reg_0248;
    42: op1_05_in20 = imem06_in[23:20];
    44: op1_05_in20 = reg_0003;
    45: op1_05_in20 = reg_1003;
    46: op1_05_in20 = reg_0783;
    48: op1_05_in20 = imem03_in[39:36];
    49: op1_05_in20 = imem07_in[63:60];
    50: op1_05_in20 = reg_0255;
    51: op1_05_in20 = imem04_in[71:68];
    52: op1_05_in20 = reg_1035;
    54: op1_05_in20 = imem04_in[119:116];
    55: op1_05_in20 = reg_0237;
    56: op1_05_in20 = reg_0333;
    57: op1_05_in20 = imem07_in[107:104];
    59: op1_05_in20 = reg_0735;
    60: op1_05_in20 = reg_0207;
    62: op1_05_in20 = reg_0192;
    63: op1_05_in20 = reg_0912;
    64: op1_05_in20 = imem05_in[67:64];
    65: op1_05_in20 = reg_0382;
    66: op1_05_in20 = reg_1011;
    67: op1_05_in20 = imem06_in[3:0];
    68: op1_05_in20 = reg_0353;
    69: op1_05_in20 = reg_0086;
    70: op1_05_in20 = reg_0693;
    71: op1_05_in20 = reg_0502;
    72: op1_05_in20 = reg_0777;
    73: op1_05_in20 = imem06_in[75:72];
    74: op1_05_in20 = reg_0403;
    76: op1_05_in20 = reg_1042;
    77: op1_05_in20 = imem01_in[103:100];
    84: op1_05_in20 = imem01_in[103:100];
    78: op1_05_in20 = reg_0886;
    79: op1_05_in20 = imem05_in[39:36];
    80: op1_05_in20 = reg_0889;
    81: op1_05_in20 = reg_0589;
    83: op1_05_in20 = reg_0823;
    85: op1_05_in20 = imem06_in[115:112];
    87: op1_05_in20 = reg_0040;
    88: op1_05_in20 = imem05_in[47:44];
    89: op1_05_in20 = reg_0521;
    90: op1_05_in20 = reg_0021;
    91: op1_05_in20 = reg_0029;
    92: op1_05_in20 = imem07_in[11:8];
    93: op1_05_in20 = reg_0514;
    94: op1_05_in20 = imem01_in[63:60];
    95: op1_05_in20 = reg_0236;
    96: op1_05_in20 = reg_0249;
    97: op1_05_in20 = reg_0449;
    default: op1_05_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv20 = 1;
    8: op1_05_inv20 = 1;
    11: op1_05_inv20 = 1;
    13: op1_05_inv20 = 1;
    14: op1_05_inv20 = 1;
    15: op1_05_inv20 = 1;
    16: op1_05_inv20 = 1;
    18: op1_05_inv20 = 1;
    20: op1_05_inv20 = 1;
    22: op1_05_inv20 = 1;
    27: op1_05_inv20 = 1;
    29: op1_05_inv20 = 1;
    31: op1_05_inv20 = 1;
    32: op1_05_inv20 = 1;
    33: op1_05_inv20 = 1;
    42: op1_05_inv20 = 1;
    46: op1_05_inv20 = 1;
    48: op1_05_inv20 = 1;
    49: op1_05_inv20 = 1;
    52: op1_05_inv20 = 1;
    55: op1_05_inv20 = 1;
    56: op1_05_inv20 = 1;
    57: op1_05_inv20 = 1;
    60: op1_05_inv20 = 1;
    63: op1_05_inv20 = 1;
    65: op1_05_inv20 = 1;
    72: op1_05_inv20 = 1;
    73: op1_05_inv20 = 1;
    78: op1_05_inv20 = 1;
    79: op1_05_inv20 = 1;
    81: op1_05_inv20 = 1;
    82: op1_05_inv20 = 1;
    83: op1_05_inv20 = 1;
    84: op1_05_inv20 = 1;
    85: op1_05_inv20 = 1;
    87: op1_05_inv20 = 1;
    89: op1_05_inv20 = 1;
    92: op1_05_inv20 = 1;
    93: op1_05_inv20 = 1;
    95: op1_05_inv20 = 1;
    default: op1_05_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in21 = reg_0516;
    6: op1_05_in21 = reg_0182;
    7: op1_05_in21 = reg_0594;
    8: op1_05_in21 = imem06_in[79:76];
    9: op1_05_in21 = imem01_in[95:92];
    10: op1_05_in21 = reg_1010;
    11: op1_05_in21 = reg_0789;
    13: op1_05_in21 = reg_0989;
    14: op1_05_in21 = imem06_in[103:100];
    16: op1_05_in21 = reg_0077;
    17: op1_05_in21 = reg_0290;
    18: op1_05_in21 = reg_0735;
    19: op1_05_in21 = reg_0949;
    20: op1_05_in21 = reg_0507;
    63: op1_05_in21 = reg_0507;
    21: op1_05_in21 = reg_0955;
    22: op1_05_in21 = reg_0213;
    23: op1_05_in21 = imem01_in[83:80];
    24: op1_05_in21 = reg_0729;
    25: op1_05_in21 = reg_0884;
    26: op1_05_in21 = reg_0774;
    27: op1_05_in21 = imem03_in[27:24];
    28: op1_05_in21 = reg_0999;
    29: op1_05_in21 = reg_0190;
    30: op1_05_in21 = imem01_in[119:116];
    31: op1_05_in21 = reg_0511;
    32: op1_05_in21 = imem07_in[23:20];
    33: op1_05_in21 = reg_0203;
    34: op1_05_in21 = reg_0049;
    36: op1_05_in21 = reg_0725;
    39: op1_05_in21 = imem01_in[43:40];
    40: op1_05_in21 = reg_0346;
    53: op1_05_in21 = reg_0346;
    41: op1_05_in21 = imem01_in[27:24];
    42: op1_05_in21 = imem06_in[63:60];
    44: op1_05_in21 = reg_0555;
    45: op1_05_in21 = reg_0799;
    46: op1_05_in21 = reg_0042;
    47: op1_05_in21 = imem01_in[47:44];
    48: op1_05_in21 = imem03_in[43:40];
    49: op1_05_in21 = imem07_in[75:72];
    50: op1_05_in21 = reg_0963;
    51: op1_05_in21 = imem04_in[75:72];
    52: op1_05_in21 = reg_0236;
    54: op1_05_in21 = reg_1004;
    55: op1_05_in21 = reg_0448;
    56: op1_05_in21 = reg_0149;
    57: op1_05_in21 = imem07_in[119:116];
    59: op1_05_in21 = reg_0534;
    80: op1_05_in21 = reg_0534;
    60: op1_05_in21 = reg_0196;
    62: op1_05_in21 = imem01_in[19:16];
    64: op1_05_in21 = imem05_in[111:108];
    65: op1_05_in21 = reg_0591;
    66: op1_05_in21 = reg_0926;
    67: op1_05_in21 = reg_1019;
    68: op1_05_in21 = reg_0350;
    69: op1_05_in21 = reg_0090;
    70: op1_05_in21 = reg_0217;
    71: op1_05_in21 = reg_0838;
    72: op1_05_in21 = reg_0044;
    73: op1_05_in21 = imem06_in[123:120];
    74: op1_05_in21 = reg_0022;
    76: op1_05_in21 = reg_0234;
    77: op1_05_in21 = reg_0969;
    78: op1_05_in21 = reg_0763;
    79: op1_05_in21 = imem05_in[55:52];
    81: op1_05_in21 = reg_0502;
    82: op1_05_in21 = reg_0755;
    83: op1_05_in21 = reg_0571;
    84: op1_05_in21 = imem01_in[123:120];
    85: op1_05_in21 = reg_0660;
    87: op1_05_in21 = reg_0767;
    88: op1_05_in21 = imem05_in[51:48];
    89: op1_05_in21 = reg_0610;
    90: op1_05_in21 = reg_0338;
    91: op1_05_in21 = reg_0719;
    92: op1_05_in21 = imem07_in[19:16];
    93: op1_05_in21 = reg_0276;
    95: op1_05_in21 = reg_0276;
    94: op1_05_in21 = imem01_in[67:64];
    96: op1_05_in21 = imem01_in[35:32];
    97: op1_05_in21 = reg_0529;
    default: op1_05_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv21 = 1;
    7: op1_05_inv21 = 1;
    9: op1_05_inv21 = 1;
    18: op1_05_inv21 = 1;
    21: op1_05_inv21 = 1;
    24: op1_05_inv21 = 1;
    25: op1_05_inv21 = 1;
    26: op1_05_inv21 = 1;
    28: op1_05_inv21 = 1;
    29: op1_05_inv21 = 1;
    30: op1_05_inv21 = 1;
    31: op1_05_inv21 = 1;
    33: op1_05_inv21 = 1;
    34: op1_05_inv21 = 1;
    40: op1_05_inv21 = 1;
    41: op1_05_inv21 = 1;
    42: op1_05_inv21 = 1;
    44: op1_05_inv21 = 1;
    45: op1_05_inv21 = 1;
    49: op1_05_inv21 = 1;
    50: op1_05_inv21 = 1;
    59: op1_05_inv21 = 1;
    62: op1_05_inv21 = 1;
    69: op1_05_inv21 = 1;
    71: op1_05_inv21 = 1;
    72: op1_05_inv21 = 1;
    73: op1_05_inv21 = 1;
    76: op1_05_inv21 = 1;
    83: op1_05_inv21 = 1;
    89: op1_05_inv21 = 1;
    90: op1_05_inv21 = 1;
    91: op1_05_inv21 = 1;
    93: op1_05_inv21 = 1;
    94: op1_05_inv21 = 1;
    95: op1_05_inv21 = 1;
    default: op1_05_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in22 = reg_0505;
    6: op1_05_in22 = reg_0160;
    7: op1_05_in22 = reg_0580;
    8: op1_05_in22 = reg_0606;
    9: op1_05_in22 = imem01_in[119:116];
    10: op1_05_in22 = reg_1011;
    11: op1_05_in22 = reg_0794;
    13: op1_05_in22 = imem04_in[55:52];
    14: op1_05_in22 = imem06_in[111:108];
    16: op1_05_in22 = reg_0079;
    17: op1_05_in22 = reg_0296;
    18: op1_05_in22 = reg_0766;
    19: op1_05_in22 = reg_0947;
    20: op1_05_in22 = reg_0869;
    21: op1_05_in22 = reg_0954;
    22: op1_05_in22 = reg_0212;
    23: op1_05_in22 = imem01_in[95:92];
    24: op1_05_in22 = reg_0427;
    25: op1_05_in22 = imem03_in[19:16];
    26: op1_05_in22 = imem05_in[11:8];
    27: op1_05_in22 = imem03_in[47:44];
    28: op1_05_in22 = reg_0981;
    29: op1_05_in22 = reg_0202;
    30: op1_05_in22 = reg_0810;
    31: op1_05_in22 = reg_0265;
    32: op1_05_in22 = imem07_in[39:36];
    33: op1_05_in22 = reg_0198;
    34: op1_05_in22 = reg_0872;
    36: op1_05_in22 = reg_0703;
    39: op1_05_in22 = imem01_in[71:68];
    40: op1_05_in22 = reg_0396;
    41: op1_05_in22 = imem01_in[55:52];
    42: op1_05_in22 = imem06_in[99:96];
    44: op1_05_in22 = reg_0249;
    45: op1_05_in22 = reg_0848;
    46: op1_05_in22 = reg_0351;
    47: op1_05_in22 = imem01_in[67:64];
    96: op1_05_in22 = imem01_in[67:64];
    48: op1_05_in22 = imem03_in[67:64];
    49: op1_05_in22 = imem07_in[83:80];
    50: op1_05_in22 = reg_0956;
    51: op1_05_in22 = imem04_in[95:92];
    52: op1_05_in22 = reg_0522;
    53: op1_05_in22 = reg_0824;
    54: op1_05_in22 = reg_1003;
    55: op1_05_in22 = reg_0148;
    56: op1_05_in22 = reg_0150;
    57: op1_05_in22 = imem07_in[123:120];
    59: op1_05_in22 = reg_0395;
    60: op1_05_in22 = imem01_in[3:0];
    62: op1_05_in22 = imem01_in[75:72];
    63: op1_05_in22 = reg_0850;
    64: op1_05_in22 = reg_0940;
    65: op1_05_in22 = reg_0863;
    66: op1_05_in22 = reg_0754;
    67: op1_05_in22 = reg_0691;
    68: op1_05_in22 = reg_0024;
    69: op1_05_in22 = reg_0049;
    70: op1_05_in22 = reg_0651;
    71: op1_05_in22 = reg_0167;
    72: op1_05_in22 = imem05_in[39:36];
    73: op1_05_in22 = reg_0344;
    74: op1_05_in22 = reg_0566;
    76: op1_05_in22 = reg_1024;
    77: op1_05_in22 = reg_0246;
    78: op1_05_in22 = reg_0908;
    79: op1_05_in22 = imem05_in[95:92];
    80: op1_05_in22 = reg_0533;
    81: op1_05_in22 = reg_0640;
    82: op1_05_in22 = reg_0022;
    83: op1_05_in22 = reg_0239;
    84: op1_05_in22 = reg_0234;
    85: op1_05_in22 = reg_0080;
    87: op1_05_in22 = reg_0385;
    88: op1_05_in22 = imem05_in[75:72];
    89: op1_05_in22 = reg_0906;
    90: op1_05_in22 = reg_0229;
    91: op1_05_in22 = reg_0380;
    92: op1_05_in22 = imem07_in[43:40];
    93: op1_05_in22 = reg_0225;
    94: op1_05_in22 = imem01_in[99:96];
    95: op1_05_in22 = reg_0544;
    97: op1_05_in22 = reg_0371;
    default: op1_05_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    16: op1_05_inv22 = 1;
    18: op1_05_inv22 = 1;
    20: op1_05_inv22 = 1;
    22: op1_05_inv22 = 1;
    24: op1_05_inv22 = 1;
    25: op1_05_inv22 = 1;
    26: op1_05_inv22 = 1;
    28: op1_05_inv22 = 1;
    30: op1_05_inv22 = 1;
    31: op1_05_inv22 = 1;
    32: op1_05_inv22 = 1;
    34: op1_05_inv22 = 1;
    39: op1_05_inv22 = 1;
    41: op1_05_inv22 = 1;
    44: op1_05_inv22 = 1;
    49: op1_05_inv22 = 1;
    50: op1_05_inv22 = 1;
    54: op1_05_inv22 = 1;
    56: op1_05_inv22 = 1;
    57: op1_05_inv22 = 1;
    59: op1_05_inv22 = 1;
    60: op1_05_inv22 = 1;
    62: op1_05_inv22 = 1;
    64: op1_05_inv22 = 1;
    66: op1_05_inv22 = 1;
    67: op1_05_inv22 = 1;
    68: op1_05_inv22 = 1;
    73: op1_05_inv22 = 1;
    76: op1_05_inv22 = 1;
    77: op1_05_inv22 = 1;
    80: op1_05_inv22 = 1;
    83: op1_05_inv22 = 1;
    85: op1_05_inv22 = 1;
    87: op1_05_inv22 = 1;
    94: op1_05_inv22 = 1;
    95: op1_05_inv22 = 1;
    default: op1_05_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in23 = reg_0235;
    6: op1_05_in23 = reg_0168;
    7: op1_05_in23 = reg_0595;
    8: op1_05_in23 = reg_0402;
    9: op1_05_in23 = reg_0512;
    10: op1_05_in23 = reg_0754;
    11: op1_05_in23 = reg_0791;
    13: op1_05_in23 = imem04_in[59:56];
    14: op1_05_in23 = reg_0629;
    16: op1_05_in23 = imem03_in[35:32];
    17: op1_05_in23 = reg_0292;
    18: op1_05_in23 = reg_0487;
    19: op1_05_in23 = reg_0953;
    20: op1_05_in23 = reg_0885;
    21: op1_05_in23 = reg_0957;
    22: op1_05_in23 = imem01_in[11:8];
    23: op1_05_in23 = reg_0013;
    24: op1_05_in23 = reg_0420;
    25: op1_05_in23 = imem03_in[47:44];
    26: op1_05_in23 = imem05_in[39:36];
    27: op1_05_in23 = imem03_in[83:80];
    28: op1_05_in23 = reg_0977;
    29: op1_05_in23 = imem01_in[63:60];
    30: op1_05_in23 = reg_0860;
    31: op1_05_in23 = reg_0277;
    54: op1_05_in23 = reg_0277;
    32: op1_05_in23 = imem07_in[43:40];
    33: op1_05_in23 = reg_0195;
    34: op1_05_in23 = imem03_in[59:56];
    36: op1_05_in23 = reg_0729;
    39: op1_05_in23 = imem01_in[79:76];
    40: op1_05_in23 = reg_0823;
    53: op1_05_in23 = reg_0823;
    41: op1_05_in23 = imem01_in[75:72];
    96: op1_05_in23 = imem01_in[75:72];
    42: op1_05_in23 = imem06_in[123:120];
    44: op1_05_in23 = reg_1039;
    45: op1_05_in23 = reg_0058;
    63: op1_05_in23 = reg_0058;
    46: op1_05_in23 = reg_0391;
    47: op1_05_in23 = imem01_in[87:84];
    48: op1_05_in23 = imem03_in[99:96];
    49: op1_05_in23 = reg_0716;
    50: op1_05_in23 = reg_0950;
    70: op1_05_in23 = reg_0950;
    51: op1_05_in23 = imem04_in[107:104];
    52: op1_05_in23 = reg_0829;
    55: op1_05_in23 = reg_0135;
    56: op1_05_in23 = reg_0151;
    57: op1_05_in23 = reg_0722;
    59: op1_05_in23 = reg_0591;
    60: op1_05_in23 = imem01_in[43:40];
    62: op1_05_in23 = imem01_in[91:88];
    64: op1_05_in23 = reg_0491;
    65: op1_05_in23 = reg_0222;
    66: op1_05_in23 = reg_0534;
    67: op1_05_in23 = reg_0262;
    68: op1_05_in23 = reg_0182;
    69: op1_05_in23 = reg_0884;
    71: op1_05_in23 = reg_0160;
    72: op1_05_in23 = imem05_in[67:64];
    73: op1_05_in23 = reg_1011;
    74: op1_05_in23 = imem07_in[51:48];
    76: op1_05_in23 = reg_0962;
    77: op1_05_in23 = reg_0973;
    78: op1_05_in23 = reg_0095;
    79: op1_05_in23 = imem05_in[99:96];
    80: op1_05_in23 = reg_0698;
    81: op1_05_in23 = reg_0838;
    82: op1_05_in23 = reg_0758;
    83: op1_05_in23 = reg_0040;
    84: op1_05_in23 = reg_0225;
    85: op1_05_in23 = reg_1019;
    87: op1_05_in23 = reg_0588;
    88: op1_05_in23 = imem05_in[87:84];
    89: op1_05_in23 = reg_1055;
    90: op1_05_in23 = reg_0889;
    91: op1_05_in23 = reg_0084;
    92: op1_05_in23 = imem07_in[47:44];
    93: op1_05_in23 = reg_0105;
    94: op1_05_in23 = imem01_in[107:104];
    95: op1_05_in23 = reg_0368;
    97: op1_05_in23 = reg_0184;
    default: op1_05_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv23 = 1;
    6: op1_05_inv23 = 1;
    7: op1_05_inv23 = 1;
    8: op1_05_inv23 = 1;
    9: op1_05_inv23 = 1;
    13: op1_05_inv23 = 1;
    20: op1_05_inv23 = 1;
    21: op1_05_inv23 = 1;
    22: op1_05_inv23 = 1;
    24: op1_05_inv23 = 1;
    28: op1_05_inv23 = 1;
    32: op1_05_inv23 = 1;
    33: op1_05_inv23 = 1;
    36: op1_05_inv23 = 1;
    39: op1_05_inv23 = 1;
    40: op1_05_inv23 = 1;
    41: op1_05_inv23 = 1;
    42: op1_05_inv23 = 1;
    45: op1_05_inv23 = 1;
    46: op1_05_inv23 = 1;
    47: op1_05_inv23 = 1;
    48: op1_05_inv23 = 1;
    49: op1_05_inv23 = 1;
    51: op1_05_inv23 = 1;
    52: op1_05_inv23 = 1;
    53: op1_05_inv23 = 1;
    54: op1_05_inv23 = 1;
    59: op1_05_inv23 = 1;
    64: op1_05_inv23 = 1;
    68: op1_05_inv23 = 1;
    76: op1_05_inv23 = 1;
    77: op1_05_inv23 = 1;
    78: op1_05_inv23 = 1;
    80: op1_05_inv23 = 1;
    82: op1_05_inv23 = 1;
    83: op1_05_inv23 = 1;
    90: op1_05_inv23 = 1;
    91: op1_05_inv23 = 1;
    94: op1_05_inv23 = 1;
    95: op1_05_inv23 = 1;
    default: op1_05_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in24 = reg_0227;
    52: op1_05_in24 = reg_0227;
    6: op1_05_in24 = reg_0157;
    68: op1_05_in24 = reg_0157;
    7: op1_05_in24 = reg_0394;
    8: op1_05_in24 = reg_0356;
    9: op1_05_in24 = reg_0503;
    10: op1_05_in24 = imem07_in[3:0];
    11: op1_05_in24 = reg_0224;
    13: op1_05_in24 = imem04_in[111:108];
    14: op1_05_in24 = reg_0624;
    16: op1_05_in24 = imem03_in[55:52];
    17: op1_05_in24 = reg_0295;
    18: op1_05_in24 = reg_0507;
    19: op1_05_in24 = reg_0865;
    20: op1_05_in24 = reg_1037;
    21: op1_05_in24 = reg_0950;
    22: op1_05_in24 = imem01_in[35:32];
    23: op1_05_in24 = reg_1051;
    24: op1_05_in24 = reg_0175;
    25: op1_05_in24 = imem03_in[51:48];
    26: op1_05_in24 = imem05_in[67:64];
    27: op1_05_in24 = imem03_in[91:88];
    28: op1_05_in24 = reg_0988;
    29: op1_05_in24 = imem01_in[79:76];
    30: op1_05_in24 = reg_0236;
    31: op1_05_in24 = reg_0306;
    32: op1_05_in24 = imem07_in[63:60];
    33: op1_05_in24 = reg_0199;
    34: op1_05_in24 = imem03_in[79:76];
    36: op1_05_in24 = reg_0418;
    39: op1_05_in24 = imem01_in[87:84];
    40: op1_05_in24 = reg_0874;
    41: op1_05_in24 = reg_0100;
    42: op1_05_in24 = reg_0883;
    44: op1_05_in24 = reg_0737;
    45: op1_05_in24 = reg_0302;
    46: op1_05_in24 = reg_0399;
    47: op1_05_in24 = imem01_in[103:100];
    48: op1_05_in24 = imem03_in[107:104];
    49: op1_05_in24 = reg_0726;
    50: op1_05_in24 = reg_0964;
    51: op1_05_in24 = imem04_in[115:112];
    53: op1_05_in24 = reg_0847;
    54: op1_05_in24 = reg_0912;
    55: op1_05_in24 = reg_0128;
    56: op1_05_in24 = reg_0128;
    57: op1_05_in24 = reg_0719;
    59: op1_05_in24 = reg_0695;
    60: op1_05_in24 = imem01_in[55:52];
    62: op1_05_in24 = reg_0779;
    63: op1_05_in24 = reg_0067;
    64: op1_05_in24 = reg_0030;
    65: op1_05_in24 = reg_0946;
    66: op1_05_in24 = reg_0556;
    67: op1_05_in24 = reg_0692;
    90: op1_05_in24 = reg_0692;
    69: op1_05_in24 = imem03_in[75:72];
    70: op1_05_in24 = reg_0343;
    71: op1_05_in24 = reg_0185;
    72: op1_05_in24 = imem05_in[91:88];
    73: op1_05_in24 = reg_1030;
    74: op1_05_in24 = imem07_in[79:76];
    76: op1_05_in24 = reg_0904;
    77: op1_05_in24 = reg_0968;
    78: op1_05_in24 = reg_0664;
    79: op1_05_in24 = reg_0145;
    80: op1_05_in24 = reg_0011;
    81: op1_05_in24 = reg_0431;
    82: op1_05_in24 = reg_0757;
    83: op1_05_in24 = reg_0773;
    84: op1_05_in24 = reg_1039;
    85: op1_05_in24 = reg_0926;
    87: op1_05_in24 = reg_0266;
    88: op1_05_in24 = reg_0215;
    89: op1_05_in24 = reg_0283;
    91: op1_05_in24 = imem07_in[15:12];
    92: op1_05_in24 = imem07_in[55:52];
    93: op1_05_in24 = reg_1023;
    94: op1_05_in24 = imem01_in[123:120];
    95: op1_05_in24 = reg_0304;
    96: op1_05_in24 = reg_0522;
    default: op1_05_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv24 = 1;
    11: op1_05_inv24 = 1;
    14: op1_05_inv24 = 1;
    21: op1_05_inv24 = 1;
    23: op1_05_inv24 = 1;
    24: op1_05_inv24 = 1;
    25: op1_05_inv24 = 1;
    27: op1_05_inv24 = 1;
    29: op1_05_inv24 = 1;
    30: op1_05_inv24 = 1;
    31: op1_05_inv24 = 1;
    32: op1_05_inv24 = 1;
    39: op1_05_inv24 = 1;
    44: op1_05_inv24 = 1;
    45: op1_05_inv24 = 1;
    47: op1_05_inv24 = 1;
    52: op1_05_inv24 = 1;
    54: op1_05_inv24 = 1;
    55: op1_05_inv24 = 1;
    56: op1_05_inv24 = 1;
    59: op1_05_inv24 = 1;
    64: op1_05_inv24 = 1;
    65: op1_05_inv24 = 1;
    69: op1_05_inv24 = 1;
    72: op1_05_inv24 = 1;
    73: op1_05_inv24 = 1;
    74: op1_05_inv24 = 1;
    77: op1_05_inv24 = 1;
    78: op1_05_inv24 = 1;
    79: op1_05_inv24 = 1;
    83: op1_05_inv24 = 1;
    84: op1_05_inv24 = 1;
    88: op1_05_inv24 = 1;
    90: op1_05_inv24 = 1;
    93: op1_05_inv24 = 1;
    95: op1_05_inv24 = 1;
    default: op1_05_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in25 = reg_0220;
    7: op1_05_in25 = reg_0384;
    85: op1_05_in25 = reg_0384;
    8: op1_05_in25 = reg_0405;
    9: op1_05_in25 = reg_0506;
    10: op1_05_in25 = imem07_in[27:24];
    11: op1_05_in25 = reg_0795;
    13: op1_05_in25 = imem04_in[119:116];
    14: op1_05_in25 = reg_0618;
    16: op1_05_in25 = imem03_in[71:68];
    17: op1_05_in25 = reg_0307;
    18: op1_05_in25 = reg_0249;
    19: op1_05_in25 = reg_0149;
    20: op1_05_in25 = reg_0227;
    21: op1_05_in25 = reg_0953;
    22: op1_05_in25 = imem01_in[47:44];
    23: op1_05_in25 = reg_1055;
    24: op1_05_in25 = reg_0165;
    25: op1_05_in25 = imem03_in[55:52];
    26: op1_05_in25 = imem05_in[107:104];
    27: op1_05_in25 = imem03_in[115:112];
    28: op1_05_in25 = reg_0976;
    29: op1_05_in25 = imem01_in[107:104];
    60: op1_05_in25 = imem01_in[107:104];
    30: op1_05_in25 = reg_0496;
    84: op1_05_in25 = reg_0496;
    31: op1_05_in25 = reg_1057;
    54: op1_05_in25 = reg_1057;
    32: op1_05_in25 = reg_0719;
    33: op1_05_in25 = reg_0197;
    34: op1_05_in25 = imem03_in[111:108];
    36: op1_05_in25 = reg_0434;
    39: op1_05_in25 = imem01_in[95:92];
    40: op1_05_in25 = reg_0543;
    41: op1_05_in25 = reg_0126;
    42: op1_05_in25 = reg_0895;
    44: op1_05_in25 = reg_1041;
    45: op1_05_in25 = reg_0808;
    46: op1_05_in25 = reg_0804;
    47: op1_05_in25 = imem01_in[111:108];
    48: op1_05_in25 = reg_0317;
    49: op1_05_in25 = reg_0717;
    50: op1_05_in25 = reg_0943;
    51: op1_05_in25 = reg_0277;
    52: op1_05_in25 = reg_1040;
    53: op1_05_in25 = reg_0784;
    55: op1_05_in25 = reg_0152;
    56: op1_05_in25 = reg_0142;
    57: op1_05_in25 = reg_0729;
    59: op1_05_in25 = reg_0780;
    62: op1_05_in25 = reg_0223;
    63: op1_05_in25 = reg_0276;
    64: op1_05_in25 = reg_0237;
    65: op1_05_in25 = reg_0257;
    66: op1_05_in25 = reg_0699;
    67: op1_05_in25 = reg_0028;
    69: op1_05_in25 = imem03_in[87:84];
    70: op1_05_in25 = reg_0259;
    71: op1_05_in25 = reg_0176;
    72: op1_05_in25 = imem05_in[119:116];
    73: op1_05_in25 = reg_0439;
    74: op1_05_in25 = imem07_in[119:116];
    76: op1_05_in25 = reg_0829;
    77: op1_05_in25 = reg_1044;
    78: op1_05_in25 = reg_0087;
    79: op1_05_in25 = reg_0252;
    80: op1_05_in25 = reg_0380;
    81: op1_05_in25 = imem07_in[31:28];
    91: op1_05_in25 = imem07_in[31:28];
    82: op1_05_in25 = reg_0710;
    83: op1_05_in25 = reg_0377;
    87: op1_05_in25 = reg_0985;
    88: op1_05_in25 = reg_0826;
    89: op1_05_in25 = reg_1033;
    90: op1_05_in25 = reg_0297;
    92: op1_05_in25 = imem07_in[67:64];
    93: op1_05_in25 = imem01_in[39:36];
    94: op1_05_in25 = reg_0905;
    95: op1_05_in25 = reg_1039;
    96: op1_05_in25 = reg_0222;
    default: op1_05_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv25 = 1;
    11: op1_05_inv25 = 1;
    13: op1_05_inv25 = 1;
    14: op1_05_inv25 = 1;
    16: op1_05_inv25 = 1;
    17: op1_05_inv25 = 1;
    18: op1_05_inv25 = 1;
    19: op1_05_inv25 = 1;
    20: op1_05_inv25 = 1;
    21: op1_05_inv25 = 1;
    22: op1_05_inv25 = 1;
    23: op1_05_inv25 = 1;
    24: op1_05_inv25 = 1;
    26: op1_05_inv25 = 1;
    30: op1_05_inv25 = 1;
    31: op1_05_inv25 = 1;
    32: op1_05_inv25 = 1;
    33: op1_05_inv25 = 1;
    34: op1_05_inv25 = 1;
    36: op1_05_inv25 = 1;
    40: op1_05_inv25 = 1;
    41: op1_05_inv25 = 1;
    50: op1_05_inv25 = 1;
    51: op1_05_inv25 = 1;
    52: op1_05_inv25 = 1;
    53: op1_05_inv25 = 1;
    54: op1_05_inv25 = 1;
    55: op1_05_inv25 = 1;
    57: op1_05_inv25 = 1;
    59: op1_05_inv25 = 1;
    62: op1_05_inv25 = 1;
    64: op1_05_inv25 = 1;
    65: op1_05_inv25 = 1;
    66: op1_05_inv25 = 1;
    67: op1_05_inv25 = 1;
    69: op1_05_inv25 = 1;
    71: op1_05_inv25 = 1;
    73: op1_05_inv25 = 1;
    76: op1_05_inv25 = 1;
    78: op1_05_inv25 = 1;
    79: op1_05_inv25 = 1;
    81: op1_05_inv25 = 1;
    82: op1_05_inv25 = 1;
    87: op1_05_inv25 = 1;
    88: op1_05_inv25 = 1;
    90: op1_05_inv25 = 1;
    92: op1_05_inv25 = 1;
    93: op1_05_inv25 = 1;
    95: op1_05_inv25 = 1;
    default: op1_05_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in26 = reg_0236;
    7: op1_05_in26 = reg_0388;
    8: op1_05_in26 = reg_0371;
    42: op1_05_in26 = reg_0371;
    9: op1_05_in26 = reg_0510;
    10: op1_05_in26 = imem07_in[31:28];
    11: op1_05_in26 = reg_0221;
    13: op1_05_in26 = reg_0530;
    14: op1_05_in26 = reg_0379;
    16: op1_05_in26 = imem03_in[107:104];
    69: op1_05_in26 = imem03_in[107:104];
    17: op1_05_in26 = reg_0078;
    18: op1_05_in26 = reg_0227;
    19: op1_05_in26 = reg_0154;
    55: op1_05_in26 = reg_0154;
    20: op1_05_in26 = reg_0216;
    21: op1_05_in26 = reg_0960;
    22: op1_05_in26 = imem01_in[95:92];
    23: op1_05_in26 = reg_1053;
    24: op1_05_in26 = reg_0166;
    25: op1_05_in26 = imem03_in[59:56];
    26: op1_05_in26 = imem05_in[127:124];
    27: op1_05_in26 = reg_0582;
    28: op1_05_in26 = imem04_in[43:40];
    29: op1_05_in26 = imem01_in[111:108];
    60: op1_05_in26 = imem01_in[111:108];
    30: op1_05_in26 = reg_1037;
    31: op1_05_in26 = reg_0760;
    32: op1_05_in26 = reg_0726;
    82: op1_05_in26 = reg_0726;
    33: op1_05_in26 = imem01_in[19:16];
    34: op1_05_in26 = imem03_in[123:120];
    36: op1_05_in26 = reg_0443;
    39: op1_05_in26 = imem01_in[103:100];
    40: op1_05_in26 = reg_0767;
    41: op1_05_in26 = imem02_in[59:56];
    44: op1_05_in26 = reg_0906;
    76: op1_05_in26 = reg_0906;
    45: op1_05_in26 = reg_0288;
    46: op1_05_in26 = reg_0332;
    47: op1_05_in26 = reg_0779;
    48: op1_05_in26 = reg_0346;
    49: op1_05_in26 = reg_0725;
    50: op1_05_in26 = reg_0953;
    51: op1_05_in26 = reg_0282;
    52: op1_05_in26 = reg_0737;
    53: op1_05_in26 = reg_0836;
    54: op1_05_in26 = reg_1020;
    56: op1_05_in26 = reg_0140;
    57: op1_05_in26 = reg_0715;
    59: op1_05_in26 = reg_0609;
    62: op1_05_in26 = reg_0928;
    63: op1_05_in26 = reg_0584;
    64: op1_05_in26 = reg_0942;
    65: op1_05_in26 = reg_0605;
    66: op1_05_in26 = reg_0632;
    67: op1_05_in26 = reg_0895;
    70: op1_05_in26 = reg_0948;
    71: op1_05_in26 = reg_0171;
    72: op1_05_in26 = reg_0950;
    73: op1_05_in26 = reg_0834;
    74: op1_05_in26 = reg_0730;
    77: op1_05_in26 = reg_0546;
    78: op1_05_in26 = reg_0644;
    79: op1_05_in26 = reg_0816;
    80: op1_05_in26 = reg_0917;
    81: op1_05_in26 = imem07_in[43:40];
    83: op1_05_in26 = reg_0581;
    84: op1_05_in26 = reg_0604;
    85: op1_05_in26 = reg_0692;
    87: op1_05_in26 = reg_0982;
    88: op1_05_in26 = reg_0063;
    89: op1_05_in26 = reg_0101;
    90: op1_05_in26 = reg_0439;
    91: op1_05_in26 = imem07_in[39:36];
    92: op1_05_in26 = imem07_in[75:72];
    93: op1_05_in26 = imem01_in[63:60];
    94: op1_05_in26 = reg_0501;
    95: op1_05_in26 = reg_0122;
    96: op1_05_in26 = reg_0524;
    default: op1_05_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_05_inv26 = 1;
    9: op1_05_inv26 = 1;
    10: op1_05_inv26 = 1;
    11: op1_05_inv26 = 1;
    14: op1_05_inv26 = 1;
    16: op1_05_inv26 = 1;
    17: op1_05_inv26 = 1;
    18: op1_05_inv26 = 1;
    20: op1_05_inv26 = 1;
    21: op1_05_inv26 = 1;
    22: op1_05_inv26 = 1;
    23: op1_05_inv26 = 1;
    25: op1_05_inv26 = 1;
    27: op1_05_inv26 = 1;
    29: op1_05_inv26 = 1;
    32: op1_05_inv26 = 1;
    33: op1_05_inv26 = 1;
    34: op1_05_inv26 = 1;
    36: op1_05_inv26 = 1;
    40: op1_05_inv26 = 1;
    42: op1_05_inv26 = 1;
    44: op1_05_inv26 = 1;
    48: op1_05_inv26 = 1;
    49: op1_05_inv26 = 1;
    52: op1_05_inv26 = 1;
    53: op1_05_inv26 = 1;
    59: op1_05_inv26 = 1;
    60: op1_05_inv26 = 1;
    62: op1_05_inv26 = 1;
    66: op1_05_inv26 = 1;
    69: op1_05_inv26 = 1;
    71: op1_05_inv26 = 1;
    72: op1_05_inv26 = 1;
    78: op1_05_inv26 = 1;
    79: op1_05_inv26 = 1;
    80: op1_05_inv26 = 1;
    81: op1_05_inv26 = 1;
    82: op1_05_inv26 = 1;
    85: op1_05_inv26 = 1;
    91: op1_05_inv26 = 1;
    93: op1_05_inv26 = 1;
    96: op1_05_inv26 = 1;
    default: op1_05_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in27 = reg_0237;
    7: op1_05_in27 = reg_0323;
    8: op1_05_in27 = reg_0375;
    9: op1_05_in27 = reg_0507;
    10: op1_05_in27 = imem07_in[39:36];
    11: op1_05_in27 = reg_0219;
    13: op1_05_in27 = reg_0542;
    14: op1_05_in27 = reg_0351;
    16: op1_05_in27 = reg_0602;
    17: op1_05_in27 = reg_0062;
    18: op1_05_in27 = reg_0123;
    19: op1_05_in27 = reg_0138;
    20: op1_05_in27 = reg_1031;
    21: op1_05_in27 = reg_0834;
    22: op1_05_in27 = imem01_in[115:112];
    23: op1_05_in27 = reg_0239;
    24: op1_05_in27 = reg_0177;
    25: op1_05_in27 = imem03_in[127:124];
    26: op1_05_in27 = reg_0949;
    27: op1_05_in27 = reg_0571;
    28: op1_05_in27 = imem04_in[51:48];
    29: op1_05_in27 = reg_0786;
    30: op1_05_in27 = reg_0871;
    31: op1_05_in27 = reg_0065;
    32: op1_05_in27 = reg_0715;
    33: op1_05_in27 = imem01_in[43:40];
    34: op1_05_in27 = reg_0343;
    36: op1_05_in27 = reg_0420;
    39: op1_05_in27 = reg_0510;
    40: op1_05_in27 = reg_0376;
    53: op1_05_in27 = reg_0376;
    41: op1_05_in27 = imem02_in[79:76];
    42: op1_05_in27 = reg_0556;
    44: op1_05_in27 = reg_0122;
    45: op1_05_in27 = reg_0283;
    46: op1_05_in27 = reg_0017;
    73: op1_05_in27 = reg_0017;
    47: op1_05_in27 = reg_0828;
    48: op1_05_in27 = reg_0807;
    49: op1_05_in27 = reg_0709;
    50: op1_05_in27 = imem05_in[47:44];
    51: op1_05_in27 = reg_0539;
    52: op1_05_in27 = reg_0906;
    54: op1_05_in27 = reg_0292;
    55: op1_05_in27 = imem06_in[3:0];
    79: op1_05_in27 = imem06_in[3:0];
    56: op1_05_in27 = imem06_in[71:68];
    57: op1_05_in27 = reg_0002;
    59: op1_05_in27 = imem07_in[7:4];
    60: op1_05_in27 = imem01_in[119:116];
    62: op1_05_in27 = reg_0242;
    63: op1_05_in27 = reg_0074;
    64: op1_05_in27 = reg_0750;
    65: op1_05_in27 = reg_0405;
    66: op1_05_in27 = reg_0915;
    67: op1_05_in27 = reg_0699;
    69: op1_05_in27 = reg_1007;
    70: op1_05_in27 = reg_0004;
    72: op1_05_in27 = reg_0945;
    74: op1_05_in27 = reg_0726;
    76: op1_05_in27 = reg_1055;
    77: op1_05_in27 = reg_0592;
    78: op1_05_in27 = reg_0335;
    80: op1_05_in27 = imem07_in[51:48];
    81: op1_05_in27 = imem07_in[67:64];
    82: op1_05_in27 = reg_0563;
    83: op1_05_in27 = reg_1001;
    84: op1_05_in27 = reg_0829;
    85: op1_05_in27 = reg_0613;
    87: op1_05_in27 = reg_0980;
    88: op1_05_in27 = reg_0964;
    89: op1_05_in27 = imem02_in[3:0];
    90: op1_05_in27 = reg_0264;
    91: op1_05_in27 = reg_0159;
    92: op1_05_in27 = imem07_in[83:80];
    93: op1_05_in27 = imem01_in[111:108];
    94: op1_05_in27 = reg_0798;
    95: op1_05_in27 = reg_0059;
    96: op1_05_in27 = reg_0409;
    default: op1_05_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv27 = 1;
    7: op1_05_inv27 = 1;
    8: op1_05_inv27 = 1;
    9: op1_05_inv27 = 1;
    16: op1_05_inv27 = 1;
    17: op1_05_inv27 = 1;
    18: op1_05_inv27 = 1;
    23: op1_05_inv27 = 1;
    26: op1_05_inv27 = 1;
    27: op1_05_inv27 = 1;
    28: op1_05_inv27 = 1;
    29: op1_05_inv27 = 1;
    30: op1_05_inv27 = 1;
    33: op1_05_inv27 = 1;
    34: op1_05_inv27 = 1;
    39: op1_05_inv27 = 1;
    41: op1_05_inv27 = 1;
    45: op1_05_inv27 = 1;
    46: op1_05_inv27 = 1;
    47: op1_05_inv27 = 1;
    49: op1_05_inv27 = 1;
    51: op1_05_inv27 = 1;
    53: op1_05_inv27 = 1;
    54: op1_05_inv27 = 1;
    55: op1_05_inv27 = 1;
    57: op1_05_inv27 = 1;
    60: op1_05_inv27 = 1;
    65: op1_05_inv27 = 1;
    77: op1_05_inv27 = 1;
    79: op1_05_inv27 = 1;
    82: op1_05_inv27 = 1;
    87: op1_05_inv27 = 1;
    91: op1_05_inv27 = 1;
    92: op1_05_inv27 = 1;
    93: op1_05_inv27 = 1;
    95: op1_05_inv27 = 1;
    default: op1_05_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in28 = reg_0238;
    7: op1_05_in28 = reg_0312;
    8: op1_05_in28 = reg_0383;
    9: op1_05_in28 = reg_0505;
    10: op1_05_in28 = imem07_in[59:56];
    80: op1_05_in28 = imem07_in[59:56];
    11: op1_05_in28 = imem01_in[115:112];
    13: op1_05_in28 = reg_0529;
    14: op1_05_in28 = reg_0337;
    16: op1_05_in28 = reg_0573;
    27: op1_05_in28 = reg_0573;
    17: op1_05_in28 = reg_0065;
    18: op1_05_in28 = imem02_in[19:16];
    19: op1_05_in28 = reg_0129;
    20: op1_05_in28 = reg_1045;
    21: op1_05_in28 = reg_0835;
    73: op1_05_in28 = reg_0835;
    22: op1_05_in28 = reg_0239;
    23: op1_05_in28 = reg_0735;
    24: op1_05_in28 = reg_0158;
    25: op1_05_in28 = reg_0582;
    26: op1_05_in28 = reg_0968;
    28: op1_05_in28 = imem04_in[71:68];
    29: op1_05_in28 = reg_0003;
    30: op1_05_in28 = reg_1038;
    31: op1_05_in28 = reg_0071;
    32: op1_05_in28 = reg_0707;
    49: op1_05_in28 = reg_0707;
    33: op1_05_in28 = imem01_in[59:56];
    34: op1_05_in28 = reg_0581;
    36: op1_05_in28 = reg_0431;
    39: op1_05_in28 = reg_0487;
    40: op1_05_in28 = reg_0844;
    41: op1_05_in28 = reg_0642;
    42: op1_05_in28 = reg_0577;
    44: op1_05_in28 = imem02_in[31:28];
    45: op1_05_in28 = reg_0528;
    46: op1_05_in28 = reg_0263;
    47: op1_05_in28 = reg_0236;
    48: op1_05_in28 = reg_0996;
    50: op1_05_in28 = imem05_in[67:64];
    51: op1_05_in28 = reg_1020;
    52: op1_05_in28 = reg_0122;
    53: op1_05_in28 = reg_0985;
    54: op1_05_in28 = reg_0050;
    55: op1_05_in28 = imem06_in[27:24];
    56: op1_05_in28 = reg_0534;
    57: op1_05_in28 = reg_0321;
    59: op1_05_in28 = imem07_in[11:8];
    60: op1_05_in28 = reg_0779;
    62: op1_05_in28 = reg_1035;
    63: op1_05_in28 = reg_0809;
    64: op1_05_in28 = reg_0508;
    65: op1_05_in28 = reg_0571;
    66: op1_05_in28 = reg_0264;
    67: op1_05_in28 = reg_0632;
    69: op1_05_in28 = reg_0661;
    70: op1_05_in28 = reg_0147;
    72: op1_05_in28 = reg_0343;
    74: op1_05_in28 = reg_0718;
    76: op1_05_in28 = reg_0112;
    77: op1_05_in28 = reg_0503;
    78: op1_05_in28 = reg_0007;
    79: op1_05_in28 = imem06_in[7:4];
    81: op1_05_in28 = imem07_in[107:104];
    82: op1_05_in28 = reg_0903;
    83: op1_05_in28 = reg_0309;
    84: op1_05_in28 = reg_0514;
    85: op1_05_in28 = reg_0392;
    87: op1_05_in28 = imem04_in[11:8];
    88: op1_05_in28 = reg_0831;
    89: op1_05_in28 = imem02_in[27:24];
    90: op1_05_in28 = reg_0822;
    91: op1_05_in28 = reg_0560;
    92: op1_05_in28 = imem07_in[119:116];
    93: op1_05_in28 = imem01_in[119:116];
    94: op1_05_in28 = reg_0619;
    95: op1_05_in28 = reg_0154;
    96: op1_05_in28 = reg_0737;
    default: op1_05_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv28 = 1;
    8: op1_05_inv28 = 1;
    9: op1_05_inv28 = 1;
    10: op1_05_inv28 = 1;
    13: op1_05_inv28 = 1;
    14: op1_05_inv28 = 1;
    16: op1_05_inv28 = 1;
    18: op1_05_inv28 = 1;
    19: op1_05_inv28 = 1;
    20: op1_05_inv28 = 1;
    21: op1_05_inv28 = 1;
    23: op1_05_inv28 = 1;
    25: op1_05_inv28 = 1;
    27: op1_05_inv28 = 1;
    30: op1_05_inv28 = 1;
    31: op1_05_inv28 = 1;
    33: op1_05_inv28 = 1;
    44: op1_05_inv28 = 1;
    45: op1_05_inv28 = 1;
    46: op1_05_inv28 = 1;
    47: op1_05_inv28 = 1;
    48: op1_05_inv28 = 1;
    50: op1_05_inv28 = 1;
    54: op1_05_inv28 = 1;
    56: op1_05_inv28 = 1;
    57: op1_05_inv28 = 1;
    60: op1_05_inv28 = 1;
    63: op1_05_inv28 = 1;
    64: op1_05_inv28 = 1;
    70: op1_05_inv28 = 1;
    73: op1_05_inv28 = 1;
    76: op1_05_inv28 = 1;
    79: op1_05_inv28 = 1;
    80: op1_05_inv28 = 1;
    81: op1_05_inv28 = 1;
    82: op1_05_inv28 = 1;
    83: op1_05_inv28 = 1;
    84: op1_05_inv28 = 1;
    87: op1_05_inv28 = 1;
    90: op1_05_inv28 = 1;
    93: op1_05_inv28 = 1;
    94: op1_05_inv28 = 1;
    default: op1_05_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in29 = reg_0119;
    7: op1_05_in29 = reg_0393;
    8: op1_05_in29 = reg_0404;
    9: op1_05_in29 = reg_0238;
    10: op1_05_in29 = imem07_in[83:80];
    11: op1_05_in29 = reg_0226;
    13: op1_05_in29 = reg_0539;
    14: op1_05_in29 = reg_0026;
    16: op1_05_in29 = reg_0568;
    17: op1_05_in29 = reg_0067;
    18: op1_05_in29 = imem02_in[35:32];
    19: op1_05_in29 = reg_0134;
    20: op1_05_in29 = reg_1034;
    21: op1_05_in29 = reg_0827;
    22: op1_05_in29 = reg_0236;
    23: op1_05_in29 = reg_0487;
    24: op1_05_in29 = reg_0173;
    25: op1_05_in29 = reg_0571;
    26: op1_05_in29 = reg_0952;
    27: op1_05_in29 = reg_0583;
    28: op1_05_in29 = imem04_in[95:92];
    29: op1_05_in29 = reg_0905;
    30: op1_05_in29 = reg_0904;
    31: op1_05_in29 = reg_0015;
    32: op1_05_in29 = reg_0434;
    33: op1_05_in29 = reg_0003;
    34: op1_05_in29 = reg_0396;
    36: op1_05_in29 = reg_0162;
    39: op1_05_in29 = reg_1039;
    40: op1_05_in29 = reg_0234;
    41: op1_05_in29 = reg_0653;
    42: op1_05_in29 = reg_0349;
    65: op1_05_in29 = reg_0349;
    44: op1_05_in29 = imem02_in[43:40];
    45: op1_05_in29 = reg_0043;
    46: op1_05_in29 = imem07_in[23:20];
    47: op1_05_in29 = reg_0274;
    62: op1_05_in29 = reg_0274;
    48: op1_05_in29 = reg_0994;
    49: op1_05_in29 = reg_0361;
    50: op1_05_in29 = reg_0147;
    51: op1_05_in29 = reg_0292;
    52: op1_05_in29 = reg_0124;
    53: op1_05_in29 = reg_0998;
    54: op1_05_in29 = reg_0802;
    55: op1_05_in29 = imem06_in[47:44];
    56: op1_05_in29 = reg_0895;
    57: op1_05_in29 = reg_0024;
    59: op1_05_in29 = imem07_in[15:12];
    60: op1_05_in29 = reg_0223;
    63: op1_05_in29 = imem05_in[7:4];
    64: op1_05_in29 = reg_0436;
    66: op1_05_in29 = reg_0399;
    67: op1_05_in29 = reg_0619;
    69: op1_05_in29 = reg_0874;
    70: op1_05_in29 = reg_0148;
    72: op1_05_in29 = reg_0486;
    73: op1_05_in29 = reg_0018;
    74: op1_05_in29 = reg_0727;
    76: op1_05_in29 = reg_0114;
    77: op1_05_in29 = reg_0829;
    78: op1_05_in29 = reg_0776;
    79: op1_05_in29 = imem06_in[55:52];
    80: op1_05_in29 = imem07_in[103:100];
    81: op1_05_in29 = imem07_in[115:112];
    82: op1_05_in29 = reg_0002;
    83: op1_05_in29 = reg_1003;
    84: op1_05_in29 = reg_0830;
    85: op1_05_in29 = reg_0617;
    87: op1_05_in29 = imem04_in[23:20];
    88: op1_05_in29 = reg_0706;
    89: op1_05_in29 = imem02_in[87:84];
    90: op1_05_in29 = reg_0320;
    91: op1_05_in29 = reg_0164;
    92: op1_05_in29 = imem07_in[127:124];
    93: op1_05_in29 = imem01_in[127:124];
    94: op1_05_in29 = reg_1056;
    95: op1_05_in29 = reg_0793;
    96: op1_05_in29 = reg_0221;
    default: op1_05_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv29 = 1;
    8: op1_05_inv29 = 1;
    13: op1_05_inv29 = 1;
    17: op1_05_inv29 = 1;
    18: op1_05_inv29 = 1;
    20: op1_05_inv29 = 1;
    21: op1_05_inv29 = 1;
    22: op1_05_inv29 = 1;
    23: op1_05_inv29 = 1;
    24: op1_05_inv29 = 1;
    25: op1_05_inv29 = 1;
    26: op1_05_inv29 = 1;
    27: op1_05_inv29 = 1;
    33: op1_05_inv29 = 1;
    40: op1_05_inv29 = 1;
    41: op1_05_inv29 = 1;
    44: op1_05_inv29 = 1;
    50: op1_05_inv29 = 1;
    51: op1_05_inv29 = 1;
    59: op1_05_inv29 = 1;
    60: op1_05_inv29 = 1;
    62: op1_05_inv29 = 1;
    63: op1_05_inv29 = 1;
    67: op1_05_inv29 = 1;
    69: op1_05_inv29 = 1;
    70: op1_05_inv29 = 1;
    72: op1_05_inv29 = 1;
    73: op1_05_inv29 = 1;
    76: op1_05_inv29 = 1;
    79: op1_05_inv29 = 1;
    81: op1_05_inv29 = 1;
    84: op1_05_inv29 = 1;
    85: op1_05_inv29 = 1;
    88: op1_05_inv29 = 1;
    89: op1_05_inv29 = 1;
    90: op1_05_inv29 = 1;
    91: op1_05_inv29 = 1;
    92: op1_05_inv29 = 1;
    95: op1_05_inv29 = 1;
    default: op1_05_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_05_in30 = reg_0120;
    9: op1_05_in30 = reg_0120;
    7: op1_05_in30 = reg_0389;
    8: op1_05_in30 = reg_0337;
    10: op1_05_in30 = reg_0719;
    11: op1_05_in30 = reg_0230;
    13: op1_05_in30 = reg_0281;
    14: op1_05_in30 = reg_0802;
    16: op1_05_in30 = reg_0584;
    17: op1_05_in30 = reg_0068;
    18: op1_05_in30 = imem02_in[67:64];
    19: op1_05_in30 = imem06_in[15:12];
    20: op1_05_in30 = reg_0103;
    21: op1_05_in30 = reg_0275;
    22: op1_05_in30 = reg_0487;
    23: op1_05_in30 = reg_1050;
    25: op1_05_in30 = reg_0599;
    26: op1_05_in30 = reg_0835;
    27: op1_05_in30 = reg_0568;
    28: op1_05_in30 = imem04_in[127:124];
    29: op1_05_in30 = reg_1042;
    39: op1_05_in30 = reg_1042;
    30: op1_05_in30 = reg_0127;
    31: op1_05_in30 = reg_0736;
    32: op1_05_in30 = reg_0435;
    33: op1_05_in30 = reg_0218;
    34: op1_05_in30 = reg_0874;
    36: op1_05_in30 = reg_0173;
    94: op1_05_in30 = reg_0173;
    40: op1_05_in30 = reg_0985;
    41: op1_05_in30 = reg_0646;
    42: op1_05_in30 = reg_0628;
    44: op1_05_in30 = imem02_in[71:68];
    45: op1_05_in30 = imem05_in[3:0];
    46: op1_05_in30 = imem07_in[63:60];
    47: op1_05_in30 = reg_0238;
    48: op1_05_in30 = imem04_in[51:48];
    49: op1_05_in30 = reg_0575;
    50: op1_05_in30 = reg_0145;
    70: op1_05_in30 = reg_0145;
    51: op1_05_in30 = reg_1016;
    52: op1_05_in30 = reg_0125;
    53: op1_05_in30 = reg_0992;
    54: op1_05_in30 = reg_0848;
    55: op1_05_in30 = imem06_in[79:76];
    56: op1_05_in30 = reg_0624;
    57: op1_05_in30 = reg_0431;
    59: op1_05_in30 = imem07_in[19:16];
    60: op1_05_in30 = reg_0936;
    62: op1_05_in30 = reg_0607;
    63: op1_05_in30 = imem05_in[59:56];
    64: op1_05_in30 = reg_0094;
    65: op1_05_in30 = imem07_in[47:44];
    66: op1_05_in30 = reg_0957;
    67: op1_05_in30 = reg_0408;
    69: op1_05_in30 = reg_0833;
    72: op1_05_in30 = reg_0963;
    73: op1_05_in30 = reg_0022;
    74: op1_05_in30 = reg_0419;
    76: op1_05_in30 = reg_0110;
    77: op1_05_in30 = reg_0830;
    78: op1_05_in30 = reg_0090;
    79: op1_05_in30 = imem06_in[87:84];
    80: op1_05_in30 = reg_0567;
    82: op1_05_in30 = reg_0421;
    83: op1_05_in30 = reg_0300;
    84: op1_05_in30 = reg_0500;
    85: op1_05_in30 = reg_0804;
    87: op1_05_in30 = imem04_in[43:40];
    88: op1_05_in30 = reg_0950;
    89: op1_05_in30 = imem02_in[115:112];
    90: op1_05_in30 = reg_0169;
    91: op1_05_in30 = reg_0247;
    92: op1_05_in30 = reg_0569;
    93: op1_05_in30 = reg_0832;
    95: op1_05_in30 = reg_1034;
    96: op1_05_in30 = reg_0225;
    default: op1_05_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_05_inv30 = 1;
    16: op1_05_inv30 = 1;
    18: op1_05_inv30 = 1;
    20: op1_05_inv30 = 1;
    21: op1_05_inv30 = 1;
    23: op1_05_inv30 = 1;
    25: op1_05_inv30 = 1;
    26: op1_05_inv30 = 1;
    27: op1_05_inv30 = 1;
    29: op1_05_inv30 = 1;
    30: op1_05_inv30 = 1;
    31: op1_05_inv30 = 1;
    33: op1_05_inv30 = 1;
    36: op1_05_inv30 = 1;
    42: op1_05_inv30 = 1;
    44: op1_05_inv30 = 1;
    45: op1_05_inv30 = 1;
    48: op1_05_inv30 = 1;
    49: op1_05_inv30 = 1;
    51: op1_05_inv30 = 1;
    52: op1_05_inv30 = 1;
    53: op1_05_inv30 = 1;
    55: op1_05_inv30 = 1;
    59: op1_05_inv30 = 1;
    62: op1_05_inv30 = 1;
    63: op1_05_inv30 = 1;
    67: op1_05_inv30 = 1;
    69: op1_05_inv30 = 1;
    70: op1_05_inv30 = 1;
    72: op1_05_inv30 = 1;
    74: op1_05_inv30 = 1;
    77: op1_05_inv30 = 1;
    80: op1_05_inv30 = 1;
    83: op1_05_inv30 = 1;
    87: op1_05_inv30 = 1;
    90: op1_05_inv30 = 1;
    94: op1_05_inv30 = 1;
    95: op1_05_inv30 = 1;
    default: op1_05_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_05_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_05_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in00 = reg_0121;
    6: op1_06_in00 = imem00_in[55:52];
    7: op1_06_in00 = reg_0991;
    8: op1_06_in00 = reg_0033;
    9: op1_06_in00 = reg_0112;
    10: op1_06_in00 = imem00_in[3:0];
    37: op1_06_in00 = imem00_in[3:0];
    43: op1_06_in00 = imem00_in[3:0];
    11: op1_06_in00 = reg_1037;
    84: op1_06_in00 = reg_1037;
    12: op1_06_in00 = imem00_in[23:20];
    4: op1_06_in00 = imem07_in[23:20];
    66: op1_06_in00 = imem07_in[23:20];
    13: op1_06_in00 = reg_0283;
    14: op1_06_in00 = reg_0753;
    15: op1_06_in00 = imem00_in[35:32];
    16: op1_06_in00 = reg_0585;
    17: op1_06_in00 = reg_0071;
    18: op1_06_in00 = imem02_in[95:92];
    19: op1_06_in00 = imem06_in[19:16];
    3: op1_06_in00 = imem07_in[47:44];
    20: op1_06_in00 = reg_0119;
    52: op1_06_in00 = reg_0119;
    21: op1_06_in00 = reg_0825;
    22: op1_06_in00 = reg_1045;
    23: op1_06_in00 = reg_0249;
    24: op1_06_in00 = reg_0694;
    25: op1_06_in00 = reg_0578;
    2: op1_06_in00 = imem07_in[115:112];
    26: op1_06_in00 = reg_0900;
    27: op1_06_in00 = reg_0592;
    28: op1_06_in00 = reg_0537;
    29: op1_06_in00 = reg_0496;
    30: op1_06_in00 = imem02_in[7:4];
    31: op1_06_in00 = reg_0053;
    83: op1_06_in00 = reg_0053;
    32: op1_06_in00 = imem00_in[7:4];
    35: op1_06_in00 = imem00_in[7:4];
    68: op1_06_in00 = imem00_in[7:4];
    86: op1_06_in00 = imem00_in[7:4];
    97: op1_06_in00 = imem00_in[7:4];
    33: op1_06_in00 = reg_0810;
    34: op1_06_in00 = reg_0543;
    36: op1_06_in00 = reg_0184;
    38: op1_06_in00 = imem00_in[11:8];
    39: op1_06_in00 = reg_1044;
    40: op1_06_in00 = reg_0992;
    41: op1_06_in00 = reg_0660;
    42: op1_06_in00 = reg_0894;
    44: op1_06_in00 = imem02_in[83:80];
    45: op1_06_in00 = imem05_in[51:48];
    46: op1_06_in00 = imem07_in[71:68];
    47: op1_06_in00 = reg_0219;
    48: op1_06_in00 = imem04_in[127:124];
    49: op1_06_in00 = reg_0419;
    50: op1_06_in00 = reg_0142;
    51: op1_06_in00 = reg_0313;
    53: op1_06_in00 = reg_0996;
    54: op1_06_in00 = reg_0850;
    55: op1_06_in00 = imem06_in[83:80];
    56: op1_06_in00 = reg_0533;
    57: op1_06_in00 = reg_0161;
    58: op1_06_in00 = imem00_in[15:12];
    59: op1_06_in00 = imem07_in[59:56];
    60: op1_06_in00 = reg_0904;
    61: op1_06_in00 = imem00_in[83:80];
    62: op1_06_in00 = reg_0304;
    63: op1_06_in00 = imem05_in[79:76];
    64: op1_06_in00 = reg_0447;
    65: op1_06_in00 = reg_0713;
    67: op1_06_in00 = reg_0241;
    69: op1_06_in00 = reg_0513;
    70: op1_06_in00 = reg_0143;
    71: op1_06_in00 = imem00_in[19:16];
    72: op1_06_in00 = reg_0147;
    73: op1_06_in00 = imem07_in[3:0];
    74: op1_06_in00 = reg_0641;
    75: op1_06_in00 = imem00_in[43:40];
    76: op1_06_in00 = imem02_in[23:20];
    77: op1_06_in00 = reg_0906;
    78: op1_06_in00 = reg_0091;
    79: op1_06_in00 = imem06_in[91:88];
    80: op1_06_in00 = reg_0569;
    81: op1_06_in00 = imem00_in[27:24];
    82: op1_06_in00 = reg_0315;
    85: op1_06_in00 = reg_0699;
    87: op1_06_in00 = imem04_in[47:44];
    88: op1_06_in00 = reg_0945;
    89: op1_06_in00 = imem02_in[127:124];
    90: op1_06_in00 = reg_0914;
    91: op1_06_in00 = reg_0718;
    92: op1_06_in00 = reg_0164;
    93: op1_06_in00 = reg_0512;
    94: op1_06_in00 = reg_1031;
    95: op1_06_in00 = imem01_in[7:4];
    96: op1_06_in00 = reg_1051;
    default: op1_06_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv00 = 1;
    6: op1_06_inv00 = 1;
    7: op1_06_inv00 = 1;
    9: op1_06_inv00 = 1;
    11: op1_06_inv00 = 1;
    15: op1_06_inv00 = 1;
    17: op1_06_inv00 = 1;
    18: op1_06_inv00 = 1;
    21: op1_06_inv00 = 1;
    24: op1_06_inv00 = 1;
    2: op1_06_inv00 = 1;
    26: op1_06_inv00 = 1;
    28: op1_06_inv00 = 1;
    29: op1_06_inv00 = 1;
    31: op1_06_inv00 = 1;
    33: op1_06_inv00 = 1;
    35: op1_06_inv00 = 1;
    38: op1_06_inv00 = 1;
    39: op1_06_inv00 = 1;
    41: op1_06_inv00 = 1;
    42: op1_06_inv00 = 1;
    44: op1_06_inv00 = 1;
    46: op1_06_inv00 = 1;
    47: op1_06_inv00 = 1;
    49: op1_06_inv00 = 1;
    51: op1_06_inv00 = 1;
    52: op1_06_inv00 = 1;
    53: op1_06_inv00 = 1;
    54: op1_06_inv00 = 1;
    58: op1_06_inv00 = 1;
    59: op1_06_inv00 = 1;
    61: op1_06_inv00 = 1;
    63: op1_06_inv00 = 1;
    67: op1_06_inv00 = 1;
    68: op1_06_inv00 = 1;
    69: op1_06_inv00 = 1;
    72: op1_06_inv00 = 1;
    74: op1_06_inv00 = 1;
    75: op1_06_inv00 = 1;
    77: op1_06_inv00 = 1;
    78: op1_06_inv00 = 1;
    80: op1_06_inv00 = 1;
    81: op1_06_inv00 = 1;
    82: op1_06_inv00 = 1;
    87: op1_06_inv00 = 1;
    88: op1_06_inv00 = 1;
    89: op1_06_inv00 = 1;
    91: op1_06_inv00 = 1;
    94: op1_06_inv00 = 1;
    96: op1_06_inv00 = 1;
    97: op1_06_inv00 = 1;
    default: op1_06_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in01 = reg_0110;
    6: op1_06_in01 = imem00_in[75:72];
    7: op1_06_in01 = reg_0995;
    8: op1_06_in01 = reg_0028;
    9: op1_06_in01 = reg_0113;
    10: op1_06_in01 = imem00_in[23:20];
    35: op1_06_in01 = imem00_in[23:20];
    71: op1_06_in01 = imem00_in[23:20];
    11: op1_06_in01 = reg_0227;
    12: op1_06_in01 = imem00_in[43:40];
    97: op1_06_in01 = imem00_in[43:40];
    4: op1_06_in01 = imem07_in[39:36];
    13: op1_06_in01 = reg_0300;
    14: op1_06_in01 = reg_0781;
    56: op1_06_in01 = reg_0781;
    15: op1_06_in01 = imem00_in[39:36];
    43: op1_06_in01 = imem00_in[39:36];
    16: op1_06_in01 = reg_0600;
    17: op1_06_in01 = imem05_in[3:0];
    18: op1_06_in01 = reg_0653;
    80: op1_06_in01 = reg_0653;
    19: op1_06_in01 = imem06_in[43:40];
    3: op1_06_in01 = imem07_in[71:68];
    20: op1_06_in01 = reg_0112;
    21: op1_06_in01 = reg_0244;
    22: op1_06_in01 = reg_1041;
    23: op1_06_in01 = reg_1033;
    24: op1_06_in01 = reg_0676;
    25: op1_06_in01 = reg_0597;
    26: op1_06_in01 = reg_0827;
    27: op1_06_in01 = reg_0589;
    28: op1_06_in01 = reg_0313;
    29: op1_06_in01 = reg_0871;
    30: op1_06_in01 = imem02_in[67:64];
    31: op1_06_in01 = reg_0285;
    32: op1_06_in01 = imem00_in[31:28];
    58: op1_06_in01 = imem00_in[31:28];
    33: op1_06_in01 = reg_0247;
    34: op1_06_in01 = reg_0795;
    37: op1_06_in01 = imem00_in[55:52];
    38: op1_06_in01 = imem00_in[59:56];
    39: op1_06_in01 = reg_1040;
    40: op1_06_in01 = reg_0979;
    41: op1_06_in01 = reg_0639;
    42: op1_06_in01 = reg_0630;
    44: op1_06_in01 = imem02_in[87:84];
    45: op1_06_in01 = imem05_in[63:60];
    46: op1_06_in01 = imem07_in[99:96];
    47: op1_06_in01 = reg_0496;
    48: op1_06_in01 = reg_0055;
    49: op1_06_in01 = reg_0180;
    50: op1_06_in01 = reg_0140;
    51: op1_06_in01 = reg_0568;
    52: op1_06_in01 = reg_0127;
    53: op1_06_in01 = reg_1001;
    54: op1_06_in01 = reg_0281;
    55: op1_06_in01 = imem06_in[99:96];
    57: op1_06_in01 = reg_0167;
    59: op1_06_in01 = imem07_in[63:60];
    60: op1_06_in01 = reg_1036;
    61: op1_06_in01 = imem00_in[87:84];
    62: op1_06_in01 = reg_0512;
    96: op1_06_in01 = reg_0512;
    63: op1_06_in01 = imem05_in[111:108];
    64: op1_06_in01 = reg_0819;
    65: op1_06_in01 = reg_0707;
    66: op1_06_in01 = imem07_in[43:40];
    67: op1_06_in01 = reg_0605;
    68: op1_06_in01 = imem00_in[47:44];
    69: op1_06_in01 = reg_0844;
    70: op1_06_in01 = reg_0137;
    72: op1_06_in01 = reg_0149;
    73: op1_06_in01 = imem07_in[27:24];
    74: op1_06_in01 = reg_0599;
    75: op1_06_in01 = imem00_in[123:120];
    76: op1_06_in01 = imem02_in[99:96];
    77: op1_06_in01 = reg_0733;
    78: op1_06_in01 = reg_0049;
    79: op1_06_in01 = imem06_in[95:92];
    81: op1_06_in01 = reg_0682;
    82: op1_06_in01 = reg_0532;
    83: op1_06_in01 = reg_0774;
    84: op1_06_in01 = reg_1031;
    85: op1_06_in01 = reg_0632;
    86: op1_06_in01 = imem00_in[11:8];
    87: op1_06_in01 = imem04_in[75:72];
    88: op1_06_in01 = reg_0965;
    89: op1_06_in01 = reg_0305;
    90: op1_06_in01 = reg_0034;
    91: op1_06_in01 = reg_0299;
    92: op1_06_in01 = reg_0959;
    93: op1_06_in01 = reg_1053;
    94: op1_06_in01 = reg_1045;
    95: op1_06_in01 = imem01_in[11:8];
    default: op1_06_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv01 = 1;
    6: op1_06_inv01 = 1;
    10: op1_06_inv01 = 1;
    14: op1_06_inv01 = 1;
    16: op1_06_inv01 = 1;
    17: op1_06_inv01 = 1;
    19: op1_06_inv01 = 1;
    20: op1_06_inv01 = 1;
    22: op1_06_inv01 = 1;
    25: op1_06_inv01 = 1;
    28: op1_06_inv01 = 1;
    29: op1_06_inv01 = 1;
    32: op1_06_inv01 = 1;
    33: op1_06_inv01 = 1;
    38: op1_06_inv01 = 1;
    39: op1_06_inv01 = 1;
    40: op1_06_inv01 = 1;
    46: op1_06_inv01 = 1;
    50: op1_06_inv01 = 1;
    52: op1_06_inv01 = 1;
    53: op1_06_inv01 = 1;
    54: op1_06_inv01 = 1;
    56: op1_06_inv01 = 1;
    57: op1_06_inv01 = 1;
    58: op1_06_inv01 = 1;
    59: op1_06_inv01 = 1;
    62: op1_06_inv01 = 1;
    63: op1_06_inv01 = 1;
    64: op1_06_inv01 = 1;
    67: op1_06_inv01 = 1;
    72: op1_06_inv01 = 1;
    75: op1_06_inv01 = 1;
    78: op1_06_inv01 = 1;
    81: op1_06_inv01 = 1;
    84: op1_06_inv01 = 1;
    85: op1_06_inv01 = 1;
    88: op1_06_inv01 = 1;
    91: op1_06_inv01 = 1;
    92: op1_06_inv01 = 1;
    94: op1_06_inv01 = 1;
    95: op1_06_inv01 = 1;
    default: op1_06_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in02 = imem02_in[3:0];
    6: op1_06_in02 = imem00_in[123:120];
    7: op1_06_in02 = reg_0986;
    8: op1_06_in02 = reg_0039;
    9: op1_06_in02 = imem02_in[23:20];
    10: op1_06_in02 = imem00_in[27:24];
    11: op1_06_in02 = reg_1036;
    12: op1_06_in02 = imem00_in[75:72];
    4: op1_06_in02 = imem07_in[83:80];
    13: op1_06_in02 = reg_0299;
    92: op1_06_in02 = reg_0299;
    14: op1_06_in02 = reg_0783;
    15: op1_06_in02 = imem00_in[83:80];
    16: op1_06_in02 = reg_0576;
    17: op1_06_in02 = imem05_in[15:12];
    31: op1_06_in02 = imem05_in[15:12];
    18: op1_06_in02 = reg_0662;
    19: op1_06_in02 = imem06_in[67:64];
    3: op1_06_in02 = imem07_in[87:84];
    20: op1_06_in02 = imem02_in[75:72];
    21: op1_06_in02 = reg_0896;
    22: op1_06_in02 = reg_1038;
    23: op1_06_in02 = reg_1038;
    24: op1_06_in02 = reg_0677;
    25: op1_06_in02 = reg_0581;
    26: op1_06_in02 = reg_0785;
    27: op1_06_in02 = reg_0580;
    28: op1_06_in02 = reg_0740;
    29: op1_06_in02 = reg_0123;
    30: op1_06_in02 = imem02_in[123:120];
    76: op1_06_in02 = imem02_in[123:120];
    32: op1_06_in02 = imem00_in[55:52];
    68: op1_06_in02 = imem00_in[55:52];
    71: op1_06_in02 = imem00_in[55:52];
    33: op1_06_in02 = reg_0544;
    34: op1_06_in02 = reg_0373;
    35: op1_06_in02 = imem00_in[35:32];
    37: op1_06_in02 = imem00_in[67:64];
    97: op1_06_in02 = imem00_in[67:64];
    38: op1_06_in02 = imem00_in[63:60];
    58: op1_06_in02 = imem00_in[63:60];
    39: op1_06_in02 = reg_1041;
    40: op1_06_in02 = reg_0999;
    53: op1_06_in02 = reg_0999;
    41: op1_06_in02 = reg_0652;
    42: op1_06_in02 = reg_0241;
    43: op1_06_in02 = imem00_in[99:96];
    44: op1_06_in02 = imem02_in[119:116];
    45: op1_06_in02 = reg_0970;
    46: op1_06_in02 = reg_0726;
    47: op1_06_in02 = reg_0216;
    48: op1_06_in02 = reg_0932;
    49: op1_06_in02 = reg_0182;
    50: op1_06_in02 = imem06_in[11:8];
    51: op1_06_in02 = reg_0015;
    52: op1_06_in02 = reg_0126;
    54: op1_06_in02 = reg_0756;
    55: op1_06_in02 = reg_0613;
    56: op1_06_in02 = reg_0619;
    57: op1_06_in02 = reg_0183;
    59: op1_06_in02 = reg_0704;
    60: op1_06_in02 = reg_1045;
    61: op1_06_in02 = reg_0825;
    62: op1_06_in02 = reg_0003;
    63: op1_06_in02 = reg_0835;
    64: op1_06_in02 = reg_0438;
    65: op1_06_in02 = reg_0706;
    66: op1_06_in02 = imem07_in[59:56];
    67: op1_06_in02 = reg_1010;
    69: op1_06_in02 = reg_0822;
    70: op1_06_in02 = reg_0134;
    72: op1_06_in02 = reg_0146;
    73: op1_06_in02 = imem07_in[43:40];
    74: op1_06_in02 = reg_0868;
    75: op1_06_in02 = reg_0001;
    77: op1_06_in02 = reg_0113;
    78: op1_06_in02 = imem03_in[11:8];
    79: op1_06_in02 = imem06_in[103:100];
    80: op1_06_in02 = reg_0002;
    81: op1_06_in02 = reg_0683;
    82: op1_06_in02 = reg_0431;
    83: op1_06_in02 = reg_0656;
    84: op1_06_in02 = reg_0610;
    85: op1_06_in02 = reg_0917;
    86: op1_06_in02 = imem00_in[19:16];
    87: op1_06_in02 = imem04_in[119:116];
    88: op1_06_in02 = imem06_in[47:44];
    89: op1_06_in02 = reg_0639;
    90: op1_06_in02 = reg_0124;
    91: op1_06_in02 = reg_0805;
    93: op1_06_in02 = reg_0273;
    94: op1_06_in02 = reg_0294;
    95: op1_06_in02 = imem01_in[47:44];
    96: op1_06_in02 = reg_0860;
    default: op1_06_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv02 = 1;
    6: op1_06_inv02 = 1;
    7: op1_06_inv02 = 1;
    8: op1_06_inv02 = 1;
    9: op1_06_inv02 = 1;
    12: op1_06_inv02 = 1;
    15: op1_06_inv02 = 1;
    17: op1_06_inv02 = 1;
    18: op1_06_inv02 = 1;
    19: op1_06_inv02 = 1;
    3: op1_06_inv02 = 1;
    21: op1_06_inv02 = 1;
    22: op1_06_inv02 = 1;
    24: op1_06_inv02 = 1;
    25: op1_06_inv02 = 1;
    26: op1_06_inv02 = 1;
    27: op1_06_inv02 = 1;
    28: op1_06_inv02 = 1;
    30: op1_06_inv02 = 1;
    35: op1_06_inv02 = 1;
    38: op1_06_inv02 = 1;
    39: op1_06_inv02 = 1;
    40: op1_06_inv02 = 1;
    41: op1_06_inv02 = 1;
    42: op1_06_inv02 = 1;
    43: op1_06_inv02 = 1;
    44: op1_06_inv02 = 1;
    45: op1_06_inv02 = 1;
    46: op1_06_inv02 = 1;
    47: op1_06_inv02 = 1;
    49: op1_06_inv02 = 1;
    50: op1_06_inv02 = 1;
    52: op1_06_inv02 = 1;
    53: op1_06_inv02 = 1;
    55: op1_06_inv02 = 1;
    56: op1_06_inv02 = 1;
    60: op1_06_inv02 = 1;
    61: op1_06_inv02 = 1;
    64: op1_06_inv02 = 1;
    67: op1_06_inv02 = 1;
    69: op1_06_inv02 = 1;
    70: op1_06_inv02 = 1;
    72: op1_06_inv02 = 1;
    73: op1_06_inv02 = 1;
    74: op1_06_inv02 = 1;
    75: op1_06_inv02 = 1;
    76: op1_06_inv02 = 1;
    77: op1_06_inv02 = 1;
    81: op1_06_inv02 = 1;
    82: op1_06_inv02 = 1;
    83: op1_06_inv02 = 1;
    84: op1_06_inv02 = 1;
    87: op1_06_inv02 = 1;
    91: op1_06_inv02 = 1;
    95: op1_06_inv02 = 1;
    97: op1_06_inv02 = 1;
    default: op1_06_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in03 = imem02_in[7:4];
    6: op1_06_in03 = reg_0681;
    7: op1_06_in03 = reg_0981;
    53: op1_06_in03 = reg_0981;
    8: op1_06_in03 = reg_0031;
    9: op1_06_in03 = imem02_in[31:28];
    10: op1_06_in03 = imem00_in[31:28];
    11: op1_06_in03 = reg_1015;
    12: op1_06_in03 = imem00_in[103:100];
    4: op1_06_in03 = imem07_in[99:96];
    13: op1_06_in03 = reg_0302;
    14: op1_06_in03 = reg_0005;
    15: op1_06_in03 = imem00_in[107:104];
    16: op1_06_in03 = reg_0395;
    17: op1_06_in03 = imem05_in[19:16];
    18: op1_06_in03 = reg_0352;
    19: op1_06_in03 = imem06_in[99:96];
    3: op1_06_in03 = imem07_in[91:88];
    20: op1_06_in03 = imem02_in[115:112];
    21: op1_06_in03 = reg_0489;
    22: op1_06_in03 = reg_0107;
    23: op1_06_in03 = reg_0123;
    24: op1_06_in03 = reg_0680;
    61: op1_06_in03 = reg_0680;
    25: op1_06_in03 = reg_0595;
    56: op1_06_in03 = reg_0595;
    26: op1_06_in03 = reg_0896;
    27: op1_06_in03 = reg_0590;
    28: op1_06_in03 = reg_0075;
    29: op1_06_in03 = reg_0100;
    30: op1_06_in03 = imem02_in[127:124];
    44: op1_06_in03 = imem02_in[127:124];
    31: op1_06_in03 = imem05_in[59:56];
    32: op1_06_in03 = imem00_in[79:76];
    33: op1_06_in03 = reg_0769;
    34: op1_06_in03 = reg_0377;
    35: op1_06_in03 = imem00_in[39:36];
    37: op1_06_in03 = imem00_in[95:92];
    38: op1_06_in03 = imem00_in[67:64];
    58: op1_06_in03 = imem00_in[67:64];
    39: op1_06_in03 = reg_1038;
    40: op1_06_in03 = reg_0988;
    41: op1_06_in03 = reg_0667;
    42: op1_06_in03 = reg_0596;
    43: op1_06_in03 = imem00_in[123:120];
    45: op1_06_in03 = reg_0955;
    46: op1_06_in03 = reg_0703;
    47: op1_06_in03 = reg_1040;
    48: op1_06_in03 = reg_0584;
    49: op1_06_in03 = reg_0177;
    50: op1_06_in03 = imem06_in[55:52];
    51: op1_06_in03 = reg_0074;
    52: op1_06_in03 = reg_0314;
    54: op1_06_in03 = reg_0578;
    55: op1_06_in03 = reg_0624;
    57: op1_06_in03 = reg_0164;
    59: op1_06_in03 = reg_0724;
    60: op1_06_in03 = reg_0487;
    62: op1_06_in03 = reg_0116;
    63: op1_06_in03 = reg_0969;
    64: op1_06_in03 = reg_0133;
    65: op1_06_in03 = reg_0361;
    66: op1_06_in03 = imem07_in[79:76];
    67: op1_06_in03 = reg_0633;
    83: op1_06_in03 = reg_0633;
    68: op1_06_in03 = reg_0843;
    69: op1_06_in03 = reg_0993;
    70: op1_06_in03 = imem06_in[7:4];
    71: op1_06_in03 = imem00_in[63:60];
    72: op1_06_in03 = imem06_in[91:88];
    73: op1_06_in03 = imem07_in[59:56];
    74: op1_06_in03 = reg_0173;
    75: op1_06_in03 = reg_0825;
    76: op1_06_in03 = reg_0803;
    77: op1_06_in03 = imem02_in[23:20];
    78: op1_06_in03 = imem03_in[127:124];
    79: op1_06_in03 = imem06_in[115:112];
    80: op1_06_in03 = reg_0250;
    81: op1_06_in03 = reg_0768;
    82: op1_06_in03 = imem07_in[3:0];
    84: op1_06_in03 = reg_0111;
    85: op1_06_in03 = reg_0289;
    86: op1_06_in03 = imem00_in[35:32];
    87: op1_06_in03 = imem04_in[123:120];
    88: op1_06_in03 = imem06_in[59:56];
    89: op1_06_in03 = reg_0091;
    90: op1_06_in03 = reg_0782;
    91: op1_06_in03 = reg_0575;
    92: op1_06_in03 = reg_0805;
    93: op1_06_in03 = reg_0827;
    94: op1_06_in03 = reg_0832;
    95: op1_06_in03 = imem01_in[51:48];
    96: op1_06_in03 = reg_0103;
    97: op1_06_in03 = imem00_in[75:72];
    default: op1_06_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv03 = 1;
    7: op1_06_inv03 = 1;
    9: op1_06_inv03 = 1;
    10: op1_06_inv03 = 1;
    11: op1_06_inv03 = 1;
    12: op1_06_inv03 = 1;
    13: op1_06_inv03 = 1;
    15: op1_06_inv03 = 1;
    18: op1_06_inv03 = 1;
    20: op1_06_inv03 = 1;
    21: op1_06_inv03 = 1;
    23: op1_06_inv03 = 1;
    24: op1_06_inv03 = 1;
    26: op1_06_inv03 = 1;
    30: op1_06_inv03 = 1;
    31: op1_06_inv03 = 1;
    34: op1_06_inv03 = 1;
    35: op1_06_inv03 = 1;
    39: op1_06_inv03 = 1;
    40: op1_06_inv03 = 1;
    41: op1_06_inv03 = 1;
    42: op1_06_inv03 = 1;
    47: op1_06_inv03 = 1;
    48: op1_06_inv03 = 1;
    51: op1_06_inv03 = 1;
    54: op1_06_inv03 = 1;
    55: op1_06_inv03 = 1;
    57: op1_06_inv03 = 1;
    59: op1_06_inv03 = 1;
    61: op1_06_inv03 = 1;
    62: op1_06_inv03 = 1;
    67: op1_06_inv03 = 1;
    69: op1_06_inv03 = 1;
    70: op1_06_inv03 = 1;
    72: op1_06_inv03 = 1;
    73: op1_06_inv03 = 1;
    75: op1_06_inv03 = 1;
    80: op1_06_inv03 = 1;
    82: op1_06_inv03 = 1;
    84: op1_06_inv03 = 1;
    90: op1_06_inv03 = 1;
    92: op1_06_inv03 = 1;
    94: op1_06_inv03 = 1;
    default: op1_06_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in04 = imem02_in[47:44];
    6: op1_06_in04 = reg_0686;
    68: op1_06_in04 = reg_0686;
    7: op1_06_in04 = imem04_in[11:8];
    8: op1_06_in04 = reg_0034;
    9: op1_06_in04 = imem02_in[51:48];
    10: op1_06_in04 = imem00_in[35:32];
    11: op1_06_in04 = reg_1041;
    12: op1_06_in04 = reg_0697;
    4: op1_06_in04 = reg_0424;
    13: op1_06_in04 = reg_0298;
    14: op1_06_in04 = imem07_in[15:12];
    15: op1_06_in04 = reg_0693;
    43: op1_06_in04 = reg_0693;
    16: op1_06_in04 = reg_0376;
    34: op1_06_in04 = reg_0376;
    17: op1_06_in04 = imem05_in[27:24];
    18: op1_06_in04 = reg_0357;
    19: op1_06_in04 = imem06_in[103:100];
    3: op1_06_in04 = imem07_in[107:104];
    20: op1_06_in04 = reg_0650;
    21: op1_06_in04 = reg_0149;
    22: op1_06_in04 = reg_0117;
    23: op1_06_in04 = reg_0103;
    24: op1_06_in04 = reg_0453;
    25: op1_06_in04 = reg_0590;
    26: op1_06_in04 = reg_0147;
    27: op1_06_in04 = reg_0395;
    56: op1_06_in04 = reg_0395;
    28: op1_06_in04 = reg_0070;
    29: op1_06_in04 = imem02_in[3:0];
    30: op1_06_in04 = reg_0658;
    31: op1_06_in04 = imem05_in[79:76];
    32: op1_06_in04 = imem00_in[111:108];
    97: op1_06_in04 = imem00_in[111:108];
    33: op1_06_in04 = reg_0905;
    35: op1_06_in04 = imem00_in[43:40];
    37: op1_06_in04 = imem00_in[107:104];
    38: op1_06_in04 = imem00_in[115:112];
    39: op1_06_in04 = reg_0104;
    40: op1_06_in04 = imem04_in[7:4];
    69: op1_06_in04 = imem04_in[7:4];
    41: op1_06_in04 = reg_0045;
    42: op1_06_in04 = reg_1010;
    44: op1_06_in04 = reg_0660;
    45: op1_06_in04 = reg_0948;
    46: op1_06_in04 = reg_0729;
    47: op1_06_in04 = reg_0616;
    48: op1_06_in04 = reg_0401;
    50: op1_06_in04 = imem06_in[67:64];
    51: op1_06_in04 = reg_0748;
    52: op1_06_in04 = reg_0566;
    53: op1_06_in04 = imem04_in[99:96];
    54: op1_06_in04 = reg_0864;
    55: op1_06_in04 = reg_0020;
    57: op1_06_in04 = reg_0168;
    58: op1_06_in04 = imem00_in[99:96];
    59: op1_06_in04 = reg_0709;
    60: op1_06_in04 = reg_1039;
    61: op1_06_in04 = reg_0454;
    62: op1_06_in04 = reg_0283;
    63: op1_06_in04 = reg_0949;
    64: op1_06_in04 = reg_0152;
    65: op1_06_in04 = reg_0325;
    66: op1_06_in04 = imem07_in[95:92];
    67: op1_06_in04 = imem07_in[75:72];
    70: op1_06_in04 = imem06_in[39:36];
    71: op1_06_in04 = imem00_in[67:64];
    72: op1_06_in04 = imem06_in[107:104];
    73: op1_06_in04 = imem07_in[63:60];
    74: op1_06_in04 = reg_0171;
    75: op1_06_in04 = reg_0842;
    76: op1_06_in04 = reg_0813;
    77: op1_06_in04 = imem02_in[59:56];
    78: op1_06_in04 = reg_1007;
    79: op1_06_in04 = reg_0625;
    80: op1_06_in04 = reg_0641;
    81: op1_06_in04 = reg_0825;
    82: op1_06_in04 = imem07_in[23:20];
    83: op1_06_in04 = reg_0932;
    84: op1_06_in04 = reg_0116;
    85: op1_06_in04 = reg_0807;
    86: op1_06_in04 = imem00_in[127:124];
    87: op1_06_in04 = reg_0405;
    88: op1_06_in04 = imem06_in[75:72];
    89: op1_06_in04 = reg_0621;
    90: op1_06_in04 = reg_0222;
    91: op1_06_in04 = reg_0002;
    92: op1_06_in04 = reg_0422;
    93: op1_06_in04 = imem02_in[11:8];
    94: op1_06_in04 = reg_1051;
    95: op1_06_in04 = imem01_in[63:60];
    96: op1_06_in04 = reg_0821;
    default: op1_06_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv04 = 1;
    8: op1_06_inv04 = 1;
    9: op1_06_inv04 = 1;
    11: op1_06_inv04 = 1;
    14: op1_06_inv04 = 1;
    15: op1_06_inv04 = 1;
    17: op1_06_inv04 = 1;
    20: op1_06_inv04 = 1;
    21: op1_06_inv04 = 1;
    24: op1_06_inv04 = 1;
    26: op1_06_inv04 = 1;
    29: op1_06_inv04 = 1;
    31: op1_06_inv04 = 1;
    32: op1_06_inv04 = 1;
    33: op1_06_inv04 = 1;
    34: op1_06_inv04 = 1;
    37: op1_06_inv04 = 1;
    38: op1_06_inv04 = 1;
    40: op1_06_inv04 = 1;
    41: op1_06_inv04 = 1;
    42: op1_06_inv04 = 1;
    43: op1_06_inv04 = 1;
    44: op1_06_inv04 = 1;
    50: op1_06_inv04 = 1;
    51: op1_06_inv04 = 1;
    56: op1_06_inv04 = 1;
    57: op1_06_inv04 = 1;
    58: op1_06_inv04 = 1;
    59: op1_06_inv04 = 1;
    60: op1_06_inv04 = 1;
    61: op1_06_inv04 = 1;
    62: op1_06_inv04 = 1;
    63: op1_06_inv04 = 1;
    64: op1_06_inv04 = 1;
    67: op1_06_inv04 = 1;
    69: op1_06_inv04 = 1;
    70: op1_06_inv04 = 1;
    72: op1_06_inv04 = 1;
    73: op1_06_inv04 = 1;
    75: op1_06_inv04 = 1;
    76: op1_06_inv04 = 1;
    77: op1_06_inv04 = 1;
    78: op1_06_inv04 = 1;
    81: op1_06_inv04 = 1;
    82: op1_06_inv04 = 1;
    83: op1_06_inv04 = 1;
    84: op1_06_inv04 = 1;
    85: op1_06_inv04 = 1;
    88: op1_06_inv04 = 1;
    89: op1_06_inv04 = 1;
    90: op1_06_inv04 = 1;
    92: op1_06_inv04 = 1;
    94: op1_06_inv04 = 1;
    default: op1_06_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in05 = imem02_in[71:68];
    9: op1_06_in05 = imem02_in[71:68];
    6: op1_06_in05 = reg_0691;
    7: op1_06_in05 = imem04_in[87:84];
    8: op1_06_in05 = reg_0035;
    10: op1_06_in05 = imem00_in[39:36];
    11: op1_06_in05 = reg_0228;
    12: op1_06_in05 = reg_0686;
    32: op1_06_in05 = reg_0686;
    4: op1_06_in05 = reg_0428;
    13: op1_06_in05 = reg_0278;
    14: op1_06_in05 = imem07_in[51:48];
    15: op1_06_in05 = reg_0683;
    16: op1_06_in05 = reg_0309;
    17: op1_06_in05 = imem05_in[51:48];
    18: op1_06_in05 = reg_0345;
    19: op1_06_in05 = imem06_in[111:108];
    3: op1_06_in05 = imem07_in[123:120];
    66: op1_06_in05 = imem07_in[123:120];
    67: op1_06_in05 = imem07_in[123:120];
    20: op1_06_in05 = reg_0655;
    21: op1_06_in05 = reg_0145;
    22: op1_06_in05 = reg_0113;
    23: op1_06_in05 = reg_0100;
    24: op1_06_in05 = reg_0476;
    25: op1_06_in05 = reg_0391;
    26: op1_06_in05 = reg_0135;
    27: op1_06_in05 = reg_0384;
    28: op1_06_in05 = reg_0047;
    29: op1_06_in05 = imem02_in[27:24];
    30: op1_06_in05 = reg_0640;
    31: op1_06_in05 = imem05_in[107:104];
    33: op1_06_in05 = reg_1042;
    34: op1_06_in05 = reg_0234;
    35: op1_06_in05 = imem00_in[51:48];
    37: op1_06_in05 = imem00_in[119:116];
    38: op1_06_in05 = imem00_in[119:116];
    39: op1_06_in05 = reg_0099;
    40: op1_06_in05 = imem04_in[31:28];
    41: op1_06_in05 = reg_0039;
    42: op1_06_in05 = reg_0531;
    43: op1_06_in05 = reg_0676;
    44: op1_06_in05 = reg_0662;
    45: op1_06_in05 = reg_0950;
    46: op1_06_in05 = reg_0718;
    47: op1_06_in05 = reg_0119;
    48: op1_06_in05 = reg_0015;
    50: op1_06_in05 = imem06_in[75:72];
    51: op1_06_in05 = reg_0444;
    52: op1_06_in05 = reg_0547;
    53: op1_06_in05 = imem04_in[111:108];
    54: op1_06_in05 = reg_0031;
    55: op1_06_in05 = reg_0781;
    56: op1_06_in05 = reg_0392;
    57: op1_06_in05 = reg_0170;
    58: op1_06_in05 = imem00_in[103:100];
    59: op1_06_in05 = reg_0321;
    60: op1_06_in05 = reg_0522;
    61: op1_06_in05 = reg_0450;
    62: op1_06_in05 = reg_1033;
    63: op1_06_in05 = reg_0272;
    64: op1_06_in05 = reg_0156;
    65: op1_06_in05 = reg_0431;
    68: op1_06_in05 = reg_0842;
    69: op1_06_in05 = imem04_in[43:40];
    70: op1_06_in05 = imem06_in[59:56];
    71: op1_06_in05 = imem00_in[75:72];
    72: op1_06_in05 = reg_0021;
    73: op1_06_in05 = imem07_in[71:68];
    75: op1_06_in05 = reg_0668;
    76: op1_06_in05 = reg_0034;
    77: op1_06_in05 = imem02_in[91:88];
    78: op1_06_in05 = reg_0327;
    79: op1_06_in05 = reg_1018;
    80: op1_06_in05 = reg_0420;
    81: op1_06_in05 = reg_0738;
    82: op1_06_in05 = imem07_in[27:24];
    83: op1_06_in05 = imem04_in[75:72];
    84: op1_06_in05 = reg_0283;
    85: op1_06_in05 = reg_0834;
    86: op1_06_in05 = reg_0519;
    87: op1_06_in05 = reg_0446;
    88: op1_06_in05 = imem06_in[83:80];
    89: op1_06_in05 = reg_0642;
    90: op1_06_in05 = reg_0566;
    91: op1_06_in05 = reg_0250;
    92: op1_06_in05 = reg_0744;
    93: op1_06_in05 = imem02_in[35:32];
    94: op1_06_in05 = reg_0555;
    95: op1_06_in05 = imem01_in[87:84];
    96: op1_06_in05 = reg_0745;
    97: op1_06_in05 = reg_0009;
    default: op1_06_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv05 = 1;
    11: op1_06_inv05 = 1;
    15: op1_06_inv05 = 1;
    18: op1_06_inv05 = 1;
    21: op1_06_inv05 = 1;
    22: op1_06_inv05 = 1;
    23: op1_06_inv05 = 1;
    24: op1_06_inv05 = 1;
    25: op1_06_inv05 = 1;
    28: op1_06_inv05 = 1;
    30: op1_06_inv05 = 1;
    32: op1_06_inv05 = 1;
    37: op1_06_inv05 = 1;
    38: op1_06_inv05 = 1;
    41: op1_06_inv05 = 1;
    42: op1_06_inv05 = 1;
    45: op1_06_inv05 = 1;
    46: op1_06_inv05 = 1;
    51: op1_06_inv05 = 1;
    53: op1_06_inv05 = 1;
    54: op1_06_inv05 = 1;
    55: op1_06_inv05 = 1;
    60: op1_06_inv05 = 1;
    62: op1_06_inv05 = 1;
    63: op1_06_inv05 = 1;
    65: op1_06_inv05 = 1;
    66: op1_06_inv05 = 1;
    67: op1_06_inv05 = 1;
    69: op1_06_inv05 = 1;
    71: op1_06_inv05 = 1;
    73: op1_06_inv05 = 1;
    75: op1_06_inv05 = 1;
    79: op1_06_inv05 = 1;
    83: op1_06_inv05 = 1;
    84: op1_06_inv05 = 1;
    85: op1_06_inv05 = 1;
    88: op1_06_inv05 = 1;
    92: op1_06_inv05 = 1;
    95: op1_06_inv05 = 1;
    97: op1_06_inv05 = 1;
    default: op1_06_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in06 = imem02_in[103:100];
    6: op1_06_in06 = reg_0680;
    7: op1_06_in06 = reg_0536;
    8: op1_06_in06 = reg_0040;
    9: op1_06_in06 = imem02_in[107:104];
    77: op1_06_in06 = imem02_in[107:104];
    10: op1_06_in06 = imem00_in[55:52];
    11: op1_06_in06 = reg_0122;
    12: op1_06_in06 = reg_0673;
    4: op1_06_in06 = reg_0434;
    13: op1_06_in06 = reg_0062;
    14: op1_06_in06 = imem07_in[79:76];
    73: op1_06_in06 = imem07_in[79:76];
    15: op1_06_in06 = reg_0685;
    86: op1_06_in06 = reg_0685;
    16: op1_06_in06 = reg_0982;
    17: op1_06_in06 = imem05_in[71:68];
    18: op1_06_in06 = reg_0363;
    19: op1_06_in06 = imem06_in[127:124];
    3: op1_06_in06 = imem07_in[127:124];
    20: op1_06_in06 = reg_0647;
    21: op1_06_in06 = reg_0151;
    22: op1_06_in06 = imem02_in[3:0];
    23: op1_06_in06 = reg_0110;
    24: op1_06_in06 = reg_0475;
    25: op1_06_in06 = reg_0397;
    26: op1_06_in06 = reg_0143;
    27: op1_06_in06 = reg_0388;
    28: op1_06_in06 = reg_0517;
    29: op1_06_in06 = imem02_in[67:64];
    30: op1_06_in06 = reg_0045;
    31: op1_06_in06 = imem05_in[119:116];
    32: op1_06_in06 = reg_0670;
    33: op1_06_in06 = reg_0830;
    60: op1_06_in06 = reg_0830;
    34: op1_06_in06 = reg_1001;
    35: op1_06_in06 = imem00_in[79:76];
    37: op1_06_in06 = imem00_in[123:120];
    38: op1_06_in06 = reg_0697;
    39: op1_06_in06 = reg_0114;
    40: op1_06_in06 = imem04_in[39:36];
    41: op1_06_in06 = reg_0007;
    42: op1_06_in06 = reg_0633;
    43: op1_06_in06 = reg_0679;
    44: op1_06_in06 = reg_0665;
    45: op1_06_in06 = reg_0947;
    46: op1_06_in06 = reg_0701;
    47: op1_06_in06 = reg_0100;
    48: op1_06_in06 = reg_0815;
    50: op1_06_in06 = imem06_in[79:76];
    51: op1_06_in06 = reg_0899;
    52: op1_06_in06 = reg_0667;
    53: op1_06_in06 = reg_0483;
    54: op1_06_in06 = imem05_in[23:20];
    55: op1_06_in06 = reg_0783;
    56: op1_06_in06 = reg_0382;
    57: op1_06_in06 = reg_0171;
    58: op1_06_in06 = reg_0841;
    59: op1_06_in06 = reg_0160;
    61: op1_06_in06 = reg_0451;
    62: op1_06_in06 = reg_0117;
    94: op1_06_in06 = reg_0117;
    63: op1_06_in06 = reg_0254;
    64: op1_06_in06 = reg_0138;
    65: op1_06_in06 = reg_0175;
    66: op1_06_in06 = reg_0722;
    67: op1_06_in06 = reg_0707;
    68: op1_06_in06 = reg_0883;
    69: op1_06_in06 = imem04_in[55:52];
    70: op1_06_in06 = imem06_in[107:104];
    71: op1_06_in06 = imem00_in[111:108];
    72: op1_06_in06 = reg_0229;
    75: op1_06_in06 = reg_0753;
    76: op1_06_in06 = reg_0887;
    78: op1_06_in06 = reg_0240;
    79: op1_06_in06 = reg_0294;
    80: op1_06_in06 = reg_0502;
    81: op1_06_in06 = reg_0463;
    82: op1_06_in06 = imem07_in[31:28];
    83: op1_06_in06 = imem04_in[79:76];
    84: op1_06_in06 = reg_0733;
    85: op1_06_in06 = reg_0573;
    87: op1_06_in06 = reg_0550;
    88: op1_06_in06 = imem06_in[99:96];
    89: op1_06_in06 = reg_0073;
    90: op1_06_in06 = imem07_in[19:16];
    91: op1_06_in06 = reg_0532;
    92: op1_06_in06 = reg_0406;
    93: op1_06_in06 = imem02_in[91:88];
    95: op1_06_in06 = imem01_in[95:92];
    96: op1_06_in06 = imem02_in[39:36];
    97: op1_06_in06 = reg_0028;
    default: op1_06_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_06_inv06 = 1;
    8: op1_06_inv06 = 1;
    10: op1_06_inv06 = 1;
    11: op1_06_inv06 = 1;
    12: op1_06_inv06 = 1;
    13: op1_06_inv06 = 1;
    14: op1_06_inv06 = 1;
    16: op1_06_inv06 = 1;
    17: op1_06_inv06 = 1;
    3: op1_06_inv06 = 1;
    23: op1_06_inv06 = 1;
    24: op1_06_inv06 = 1;
    26: op1_06_inv06 = 1;
    29: op1_06_inv06 = 1;
    33: op1_06_inv06 = 1;
    34: op1_06_inv06 = 1;
    37: op1_06_inv06 = 1;
    38: op1_06_inv06 = 1;
    39: op1_06_inv06 = 1;
    40: op1_06_inv06 = 1;
    42: op1_06_inv06 = 1;
    44: op1_06_inv06 = 1;
    45: op1_06_inv06 = 1;
    46: op1_06_inv06 = 1;
    50: op1_06_inv06 = 1;
    52: op1_06_inv06 = 1;
    53: op1_06_inv06 = 1;
    55: op1_06_inv06 = 1;
    59: op1_06_inv06 = 1;
    63: op1_06_inv06 = 1;
    65: op1_06_inv06 = 1;
    66: op1_06_inv06 = 1;
    67: op1_06_inv06 = 1;
    68: op1_06_inv06 = 1;
    69: op1_06_inv06 = 1;
    70: op1_06_inv06 = 1;
    75: op1_06_inv06 = 1;
    76: op1_06_inv06 = 1;
    82: op1_06_inv06 = 1;
    87: op1_06_inv06 = 1;
    90: op1_06_inv06 = 1;
    91: op1_06_inv06 = 1;
    94: op1_06_inv06 = 1;
    96: op1_06_inv06 = 1;
    97: op1_06_inv06 = 1;
    default: op1_06_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in07 = imem02_in[111:108];
    93: op1_06_in07 = imem02_in[111:108];
    6: op1_06_in07 = reg_0687;
    12: op1_06_in07 = reg_0687;
    7: op1_06_in07 = reg_0550;
    8: op1_06_in07 = reg_0030;
    9: op1_06_in07 = imem02_in[115:112];
    10: op1_06_in07 = reg_0463;
    68: op1_06_in07 = reg_0463;
    11: op1_06_in07 = reg_0120;
    4: op1_06_in07 = reg_0435;
    13: op1_06_in07 = reg_0065;
    14: op1_06_in07 = imem07_in[99:96];
    15: op1_06_in07 = reg_0698;
    16: op1_06_in07 = reg_0993;
    17: op1_06_in07 = imem05_in[99:96];
    18: op1_06_in07 = reg_0338;
    19: op1_06_in07 = reg_0614;
    3: op1_06_in07 = reg_0174;
    20: op1_06_in07 = reg_0643;
    76: op1_06_in07 = reg_0643;
    21: op1_06_in07 = reg_0129;
    64: op1_06_in07 = reg_0129;
    22: op1_06_in07 = imem02_in[11:8];
    23: op1_06_in07 = imem02_in[23:20];
    24: op1_06_in07 = reg_0472;
    61: op1_06_in07 = reg_0472;
    25: op1_06_in07 = reg_0393;
    79: op1_06_in07 = reg_0393;
    26: op1_06_in07 = imem06_in[7:4];
    27: op1_06_in07 = reg_0385;
    28: op1_06_in07 = reg_0774;
    29: op1_06_in07 = imem02_in[75:72];
    30: op1_06_in07 = reg_0039;
    31: op1_06_in07 = reg_0956;
    32: op1_06_in07 = reg_0679;
    33: op1_06_in07 = reg_0216;
    34: op1_06_in07 = reg_0989;
    35: op1_06_in07 = imem00_in[87:84];
    37: op1_06_in07 = reg_0697;
    38: op1_06_in07 = reg_0685;
    39: op1_06_in07 = imem02_in[47:44];
    40: op1_06_in07 = imem04_in[75:72];
    41: op1_06_in07 = reg_0310;
    42: op1_06_in07 = reg_0029;
    43: op1_06_in07 = reg_0674;
    44: op1_06_in07 = reg_0667;
    45: op1_06_in07 = reg_0256;
    46: op1_06_in07 = reg_0250;
    47: op1_06_in07 = reg_0110;
    62: op1_06_in07 = reg_0110;
    48: op1_06_in07 = reg_0308;
    50: op1_06_in07 = imem06_in[103:100];
    51: op1_06_in07 = reg_0554;
    52: op1_06_in07 = reg_0650;
    53: op1_06_in07 = reg_0301;
    54: op1_06_in07 = imem05_in[43:40];
    55: op1_06_in07 = reg_0754;
    56: op1_06_in07 = reg_0894;
    58: op1_06_in07 = reg_0519;
    71: op1_06_in07 = reg_0519;
    59: op1_06_in07 = reg_0183;
    60: op1_06_in07 = reg_0737;
    63: op1_06_in07 = reg_0252;
    65: op1_06_in07 = reg_0167;
    66: op1_06_in07 = reg_0721;
    67: op1_06_in07 = reg_0727;
    69: op1_06_in07 = imem04_in[63:60];
    70: op1_06_in07 = reg_0080;
    72: op1_06_in07 = reg_0735;
    73: op1_06_in07 = imem07_in[83:80];
    75: op1_06_in07 = reg_0450;
    77: op1_06_in07 = imem02_in[123:120];
    78: op1_06_in07 = reg_0238;
    80: op1_06_in07 = reg_0640;
    81: op1_06_in07 = reg_0457;
    82: op1_06_in07 = imem07_in[43:40];
    83: op1_06_in07 = imem04_in[123:120];
    84: op1_06_in07 = reg_0821;
    85: op1_06_in07 = imem07_in[39:36];
    86: op1_06_in07 = reg_0900;
    87: op1_06_in07 = reg_0430;
    88: op1_06_in07 = reg_0351;
    89: op1_06_in07 = reg_0644;
    90: op1_06_in07 = imem07_in[31:28];
    91: op1_06_in07 = reg_0868;
    92: op1_06_in07 = reg_0420;
    94: op1_06_in07 = reg_0113;
    95: op1_06_in07 = imem01_in[111:108];
    96: op1_06_in07 = imem02_in[103:100];
    97: op1_06_in07 = reg_0810;
    default: op1_06_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_06_inv07 = 1;
    11: op1_06_inv07 = 1;
    12: op1_06_inv07 = 1;
    16: op1_06_inv07 = 1;
    17: op1_06_inv07 = 1;
    19: op1_06_inv07 = 1;
    21: op1_06_inv07 = 1;
    22: op1_06_inv07 = 1;
    25: op1_06_inv07 = 1;
    26: op1_06_inv07 = 1;
    27: op1_06_inv07 = 1;
    29: op1_06_inv07 = 1;
    30: op1_06_inv07 = 1;
    31: op1_06_inv07 = 1;
    32: op1_06_inv07 = 1;
    33: op1_06_inv07 = 1;
    34: op1_06_inv07 = 1;
    35: op1_06_inv07 = 1;
    38: op1_06_inv07 = 1;
    40: op1_06_inv07 = 1;
    41: op1_06_inv07 = 1;
    42: op1_06_inv07 = 1;
    43: op1_06_inv07 = 1;
    48: op1_06_inv07 = 1;
    51: op1_06_inv07 = 1;
    53: op1_06_inv07 = 1;
    56: op1_06_inv07 = 1;
    58: op1_06_inv07 = 1;
    64: op1_06_inv07 = 1;
    66: op1_06_inv07 = 1;
    72: op1_06_inv07 = 1;
    78: op1_06_inv07 = 1;
    81: op1_06_inv07 = 1;
    82: op1_06_inv07 = 1;
    85: op1_06_inv07 = 1;
    87: op1_06_inv07 = 1;
    88: op1_06_inv07 = 1;
    89: op1_06_inv07 = 1;
    90: op1_06_inv07 = 1;
    91: op1_06_inv07 = 1;
    92: op1_06_inv07 = 1;
    93: op1_06_inv07 = 1;
    95: op1_06_inv07 = 1;
    97: op1_06_inv07 = 1;
    default: op1_06_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in08 = imem02_in[127:124];
    6: op1_06_in08 = reg_0454;
    7: op1_06_in08 = reg_0529;
    8: op1_06_in08 = imem07_in[15:12];
    9: op1_06_in08 = imem02_in[123:120];
    10: op1_06_in08 = reg_0457;
    11: op1_06_in08 = reg_0114;
    12: op1_06_in08 = reg_0453;
    4: op1_06_in08 = reg_0161;
    13: op1_06_in08 = reg_0067;
    14: op1_06_in08 = imem07_in[107:104];
    15: op1_06_in08 = reg_0691;
    70: op1_06_in08 = reg_0691;
    16: op1_06_in08 = reg_0986;
    17: op1_06_in08 = imem05_in[103:100];
    18: op1_06_in08 = reg_0335;
    19: op1_06_in08 = reg_0607;
    3: op1_06_in08 = reg_0175;
    20: op1_06_in08 = reg_0659;
    21: op1_06_in08 = reg_0130;
    64: op1_06_in08 = reg_0130;
    22: op1_06_in08 = imem02_in[15:12];
    23: op1_06_in08 = imem02_in[31:28];
    94: op1_06_in08 = imem02_in[31:28];
    24: op1_06_in08 = reg_0467;
    25: op1_06_in08 = reg_0396;
    26: op1_06_in08 = imem06_in[71:68];
    27: op1_06_in08 = reg_0984;
    28: op1_06_in08 = reg_0777;
    29: op1_06_in08 = imem02_in[91:88];
    30: op1_06_in08 = reg_0096;
    31: op1_06_in08 = reg_0948;
    32: op1_06_in08 = reg_0674;
    33: op1_06_in08 = reg_1036;
    34: op1_06_in08 = reg_0981;
    35: op1_06_in08 = imem00_in[99:96];
    37: op1_06_in08 = reg_0698;
    38: op1_06_in08 = reg_0676;
    39: op1_06_in08 = imem02_in[71:68];
    40: op1_06_in08 = imem04_in[91:88];
    41: op1_06_in08 = reg_0016;
    42: op1_06_in08 = reg_0926;
    43: op1_06_in08 = reg_0460;
    44: op1_06_in08 = reg_0916;
    45: op1_06_in08 = reg_0251;
    46: op1_06_in08 = reg_0426;
    47: op1_06_in08 = imem02_in[51:48];
    48: op1_06_in08 = reg_0763;
    50: op1_06_in08 = imem06_in[107:104];
    51: op1_06_in08 = reg_0816;
    52: op1_06_in08 = reg_0657;
    53: op1_06_in08 = reg_1003;
    54: op1_06_in08 = imem05_in[55:52];
    55: op1_06_in08 = reg_0348;
    56: op1_06_in08 = reg_0780;
    58: op1_06_in08 = reg_0671;
    59: op1_06_in08 = reg_0166;
    60: op1_06_in08 = reg_0740;
    61: op1_06_in08 = reg_0474;
    62: op1_06_in08 = imem02_in[7:4];
    63: op1_06_in08 = reg_0023;
    65: op1_06_in08 = reg_0159;
    66: op1_06_in08 = reg_0303;
    67: op1_06_in08 = reg_0805;
    68: op1_06_in08 = reg_0455;
    69: op1_06_in08 = imem04_in[67:64];
    71: op1_06_in08 = reg_0768;
    72: op1_06_in08 = reg_0392;
    73: op1_06_in08 = imem07_in[119:116];
    75: op1_06_in08 = reg_0464;
    81: op1_06_in08 = reg_0464;
    76: op1_06_in08 = reg_0644;
    77: op1_06_in08 = reg_0907;
    78: op1_06_in08 = reg_0756;
    79: op1_06_in08 = reg_0025;
    80: op1_06_in08 = reg_0180;
    83: op1_06_in08 = reg_0850;
    84: op1_06_in08 = reg_0110;
    85: op1_06_in08 = imem07_in[51:48];
    90: op1_06_in08 = imem07_in[51:48];
    86: op1_06_in08 = reg_0684;
    87: op1_06_in08 = reg_0864;
    88: op1_06_in08 = reg_0754;
    89: op1_06_in08 = imem03_in[43:40];
    91: op1_06_in08 = reg_0181;
    92: op1_06_in08 = reg_0640;
    93: op1_06_in08 = reg_0750;
    95: op1_06_in08 = reg_0003;
    96: op1_06_in08 = reg_0844;
    97: op1_06_in08 = reg_0477;
    default: op1_06_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv08 = 1;
    7: op1_06_inv08 = 1;
    10: op1_06_inv08 = 1;
    11: op1_06_inv08 = 1;
    15: op1_06_inv08 = 1;
    18: op1_06_inv08 = 1;
    21: op1_06_inv08 = 1;
    24: op1_06_inv08 = 1;
    27: op1_06_inv08 = 1;
    28: op1_06_inv08 = 1;
    32: op1_06_inv08 = 1;
    33: op1_06_inv08 = 1;
    34: op1_06_inv08 = 1;
    38: op1_06_inv08 = 1;
    39: op1_06_inv08 = 1;
    40: op1_06_inv08 = 1;
    41: op1_06_inv08 = 1;
    43: op1_06_inv08 = 1;
    45: op1_06_inv08 = 1;
    50: op1_06_inv08 = 1;
    52: op1_06_inv08 = 1;
    53: op1_06_inv08 = 1;
    54: op1_06_inv08 = 1;
    55: op1_06_inv08 = 1;
    56: op1_06_inv08 = 1;
    58: op1_06_inv08 = 1;
    59: op1_06_inv08 = 1;
    60: op1_06_inv08 = 1;
    62: op1_06_inv08 = 1;
    66: op1_06_inv08 = 1;
    69: op1_06_inv08 = 1;
    70: op1_06_inv08 = 1;
    72: op1_06_inv08 = 1;
    73: op1_06_inv08 = 1;
    77: op1_06_inv08 = 1;
    79: op1_06_inv08 = 1;
    80: op1_06_inv08 = 1;
    87: op1_06_inv08 = 1;
    88: op1_06_inv08 = 1;
    90: op1_06_inv08 = 1;
    91: op1_06_inv08 = 1;
    92: op1_06_inv08 = 1;
    97: op1_06_inv08 = 1;
    default: op1_06_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in09 = reg_0650;
    6: op1_06_in09 = reg_0451;
    7: op1_06_in09 = reg_0555;
    8: op1_06_in09 = imem07_in[63:60];
    9: op1_06_in09 = reg_0642;
    10: op1_06_in09 = reg_0469;
    11: op1_06_in09 = reg_0109;
    12: op1_06_in09 = reg_0464;
    4: op1_06_in09 = reg_0159;
    13: op1_06_in09 = reg_0068;
    14: op1_06_in09 = reg_0721;
    15: op1_06_in09 = reg_0692;
    16: op1_06_in09 = reg_0977;
    34: op1_06_in09 = reg_0977;
    17: op1_06_in09 = imem05_in[107:104];
    18: op1_06_in09 = imem03_in[7:4];
    19: op1_06_in09 = reg_0605;
    3: op1_06_in09 = reg_0165;
    20: op1_06_in09 = reg_0325;
    21: op1_06_in09 = reg_0140;
    22: op1_06_in09 = imem02_in[31:28];
    23: op1_06_in09 = imem02_in[47:44];
    24: op1_06_in09 = reg_0468;
    25: op1_06_in09 = reg_0986;
    26: op1_06_in09 = imem06_in[75:72];
    27: op1_06_in09 = reg_1001;
    28: op1_06_in09 = imem05_in[3:0];
    29: op1_06_in09 = imem02_in[99:96];
    30: op1_06_in09 = reg_0857;
    31: op1_06_in09 = reg_0964;
    32: op1_06_in09 = reg_0678;
    33: op1_06_in09 = reg_0871;
    35: op1_06_in09 = imem00_in[103:100];
    37: op1_06_in09 = reg_0670;
    38: op1_06_in09 = reg_0674;
    39: op1_06_in09 = imem02_in[87:84];
    40: op1_06_in09 = imem04_in[115:112];
    41: op1_06_in09 = imem03_in[47:44];
    42: op1_06_in09 = reg_0622;
    43: op1_06_in09 = reg_0210;
    44: op1_06_in09 = reg_0842;
    45: op1_06_in09 = reg_0145;
    46: op1_06_in09 = reg_0321;
    66: op1_06_in09 = reg_0321;
    47: op1_06_in09 = imem02_in[95:92];
    48: op1_06_in09 = reg_0367;
    50: op1_06_in09 = reg_0613;
    51: op1_06_in09 = imem05_in[19:16];
    52: op1_06_in09 = reg_0326;
    53: op1_06_in09 = reg_0937;
    54: op1_06_in09 = reg_0962;
    55: op1_06_in09 = reg_0344;
    56: op1_06_in09 = reg_0008;
    87: op1_06_in09 = reg_0008;
    58: op1_06_in09 = reg_0684;
    59: op1_06_in09 = reg_0184;
    60: op1_06_in09 = reg_1017;
    61: op1_06_in09 = reg_0452;
    62: op1_06_in09 = imem02_in[75:72];
    63: op1_06_in09 = reg_0133;
    64: op1_06_in09 = imem06_in[3:0];
    67: op1_06_in09 = reg_0361;
    68: op1_06_in09 = reg_0474;
    69: op1_06_in09 = reg_1006;
    70: op1_06_in09 = reg_0351;
    71: op1_06_in09 = reg_0738;
    72: op1_06_in09 = reg_0632;
    73: op1_06_in09 = reg_0710;
    75: op1_06_in09 = reg_0477;
    81: op1_06_in09 = reg_0477;
    76: op1_06_in09 = reg_0037;
    77: op1_06_in09 = reg_0082;
    78: op1_06_in09 = reg_0038;
    79: op1_06_in09 = reg_1011;
    80: op1_06_in09 = reg_0182;
    83: op1_06_in09 = reg_0401;
    84: op1_06_in09 = reg_0352;
    85: op1_06_in09 = imem07_in[83:80];
    86: op1_06_in09 = reg_0883;
    88: op1_06_in09 = reg_0384;
    89: op1_06_in09 = imem03_in[55:52];
    90: op1_06_in09 = imem07_in[59:56];
    91: op1_06_in09 = reg_0714;
    92: op1_06_in09 = reg_0183;
    93: op1_06_in09 = reg_0285;
    94: op1_06_in09 = imem02_in[51:48];
    95: op1_06_in09 = reg_0273;
    96: op1_06_in09 = reg_0348;
    97: op1_06_in09 = reg_0481;
    default: op1_06_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_06_inv09 = 1;
    8: op1_06_inv09 = 1;
    9: op1_06_inv09 = 1;
    10: op1_06_inv09 = 1;
    11: op1_06_inv09 = 1;
    4: op1_06_inv09 = 1;
    15: op1_06_inv09 = 1;
    18: op1_06_inv09 = 1;
    19: op1_06_inv09 = 1;
    3: op1_06_inv09 = 1;
    21: op1_06_inv09 = 1;
    22: op1_06_inv09 = 1;
    24: op1_06_inv09 = 1;
    28: op1_06_inv09 = 1;
    32: op1_06_inv09 = 1;
    37: op1_06_inv09 = 1;
    39: op1_06_inv09 = 1;
    40: op1_06_inv09 = 1;
    41: op1_06_inv09 = 1;
    42: op1_06_inv09 = 1;
    45: op1_06_inv09 = 1;
    46: op1_06_inv09 = 1;
    47: op1_06_inv09 = 1;
    48: op1_06_inv09 = 1;
    51: op1_06_inv09 = 1;
    54: op1_06_inv09 = 1;
    55: op1_06_inv09 = 1;
    56: op1_06_inv09 = 1;
    58: op1_06_inv09 = 1;
    59: op1_06_inv09 = 1;
    60: op1_06_inv09 = 1;
    61: op1_06_inv09 = 1;
    62: op1_06_inv09 = 1;
    63: op1_06_inv09 = 1;
    67: op1_06_inv09 = 1;
    69: op1_06_inv09 = 1;
    72: op1_06_inv09 = 1;
    73: op1_06_inv09 = 1;
    77: op1_06_inv09 = 1;
    79: op1_06_inv09 = 1;
    80: op1_06_inv09 = 1;
    81: op1_06_inv09 = 1;
    83: op1_06_inv09 = 1;
    84: op1_06_inv09 = 1;
    85: op1_06_inv09 = 1;
    88: op1_06_inv09 = 1;
    89: op1_06_inv09 = 1;
    94: op1_06_inv09 = 1;
    95: op1_06_inv09 = 1;
    default: op1_06_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in10 = reg_0637;
    6: op1_06_in10 = reg_0470;
    7: op1_06_in10 = reg_0556;
    8: op1_06_in10 = imem07_in[67:64];
    9: op1_06_in10 = reg_0646;
    10: op1_06_in10 = reg_0476;
    11: op1_06_in10 = reg_0110;
    12: op1_06_in10 = reg_0469;
    75: op1_06_in10 = reg_0469;
    4: op1_06_in10 = reg_0171;
    13: op1_06_in10 = reg_0048;
    14: op1_06_in10 = reg_0703;
    15: op1_06_in10 = reg_0463;
    16: op1_06_in10 = reg_0988;
    17: op1_06_in10 = imem05_in[111:108];
    18: op1_06_in10 = imem03_in[31:28];
    19: op1_06_in10 = reg_0621;
    3: op1_06_in10 = reg_0185;
    80: op1_06_in10 = reg_0185;
    92: op1_06_in10 = reg_0185;
    20: op1_06_in10 = reg_0354;
    21: op1_06_in10 = imem06_in[3:0];
    22: op1_06_in10 = imem02_in[63:60];
    23: op1_06_in10 = imem02_in[51:48];
    24: op1_06_in10 = reg_0200;
    25: op1_06_in10 = reg_0989;
    26: op1_06_in10 = reg_0614;
    27: op1_06_in10 = reg_0999;
    28: op1_06_in10 = imem05_in[15:12];
    29: op1_06_in10 = imem02_in[107:104];
    30: op1_06_in10 = reg_0088;
    31: op1_06_in10 = reg_0952;
    32: op1_06_in10 = reg_0688;
    33: op1_06_in10 = reg_0111;
    34: op1_06_in10 = reg_0975;
    35: op1_06_in10 = reg_0681;
    37: op1_06_in10 = reg_0690;
    38: op1_06_in10 = reg_0671;
    39: op1_06_in10 = reg_0642;
    40: op1_06_in10 = reg_0277;
    41: op1_06_in10 = imem03_in[83:80];
    42: op1_06_in10 = imem07_in[27:24];
    56: op1_06_in10 = imem07_in[27:24];
    43: op1_06_in10 = reg_0187;
    44: op1_06_in10 = reg_0339;
    45: op1_06_in10 = reg_0142;
    46: op1_06_in10 = reg_0641;
    66: op1_06_in10 = reg_0641;
    47: op1_06_in10 = imem02_in[115:112];
    48: op1_06_in10 = reg_0057;
    50: op1_06_in10 = reg_0624;
    51: op1_06_in10 = imem05_in[23:20];
    52: op1_06_in10 = imem02_in[3:0];
    53: op1_06_in10 = reg_0306;
    54: op1_06_in10 = reg_0973;
    55: op1_06_in10 = reg_0351;
    58: op1_06_in10 = reg_0356;
    60: op1_06_in10 = reg_0232;
    61: op1_06_in10 = reg_0478;
    62: op1_06_in10 = imem02_in[79:76];
    63: op1_06_in10 = reg_0138;
    64: op1_06_in10 = imem06_in[87:84];
    67: op1_06_in10 = reg_0325;
    68: op1_06_in10 = reg_0471;
    69: op1_06_in10 = reg_0536;
    70: op1_06_in10 = reg_0926;
    71: op1_06_in10 = reg_0674;
    72: op1_06_in10 = reg_0222;
    73: op1_06_in10 = reg_0726;
    76: op1_06_in10 = reg_0083;
    77: op1_06_in10 = reg_0886;
    78: op1_06_in10 = reg_1008;
    79: op1_06_in10 = reg_0735;
    81: op1_06_in10 = reg_0460;
    83: op1_06_in10 = reg_0808;
    84: op1_06_in10 = reg_0634;
    85: op1_06_in10 = reg_0720;
    86: op1_06_in10 = reg_0828;
    87: op1_06_in10 = reg_0031;
    88: op1_06_in10 = reg_0895;
    89: op1_06_in10 = imem03_in[123:120];
    90: op1_06_in10 = imem07_in[111:108];
    91: op1_06_in10 = reg_0539;
    93: op1_06_in10 = reg_0639;
    94: op1_06_in10 = imem02_in[75:72];
    95: op1_06_in10 = reg_0555;
    96: op1_06_in10 = reg_0483;
    97: op1_06_in10 = reg_0473;
    default: op1_06_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv10 = 1;
    6: op1_06_inv10 = 1;
    8: op1_06_inv10 = 1;
    11: op1_06_inv10 = 1;
    12: op1_06_inv10 = 1;
    4: op1_06_inv10 = 1;
    13: op1_06_inv10 = 1;
    14: op1_06_inv10 = 1;
    15: op1_06_inv10 = 1;
    16: op1_06_inv10 = 1;
    20: op1_06_inv10 = 1;
    21: op1_06_inv10 = 1;
    22: op1_06_inv10 = 1;
    28: op1_06_inv10 = 1;
    29: op1_06_inv10 = 1;
    30: op1_06_inv10 = 1;
    32: op1_06_inv10 = 1;
    33: op1_06_inv10 = 1;
    34: op1_06_inv10 = 1;
    38: op1_06_inv10 = 1;
    40: op1_06_inv10 = 1;
    42: op1_06_inv10 = 1;
    44: op1_06_inv10 = 1;
    46: op1_06_inv10 = 1;
    48: op1_06_inv10 = 1;
    54: op1_06_inv10 = 1;
    55: op1_06_inv10 = 1;
    56: op1_06_inv10 = 1;
    60: op1_06_inv10 = 1;
    62: op1_06_inv10 = 1;
    63: op1_06_inv10 = 1;
    69: op1_06_inv10 = 1;
    70: op1_06_inv10 = 1;
    72: op1_06_inv10 = 1;
    73: op1_06_inv10 = 1;
    75: op1_06_inv10 = 1;
    76: op1_06_inv10 = 1;
    84: op1_06_inv10 = 1;
    85: op1_06_inv10 = 1;
    90: op1_06_inv10 = 1;
    91: op1_06_inv10 = 1;
    92: op1_06_inv10 = 1;
    93: op1_06_inv10 = 1;
    94: op1_06_inv10 = 1;
    95: op1_06_inv10 = 1;
    96: op1_06_inv10 = 1;
    default: op1_06_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in11 = reg_0660;
    22: op1_06_in11 = reg_0660;
    6: op1_06_in11 = reg_0208;
    24: op1_06_in11 = reg_0208;
    7: op1_06_in11 = reg_0304;
    8: op1_06_in11 = imem07_in[75:72];
    9: op1_06_in11 = reg_0661;
    10: op1_06_in11 = reg_0198;
    11: op1_06_in11 = imem02_in[47:44];
    12: op1_06_in11 = reg_0460;
    13: op1_06_in11 = reg_0050;
    14: op1_06_in11 = reg_0712;
    73: op1_06_in11 = reg_0712;
    15: op1_06_in11 = reg_0477;
    16: op1_06_in11 = reg_1000;
    34: op1_06_in11 = reg_1000;
    17: op1_06_in11 = reg_0963;
    18: op1_06_in11 = imem03_in[39:36];
    19: op1_06_in11 = reg_0619;
    20: op1_06_in11 = reg_0345;
    21: op1_06_in11 = imem06_in[15:12];
    23: op1_06_in11 = imem02_in[111:108];
    25: op1_06_in11 = reg_0977;
    26: op1_06_in11 = reg_0613;
    27: op1_06_in11 = reg_0989;
    28: op1_06_in11 = imem05_in[31:28];
    29: op1_06_in11 = reg_0658;
    30: op1_06_in11 = reg_0079;
    31: op1_06_in11 = reg_0806;
    32: op1_06_in11 = reg_0687;
    33: op1_06_in11 = reg_0116;
    35: op1_06_in11 = reg_0696;
    37: op1_06_in11 = reg_0699;
    38: op1_06_in11 = reg_0668;
    39: op1_06_in11 = reg_0645;
    40: op1_06_in11 = reg_0306;
    41: op1_06_in11 = imem03_in[99:96];
    42: op1_06_in11 = imem07_in[79:76];
    43: op1_06_in11 = reg_0211;
    44: op1_06_in11 = reg_0865;
    45: op1_06_in11 = reg_0143;
    46: op1_06_in11 = reg_0589;
    47: op1_06_in11 = reg_0639;
    48: op1_06_in11 = reg_0448;
    50: op1_06_in11 = reg_0611;
    51: op1_06_in11 = imem05_in[63:60];
    52: op1_06_in11 = imem02_in[35:32];
    53: op1_06_in11 = reg_1020;
    54: op1_06_in11 = reg_0955;
    55: op1_06_in11 = reg_0393;
    56: op1_06_in11 = imem07_in[51:48];
    58: op1_06_in11 = reg_0674;
    60: op1_06_in11 = reg_1053;
    61: op1_06_in11 = reg_0214;
    62: op1_06_in11 = imem02_in[115:112];
    63: op1_06_in11 = imem06_in[91:88];
    64: op1_06_in11 = reg_0080;
    66: op1_06_in11 = reg_0599;
    67: op1_06_in11 = reg_0422;
    68: op1_06_in11 = reg_0210;
    69: op1_06_in11 = reg_1009;
    70: op1_06_in11 = reg_1030;
    71: op1_06_in11 = reg_0828;
    72: op1_06_in11 = reg_0695;
    75: op1_06_in11 = reg_0468;
    76: op1_06_in11 = reg_0761;
    77: op1_06_in11 = reg_0095;
    78: op1_06_in11 = reg_0779;
    79: op1_06_in11 = reg_0384;
    81: op1_06_in11 = reg_0473;
    83: op1_06_in11 = reg_0072;
    84: op1_06_in11 = reg_0261;
    85: op1_06_in11 = reg_0721;
    86: op1_06_in11 = reg_0465;
    87: op1_06_in11 = reg_0586;
    88: op1_06_in11 = reg_1028;
    89: op1_06_in11 = imem03_in[127:124];
    90: op1_06_in11 = reg_0717;
    91: op1_06_in11 = reg_0701;
    93: op1_06_in11 = reg_0055;
    94: op1_06_in11 = imem02_in[79:76];
    95: op1_06_in11 = reg_0101;
    96: op1_06_in11 = reg_0052;
    97: op1_06_in11 = reg_0474;
    default: op1_06_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_06_inv11 = 1;
    8: op1_06_inv11 = 1;
    9: op1_06_inv11 = 1;
    11: op1_06_inv11 = 1;
    15: op1_06_inv11 = 1;
    17: op1_06_inv11 = 1;
    19: op1_06_inv11 = 1;
    22: op1_06_inv11 = 1;
    23: op1_06_inv11 = 1;
    24: op1_06_inv11 = 1;
    26: op1_06_inv11 = 1;
    30: op1_06_inv11 = 1;
    33: op1_06_inv11 = 1;
    37: op1_06_inv11 = 1;
    39: op1_06_inv11 = 1;
    40: op1_06_inv11 = 1;
    41: op1_06_inv11 = 1;
    44: op1_06_inv11 = 1;
    48: op1_06_inv11 = 1;
    50: op1_06_inv11 = 1;
    51: op1_06_inv11 = 1;
    53: op1_06_inv11 = 1;
    55: op1_06_inv11 = 1;
    56: op1_06_inv11 = 1;
    58: op1_06_inv11 = 1;
    60: op1_06_inv11 = 1;
    61: op1_06_inv11 = 1;
    64: op1_06_inv11 = 1;
    66: op1_06_inv11 = 1;
    68: op1_06_inv11 = 1;
    70: op1_06_inv11 = 1;
    77: op1_06_inv11 = 1;
    81: op1_06_inv11 = 1;
    83: op1_06_inv11 = 1;
    89: op1_06_inv11 = 1;
    90: op1_06_inv11 = 1;
    93: op1_06_inv11 = 1;
    96: op1_06_inv11 = 1;
    default: op1_06_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in12 = reg_0661;
    6: op1_06_in12 = reg_0210;
    61: op1_06_in12 = reg_0210;
    7: op1_06_in12 = reg_0294;
    8: op1_06_in12 = imem07_in[91:88];
    9: op1_06_in12 = reg_0648;
    47: op1_06_in12 = reg_0648;
    10: op1_06_in12 = reg_0788;
    11: op1_06_in12 = imem02_in[55:52];
    12: op1_06_in12 = reg_0481;
    13: op1_06_in12 = reg_0963;
    14: op1_06_in12 = reg_0715;
    15: op1_06_in12 = reg_0469;
    86: op1_06_in12 = reg_0469;
    16: op1_06_in12 = imem04_in[3:0];
    17: op1_06_in12 = reg_0966;
    18: op1_06_in12 = imem03_in[79:76];
    19: op1_06_in12 = reg_0615;
    20: op1_06_in12 = reg_0355;
    21: op1_06_in12 = imem06_in[35:32];
    22: op1_06_in12 = reg_0656;
    23: op1_06_in12 = imem02_in[115:112];
    24: op1_06_in12 = reg_0207;
    25: op1_06_in12 = reg_0988;
    26: op1_06_in12 = reg_0605;
    27: op1_06_in12 = reg_0975;
    28: op1_06_in12 = imem05_in[39:36];
    29: op1_06_in12 = reg_0664;
    30: op1_06_in12 = imem03_in[15:12];
    31: op1_06_in12 = reg_0251;
    32: op1_06_in12 = reg_0454;
    33: op1_06_in12 = reg_0114;
    34: op1_06_in12 = imem04_in[7:4];
    35: op1_06_in12 = reg_0677;
    37: op1_06_in12 = reg_0463;
    38: op1_06_in12 = reg_0669;
    39: op1_06_in12 = reg_0651;
    40: op1_06_in12 = reg_0540;
    41: op1_06_in12 = imem03_in[127:124];
    42: op1_06_in12 = imem07_in[115:112];
    43: op1_06_in12 = reg_0186;
    44: op1_06_in12 = reg_0098;
    45: op1_06_in12 = reg_0140;
    46: op1_06_in12 = reg_0180;
    48: op1_06_in12 = imem05_in[31:28];
    50: op1_06_in12 = reg_0754;
    51: op1_06_in12 = imem05_in[71:68];
    52: op1_06_in12 = imem02_in[79:76];
    53: op1_06_in12 = reg_0292;
    54: op1_06_in12 = reg_0954;
    55: op1_06_in12 = reg_0264;
    56: op1_06_in12 = imem07_in[59:56];
    58: op1_06_in12 = reg_0476;
    60: op1_06_in12 = reg_0273;
    62: op1_06_in12 = reg_0657;
    63: op1_06_in12 = imem06_in[123:120];
    64: op1_06_in12 = reg_0696;
    66: op1_06_in12 = reg_0640;
    67: op1_06_in12 = reg_0433;
    68: op1_06_in12 = reg_0194;
    69: op1_06_in12 = reg_0055;
    70: op1_06_in12 = reg_0011;
    71: op1_06_in12 = reg_0687;
    72: op1_06_in12 = reg_0289;
    73: op1_06_in12 = reg_0724;
    75: op1_06_in12 = reg_0479;
    81: op1_06_in12 = reg_0479;
    76: op1_06_in12 = reg_0876;
    77: op1_06_in12 = reg_0248;
    78: op1_06_in12 = reg_0767;
    79: op1_06_in12 = reg_1030;
    83: op1_06_in12 = reg_0432;
    84: op1_06_in12 = imem02_in[19:16];
    85: op1_06_in12 = reg_0442;
    87: op1_06_in12 = reg_0537;
    88: op1_06_in12 = reg_0698;
    89: op1_06_in12 = reg_0976;
    90: op1_06_in12 = reg_0744;
    91: op1_06_in12 = reg_0449;
    93: op1_06_in12 = reg_0279;
    94: op1_06_in12 = imem02_in[103:100];
    95: op1_06_in12 = reg_0115;
    96: op1_06_in12 = reg_0423;
    97: op1_06_in12 = reg_0478;
    default: op1_06_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv12 = 1;
    7: op1_06_inv12 = 1;
    8: op1_06_inv12 = 1;
    9: op1_06_inv12 = 1;
    13: op1_06_inv12 = 1;
    17: op1_06_inv12 = 1;
    19: op1_06_inv12 = 1;
    23: op1_06_inv12 = 1;
    24: op1_06_inv12 = 1;
    25: op1_06_inv12 = 1;
    28: op1_06_inv12 = 1;
    29: op1_06_inv12 = 1;
    31: op1_06_inv12 = 1;
    35: op1_06_inv12 = 1;
    38: op1_06_inv12 = 1;
    40: op1_06_inv12 = 1;
    41: op1_06_inv12 = 1;
    43: op1_06_inv12 = 1;
    45: op1_06_inv12 = 1;
    54: op1_06_inv12 = 1;
    60: op1_06_inv12 = 1;
    63: op1_06_inv12 = 1;
    66: op1_06_inv12 = 1;
    67: op1_06_inv12 = 1;
    68: op1_06_inv12 = 1;
    73: op1_06_inv12 = 1;
    75: op1_06_inv12 = 1;
    81: op1_06_inv12 = 1;
    86: op1_06_inv12 = 1;
    90: op1_06_inv12 = 1;
    93: op1_06_inv12 = 1;
    95: op1_06_inv12 = 1;
    default: op1_06_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in13 = reg_0639;
    6: op1_06_in13 = reg_0204;
    7: op1_06_in13 = reg_0277;
    8: op1_06_in13 = imem07_in[95:92];
    9: op1_06_in13 = reg_0638;
    10: op1_06_in13 = reg_0779;
    11: op1_06_in13 = imem02_in[63:60];
    12: op1_06_in13 = reg_0473;
    13: op1_06_in13 = reg_0970;
    14: op1_06_in13 = reg_0701;
    15: op1_06_in13 = reg_0466;
    86: op1_06_in13 = reg_0466;
    16: op1_06_in13 = imem04_in[75:72];
    17: op1_06_in13 = reg_0949;
    18: op1_06_in13 = imem03_in[115:112];
    19: op1_06_in13 = reg_0601;
    20: op1_06_in13 = reg_0314;
    21: op1_06_in13 = imem06_in[39:36];
    22: op1_06_in13 = reg_0641;
    23: op1_06_in13 = imem02_in[123:120];
    24: op1_06_in13 = reg_0211;
    75: op1_06_in13 = reg_0211;
    25: op1_06_in13 = imem04_in[3:0];
    26: op1_06_in13 = reg_0616;
    27: op1_06_in13 = reg_0994;
    28: op1_06_in13 = imem05_in[63:60];
    29: op1_06_in13 = reg_0647;
    30: op1_06_in13 = imem03_in[43:40];
    31: op1_06_in13 = reg_0275;
    32: op1_06_in13 = reg_0469;
    33: op1_06_in13 = reg_0100;
    34: op1_06_in13 = imem04_in[11:8];
    35: op1_06_in13 = reg_0691;
    64: op1_06_in13 = reg_0691;
    37: op1_06_in13 = reg_0450;
    38: op1_06_in13 = reg_0465;
    39: op1_06_in13 = reg_0842;
    40: op1_06_in13 = reg_0537;
    69: op1_06_in13 = reg_0537;
    41: op1_06_in13 = reg_0006;
    42: op1_06_in13 = reg_0722;
    43: op1_06_in13 = reg_0201;
    44: op1_06_in13 = reg_0482;
    45: op1_06_in13 = imem06_in[31:28];
    46: op1_06_in13 = reg_0167;
    47: op1_06_in13 = reg_0096;
    48: op1_06_in13 = imem05_in[67:64];
    50: op1_06_in13 = reg_0344;
    51: op1_06_in13 = imem05_in[87:84];
    52: op1_06_in13 = imem02_in[91:88];
    53: op1_06_in13 = reg_0848;
    54: op1_06_in13 = reg_0956;
    55: op1_06_in13 = reg_0332;
    56: op1_06_in13 = imem07_in[99:96];
    58: op1_06_in13 = reg_0480;
    60: op1_06_in13 = reg_0112;
    61: op1_06_in13 = reg_0188;
    62: op1_06_in13 = reg_0326;
    63: op1_06_in13 = reg_0625;
    66: op1_06_in13 = reg_0431;
    67: op1_06_in13 = reg_0350;
    68: op1_06_in13 = imem01_in[15:12];
    70: op1_06_in13 = reg_0816;
    71: op1_06_in13 = reg_0464;
    72: op1_06_in13 = reg_0403;
    73: op1_06_in13 = reg_0713;
    76: op1_06_in13 = reg_0091;
    77: op1_06_in13 = reg_0331;
    78: op1_06_in13 = reg_0376;
    79: op1_06_in13 = reg_0624;
    81: op1_06_in13 = reg_0186;
    83: op1_06_in13 = reg_0243;
    84: op1_06_in13 = imem02_in[35:32];
    85: op1_06_in13 = reg_0575;
    87: op1_06_in13 = reg_0123;
    88: op1_06_in13 = reg_0928;
    89: op1_06_in13 = reg_0342;
    90: op1_06_in13 = reg_0406;
    93: op1_06_in13 = reg_0664;
    94: op1_06_in13 = imem02_in[111:108];
    95: op1_06_in13 = reg_0113;
    96: op1_06_in13 = reg_0248;
    97: op1_06_in13 = reg_0212;
    default: op1_06_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv13 = 1;
    6: op1_06_inv13 = 1;
    8: op1_06_inv13 = 1;
    11: op1_06_inv13 = 1;
    14: op1_06_inv13 = 1;
    19: op1_06_inv13 = 1;
    20: op1_06_inv13 = 1;
    21: op1_06_inv13 = 1;
    23: op1_06_inv13 = 1;
    24: op1_06_inv13 = 1;
    25: op1_06_inv13 = 1;
    29: op1_06_inv13 = 1;
    31: op1_06_inv13 = 1;
    35: op1_06_inv13 = 1;
    38: op1_06_inv13 = 1;
    39: op1_06_inv13 = 1;
    40: op1_06_inv13 = 1;
    41: op1_06_inv13 = 1;
    42: op1_06_inv13 = 1;
    47: op1_06_inv13 = 1;
    50: op1_06_inv13 = 1;
    52: op1_06_inv13 = 1;
    53: op1_06_inv13 = 1;
    55: op1_06_inv13 = 1;
    56: op1_06_inv13 = 1;
    58: op1_06_inv13 = 1;
    64: op1_06_inv13 = 1;
    66: op1_06_inv13 = 1;
    67: op1_06_inv13 = 1;
    69: op1_06_inv13 = 1;
    73: op1_06_inv13 = 1;
    75: op1_06_inv13 = 1;
    76: op1_06_inv13 = 1;
    77: op1_06_inv13 = 1;
    78: op1_06_inv13 = 1;
    83: op1_06_inv13 = 1;
    85: op1_06_inv13 = 1;
    86: op1_06_inv13 = 1;
    88: op1_06_inv13 = 1;
    90: op1_06_inv13 = 1;
    94: op1_06_inv13 = 1;
    95: op1_06_inv13 = 1;
    97: op1_06_inv13 = 1;
    default: op1_06_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in14 = reg_0640;
    6: op1_06_in14 = reg_0203;
    7: op1_06_in14 = reg_0059;
    8: op1_06_in14 = imem07_in[111:108];
    56: op1_06_in14 = imem07_in[111:108];
    9: op1_06_in14 = reg_0659;
    10: op1_06_in14 = reg_0765;
    11: op1_06_in14 = reg_0642;
    12: op1_06_in14 = reg_0467;
    13: op1_06_in14 = reg_0959;
    14: op1_06_in14 = reg_0700;
    15: op1_06_in14 = reg_0468;
    16: op1_06_in14 = imem04_in[99:96];
    17: op1_06_in14 = reg_0968;
    18: op1_06_in14 = reg_0602;
    19: op1_06_in14 = reg_0402;
    20: op1_06_in14 = reg_0096;
    21: op1_06_in14 = reg_0628;
    22: op1_06_in14 = reg_0345;
    23: op1_06_in14 = reg_0666;
    24: op1_06_in14 = imem01_in[23:20];
    25: op1_06_in14 = imem04_in[15:12];
    26: op1_06_in14 = reg_0619;
    27: op1_06_in14 = imem04_in[71:68];
    28: op1_06_in14 = imem05_in[115:112];
    29: op1_06_in14 = reg_0667;
    30: op1_06_in14 = reg_0598;
    31: op1_06_in14 = reg_0825;
    32: op1_06_in14 = reg_0472;
    33: op1_06_in14 = imem02_in[11:8];
    34: op1_06_in14 = imem04_in[19:16];
    35: op1_06_in14 = reg_0688;
    37: op1_06_in14 = reg_0455;
    38: op1_06_in14 = reg_0450;
    39: op1_06_in14 = reg_0095;
    40: op1_06_in14 = reg_0763;
    41: op1_06_in14 = reg_0940;
    42: op1_06_in14 = reg_0719;
    43: op1_06_in14 = reg_0212;
    44: op1_06_in14 = reg_0761;
    45: op1_06_in14 = imem06_in[79:76];
    46: op1_06_in14 = reg_0160;
    47: op1_06_in14 = reg_0318;
    48: op1_06_in14 = imem05_in[71:68];
    50: op1_06_in14 = reg_0395;
    51: op1_06_in14 = imem05_in[111:108];
    52: op1_06_in14 = imem02_in[127:124];
    53: op1_06_in14 = reg_0076;
    54: op1_06_in14 = reg_0951;
    55: op1_06_in14 = reg_0629;
    58: op1_06_in14 = reg_0214;
    60: op1_06_in14 = reg_0860;
    61: op1_06_in14 = reg_0213;
    62: op1_06_in14 = reg_0649;
    63: op1_06_in14 = reg_0694;
    64: op1_06_in14 = reg_0626;
    66: op1_06_in14 = reg_0162;
    67: op1_06_in14 = reg_0589;
    68: op1_06_in14 = reg_0586;
    69: op1_06_in14 = reg_0568;
    70: op1_06_in14 = reg_0630;
    71: op1_06_in14 = reg_0461;
    72: op1_06_in14 = imem07_in[11:8];
    73: op1_06_in14 = reg_0422;
    75: op1_06_in14 = reg_0201;
    76: op1_06_in14 = reg_0484;
    77: op1_06_in14 = reg_0347;
    78: op1_06_in14 = reg_0597;
    79: op1_06_in14 = reg_0863;
    81: op1_06_in14 = reg_0198;
    83: op1_06_in14 = reg_0108;
    84: op1_06_in14 = imem02_in[39:36];
    85: op1_06_in14 = reg_0002;
    86: op1_06_in14 = reg_0475;
    87: op1_06_in14 = reg_0752;
    88: op1_06_in14 = reg_0382;
    89: op1_06_in14 = reg_0051;
    90: op1_06_in14 = reg_0419;
    93: op1_06_in14 = reg_0359;
    94: op1_06_in14 = imem02_in[115:112];
    95: op1_06_in14 = reg_0110;
    96: op1_06_in14 = reg_0054;
    97: op1_06_in14 = imem01_in[11:8];
    default: op1_06_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv14 = 1;
    7: op1_06_inv14 = 1;
    11: op1_06_inv14 = 1;
    15: op1_06_inv14 = 1;
    16: op1_06_inv14 = 1;
    19: op1_06_inv14 = 1;
    22: op1_06_inv14 = 1;
    24: op1_06_inv14 = 1;
    26: op1_06_inv14 = 1;
    29: op1_06_inv14 = 1;
    32: op1_06_inv14 = 1;
    33: op1_06_inv14 = 1;
    35: op1_06_inv14 = 1;
    42: op1_06_inv14 = 1;
    43: op1_06_inv14 = 1;
    44: op1_06_inv14 = 1;
    45: op1_06_inv14 = 1;
    48: op1_06_inv14 = 1;
    52: op1_06_inv14 = 1;
    56: op1_06_inv14 = 1;
    60: op1_06_inv14 = 1;
    61: op1_06_inv14 = 1;
    62: op1_06_inv14 = 1;
    67: op1_06_inv14 = 1;
    75: op1_06_inv14 = 1;
    76: op1_06_inv14 = 1;
    78: op1_06_inv14 = 1;
    79: op1_06_inv14 = 1;
    81: op1_06_inv14 = 1;
    83: op1_06_inv14 = 1;
    84: op1_06_inv14 = 1;
    85: op1_06_inv14 = 1;
    87: op1_06_inv14 = 1;
    88: op1_06_inv14 = 1;
    89: op1_06_inv14 = 1;
    90: op1_06_inv14 = 1;
    94: op1_06_inv14 = 1;
    95: op1_06_inv14 = 1;
    96: op1_06_inv14 = 1;
    97: op1_06_inv14 = 1;
    default: op1_06_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in15 = reg_0641;
    90: op1_06_in15 = reg_0641;
    6: op1_06_in15 = reg_0213;
    81: op1_06_in15 = reg_0213;
    7: op1_06_in15 = reg_0062;
    8: op1_06_in15 = reg_0723;
    9: op1_06_in15 = reg_0636;
    10: op1_06_in15 = reg_0789;
    11: op1_06_in15 = reg_0654;
    12: op1_06_in15 = reg_0474;
    13: op1_06_in15 = reg_0947;
    14: op1_06_in15 = reg_0441;
    15: op1_06_in15 = reg_0459;
    16: op1_06_in15 = reg_0544;
    17: op1_06_in15 = reg_0943;
    18: op1_06_in15 = reg_0591;
    19: op1_06_in15 = reg_0332;
    20: op1_06_in15 = reg_0097;
    21: op1_06_in15 = reg_0632;
    22: op1_06_in15 = reg_0318;
    23: op1_06_in15 = reg_0646;
    24: op1_06_in15 = imem01_in[107:104];
    25: op1_06_in15 = imem04_in[59:56];
    26: op1_06_in15 = reg_0601;
    27: op1_06_in15 = imem04_in[79:76];
    28: op1_06_in15 = reg_0973;
    29: op1_06_in15 = reg_0081;
    30: op1_06_in15 = reg_0582;
    31: op1_06_in15 = reg_0142;
    32: op1_06_in15 = reg_0189;
    33: op1_06_in15 = imem02_in[35:32];
    34: op1_06_in15 = imem04_in[23:20];
    35: op1_06_in15 = reg_0453;
    37: op1_06_in15 = reg_0466;
    38: op1_06_in15 = reg_0208;
    58: op1_06_in15 = reg_0208;
    39: op1_06_in15 = reg_0096;
    40: op1_06_in15 = reg_0268;
    41: op1_06_in15 = reg_0573;
    42: op1_06_in15 = reg_0710;
    43: op1_06_in15 = reg_0190;
    44: op1_06_in15 = reg_0867;
    45: op1_06_in15 = imem06_in[87:84];
    46: op1_06_in15 = reg_0183;
    47: op1_06_in15 = reg_0857;
    48: op1_06_in15 = imem05_in[79:76];
    50: op1_06_in15 = reg_0391;
    51: op1_06_in15 = imem05_in[119:116];
    52: op1_06_in15 = reg_0083;
    53: op1_06_in15 = reg_0584;
    54: op1_06_in15 = reg_0953;
    55: op1_06_in15 = reg_0630;
    56: op1_06_in15 = imem07_in[123:120];
    60: op1_06_in15 = reg_0101;
    61: op1_06_in15 = reg_0205;
    62: op1_06_in15 = reg_0645;
    63: op1_06_in15 = reg_0262;
    64: op1_06_in15 = reg_0895;
    67: op1_06_in15 = reg_0868;
    68: op1_06_in15 = reg_0762;
    69: op1_06_in15 = reg_0524;
    87: op1_06_in15 = reg_0524;
    70: op1_06_in15 = reg_0957;
    71: op1_06_in15 = reg_0473;
    72: op1_06_in15 = imem07_in[27:24];
    73: op1_06_in15 = reg_0406;
    75: op1_06_in15 = imem01_in[39:36];
    76: op1_06_in15 = imem03_in[7:4];
    77: op1_06_in15 = reg_0772;
    78: op1_06_in15 = reg_0385;
    79: op1_06_in15 = reg_0380;
    83: op1_06_in15 = reg_0542;
    84: op1_06_in15 = imem02_in[71:68];
    85: op1_06_in15 = reg_0250;
    86: op1_06_in15 = reg_0472;
    88: op1_06_in15 = reg_0921;
    89: op1_06_in15 = reg_0672;
    93: op1_06_in15 = reg_0408;
    94: op1_06_in15 = reg_0750;
    95: op1_06_in15 = imem02_in[103:100];
    96: op1_06_in15 = reg_0347;
    97: op1_06_in15 = imem01_in[67:64];
    default: op1_06_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_06_inv15 = 1;
    9: op1_06_inv15 = 1;
    10: op1_06_inv15 = 1;
    12: op1_06_inv15 = 1;
    13: op1_06_inv15 = 1;
    15: op1_06_inv15 = 1;
    20: op1_06_inv15 = 1;
    21: op1_06_inv15 = 1;
    25: op1_06_inv15 = 1;
    26: op1_06_inv15 = 1;
    27: op1_06_inv15 = 1;
    28: op1_06_inv15 = 1;
    29: op1_06_inv15 = 1;
    32: op1_06_inv15 = 1;
    37: op1_06_inv15 = 1;
    38: op1_06_inv15 = 1;
    40: op1_06_inv15 = 1;
    41: op1_06_inv15 = 1;
    43: op1_06_inv15 = 1;
    44: op1_06_inv15 = 1;
    47: op1_06_inv15 = 1;
    48: op1_06_inv15 = 1;
    50: op1_06_inv15 = 1;
    51: op1_06_inv15 = 1;
    52: op1_06_inv15 = 1;
    53: op1_06_inv15 = 1;
    54: op1_06_inv15 = 1;
    56: op1_06_inv15 = 1;
    58: op1_06_inv15 = 1;
    60: op1_06_inv15 = 1;
    63: op1_06_inv15 = 1;
    71: op1_06_inv15 = 1;
    73: op1_06_inv15 = 1;
    76: op1_06_inv15 = 1;
    77: op1_06_inv15 = 1;
    78: op1_06_inv15 = 1;
    79: op1_06_inv15 = 1;
    81: op1_06_inv15 = 1;
    88: op1_06_inv15 = 1;
    89: op1_06_inv15 = 1;
    90: op1_06_inv15 = 1;
    95: op1_06_inv15 = 1;
    97: op1_06_inv15 = 1;
    default: op1_06_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in16 = reg_0333;
    6: op1_06_in16 = reg_0202;
    43: op1_06_in16 = reg_0202;
    7: op1_06_in16 = reg_0058;
    8: op1_06_in16 = reg_0430;
    9: op1_06_in16 = reg_0358;
    41: op1_06_in16 = reg_0358;
    10: op1_06_in16 = reg_0218;
    93: op1_06_in16 = reg_0218;
    11: op1_06_in16 = reg_0646;
    12: op1_06_in16 = reg_0471;
    13: op1_06_in16 = reg_0217;
    14: op1_06_in16 = reg_0422;
    15: op1_06_in16 = reg_0204;
    16: op1_06_in16 = reg_0536;
    17: op1_06_in16 = reg_0953;
    18: op1_06_in16 = reg_0570;
    19: op1_06_in16 = reg_0372;
    20: op1_06_in16 = imem03_in[7:4];
    21: op1_06_in16 = reg_0402;
    22: op1_06_in16 = reg_0330;
    23: op1_06_in16 = reg_0648;
    24: op1_06_in16 = imem01_in[115:112];
    25: op1_06_in16 = imem04_in[67:64];
    26: op1_06_in16 = reg_0379;
    27: op1_06_in16 = imem04_in[111:108];
    28: op1_06_in16 = reg_0943;
    29: op1_06_in16 = reg_0097;
    30: op1_06_in16 = reg_0596;
    55: op1_06_in16 = reg_0596;
    31: op1_06_in16 = reg_0139;
    32: op1_06_in16 = reg_0193;
    33: op1_06_in16 = imem02_in[43:40];
    34: op1_06_in16 = imem04_in[35:32];
    35: op1_06_in16 = reg_0451;
    37: op1_06_in16 = reg_0459;
    38: op1_06_in16 = reg_0203;
    39: op1_06_in16 = reg_0290;
    40: op1_06_in16 = reg_0296;
    42: op1_06_in16 = reg_0731;
    44: op1_06_in16 = reg_0876;
    52: op1_06_in16 = reg_0876;
    45: op1_06_in16 = imem06_in[107:104];
    46: op1_06_in16 = reg_0177;
    47: op1_06_in16 = reg_0772;
    48: op1_06_in16 = imem05_in[83:80];
    50: op1_06_in16 = reg_0386;
    51: op1_06_in16 = reg_0958;
    53: op1_06_in16 = reg_0815;
    54: op1_06_in16 = reg_0063;
    56: op1_06_in16 = reg_0720;
    58: op1_06_in16 = reg_0195;
    60: op1_06_in16 = reg_0110;
    61: op1_06_in16 = reg_0190;
    62: op1_06_in16 = reg_0052;
    63: op1_06_in16 = reg_0384;
    64: op1_06_in16 = reg_0533;
    67: op1_06_in16 = reg_0640;
    68: op1_06_in16 = reg_0236;
    69: op1_06_in16 = reg_0076;
    70: op1_06_in16 = reg_0219;
    71: op1_06_in16 = reg_0470;
    72: op1_06_in16 = imem07_in[43:40];
    73: op1_06_in16 = reg_0181;
    75: op1_06_in16 = imem01_in[59:56];
    76: op1_06_in16 = imem03_in[39:36];
    77: op1_06_in16 = reg_0482;
    78: op1_06_in16 = reg_0987;
    79: op1_06_in16 = reg_0695;
    81: op1_06_in16 = reg_0196;
    83: op1_06_in16 = reg_0044;
    84: op1_06_in16 = imem02_in[111:108];
    95: op1_06_in16 = imem02_in[111:108];
    85: op1_06_in16 = reg_0325;
    86: op1_06_in16 = reg_0456;
    87: op1_06_in16 = reg_0074;
    88: op1_06_in16 = reg_0026;
    89: op1_06_in16 = reg_0376;
    90: op1_06_in16 = reg_0599;
    94: op1_06_in16 = reg_0666;
    96: op1_06_in16 = reg_0776;
    97: op1_06_in16 = imem01_in[71:68];
    default: op1_06_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv16 = 1;
    7: op1_06_inv16 = 1;
    8: op1_06_inv16 = 1;
    11: op1_06_inv16 = 1;
    12: op1_06_inv16 = 1;
    14: op1_06_inv16 = 1;
    16: op1_06_inv16 = 1;
    22: op1_06_inv16 = 1;
    24: op1_06_inv16 = 1;
    25: op1_06_inv16 = 1;
    37: op1_06_inv16 = 1;
    38: op1_06_inv16 = 1;
    41: op1_06_inv16 = 1;
    43: op1_06_inv16 = 1;
    45: op1_06_inv16 = 1;
    46: op1_06_inv16 = 1;
    47: op1_06_inv16 = 1;
    52: op1_06_inv16 = 1;
    55: op1_06_inv16 = 1;
    56: op1_06_inv16 = 1;
    58: op1_06_inv16 = 1;
    60: op1_06_inv16 = 1;
    62: op1_06_inv16 = 1;
    71: op1_06_inv16 = 1;
    78: op1_06_inv16 = 1;
    79: op1_06_inv16 = 1;
    83: op1_06_inv16 = 1;
    84: op1_06_inv16 = 1;
    86: op1_06_inv16 = 1;
    93: op1_06_inv16 = 1;
    94: op1_06_inv16 = 1;
    97: op1_06_inv16 = 1;
    default: op1_06_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in17 = reg_0345;
    6: op1_06_in17 = imem01_in[35:32];
    7: op1_06_in17 = reg_0066;
    8: op1_06_in17 = reg_0445;
    9: op1_06_in17 = reg_0364;
    10: op1_06_in17 = reg_0224;
    11: op1_06_in17 = reg_0656;
    96: op1_06_in17 = reg_0656;
    12: op1_06_in17 = reg_0468;
    13: op1_06_in17 = reg_0250;
    14: op1_06_in17 = reg_0447;
    15: op1_06_in17 = reg_0198;
    16: op1_06_in17 = reg_0542;
    17: op1_06_in17 = reg_0215;
    18: op1_06_in17 = reg_0590;
    19: op1_06_in17 = reg_0408;
    20: op1_06_in17 = imem03_in[11:8];
    21: op1_06_in17 = reg_0348;
    22: op1_06_in17 = reg_0482;
    23: op1_06_in17 = reg_0636;
    24: op1_06_in17 = reg_1055;
    25: op1_06_in17 = imem04_in[107:104];
    26: op1_06_in17 = reg_0381;
    27: op1_06_in17 = imem04_in[119:116];
    28: op1_06_in17 = reg_0834;
    29: op1_06_in17 = reg_0886;
    30: op1_06_in17 = reg_0599;
    31: op1_06_in17 = reg_0129;
    32: op1_06_in17 = reg_0194;
    33: op1_06_in17 = imem02_in[63:60];
    34: op1_06_in17 = imem04_in[43:40];
    35: op1_06_in17 = reg_0466;
    37: op1_06_in17 = reg_0452;
    38: op1_06_in17 = reg_0193;
    39: op1_06_in17 = reg_0772;
    40: op1_06_in17 = reg_0074;
    41: op1_06_in17 = reg_0004;
    42: op1_06_in17 = reg_0723;
    43: op1_06_in17 = reg_0195;
    44: op1_06_in17 = reg_0792;
    45: op1_06_in17 = imem06_in[115:112];
    46: op1_06_in17 = reg_0158;
    47: op1_06_in17 = reg_0007;
    48: op1_06_in17 = imem05_in[111:108];
    50: op1_06_in17 = reg_0804;
    51: op1_06_in17 = reg_0955;
    52: op1_06_in17 = reg_0291;
    53: op1_06_in17 = reg_0061;
    54: op1_06_in17 = reg_0774;
    55: op1_06_in17 = reg_0926;
    56: op1_06_in17 = reg_0721;
    58: op1_06_in17 = reg_0192;
    81: op1_06_in17 = reg_0192;
    60: op1_06_in17 = imem02_in[7:4];
    61: op1_06_in17 = imem01_in[39:36];
    62: op1_06_in17 = reg_0516;
    63: op1_06_in17 = reg_1030;
    64: op1_06_in17 = reg_0611;
    67: op1_06_in17 = reg_0431;
    68: op1_06_in17 = reg_0869;
    69: op1_06_in17 = reg_0015;
    70: op1_06_in17 = imem07_in[95:92];
    71: op1_06_in17 = reg_0478;
    72: op1_06_in17 = imem07_in[55:52];
    73: op1_06_in17 = reg_0179;
    75: op1_06_in17 = reg_0106;
    76: op1_06_in17 = imem03_in[95:92];
    77: op1_06_in17 = reg_0090;
    78: op1_06_in17 = reg_0995;
    79: op1_06_in17 = reg_0619;
    83: op1_06_in17 = imem05_in[107:104];
    84: op1_06_in17 = imem02_in[127:124];
    85: op1_06_in17 = reg_0172;
    86: op1_06_in17 = reg_0458;
    87: op1_06_in17 = reg_0893;
    88: op1_06_in17 = reg_0270;
    89: op1_06_in17 = reg_0233;
    90: op1_06_in17 = reg_0420;
    93: op1_06_in17 = reg_0365;
    94: op1_06_in17 = reg_0543;
    95: op1_06_in17 = imem02_in[119:116];
    97: op1_06_in17 = imem01_in[107:104];
    default: op1_06_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv17 = 1;
    12: op1_06_inv17 = 1;
    15: op1_06_inv17 = 1;
    18: op1_06_inv17 = 1;
    19: op1_06_inv17 = 1;
    20: op1_06_inv17 = 1;
    24: op1_06_inv17 = 1;
    25: op1_06_inv17 = 1;
    26: op1_06_inv17 = 1;
    29: op1_06_inv17 = 1;
    31: op1_06_inv17 = 1;
    34: op1_06_inv17 = 1;
    38: op1_06_inv17 = 1;
    39: op1_06_inv17 = 1;
    40: op1_06_inv17 = 1;
    42: op1_06_inv17 = 1;
    43: op1_06_inv17 = 1;
    46: op1_06_inv17 = 1;
    48: op1_06_inv17 = 1;
    52: op1_06_inv17 = 1;
    53: op1_06_inv17 = 1;
    67: op1_06_inv17 = 1;
    68: op1_06_inv17 = 1;
    69: op1_06_inv17 = 1;
    72: op1_06_inv17 = 1;
    73: op1_06_inv17 = 1;
    75: op1_06_inv17 = 1;
    78: op1_06_inv17 = 1;
    79: op1_06_inv17 = 1;
    86: op1_06_inv17 = 1;
    88: op1_06_inv17 = 1;
    89: op1_06_inv17 = 1;
    90: op1_06_inv17 = 1;
    93: op1_06_inv17 = 1;
    97: op1_06_inv17 = 1;
    default: op1_06_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in18 = reg_0346;
    6: op1_06_in18 = imem01_in[103:100];
    7: op1_06_in18 = reg_0043;
    8: op1_06_in18 = reg_0167;
    9: op1_06_in18 = reg_0326;
    10: op1_06_in18 = reg_0792;
    11: op1_06_in18 = reg_0662;
    12: op1_06_in18 = reg_0478;
    13: op1_06_in18 = reg_0836;
    17: op1_06_in18 = reg_0836;
    14: op1_06_in18 = reg_0445;
    15: op1_06_in18 = reg_0212;
    16: op1_06_in18 = reg_0558;
    18: op1_06_in18 = reg_0395;
    19: op1_06_in18 = reg_0351;
    20: op1_06_in18 = imem03_in[31:28];
    21: op1_06_in18 = reg_0356;
    22: op1_06_in18 = reg_0814;
    44: op1_06_in18 = reg_0814;
    23: op1_06_in18 = reg_0663;
    24: op1_06_in18 = reg_0246;
    25: op1_06_in18 = imem04_in[127:124];
    27: op1_06_in18 = imem04_in[127:124];
    26: op1_06_in18 = reg_0392;
    28: op1_06_in18 = reg_0826;
    29: op1_06_in18 = reg_0037;
    30: op1_06_in18 = reg_0583;
    31: op1_06_in18 = reg_0141;
    32: op1_06_in18 = reg_0198;
    33: op1_06_in18 = imem02_in[95:92];
    34: op1_06_in18 = imem04_in[115:112];
    35: op1_06_in18 = reg_0472;
    37: op1_06_in18 = reg_0456;
    38: op1_06_in18 = reg_0194;
    71: op1_06_in18 = reg_0194;
    39: op1_06_in18 = reg_0088;
    40: op1_06_in18 = reg_0059;
    41: op1_06_in18 = reg_0765;
    42: op1_06_in18 = reg_0725;
    43: op1_06_in18 = imem01_in[11:8];
    45: op1_06_in18 = reg_0020;
    47: op1_06_in18 = reg_0089;
    48: op1_06_in18 = imem05_in[123:120];
    50: op1_06_in18 = reg_0349;
    51: op1_06_in18 = reg_0964;
    52: op1_06_in18 = reg_0079;
    53: op1_06_in18 = reg_0554;
    54: op1_06_in18 = reg_0493;
    55: op1_06_in18 = imem07_in[3:0];
    56: op1_06_in18 = reg_0723;
    58: op1_06_in18 = imem01_in[19:16];
    60: op1_06_in18 = imem02_in[15:12];
    61: op1_06_in18 = imem01_in[43:40];
    62: op1_06_in18 = reg_0007;
    63: op1_06_in18 = reg_0297;
    64: op1_06_in18 = reg_0380;
    67: op1_06_in18 = reg_0174;
    68: op1_06_in18 = reg_1043;
    69: op1_06_in18 = reg_0732;
    70: op1_06_in18 = imem07_in[107:104];
    72: op1_06_in18 = imem07_in[71:68];
    73: op1_06_in18 = reg_0161;
    75: op1_06_in18 = reg_0973;
    76: op1_06_in18 = reg_0322;
    77: op1_06_in18 = imem03_in[39:36];
    78: op1_06_in18 = reg_0979;
    79: op1_06_in18 = reg_0857;
    81: op1_06_in18 = imem01_in[3:0];
    83: op1_06_in18 = imem05_in[119:116];
    84: op1_06_in18 = reg_0645;
    85: op1_06_in18 = reg_0179;
    86: op1_06_in18 = reg_0214;
    87: op1_06_in18 = reg_0432;
    88: op1_06_in18 = reg_0915;
    89: op1_06_in18 = reg_0998;
    90: op1_06_in18 = reg_0024;
    93: op1_06_in18 = reg_0367;
    94: op1_06_in18 = reg_0639;
    95: op1_06_in18 = imem02_in[127:124];
    96: op1_06_in18 = reg_0788;
    97: op1_06_in18 = imem01_in[111:108];
    default: op1_06_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv18 = 1;
    6: op1_06_inv18 = 1;
    9: op1_06_inv18 = 1;
    11: op1_06_inv18 = 1;
    12: op1_06_inv18 = 1;
    14: op1_06_inv18 = 1;
    15: op1_06_inv18 = 1;
    16: op1_06_inv18 = 1;
    19: op1_06_inv18 = 1;
    20: op1_06_inv18 = 1;
    21: op1_06_inv18 = 1;
    24: op1_06_inv18 = 1;
    25: op1_06_inv18 = 1;
    26: op1_06_inv18 = 1;
    29: op1_06_inv18 = 1;
    30: op1_06_inv18 = 1;
    31: op1_06_inv18 = 1;
    33: op1_06_inv18 = 1;
    34: op1_06_inv18 = 1;
    35: op1_06_inv18 = 1;
    39: op1_06_inv18 = 1;
    41: op1_06_inv18 = 1;
    42: op1_06_inv18 = 1;
    43: op1_06_inv18 = 1;
    44: op1_06_inv18 = 1;
    51: op1_06_inv18 = 1;
    52: op1_06_inv18 = 1;
    56: op1_06_inv18 = 1;
    58: op1_06_inv18 = 1;
    60: op1_06_inv18 = 1;
    61: op1_06_inv18 = 1;
    62: op1_06_inv18 = 1;
    63: op1_06_inv18 = 1;
    67: op1_06_inv18 = 1;
    69: op1_06_inv18 = 1;
    72: op1_06_inv18 = 1;
    73: op1_06_inv18 = 1;
    75: op1_06_inv18 = 1;
    77: op1_06_inv18 = 1;
    81: op1_06_inv18 = 1;
    86: op1_06_inv18 = 1;
    88: op1_06_inv18 = 1;
    89: op1_06_inv18 = 1;
    90: op1_06_inv18 = 1;
    96: op1_06_inv18 = 1;
    default: op1_06_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in19 = reg_0347;
    6: op1_06_in19 = reg_0500;
    7: op1_06_in19 = reg_0053;
    8: op1_06_in19 = reg_0169;
    9: op1_06_in19 = reg_0329;
    10: op1_06_in19 = reg_0219;
    11: op1_06_in19 = reg_0358;
    12: op1_06_in19 = reg_0204;
    13: op1_06_in19 = reg_0865;
    17: op1_06_in19 = reg_0865;
    14: op1_06_in19 = reg_0428;
    15: op1_06_in19 = reg_0190;
    16: op1_06_in19 = reg_0533;
    18: op1_06_in19 = reg_0384;
    19: op1_06_in19 = reg_0405;
    20: op1_06_in19 = imem03_in[55:52];
    21: op1_06_in19 = reg_0382;
    63: op1_06_in19 = reg_0382;
    22: op1_06_in19 = imem03_in[59:56];
    23: op1_06_in19 = reg_0352;
    24: op1_06_in19 = reg_1043;
    25: op1_06_in19 = reg_1003;
    26: op1_06_in19 = reg_0383;
    27: op1_06_in19 = reg_0483;
    28: op1_06_in19 = reg_0757;
    29: op1_06_in19 = reg_0335;
    30: op1_06_in19 = reg_0592;
    31: op1_06_in19 = imem06_in[47:44];
    32: op1_06_in19 = imem01_in[31:28];
    43: op1_06_in19 = imem01_in[31:28];
    58: op1_06_in19 = imem01_in[31:28];
    33: op1_06_in19 = imem02_in[107:104];
    34: op1_06_in19 = reg_0541;
    35: op1_06_in19 = reg_0470;
    37: op1_06_in19 = reg_0187;
    38: op1_06_in19 = reg_0201;
    39: op1_06_in19 = reg_0876;
    40: op1_06_in19 = reg_0054;
    41: op1_06_in19 = reg_0795;
    42: op1_06_in19 = reg_0703;
    44: op1_06_in19 = reg_0086;
    45: op1_06_in19 = reg_0556;
    47: op1_06_in19 = reg_0814;
    48: op1_06_in19 = reg_0963;
    50: op1_06_in19 = reg_0332;
    51: op1_06_in19 = reg_0968;
    52: op1_06_in19 = imem03_in[7:4];
    53: op1_06_in19 = reg_0528;
    54: op1_06_in19 = reg_0094;
    55: op1_06_in19 = imem07_in[19:16];
    56: op1_06_in19 = reg_0717;
    60: op1_06_in19 = imem02_in[27:24];
    61: op1_06_in19 = imem01_in[91:88];
    62: op1_06_in19 = reg_0776;
    64: op1_06_in19 = reg_0619;
    67: op1_06_in19 = reg_0172;
    68: op1_06_in19 = reg_0113;
    69: op1_06_in19 = reg_0432;
    70: op1_06_in19 = imem07_in[111:108];
    71: op1_06_in19 = imem01_in[11:8];
    72: op1_06_in19 = imem07_in[123:120];
    73: op1_06_in19 = reg_0167;
    75: op1_06_in19 = reg_0793;
    76: op1_06_in19 = reg_0547;
    77: op1_06_in19 = imem03_in[71:68];
    78: op1_06_in19 = reg_0984;
    79: op1_06_in19 = reg_0220;
    81: op1_06_in19 = imem01_in[7:4];
    83: op1_06_in19 = reg_1021;
    84: op1_06_in19 = reg_0664;
    85: op1_06_in19 = reg_0185;
    86: op1_06_in19 = reg_0191;
    87: op1_06_in19 = reg_0517;
    88: op1_06_in19 = reg_0755;
    89: op1_06_in19 = reg_0995;
    90: op1_06_in19 = reg_0179;
    93: op1_06_in19 = imem03_in[31:28];
    94: op1_06_in19 = reg_0887;
    95: op1_06_in19 = reg_0277;
    96: op1_06_in19 = reg_0493;
    97: op1_06_in19 = reg_0798;
    default: op1_06_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv19 = 1;
    8: op1_06_inv19 = 1;
    9: op1_06_inv19 = 1;
    10: op1_06_inv19 = 1;
    12: op1_06_inv19 = 1;
    13: op1_06_inv19 = 1;
    15: op1_06_inv19 = 1;
    19: op1_06_inv19 = 1;
    20: op1_06_inv19 = 1;
    21: op1_06_inv19 = 1;
    24: op1_06_inv19 = 1;
    25: op1_06_inv19 = 1;
    26: op1_06_inv19 = 1;
    29: op1_06_inv19 = 1;
    37: op1_06_inv19 = 1;
    39: op1_06_inv19 = 1;
    40: op1_06_inv19 = 1;
    41: op1_06_inv19 = 1;
    44: op1_06_inv19 = 1;
    53: op1_06_inv19 = 1;
    54: op1_06_inv19 = 1;
    56: op1_06_inv19 = 1;
    60: op1_06_inv19 = 1;
    61: op1_06_inv19 = 1;
    62: op1_06_inv19 = 1;
    67: op1_06_inv19 = 1;
    71: op1_06_inv19 = 1;
    77: op1_06_inv19 = 1;
    79: op1_06_inv19 = 1;
    83: op1_06_inv19 = 1;
    84: op1_06_inv19 = 1;
    85: op1_06_inv19 = 1;
    86: op1_06_inv19 = 1;
    88: op1_06_inv19 = 1;
    94: op1_06_inv19 = 1;
    96: op1_06_inv19 = 1;
    97: op1_06_inv19 = 1;
    default: op1_06_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in20 = reg_0092;
    6: op1_06_in20 = reg_0519;
    7: op1_06_in20 = reg_0071;
    8: op1_06_in20 = reg_0160;
    9: op1_06_in20 = reg_0339;
    10: op1_06_in20 = reg_0225;
    11: op1_06_in20 = reg_0353;
    12: op1_06_in20 = reg_0198;
    13: op1_06_in20 = reg_0896;
    14: op1_06_in20 = reg_0444;
    15: op1_06_in20 = reg_0197;
    16: op1_06_in20 = reg_0531;
    17: op1_06_in20 = reg_0828;
    18: op1_06_in20 = reg_0360;
    19: op1_06_in20 = reg_0371;
    20: op1_06_in20 = imem03_in[103:100];
    21: op1_06_in20 = reg_0315;
    22: op1_06_in20 = imem03_in[91:88];
    23: op1_06_in20 = reg_0364;
    24: op1_06_in20 = reg_0122;
    25: op1_06_in20 = reg_0937;
    26: op1_06_in20 = reg_0404;
    27: op1_06_in20 = reg_0301;
    28: op1_06_in20 = reg_0491;
    29: op1_06_in20 = reg_0876;
    30: op1_06_in20 = reg_0591;
    31: op1_06_in20 = imem06_in[63:60];
    32: op1_06_in20 = imem01_in[35:32];
    58: op1_06_in20 = imem01_in[35:32];
    33: op1_06_in20 = reg_0661;
    34: op1_06_in20 = reg_0733;
    35: op1_06_in20 = reg_0474;
    37: op1_06_in20 = reg_0203;
    38: op1_06_in20 = reg_0190;
    39: op1_06_in20 = reg_0792;
    40: op1_06_in20 = reg_0528;
    41: op1_06_in20 = reg_0369;
    88: op1_06_in20 = reg_0369;
    42: op1_06_in20 = reg_0729;
    43: op1_06_in20 = imem01_in[43:40];
    44: op1_06_in20 = imem03_in[11:8];
    45: op1_06_in20 = reg_0619;
    47: op1_06_in20 = reg_0090;
    48: op1_06_in20 = reg_0973;
    50: op1_06_in20 = reg_0630;
    51: op1_06_in20 = reg_0945;
    52: op1_06_in20 = imem03_in[75:72];
    53: op1_06_in20 = reg_0043;
    54: op1_06_in20 = reg_0448;
    55: op1_06_in20 = imem07_in[27:24];
    56: op1_06_in20 = reg_0725;
    60: op1_06_in20 = imem02_in[35:32];
    61: op1_06_in20 = imem01_in[123:120];
    62: op1_06_in20 = reg_0085;
    63: op1_06_in20 = reg_0222;
    64: op1_06_in20 = reg_0257;
    67: op1_06_in20 = reg_0179;
    68: op1_06_in20 = reg_0821;
    69: op1_06_in20 = reg_0409;
    70: op1_06_in20 = reg_0718;
    71: op1_06_in20 = imem01_in[67:64];
    72: op1_06_in20 = reg_0721;
    75: op1_06_in20 = reg_0862;
    76: op1_06_in20 = reg_0571;
    77: op1_06_in20 = imem03_in[87:84];
    78: op1_06_in20 = imem04_in[75:72];
    79: op1_06_in20 = reg_0612;
    81: op1_06_in20 = imem01_in[31:28];
    83: op1_06_in20 = reg_0319;
    84: op1_06_in20 = reg_0423;
    86: op1_06_in20 = reg_0210;
    87: op1_06_in20 = reg_0777;
    89: op1_06_in20 = reg_1001;
    90: op1_06_in20 = reg_0714;
    93: op1_06_in20 = imem03_in[67:64];
    94: op1_06_in20 = reg_0855;
    95: op1_06_in20 = reg_0073;
    96: op1_06_in20 = imem03_in[31:28];
    97: op1_06_in20 = reg_0246;
    default: op1_06_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv20 = 1;
    8: op1_06_inv20 = 1;
    9: op1_06_inv20 = 1;
    10: op1_06_inv20 = 1;
    12: op1_06_inv20 = 1;
    13: op1_06_inv20 = 1;
    16: op1_06_inv20 = 1;
    18: op1_06_inv20 = 1;
    19: op1_06_inv20 = 1;
    21: op1_06_inv20 = 1;
    23: op1_06_inv20 = 1;
    25: op1_06_inv20 = 1;
    27: op1_06_inv20 = 1;
    30: op1_06_inv20 = 1;
    32: op1_06_inv20 = 1;
    33: op1_06_inv20 = 1;
    37: op1_06_inv20 = 1;
    38: op1_06_inv20 = 1;
    39: op1_06_inv20 = 1;
    41: op1_06_inv20 = 1;
    48: op1_06_inv20 = 1;
    52: op1_06_inv20 = 1;
    60: op1_06_inv20 = 1;
    72: op1_06_inv20 = 1;
    76: op1_06_inv20 = 1;
    77: op1_06_inv20 = 1;
    78: op1_06_inv20 = 1;
    81: op1_06_inv20 = 1;
    86: op1_06_inv20 = 1;
    87: op1_06_inv20 = 1;
    89: op1_06_inv20 = 1;
    90: op1_06_inv20 = 1;
    95: op1_06_inv20 = 1;
    97: op1_06_inv20 = 1;
    default: op1_06_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in21 = reg_0051;
    6: op1_06_in21 = reg_0499;
    7: op1_06_in21 = reg_0064;
    8: op1_06_in21 = reg_0166;
    9: op1_06_in21 = reg_0355;
    10: op1_06_in21 = reg_0522;
    11: op1_06_in21 = reg_0342;
    12: op1_06_in21 = reg_0205;
    13: op1_06_in21 = reg_0894;
    14: op1_06_in21 = reg_0442;
    15: op1_06_in21 = imem01_in[27:24];
    16: op1_06_in21 = reg_0305;
    17: op1_06_in21 = reg_0255;
    18: op1_06_in21 = reg_0370;
    19: op1_06_in21 = reg_0313;
    20: op1_06_in21 = imem03_in[127:124];
    21: op1_06_in21 = reg_0808;
    22: op1_06_in21 = reg_0582;
    23: op1_06_in21 = reg_0339;
    24: op1_06_in21 = reg_0125;
    25: op1_06_in21 = reg_0277;
    26: op1_06_in21 = reg_0368;
    27: op1_06_in21 = reg_0530;
    28: op1_06_in21 = reg_0260;
    29: op1_06_in21 = reg_0291;
    30: op1_06_in21 = reg_0589;
    31: op1_06_in21 = imem06_in[115:112];
    32: op1_06_in21 = imem01_in[43:40];
    33: op1_06_in21 = reg_0639;
    34: op1_06_in21 = reg_0763;
    35: op1_06_in21 = reg_0459;
    37: op1_06_in21 = reg_0207;
    38: op1_06_in21 = imem01_in[11:8];
    39: op1_06_in21 = imem03_in[35:32];
    40: op1_06_in21 = reg_0517;
    41: op1_06_in21 = reg_0377;
    42: op1_06_in21 = reg_0718;
    43: op1_06_in21 = imem01_in[47:44];
    44: op1_06_in21 = imem03_in[27:24];
    45: op1_06_in21 = reg_0632;
    47: op1_06_in21 = reg_0084;
    48: op1_06_in21 = reg_0968;
    50: op1_06_in21 = reg_0241;
    51: op1_06_in21 = reg_0952;
    52: op1_06_in21 = imem03_in[87:84];
    93: op1_06_in21 = imem03_in[87:84];
    53: op1_06_in21 = reg_0429;
    54: op1_06_in21 = reg_0404;
    55: op1_06_in21 = imem07_in[43:40];
    56: op1_06_in21 = reg_0709;
    58: op1_06_in21 = imem01_in[39:36];
    60: op1_06_in21 = imem02_in[75:72];
    61: op1_06_in21 = reg_0936;
    62: op1_06_in21 = imem03_in[43:40];
    63: op1_06_in21 = reg_1029;
    64: op1_06_in21 = reg_0630;
    67: op1_06_in21 = reg_0160;
    68: op1_06_in21 = reg_0110;
    69: op1_06_in21 = reg_0824;
    70: op1_06_in21 = reg_0002;
    71: op1_06_in21 = imem01_in[75:72];
    72: op1_06_in21 = reg_0717;
    75: op1_06_in21 = reg_1031;
    76: op1_06_in21 = reg_0767;
    77: op1_06_in21 = imem03_in[107:104];
    78: op1_06_in21 = imem04_in[83:80];
    79: op1_06_in21 = reg_0915;
    81: op1_06_in21 = imem01_in[55:52];
    83: op1_06_in21 = reg_0143;
    84: op1_06_in21 = reg_0394;
    86: op1_06_in21 = imem01_in[3:0];
    87: op1_06_in21 = reg_0020;
    88: op1_06_in21 = imem07_in[7:4];
    89: op1_06_in21 = reg_0997;
    90: op1_06_in21 = reg_0184;
    94: op1_06_in21 = reg_0645;
    95: op1_06_in21 = reg_0095;
    96: op1_06_in21 = imem03_in[63:60];
    97: op1_06_in21 = reg_0070;
    default: op1_06_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv21 = 1;
    8: op1_06_inv21 = 1;
    9: op1_06_inv21 = 1;
    10: op1_06_inv21 = 1;
    12: op1_06_inv21 = 1;
    13: op1_06_inv21 = 1;
    14: op1_06_inv21 = 1;
    15: op1_06_inv21 = 1;
    16: op1_06_inv21 = 1;
    17: op1_06_inv21 = 1;
    20: op1_06_inv21 = 1;
    22: op1_06_inv21 = 1;
    23: op1_06_inv21 = 1;
    25: op1_06_inv21 = 1;
    27: op1_06_inv21 = 1;
    28: op1_06_inv21 = 1;
    30: op1_06_inv21 = 1;
    34: op1_06_inv21 = 1;
    35: op1_06_inv21 = 1;
    37: op1_06_inv21 = 1;
    38: op1_06_inv21 = 1;
    40: op1_06_inv21 = 1;
    42: op1_06_inv21 = 1;
    43: op1_06_inv21 = 1;
    44: op1_06_inv21 = 1;
    47: op1_06_inv21 = 1;
    48: op1_06_inv21 = 1;
    50: op1_06_inv21 = 1;
    51: op1_06_inv21 = 1;
    54: op1_06_inv21 = 1;
    56: op1_06_inv21 = 1;
    62: op1_06_inv21 = 1;
    63: op1_06_inv21 = 1;
    68: op1_06_inv21 = 1;
    69: op1_06_inv21 = 1;
    72: op1_06_inv21 = 1;
    77: op1_06_inv21 = 1;
    83: op1_06_inv21 = 1;
    86: op1_06_inv21 = 1;
    96: op1_06_inv21 = 1;
    97: op1_06_inv21 = 1;
    default: op1_06_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in22 = reg_0084;
    6: op1_06_in22 = reg_0507;
    7: op1_06_in22 = reg_0050;
    8: op1_06_in22 = reg_0177;
    67: op1_06_in22 = reg_0177;
    9: op1_06_in22 = reg_0097;
    10: op1_06_in22 = reg_0520;
    11: op1_06_in22 = reg_0082;
    12: op1_06_in22 = reg_0202;
    13: op1_06_in22 = reg_0132;
    14: op1_06_in22 = reg_0175;
    15: op1_06_in22 = imem01_in[35:32];
    16: op1_06_in22 = reg_0290;
    17: op1_06_in22 = reg_0832;
    18: op1_06_in22 = reg_0312;
    19: op1_06_in22 = reg_0406;
    20: op1_06_in22 = reg_0586;
    21: op1_06_in22 = reg_0017;
    50: op1_06_in22 = reg_0017;
    22: op1_06_in22 = reg_0599;
    23: op1_06_in22 = reg_0776;
    24: op1_06_in22 = reg_0108;
    25: op1_06_in22 = reg_0282;
    26: op1_06_in22 = reg_1029;
    27: op1_06_in22 = reg_0277;
    28: op1_06_in22 = reg_0785;
    29: op1_06_in22 = imem03_in[39:36];
    30: op1_06_in22 = reg_0593;
    31: op1_06_in22 = reg_0625;
    32: op1_06_in22 = imem01_in[111:108];
    33: op1_06_in22 = reg_0651;
    34: op1_06_in22 = reg_0296;
    35: op1_06_in22 = reg_0478;
    37: op1_06_in22 = reg_0211;
    38: op1_06_in22 = imem01_in[15:12];
    39: op1_06_in22 = imem03_in[63:60];
    62: op1_06_in22 = imem03_in[63:60];
    40: op1_06_in22 = reg_0855;
    41: op1_06_in22 = reg_0767;
    42: op1_06_in22 = reg_0449;
    43: op1_06_in22 = imem01_in[59:56];
    58: op1_06_in22 = imem01_in[59:56];
    44: op1_06_in22 = imem03_in[75:72];
    45: op1_06_in22 = reg_0612;
    47: op1_06_in22 = reg_0016;
    48: op1_06_in22 = reg_0961;
    51: op1_06_in22 = reg_0953;
    52: op1_06_in22 = reg_1008;
    53: op1_06_in22 = reg_0777;
    54: op1_06_in22 = reg_0447;
    55: op1_06_in22 = imem07_in[51:48];
    56: op1_06_in22 = reg_0705;
    60: op1_06_in22 = imem02_in[83:80];
    61: op1_06_in22 = reg_1044;
    63: op1_06_in22 = reg_0946;
    64: op1_06_in22 = reg_0408;
    68: op1_06_in22 = imem02_in[3:0];
    69: op1_06_in22 = reg_0542;
    70: op1_06_in22 = reg_0353;
    71: op1_06_in22 = reg_0969;
    97: op1_06_in22 = reg_0969;
    72: op1_06_in22 = reg_0729;
    75: op1_06_in22 = reg_0737;
    76: op1_06_in22 = reg_0233;
    77: op1_06_in22 = reg_0620;
    78: op1_06_in22 = imem04_in[87:84];
    79: op1_06_in22 = reg_0755;
    81: op1_06_in22 = imem01_in[63:60];
    83: op1_06_in22 = reg_0365;
    84: op1_06_in22 = reg_0248;
    86: op1_06_in22 = imem01_in[55:52];
    87: op1_06_in22 = reg_0673;
    88: op1_06_in22 = imem07_in[19:16];
    89: op1_06_in22 = imem04_in[3:0];
    93: op1_06_in22 = imem03_in[95:92];
    94: op1_06_in22 = reg_0664;
    95: op1_06_in22 = reg_0279;
    96: op1_06_in22 = reg_0631;
    default: op1_06_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_06_inv22 = 1;
    10: op1_06_inv22 = 1;
    12: op1_06_inv22 = 1;
    14: op1_06_inv22 = 1;
    15: op1_06_inv22 = 1;
    20: op1_06_inv22 = 1;
    21: op1_06_inv22 = 1;
    25: op1_06_inv22 = 1;
    26: op1_06_inv22 = 1;
    31: op1_06_inv22 = 1;
    32: op1_06_inv22 = 1;
    33: op1_06_inv22 = 1;
    34: op1_06_inv22 = 1;
    39: op1_06_inv22 = 1;
    43: op1_06_inv22 = 1;
    47: op1_06_inv22 = 1;
    51: op1_06_inv22 = 1;
    52: op1_06_inv22 = 1;
    53: op1_06_inv22 = 1;
    58: op1_06_inv22 = 1;
    60: op1_06_inv22 = 1;
    61: op1_06_inv22 = 1;
    63: op1_06_inv22 = 1;
    64: op1_06_inv22 = 1;
    68: op1_06_inv22 = 1;
    72: op1_06_inv22 = 1;
    75: op1_06_inv22 = 1;
    76: op1_06_inv22 = 1;
    81: op1_06_inv22 = 1;
    83: op1_06_inv22 = 1;
    84: op1_06_inv22 = 1;
    87: op1_06_inv22 = 1;
    88: op1_06_inv22 = 1;
    89: op1_06_inv22 = 1;
    93: op1_06_inv22 = 1;
    96: op1_06_inv22 = 1;
    default: op1_06_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in23 = reg_0093;
    6: op1_06_in23 = reg_0235;
    7: op1_06_in23 = imem05_in[91:88];
    8: op1_06_in23 = reg_0185;
    9: op1_06_in23 = reg_0091;
    10: op1_06_in23 = reg_0514;
    11: op1_06_in23 = reg_0073;
    12: op1_06_in23 = reg_0195;
    13: op1_06_in23 = reg_0148;
    17: op1_06_in23 = reg_0148;
    14: op1_06_in23 = reg_0169;
    15: op1_06_in23 = imem01_in[39:36];
    16: op1_06_in23 = reg_0295;
    69: op1_06_in23 = reg_0295;
    18: op1_06_in23 = reg_1002;
    19: op1_06_in23 = reg_0799;
    20: op1_06_in23 = reg_0579;
    22: op1_06_in23 = reg_0579;
    21: op1_06_in23 = reg_0803;
    23: op1_06_in23 = imem03_in[7:4];
    24: op1_06_in23 = imem02_in[15:12];
    25: op1_06_in23 = reg_0048;
    26: op1_06_in23 = reg_1028;
    27: op1_06_in23 = reg_0537;
    28: op1_06_in23 = reg_0896;
    29: op1_06_in23 = imem03_in[63:60];
    30: op1_06_in23 = reg_0595;
    31: op1_06_in23 = reg_0604;
    32: op1_06_in23 = imem01_in[119:116];
    33: op1_06_in23 = reg_0647;
    34: op1_06_in23 = reg_0074;
    35: op1_06_in23 = reg_0200;
    37: op1_06_in23 = reg_0194;
    38: op1_06_in23 = imem01_in[19:16];
    39: op1_06_in23 = reg_0343;
    40: op1_06_in23 = reg_0044;
    41: op1_06_in23 = reg_0820;
    42: op1_06_in23 = reg_0444;
    43: op1_06_in23 = imem01_in[103:100];
    44: op1_06_in23 = imem03_in[91:88];
    45: op1_06_in23 = reg_0387;
    47: op1_06_in23 = imem03_in[39:36];
    48: op1_06_in23 = reg_0900;
    50: op1_06_in23 = reg_0609;
    51: op1_06_in23 = reg_0972;
    52: op1_06_in23 = reg_0580;
    53: op1_06_in23 = reg_0070;
    54: op1_06_in23 = reg_0269;
    55: op1_06_in23 = imem07_in[55:52];
    56: op1_06_in23 = reg_0707;
    72: op1_06_in23 = reg_0707;
    58: op1_06_in23 = imem01_in[87:84];
    60: op1_06_in23 = reg_0642;
    61: op1_06_in23 = reg_0242;
    62: op1_06_in23 = imem03_in[95:92];
    63: op1_06_in23 = reg_0408;
    64: op1_06_in23 = reg_0780;
    67: op1_06_in23 = reg_0157;
    68: op1_06_in23 = imem02_in[19:16];
    70: op1_06_in23 = reg_0589;
    71: op1_06_in23 = reg_1044;
    75: op1_06_in23 = reg_0740;
    76: op1_06_in23 = reg_0987;
    77: op1_06_in23 = reg_1007;
    78: op1_06_in23 = imem04_in[111:108];
    79: op1_06_in23 = reg_0730;
    81: op1_06_in23 = reg_0105;
    83: op1_06_in23 = reg_0314;
    84: op1_06_in23 = reg_0087;
    86: op1_06_in23 = imem01_in[83:80];
    87: op1_06_in23 = reg_0946;
    88: op1_06_in23 = imem07_in[31:28];
    89: op1_06_in23 = reg_0395;
    93: op1_06_in23 = imem03_in[107:104];
    94: op1_06_in23 = reg_0394;
    95: op1_06_in23 = reg_0358;
    96: op1_06_in23 = reg_0761;
    97: op1_06_in23 = reg_0222;
    default: op1_06_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv23 = 1;
    7: op1_06_inv23 = 1;
    8: op1_06_inv23 = 1;
    9: op1_06_inv23 = 1;
    10: op1_06_inv23 = 1;
    12: op1_06_inv23 = 1;
    14: op1_06_inv23 = 1;
    15: op1_06_inv23 = 1;
    16: op1_06_inv23 = 1;
    19: op1_06_inv23 = 1;
    20: op1_06_inv23 = 1;
    23: op1_06_inv23 = 1;
    24: op1_06_inv23 = 1;
    25: op1_06_inv23 = 1;
    28: op1_06_inv23 = 1;
    30: op1_06_inv23 = 1;
    32: op1_06_inv23 = 1;
    33: op1_06_inv23 = 1;
    35: op1_06_inv23 = 1;
    37: op1_06_inv23 = 1;
    38: op1_06_inv23 = 1;
    41: op1_06_inv23 = 1;
    42: op1_06_inv23 = 1;
    48: op1_06_inv23 = 1;
    51: op1_06_inv23 = 1;
    53: op1_06_inv23 = 1;
    54: op1_06_inv23 = 1;
    58: op1_06_inv23 = 1;
    60: op1_06_inv23 = 1;
    62: op1_06_inv23 = 1;
    64: op1_06_inv23 = 1;
    67: op1_06_inv23 = 1;
    68: op1_06_inv23 = 1;
    72: op1_06_inv23 = 1;
    75: op1_06_inv23 = 1;
    76: op1_06_inv23 = 1;
    78: op1_06_inv23 = 1;
    79: op1_06_inv23 = 1;
    84: op1_06_inv23 = 1;
    86: op1_06_inv23 = 1;
    87: op1_06_inv23 = 1;
    89: op1_06_inv23 = 1;
    93: op1_06_inv23 = 1;
    96: op1_06_inv23 = 1;
    97: op1_06_inv23 = 1;
    default: op1_06_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in24 = imem03_in[59:56];
    6: op1_06_in24 = reg_0222;
    7: op1_06_in24 = imem05_in[99:96];
    8: op1_06_in24 = reg_0168;
    9: op1_06_in24 = reg_0084;
    10: op1_06_in24 = reg_0521;
    11: op1_06_in24 = imem03_in[3:0];
    12: op1_06_in24 = reg_0199;
    13: op1_06_in24 = reg_0154;
    14: op1_06_in24 = reg_0163;
    15: op1_06_in24 = imem01_in[55:52];
    16: op1_06_in24 = reg_0059;
    17: op1_06_in24 = reg_0152;
    18: op1_06_in24 = reg_0974;
    19: op1_06_in24 = reg_0787;
    20: op1_06_in24 = reg_0585;
    21: op1_06_in24 = reg_0754;
    22: op1_06_in24 = reg_0572;
    23: op1_06_in24 = imem03_in[43:40];
    24: op1_06_in24 = imem02_in[31:28];
    25: op1_06_in24 = reg_1057;
    26: op1_06_in24 = reg_0017;
    27: op1_06_in24 = reg_0313;
    28: op1_06_in24 = reg_0497;
    29: op1_06_in24 = imem03_in[87:84];
    30: op1_06_in24 = reg_0588;
    31: op1_06_in24 = reg_0605;
    32: op1_06_in24 = imem01_in[123:120];
    33: op1_06_in24 = reg_0638;
    34: op1_06_in24 = reg_0064;
    35: op1_06_in24 = reg_0193;
    37: op1_06_in24 = imem01_in[23:20];
    38: op1_06_in24 = imem01_in[43:40];
    39: op1_06_in24 = reg_0938;
    40: op1_06_in24 = imem05_in[7:4];
    41: op1_06_in24 = reg_0984;
    42: op1_06_in24 = reg_0442;
    43: op1_06_in24 = imem01_in[127:124];
    44: op1_06_in24 = reg_0571;
    45: op1_06_in24 = reg_0344;
    47: op1_06_in24 = imem03_in[47:44];
    48: op1_06_in24 = reg_0260;
    50: op1_06_in24 = reg_0633;
    51: op1_06_in24 = reg_0259;
    52: op1_06_in24 = reg_0396;
    53: op1_06_in24 = reg_0864;
    54: op1_06_in24 = reg_0147;
    55: op1_06_in24 = imem07_in[83:80];
    56: op1_06_in24 = reg_0701;
    58: op1_06_in24 = imem01_in[95:92];
    60: op1_06_in24 = reg_0657;
    61: op1_06_in24 = reg_0933;
    62: op1_06_in24 = imem03_in[107:104];
    63: op1_06_in24 = reg_0241;
    64: op1_06_in24 = reg_0241;
    68: op1_06_in24 = imem02_in[79:76];
    69: op1_06_in24 = reg_0531;
    70: op1_06_in24 = reg_0172;
    71: op1_06_in24 = reg_0120;
    81: op1_06_in24 = reg_0120;
    72: op1_06_in24 = reg_0706;
    75: op1_06_in24 = reg_1017;
    76: op1_06_in24 = reg_0998;
    77: op1_06_in24 = reg_0445;
    78: op1_06_in24 = imem04_in[115:112];
    79: op1_06_in24 = reg_0158;
    83: op1_06_in24 = reg_0948;
    84: op1_06_in24 = reg_0335;
    86: op1_06_in24 = imem01_in[107:104];
    87: op1_06_in24 = reg_0319;
    88: op1_06_in24 = imem07_in[35:32];
    89: op1_06_in24 = reg_0511;
    93: op1_06_in24 = imem03_in[119:116];
    94: op1_06_in24 = reg_0248;
    95: op1_06_in24 = reg_0739;
    96: op1_06_in24 = reg_0578;
    97: op1_06_in24 = reg_0604;
    default: op1_06_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv24 = 1;
    7: op1_06_inv24 = 1;
    8: op1_06_inv24 = 1;
    9: op1_06_inv24 = 1;
    13: op1_06_inv24 = 1;
    18: op1_06_inv24 = 1;
    20: op1_06_inv24 = 1;
    21: op1_06_inv24 = 1;
    22: op1_06_inv24 = 1;
    23: op1_06_inv24 = 1;
    24: op1_06_inv24 = 1;
    26: op1_06_inv24 = 1;
    28: op1_06_inv24 = 1;
    29: op1_06_inv24 = 1;
    30: op1_06_inv24 = 1;
    31: op1_06_inv24 = 1;
    32: op1_06_inv24 = 1;
    33: op1_06_inv24 = 1;
    34: op1_06_inv24 = 1;
    40: op1_06_inv24 = 1;
    41: op1_06_inv24 = 1;
    42: op1_06_inv24 = 1;
    44: op1_06_inv24 = 1;
    47: op1_06_inv24 = 1;
    50: op1_06_inv24 = 1;
    52: op1_06_inv24 = 1;
    53: op1_06_inv24 = 1;
    54: op1_06_inv24 = 1;
    56: op1_06_inv24 = 1;
    58: op1_06_inv24 = 1;
    60: op1_06_inv24 = 1;
    61: op1_06_inv24 = 1;
    70: op1_06_inv24 = 1;
    75: op1_06_inv24 = 1;
    76: op1_06_inv24 = 1;
    77: op1_06_inv24 = 1;
    78: op1_06_inv24 = 1;
    79: op1_06_inv24 = 1;
    81: op1_06_inv24 = 1;
    83: op1_06_inv24 = 1;
    86: op1_06_inv24 = 1;
    87: op1_06_inv24 = 1;
    88: op1_06_inv24 = 1;
    89: op1_06_inv24 = 1;
    93: op1_06_inv24 = 1;
    94: op1_06_inv24 = 1;
    95: op1_06_inv24 = 1;
    96: op1_06_inv24 = 1;
    97: op1_06_inv24 = 1;
    default: op1_06_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in25 = imem03_in[95:92];
    23: op1_06_in25 = imem03_in[95:92];
    6: op1_06_in25 = reg_0240;
    7: op1_06_in25 = imem05_in[123:120];
    9: op1_06_in25 = reg_0055;
    10: op1_06_in25 = reg_0518;
    11: op1_06_in25 = imem03_in[115:112];
    12: op1_06_in25 = reg_0197;
    35: op1_06_in25 = reg_0197;
    13: op1_06_in25 = reg_0153;
    15: op1_06_in25 = imem01_in[59:56];
    16: op1_06_in25 = reg_0054;
    17: op1_06_in25 = reg_0142;
    18: op1_06_in25 = reg_0281;
    19: op1_06_in25 = reg_0808;
    20: op1_06_in25 = reg_0578;
    21: op1_06_in25 = imem07_in[11:8];
    50: op1_06_in25 = imem07_in[11:8];
    22: op1_06_in25 = reg_0593;
    24: op1_06_in25 = imem02_in[39:36];
    25: op1_06_in25 = reg_0888;
    26: op1_06_in25 = imem07_in[71:68];
    27: op1_06_in25 = reg_0067;
    28: op1_06_in25 = reg_0132;
    29: op1_06_in25 = imem03_in[123:120];
    30: op1_06_in25 = reg_0051;
    31: op1_06_in25 = reg_0616;
    32: op1_06_in25 = reg_0560;
    33: op1_06_in25 = reg_0636;
    34: op1_06_in25 = reg_0748;
    37: op1_06_in25 = imem01_in[115:112];
    86: op1_06_in25 = imem01_in[115:112];
    38: op1_06_in25 = imem01_in[63:60];
    39: op1_06_in25 = reg_0396;
    40: op1_06_in25 = imem05_in[35:32];
    41: op1_06_in25 = reg_0975;
    42: op1_06_in25 = reg_0443;
    43: op1_06_in25 = reg_0236;
    44: op1_06_in25 = reg_1050;
    45: op1_06_in25 = reg_0914;
    47: op1_06_in25 = imem03_in[59:56];
    48: op1_06_in25 = reg_1046;
    51: op1_06_in25 = reg_0446;
    52: op1_06_in25 = reg_0833;
    53: op1_06_in25 = reg_0882;
    54: op1_06_in25 = reg_0129;
    55: op1_06_in25 = reg_0704;
    56: op1_06_in25 = reg_0700;
    58: op1_06_in25 = reg_0786;
    60: op1_06_in25 = reg_0647;
    61: op1_06_in25 = reg_0870;
    62: op1_06_in25 = imem03_in[111:108];
    63: op1_06_in25 = reg_0571;
    64: op1_06_in25 = reg_0386;
    68: op1_06_in25 = imem02_in[95:92];
    69: op1_06_in25 = imem05_in[23:20];
    70: op1_06_in25 = reg_0161;
    71: op1_06_in25 = reg_1023;
    72: op1_06_in25 = reg_0426;
    75: op1_06_in25 = reg_1055;
    76: op1_06_in25 = reg_1001;
    77: op1_06_in25 = reg_1049;
    78: op1_06_in25 = reg_0292;
    89: op1_06_in25 = reg_0292;
    79: op1_06_in25 = reg_0789;
    81: op1_06_in25 = reg_0546;
    83: op1_06_in25 = reg_0154;
    84: op1_06_in25 = reg_0840;
    87: op1_06_in25 = imem05_in[11:8];
    88: op1_06_in25 = reg_0162;
    93: op1_06_in25 = reg_0631;
    94: op1_06_in25 = reg_0037;
    95: op1_06_in25 = reg_0650;
    96: op1_06_in25 = reg_0278;
    97: op1_06_in25 = reg_0089;
    default: op1_06_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv25 = 1;
    6: op1_06_inv25 = 1;
    7: op1_06_inv25 = 1;
    9: op1_06_inv25 = 1;
    15: op1_06_inv25 = 1;
    22: op1_06_inv25 = 1;
    23: op1_06_inv25 = 1;
    25: op1_06_inv25 = 1;
    29: op1_06_inv25 = 1;
    30: op1_06_inv25 = 1;
    31: op1_06_inv25 = 1;
    32: op1_06_inv25 = 1;
    33: op1_06_inv25 = 1;
    39: op1_06_inv25 = 1;
    40: op1_06_inv25 = 1;
    42: op1_06_inv25 = 1;
    43: op1_06_inv25 = 1;
    45: op1_06_inv25 = 1;
    48: op1_06_inv25 = 1;
    50: op1_06_inv25 = 1;
    52: op1_06_inv25 = 1;
    53: op1_06_inv25 = 1;
    54: op1_06_inv25 = 1;
    56: op1_06_inv25 = 1;
    62: op1_06_inv25 = 1;
    70: op1_06_inv25 = 1;
    71: op1_06_inv25 = 1;
    75: op1_06_inv25 = 1;
    76: op1_06_inv25 = 1;
    77: op1_06_inv25 = 1;
    79: op1_06_inv25 = 1;
    83: op1_06_inv25 = 1;
    89: op1_06_inv25 = 1;
    95: op1_06_inv25 = 1;
    default: op1_06_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in26 = reg_0563;
    6: op1_06_in26 = reg_0216;
    7: op1_06_in26 = reg_0954;
    9: op1_06_in26 = imem03_in[7:4];
    10: op1_06_in26 = reg_0515;
    11: op1_06_in26 = reg_0582;
    12: op1_06_in26 = imem01_in[11:8];
    13: op1_06_in26 = reg_0131;
    15: op1_06_in26 = reg_1053;
    16: op1_06_in26 = reg_0058;
    17: op1_06_in26 = reg_0138;
    18: op1_06_in26 = reg_0260;
    19: op1_06_in26 = reg_0801;
    20: op1_06_in26 = reg_0360;
    21: op1_06_in26 = imem07_in[15:12];
    22: op1_06_in26 = reg_0394;
    23: op1_06_in26 = imem03_in[99:96];
    24: op1_06_in26 = imem02_in[43:40];
    25: op1_06_in26 = reg_0537;
    26: op1_06_in26 = imem07_in[99:96];
    27: op1_06_in26 = reg_0014;
    28: op1_06_in26 = reg_0149;
    29: op1_06_in26 = reg_0585;
    30: op1_06_in26 = imem04_in[35:32];
    31: op1_06_in26 = reg_0606;
    32: op1_06_in26 = reg_0218;
    33: op1_06_in26 = reg_0652;
    34: op1_06_in26 = reg_0854;
    35: op1_06_in26 = imem01_in[55:52];
    37: op1_06_in26 = reg_0235;
    38: op1_06_in26 = imem01_in[67:64];
    39: op1_06_in26 = reg_0824;
    40: op1_06_in26 = imem05_in[75:72];
    41: op1_06_in26 = reg_0997;
    42: op1_06_in26 = reg_0448;
    43: op1_06_in26 = reg_0544;
    44: op1_06_in26 = reg_0327;
    45: op1_06_in26 = reg_0042;
    47: op1_06_in26 = imem03_in[67:64];
    48: op1_06_in26 = reg_0132;
    50: op1_06_in26 = imem07_in[23:20];
    51: op1_06_in26 = reg_0336;
    52: op1_06_in26 = reg_0373;
    53: op1_06_in26 = reg_0764;
    54: op1_06_in26 = reg_0144;
    55: op1_06_in26 = reg_0719;
    56: op1_06_in26 = reg_0805;
    58: op1_06_in26 = reg_0779;
    60: op1_06_in26 = reg_0643;
    61: op1_06_in26 = reg_0236;
    62: op1_06_in26 = imem03_in[119:116];
    63: op1_06_in26 = imem07_in[67:64];
    64: op1_06_in26 = reg_0371;
    68: op1_06_in26 = reg_0914;
    69: op1_06_in26 = imem05_in[51:48];
    70: op1_06_in26 = reg_0182;
    71: op1_06_in26 = reg_0592;
    72: op1_06_in26 = reg_0419;
    75: op1_06_in26 = reg_0733;
    76: op1_06_in26 = reg_0978;
    77: op1_06_in26 = reg_0051;
    78: op1_06_in26 = reg_0050;
    79: op1_06_in26 = imem07_in[3:0];
    81: op1_06_in26 = reg_0904;
    83: op1_06_in26 = reg_0957;
    84: op1_06_in26 = reg_0484;
    86: op1_06_in26 = reg_0968;
    87: op1_06_in26 = imem05_in[15:12];
    88: op1_06_in26 = reg_0374;
    89: op1_06_in26 = reg_0799;
    93: op1_06_in26 = reg_0662;
    94: op1_06_in26 = reg_0045;
    95: op1_06_in26 = reg_0730;
    96: op1_06_in26 = reg_0672;
    97: op1_06_in26 = reg_0409;
    default: op1_06_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv26 = 1;
    6: op1_06_inv26 = 1;
    9: op1_06_inv26 = 1;
    11: op1_06_inv26 = 1;
    12: op1_06_inv26 = 1;
    18: op1_06_inv26 = 1;
    19: op1_06_inv26 = 1;
    22: op1_06_inv26 = 1;
    24: op1_06_inv26 = 1;
    25: op1_06_inv26 = 1;
    27: op1_06_inv26 = 1;
    28: op1_06_inv26 = 1;
    34: op1_06_inv26 = 1;
    39: op1_06_inv26 = 1;
    44: op1_06_inv26 = 1;
    56: op1_06_inv26 = 1;
    63: op1_06_inv26 = 1;
    68: op1_06_inv26 = 1;
    69: op1_06_inv26 = 1;
    71: op1_06_inv26 = 1;
    75: op1_06_inv26 = 1;
    77: op1_06_inv26 = 1;
    83: op1_06_inv26 = 1;
    84: op1_06_inv26 = 1;
    86: op1_06_inv26 = 1;
    88: op1_06_inv26 = 1;
    89: op1_06_inv26 = 1;
    94: op1_06_inv26 = 1;
    96: op1_06_inv26 = 1;
    97: op1_06_inv26 = 1;
    default: op1_06_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in27 = reg_0322;
    6: op1_06_in27 = reg_0123;
    7: op1_06_in27 = reg_0969;
    9: op1_06_in27 = imem03_in[11:8];
    10: op1_06_in27 = reg_0516;
    11: op1_06_in27 = reg_0573;
    12: op1_06_in27 = imem01_in[27:24];
    13: op1_06_in27 = imem06_in[47:44];
    15: op1_06_in27 = reg_0735;
    16: op1_06_in27 = reg_0076;
    17: op1_06_in27 = reg_0153;
    18: op1_06_in27 = reg_0776;
    19: op1_06_in27 = reg_1010;
    20: op1_06_in27 = reg_0311;
    21: op1_06_in27 = imem07_in[19:16];
    22: op1_06_in27 = reg_0395;
    23: op1_06_in27 = imem03_in[127:124];
    62: op1_06_in27 = imem03_in[127:124];
    24: op1_06_in27 = imem02_in[67:64];
    25: op1_06_in27 = reg_0061;
    26: op1_06_in27 = imem07_in[107:104];
    27: op1_06_in27 = reg_0075;
    28: op1_06_in27 = reg_0145;
    29: op1_06_in27 = reg_0578;
    30: op1_06_in27 = imem04_in[63:60];
    31: op1_06_in27 = reg_0627;
    32: op1_06_in27 = reg_1032;
    33: op1_06_in27 = reg_0663;
    34: op1_06_in27 = reg_0875;
    35: op1_06_in27 = imem01_in[59:56];
    37: op1_06_in27 = reg_0560;
    38: op1_06_in27 = imem01_in[87:84];
    39: op1_06_in27 = reg_0823;
    40: op1_06_in27 = imem05_in[83:80];
    41: op1_06_in27 = imem04_in[3:0];
    42: op1_06_in27 = reg_0160;
    43: op1_06_in27 = reg_0830;
    44: op1_06_in27 = reg_0389;
    45: op1_06_in27 = reg_0294;
    47: op1_06_in27 = imem03_in[83:80];
    48: op1_06_in27 = reg_0133;
    50: op1_06_in27 = imem07_in[35:32];
    51: op1_06_in27 = reg_0404;
    52: op1_06_in27 = reg_0982;
    53: op1_06_in27 = imem05_in[27:24];
    87: op1_06_in27 = imem05_in[27:24];
    54: op1_06_in27 = reg_0613;
    55: op1_06_in27 = reg_0721;
    56: op1_06_in27 = reg_0361;
    58: op1_06_in27 = reg_0223;
    60: op1_06_in27 = reg_0648;
    61: op1_06_in27 = reg_1039;
    63: op1_06_in27 = imem07_in[127:124];
    64: op1_06_in27 = reg_0955;
    68: op1_06_in27 = reg_0647;
    69: op1_06_in27 = imem05_in[71:68];
    71: op1_06_in27 = reg_0831;
    72: op1_06_in27 = reg_0350;
    75: op1_06_in27 = reg_0114;
    76: op1_06_in27 = reg_0981;
    77: op1_06_in27 = reg_0998;
    78: op1_06_in27 = reg_0541;
    79: op1_06_in27 = imem07_in[11:8];
    81: op1_06_in27 = reg_0522;
    83: op1_06_in27 = reg_0707;
    84: op1_06_in27 = reg_0884;
    86: op1_06_in27 = reg_0546;
    88: op1_06_in27 = reg_0515;
    89: op1_06_in27 = reg_0848;
    93: op1_06_in27 = reg_0623;
    94: op1_06_in27 = reg_0341;
    95: op1_06_in27 = imem03_in[3:0];
    96: op1_06_in27 = reg_0373;
    97: op1_06_in27 = reg_0232;
    default: op1_06_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv27 = 1;
    6: op1_06_inv27 = 1;
    10: op1_06_inv27 = 1;
    11: op1_06_inv27 = 1;
    12: op1_06_inv27 = 1;
    13: op1_06_inv27 = 1;
    18: op1_06_inv27 = 1;
    19: op1_06_inv27 = 1;
    20: op1_06_inv27 = 1;
    23: op1_06_inv27 = 1;
    25: op1_06_inv27 = 1;
    26: op1_06_inv27 = 1;
    27: op1_06_inv27 = 1;
    29: op1_06_inv27 = 1;
    30: op1_06_inv27 = 1;
    31: op1_06_inv27 = 1;
    32: op1_06_inv27 = 1;
    34: op1_06_inv27 = 1;
    37: op1_06_inv27 = 1;
    47: op1_06_inv27 = 1;
    51: op1_06_inv27 = 1;
    53: op1_06_inv27 = 1;
    54: op1_06_inv27 = 1;
    55: op1_06_inv27 = 1;
    60: op1_06_inv27 = 1;
    63: op1_06_inv27 = 1;
    69: op1_06_inv27 = 1;
    71: op1_06_inv27 = 1;
    75: op1_06_inv27 = 1;
    76: op1_06_inv27 = 1;
    77: op1_06_inv27 = 1;
    83: op1_06_inv27 = 1;
    87: op1_06_inv27 = 1;
    89: op1_06_inv27 = 1;
    95: op1_06_inv27 = 1;
    96: op1_06_inv27 = 1;
    97: op1_06_inv27 = 1;
    default: op1_06_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in28 = reg_0323;
    6: op1_06_in28 = reg_0105;
    7: op1_06_in28 = reg_0950;
    9: op1_06_in28 = imem03_in[43:40];
    10: op1_06_in28 = imem01_in[19:16];
    11: op1_06_in28 = reg_0578;
    12: op1_06_in28 = imem01_in[35:32];
    13: op1_06_in28 = imem06_in[71:68];
    15: op1_06_in28 = reg_0503;
    16: op1_06_in28 = imem05_in[3:0];
    34: op1_06_in28 = imem05_in[3:0];
    17: op1_06_in28 = imem06_in[43:40];
    18: op1_06_in28 = reg_0857;
    19: op1_06_in28 = reg_0011;
    20: op1_06_in28 = reg_0374;
    21: op1_06_in28 = imem07_in[51:48];
    22: op1_06_in28 = reg_0369;
    23: op1_06_in28 = reg_0592;
    24: op1_06_in28 = imem02_in[75:72];
    25: op1_06_in28 = reg_0763;
    26: op1_06_in28 = imem07_in[115:112];
    27: op1_06_in28 = reg_0064;
    28: op1_06_in28 = reg_0136;
    29: op1_06_in28 = reg_0795;
    30: op1_06_in28 = imem04_in[123:120];
    31: op1_06_in28 = reg_0615;
    32: op1_06_in28 = reg_0830;
    33: op1_06_in28 = reg_0095;
    35: op1_06_in28 = imem01_in[71:68];
    37: op1_06_in28 = reg_0239;
    38: op1_06_in28 = imem01_in[111:108];
    39: op1_06_in28 = reg_0923;
    44: op1_06_in28 = reg_0923;
    40: op1_06_in28 = imem05_in[87:84];
    41: op1_06_in28 = imem04_in[107:104];
    42: op1_06_in28 = reg_0183;
    43: op1_06_in28 = reg_0123;
    45: op1_06_in28 = reg_0349;
    47: op1_06_in28 = imem03_in[99:96];
    48: op1_06_in28 = reg_0144;
    50: op1_06_in28 = imem07_in[39:36];
    51: op1_06_in28 = reg_0819;
    52: op1_06_in28 = reg_0991;
    53: op1_06_in28 = imem05_in[31:28];
    54: op1_06_in28 = reg_0073;
    55: op1_06_in28 = reg_0726;
    56: op1_06_in28 = reg_0303;
    58: op1_06_in28 = reg_0936;
    60: op1_06_in28 = reg_0652;
    61: op1_06_in28 = reg_0496;
    62: op1_06_in28 = reg_0006;
    63: op1_06_in28 = reg_0728;
    64: op1_06_in28 = reg_0957;
    68: op1_06_in28 = reg_0224;
    69: op1_06_in28 = imem05_in[95:92];
    71: op1_06_in28 = reg_0904;
    72: op1_06_in28 = reg_0174;
    75: op1_06_in28 = reg_0115;
    76: op1_06_in28 = reg_0975;
    77: op1_06_in28 = reg_0984;
    78: op1_06_in28 = reg_0537;
    79: op1_06_in28 = imem07_in[47:44];
    81: op1_06_in28 = reg_0733;
    83: op1_06_in28 = reg_0780;
    84: op1_06_in28 = imem03_in[39:36];
    86: op1_06_in28 = reg_0234;
    87: op1_06_in28 = imem05_in[71:68];
    88: op1_06_in28 = reg_0299;
    89: op1_06_in28 = reg_0752;
    93: op1_06_in28 = reg_0238;
    94: op1_06_in28 = imem03_in[11:8];
    95: op1_06_in28 = imem03_in[55:52];
    96: op1_06_in28 = reg_0986;
    97: op1_06_in28 = reg_0832;
    default: op1_06_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_06_inv28 = 1;
    11: op1_06_inv28 = 1;
    19: op1_06_inv28 = 1;
    22: op1_06_inv28 = 1;
    23: op1_06_inv28 = 1;
    24: op1_06_inv28 = 1;
    26: op1_06_inv28 = 1;
    27: op1_06_inv28 = 1;
    28: op1_06_inv28 = 1;
    30: op1_06_inv28 = 1;
    31: op1_06_inv28 = 1;
    33: op1_06_inv28 = 1;
    38: op1_06_inv28 = 1;
    40: op1_06_inv28 = 1;
    41: op1_06_inv28 = 1;
    42: op1_06_inv28 = 1;
    43: op1_06_inv28 = 1;
    47: op1_06_inv28 = 1;
    48: op1_06_inv28 = 1;
    50: op1_06_inv28 = 1;
    51: op1_06_inv28 = 1;
    52: op1_06_inv28 = 1;
    55: op1_06_inv28 = 1;
    56: op1_06_inv28 = 1;
    58: op1_06_inv28 = 1;
    61: op1_06_inv28 = 1;
    68: op1_06_inv28 = 1;
    69: op1_06_inv28 = 1;
    76: op1_06_inv28 = 1;
    83: op1_06_inv28 = 1;
    86: op1_06_inv28 = 1;
    88: op1_06_inv28 = 1;
    89: op1_06_inv28 = 1;
    94: op1_06_inv28 = 1;
    default: op1_06_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in29 = reg_0006;
    6: op1_06_in29 = reg_0124;
    43: op1_06_in29 = reg_0124;
    7: op1_06_in29 = reg_0965;
    9: op1_06_in29 = imem03_in[55:52];
    10: op1_06_in29 = imem01_in[75:72];
    11: op1_06_in29 = reg_0581;
    12: op1_06_in29 = imem01_in[127:124];
    13: op1_06_in29 = imem06_in[115:112];
    15: op1_06_in29 = reg_0507;
    16: op1_06_in29 = imem05_in[7:4];
    17: op1_06_in29 = imem06_in[67:64];
    18: op1_06_in29 = reg_0485;
    19: op1_06_in29 = imem07_in[3:0];
    20: op1_06_in29 = reg_0389;
    21: op1_06_in29 = imem07_in[63:60];
    79: op1_06_in29 = imem07_in[63:60];
    22: op1_06_in29 = reg_0985;
    23: op1_06_in29 = reg_0591;
    24: op1_06_in29 = imem02_in[79:76];
    25: op1_06_in29 = reg_0078;
    26: op1_06_in29 = reg_0716;
    63: op1_06_in29 = reg_0716;
    27: op1_06_in29 = reg_0047;
    28: op1_06_in29 = reg_0133;
    29: op1_06_in29 = reg_0373;
    30: op1_06_in29 = reg_0483;
    31: op1_06_in29 = reg_0348;
    32: op1_06_in29 = reg_1040;
    33: op1_06_in29 = reg_0098;
    34: op1_06_in29 = imem05_in[23:20];
    35: op1_06_in29 = imem01_in[87:84];
    37: op1_06_in29 = reg_0274;
    38: op1_06_in29 = imem01_in[115:112];
    39: op1_06_in29 = reg_0369;
    40: op1_06_in29 = reg_0954;
    41: op1_06_in29 = imem04_in[111:108];
    42: op1_06_in29 = reg_0164;
    44: op1_06_in29 = reg_0784;
    45: op1_06_in29 = reg_0629;
    47: op1_06_in29 = reg_0357;
    48: op1_06_in29 = imem06_in[43:40];
    50: op1_06_in29 = imem07_in[83:80];
    51: op1_06_in29 = reg_0489;
    52: op1_06_in29 = reg_0992;
    53: op1_06_in29 = imem05_in[39:36];
    54: op1_06_in29 = reg_0895;
    55: op1_06_in29 = reg_0717;
    56: op1_06_in29 = reg_0744;
    58: op1_06_in29 = reg_0218;
    60: op1_06_in29 = reg_0081;
    61: op1_06_in29 = reg_0604;
    62: op1_06_in29 = reg_0535;
    64: op1_06_in29 = imem07_in[7:4];
    68: op1_06_in29 = reg_0894;
    69: op1_06_in29 = imem05_in[99:96];
    71: op1_06_in29 = reg_0225;
    72: op1_06_in29 = reg_0181;
    75: op1_06_in29 = reg_0110;
    76: op1_06_in29 = imem04_in[7:4];
    77: op1_06_in29 = reg_0993;
    78: op1_06_in29 = reg_0014;
    81: op1_06_in29 = reg_0114;
    97: op1_06_in29 = reg_0114;
    83: op1_06_in29 = reg_0508;
    84: op1_06_in29 = imem03_in[43:40];
    86: op1_06_in29 = reg_1024;
    87: op1_06_in29 = imem05_in[87:84];
    88: op1_06_in29 = reg_0727;
    89: op1_06_in29 = reg_0732;
    93: op1_06_in29 = reg_0278;
    94: op1_06_in29 = imem03_in[123:120];
    95: op1_06_in29 = imem03_in[79:76];
    96: op1_06_in29 = reg_0978;
    default: op1_06_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv29 = 1;
    6: op1_06_inv29 = 1;
    7: op1_06_inv29 = 1;
    10: op1_06_inv29 = 1;
    11: op1_06_inv29 = 1;
    12: op1_06_inv29 = 1;
    13: op1_06_inv29 = 1;
    15: op1_06_inv29 = 1;
    17: op1_06_inv29 = 1;
    19: op1_06_inv29 = 1;
    21: op1_06_inv29 = 1;
    22: op1_06_inv29 = 1;
    23: op1_06_inv29 = 1;
    24: op1_06_inv29 = 1;
    29: op1_06_inv29 = 1;
    30: op1_06_inv29 = 1;
    31: op1_06_inv29 = 1;
    34: op1_06_inv29 = 1;
    38: op1_06_inv29 = 1;
    40: op1_06_inv29 = 1;
    42: op1_06_inv29 = 1;
    45: op1_06_inv29 = 1;
    47: op1_06_inv29 = 1;
    48: op1_06_inv29 = 1;
    52: op1_06_inv29 = 1;
    53: op1_06_inv29 = 1;
    54: op1_06_inv29 = 1;
    56: op1_06_inv29 = 1;
    58: op1_06_inv29 = 1;
    60: op1_06_inv29 = 1;
    61: op1_06_inv29 = 1;
    62: op1_06_inv29 = 1;
    64: op1_06_inv29 = 1;
    69: op1_06_inv29 = 1;
    71: op1_06_inv29 = 1;
    72: op1_06_inv29 = 1;
    76: op1_06_inv29 = 1;
    77: op1_06_inv29 = 1;
    78: op1_06_inv29 = 1;
    79: op1_06_inv29 = 1;
    81: op1_06_inv29 = 1;
    86: op1_06_inv29 = 1;
    87: op1_06_inv29 = 1;
    88: op1_06_inv29 = 1;
    89: op1_06_inv29 = 1;
    93: op1_06_inv29 = 1;
    95: op1_06_inv29 = 1;
    97: op1_06_inv29 = 1;
    default: op1_06_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_06_in30 = reg_0001;
    6: op1_06_in30 = reg_0125;
    7: op1_06_in30 = reg_0961;
    9: op1_06_in30 = imem03_in[59:56];
    10: op1_06_in30 = imem01_in[79:76];
    11: op1_06_in30 = reg_0398;
    12: op1_06_in30 = reg_0240;
    38: op1_06_in30 = reg_0240;
    13: op1_06_in30 = reg_0621;
    15: op1_06_in30 = reg_0249;
    16: op1_06_in30 = imem05_in[27:24];
    17: op1_06_in30 = imem06_in[95:92];
    48: op1_06_in30 = imem06_in[95:92];
    18: op1_06_in30 = reg_0552;
    19: op1_06_in30 = imem07_in[27:24];
    20: op1_06_in30 = reg_0995;
    21: op1_06_in30 = imem07_in[75:72];
    22: op1_06_in30 = reg_0991;
    23: op1_06_in30 = reg_0593;
    24: op1_06_in30 = reg_0656;
    25: op1_06_in30 = reg_0067;
    26: op1_06_in30 = reg_0704;
    27: op1_06_in30 = reg_0864;
    28: op1_06_in30 = reg_0131;
    29: op1_06_in30 = reg_0369;
    30: op1_06_in30 = reg_0511;
    31: op1_06_in30 = reg_0344;
    32: op1_06_in30 = reg_1035;
    33: op1_06_in30 = reg_0857;
    34: op1_06_in30 = imem05_in[95:92];
    35: op1_06_in30 = reg_0013;
    37: op1_06_in30 = reg_1039;
    71: op1_06_in30 = reg_1039;
    39: op1_06_in30 = reg_0820;
    40: op1_06_in30 = reg_0956;
    41: op1_06_in30 = imem04_in[115:112];
    43: op1_06_in30 = reg_0119;
    44: op1_06_in30 = reg_0509;
    45: op1_06_in30 = reg_0241;
    47: op1_06_in30 = reg_1007;
    50: op1_06_in30 = reg_0722;
    51: op1_06_in30 = reg_0137;
    52: op1_06_in30 = reg_0979;
    53: op1_06_in30 = imem05_in[75:72];
    54: op1_06_in30 = reg_0624;
    55: op1_06_in30 = reg_0702;
    56: op1_06_in30 = reg_0641;
    58: op1_06_in30 = reg_0919;
    60: op1_06_in30 = reg_0424;
    61: op1_06_in30 = reg_0520;
    62: op1_06_in30 = reg_0099;
    63: op1_06_in30 = reg_0710;
    64: op1_06_in30 = imem07_in[67:64];
    68: op1_06_in30 = reg_0648;
    69: op1_06_in30 = reg_0650;
    72: op1_06_in30 = reg_0160;
    75: op1_06_in30 = imem02_in[7:4];
    76: op1_06_in30 = imem04_in[11:8];
    77: op1_06_in30 = reg_0980;
    78: op1_06_in30 = reg_0068;
    79: op1_06_in30 = imem07_in[95:92];
    81: op1_06_in30 = imem02_in[23:20];
    83: op1_06_in30 = imem06_in[19:16];
    84: op1_06_in30 = imem03_in[99:96];
    86: op1_06_in30 = reg_0962;
    87: op1_06_in30 = imem05_in[115:112];
    88: op1_06_in30 = reg_0422;
    89: op1_06_in30 = reg_0108;
    93: op1_06_in30 = reg_0281;
    94: op1_06_in30 = reg_0784;
    95: op1_06_in30 = reg_0758;
    96: op1_06_in30 = reg_0989;
    97: op1_06_in30 = imem02_in[27:24];
    default: op1_06_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv30 = 1;
    6: op1_06_inv30 = 1;
    9: op1_06_inv30 = 1;
    11: op1_06_inv30 = 1;
    12: op1_06_inv30 = 1;
    13: op1_06_inv30 = 1;
    15: op1_06_inv30 = 1;
    17: op1_06_inv30 = 1;
    18: op1_06_inv30 = 1;
    20: op1_06_inv30 = 1;
    21: op1_06_inv30 = 1;
    24: op1_06_inv30 = 1;
    27: op1_06_inv30 = 1;
    30: op1_06_inv30 = 1;
    32: op1_06_inv30 = 1;
    33: op1_06_inv30 = 1;
    39: op1_06_inv30 = 1;
    40: op1_06_inv30 = 1;
    44: op1_06_inv30 = 1;
    45: op1_06_inv30 = 1;
    47: op1_06_inv30 = 1;
    50: op1_06_inv30 = 1;
    51: op1_06_inv30 = 1;
    52: op1_06_inv30 = 1;
    53: op1_06_inv30 = 1;
    55: op1_06_inv30 = 1;
    56: op1_06_inv30 = 1;
    58: op1_06_inv30 = 1;
    63: op1_06_inv30 = 1;
    68: op1_06_inv30 = 1;
    69: op1_06_inv30 = 1;
    76: op1_06_inv30 = 1;
    86: op1_06_inv30 = 1;
    89: op1_06_inv30 = 1;
    94: op1_06_inv30 = 1;
    95: op1_06_inv30 = 1;
    96: op1_06_inv30 = 1;
    default: op1_06_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_06_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_06_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in00 = reg_0007;
    6: op1_07_in00 = reg_0102;
    7: op1_07_in00 = reg_0947;
    8: op1_07_in00 = imem00_in[23:20];
    67: op1_07_in00 = imem00_in[23:20];
    85: op1_07_in00 = imem00_in[23:20];
    9: op1_07_in00 = imem03_in[83:80];
    10: op1_07_in00 = imem01_in[91:88];
    11: op1_07_in00 = reg_0397;
    12: op1_07_in00 = reg_0502;
    56: op1_07_in00 = reg_0502;
    13: op1_07_in00 = reg_0606;
    14: op1_07_in00 = imem00_in[11:8];
    46: op1_07_in00 = imem00_in[11:8];
    57: op1_07_in00 = imem00_in[11:8];
    4: op1_07_in00 = imem07_in[91:88];
    15: op1_07_in00 = reg_1040;
    16: op1_07_in00 = imem05_in[31:28];
    17: op1_07_in00 = imem06_in[123:120];
    18: op1_07_in00 = reg_0534;
    19: op1_07_in00 = imem07_in[35:32];
    20: op1_07_in00 = imem04_in[3:0];
    21: op1_07_in00 = imem07_in[87:84];
    3: op1_07_in00 = imem07_in[55:52];
    2: op1_07_in00 = imem07_in[55:52];
    22: op1_07_in00 = reg_0979;
    23: op1_07_in00 = reg_0580;
    24: op1_07_in00 = reg_0651;
    25: op1_07_in00 = reg_0014;
    26: op1_07_in00 = imem00_in[43:40];
    36: op1_07_in00 = imem00_in[43:40];
    27: op1_07_in00 = imem05_in[11:8];
    28: op1_07_in00 = imem06_in[43:40];
    83: op1_07_in00 = imem06_in[43:40];
    29: op1_07_in00 = reg_0051;
    30: op1_07_in00 = reg_0541;
    31: op1_07_in00 = reg_0914;
    32: op1_07_in00 = reg_1015;
    33: op1_07_in00 = reg_0817;
    34: op1_07_in00 = imem05_in[115:112];
    35: op1_07_in00 = reg_0786;
    37: op1_07_in00 = reg_0869;
    38: op1_07_in00 = reg_0860;
    39: op1_07_in00 = reg_0518;
    40: op1_07_in00 = reg_0950;
    41: op1_07_in00 = imem04_in[123:120];
    42: op1_07_in00 = imem00_in[99:96];
    92: op1_07_in00 = imem00_in[99:96];
    43: op1_07_in00 = reg_0100;
    44: op1_07_in00 = reg_0820;
    45: op1_07_in00 = reg_0029;
    47: op1_07_in00 = reg_1019;
    48: op1_07_in00 = imem06_in[99:96];
    49: op1_07_in00 = imem00_in[7:4];
    70: op1_07_in00 = imem00_in[7:4];
    50: op1_07_in00 = reg_0717;
    51: op1_07_in00 = imem06_in[3:0];
    52: op1_07_in00 = reg_1000;
    53: op1_07_in00 = reg_0969;
    54: op1_07_in00 = reg_0486;
    55: op1_07_in00 = reg_0703;
    58: op1_07_in00 = reg_1056;
    59: op1_07_in00 = imem00_in[31:28];
    73: op1_07_in00 = imem00_in[31:28];
    74: op1_07_in00 = imem00_in[31:28];
    60: op1_07_in00 = reg_0664;
    61: op1_07_in00 = reg_0514;
    62: op1_07_in00 = reg_0662;
    63: op1_07_in00 = reg_0726;
    64: op1_07_in00 = imem07_in[83:80];
    65: op1_07_in00 = imem00_in[27:24];
    66: op1_07_in00 = imem00_in[39:36];
    68: op1_07_in00 = reg_0908;
    69: op1_07_in00 = reg_0944;
    71: op1_07_in00 = reg_0798;
    72: op1_07_in00 = reg_0163;
    75: op1_07_in00 = imem02_in[15:12];
    76: op1_07_in00 = imem04_in[51:48];
    77: op1_07_in00 = reg_0978;
    78: op1_07_in00 = reg_0658;
    79: op1_07_in00 = imem07_in[103:100];
    80: op1_07_in00 = imem00_in[59:56];
    81: op1_07_in00 = imem02_in[31:28];
    82: op1_07_in00 = imem00_in[3:0];
    84: op1_07_in00 = imem03_in[107:104];
    86: op1_07_in00 = reg_0520;
    87: op1_07_in00 = reg_0508;
    88: op1_07_in00 = reg_0532;
    89: op1_07_in00 = reg_0824;
    90: op1_07_in00 = imem00_in[15:12];
    91: op1_07_in00 = reg_0513;
    93: op1_07_in00 = reg_0230;
    94: op1_07_in00 = reg_0836;
    95: op1_07_in00 = reg_0049;
    96: op1_07_in00 = reg_0981;
    97: op1_07_in00 = imem02_in[123:120];
    default: op1_07_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_07_inv00 = 1;
    9: op1_07_inv00 = 1;
    11: op1_07_inv00 = 1;
    12: op1_07_inv00 = 1;
    4: op1_07_inv00 = 1;
    16: op1_07_inv00 = 1;
    17: op1_07_inv00 = 1;
    19: op1_07_inv00 = 1;
    20: op1_07_inv00 = 1;
    21: op1_07_inv00 = 1;
    22: op1_07_inv00 = 1;
    24: op1_07_inv00 = 1;
    26: op1_07_inv00 = 1;
    31: op1_07_inv00 = 1;
    32: op1_07_inv00 = 1;
    34: op1_07_inv00 = 1;
    35: op1_07_inv00 = 1;
    37: op1_07_inv00 = 1;
    38: op1_07_inv00 = 1;
    40: op1_07_inv00 = 1;
    45: op1_07_inv00 = 1;
    48: op1_07_inv00 = 1;
    49: op1_07_inv00 = 1;
    50: op1_07_inv00 = 1;
    51: op1_07_inv00 = 1;
    53: op1_07_inv00 = 1;
    58: op1_07_inv00 = 1;
    62: op1_07_inv00 = 1;
    66: op1_07_inv00 = 1;
    71: op1_07_inv00 = 1;
    74: op1_07_inv00 = 1;
    75: op1_07_inv00 = 1;
    77: op1_07_inv00 = 1;
    78: op1_07_inv00 = 1;
    79: op1_07_inv00 = 1;
    80: op1_07_inv00 = 1;
    83: op1_07_inv00 = 1;
    91: op1_07_inv00 = 1;
    92: op1_07_inv00 = 1;
    93: op1_07_inv00 = 1;
    94: op1_07_inv00 = 1;
    96: op1_07_inv00 = 1;
    97: op1_07_inv00 = 1;
    default: op1_07_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in01 = reg_0008;
    6: op1_07_in01 = reg_0115;
    7: op1_07_in01 = reg_0259;
    8: op1_07_in01 = imem00_in[27:24];
    67: op1_07_in01 = imem00_in[27:24];
    9: op1_07_in01 = imem03_in[87:84];
    10: op1_07_in01 = imem01_in[111:108];
    11: op1_07_in01 = reg_0361;
    12: op1_07_in01 = reg_0248;
    13: op1_07_in01 = reg_0609;
    14: op1_07_in01 = imem00_in[15:12];
    49: op1_07_in01 = imem00_in[15:12];
    4: op1_07_in01 = reg_0443;
    15: op1_07_in01 = reg_0913;
    16: op1_07_in01 = imem05_in[63:60];
    17: op1_07_in01 = reg_0610;
    18: op1_07_in01 = reg_0535;
    19: op1_07_in01 = imem07_in[63:60];
    2: op1_07_in01 = imem07_in[63:60];
    20: op1_07_in01 = imem04_in[47:44];
    21: op1_07_in01 = imem07_in[99:96];
    3: op1_07_in01 = imem07_in[103:100];
    22: op1_07_in01 = reg_0975;
    23: op1_07_in01 = reg_0384;
    24: op1_07_in01 = reg_0652;
    25: op1_07_in01 = reg_0068;
    26: op1_07_in01 = imem00_in[95:92];
    57: op1_07_in01 = imem00_in[95:92];
    27: op1_07_in01 = imem05_in[23:20];
    28: op1_07_in01 = imem06_in[71:68];
    29: op1_07_in01 = reg_0987;
    39: op1_07_in01 = reg_0987;
    30: op1_07_in01 = reg_0763;
    31: op1_07_in01 = reg_0399;
    32: op1_07_in01 = reg_0228;
    33: op1_07_in01 = reg_0090;
    34: op1_07_in01 = imem05_in[123:120];
    35: op1_07_in01 = reg_0779;
    36: op1_07_in01 = imem00_in[63:60];
    37: op1_07_in01 = reg_0227;
    38: op1_07_in01 = reg_0247;
    40: op1_07_in01 = reg_0964;
    41: op1_07_in01 = reg_0301;
    42: op1_07_in01 = imem00_in[119:116];
    43: op1_07_in01 = reg_0107;
    44: op1_07_in01 = reg_1002;
    45: op1_07_in01 = imem07_in[11:8];
    46: op1_07_in01 = imem00_in[31:28];
    85: op1_07_in01 = imem00_in[31:28];
    47: op1_07_in01 = reg_0824;
    48: op1_07_in01 = imem06_in[119:116];
    50: op1_07_in01 = reg_0718;
    51: op1_07_in01 = imem06_in[15:12];
    52: op1_07_in01 = reg_0997;
    53: op1_07_in01 = reg_0951;
    54: op1_07_in01 = reg_0892;
    55: op1_07_in01 = reg_0724;
    56: op1_07_in01 = reg_0180;
    58: op1_07_in01 = reg_0592;
    59: op1_07_in01 = imem00_in[87:84];
    60: op1_07_in01 = reg_0389;
    61: op1_07_in01 = reg_0500;
    62: op1_07_in01 = reg_0823;
    63: op1_07_in01 = reg_0725;
    64: op1_07_in01 = imem07_in[123:120];
    65: op1_07_in01 = imem00_in[51:48];
    66: op1_07_in01 = imem00_in[43:40];
    73: op1_07_in01 = imem00_in[43:40];
    68: op1_07_in01 = reg_0233;
    69: op1_07_in01 = reg_0673;
    70: op1_07_in01 = imem00_in[107:104];
    71: op1_07_in01 = reg_0737;
    72: op1_07_in01 = reg_0166;
    74: op1_07_in01 = imem00_in[39:36];
    75: op1_07_in01 = imem02_in[19:16];
    76: op1_07_in01 = imem04_in[67:64];
    77: op1_07_in01 = reg_0999;
    78: op1_07_in01 = reg_0065;
    79: op1_07_in01 = imem07_in[107:104];
    80: op1_07_in01 = reg_0523;
    81: op1_07_in01 = imem02_in[63:60];
    82: op1_07_in01 = imem00_in[67:64];
    83: op1_07_in01 = imem06_in[51:48];
    84: op1_07_in01 = imem03_in[115:112];
    86: op1_07_in01 = reg_0514;
    87: op1_07_in01 = reg_0528;
    88: op1_07_in01 = reg_0599;
    89: op1_07_in01 = reg_0332;
    90: op1_07_in01 = imem00_in[75:72];
    91: op1_07_in01 = reg_0753;
    92: op1_07_in01 = imem00_in[123:120];
    93: op1_07_in01 = reg_0773;
    94: op1_07_in01 = reg_0307;
    95: op1_07_in01 = reg_0363;
    96: op1_07_in01 = imem04_in[15:12];
    97: op1_07_in01 = reg_0750;
    default: op1_07_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv01 = 1;
    6: op1_07_inv01 = 1;
    9: op1_07_inv01 = 1;
    12: op1_07_inv01 = 1;
    14: op1_07_inv01 = 1;
    4: op1_07_inv01 = 1;
    16: op1_07_inv01 = 1;
    18: op1_07_inv01 = 1;
    20: op1_07_inv01 = 1;
    23: op1_07_inv01 = 1;
    24: op1_07_inv01 = 1;
    2: op1_07_inv01 = 1;
    27: op1_07_inv01 = 1;
    34: op1_07_inv01 = 1;
    35: op1_07_inv01 = 1;
    36: op1_07_inv01 = 1;
    37: op1_07_inv01 = 1;
    39: op1_07_inv01 = 1;
    40: op1_07_inv01 = 1;
    41: op1_07_inv01 = 1;
    42: op1_07_inv01 = 1;
    44: op1_07_inv01 = 1;
    46: op1_07_inv01 = 1;
    48: op1_07_inv01 = 1;
    49: op1_07_inv01 = 1;
    50: op1_07_inv01 = 1;
    51: op1_07_inv01 = 1;
    52: op1_07_inv01 = 1;
    53: op1_07_inv01 = 1;
    55: op1_07_inv01 = 1;
    58: op1_07_inv01 = 1;
    61: op1_07_inv01 = 1;
    67: op1_07_inv01 = 1;
    68: op1_07_inv01 = 1;
    70: op1_07_inv01 = 1;
    73: op1_07_inv01 = 1;
    74: op1_07_inv01 = 1;
    75: op1_07_inv01 = 1;
    76: op1_07_inv01 = 1;
    77: op1_07_inv01 = 1;
    80: op1_07_inv01 = 1;
    81: op1_07_inv01 = 1;
    86: op1_07_inv01 = 1;
    87: op1_07_inv01 = 1;
    88: op1_07_inv01 = 1;
    92: op1_07_inv01 = 1;
    93: op1_07_inv01 = 1;
    94: op1_07_inv01 = 1;
    96: op1_07_inv01 = 1;
    default: op1_07_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in02 = reg_0009;
    6: op1_07_in02 = reg_0109;
    7: op1_07_in02 = reg_0241;
    8: op1_07_in02 = imem00_in[35:32];
    46: op1_07_in02 = imem00_in[35:32];
    67: op1_07_in02 = imem00_in[35:32];
    9: op1_07_in02 = imem03_in[107:104];
    10: op1_07_in02 = imem01_in[115:112];
    11: op1_07_in02 = reg_0992;
    44: op1_07_in02 = reg_0992;
    12: op1_07_in02 = reg_0237;
    13: op1_07_in02 = reg_0623;
    14: op1_07_in02 = imem00_in[55:52];
    4: op1_07_in02 = reg_0438;
    15: op1_07_in02 = reg_1036;
    16: op1_07_in02 = imem05_in[87:84];
    17: op1_07_in02 = reg_0604;
    18: op1_07_in02 = reg_0539;
    19: op1_07_in02 = imem07_in[75:72];
    20: op1_07_in02 = imem04_in[51:48];
    21: op1_07_in02 = imem07_in[119:116];
    79: op1_07_in02 = imem07_in[119:116];
    3: op1_07_in02 = imem07_in[111:108];
    22: op1_07_in02 = reg_0983;
    23: op1_07_in02 = reg_0391;
    24: op1_07_in02 = reg_0352;
    25: op1_07_in02 = reg_0071;
    2: op1_07_in02 = imem07_in[83:80];
    26: op1_07_in02 = imem00_in[127:124];
    42: op1_07_in02 = imem00_in[127:124];
    27: op1_07_in02 = imem05_in[47:44];
    28: op1_07_in02 = imem06_in[103:100];
    29: op1_07_in02 = reg_1002;
    30: op1_07_in02 = reg_0268;
    31: op1_07_in02 = reg_0804;
    32: op1_07_in02 = reg_0105;
    33: op1_07_in02 = reg_0506;
    34: op1_07_in02 = reg_0955;
    35: op1_07_in02 = reg_0560;
    36: op1_07_in02 = imem00_in[107:104];
    37: op1_07_in02 = reg_0119;
    38: op1_07_in02 = reg_0274;
    39: op1_07_in02 = reg_0982;
    40: op1_07_in02 = reg_0965;
    41: op1_07_in02 = reg_1003;
    43: op1_07_in02 = imem02_in[3:0];
    45: op1_07_in02 = imem07_in[55:52];
    47: op1_07_in02 = reg_0543;
    48: op1_07_in02 = reg_0356;
    49: op1_07_in02 = imem00_in[71:68];
    50: op1_07_in02 = reg_0707;
    51: op1_07_in02 = imem06_in[23:20];
    52: op1_07_in02 = imem04_in[11:8];
    53: op1_07_in02 = reg_0968;
    54: op1_07_in02 = reg_0371;
    55: op1_07_in02 = reg_0715;
    56: op1_07_in02 = reg_0178;
    57: op1_07_in02 = imem00_in[119:116];
    58: op1_07_in02 = reg_0503;
    59: op1_07_in02 = reg_0683;
    60: op1_07_in02 = reg_0425;
    61: op1_07_in02 = reg_1031;
    62: op1_07_in02 = reg_0370;
    63: op1_07_in02 = reg_0705;
    64: op1_07_in02 = reg_0728;
    65: op1_07_in02 = imem00_in[59:56];
    66: op1_07_in02 = imem00_in[83:80];
    85: op1_07_in02 = imem00_in[83:80];
    68: op1_07_in02 = reg_0423;
    69: op1_07_in02 = reg_0656;
    70: op1_07_in02 = imem00_in[111:108];
    71: op1_07_in02 = reg_0616;
    73: op1_07_in02 = imem00_in[91:88];
    74: op1_07_in02 = imem00_in[51:48];
    75: op1_07_in02 = imem02_in[23:20];
    76: op1_07_in02 = imem04_in[91:88];
    77: op1_07_in02 = reg_0981;
    78: op1_07_in02 = reg_0777;
    80: op1_07_in02 = reg_0738;
    81: op1_07_in02 = reg_0844;
    82: op1_07_in02 = imem00_in[103:100];
    83: op1_07_in02 = imem06_in[115:112];
    84: op1_07_in02 = reg_0620;
    86: op1_07_in02 = reg_1037;
    87: op1_07_in02 = reg_0816;
    88: op1_07_in02 = reg_0589;
    89: op1_07_in02 = imem05_in[19:16];
    90: op1_07_in02 = imem00_in[95:92];
    91: op1_07_in02 = imem00_in[11:8];
    92: op1_07_in02 = reg_0166;
    93: op1_07_in02 = reg_0767;
    94: op1_07_in02 = reg_0007;
    95: op1_07_in02 = reg_0346;
    96: op1_07_in02 = imem04_in[107:104];
    97: op1_07_in02 = reg_0536;
    default: op1_07_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_07_inv02 = 1;
    14: op1_07_inv02 = 1;
    16: op1_07_inv02 = 1;
    18: op1_07_inv02 = 1;
    19: op1_07_inv02 = 1;
    20: op1_07_inv02 = 1;
    21: op1_07_inv02 = 1;
    23: op1_07_inv02 = 1;
    24: op1_07_inv02 = 1;
    27: op1_07_inv02 = 1;
    28: op1_07_inv02 = 1;
    30: op1_07_inv02 = 1;
    34: op1_07_inv02 = 1;
    35: op1_07_inv02 = 1;
    38: op1_07_inv02 = 1;
    46: op1_07_inv02 = 1;
    52: op1_07_inv02 = 1;
    53: op1_07_inv02 = 1;
    55: op1_07_inv02 = 1;
    57: op1_07_inv02 = 1;
    58: op1_07_inv02 = 1;
    60: op1_07_inv02 = 1;
    63: op1_07_inv02 = 1;
    64: op1_07_inv02 = 1;
    65: op1_07_inv02 = 1;
    67: op1_07_inv02 = 1;
    69: op1_07_inv02 = 1;
    71: op1_07_inv02 = 1;
    74: op1_07_inv02 = 1;
    78: op1_07_inv02 = 1;
    82: op1_07_inv02 = 1;
    85: op1_07_inv02 = 1;
    93: op1_07_inv02 = 1;
    94: op1_07_inv02 = 1;
    95: op1_07_inv02 = 1;
    default: op1_07_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in03 = reg_0010;
    6: op1_07_in03 = imem02_in[67:64];
    7: op1_07_in03 = reg_0264;
    8: op1_07_in03 = imem00_in[95:92];
    14: op1_07_in03 = imem00_in[95:92];
    9: op1_07_in03 = reg_0579;
    10: op1_07_in03 = imem01_in[123:120];
    11: op1_07_in03 = reg_0978;
    12: op1_07_in03 = reg_0508;
    22: op1_07_in03 = reg_0508;
    13: op1_07_in03 = reg_0612;
    4: op1_07_in03 = reg_0159;
    15: op1_07_in03 = reg_1017;
    16: op1_07_in03 = imem05_in[115:112];
    17: op1_07_in03 = reg_0605;
    18: op1_07_in03 = reg_0546;
    19: op1_07_in03 = imem07_in[115:112];
    20: op1_07_in03 = imem04_in[71:68];
    52: op1_07_in03 = imem04_in[71:68];
    21: op1_07_in03 = reg_0720;
    3: op1_07_in03 = reg_0179;
    23: op1_07_in03 = reg_0343;
    24: op1_07_in03 = reg_0333;
    25: op1_07_in03 = reg_0070;
    2: op1_07_in03 = imem07_in[111:108];
    26: op1_07_in03 = reg_0679;
    27: op1_07_in03 = imem05_in[83:80];
    28: op1_07_in03 = imem06_in[111:108];
    29: op1_07_in03 = reg_0991;
    30: op1_07_in03 = reg_0067;
    31: op1_07_in03 = reg_0917;
    32: op1_07_in03 = reg_0114;
    33: op1_07_in03 = reg_0084;
    34: op1_07_in03 = reg_0956;
    35: op1_07_in03 = reg_0239;
    36: op1_07_in03 = imem00_in[115:112];
    37: op1_07_in03 = reg_0102;
    38: op1_07_in03 = reg_0544;
    39: op1_07_in03 = reg_0979;
    40: op1_07_in03 = reg_0943;
    41: op1_07_in03 = reg_1009;
    42: op1_07_in03 = reg_0695;
    43: op1_07_in03 = imem02_in[15:12];
    44: op1_07_in03 = reg_0989;
    45: op1_07_in03 = imem07_in[123:120];
    46: op1_07_in03 = imem00_in[59:56];
    47: op1_07_in03 = reg_0795;
    48: op1_07_in03 = reg_0381;
    49: op1_07_in03 = imem00_in[111:108];
    50: op1_07_in03 = reg_0727;
    51: op1_07_in03 = imem06_in[55:52];
    53: op1_07_in03 = reg_0961;
    54: op1_07_in03 = reg_0889;
    55: op1_07_in03 = reg_0706;
    56: op1_07_in03 = reg_0170;
    57: op1_07_in03 = reg_0768;
    58: op1_07_in03 = reg_1045;
    59: op1_07_in03 = reg_0843;
    60: op1_07_in03 = reg_0372;
    61: op1_07_in03 = reg_1051;
    62: op1_07_in03 = reg_0038;
    63: op1_07_in03 = reg_0047;
    64: op1_07_in03 = reg_0716;
    65: op1_07_in03 = imem00_in[107:104];
    66: op1_07_in03 = imem00_in[103:100];
    73: op1_07_in03 = imem00_in[103:100];
    85: op1_07_in03 = imem00_in[103:100];
    67: op1_07_in03 = imem00_in[39:36];
    91: op1_07_in03 = imem00_in[39:36];
    68: op1_07_in03 = reg_0608;
    69: op1_07_in03 = reg_0953;
    70: op1_07_in03 = reg_0842;
    71: op1_07_in03 = reg_0354;
    74: op1_07_in03 = imem00_in[99:96];
    75: op1_07_in03 = imem02_in[31:28];
    76: op1_07_in03 = imem04_in[95:92];
    77: op1_07_in03 = reg_0983;
    78: op1_07_in03 = reg_0044;
    79: op1_07_in03 = reg_0361;
    80: op1_07_in03 = reg_0668;
    81: op1_07_in03 = reg_0096;
    82: op1_07_in03 = imem00_in[123:120];
    83: op1_07_in03 = imem06_in[127:124];
    84: op1_07_in03 = reg_0012;
    86: op1_07_in03 = reg_0216;
    87: op1_07_in03 = reg_0657;
    88: op1_07_in03 = reg_0427;
    89: op1_07_in03 = imem05_in[47:44];
    90: op1_07_in03 = reg_0685;
    92: op1_07_in03 = reg_0186;
    93: op1_07_in03 = reg_0060;
    94: op1_07_in03 = reg_0346;
    95: op1_07_in03 = reg_0558;
    96: op1_07_in03 = imem04_in[123:120];
    97: op1_07_in03 = reg_0305;
    default: op1_07_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv03 = 1;
    8: op1_07_inv03 = 1;
    9: op1_07_inv03 = 1;
    11: op1_07_inv03 = 1;
    12: op1_07_inv03 = 1;
    13: op1_07_inv03 = 1;
    14: op1_07_inv03 = 1;
    4: op1_07_inv03 = 1;
    15: op1_07_inv03 = 1;
    16: op1_07_inv03 = 1;
    17: op1_07_inv03 = 1;
    18: op1_07_inv03 = 1;
    19: op1_07_inv03 = 1;
    20: op1_07_inv03 = 1;
    3: op1_07_inv03 = 1;
    23: op1_07_inv03 = 1;
    25: op1_07_inv03 = 1;
    2: op1_07_inv03 = 1;
    26: op1_07_inv03 = 1;
    28: op1_07_inv03 = 1;
    31: op1_07_inv03 = 1;
    34: op1_07_inv03 = 1;
    36: op1_07_inv03 = 1;
    37: op1_07_inv03 = 1;
    40: op1_07_inv03 = 1;
    41: op1_07_inv03 = 1;
    43: op1_07_inv03 = 1;
    48: op1_07_inv03 = 1;
    50: op1_07_inv03 = 1;
    51: op1_07_inv03 = 1;
    52: op1_07_inv03 = 1;
    55: op1_07_inv03 = 1;
    56: op1_07_inv03 = 1;
    60: op1_07_inv03 = 1;
    61: op1_07_inv03 = 1;
    62: op1_07_inv03 = 1;
    63: op1_07_inv03 = 1;
    64: op1_07_inv03 = 1;
    66: op1_07_inv03 = 1;
    67: op1_07_inv03 = 1;
    69: op1_07_inv03 = 1;
    70: op1_07_inv03 = 1;
    71: op1_07_inv03 = 1;
    76: op1_07_inv03 = 1;
    78: op1_07_inv03 = 1;
    80: op1_07_inv03 = 1;
    81: op1_07_inv03 = 1;
    82: op1_07_inv03 = 1;
    83: op1_07_inv03 = 1;
    84: op1_07_inv03 = 1;
    85: op1_07_inv03 = 1;
    86: op1_07_inv03 = 1;
    88: op1_07_inv03 = 1;
    90: op1_07_inv03 = 1;
    96: op1_07_inv03 = 1;
    default: op1_07_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in04 = reg_0004;
    6: op1_07_in04 = imem02_in[91:88];
    7: op1_07_in04 = reg_0251;
    8: op1_07_in04 = reg_0682;
    9: op1_07_in04 = reg_0572;
    10: op1_07_in04 = reg_0108;
    11: op1_07_in04 = reg_0975;
    12: op1_07_in04 = reg_1039;
    13: op1_07_in04 = reg_0344;
    83: op1_07_in04 = reg_0344;
    14: op1_07_in04 = reg_0679;
    4: op1_07_in04 = reg_0173;
    15: op1_07_in04 = reg_1018;
    16: op1_07_in04 = imem05_in[119:116];
    27: op1_07_in04 = imem05_in[119:116];
    17: op1_07_in04 = reg_0621;
    18: op1_07_in04 = reg_0532;
    19: op1_07_in04 = imem07_in[123:120];
    20: op1_07_in04 = imem04_in[111:108];
    21: op1_07_in04 = reg_0701;
    3: op1_07_in04 = reg_0183;
    22: op1_07_in04 = reg_0536;
    23: op1_07_in04 = reg_0362;
    24: op1_07_in04 = reg_0359;
    25: op1_07_in04 = reg_0072;
    26: op1_07_in04 = reg_0668;
    28: op1_07_in04 = reg_0577;
    29: op1_07_in04 = reg_0980;
    30: op1_07_in04 = reg_0071;
    31: op1_07_in04 = reg_0017;
    32: op1_07_in04 = reg_0106;
    33: op1_07_in04 = imem03_in[3:0];
    34: op1_07_in04 = reg_0948;
    35: op1_07_in04 = reg_0299;
    36: op1_07_in04 = imem00_in[119:116];
    85: op1_07_in04 = imem00_in[119:116];
    37: op1_07_in04 = reg_0114;
    38: op1_07_in04 = reg_0811;
    39: op1_07_in04 = reg_0993;
    40: op1_07_in04 = reg_0022;
    41: op1_07_in04 = reg_0313;
    42: op1_07_in04 = reg_0670;
    57: op1_07_in04 = reg_0670;
    90: op1_07_in04 = reg_0670;
    43: op1_07_in04 = imem02_in[31:28];
    44: op1_07_in04 = reg_0977;
    45: op1_07_in04 = reg_0716;
    46: op1_07_in04 = imem00_in[63:60];
    47: op1_07_in04 = reg_0040;
    48: op1_07_in04 = reg_0294;
    49: op1_07_in04 = reg_0681;
    50: op1_07_in04 = reg_0422;
    51: op1_07_in04 = imem06_in[59:56];
    52: op1_07_in04 = imem04_in[107:104];
    53: op1_07_in04 = reg_0953;
    54: op1_07_in04 = reg_0387;
    55: op1_07_in04 = reg_0361;
    56: op1_07_in04 = reg_0176;
    58: op1_07_in04 = reg_0253;
    59: op1_07_in04 = reg_0669;
    60: op1_07_in04 = reg_0037;
    61: op1_07_in04 = reg_0512;
    62: op1_07_in04 = reg_0051;
    63: op1_07_in04 = reg_0406;
    64: op1_07_in04 = reg_0731;
    65: op1_07_in04 = reg_0841;
    66: op1_07_in04 = imem00_in[111:108];
    67: op1_07_in04 = imem00_in[51:48];
    68: op1_07_in04 = reg_0758;
    69: op1_07_in04 = reg_0583;
    70: op1_07_in04 = reg_0069;
    71: op1_07_in04 = reg_0610;
    73: op1_07_in04 = reg_0001;
    74: op1_07_in04 = imem00_in[123:120];
    75: op1_07_in04 = imem02_in[47:44];
    76: op1_07_in04 = imem04_in[103:100];
    77: op1_07_in04 = reg_0976;
    78: op1_07_in04 = imem05_in[91:88];
    79: op1_07_in04 = reg_0175;
    80: op1_07_in04 = reg_0663;
    81: op1_07_in04 = reg_0341;
    82: op1_07_in04 = reg_0843;
    84: op1_07_in04 = reg_0099;
    86: op1_07_in04 = reg_0521;
    87: op1_07_in04 = imem06_in[55:52];
    88: op1_07_in04 = reg_0838;
    89: op1_07_in04 = reg_0636;
    91: op1_07_in04 = imem00_in[59:56];
    92: op1_07_in04 = reg_0760;
    93: op1_07_in04 = reg_0290;
    94: op1_07_in04 = reg_0342;
    95: op1_07_in04 = reg_0823;
    96: op1_07_in04 = reg_0937;
    97: op1_07_in04 = reg_0639;
    default: op1_07_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv04 = 1;
    6: op1_07_inv04 = 1;
    8: op1_07_inv04 = 1;
    12: op1_07_inv04 = 1;
    13: op1_07_inv04 = 1;
    4: op1_07_inv04 = 1;
    15: op1_07_inv04 = 1;
    16: op1_07_inv04 = 1;
    18: op1_07_inv04 = 1;
    20: op1_07_inv04 = 1;
    21: op1_07_inv04 = 1;
    3: op1_07_inv04 = 1;
    23: op1_07_inv04 = 1;
    25: op1_07_inv04 = 1;
    29: op1_07_inv04 = 1;
    30: op1_07_inv04 = 1;
    31: op1_07_inv04 = 1;
    33: op1_07_inv04 = 1;
    34: op1_07_inv04 = 1;
    37: op1_07_inv04 = 1;
    40: op1_07_inv04 = 1;
    42: op1_07_inv04 = 1;
    43: op1_07_inv04 = 1;
    45: op1_07_inv04 = 1;
    47: op1_07_inv04 = 1;
    48: op1_07_inv04 = 1;
    51: op1_07_inv04 = 1;
    57: op1_07_inv04 = 1;
    58: op1_07_inv04 = 1;
    59: op1_07_inv04 = 1;
    60: op1_07_inv04 = 1;
    62: op1_07_inv04 = 1;
    68: op1_07_inv04 = 1;
    70: op1_07_inv04 = 1;
    71: op1_07_inv04 = 1;
    73: op1_07_inv04 = 1;
    76: op1_07_inv04 = 1;
    79: op1_07_inv04 = 1;
    82: op1_07_inv04 = 1;
    85: op1_07_inv04 = 1;
    87: op1_07_inv04 = 1;
    93: op1_07_inv04 = 1;
    95: op1_07_inv04 = 1;
    default: op1_07_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in05 = imem04_in[11:8];
    6: op1_07_in05 = imem02_in[99:96];
    7: op1_07_in05 = reg_0254;
    8: op1_07_in05 = reg_0697;
    9: op1_07_in05 = reg_0569;
    10: op1_07_in05 = reg_0115;
    11: op1_07_in05 = imem04_in[43:40];
    12: op1_07_in05 = reg_0496;
    58: op1_07_in05 = reg_0496;
    13: op1_07_in05 = reg_0392;
    14: op1_07_in05 = reg_0463;
    80: op1_07_in05 = reg_0463;
    15: op1_07_in05 = reg_0123;
    16: op1_07_in05 = imem05_in[123:120];
    17: op1_07_in05 = reg_0616;
    18: op1_07_in05 = reg_0533;
    19: op1_07_in05 = reg_0722;
    20: op1_07_in05 = imem04_in[115:112];
    52: op1_07_in05 = imem04_in[115:112];
    21: op1_07_in05 = reg_0423;
    3: op1_07_in05 = reg_0178;
    22: op1_07_in05 = reg_0511;
    23: op1_07_in05 = reg_0385;
    24: op1_07_in05 = reg_0330;
    25: op1_07_in05 = reg_0015;
    26: op1_07_in05 = reg_0699;
    27: op1_07_in05 = reg_0967;
    28: op1_07_in05 = reg_0622;
    29: op1_07_in05 = reg_0974;
    30: op1_07_in05 = reg_0063;
    31: op1_07_in05 = reg_0802;
    32: op1_07_in05 = reg_0126;
    33: op1_07_in05 = imem03_in[7:4];
    34: op1_07_in05 = reg_0946;
    35: op1_07_in05 = reg_0242;
    36: op1_07_in05 = reg_0689;
    37: op1_07_in05 = reg_0107;
    38: op1_07_in05 = reg_0249;
    39: op1_07_in05 = reg_0980;
    40: op1_07_in05 = reg_0835;
    41: op1_07_in05 = reg_0078;
    42: op1_07_in05 = reg_0678;
    43: op1_07_in05 = reg_0655;
    44: op1_07_in05 = imem04_in[35:32];
    45: op1_07_in05 = reg_0731;
    46: op1_07_in05 = imem00_in[107:104];
    47: op1_07_in05 = reg_0051;
    48: op1_07_in05 = reg_0594;
    49: op1_07_in05 = reg_0686;
    85: op1_07_in05 = reg_0686;
    50: op1_07_in05 = reg_0047;
    51: op1_07_in05 = imem06_in[71:68];
    53: op1_07_in05 = reg_0972;
    54: op1_07_in05 = reg_0344;
    55: op1_07_in05 = reg_0250;
    57: op1_07_in05 = reg_0738;
    59: op1_07_in05 = reg_0476;
    60: op1_07_in05 = reg_0482;
    61: op1_07_in05 = reg_0283;
    62: op1_07_in05 = reg_0998;
    63: op1_07_in05 = reg_0532;
    64: op1_07_in05 = reg_0718;
    65: op1_07_in05 = reg_0523;
    66: op1_07_in05 = reg_0768;
    67: op1_07_in05 = imem00_in[67:64];
    68: op1_07_in05 = imem03_in[3:0];
    69: op1_07_in05 = reg_0963;
    70: op1_07_in05 = reg_0668;
    71: op1_07_in05 = reg_0740;
    73: op1_07_in05 = reg_0748;
    74: op1_07_in05 = reg_0685;
    75: op1_07_in05 = imem02_in[83:80];
    76: op1_07_in05 = reg_1006;
    77: op1_07_in05 = reg_0997;
    78: op1_07_in05 = imem05_in[99:96];
    79: op1_07_in05 = reg_0169;
    81: op1_07_in05 = reg_0279;
    82: op1_07_in05 = reg_0883;
    83: op1_07_in05 = reg_1011;
    84: op1_07_in05 = reg_0760;
    86: op1_07_in05 = reg_1017;
    87: op1_07_in05 = imem06_in[99:96];
    88: op1_07_in05 = reg_0174;
    89: op1_07_in05 = reg_0652;
    90: op1_07_in05 = reg_0356;
    91: op1_07_in05 = imem00_in[75:72];
    92: op1_07_in05 = reg_0028;
    93: op1_07_in05 = reg_0988;
    94: op1_07_in05 = reg_0756;
    95: op1_07_in05 = reg_0397;
    96: op1_07_in05 = reg_0913;
    97: op1_07_in05 = reg_0073;
    default: op1_07_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_07_inv05 = 1;
    11: op1_07_inv05 = 1;
    12: op1_07_inv05 = 1;
    15: op1_07_inv05 = 1;
    16: op1_07_inv05 = 1;
    17: op1_07_inv05 = 1;
    18: op1_07_inv05 = 1;
    19: op1_07_inv05 = 1;
    20: op1_07_inv05 = 1;
    22: op1_07_inv05 = 1;
    23: op1_07_inv05 = 1;
    24: op1_07_inv05 = 1;
    27: op1_07_inv05 = 1;
    28: op1_07_inv05 = 1;
    30: op1_07_inv05 = 1;
    31: op1_07_inv05 = 1;
    32: op1_07_inv05 = 1;
    34: op1_07_inv05 = 1;
    35: op1_07_inv05 = 1;
    36: op1_07_inv05 = 1;
    37: op1_07_inv05 = 1;
    38: op1_07_inv05 = 1;
    42: op1_07_inv05 = 1;
    43: op1_07_inv05 = 1;
    46: op1_07_inv05 = 1;
    50: op1_07_inv05 = 1;
    51: op1_07_inv05 = 1;
    52: op1_07_inv05 = 1;
    54: op1_07_inv05 = 1;
    59: op1_07_inv05 = 1;
    60: op1_07_inv05 = 1;
    64: op1_07_inv05 = 1;
    65: op1_07_inv05 = 1;
    66: op1_07_inv05 = 1;
    67: op1_07_inv05 = 1;
    70: op1_07_inv05 = 1;
    73: op1_07_inv05 = 1;
    76: op1_07_inv05 = 1;
    79: op1_07_inv05 = 1;
    80: op1_07_inv05 = 1;
    81: op1_07_inv05 = 1;
    82: op1_07_inv05 = 1;
    85: op1_07_inv05 = 1;
    90: op1_07_inv05 = 1;
    92: op1_07_inv05 = 1;
    93: op1_07_inv05 = 1;
    96: op1_07_inv05 = 1;
    97: op1_07_inv05 = 1;
    default: op1_07_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in06 = imem04_in[31:28];
    6: op1_07_in06 = imem02_in[119:116];
    7: op1_07_in06 = reg_0148;
    8: op1_07_in06 = reg_0681;
    9: op1_07_in06 = reg_0600;
    10: op1_07_in06 = reg_0109;
    11: op1_07_in06 = reg_0536;
    52: op1_07_in06 = reg_0536;
    12: op1_07_in06 = reg_1043;
    13: op1_07_in06 = reg_0390;
    14: op1_07_in06 = reg_0461;
    15: op1_07_in06 = reg_0124;
    16: op1_07_in06 = reg_0971;
    17: op1_07_in06 = reg_0626;
    18: op1_07_in06 = reg_0531;
    19: op1_07_in06 = reg_0719;
    20: op1_07_in06 = reg_0545;
    21: op1_07_in06 = reg_0428;
    22: op1_07_in06 = reg_0277;
    23: op1_07_in06 = reg_0322;
    24: op1_07_in06 = reg_0346;
    25: op1_07_in06 = reg_0054;
    26: op1_07_in06 = reg_0455;
    27: op1_07_in06 = reg_0957;
    28: op1_07_in06 = reg_0601;
    29: op1_07_in06 = reg_0975;
    30: op1_07_in06 = reg_0072;
    31: op1_07_in06 = imem07_in[71:68];
    32: op1_07_in06 = imem02_in[75:72];
    33: op1_07_in06 = imem03_in[27:24];
    34: op1_07_in06 = reg_0947;
    35: op1_07_in06 = reg_0555;
    36: op1_07_in06 = reg_0684;
    74: op1_07_in06 = reg_0684;
    37: op1_07_in06 = reg_0121;
    38: op1_07_in06 = reg_1042;
    39: op1_07_in06 = imem04_in[19:16];
    40: op1_07_in06 = reg_0900;
    41: op1_07_in06 = reg_0070;
    42: op1_07_in06 = reg_0688;
    43: op1_07_in06 = reg_0653;
    44: op1_07_in06 = imem04_in[83:80];
    45: op1_07_in06 = reg_0714;
    46: op1_07_in06 = imem00_in[111:108];
    47: op1_07_in06 = reg_0312;
    48: op1_07_in06 = reg_0241;
    49: op1_07_in06 = reg_0677;
    50: op1_07_in06 = reg_0744;
    64: op1_07_in06 = reg_0744;
    51: op1_07_in06 = imem06_in[87:84];
    53: op1_07_in06 = reg_0032;
    54: op1_07_in06 = reg_0381;
    55: op1_07_in06 = reg_0419;
    57: op1_07_in06 = reg_0883;
    58: op1_07_in06 = reg_0798;
    59: op1_07_in06 = reg_0466;
    60: op1_07_in06 = reg_0758;
    61: op1_07_in06 = reg_0117;
    62: op1_07_in06 = reg_0992;
    63: op1_07_in06 = reg_0589;
    65: op1_07_in06 = reg_0753;
    66: op1_07_in06 = reg_0523;
    67: op1_07_in06 = imem00_in[83:80];
    68: op1_07_in06 = imem03_in[11:8];
    69: op1_07_in06 = reg_0940;
    70: op1_07_in06 = reg_0477;
    71: op1_07_in06 = reg_0832;
    73: op1_07_in06 = reg_0738;
    75: op1_07_in06 = imem02_in[127:124];
    76: op1_07_in06 = reg_0511;
    77: op1_07_in06 = imem04_in[67:64];
    78: op1_07_in06 = reg_1021;
    79: op1_07_in06 = reg_0177;
    80: op1_07_in06 = reg_0450;
    81: op1_07_in06 = reg_0441;
    82: op1_07_in06 = reg_0069;
    83: op1_07_in06 = reg_0392;
    84: op1_07_in06 = reg_0228;
    85: op1_07_in06 = reg_0828;
    86: op1_07_in06 = reg_1033;
    87: op1_07_in06 = imem06_in[103:100];
    88: op1_07_in06 = reg_0172;
    89: op1_07_in06 = reg_0013;
    90: op1_07_in06 = reg_0451;
    91: op1_07_in06 = imem00_in[87:84];
    92: op1_07_in06 = reg_0460;
    93: op1_07_in06 = imem04_in[11:8];
    94: op1_07_in06 = reg_0397;
    95: op1_07_in06 = reg_0596;
    96: op1_07_in06 = reg_0123;
    97: op1_07_in06 = reg_0855;
    default: op1_07_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv06 = 1;
    6: op1_07_inv06 = 1;
    8: op1_07_inv06 = 1;
    9: op1_07_inv06 = 1;
    10: op1_07_inv06 = 1;
    12: op1_07_inv06 = 1;
    13: op1_07_inv06 = 1;
    14: op1_07_inv06 = 1;
    16: op1_07_inv06 = 1;
    17: op1_07_inv06 = 1;
    19: op1_07_inv06 = 1;
    20: op1_07_inv06 = 1;
    24: op1_07_inv06 = 1;
    25: op1_07_inv06 = 1;
    30: op1_07_inv06 = 1;
    31: op1_07_inv06 = 1;
    32: op1_07_inv06 = 1;
    33: op1_07_inv06 = 1;
    34: op1_07_inv06 = 1;
    36: op1_07_inv06 = 1;
    37: op1_07_inv06 = 1;
    38: op1_07_inv06 = 1;
    40: op1_07_inv06 = 1;
    42: op1_07_inv06 = 1;
    43: op1_07_inv06 = 1;
    45: op1_07_inv06 = 1;
    48: op1_07_inv06 = 1;
    51: op1_07_inv06 = 1;
    52: op1_07_inv06 = 1;
    53: op1_07_inv06 = 1;
    58: op1_07_inv06 = 1;
    59: op1_07_inv06 = 1;
    60: op1_07_inv06 = 1;
    61: op1_07_inv06 = 1;
    63: op1_07_inv06 = 1;
    66: op1_07_inv06 = 1;
    67: op1_07_inv06 = 1;
    68: op1_07_inv06 = 1;
    70: op1_07_inv06 = 1;
    73: op1_07_inv06 = 1;
    75: op1_07_inv06 = 1;
    81: op1_07_inv06 = 1;
    82: op1_07_inv06 = 1;
    83: op1_07_inv06 = 1;
    84: op1_07_inv06 = 1;
    85: op1_07_inv06 = 1;
    87: op1_07_inv06 = 1;
    88: op1_07_inv06 = 1;
    90: op1_07_inv06 = 1;
    91: op1_07_inv06 = 1;
    93: op1_07_inv06 = 1;
    94: op1_07_inv06 = 1;
    95: op1_07_inv06 = 1;
    97: op1_07_inv06 = 1;
    default: op1_07_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in07 = imem04_in[59:56];
    6: op1_07_in07 = reg_0658;
    7: op1_07_in07 = reg_0145;
    8: op1_07_in07 = reg_0698;
    9: op1_07_in07 = reg_0581;
    10: op1_07_in07 = reg_0126;
    11: op1_07_in07 = reg_0553;
    12: op1_07_in07 = reg_1033;
    13: op1_07_in07 = reg_1010;
    14: op1_07_in07 = reg_0466;
    15: op1_07_in07 = reg_0116;
    16: op1_07_in07 = reg_0944;
    17: op1_07_in07 = reg_0619;
    18: op1_07_in07 = reg_0556;
    19: op1_07_in07 = reg_0720;
    20: op1_07_in07 = reg_0542;
    21: op1_07_in07 = reg_0434;
    22: op1_07_in07 = imem04_in[19:16];
    93: op1_07_in07 = imem04_in[19:16];
    23: op1_07_in07 = reg_0323;
    24: op1_07_in07 = reg_0338;
    25: op1_07_in07 = reg_0047;
    26: op1_07_in07 = reg_0472;
    27: op1_07_in07 = reg_0948;
    28: op1_07_in07 = reg_0402;
    29: op1_07_in07 = reg_0994;
    30: op1_07_in07 = reg_0058;
    31: op1_07_in07 = imem07_in[91:88];
    32: op1_07_in07 = imem02_in[79:76];
    33: op1_07_in07 = imem03_in[35:32];
    34: op1_07_in07 = reg_0943;
    35: op1_07_in07 = reg_0860;
    36: op1_07_in07 = reg_0679;
    37: op1_07_in07 = imem02_in[39:36];
    38: op1_07_in07 = reg_0869;
    39: op1_07_in07 = imem04_in[27:24];
    40: op1_07_in07 = reg_0806;
    41: op1_07_in07 = reg_0044;
    42: op1_07_in07 = reg_0692;
    43: op1_07_in07 = reg_0661;
    44: op1_07_in07 = reg_0530;
    45: op1_07_in07 = reg_0724;
    46: op1_07_in07 = reg_0682;
    47: op1_07_in07 = reg_0844;
    48: op1_07_in07 = imem07_in[7:4];
    49: op1_07_in07 = reg_0671;
    50: op1_07_in07 = reg_0315;
    51: op1_07_in07 = reg_0883;
    66: op1_07_in07 = reg_0883;
    52: op1_07_in07 = reg_0301;
    53: op1_07_in07 = reg_0774;
    54: op1_07_in07 = reg_0388;
    55: op1_07_in07 = reg_0420;
    57: op1_07_in07 = reg_0680;
    58: op1_07_in07 = reg_0514;
    59: op1_07_in07 = reg_0467;
    60: op1_07_in07 = reg_0088;
    61: op1_07_in07 = imem02_in[19:16];
    62: op1_07_in07 = reg_0980;
    63: op1_07_in07 = reg_0180;
    64: op1_07_in07 = reg_0640;
    65: op1_07_in07 = reg_0455;
    67: op1_07_in07 = imem00_in[99:96];
    91: op1_07_in07 = imem00_in[99:96];
    68: op1_07_in07 = imem03_in[67:64];
    69: op1_07_in07 = reg_0274;
    70: op1_07_in07 = reg_0476;
    80: op1_07_in07 = reg_0476;
    71: op1_07_in07 = reg_0111;
    73: op1_07_in07 = reg_0477;
    74: op1_07_in07 = reg_0499;
    75: op1_07_in07 = reg_0637;
    76: op1_07_in07 = reg_0912;
    77: op1_07_in07 = imem04_in[83:80];
    78: op1_07_in07 = reg_0655;
    79: op1_07_in07 = reg_0168;
    81: op1_07_in07 = reg_0664;
    82: op1_07_in07 = reg_0687;
    83: op1_07_in07 = reg_0863;
    84: op1_07_in07 = reg_0445;
    85: op1_07_in07 = reg_0669;
    86: op1_07_in07 = reg_0101;
    87: op1_07_in07 = reg_0010;
    88: op1_07_in07 = reg_0731;
    89: op1_07_in07 = reg_0137;
    90: op1_07_in07 = reg_0470;
    92: op1_07_in07 = reg_0480;
    94: op1_07_in07 = reg_0060;
    95: op1_07_in07 = reg_0773;
    96: op1_07_in07 = reg_0066;
    97: op1_07_in07 = reg_0095;
    default: op1_07_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv07 = 1;
    12: op1_07_inv07 = 1;
    13: op1_07_inv07 = 1;
    16: op1_07_inv07 = 1;
    20: op1_07_inv07 = 1;
    23: op1_07_inv07 = 1;
    26: op1_07_inv07 = 1;
    28: op1_07_inv07 = 1;
    30: op1_07_inv07 = 1;
    32: op1_07_inv07 = 1;
    33: op1_07_inv07 = 1;
    35: op1_07_inv07 = 1;
    37: op1_07_inv07 = 1;
    41: op1_07_inv07 = 1;
    45: op1_07_inv07 = 1;
    46: op1_07_inv07 = 1;
    47: op1_07_inv07 = 1;
    49: op1_07_inv07 = 1;
    51: op1_07_inv07 = 1;
    54: op1_07_inv07 = 1;
    58: op1_07_inv07 = 1;
    62: op1_07_inv07 = 1;
    63: op1_07_inv07 = 1;
    68: op1_07_inv07 = 1;
    71: op1_07_inv07 = 1;
    73: op1_07_inv07 = 1;
    76: op1_07_inv07 = 1;
    79: op1_07_inv07 = 1;
    80: op1_07_inv07 = 1;
    81: op1_07_inv07 = 1;
    83: op1_07_inv07 = 1;
    85: op1_07_inv07 = 1;
    91: op1_07_inv07 = 1;
    93: op1_07_inv07 = 1;
    96: op1_07_inv07 = 1;
    default: op1_07_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in08 = imem04_in[67:64];
    6: op1_07_in08 = reg_0654;
    7: op1_07_in08 = reg_0143;
    8: op1_07_in08 = reg_0670;
    9: op1_07_in08 = reg_0595;
    10: op1_07_in08 = reg_0110;
    11: op1_07_in08 = reg_0550;
    12: op1_07_in08 = reg_1015;
    13: op1_07_in08 = reg_1011;
    14: op1_07_in08 = reg_0460;
    80: op1_07_in08 = reg_0460;
    15: op1_07_in08 = reg_0101;
    16: op1_07_in08 = reg_0972;
    17: op1_07_in08 = reg_0608;
    18: op1_07_in08 = reg_0303;
    19: op1_07_in08 = reg_0729;
    45: op1_07_in08 = reg_0729;
    20: op1_07_in08 = reg_0554;
    21: op1_07_in08 = reg_0444;
    22: op1_07_in08 = imem04_in[27:24];
    23: op1_07_in08 = reg_0998;
    24: op1_07_in08 = reg_0355;
    25: op1_07_in08 = reg_0517;
    26: op1_07_in08 = reg_0467;
    92: op1_07_in08 = reg_0467;
    27: op1_07_in08 = reg_0949;
    28: op1_07_in08 = reg_0404;
    29: op1_07_in08 = imem04_in[11:8];
    30: op1_07_in08 = reg_0286;
    31: op1_07_in08 = imem07_in[95:92];
    32: op1_07_in08 = imem02_in[91:88];
    33: op1_07_in08 = imem03_in[39:36];
    34: op1_07_in08 = reg_0834;
    35: op1_07_in08 = reg_0248;
    36: op1_07_in08 = reg_0463;
    57: op1_07_in08 = reg_0463;
    37: op1_07_in08 = imem02_in[47:44];
    38: op1_07_in08 = reg_0885;
    39: op1_07_in08 = imem04_in[55:52];
    40: op1_07_in08 = reg_0252;
    41: op1_07_in08 = imem05_in[55:52];
    42: op1_07_in08 = reg_0455;
    82: op1_07_in08 = reg_0455;
    43: op1_07_in08 = reg_0656;
    44: op1_07_in08 = reg_0265;
    46: op1_07_in08 = reg_0693;
    47: op1_07_in08 = reg_0822;
    48: op1_07_in08 = imem07_in[15:12];
    49: op1_07_in08 = reg_0454;
    50: op1_07_in08 = reg_0641;
    51: op1_07_in08 = reg_0895;
    52: op1_07_in08 = reg_0530;
    53: op1_07_in08 = reg_0436;
    54: op1_07_in08 = reg_0628;
    55: op1_07_in08 = reg_0427;
    58: op1_07_in08 = reg_0830;
    59: op1_07_in08 = reg_0200;
    60: op1_07_in08 = reg_0761;
    61: op1_07_in08 = imem02_in[43:40];
    62: op1_07_in08 = reg_0989;
    63: op1_07_in08 = reg_0181;
    64: op1_07_in08 = reg_0180;
    65: op1_07_in08 = reg_0461;
    66: op1_07_in08 = reg_0499;
    67: op1_07_in08 = reg_0843;
    68: op1_07_in08 = imem03_in[91:88];
    69: op1_07_in08 = reg_0819;
    70: op1_07_in08 = reg_0475;
    71: op1_07_in08 = reg_0555;
    73: op1_07_in08 = reg_0452;
    74: op1_07_in08 = reg_0477;
    75: op1_07_in08 = reg_0649;
    76: op1_07_in08 = reg_0539;
    77: op1_07_in08 = imem04_in[99:96];
    78: op1_07_in08 = reg_0935;
    79: op1_07_in08 = reg_0170;
    81: op1_07_in08 = reg_0329;
    83: op1_07_in08 = reg_0804;
    84: op1_07_in08 = reg_0346;
    85: op1_07_in08 = reg_0457;
    86: op1_07_in08 = reg_0115;
    87: op1_07_in08 = reg_1019;
    88: op1_07_in08 = reg_0182;
    89: op1_07_in08 = reg_0256;
    90: op1_07_in08 = reg_0189;
    91: op1_07_in08 = imem00_in[115:112];
    93: op1_07_in08 = imem04_in[51:48];
    94: op1_07_in08 = reg_0987;
    95: op1_07_in08 = reg_0377;
    96: op1_07_in08 = reg_0401;
    97: op1_07_in08 = reg_0418;
    default: op1_07_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_07_inv08 = 1;
    8: op1_07_inv08 = 1;
    12: op1_07_inv08 = 1;
    13: op1_07_inv08 = 1;
    14: op1_07_inv08 = 1;
    15: op1_07_inv08 = 1;
    16: op1_07_inv08 = 1;
    18: op1_07_inv08 = 1;
    21: op1_07_inv08 = 1;
    24: op1_07_inv08 = 1;
    25: op1_07_inv08 = 1;
    34: op1_07_inv08 = 1;
    36: op1_07_inv08 = 1;
    37: op1_07_inv08 = 1;
    38: op1_07_inv08 = 1;
    39: op1_07_inv08 = 1;
    40: op1_07_inv08 = 1;
    44: op1_07_inv08 = 1;
    45: op1_07_inv08 = 1;
    48: op1_07_inv08 = 1;
    50: op1_07_inv08 = 1;
    51: op1_07_inv08 = 1;
    52: op1_07_inv08 = 1;
    53: op1_07_inv08 = 1;
    57: op1_07_inv08 = 1;
    58: op1_07_inv08 = 1;
    59: op1_07_inv08 = 1;
    65: op1_07_inv08 = 1;
    66: op1_07_inv08 = 1;
    71: op1_07_inv08 = 1;
    74: op1_07_inv08 = 1;
    75: op1_07_inv08 = 1;
    76: op1_07_inv08 = 1;
    77: op1_07_inv08 = 1;
    80: op1_07_inv08 = 1;
    82: op1_07_inv08 = 1;
    85: op1_07_inv08 = 1;
    86: op1_07_inv08 = 1;
    88: op1_07_inv08 = 1;
    91: op1_07_inv08 = 1;
    94: op1_07_inv08 = 1;
    default: op1_07_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in09 = imem04_in[79:76];
    6: op1_07_in09 = reg_0637;
    7: op1_07_in09 = imem06_in[35:32];
    8: op1_07_in09 = reg_0677;
    9: op1_07_in09 = reg_0360;
    10: op1_07_in09 = imem02_in[3:0];
    11: op1_07_in09 = reg_0531;
    12: op1_07_in09 = reg_0871;
    13: op1_07_in09 = reg_0754;
    14: op1_07_in09 = reg_0481;
    70: op1_07_in09 = reg_0481;
    85: op1_07_in09 = reg_0481;
    15: op1_07_in09 = reg_0109;
    86: op1_07_in09 = reg_0109;
    16: op1_07_in09 = reg_0863;
    17: op1_07_in09 = reg_0622;
    18: op1_07_in09 = reg_0305;
    19: op1_07_in09 = reg_0713;
    20: op1_07_in09 = reg_0551;
    21: op1_07_in09 = reg_0438;
    22: op1_07_in09 = imem04_in[51:48];
    23: op1_07_in09 = reg_0996;
    24: op1_07_in09 = reg_0347;
    25: op1_07_in09 = reg_0286;
    26: op1_07_in09 = reg_0479;
    27: op1_07_in09 = reg_0945;
    28: op1_07_in09 = reg_0401;
    29: op1_07_in09 = imem04_in[47:44];
    30: op1_07_in09 = imem05_in[103:100];
    31: op1_07_in09 = imem07_in[127:124];
    32: op1_07_in09 = imem02_in[127:124];
    33: op1_07_in09 = imem03_in[51:48];
    34: op1_07_in09 = reg_0215;
    35: op1_07_in09 = reg_0274;
    36: op1_07_in09 = reg_0464;
    37: op1_07_in09 = imem02_in[87:84];
    38: op1_07_in09 = reg_1044;
    39: op1_07_in09 = imem04_in[127:124];
    40: op1_07_in09 = reg_0813;
    41: op1_07_in09 = imem05_in[87:84];
    42: op1_07_in09 = reg_0466;
    43: op1_07_in09 = reg_0648;
    44: op1_07_in09 = reg_1009;
    45: op1_07_in09 = reg_0711;
    46: op1_07_in09 = reg_0683;
    47: op1_07_in09 = reg_0987;
    48: op1_07_in09 = imem07_in[31:28];
    49: op1_07_in09 = reg_0457;
    50: op1_07_in09 = reg_0350;
    51: op1_07_in09 = reg_0220;
    52: op1_07_in09 = reg_0937;
    53: op1_07_in09 = reg_0333;
    54: op1_07_in09 = reg_0894;
    55: op1_07_in09 = reg_0502;
    57: op1_07_in09 = reg_0450;
    58: op1_07_in09 = reg_0216;
    59: op1_07_in09 = reg_0210;
    60: op1_07_in09 = reg_0085;
    61: op1_07_in09 = imem02_in[51:48];
    62: op1_07_in09 = reg_0976;
    63: op1_07_in09 = reg_0179;
    64: op1_07_in09 = reg_0172;
    65: op1_07_in09 = reg_0469;
    82: op1_07_in09 = reg_0469;
    66: op1_07_in09 = reg_0102;
    67: op1_07_in09 = reg_0738;
    68: op1_07_in09 = imem03_in[95:92];
    69: op1_07_in09 = reg_0132;
    71: op1_07_in09 = reg_0860;
    73: op1_07_in09 = reg_0456;
    74: op1_07_in09 = reg_0473;
    75: op1_07_in09 = reg_0907;
    76: op1_07_in09 = reg_0048;
    77: op1_07_in09 = reg_1004;
    78: op1_07_in09 = reg_0956;
    79: op1_07_in09 = reg_0173;
    80: op1_07_in09 = reg_0208;
    81: op1_07_in09 = reg_0368;
    83: op1_07_in09 = reg_0857;
    84: op1_07_in09 = reg_0662;
    87: op1_07_in09 = reg_0691;
    88: op1_07_in09 = reg_0371;
    89: op1_07_in09 = reg_0259;
    90: op1_07_in09 = reg_0204;
    91: op1_07_in09 = reg_0455;
    92: op1_07_in09 = reg_0474;
    93: op1_07_in09 = imem04_in[55:52];
    94: op1_07_in09 = reg_0373;
    95: op1_07_in09 = reg_0376;
    96: op1_07_in09 = reg_0296;
    97: op1_07_in09 = reg_0837;
    default: op1_07_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv09 = 1;
    14: op1_07_inv09 = 1;
    15: op1_07_inv09 = 1;
    18: op1_07_inv09 = 1;
    21: op1_07_inv09 = 1;
    23: op1_07_inv09 = 1;
    24: op1_07_inv09 = 1;
    25: op1_07_inv09 = 1;
    26: op1_07_inv09 = 1;
    27: op1_07_inv09 = 1;
    28: op1_07_inv09 = 1;
    31: op1_07_inv09 = 1;
    32: op1_07_inv09 = 1;
    35: op1_07_inv09 = 1;
    36: op1_07_inv09 = 1;
    37: op1_07_inv09 = 1;
    39: op1_07_inv09 = 1;
    41: op1_07_inv09 = 1;
    44: op1_07_inv09 = 1;
    45: op1_07_inv09 = 1;
    46: op1_07_inv09 = 1;
    47: op1_07_inv09 = 1;
    48: op1_07_inv09 = 1;
    49: op1_07_inv09 = 1;
    50: op1_07_inv09 = 1;
    51: op1_07_inv09 = 1;
    52: op1_07_inv09 = 1;
    53: op1_07_inv09 = 1;
    55: op1_07_inv09 = 1;
    58: op1_07_inv09 = 1;
    59: op1_07_inv09 = 1;
    64: op1_07_inv09 = 1;
    65: op1_07_inv09 = 1;
    67: op1_07_inv09 = 1;
    69: op1_07_inv09 = 1;
    70: op1_07_inv09 = 1;
    73: op1_07_inv09 = 1;
    78: op1_07_inv09 = 1;
    79: op1_07_inv09 = 1;
    80: op1_07_inv09 = 1;
    82: op1_07_inv09 = 1;
    83: op1_07_inv09 = 1;
    85: op1_07_inv09 = 1;
    90: op1_07_inv09 = 1;
    92: op1_07_inv09 = 1;
    93: op1_07_inv09 = 1;
    94: op1_07_inv09 = 1;
    96: op1_07_inv09 = 1;
    default: op1_07_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in10 = imem04_in[99:96];
    6: op1_07_in10 = reg_0649;
    43: op1_07_in10 = reg_0649;
    7: op1_07_in10 = imem06_in[67:64];
    8: op1_07_in10 = reg_0691;
    9: op1_07_in10 = reg_0311;
    10: op1_07_in10 = imem02_in[67:64];
    11: op1_07_in10 = reg_0541;
    20: op1_07_in10 = reg_0541;
    12: op1_07_in10 = reg_1018;
    13: op1_07_in10 = imem07_in[7:4];
    14: op1_07_in10 = reg_0480;
    70: op1_07_in10 = reg_0480;
    15: op1_07_in10 = reg_0110;
    16: op1_07_in10 = reg_0215;
    17: op1_07_in10 = reg_0601;
    18: op1_07_in10 = imem04_in[31:28];
    19: op1_07_in10 = reg_0425;
    21: op1_07_in10 = reg_0448;
    22: op1_07_in10 = imem04_in[87:84];
    23: op1_07_in10 = reg_0993;
    24: op1_07_in10 = reg_0792;
    25: op1_07_in10 = imem05_in[23:20];
    26: op1_07_in10 = reg_0478;
    27: op1_07_in10 = reg_0946;
    28: op1_07_in10 = reg_1030;
    29: op1_07_in10 = imem04_in[103:100];
    30: op1_07_in10 = reg_0948;
    31: op1_07_in10 = reg_0704;
    32: op1_07_in10 = reg_0658;
    33: op1_07_in10 = imem03_in[59:56];
    34: op1_07_in10 = reg_0835;
    35: op1_07_in10 = reg_0544;
    36: op1_07_in10 = reg_0466;
    37: op1_07_in10 = imem02_in[111:108];
    38: op1_07_in10 = reg_1037;
    39: op1_07_in10 = reg_0530;
    40: op1_07_in10 = reg_0152;
    41: op1_07_in10 = imem05_in[115:112];
    42: op1_07_in10 = reg_0472;
    85: op1_07_in10 = reg_0472;
    44: op1_07_in10 = reg_0931;
    45: op1_07_in10 = reg_0727;
    46: op1_07_in10 = reg_0685;
    47: op1_07_in10 = reg_0981;
    48: op1_07_in10 = imem07_in[43:40];
    49: op1_07_in10 = reg_0470;
    65: op1_07_in10 = reg_0470;
    50: op1_07_in10 = reg_0427;
    51: op1_07_in10 = reg_0533;
    52: op1_07_in10 = reg_0055;
    53: op1_07_in10 = reg_0142;
    54: op1_07_in10 = reg_0596;
    55: op1_07_in10 = reg_0160;
    57: op1_07_in10 = reg_0474;
    58: op1_07_in10 = reg_1040;
    59: op1_07_in10 = reg_0203;
    60: op1_07_in10 = reg_0016;
    61: op1_07_in10 = imem02_in[99:96];
    62: op1_07_in10 = imem04_in[7:4];
    63: op1_07_in10 = reg_0169;
    64: op1_07_in10 = reg_0181;
    66: op1_07_in10 = reg_0464;
    67: op1_07_in10 = reg_0356;
    68: op1_07_in10 = imem03_in[103:100];
    69: op1_07_in10 = reg_0136;
    71: op1_07_in10 = reg_0109;
    73: op1_07_in10 = reg_0201;
    74: op1_07_in10 = reg_0467;
    75: op1_07_in10 = reg_0095;
    76: op1_07_in10 = reg_0848;
    77: op1_07_in10 = reg_0536;
    78: op1_07_in10 = reg_0135;
    80: op1_07_in10 = reg_0194;
    81: op1_07_in10 = reg_0372;
    82: op1_07_in10 = reg_0475;
    83: op1_07_in10 = reg_0381;
    84: op1_07_in10 = reg_0278;
    86: op1_07_in10 = reg_0103;
    87: op1_07_in10 = reg_0294;
    89: op1_07_in10 = reg_0956;
    90: op1_07_in10 = reg_0198;
    91: op1_07_in10 = reg_0457;
    92: op1_07_in10 = reg_0471;
    93: op1_07_in10 = imem04_in[71:68];
    94: op1_07_in10 = reg_0445;
    95: op1_07_in10 = reg_0597;
    96: op1_07_in10 = reg_0432;
    97: op1_07_in10 = reg_0323;
    default: op1_07_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv10 = 1;
    11: op1_07_inv10 = 1;
    14: op1_07_inv10 = 1;
    15: op1_07_inv10 = 1;
    16: op1_07_inv10 = 1;
    17: op1_07_inv10 = 1;
    18: op1_07_inv10 = 1;
    20: op1_07_inv10 = 1;
    22: op1_07_inv10 = 1;
    23: op1_07_inv10 = 1;
    24: op1_07_inv10 = 1;
    25: op1_07_inv10 = 1;
    27: op1_07_inv10 = 1;
    28: op1_07_inv10 = 1;
    30: op1_07_inv10 = 1;
    31: op1_07_inv10 = 1;
    32: op1_07_inv10 = 1;
    35: op1_07_inv10 = 1;
    38: op1_07_inv10 = 1;
    41: op1_07_inv10 = 1;
    42: op1_07_inv10 = 1;
    43: op1_07_inv10 = 1;
    47: op1_07_inv10 = 1;
    48: op1_07_inv10 = 1;
    49: op1_07_inv10 = 1;
    50: op1_07_inv10 = 1;
    51: op1_07_inv10 = 1;
    57: op1_07_inv10 = 1;
    58: op1_07_inv10 = 1;
    63: op1_07_inv10 = 1;
    64: op1_07_inv10 = 1;
    65: op1_07_inv10 = 1;
    66: op1_07_inv10 = 1;
    67: op1_07_inv10 = 1;
    69: op1_07_inv10 = 1;
    77: op1_07_inv10 = 1;
    78: op1_07_inv10 = 1;
    80: op1_07_inv10 = 1;
    82: op1_07_inv10 = 1;
    85: op1_07_inv10 = 1;
    86: op1_07_inv10 = 1;
    87: op1_07_inv10 = 1;
    90: op1_07_inv10 = 1;
    91: op1_07_inv10 = 1;
    94: op1_07_inv10 = 1;
    97: op1_07_inv10 = 1;
    default: op1_07_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in11 = imem04_in[103:100];
    93: op1_07_in11 = imem04_in[103:100];
    6: op1_07_in11 = reg_0643;
    7: op1_07_in11 = imem06_in[75:72];
    8: op1_07_in11 = reg_0450;
    9: op1_07_in11 = reg_0385;
    10: op1_07_in11 = imem02_in[111:108];
    11: op1_07_in11 = reg_0301;
    12: op1_07_in11 = reg_0123;
    13: op1_07_in11 = imem07_in[27:24];
    14: op1_07_in11 = reg_0467;
    15: op1_07_in11 = imem02_in[31:28];
    16: op1_07_in11 = reg_0835;
    17: op1_07_in11 = reg_0379;
    18: op1_07_in11 = imem04_in[43:40];
    19: op1_07_in11 = reg_0429;
    20: op1_07_in11 = reg_0259;
    21: op1_07_in11 = reg_0166;
    22: op1_07_in11 = imem04_in[91:88];
    23: op1_07_in11 = imem04_in[51:48];
    24: op1_07_in11 = reg_0084;
    25: op1_07_in11 = reg_0967;
    26: op1_07_in11 = reg_0204;
    27: op1_07_in11 = reg_0953;
    28: op1_07_in11 = reg_0027;
    29: op1_07_in11 = reg_0536;
    30: op1_07_in11 = reg_0215;
    31: op1_07_in11 = reg_0714;
    32: op1_07_in11 = reg_0666;
    33: op1_07_in11 = imem03_in[103:100];
    34: op1_07_in11 = reg_0831;
    35: op1_07_in11 = reg_0221;
    36: op1_07_in11 = reg_0480;
    37: op1_07_in11 = imem02_in[115:112];
    38: op1_07_in11 = reg_0227;
    39: op1_07_in11 = reg_0306;
    40: op1_07_in11 = reg_0146;
    53: op1_07_in11 = reg_0146;
    41: op1_07_in11 = reg_0970;
    42: op1_07_in11 = reg_0459;
    49: op1_07_in11 = reg_0459;
    43: op1_07_in11 = reg_0662;
    44: op1_07_in11 = reg_0507;
    45: op1_07_in11 = reg_0002;
    46: op1_07_in11 = reg_0672;
    47: op1_07_in11 = reg_0975;
    48: op1_07_in11 = imem07_in[51:48];
    50: op1_07_in11 = reg_0161;
    64: op1_07_in11 = reg_0161;
    51: op1_07_in11 = reg_0348;
    52: op1_07_in11 = reg_0778;
    54: op1_07_in11 = reg_0631;
    55: op1_07_in11 = reg_0185;
    57: op1_07_in11 = reg_0479;
    85: op1_07_in11 = reg_0479;
    58: op1_07_in11 = reg_0902;
    59: op1_07_in11 = reg_0207;
    60: op1_07_in11 = imem03_in[31:28];
    61: op1_07_in11 = reg_0639;
    62: op1_07_in11 = imem04_in[39:36];
    63: op1_07_in11 = reg_0163;
    65: op1_07_in11 = reg_0474;
    66: op1_07_in11 = reg_0462;
    67: op1_07_in11 = reg_0069;
    68: op1_07_in11 = imem03_in[107:104];
    69: op1_07_in11 = reg_0140;
    70: op1_07_in11 = reg_0208;
    71: op1_07_in11 = reg_0117;
    73: op1_07_in11 = imem01_in[27:24];
    74: op1_07_in11 = reg_0470;
    75: op1_07_in11 = reg_0279;
    76: op1_07_in11 = reg_0524;
    77: op1_07_in11 = reg_0282;
    78: op1_07_in11 = reg_0252;
    80: op1_07_in11 = reg_0196;
    81: op1_07_in11 = reg_0608;
    82: op1_07_in11 = reg_0481;
    83: op1_07_in11 = reg_0220;
    84: op1_07_in11 = reg_0239;
    86: op1_07_in11 = reg_0821;
    87: op1_07_in11 = reg_0391;
    89: op1_07_in11 = reg_0892;
    90: op1_07_in11 = reg_0190;
    91: op1_07_in11 = reg_0461;
    92: op1_07_in11 = reg_0203;
    94: op1_07_in11 = reg_0825;
    95: op1_07_in11 = reg_0581;
    96: op1_07_in11 = reg_0552;
    97: op1_07_in11 = reg_0358;
    default: op1_07_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_07_inv11 = 1;
    9: op1_07_inv11 = 1;
    10: op1_07_inv11 = 1;
    13: op1_07_inv11 = 1;
    14: op1_07_inv11 = 1;
    17: op1_07_inv11 = 1;
    18: op1_07_inv11 = 1;
    19: op1_07_inv11 = 1;
    20: op1_07_inv11 = 1;
    22: op1_07_inv11 = 1;
    24: op1_07_inv11 = 1;
    26: op1_07_inv11 = 1;
    27: op1_07_inv11 = 1;
    29: op1_07_inv11 = 1;
    30: op1_07_inv11 = 1;
    31: op1_07_inv11 = 1;
    32: op1_07_inv11 = 1;
    35: op1_07_inv11 = 1;
    36: op1_07_inv11 = 1;
    38: op1_07_inv11 = 1;
    44: op1_07_inv11 = 1;
    46: op1_07_inv11 = 1;
    47: op1_07_inv11 = 1;
    48: op1_07_inv11 = 1;
    50: op1_07_inv11 = 1;
    58: op1_07_inv11 = 1;
    59: op1_07_inv11 = 1;
    60: op1_07_inv11 = 1;
    61: op1_07_inv11 = 1;
    63: op1_07_inv11 = 1;
    64: op1_07_inv11 = 1;
    67: op1_07_inv11 = 1;
    71: op1_07_inv11 = 1;
    75: op1_07_inv11 = 1;
    80: op1_07_inv11 = 1;
    81: op1_07_inv11 = 1;
    90: op1_07_inv11 = 1;
    93: op1_07_inv11 = 1;
    94: op1_07_inv11 = 1;
    96: op1_07_inv11 = 1;
    97: op1_07_inv11 = 1;
    default: op1_07_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in12 = imem04_in[127:124];
    22: op1_07_in12 = imem04_in[127:124];
    6: op1_07_in12 = reg_0357;
    7: op1_07_in12 = imem06_in[79:76];
    8: op1_07_in12 = reg_0461;
    9: op1_07_in12 = reg_0393;
    10: op1_07_in12 = imem02_in[119:116];
    37: op1_07_in12 = imem02_in[119:116];
    11: op1_07_in12 = reg_0285;
    12: op1_07_in12 = reg_0103;
    13: op1_07_in12 = imem07_in[51:48];
    14: op1_07_in12 = reg_0479;
    15: op1_07_in12 = imem02_in[47:44];
    16: op1_07_in12 = reg_0827;
    17: op1_07_in12 = reg_0375;
    18: op1_07_in12 = imem04_in[51:48];
    62: op1_07_in12 = imem04_in[51:48];
    19: op1_07_in12 = reg_0433;
    20: op1_07_in12 = reg_0748;
    21: op1_07_in12 = reg_0171;
    23: op1_07_in12 = imem04_in[99:96];
    24: op1_07_in12 = reg_0310;
    25: op1_07_in12 = reg_0948;
    26: op1_07_in12 = reg_0196;
    59: op1_07_in12 = reg_0196;
    70: op1_07_in12 = reg_0196;
    27: op1_07_in12 = reg_0960;
    28: op1_07_in12 = reg_0486;
    29: op1_07_in12 = reg_0265;
    30: op1_07_in12 = reg_0816;
    31: op1_07_in12 = reg_0712;
    32: op1_07_in12 = reg_0646;
    33: op1_07_in12 = imem03_in[111:108];
    34: op1_07_in12 = reg_0497;
    35: op1_07_in12 = reg_1039;
    36: op1_07_in12 = reg_0208;
    38: op1_07_in12 = reg_1035;
    39: op1_07_in12 = reg_1005;
    40: op1_07_in12 = reg_0140;
    41: op1_07_in12 = reg_0966;
    42: op1_07_in12 = reg_0211;
    43: op1_07_in12 = reg_0665;
    44: op1_07_in12 = reg_0799;
    45: op1_07_in12 = reg_0744;
    46: op1_07_in12 = reg_0689;
    47: op1_07_in12 = reg_0990;
    48: op1_07_in12 = imem07_in[55:52];
    49: op1_07_in12 = reg_0452;
    85: op1_07_in12 = reg_0452;
    50: op1_07_in12 = reg_0162;
    51: op1_07_in12 = reg_0391;
    52: op1_07_in12 = reg_0568;
    53: op1_07_in12 = imem06_in[11:8];
    54: op1_07_in12 = reg_0609;
    55: op1_07_in12 = reg_0168;
    57: op1_07_in12 = reg_0459;
    58: op1_07_in12 = reg_0737;
    60: op1_07_in12 = imem03_in[43:40];
    61: op1_07_in12 = reg_0648;
    63: op1_07_in12 = reg_0166;
    64: op1_07_in12 = reg_0166;
    65: op1_07_in12 = reg_0186;
    66: op1_07_in12 = reg_0480;
    91: op1_07_in12 = reg_0480;
    67: op1_07_in12 = reg_0210;
    68: op1_07_in12 = reg_0012;
    69: op1_07_in12 = imem06_in[27:24];
    71: op1_07_in12 = reg_0113;
    73: op1_07_in12 = imem01_in[51:48];
    74: op1_07_in12 = reg_0474;
    75: op1_07_in12 = reg_0359;
    76: op1_07_in12 = reg_0850;
    77: op1_07_in12 = reg_0292;
    78: op1_07_in12 = reg_0965;
    80: op1_07_in12 = reg_0205;
    81: op1_07_in12 = reg_0054;
    82: op1_07_in12 = reg_0473;
    83: op1_07_in12 = reg_1010;
    84: op1_07_in12 = reg_0551;
    86: op1_07_in12 = imem02_in[63:60];
    87: op1_07_in12 = reg_0267;
    89: op1_07_in12 = reg_0437;
    90: op1_07_in12 = reg_0202;
    92: op1_07_in12 = reg_0193;
    93: op1_07_in12 = imem04_in[107:104];
    94: op1_07_in12 = imem04_in[11:8];
    95: op1_07_in12 = reg_0385;
    96: op1_07_in12 = reg_0495;
    97: op1_07_in12 = reg_0424;
    default: op1_07_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv12 = 1;
    6: op1_07_inv12 = 1;
    7: op1_07_inv12 = 1;
    9: op1_07_inv12 = 1;
    10: op1_07_inv12 = 1;
    11: op1_07_inv12 = 1;
    13: op1_07_inv12 = 1;
    16: op1_07_inv12 = 1;
    17: op1_07_inv12 = 1;
    18: op1_07_inv12 = 1;
    19: op1_07_inv12 = 1;
    21: op1_07_inv12 = 1;
    29: op1_07_inv12 = 1;
    31: op1_07_inv12 = 1;
    33: op1_07_inv12 = 1;
    34: op1_07_inv12 = 1;
    35: op1_07_inv12 = 1;
    36: op1_07_inv12 = 1;
    38: op1_07_inv12 = 1;
    39: op1_07_inv12 = 1;
    41: op1_07_inv12 = 1;
    43: op1_07_inv12 = 1;
    48: op1_07_inv12 = 1;
    50: op1_07_inv12 = 1;
    52: op1_07_inv12 = 1;
    53: op1_07_inv12 = 1;
    54: op1_07_inv12 = 1;
    57: op1_07_inv12 = 1;
    58: op1_07_inv12 = 1;
    60: op1_07_inv12 = 1;
    61: op1_07_inv12 = 1;
    62: op1_07_inv12 = 1;
    63: op1_07_inv12 = 1;
    66: op1_07_inv12 = 1;
    69: op1_07_inv12 = 1;
    73: op1_07_inv12 = 1;
    74: op1_07_inv12 = 1;
    76: op1_07_inv12 = 1;
    77: op1_07_inv12 = 1;
    78: op1_07_inv12 = 1;
    82: op1_07_inv12 = 1;
    83: op1_07_inv12 = 1;
    89: op1_07_inv12 = 1;
    92: op1_07_inv12 = 1;
    93: op1_07_inv12 = 1;
    94: op1_07_inv12 = 1;
    95: op1_07_inv12 = 1;
    default: op1_07_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in13 = reg_0548;
    6: op1_07_in13 = reg_0358;
    7: op1_07_in13 = imem06_in[111:108];
    8: op1_07_in13 = reg_0477;
    9: op1_07_in13 = reg_0991;
    10: op1_07_in13 = reg_0642;
    37: op1_07_in13 = reg_0642;
    11: op1_07_in13 = reg_0059;
    12: op1_07_in13 = reg_0116;
    13: op1_07_in13 = imem07_in[63:60];
    14: op1_07_in13 = reg_0208;
    49: op1_07_in13 = reg_0208;
    15: op1_07_in13 = imem02_in[51:48];
    16: op1_07_in13 = reg_0908;
    17: op1_07_in13 = reg_0315;
    18: op1_07_in13 = imem04_in[59:56];
    19: op1_07_in13 = reg_0423;
    20: op1_07_in13 = reg_0047;
    22: op1_07_in13 = reg_0276;
    23: op1_07_in13 = imem04_in[119:116];
    24: op1_07_in13 = reg_0077;
    25: op1_07_in13 = reg_0964;
    26: op1_07_in13 = reg_0205;
    27: op1_07_in13 = reg_0252;
    28: op1_07_in13 = reg_0005;
    29: op1_07_in13 = reg_0277;
    30: op1_07_in13 = reg_0785;
    31: op1_07_in13 = reg_0707;
    32: op1_07_in13 = reg_0639;
    33: op1_07_in13 = imem03_in[127:124];
    34: op1_07_in13 = reg_0151;
    35: op1_07_in13 = reg_0230;
    36: op1_07_in13 = reg_0210;
    38: op1_07_in13 = reg_1041;
    39: op1_07_in13 = reg_0066;
    40: op1_07_in13 = imem06_in[51:48];
    41: op1_07_in13 = reg_0957;
    42: op1_07_in13 = reg_0201;
    43: op1_07_in13 = reg_0652;
    44: op1_07_in13 = reg_0302;
    45: op1_07_in13 = reg_0641;
    46: op1_07_in13 = reg_0670;
    47: op1_07_in13 = imem04_in[7:4];
    48: op1_07_in13 = imem07_in[59:56];
    50: op1_07_in13 = reg_0159;
    51: op1_07_in13 = reg_0388;
    52: op1_07_in13 = reg_0850;
    53: op1_07_in13 = imem06_in[23:20];
    54: op1_07_in13 = reg_1010;
    57: op1_07_in13 = reg_0214;
    58: op1_07_in13 = reg_1017;
    59: op1_07_in13 = imem01_in[47:44];
    60: op1_07_in13 = imem03_in[59:56];
    61: op1_07_in13 = reg_0837;
    62: op1_07_in13 = imem04_in[67:64];
    63: op1_07_in13 = reg_0185;
    64: op1_07_in13 = reg_0164;
    65: op1_07_in13 = reg_0213;
    66: op1_07_in13 = reg_0471;
    74: op1_07_in13 = reg_0471;
    67: op1_07_in13 = reg_0203;
    68: op1_07_in13 = reg_0357;
    69: op1_07_in13 = imem06_in[63:60];
    70: op1_07_in13 = reg_0195;
    85: op1_07_in13 = reg_0195;
    71: op1_07_in13 = imem02_in[55:52];
    73: op1_07_in13 = imem01_in[67:64];
    75: op1_07_in13 = reg_0389;
    76: op1_07_in13 = reg_0014;
    77: op1_07_in13 = reg_0540;
    78: op1_07_in13 = reg_0741;
    80: op1_07_in13 = reg_0192;
    81: op1_07_in13 = reg_0776;
    82: op1_07_in13 = reg_0187;
    83: op1_07_in13 = reg_0403;
    84: op1_07_in13 = reg_0985;
    86: op1_07_in13 = imem02_in[71:68];
    87: op1_07_in13 = reg_0393;
    89: op1_07_in13 = reg_0780;
    90: op1_07_in13 = reg_0206;
    91: op1_07_in13 = reg_0470;
    92: op1_07_in13 = reg_0198;
    93: op1_07_in13 = reg_0147;
    94: op1_07_in13 = imem04_in[19:16];
    95: op1_07_in13 = reg_0373;
    96: op1_07_in13 = reg_0777;
    97: op1_07_in13 = reg_0248;
    default: op1_07_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv13 = 1;
    6: op1_07_inv13 = 1;
    7: op1_07_inv13 = 1;
    8: op1_07_inv13 = 1;
    13: op1_07_inv13 = 1;
    14: op1_07_inv13 = 1;
    15: op1_07_inv13 = 1;
    17: op1_07_inv13 = 1;
    18: op1_07_inv13 = 1;
    20: op1_07_inv13 = 1;
    22: op1_07_inv13 = 1;
    24: op1_07_inv13 = 1;
    25: op1_07_inv13 = 1;
    27: op1_07_inv13 = 1;
    28: op1_07_inv13 = 1;
    31: op1_07_inv13 = 1;
    32: op1_07_inv13 = 1;
    34: op1_07_inv13 = 1;
    36: op1_07_inv13 = 1;
    38: op1_07_inv13 = 1;
    40: op1_07_inv13 = 1;
    41: op1_07_inv13 = 1;
    42: op1_07_inv13 = 1;
    43: op1_07_inv13 = 1;
    48: op1_07_inv13 = 1;
    49: op1_07_inv13 = 1;
    50: op1_07_inv13 = 1;
    51: op1_07_inv13 = 1;
    52: op1_07_inv13 = 1;
    59: op1_07_inv13 = 1;
    60: op1_07_inv13 = 1;
    63: op1_07_inv13 = 1;
    64: op1_07_inv13 = 1;
    65: op1_07_inv13 = 1;
    66: op1_07_inv13 = 1;
    67: op1_07_inv13 = 1;
    73: op1_07_inv13 = 1;
    76: op1_07_inv13 = 1;
    78: op1_07_inv13 = 1;
    80: op1_07_inv13 = 1;
    83: op1_07_inv13 = 1;
    84: op1_07_inv13 = 1;
    85: op1_07_inv13 = 1;
    86: op1_07_inv13 = 1;
    89: op1_07_inv13 = 1;
    90: op1_07_inv13 = 1;
    91: op1_07_inv13 = 1;
    92: op1_07_inv13 = 1;
    93: op1_07_inv13 = 1;
    97: op1_07_inv13 = 1;
    default: op1_07_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in14 = reg_0549;
    6: op1_07_in14 = reg_0318;
    7: op1_07_in14 = reg_0625;
    8: op1_07_in14 = reg_0460;
    9: op1_07_in14 = reg_0983;
    10: op1_07_in14 = reg_0637;
    11: op1_07_in14 = reg_0066;
    12: op1_07_in14 = reg_0108;
    13: op1_07_in14 = imem07_in[111:108];
    14: op1_07_in14 = reg_0196;
    42: op1_07_in14 = reg_0196;
    15: op1_07_in14 = imem02_in[67:64];
    16: op1_07_in14 = reg_0252;
    17: op1_07_in14 = reg_0367;
    18: op1_07_in14 = imem04_in[67:64];
    19: op1_07_in14 = reg_0175;
    20: op1_07_in14 = reg_0043;
    22: op1_07_in14 = reg_0732;
    23: op1_07_in14 = reg_0534;
    24: op1_07_in14 = imem03_in[7:4];
    25: op1_07_in14 = reg_0968;
    26: op1_07_in14 = imem01_in[15:12];
    27: op1_07_in14 = reg_0257;
    28: op1_07_in14 = reg_0011;
    29: op1_07_in14 = reg_0292;
    30: op1_07_in14 = reg_0832;
    31: op1_07_in14 = reg_0727;
    32: op1_07_in14 = reg_0651;
    33: op1_07_in14 = reg_0940;
    34: op1_07_in14 = reg_0142;
    35: op1_07_in14 = reg_1033;
    36: op1_07_in14 = reg_0194;
    37: op1_07_in14 = reg_0645;
    61: op1_07_in14 = reg_0645;
    38: op1_07_in14 = reg_0871;
    39: op1_07_in14 = reg_0296;
    40: op1_07_in14 = imem06_in[91:88];
    41: op1_07_in14 = reg_0948;
    43: op1_07_in14 = reg_0842;
    44: op1_07_in14 = reg_0748;
    45: op1_07_in14 = reg_0420;
    46: op1_07_in14 = reg_0687;
    47: op1_07_in14 = imem04_in[55:52];
    48: op1_07_in14 = imem07_in[79:76];
    49: op1_07_in14 = reg_0191;
    50: op1_07_in14 = reg_0185;
    51: op1_07_in14 = reg_0390;
    52: op1_07_in14 = reg_0014;
    53: op1_07_in14 = imem06_in[31:28];
    54: op1_07_in14 = reg_0531;
    57: op1_07_in14 = reg_0189;
    58: op1_07_in14 = reg_0615;
    59: op1_07_in14 = imem01_in[67:64];
    60: op1_07_in14 = imem03_in[63:60];
    62: op1_07_in14 = imem04_in[71:68];
    63: op1_07_in14 = reg_0157;
    64: op1_07_in14 = reg_0157;
    65: op1_07_in14 = imem01_in[75:72];
    66: op1_07_in14 = reg_0200;
    91: op1_07_in14 = reg_0200;
    67: op1_07_in14 = reg_0207;
    68: op1_07_in14 = reg_0445;
    69: op1_07_in14 = imem06_in[67:64];
    70: op1_07_in14 = imem01_in[23:20];
    71: op1_07_in14 = imem02_in[99:96];
    73: op1_07_in14 = imem01_in[91:88];
    74: op1_07_in14 = reg_0468;
    75: op1_07_in14 = reg_0335;
    97: op1_07_in14 = reg_0335;
    76: op1_07_in14 = reg_0809;
    77: op1_07_in14 = reg_0313;
    78: op1_07_in14 = imem06_in[43:40];
    80: op1_07_in14 = reg_0197;
    81: op1_07_in14 = reg_0876;
    82: op1_07_in14 = reg_0192;
    83: op1_07_in14 = reg_0782;
    84: op1_07_in14 = reg_0982;
    95: op1_07_in14 = reg_0982;
    85: op1_07_in14 = imem01_in[31:28];
    86: op1_07_in14 = imem02_in[107:104];
    87: op1_07_in14 = reg_0025;
    89: op1_07_in14 = reg_0949;
    90: op1_07_in14 = imem01_in[43:40];
    92: op1_07_in14 = reg_0213;
    93: op1_07_in14 = reg_0511;
    94: op1_07_in14 = imem04_in[27:24];
    96: op1_07_in14 = reg_0824;
    default: op1_07_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv14 = 1;
    7: op1_07_inv14 = 1;
    9: op1_07_inv14 = 1;
    13: op1_07_inv14 = 1;
    14: op1_07_inv14 = 1;
    15: op1_07_inv14 = 1;
    16: op1_07_inv14 = 1;
    18: op1_07_inv14 = 1;
    23: op1_07_inv14 = 1;
    24: op1_07_inv14 = 1;
    26: op1_07_inv14 = 1;
    28: op1_07_inv14 = 1;
    29: op1_07_inv14 = 1;
    31: op1_07_inv14 = 1;
    33: op1_07_inv14 = 1;
    34: op1_07_inv14 = 1;
    41: op1_07_inv14 = 1;
    42: op1_07_inv14 = 1;
    44: op1_07_inv14 = 1;
    47: op1_07_inv14 = 1;
    48: op1_07_inv14 = 1;
    52: op1_07_inv14 = 1;
    54: op1_07_inv14 = 1;
    57: op1_07_inv14 = 1;
    60: op1_07_inv14 = 1;
    62: op1_07_inv14 = 1;
    64: op1_07_inv14 = 1;
    66: op1_07_inv14 = 1;
    67: op1_07_inv14 = 1;
    68: op1_07_inv14 = 1;
    81: op1_07_inv14 = 1;
    84: op1_07_inv14 = 1;
    86: op1_07_inv14 = 1;
    87: op1_07_inv14 = 1;
    93: op1_07_inv14 = 1;
    94: op1_07_inv14 = 1;
    97: op1_07_inv14 = 1;
    default: op1_07_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in15 = reg_0546;
    6: op1_07_in15 = reg_0330;
    7: op1_07_in15 = reg_0626;
    87: op1_07_in15 = reg_0626;
    8: op1_07_in15 = reg_0472;
    9: op1_07_in15 = imem04_in[27:24];
    10: op1_07_in15 = reg_0656;
    11: op1_07_in15 = reg_0076;
    12: op1_07_in15 = reg_0114;
    13: op1_07_in15 = reg_0722;
    14: op1_07_in15 = reg_0205;
    15: op1_07_in15 = imem02_in[71:68];
    16: op1_07_in15 = reg_0865;
    17: op1_07_in15 = reg_0337;
    18: op1_07_in15 = imem04_in[71:68];
    19: op1_07_in15 = reg_0165;
    20: op1_07_in15 = reg_0057;
    22: op1_07_in15 = reg_0283;
    23: op1_07_in15 = reg_0302;
    24: op1_07_in15 = imem03_in[11:8];
    25: op1_07_in15 = reg_0946;
    26: op1_07_in15 = imem01_in[19:16];
    27: op1_07_in15 = reg_0831;
    28: op1_07_in15 = imem07_in[23:20];
    29: op1_07_in15 = reg_0050;
    30: op1_07_in15 = reg_0489;
    31: op1_07_in15 = reg_0430;
    32: op1_07_in15 = reg_0641;
    33: op1_07_in15 = reg_0492;
    34: op1_07_in15 = reg_0138;
    35: op1_07_in15 = reg_0227;
    36: op1_07_in15 = reg_0213;
    37: op1_07_in15 = reg_0664;
    38: op1_07_in15 = reg_0111;
    39: op1_07_in15 = reg_0882;
    40: op1_07_in15 = imem06_in[123:120];
    41: op1_07_in15 = reg_0968;
    42: op1_07_in15 = reg_0212;
    43: op1_07_in15 = reg_0290;
    44: op1_07_in15 = reg_0043;
    45: op1_07_in15 = reg_0024;
    46: op1_07_in15 = reg_0475;
    47: op1_07_in15 = imem04_in[59:56];
    48: op1_07_in15 = imem07_in[83:80];
    49: op1_07_in15 = reg_0210;
    50: op1_07_in15 = reg_0176;
    64: op1_07_in15 = reg_0176;
    51: op1_07_in15 = reg_0349;
    52: op1_07_in15 = reg_0074;
    53: op1_07_in15 = imem06_in[47:44];
    54: op1_07_in15 = reg_0008;
    57: op1_07_in15 = reg_0190;
    92: op1_07_in15 = reg_0190;
    58: op1_07_in15 = reg_0232;
    59: op1_07_in15 = imem01_in[75:72];
    60: op1_07_in15 = imem03_in[75:72];
    61: op1_07_in15 = reg_0039;
    62: op1_07_in15 = imem04_in[95:92];
    65: op1_07_in15 = imem01_in[87:84];
    66: op1_07_in15 = reg_0208;
    67: op1_07_in15 = imem01_in[27:24];
    70: op1_07_in15 = imem01_in[27:24];
    68: op1_07_in15 = reg_0322;
    69: op1_07_in15 = imem06_in[71:68];
    78: op1_07_in15 = imem06_in[71:68];
    71: op1_07_in15 = imem02_in[119:116];
    73: op1_07_in15 = imem01_in[115:112];
    74: op1_07_in15 = reg_0452;
    75: op1_07_in15 = reg_0776;
    76: op1_07_in15 = reg_0288;
    77: op1_07_in15 = reg_0850;
    80: op1_07_in15 = imem01_in[55:52];
    81: op1_07_in15 = imem03_in[7:4];
    82: op1_07_in15 = reg_0197;
    83: op1_07_in15 = reg_0369;
    84: op1_07_in15 = reg_0984;
    85: op1_07_in15 = imem01_in[67:64];
    86: op1_07_in15 = reg_0605;
    89: op1_07_in15 = reg_0851;
    90: op1_07_in15 = imem01_in[91:88];
    91: op1_07_in15 = reg_0204;
    93: op1_07_in15 = reg_0390;
    94: op1_07_in15 = imem04_in[31:28];
    95: op1_07_in15 = reg_0242;
    96: op1_07_in15 = reg_0542;
    97: op1_07_in15 = reg_0516;
    default: op1_07_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv15 = 1;
    8: op1_07_inv15 = 1;
    11: op1_07_inv15 = 1;
    12: op1_07_inv15 = 1;
    16: op1_07_inv15 = 1;
    18: op1_07_inv15 = 1;
    24: op1_07_inv15 = 1;
    26: op1_07_inv15 = 1;
    27: op1_07_inv15 = 1;
    30: op1_07_inv15 = 1;
    33: op1_07_inv15 = 1;
    37: op1_07_inv15 = 1;
    38: op1_07_inv15 = 1;
    43: op1_07_inv15 = 1;
    45: op1_07_inv15 = 1;
    46: op1_07_inv15 = 1;
    48: op1_07_inv15 = 1;
    49: op1_07_inv15 = 1;
    50: op1_07_inv15 = 1;
    51: op1_07_inv15 = 1;
    54: op1_07_inv15 = 1;
    57: op1_07_inv15 = 1;
    59: op1_07_inv15 = 1;
    64: op1_07_inv15 = 1;
    65: op1_07_inv15 = 1;
    66: op1_07_inv15 = 1;
    67: op1_07_inv15 = 1;
    69: op1_07_inv15 = 1;
    70: op1_07_inv15 = 1;
    71: op1_07_inv15 = 1;
    73: op1_07_inv15 = 1;
    74: op1_07_inv15 = 1;
    80: op1_07_inv15 = 1;
    83: op1_07_inv15 = 1;
    89: op1_07_inv15 = 1;
    90: op1_07_inv15 = 1;
    91: op1_07_inv15 = 1;
    94: op1_07_inv15 = 1;
    95: op1_07_inv15 = 1;
    97: op1_07_inv15 = 1;
    default: op1_07_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in16 = reg_0301;
    6: op1_07_in16 = reg_0310;
    7: op1_07_in16 = reg_0633;
    8: op1_07_in16 = reg_0208;
    9: op1_07_in16 = imem04_in[31:28];
    10: op1_07_in16 = reg_0641;
    11: op1_07_in16 = reg_0048;
    12: op1_07_in16 = reg_0101;
    13: op1_07_in16 = reg_0723;
    14: op1_07_in16 = reg_0195;
    57: op1_07_in16 = reg_0195;
    15: op1_07_in16 = imem02_in[79:76];
    16: op1_07_in16 = reg_0832;
    17: op1_07_in16 = reg_0780;
    18: op1_07_in16 = imem05_in[23:20];
    19: op1_07_in16 = reg_0181;
    20: op1_07_in16 = reg_0286;
    22: op1_07_in16 = reg_0736;
    23: op1_07_in16 = reg_0829;
    24: op1_07_in16 = imem03_in[19:16];
    25: op1_07_in16 = reg_0961;
    26: op1_07_in16 = imem01_in[31:28];
    27: op1_07_in16 = reg_0132;
    28: op1_07_in16 = imem07_in[47:44];
    29: op1_07_in16 = reg_0313;
    30: op1_07_in16 = reg_0145;
    31: op1_07_in16 = reg_0426;
    32: op1_07_in16 = reg_0318;
    33: op1_07_in16 = reg_0317;
    34: op1_07_in16 = reg_0130;
    35: op1_07_in16 = reg_1017;
    36: op1_07_in16 = imem01_in[39:36];
    82: op1_07_in16 = imem01_in[39:36];
    37: op1_07_in16 = reg_0661;
    38: op1_07_in16 = reg_0125;
    39: op1_07_in16 = reg_0009;
    40: op1_07_in16 = reg_0614;
    41: op1_07_in16 = reg_0960;
    42: op1_07_in16 = reg_0197;
    43: op1_07_in16 = reg_0225;
    44: op1_07_in16 = imem05_in[3:0];
    96: op1_07_in16 = imem05_in[3:0];
    45: op1_07_in16 = reg_0175;
    46: op1_07_in16 = reg_0460;
    47: op1_07_in16 = imem04_in[71:68];
    48: op1_07_in16 = reg_0730;
    49: op1_07_in16 = reg_0204;
    66: op1_07_in16 = reg_0204;
    51: op1_07_in16 = reg_0222;
    52: op1_07_in16 = reg_0288;
    53: op1_07_in16 = imem06_in[63:60];
    54: op1_07_in16 = reg_0029;
    58: op1_07_in16 = reg_1055;
    59: op1_07_in16 = reg_0218;
    60: op1_07_in16 = imem03_in[83:80];
    61: op1_07_in16 = reg_0052;
    62: op1_07_in16 = imem04_in[123:120];
    65: op1_07_in16 = imem01_in[95:92];
    67: op1_07_in16 = imem01_in[51:48];
    68: op1_07_in16 = reg_0346;
    69: op1_07_in16 = imem06_in[111:108];
    70: op1_07_in16 = imem01_in[35:32];
    71: op1_07_in16 = reg_0905;
    73: op1_07_in16 = imem01_in[119:116];
    74: op1_07_in16 = reg_0456;
    75: op1_07_in16 = reg_0084;
    76: op1_07_in16 = reg_0407;
    77: op1_07_in16 = reg_0014;
    78: op1_07_in16 = imem06_in[79:76];
    80: op1_07_in16 = imem01_in[99:96];
    81: op1_07_in16 = imem03_in[11:8];
    83: op1_07_in16 = imem07_in[31:28];
    84: op1_07_in16 = reg_0988;
    85: op1_07_in16 = imem01_in[79:76];
    86: op1_07_in16 = reg_0305;
    87: op1_07_in16 = reg_1011;
    89: op1_07_in16 = reg_0688;
    90: op1_07_in16 = reg_0969;
    91: op1_07_in16 = reg_0193;
    92: op1_07_in16 = reg_0199;
    93: op1_07_in16 = reg_0008;
    94: op1_07_in16 = imem04_in[39:36];
    95: op1_07_in16 = reg_0986;
    97: op1_07_in16 = reg_0772;
    default: op1_07_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_07_inv16 = 1;
    8: op1_07_inv16 = 1;
    10: op1_07_inv16 = 1;
    12: op1_07_inv16 = 1;
    14: op1_07_inv16 = 1;
    15: op1_07_inv16 = 1;
    18: op1_07_inv16 = 1;
    19: op1_07_inv16 = 1;
    23: op1_07_inv16 = 1;
    24: op1_07_inv16 = 1;
    25: op1_07_inv16 = 1;
    28: op1_07_inv16 = 1;
    29: op1_07_inv16 = 1;
    30: op1_07_inv16 = 1;
    31: op1_07_inv16 = 1;
    32: op1_07_inv16 = 1;
    35: op1_07_inv16 = 1;
    36: op1_07_inv16 = 1;
    37: op1_07_inv16 = 1;
    47: op1_07_inv16 = 1;
    49: op1_07_inv16 = 1;
    51: op1_07_inv16 = 1;
    52: op1_07_inv16 = 1;
    58: op1_07_inv16 = 1;
    62: op1_07_inv16 = 1;
    68: op1_07_inv16 = 1;
    69: op1_07_inv16 = 1;
    70: op1_07_inv16 = 1;
    71: op1_07_inv16 = 1;
    76: op1_07_inv16 = 1;
    78: op1_07_inv16 = 1;
    80: op1_07_inv16 = 1;
    81: op1_07_inv16 = 1;
    85: op1_07_inv16 = 1;
    87: op1_07_inv16 = 1;
    89: op1_07_inv16 = 1;
    91: op1_07_inv16 = 1;
    default: op1_07_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in17 = reg_0289;
    6: op1_07_in17 = reg_0336;
    7: op1_07_in17 = reg_0615;
    8: op1_07_in17 = reg_0210;
    9: op1_07_in17 = imem04_in[95:92];
    10: op1_07_in17 = reg_0662;
    11: op1_07_in17 = reg_0063;
    12: op1_07_in17 = reg_0126;
    13: op1_07_in17 = reg_0703;
    14: op1_07_in17 = imem01_in[27:24];
    15: op1_07_in17 = imem02_in[91:88];
    16: op1_07_in17 = reg_0894;
    17: op1_07_in17 = reg_0801;
    18: op1_07_in17 = imem05_in[63:60];
    19: op1_07_in17 = reg_0161;
    20: op1_07_in17 = reg_0270;
    22: op1_07_in17 = reg_0279;
    23: op1_07_in17 = reg_0824;
    24: op1_07_in17 = imem03_in[47:44];
    25: op1_07_in17 = reg_0215;
    41: op1_07_in17 = reg_0215;
    26: op1_07_in17 = imem01_in[47:44];
    27: op1_07_in17 = reg_0135;
    28: op1_07_in17 = imem07_in[111:108];
    29: op1_07_in17 = reg_0740;
    30: op1_07_in17 = reg_0151;
    31: op1_07_in17 = reg_0445;
    32: op1_07_in17 = reg_0339;
    33: op1_07_in17 = reg_0938;
    34: op1_07_in17 = reg_0140;
    35: op1_07_in17 = reg_0104;
    36: op1_07_in17 = imem01_in[79:76];
    37: op1_07_in17 = reg_0644;
    38: op1_07_in17 = reg_0112;
    39: op1_07_in17 = reg_0283;
    40: op1_07_in17 = reg_0895;
    42: op1_07_in17 = imem01_in[3:0];
    43: op1_07_in17 = reg_0817;
    44: op1_07_in17 = imem05_in[7:4];
    96: op1_07_in17 = imem05_in[7:4];
    45: op1_07_in17 = reg_0163;
    46: op1_07_in17 = reg_0473;
    47: op1_07_in17 = imem04_in[91:88];
    48: op1_07_in17 = reg_0731;
    49: op1_07_in17 = reg_0188;
    51: op1_07_in17 = reg_1029;
    52: op1_07_in17 = reg_0061;
    53: op1_07_in17 = imem06_in[115:112];
    54: op1_07_in17 = imem07_in[23:20];
    57: op1_07_in17 = imem01_in[11:8];
    58: op1_07_in17 = reg_0273;
    59: op1_07_in17 = reg_0242;
    65: op1_07_in17 = reg_0242;
    60: op1_07_in17 = imem03_in[95:92];
    61: op1_07_in17 = reg_0394;
    62: op1_07_in17 = reg_0277;
    66: op1_07_in17 = reg_0193;
    67: op1_07_in17 = imem01_in[59:56];
    68: op1_07_in17 = reg_0823;
    69: op1_07_in17 = imem06_in[127:124];
    70: op1_07_in17 = imem01_in[55:52];
    71: op1_07_in17 = reg_0654;
    73: op1_07_in17 = reg_1032;
    74: op1_07_in17 = reg_0208;
    75: op1_07_in17 = reg_0310;
    76: op1_07_in17 = reg_0627;
    77: op1_07_in17 = reg_0854;
    78: op1_07_in17 = imem06_in[107:104];
    80: op1_07_in17 = imem01_in[103:100];
    81: op1_07_in17 = imem03_in[27:24];
    82: op1_07_in17 = imem01_in[43:40];
    83: op1_07_in17 = imem07_in[67:64];
    84: op1_07_in17 = imem04_in[43:40];
    85: op1_07_in17 = imem01_in[99:96];
    86: op1_07_in17 = reg_0090;
    87: op1_07_in17 = reg_0926;
    89: op1_07_in17 = reg_0705;
    90: op1_07_in17 = reg_0122;
    91: op1_07_in17 = reg_0211;
    92: op1_07_in17 = imem01_in[67:64];
    93: op1_07_in17 = reg_0882;
    94: op1_07_in17 = imem04_in[67:64];
    95: op1_07_in17 = reg_0989;
    97: op1_07_in17 = reg_0086;
    default: op1_07_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_07_inv17 = 1;
    7: op1_07_inv17 = 1;
    8: op1_07_inv17 = 1;
    12: op1_07_inv17 = 1;
    13: op1_07_inv17 = 1;
    14: op1_07_inv17 = 1;
    15: op1_07_inv17 = 1;
    17: op1_07_inv17 = 1;
    19: op1_07_inv17 = 1;
    22: op1_07_inv17 = 1;
    25: op1_07_inv17 = 1;
    26: op1_07_inv17 = 1;
    34: op1_07_inv17 = 1;
    36: op1_07_inv17 = 1;
    37: op1_07_inv17 = 1;
    38: op1_07_inv17 = 1;
    39: op1_07_inv17 = 1;
    43: op1_07_inv17 = 1;
    44: op1_07_inv17 = 1;
    45: op1_07_inv17 = 1;
    46: op1_07_inv17 = 1;
    48: op1_07_inv17 = 1;
    49: op1_07_inv17 = 1;
    54: op1_07_inv17 = 1;
    59: op1_07_inv17 = 1;
    61: op1_07_inv17 = 1;
    66: op1_07_inv17 = 1;
    68: op1_07_inv17 = 1;
    75: op1_07_inv17 = 1;
    77: op1_07_inv17 = 1;
    80: op1_07_inv17 = 1;
    82: op1_07_inv17 = 1;
    84: op1_07_inv17 = 1;
    85: op1_07_inv17 = 1;
    87: op1_07_inv17 = 1;
    90: op1_07_inv17 = 1;
    91: op1_07_inv17 = 1;
    94: op1_07_inv17 = 1;
    96: op1_07_inv17 = 1;
    default: op1_07_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in18 = reg_0290;
    6: op1_07_in18 = reg_0083;
    7: op1_07_in18 = reg_0348;
    8: op1_07_in18 = reg_0203;
    9: op1_07_in18 = imem04_in[107:104];
    10: op1_07_in18 = reg_0358;
    11: op1_07_in18 = reg_0075;
    12: op1_07_in18 = imem02_in[63:60];
    13: op1_07_in18 = reg_0705;
    14: op1_07_in18 = imem01_in[35:32];
    15: op1_07_in18 = reg_0657;
    16: op1_07_in18 = reg_0134;
    17: op1_07_in18 = reg_0017;
    18: op1_07_in18 = imem05_in[111:108];
    19: op1_07_in18 = reg_0167;
    20: op1_07_in18 = reg_0509;
    22: op1_07_in18 = reg_0058;
    23: op1_07_in18 = reg_0060;
    24: op1_07_in18 = reg_0596;
    25: op1_07_in18 = reg_0821;
    26: op1_07_in18 = imem01_in[91:88];
    27: op1_07_in18 = reg_0136;
    28: op1_07_in18 = imem07_in[127:124];
    29: op1_07_in18 = reg_0763;
    30: op1_07_in18 = reg_0155;
    31: op1_07_in18 = reg_0160;
    32: op1_07_in18 = reg_0098;
    33: op1_07_in18 = reg_1007;
    34: op1_07_in18 = imem06_in[39:36];
    35: op1_07_in18 = reg_0119;
    36: op1_07_in18 = imem01_in[83:80];
    37: op1_07_in18 = reg_0659;
    38: op1_07_in18 = reg_0100;
    39: op1_07_in18 = reg_0043;
    40: op1_07_in18 = reg_0624;
    41: op1_07_in18 = reg_0900;
    42: op1_07_in18 = imem01_in[15:12];
    43: op1_07_in18 = reg_0516;
    44: op1_07_in18 = imem05_in[27:24];
    45: op1_07_in18 = reg_0184;
    46: op1_07_in18 = reg_0458;
    47: op1_07_in18 = imem04_in[127:124];
    48: op1_07_in18 = reg_0714;
    49: op1_07_in18 = reg_0196;
    66: op1_07_in18 = reg_0196;
    51: op1_07_in18 = reg_0628;
    52: op1_07_in18 = reg_0834;
    53: op1_07_in18 = imem06_in[123:120];
    54: op1_07_in18 = imem07_in[39:36];
    57: op1_07_in18 = imem01_in[43:40];
    58: op1_07_in18 = reg_0112;
    59: op1_07_in18 = reg_0285;
    60: op1_07_in18 = reg_0572;
    61: op1_07_in18 = reg_0389;
    62: op1_07_in18 = reg_0539;
    65: op1_07_in18 = reg_0933;
    67: op1_07_in18 = imem01_in[111:108];
    85: op1_07_in18 = imem01_in[111:108];
    68: op1_07_in18 = reg_0874;
    69: op1_07_in18 = reg_0694;
    70: op1_07_in18 = imem01_in[95:92];
    71: op1_07_in18 = reg_0855;
    73: op1_07_in18 = reg_1014;
    74: op1_07_in18 = reg_0211;
    75: op1_07_in18 = reg_0077;
    76: op1_07_in18 = reg_0854;
    77: op1_07_in18 = reg_0108;
    78: op1_07_in18 = imem06_in[111:108];
    80: op1_07_in18 = imem01_in[107:104];
    81: op1_07_in18 = imem03_in[39:36];
    82: op1_07_in18 = imem01_in[115:112];
    83: op1_07_in18 = imem07_in[71:68];
    84: op1_07_in18 = imem04_in[59:56];
    86: op1_07_in18 = reg_0639;
    87: op1_07_in18 = reg_0889;
    89: op1_07_in18 = reg_0955;
    90: op1_07_in18 = reg_0973;
    91: op1_07_in18 = reg_0213;
    92: op1_07_in18 = reg_0122;
    93: op1_07_in18 = reg_0537;
    94: op1_07_in18 = imem04_in[87:84];
    95: op1_07_in18 = reg_0547;
    96: op1_07_in18 = imem05_in[55:52];
    97: op1_07_in18 = reg_0218;
    default: op1_07_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_07_inv18 = 1;
    8: op1_07_inv18 = 1;
    10: op1_07_inv18 = 1;
    11: op1_07_inv18 = 1;
    13: op1_07_inv18 = 1;
    17: op1_07_inv18 = 1;
    18: op1_07_inv18 = 1;
    22: op1_07_inv18 = 1;
    24: op1_07_inv18 = 1;
    25: op1_07_inv18 = 1;
    27: op1_07_inv18 = 1;
    33: op1_07_inv18 = 1;
    35: op1_07_inv18 = 1;
    38: op1_07_inv18 = 1;
    40: op1_07_inv18 = 1;
    42: op1_07_inv18 = 1;
    43: op1_07_inv18 = 1;
    44: op1_07_inv18 = 1;
    45: op1_07_inv18 = 1;
    46: op1_07_inv18 = 1;
    47: op1_07_inv18 = 1;
    49: op1_07_inv18 = 1;
    52: op1_07_inv18 = 1;
    53: op1_07_inv18 = 1;
    58: op1_07_inv18 = 1;
    59: op1_07_inv18 = 1;
    61: op1_07_inv18 = 1;
    62: op1_07_inv18 = 1;
    65: op1_07_inv18 = 1;
    66: op1_07_inv18 = 1;
    68: op1_07_inv18 = 1;
    69: op1_07_inv18 = 1;
    75: op1_07_inv18 = 1;
    77: op1_07_inv18 = 1;
    78: op1_07_inv18 = 1;
    81: op1_07_inv18 = 1;
    83: op1_07_inv18 = 1;
    85: op1_07_inv18 = 1;
    87: op1_07_inv18 = 1;
    89: op1_07_inv18 = 1;
    91: op1_07_inv18 = 1;
    93: op1_07_inv18 = 1;
    94: op1_07_inv18 = 1;
    97: op1_07_inv18 = 1;
    default: op1_07_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in19 = reg_0291;
    6: op1_07_in19 = reg_0092;
    7: op1_07_in19 = reg_0372;
    8: op1_07_in19 = reg_0207;
    9: op1_07_in19 = reg_0552;
    10: op1_07_in19 = reg_0359;
    11: op1_07_in19 = imem05_in[39:36];
    12: op1_07_in19 = imem02_in[75:72];
    13: op1_07_in19 = reg_0424;
    14: op1_07_in19 = imem01_in[47:44];
    15: op1_07_in19 = reg_0639;
    16: op1_07_in19 = imem06_in[15:12];
    17: op1_07_in19 = reg_0018;
    18: op1_07_in19 = imem05_in[115:112];
    19: op1_07_in19 = reg_0159;
    20: op1_07_in19 = reg_0529;
    22: op1_07_in19 = reg_0875;
    23: op1_07_in19 = reg_0779;
    24: op1_07_in19 = reg_0583;
    25: op1_07_in19 = reg_0757;
    26: op1_07_in19 = imem01_in[95:92];
    36: op1_07_in19 = imem01_in[95:92];
    27: op1_07_in19 = reg_0133;
    28: op1_07_in19 = reg_0724;
    29: op1_07_in19 = reg_0760;
    30: op1_07_in19 = imem06_in[35:32];
    31: op1_07_in19 = reg_0183;
    32: op1_07_in19 = reg_0818;
    33: op1_07_in19 = reg_1019;
    78: op1_07_in19 = reg_1019;
    34: op1_07_in19 = imem06_in[43:40];
    35: op1_07_in19 = reg_0102;
    37: op1_07_in19 = reg_0663;
    38: op1_07_in19 = reg_0106;
    39: op1_07_in19 = reg_0044;
    40: op1_07_in19 = reg_0486;
    41: op1_07_in19 = reg_1046;
    42: op1_07_in19 = imem01_in[43:40];
    43: op1_07_in19 = reg_0772;
    44: op1_07_in19 = imem05_in[31:28];
    46: op1_07_in19 = reg_0187;
    47: op1_07_in19 = reg_0511;
    48: op1_07_in19 = reg_0713;
    49: op1_07_in19 = reg_0205;
    66: op1_07_in19 = reg_0205;
    51: op1_07_in19 = reg_0609;
    52: op1_07_in19 = reg_0031;
    53: op1_07_in19 = reg_0614;
    54: op1_07_in19 = imem07_in[59:56];
    57: op1_07_in19 = imem01_in[63:60];
    58: op1_07_in19 = reg_0733;
    59: op1_07_in19 = reg_0249;
    60: op1_07_in19 = reg_0346;
    61: op1_07_in19 = reg_0087;
    62: op1_07_in19 = reg_0055;
    65: op1_07_in19 = reg_0870;
    67: op1_07_in19 = reg_1056;
    68: op1_07_in19 = reg_0795;
    69: op1_07_in19 = reg_0344;
    70: op1_07_in19 = reg_0968;
    85: op1_07_in19 = reg_0968;
    71: op1_07_in19 = reg_0441;
    73: op1_07_in19 = reg_1023;
    82: op1_07_in19 = reg_1023;
    74: op1_07_in19 = reg_0212;
    75: op1_07_in19 = imem03_in[115:112];
    76: op1_07_in19 = imem05_in[15:12];
    77: op1_07_in19 = reg_0542;
    80: op1_07_in19 = reg_1044;
    81: op1_07_in19 = imem03_in[87:84];
    83: op1_07_in19 = reg_0567;
    84: op1_07_in19 = imem04_in[71:68];
    86: op1_07_in19 = reg_0331;
    87: op1_07_in19 = reg_0440;
    89: op1_07_in19 = reg_0093;
    90: op1_07_in19 = reg_0337;
    91: op1_07_in19 = reg_0199;
    92: op1_07_in19 = reg_1042;
    93: op1_07_in19 = reg_0067;
    94: op1_07_in19 = imem04_in[119:116];
    95: op1_07_in19 = imem04_in[47:44];
    96: op1_07_in19 = reg_0275;
    97: op1_07_in19 = reg_0082;
    default: op1_07_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_07_inv19 = 1;
    9: op1_07_inv19 = 1;
    10: op1_07_inv19 = 1;
    13: op1_07_inv19 = 1;
    15: op1_07_inv19 = 1;
    16: op1_07_inv19 = 1;
    17: op1_07_inv19 = 1;
    18: op1_07_inv19 = 1;
    22: op1_07_inv19 = 1;
    24: op1_07_inv19 = 1;
    25: op1_07_inv19 = 1;
    26: op1_07_inv19 = 1;
    27: op1_07_inv19 = 1;
    28: op1_07_inv19 = 1;
    29: op1_07_inv19 = 1;
    31: op1_07_inv19 = 1;
    35: op1_07_inv19 = 1;
    36: op1_07_inv19 = 1;
    38: op1_07_inv19 = 1;
    39: op1_07_inv19 = 1;
    40: op1_07_inv19 = 1;
    44: op1_07_inv19 = 1;
    48: op1_07_inv19 = 1;
    51: op1_07_inv19 = 1;
    52: op1_07_inv19 = 1;
    53: op1_07_inv19 = 1;
    54: op1_07_inv19 = 1;
    57: op1_07_inv19 = 1;
    59: op1_07_inv19 = 1;
    60: op1_07_inv19 = 1;
    61: op1_07_inv19 = 1;
    65: op1_07_inv19 = 1;
    69: op1_07_inv19 = 1;
    71: op1_07_inv19 = 1;
    73: op1_07_inv19 = 1;
    75: op1_07_inv19 = 1;
    76: op1_07_inv19 = 1;
    77: op1_07_inv19 = 1;
    83: op1_07_inv19 = 1;
    84: op1_07_inv19 = 1;
    85: op1_07_inv19 = 1;
    87: op1_07_inv19 = 1;
    91: op1_07_inv19 = 1;
    92: op1_07_inv19 = 1;
    93: op1_07_inv19 = 1;
    94: op1_07_inv19 = 1;
    default: op1_07_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in20 = reg_0292;
    6: op1_07_in20 = reg_0089;
    7: op1_07_in20 = reg_0349;
    8: op1_07_in20 = reg_0198;
    9: op1_07_in20 = reg_0542;
    10: op1_07_in20 = reg_0330;
    11: op1_07_in20 = imem05_in[51:48];
    12: op1_07_in20 = imem02_in[87:84];
    13: op1_07_in20 = reg_0432;
    14: op1_07_in20 = imem01_in[87:84];
    15: op1_07_in20 = reg_0638;
    16: op1_07_in20 = imem06_in[35:32];
    17: op1_07_in20 = reg_0803;
    18: op1_07_in20 = reg_0963;
    19: op1_07_in20 = reg_0160;
    20: op1_07_in20 = reg_0272;
    22: op1_07_in20 = imem05_in[43:40];
    23: op1_07_in20 = reg_0533;
    24: op1_07_in20 = reg_0387;
    25: op1_07_in20 = reg_0275;
    26: op1_07_in20 = reg_0779;
    27: op1_07_in20 = reg_0151;
    28: op1_07_in20 = reg_0709;
    29: op1_07_in20 = reg_0014;
    30: op1_07_in20 = imem06_in[39:36];
    31: op1_07_in20 = reg_0178;
    32: op1_07_in20 = reg_0007;
    33: op1_07_in20 = reg_0327;
    34: op1_07_in20 = reg_0616;
    35: op1_07_in20 = reg_0127;
    36: op1_07_in20 = imem01_in[99:96];
    37: op1_07_in20 = reg_0039;
    71: op1_07_in20 = reg_0039;
    38: op1_07_in20 = reg_0109;
    39: op1_07_in20 = reg_0021;
    40: op1_07_in20 = reg_0407;
    41: op1_07_in20 = reg_0136;
    42: op1_07_in20 = imem01_in[51:48];
    43: op1_07_in20 = reg_0758;
    44: op1_07_in20 = imem05_in[83:80];
    46: op1_07_in20 = reg_0194;
    47: op1_07_in20 = reg_1057;
    48: op1_07_in20 = reg_0002;
    49: op1_07_in20 = reg_0190;
    51: op1_07_in20 = reg_1010;
    52: op1_07_in20 = imem05_in[15:12];
    53: op1_07_in20 = reg_0883;
    54: op1_07_in20 = imem07_in[67:64];
    57: op1_07_in20 = imem01_in[107:104];
    58: op1_07_in20 = reg_0860;
    59: op1_07_in20 = reg_1034;
    60: op1_07_in20 = reg_0040;
    68: op1_07_in20 = reg_0040;
    61: op1_07_in20 = reg_0608;
    62: op1_07_in20 = reg_0313;
    65: op1_07_in20 = reg_0919;
    66: op1_07_in20 = reg_0199;
    67: op1_07_in20 = reg_1045;
    69: op1_07_in20 = reg_0244;
    70: op1_07_in20 = reg_0546;
    73: op1_07_in20 = reg_0522;
    74: op1_07_in20 = imem01_in[3:0];
    75: op1_07_in20 = imem03_in[123:120];
    76: op1_07_in20 = imem05_in[39:36];
    77: op1_07_in20 = reg_0856;
    78: op1_07_in20 = reg_0691;
    80: op1_07_in20 = reg_1056;
    85: op1_07_in20 = reg_1056;
    81: op1_07_in20 = imem03_in[95:92];
    82: op1_07_in20 = reg_1039;
    83: op1_07_in20 = reg_0721;
    84: op1_07_in20 = imem04_in[87:84];
    86: op1_07_in20 = reg_0355;
    87: op1_07_in20 = reg_0895;
    89: op1_07_in20 = reg_0725;
    90: op1_07_in20 = reg_0120;
    91: op1_07_in20 = reg_0192;
    92: op1_07_in20 = reg_0973;
    93: op1_07_in20 = reg_0302;
    94: op1_07_in20 = imem04_in[123:120];
    95: op1_07_in20 = imem04_in[63:60];
    96: op1_07_in20 = reg_0226;
    97: op1_07_in20 = imem03_in[59:56];
    default: op1_07_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv20 = 1;
    7: op1_07_inv20 = 1;
    8: op1_07_inv20 = 1;
    9: op1_07_inv20 = 1;
    11: op1_07_inv20 = 1;
    12: op1_07_inv20 = 1;
    16: op1_07_inv20 = 1;
    20: op1_07_inv20 = 1;
    22: op1_07_inv20 = 1;
    24: op1_07_inv20 = 1;
    30: op1_07_inv20 = 1;
    31: op1_07_inv20 = 1;
    32: op1_07_inv20 = 1;
    33: op1_07_inv20 = 1;
    35: op1_07_inv20 = 1;
    36: op1_07_inv20 = 1;
    37: op1_07_inv20 = 1;
    38: op1_07_inv20 = 1;
    41: op1_07_inv20 = 1;
    44: op1_07_inv20 = 1;
    46: op1_07_inv20 = 1;
    47: op1_07_inv20 = 1;
    48: op1_07_inv20 = 1;
    52: op1_07_inv20 = 1;
    54: op1_07_inv20 = 1;
    57: op1_07_inv20 = 1;
    59: op1_07_inv20 = 1;
    60: op1_07_inv20 = 1;
    65: op1_07_inv20 = 1;
    67: op1_07_inv20 = 1;
    69: op1_07_inv20 = 1;
    70: op1_07_inv20 = 1;
    71: op1_07_inv20 = 1;
    74: op1_07_inv20 = 1;
    80: op1_07_inv20 = 1;
    83: op1_07_inv20 = 1;
    85: op1_07_inv20 = 1;
    90: op1_07_inv20 = 1;
    93: op1_07_inv20 = 1;
    94: op1_07_inv20 = 1;
    default: op1_07_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in21 = reg_0288;
    6: op1_07_in21 = reg_0049;
    7: op1_07_in21 = reg_0404;
    8: op1_07_in21 = reg_0201;
    9: op1_07_in21 = reg_0555;
    10: op1_07_in21 = reg_0339;
    11: op1_07_in21 = imem05_in[63:60];
    12: op1_07_in21 = imem02_in[99:96];
    13: op1_07_in21 = reg_0422;
    14: op1_07_in21 = imem01_in[103:100];
    15: op1_07_in21 = reg_0644;
    16: op1_07_in21 = imem06_in[55:52];
    17: op1_07_in21 = reg_0011;
    18: op1_07_in21 = reg_0970;
    19: op1_07_in21 = reg_0183;
    20: op1_07_in21 = reg_0269;
    22: op1_07_in21 = imem05_in[55:52];
    76: op1_07_in21 = imem05_in[55:52];
    23: op1_07_in21 = reg_0740;
    24: op1_07_in21 = reg_1001;
    25: op1_07_in21 = reg_0896;
    26: op1_07_in21 = reg_0223;
    27: op1_07_in21 = imem06_in[7:4];
    41: op1_07_in21 = imem06_in[7:4];
    28: op1_07_in21 = reg_0715;
    29: op1_07_in21 = reg_0063;
    30: op1_07_in21 = imem06_in[59:56];
    31: op1_07_in21 = reg_0157;
    32: op1_07_in21 = reg_0482;
    61: op1_07_in21 = reg_0482;
    33: op1_07_in21 = reg_0398;
    34: op1_07_in21 = reg_0631;
    35: op1_07_in21 = reg_0126;
    36: op1_07_in21 = imem01_in[107:104];
    37: op1_07_in21 = reg_0817;
    38: op1_07_in21 = reg_0107;
    39: op1_07_in21 = imem05_in[3:0];
    40: op1_07_in21 = reg_0856;
    42: op1_07_in21 = imem01_in[75:72];
    43: op1_07_in21 = reg_0867;
    44: op1_07_in21 = imem05_in[103:100];
    46: op1_07_in21 = reg_0192;
    47: op1_07_in21 = reg_1020;
    48: op1_07_in21 = reg_0421;
    49: op1_07_in21 = reg_0206;
    51: op1_07_in21 = reg_0029;
    52: op1_07_in21 = imem05_in[23:20];
    53: op1_07_in21 = reg_0624;
    54: op1_07_in21 = imem07_in[103:100];
    57: op1_07_in21 = imem01_in[115:112];
    58: op1_07_in21 = reg_0103;
    59: op1_07_in21 = reg_0607;
    60: op1_07_in21 = reg_0784;
    62: op1_07_in21 = reg_0799;
    65: op1_07_in21 = reg_1056;
    66: op1_07_in21 = imem01_in[39:36];
    91: op1_07_in21 = imem01_in[39:36];
    67: op1_07_in21 = reg_0487;
    68: op1_07_in21 = reg_0767;
    69: op1_07_in21 = reg_0025;
    70: op1_07_in21 = reg_1023;
    90: op1_07_in21 = reg_1023;
    71: op1_07_in21 = reg_0394;
    73: op1_07_in21 = reg_0906;
    74: op1_07_in21 = imem01_in[7:4];
    75: op1_07_in21 = reg_0006;
    77: op1_07_in21 = reg_0531;
    78: op1_07_in21 = reg_0262;
    80: op1_07_in21 = reg_0503;
    81: op1_07_in21 = reg_0099;
    82: op1_07_in21 = reg_0869;
    83: op1_07_in21 = reg_0159;
    84: op1_07_in21 = reg_0147;
    85: op1_07_in21 = reg_0592;
    86: op1_07_in21 = reg_0700;
    87: op1_07_in21 = reg_1028;
    89: op1_07_in21 = reg_0625;
    92: op1_07_in21 = reg_0793;
    93: op1_07_in21 = reg_0401;
    94: op1_07_in21 = imem04_in[127:124];
    95: op1_07_in21 = imem04_in[79:76];
    96: op1_07_in21 = reg_0583;
    97: op1_07_in21 = imem03_in[83:80];
    default: op1_07_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv21 = 1;
    7: op1_07_inv21 = 1;
    11: op1_07_inv21 = 1;
    12: op1_07_inv21 = 1;
    13: op1_07_inv21 = 1;
    14: op1_07_inv21 = 1;
    15: op1_07_inv21 = 1;
    18: op1_07_inv21 = 1;
    19: op1_07_inv21 = 1;
    22: op1_07_inv21 = 1;
    23: op1_07_inv21 = 1;
    24: op1_07_inv21 = 1;
    25: op1_07_inv21 = 1;
    26: op1_07_inv21 = 1;
    27: op1_07_inv21 = 1;
    34: op1_07_inv21 = 1;
    35: op1_07_inv21 = 1;
    36: op1_07_inv21 = 1;
    37: op1_07_inv21 = 1;
    38: op1_07_inv21 = 1;
    39: op1_07_inv21 = 1;
    40: op1_07_inv21 = 1;
    41: op1_07_inv21 = 1;
    42: op1_07_inv21 = 1;
    43: op1_07_inv21 = 1;
    44: op1_07_inv21 = 1;
    47: op1_07_inv21 = 1;
    48: op1_07_inv21 = 1;
    49: op1_07_inv21 = 1;
    53: op1_07_inv21 = 1;
    54: op1_07_inv21 = 1;
    61: op1_07_inv21 = 1;
    65: op1_07_inv21 = 1;
    67: op1_07_inv21 = 1;
    69: op1_07_inv21 = 1;
    73: op1_07_inv21 = 1;
    74: op1_07_inv21 = 1;
    77: op1_07_inv21 = 1;
    78: op1_07_inv21 = 1;
    81: op1_07_inv21 = 1;
    82: op1_07_inv21 = 1;
    84: op1_07_inv21 = 1;
    86: op1_07_inv21 = 1;
    87: op1_07_inv21 = 1;
    92: op1_07_inv21 = 1;
    93: op1_07_inv21 = 1;
    94: op1_07_inv21 = 1;
    95: op1_07_inv21 = 1;
    96: op1_07_inv21 = 1;
    default: op1_07_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in22 = reg_0047;
    6: op1_07_in22 = reg_0817;
    78: op1_07_in22 = reg_0817;
    7: op1_07_in22 = reg_0380;
    8: op1_07_in22 = reg_0212;
    9: op1_07_in22 = reg_0546;
    10: op1_07_in22 = reg_0353;
    11: op1_07_in22 = imem05_in[83:80];
    12: op1_07_in22 = imem02_in[119:116];
    13: op1_07_in22 = reg_0421;
    14: op1_07_in22 = imem01_in[111:108];
    36: op1_07_in22 = imem01_in[111:108];
    15: op1_07_in22 = reg_0329;
    16: op1_07_in22 = imem06_in[79:76];
    17: op1_07_in22 = imem07_in[23:20];
    18: op1_07_in22 = reg_0958;
    19: op1_07_in22 = reg_0184;
    20: op1_07_in22 = reg_0956;
    22: op1_07_in22 = imem05_in[107:104];
    23: op1_07_in22 = reg_0066;
    24: op1_07_in22 = reg_0989;
    25: op1_07_in22 = reg_0150;
    26: op1_07_in22 = reg_0218;
    86: op1_07_in22 = reg_0218;
    27: op1_07_in22 = imem06_in[39:36];
    41: op1_07_in22 = imem06_in[39:36];
    28: op1_07_in22 = reg_0424;
    29: op1_07_in22 = reg_0296;
    30: op1_07_in22 = reg_0624;
    32: op1_07_in22 = reg_0876;
    33: op1_07_in22 = reg_0346;
    34: op1_07_in22 = reg_0633;
    35: op1_07_in22 = imem02_in[3:0];
    37: op1_07_in22 = reg_0338;
    38: op1_07_in22 = imem02_in[15:12];
    39: op1_07_in22 = imem05_in[35:32];
    40: op1_07_in22 = reg_0782;
    42: op1_07_in22 = imem01_in[127:124];
    43: op1_07_in22 = reg_0090;
    44: op1_07_in22 = imem05_in[119:116];
    76: op1_07_in22 = imem05_in[119:116];
    46: op1_07_in22 = imem01_in[87:84];
    47: op1_07_in22 = reg_0778;
    48: op1_07_in22 = reg_0426;
    49: op1_07_in22 = reg_0885;
    51: op1_07_in22 = reg_0545;
    52: op1_07_in22 = imem05_in[47:44];
    53: op1_07_in22 = reg_0220;
    54: op1_07_in22 = imem07_in[123:120];
    57: op1_07_in22 = reg_0918;
    58: op1_07_in22 = reg_0110;
    59: op1_07_in22 = reg_0830;
    60: op1_07_in22 = reg_0373;
    61: op1_07_in22 = reg_0261;
    62: op1_07_in22 = reg_0848;
    65: op1_07_in22 = reg_0592;
    66: op1_07_in22 = imem01_in[59:56];
    67: op1_07_in22 = reg_1043;
    68: op1_07_in22 = reg_0376;
    69: op1_07_in22 = reg_0735;
    70: op1_07_in22 = reg_1039;
    71: op1_07_in22 = reg_0083;
    73: op1_07_in22 = reg_0273;
    74: op1_07_in22 = imem01_in[75:72];
    75: op1_07_in22 = reg_0099;
    77: op1_07_in22 = imem05_in[39:36];
    80: op1_07_in22 = reg_0962;
    81: op1_07_in22 = reg_0572;
    82: op1_07_in22 = reg_0514;
    83: op1_07_in22 = reg_0903;
    84: op1_07_in22 = reg_0577;
    85: op1_07_in22 = reg_0225;
    87: op1_07_in22 = reg_0439;
    89: op1_07_in22 = reg_1019;
    90: op1_07_in22 = reg_1056;
    91: op1_07_in22 = imem01_in[55:52];
    92: op1_07_in22 = reg_1037;
    93: op1_07_in22 = reg_0041;
    94: op1_07_in22 = reg_0511;
    95: op1_07_in22 = imem04_in[83:80];
    96: op1_07_in22 = reg_0268;
    97: op1_07_in22 = reg_0836;
    default: op1_07_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_07_inv22 = 1;
    12: op1_07_inv22 = 1;
    13: op1_07_inv22 = 1;
    14: op1_07_inv22 = 1;
    15: op1_07_inv22 = 1;
    16: op1_07_inv22 = 1;
    19: op1_07_inv22 = 1;
    20: op1_07_inv22 = 1;
    22: op1_07_inv22 = 1;
    25: op1_07_inv22 = 1;
    27: op1_07_inv22 = 1;
    29: op1_07_inv22 = 1;
    32: op1_07_inv22 = 1;
    36: op1_07_inv22 = 1;
    37: op1_07_inv22 = 1;
    38: op1_07_inv22 = 1;
    39: op1_07_inv22 = 1;
    40: op1_07_inv22 = 1;
    41: op1_07_inv22 = 1;
    42: op1_07_inv22 = 1;
    44: op1_07_inv22 = 1;
    47: op1_07_inv22 = 1;
    48: op1_07_inv22 = 1;
    53: op1_07_inv22 = 1;
    57: op1_07_inv22 = 1;
    60: op1_07_inv22 = 1;
    61: op1_07_inv22 = 1;
    62: op1_07_inv22 = 1;
    65: op1_07_inv22 = 1;
    66: op1_07_inv22 = 1;
    67: op1_07_inv22 = 1;
    69: op1_07_inv22 = 1;
    70: op1_07_inv22 = 1;
    71: op1_07_inv22 = 1;
    75: op1_07_inv22 = 1;
    78: op1_07_inv22 = 1;
    81: op1_07_inv22 = 1;
    85: op1_07_inv22 = 1;
    86: op1_07_inv22 = 1;
    87: op1_07_inv22 = 1;
    89: op1_07_inv22 = 1;
    91: op1_07_inv22 = 1;
    93: op1_07_inv22 = 1;
    96: op1_07_inv22 = 1;
    97: op1_07_inv22 = 1;
    default: op1_07_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in23 = reg_0065;
    6: op1_07_in23 = reg_0830;
    7: op1_07_in23 = reg_0368;
    8: op1_07_in23 = reg_0205;
    9: op1_07_in23 = reg_0551;
    10: op1_07_in23 = reg_0350;
    11: op1_07_in23 = imem05_in[87:84];
    12: op1_07_in23 = imem02_in[123:120];
    13: op1_07_in23 = reg_0426;
    14: op1_07_in23 = reg_0013;
    36: op1_07_in23 = reg_0013;
    15: op1_07_in23 = reg_0086;
    32: op1_07_in23 = reg_0086;
    16: op1_07_in23 = reg_0614;
    17: op1_07_in23 = imem07_in[55:52];
    18: op1_07_in23 = reg_0967;
    20: op1_07_in23 = reg_0946;
    22: op1_07_in23 = imem05_in[111:108];
    23: op1_07_in23 = reg_0068;
    24: op1_07_in23 = reg_0543;
    25: op1_07_in23 = reg_0152;
    26: op1_07_in23 = reg_0274;
    27: op1_07_in23 = imem06_in[51:48];
    28: op1_07_in23 = reg_0429;
    29: op1_07_in23 = reg_0054;
    30: op1_07_in23 = reg_0617;
    33: op1_07_in23 = reg_0581;
    34: op1_07_in23 = reg_0344;
    35: op1_07_in23 = imem02_in[11:8];
    37: op1_07_in23 = reg_0037;
    38: op1_07_in23 = imem02_in[43:40];
    39: op1_07_in23 = imem05_in[47:44];
    40: op1_07_in23 = reg_0783;
    87: op1_07_in23 = reg_0783;
    41: op1_07_in23 = imem06_in[91:88];
    42: op1_07_in23 = reg_0223;
    43: op1_07_in23 = reg_0310;
    44: op1_07_in23 = imem05_in[123:120];
    46: op1_07_in23 = imem01_in[111:108];
    47: op1_07_in23 = reg_1016;
    48: op1_07_in23 = reg_0427;
    49: op1_07_in23 = reg_0735;
    51: op1_07_in23 = imem07_in[23:20];
    52: op1_07_in23 = imem05_in[95:92];
    53: op1_07_in23 = reg_0533;
    69: op1_07_in23 = reg_0533;
    54: op1_07_in23 = reg_0704;
    57: op1_07_in23 = reg_0762;
    58: op1_07_in23 = imem02_in[27:24];
    59: op1_07_in23 = reg_0227;
    60: op1_07_in23 = reg_0312;
    61: op1_07_in23 = reg_0291;
    62: op1_07_in23 = reg_0067;
    65: op1_07_in23 = reg_0503;
    66: op1_07_in23 = imem01_in[83:80];
    67: op1_07_in23 = reg_1037;
    68: op1_07_in23 = reg_0820;
    70: op1_07_in23 = reg_0496;
    71: op1_07_in23 = reg_0884;
    73: op1_07_in23 = imem02_in[15:12];
    74: op1_07_in23 = reg_0969;
    75: op1_07_in23 = reg_0307;
    76: op1_07_in23 = reg_0217;
    77: op1_07_in23 = imem05_in[43:40];
    78: op1_07_in23 = reg_0926;
    80: op1_07_in23 = reg_0831;
    81: op1_07_in23 = reg_0580;
    82: op1_07_in23 = reg_1031;
    83: op1_07_in23 = reg_0727;
    84: op1_07_in23 = reg_0550;
    85: op1_07_in23 = reg_0522;
    86: op1_07_in23 = reg_0713;
    89: op1_07_in23 = reg_0025;
    90: op1_07_in23 = reg_0234;
    91: op1_07_in23 = imem01_in[75:72];
    92: op1_07_in23 = reg_1040;
    93: op1_07_in23 = reg_0071;
    94: op1_07_in23 = reg_0390;
    95: op1_07_in23 = imem04_in[111:108];
    96: op1_07_in23 = reg_0646;
    97: op1_07_in23 = reg_0363;
    default: op1_07_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv23 = 1;
    6: op1_07_inv23 = 1;
    8: op1_07_inv23 = 1;
    9: op1_07_inv23 = 1;
    11: op1_07_inv23 = 1;
    13: op1_07_inv23 = 1;
    15: op1_07_inv23 = 1;
    16: op1_07_inv23 = 1;
    17: op1_07_inv23 = 1;
    18: op1_07_inv23 = 1;
    22: op1_07_inv23 = 1;
    23: op1_07_inv23 = 1;
    26: op1_07_inv23 = 1;
    27: op1_07_inv23 = 1;
    28: op1_07_inv23 = 1;
    30: op1_07_inv23 = 1;
    32: op1_07_inv23 = 1;
    38: op1_07_inv23 = 1;
    43: op1_07_inv23 = 1;
    44: op1_07_inv23 = 1;
    47: op1_07_inv23 = 1;
    51: op1_07_inv23 = 1;
    52: op1_07_inv23 = 1;
    53: op1_07_inv23 = 1;
    54: op1_07_inv23 = 1;
    59: op1_07_inv23 = 1;
    60: op1_07_inv23 = 1;
    61: op1_07_inv23 = 1;
    65: op1_07_inv23 = 1;
    67: op1_07_inv23 = 1;
    68: op1_07_inv23 = 1;
    69: op1_07_inv23 = 1;
    71: op1_07_inv23 = 1;
    73: op1_07_inv23 = 1;
    75: op1_07_inv23 = 1;
    76: op1_07_inv23 = 1;
    77: op1_07_inv23 = 1;
    81: op1_07_inv23 = 1;
    83: op1_07_inv23 = 1;
    84: op1_07_inv23 = 1;
    85: op1_07_inv23 = 1;
    89: op1_07_inv23 = 1;
    90: op1_07_inv23 = 1;
    92: op1_07_inv23 = 1;
    93: op1_07_inv23 = 1;
    96: op1_07_inv23 = 1;
    97: op1_07_inv23 = 1;
    default: op1_07_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in24 = reg_0066;
    6: op1_07_in24 = reg_0831;
    7: op1_07_in24 = reg_0027;
    8: op1_07_in24 = reg_0206;
    9: op1_07_in24 = reg_0277;
    10: op1_07_in24 = reg_0095;
    11: op1_07_in24 = imem05_in[103:100];
    12: op1_07_in24 = reg_0646;
    13: op1_07_in24 = reg_0165;
    14: op1_07_in24 = reg_1055;
    15: op1_07_in24 = reg_0087;
    16: op1_07_in24 = reg_0624;
    17: op1_07_in24 = imem07_in[59:56];
    18: op1_07_in24 = reg_0945;
    20: op1_07_in24 = reg_0953;
    22: op1_07_in24 = imem05_in[115:112];
    23: op1_07_in24 = reg_0736;
    24: op1_07_in24 = reg_0557;
    25: op1_07_in24 = reg_0153;
    26: op1_07_in24 = reg_0811;
    42: op1_07_in24 = reg_0811;
    27: op1_07_in24 = reg_0625;
    28: op1_07_in24 = reg_0419;
    29: op1_07_in24 = reg_0738;
    30: op1_07_in24 = reg_0381;
    32: op1_07_in24 = reg_0261;
    33: op1_07_in24 = reg_0823;
    34: op1_07_in24 = reg_0295;
    35: op1_07_in24 = imem02_in[19:16];
    36: op1_07_in24 = reg_0510;
    37: op1_07_in24 = reg_0762;
    38: op1_07_in24 = imem02_in[55:52];
    39: op1_07_in24 = imem05_in[59:56];
    40: op1_07_in24 = reg_0387;
    41: op1_07_in24 = imem06_in[107:104];
    43: op1_07_in24 = reg_0077;
    44: op1_07_in24 = reg_0963;
    46: op1_07_in24 = reg_0786;
    47: op1_07_in24 = reg_0507;
    48: op1_07_in24 = reg_0640;
    49: op1_07_in24 = reg_0791;
    51: op1_07_in24 = imem07_in[67:64];
    52: op1_07_in24 = imem05_in[111:108];
    53: op1_07_in24 = reg_0627;
    54: op1_07_in24 = reg_0719;
    87: op1_07_in24 = reg_0719;
    57: op1_07_in24 = reg_0218;
    58: op1_07_in24 = imem02_in[123:120];
    59: op1_07_in24 = reg_0304;
    60: op1_07_in24 = reg_0820;
    61: op1_07_in24 = imem03_in[31:28];
    62: op1_07_in24 = reg_0809;
    65: op1_07_in24 = reg_0487;
    66: op1_07_in24 = imem01_in[99:96];
    67: op1_07_in24 = reg_1040;
    68: op1_07_in24 = reg_0822;
    69: op1_07_in24 = reg_0698;
    70: op1_07_in24 = reg_0798;
    85: op1_07_in24 = reg_0798;
    71: op1_07_in24 = imem03_in[19:16];
    73: op1_07_in24 = imem02_in[27:24];
    74: op1_07_in24 = reg_1044;
    75: op1_07_in24 = reg_0547;
    76: op1_07_in24 = reg_0655;
    77: op1_07_in24 = imem05_in[79:76];
    78: op1_07_in24 = reg_0439;
    80: op1_07_in24 = reg_0501;
    81: op1_07_in24 = reg_0445;
    82: op1_07_in24 = reg_1041;
    83: op1_07_in24 = reg_0805;
    84: op1_07_in24 = reg_0870;
    86: op1_07_in24 = reg_0341;
    89: op1_07_in24 = reg_0338;
    90: op1_07_in24 = reg_0225;
    91: op1_07_in24 = imem01_in[91:88];
    92: op1_07_in24 = reg_0737;
    93: op1_07_in24 = reg_0542;
    94: op1_07_in24 = reg_0913;
    95: op1_07_in24 = imem04_in[119:116];
    96: op1_07_in24 = reg_0675;
    97: op1_07_in24 = reg_0301;
    default: op1_07_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv24 = 1;
    9: op1_07_inv24 = 1;
    10: op1_07_inv24 = 1;
    11: op1_07_inv24 = 1;
    12: op1_07_inv24 = 1;
    18: op1_07_inv24 = 1;
    20: op1_07_inv24 = 1;
    22: op1_07_inv24 = 1;
    24: op1_07_inv24 = 1;
    25: op1_07_inv24 = 1;
    27: op1_07_inv24 = 1;
    30: op1_07_inv24 = 1;
    40: op1_07_inv24 = 1;
    42: op1_07_inv24 = 1;
    43: op1_07_inv24 = 1;
    44: op1_07_inv24 = 1;
    49: op1_07_inv24 = 1;
    51: op1_07_inv24 = 1;
    53: op1_07_inv24 = 1;
    59: op1_07_inv24 = 1;
    60: op1_07_inv24 = 1;
    62: op1_07_inv24 = 1;
    65: op1_07_inv24 = 1;
    68: op1_07_inv24 = 1;
    70: op1_07_inv24 = 1;
    71: op1_07_inv24 = 1;
    73: op1_07_inv24 = 1;
    76: op1_07_inv24 = 1;
    81: op1_07_inv24 = 1;
    83: op1_07_inv24 = 1;
    89: op1_07_inv24 = 1;
    94: op1_07_inv24 = 1;
    default: op1_07_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in25 = reg_0067;
    6: op1_07_in25 = reg_0824;
    7: op1_07_in25 = reg_0026;
    8: op1_07_in25 = imem01_in[47:44];
    9: op1_07_in25 = reg_0285;
    10: op1_07_in25 = reg_0090;
    11: op1_07_in25 = imem05_in[111:108];
    12: op1_07_in25 = reg_0651;
    13: op1_07_in25 = reg_0161;
    14: op1_07_in25 = reg_0233;
    15: op1_07_in25 = imem03_in[19:16];
    16: op1_07_in25 = reg_0621;
    17: op1_07_in25 = imem07_in[103:100];
    18: op1_07_in25 = reg_0947;
    20: op1_07_in25 = reg_0972;
    22: op1_07_in25 = reg_0958;
    23: op1_07_in25 = reg_0058;
    24: op1_07_in25 = reg_0550;
    25: op1_07_in25 = reg_0144;
    26: op1_07_in25 = reg_0221;
    27: op1_07_in25 = reg_0624;
    28: op1_07_in25 = reg_0434;
    29: op1_07_in25 = reg_0053;
    30: op1_07_in25 = reg_0042;
    32: op1_07_in25 = reg_0884;
    43: op1_07_in25 = reg_0884;
    33: op1_07_in25 = reg_0765;
    34: op1_07_in25 = reg_0399;
    35: op1_07_in25 = imem02_in[27:24];
    36: op1_07_in25 = reg_0230;
    37: op1_07_in25 = reg_0776;
    38: op1_07_in25 = imem02_in[91:88];
    39: op1_07_in25 = imem05_in[75:72];
    40: op1_07_in25 = reg_0390;
    41: op1_07_in25 = reg_0533;
    42: op1_07_in25 = reg_0219;
    44: op1_07_in25 = reg_0966;
    46: op1_07_in25 = reg_0779;
    47: op1_07_in25 = reg_0909;
    48: op1_07_in25 = reg_0431;
    49: op1_07_in25 = imem01_in[63:60];
    51: op1_07_in25 = imem07_in[71:68];
    52: op1_07_in25 = reg_0951;
    53: op1_07_in25 = reg_0595;
    54: op1_07_in25 = reg_0723;
    57: op1_07_in25 = reg_1056;
    58: op1_07_in25 = reg_0341;
    59: op1_07_in25 = reg_0232;
    60: op1_07_in25 = reg_0513;
    61: op1_07_in25 = imem03_in[63:60];
    62: op1_07_in25 = reg_0732;
    65: op1_07_in25 = reg_1052;
    66: op1_07_in25 = imem01_in[103:100];
    67: op1_07_in25 = reg_0304;
    68: op1_07_in25 = reg_0985;
    69: op1_07_in25 = reg_0632;
    70: op1_07_in25 = reg_0604;
    71: op1_07_in25 = imem03_in[35:32];
    73: op1_07_in25 = imem02_in[75:72];
    74: op1_07_in25 = reg_0962;
    75: op1_07_in25 = reg_0298;
    76: op1_07_in25 = reg_0140;
    77: op1_07_in25 = imem05_in[87:84];
    78: op1_07_in25 = reg_0863;
    80: op1_07_in25 = reg_0111;
    81: op1_07_in25 = reg_0307;
    82: op1_07_in25 = reg_0555;
    83: op1_07_in25 = reg_0532;
    84: op1_07_in25 = reg_0430;
    85: op1_07_in25 = reg_0869;
    86: op1_07_in25 = imem03_in[3:0];
    87: op1_07_in25 = reg_0857;
    89: op1_07_in25 = reg_0926;
    90: op1_07_in25 = reg_1039;
    91: op1_07_in25 = imem01_in[119:116];
    92: op1_07_in25 = reg_0616;
    93: op1_07_in25 = reg_0856;
    94: op1_07_in25 = reg_0586;
    95: op1_07_in25 = reg_0405;
    96: op1_07_in25 = reg_0695;
    97: op1_07_in25 = reg_0763;
    default: op1_07_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_07_inv25 = 1;
    9: op1_07_inv25 = 1;
    11: op1_07_inv25 = 1;
    15: op1_07_inv25 = 1;
    18: op1_07_inv25 = 1;
    23: op1_07_inv25 = 1;
    24: op1_07_inv25 = 1;
    25: op1_07_inv25 = 1;
    26: op1_07_inv25 = 1;
    28: op1_07_inv25 = 1;
    29: op1_07_inv25 = 1;
    30: op1_07_inv25 = 1;
    32: op1_07_inv25 = 1;
    35: op1_07_inv25 = 1;
    37: op1_07_inv25 = 1;
    44: op1_07_inv25 = 1;
    46: op1_07_inv25 = 1;
    48: op1_07_inv25 = 1;
    49: op1_07_inv25 = 1;
    52: op1_07_inv25 = 1;
    53: op1_07_inv25 = 1;
    59: op1_07_inv25 = 1;
    61: op1_07_inv25 = 1;
    65: op1_07_inv25 = 1;
    66: op1_07_inv25 = 1;
    70: op1_07_inv25 = 1;
    71: op1_07_inv25 = 1;
    73: op1_07_inv25 = 1;
    80: op1_07_inv25 = 1;
    81: op1_07_inv25 = 1;
    84: op1_07_inv25 = 1;
    87: op1_07_inv25 = 1;
    89: op1_07_inv25 = 1;
    91: op1_07_inv25 = 1;
    92: op1_07_inv25 = 1;
    93: op1_07_inv25 = 1;
    94: op1_07_inv25 = 1;
    95: op1_07_inv25 = 1;
    96: op1_07_inv25 = 1;
    default: op1_07_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in26 = reg_0068;
    6: op1_07_in26 = reg_0569;
    7: op1_07_in26 = reg_0036;
    8: op1_07_in26 = imem01_in[51:48];
    9: op1_07_in26 = reg_0046;
    10: op1_07_in26 = reg_0093;
    11: op1_07_in26 = imem05_in[123:120];
    12: op1_07_in26 = reg_0652;
    13: op1_07_in26 = reg_0167;
    14: op1_07_in26 = reg_0242;
    15: op1_07_in26 = imem03_in[43:40];
    16: op1_07_in26 = reg_0609;
    17: op1_07_in26 = reg_0722;
    18: op1_07_in26 = reg_0863;
    20: op1_07_in26 = imem05_in[15:12];
    22: op1_07_in26 = reg_0956;
    23: op1_07_in26 = reg_0875;
    24: op1_07_in26 = reg_0877;
    25: op1_07_in26 = imem06_in[35:32];
    26: op1_07_in26 = reg_0249;
    27: op1_07_in26 = reg_0622;
    28: op1_07_in26 = reg_0446;
    29: op1_07_in26 = reg_0864;
    30: op1_07_in26 = reg_0384;
    32: op1_07_in26 = reg_0872;
    33: op1_07_in26 = reg_0767;
    34: op1_07_in26 = reg_0349;
    35: op1_07_in26 = imem02_in[43:40];
    36: op1_07_in26 = reg_1036;
    37: op1_07_in26 = reg_0261;
    38: op1_07_in26 = imem02_in[107:104];
    39: op1_07_in26 = imem05_in[79:76];
    40: op1_07_in26 = reg_0380;
    41: op1_07_in26 = reg_0020;
    42: op1_07_in26 = reg_0607;
    49: op1_07_in26 = reg_0607;
    43: op1_07_in26 = imem03_in[3:0];
    44: op1_07_in26 = reg_0967;
    46: op1_07_in26 = reg_0223;
    47: op1_07_in26 = reg_0302;
    48: op1_07_in26 = reg_0180;
    51: op1_07_in26 = imem07_in[79:76];
    52: op1_07_in26 = reg_0946;
    53: op1_07_in26 = reg_0387;
    54: op1_07_in26 = reg_0726;
    57: op1_07_in26 = reg_1035;
    58: op1_07_in26 = reg_0656;
    59: op1_07_in26 = reg_0111;
    60: op1_07_in26 = reg_0844;
    61: op1_07_in26 = imem03_in[83:80];
    62: op1_07_in26 = reg_0332;
    65: op1_07_in26 = reg_0830;
    66: op1_07_in26 = imem01_in[111:108];
    67: op1_07_in26 = reg_0116;
    80: op1_07_in26 = reg_0116;
    68: op1_07_in26 = reg_0976;
    69: op1_07_in26 = reg_0222;
    70: op1_07_in26 = reg_0737;
    71: op1_07_in26 = imem03_in[39:36];
    73: op1_07_in26 = imem02_in[123:120];
    74: op1_07_in26 = reg_0514;
    85: op1_07_in26 = reg_0514;
    90: op1_07_in26 = reg_0514;
    75: op1_07_in26 = reg_0661;
    76: op1_07_in26 = reg_0269;
    77: op1_07_in26 = reg_0944;
    78: op1_07_in26 = reg_0011;
    81: op1_07_in26 = reg_0245;
    82: op1_07_in26 = reg_0114;
    83: op1_07_in26 = reg_0431;
    84: op1_07_in26 = reg_0586;
    86: op1_07_in26 = imem03_in[15:12];
    87: op1_07_in26 = reg_0807;
    89: op1_07_in26 = reg_0889;
    91: op1_07_in26 = imem01_in[123:120];
    92: op1_07_in26 = reg_1017;
    93: op1_07_in26 = imem05_in[11:8];
    94: op1_07_in26 = reg_0909;
    95: op1_07_in26 = reg_0937;
    96: op1_07_in26 = reg_0892;
    97: op1_07_in26 = reg_0331;
    default: op1_07_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_07_inv26 = 1;
    12: op1_07_inv26 = 1;
    14: op1_07_inv26 = 1;
    15: op1_07_inv26 = 1;
    17: op1_07_inv26 = 1;
    22: op1_07_inv26 = 1;
    24: op1_07_inv26 = 1;
    25: op1_07_inv26 = 1;
    34: op1_07_inv26 = 1;
    35: op1_07_inv26 = 1;
    37: op1_07_inv26 = 1;
    41: op1_07_inv26 = 1;
    43: op1_07_inv26 = 1;
    46: op1_07_inv26 = 1;
    47: op1_07_inv26 = 1;
    48: op1_07_inv26 = 1;
    49: op1_07_inv26 = 1;
    51: op1_07_inv26 = 1;
    52: op1_07_inv26 = 1;
    57: op1_07_inv26 = 1;
    62: op1_07_inv26 = 1;
    65: op1_07_inv26 = 1;
    66: op1_07_inv26 = 1;
    69: op1_07_inv26 = 1;
    71: op1_07_inv26 = 1;
    74: op1_07_inv26 = 1;
    76: op1_07_inv26 = 1;
    77: op1_07_inv26 = 1;
    80: op1_07_inv26 = 1;
    82: op1_07_inv26 = 1;
    86: op1_07_inv26 = 1;
    87: op1_07_inv26 = 1;
    93: op1_07_inv26 = 1;
    94: op1_07_inv26 = 1;
    default: op1_07_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in27 = reg_0063;
    6: op1_07_in27 = reg_0591;
    7: op1_07_in27 = reg_0030;
    8: op1_07_in27 = imem01_in[91:88];
    9: op1_07_in27 = reg_0054;
    10: op1_07_in27 = imem03_in[55:52];
    11: op1_07_in27 = reg_0962;
    12: op1_07_in27 = reg_0325;
    13: op1_07_in27 = reg_0169;
    14: op1_07_in27 = reg_0240;
    15: op1_07_in27 = imem03_in[51:48];
    16: op1_07_in27 = reg_0619;
    17: op1_07_in27 = reg_0704;
    18: op1_07_in27 = reg_0215;
    20: op1_07_in27 = imem05_in[35:32];
    22: op1_07_in27 = reg_0949;
    44: op1_07_in27 = reg_0949;
    23: op1_07_in27 = reg_0777;
    24: op1_07_in27 = reg_0289;
    25: op1_07_in27 = imem06_in[43:40];
    26: op1_07_in27 = reg_0769;
    27: op1_07_in27 = reg_0379;
    28: op1_07_in27 = reg_0438;
    29: op1_07_in27 = reg_0044;
    62: op1_07_in27 = reg_0044;
    30: op1_07_in27 = reg_1029;
    32: op1_07_in27 = imem03_in[87:84];
    61: op1_07_in27 = imem03_in[87:84];
    33: op1_07_in27 = reg_0312;
    34: op1_07_in27 = reg_0402;
    35: op1_07_in27 = imem02_in[51:48];
    36: op1_07_in27 = reg_0871;
    37: op1_07_in27 = reg_0484;
    38: op1_07_in27 = imem02_in[111:108];
    39: op1_07_in27 = imem05_in[111:108];
    40: op1_07_in27 = reg_0332;
    41: op1_07_in27 = reg_0371;
    42: op1_07_in27 = reg_1039;
    43: op1_07_in27 = imem03_in[7:4];
    46: op1_07_in27 = reg_0247;
    47: op1_07_in27 = reg_0064;
    48: op1_07_in27 = reg_0161;
    49: op1_07_in27 = reg_0501;
    51: op1_07_in27 = imem07_in[115:112];
    52: op1_07_in27 = reg_0774;
    53: op1_07_in27 = reg_0356;
    54: op1_07_in27 = reg_0724;
    57: op1_07_in27 = reg_1052;
    58: op1_07_in27 = reg_0026;
    59: op1_07_in27 = reg_0512;
    60: op1_07_in27 = reg_0374;
    65: op1_07_in27 = reg_0227;
    66: op1_07_in27 = reg_0933;
    67: op1_07_in27 = reg_0733;
    68: op1_07_in27 = reg_0997;
    69: op1_07_in27 = reg_0915;
    70: op1_07_in27 = reg_0740;
    71: op1_07_in27 = imem03_in[75:72];
    73: op1_07_in27 = reg_0650;
    74: op1_07_in27 = reg_1037;
    75: op1_07_in27 = reg_1008;
    76: op1_07_in27 = reg_0583;
    77: op1_07_in27 = reg_0217;
    78: op1_07_in27 = reg_0293;
    80: op1_07_in27 = reg_1033;
    81: op1_07_in27 = reg_0585;
    82: op1_07_in27 = imem02_in[19:16];
    83: op1_07_in27 = reg_0185;
    84: op1_07_in27 = reg_0507;
    85: op1_07_in27 = reg_0737;
    86: op1_07_in27 = imem03_in[23:20];
    87: op1_07_in27 = reg_0370;
    89: op1_07_in27 = reg_0440;
    90: op1_07_in27 = reg_0830;
    91: op1_07_in27 = reg_0105;
    92: op1_07_in27 = reg_0925;
    93: op1_07_in27 = imem05_in[63:60];
    94: op1_07_in27 = reg_0809;
    95: op1_07_in27 = reg_1009;
    96: op1_07_in27 = reg_0972;
    97: op1_07_in27 = reg_1049;
    default: op1_07_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_07_inv27 = 1;
    8: op1_07_inv27 = 1;
    10: op1_07_inv27 = 1;
    12: op1_07_inv27 = 1;
    13: op1_07_inv27 = 1;
    14: op1_07_inv27 = 1;
    15: op1_07_inv27 = 1;
    17: op1_07_inv27 = 1;
    18: op1_07_inv27 = 1;
    22: op1_07_inv27 = 1;
    23: op1_07_inv27 = 1;
    25: op1_07_inv27 = 1;
    26: op1_07_inv27 = 1;
    28: op1_07_inv27 = 1;
    30: op1_07_inv27 = 1;
    34: op1_07_inv27 = 1;
    35: op1_07_inv27 = 1;
    36: op1_07_inv27 = 1;
    37: op1_07_inv27 = 1;
    40: op1_07_inv27 = 1;
    41: op1_07_inv27 = 1;
    44: op1_07_inv27 = 1;
    53: op1_07_inv27 = 1;
    54: op1_07_inv27 = 1;
    57: op1_07_inv27 = 1;
    60: op1_07_inv27 = 1;
    66: op1_07_inv27 = 1;
    67: op1_07_inv27 = 1;
    68: op1_07_inv27 = 1;
    70: op1_07_inv27 = 1;
    74: op1_07_inv27 = 1;
    75: op1_07_inv27 = 1;
    76: op1_07_inv27 = 1;
    77: op1_07_inv27 = 1;
    78: op1_07_inv27 = 1;
    82: op1_07_inv27 = 1;
    86: op1_07_inv27 = 1;
    89: op1_07_inv27 = 1;
    91: op1_07_inv27 = 1;
    92: op1_07_inv27 = 1;
    93: op1_07_inv27 = 1;
    94: op1_07_inv27 = 1;
    95: op1_07_inv27 = 1;
    default: op1_07_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in28 = reg_0069;
    6: op1_07_in28 = reg_0588;
    7: op1_07_in28 = imem07_in[11:8];
    8: op1_07_in28 = reg_0523;
    9: op1_07_in28 = reg_0078;
    10: op1_07_in28 = imem03_in[75:72];
    11: op1_07_in28 = reg_0968;
    12: op1_07_in28 = reg_0310;
    13: op1_07_in28 = reg_0164;
    14: op1_07_in28 = reg_1056;
    15: op1_07_in28 = imem03_in[67:64];
    16: op1_07_in28 = reg_0615;
    17: op1_07_in28 = reg_0720;
    18: op1_07_in28 = reg_0900;
    20: op1_07_in28 = reg_0130;
    22: op1_07_in28 = reg_0965;
    23: op1_07_in28 = reg_0855;
    24: op1_07_in28 = reg_0290;
    25: op1_07_in28 = imem06_in[47:44];
    26: op1_07_in28 = reg_0226;
    27: op1_07_in28 = reg_0392;
    28: op1_07_in28 = reg_0174;
    29: op1_07_in28 = reg_0021;
    30: op1_07_in28 = reg_0808;
    32: op1_07_in28 = imem03_in[95:92];
    86: op1_07_in28 = imem03_in[95:92];
    33: op1_07_in28 = reg_0844;
    34: op1_07_in28 = reg_0031;
    35: op1_07_in28 = imem02_in[63:60];
    36: op1_07_in28 = reg_1018;
    37: op1_07_in28 = imem03_in[79:76];
    38: op1_07_in28 = imem02_in[127:124];
    39: op1_07_in28 = reg_0973;
    40: op1_07_in28 = reg_0241;
    41: op1_07_in28 = reg_0782;
    42: op1_07_in28 = reg_0501;
    43: op1_07_in28 = imem03_in[71:68];
    44: op1_07_in28 = reg_0821;
    46: op1_07_in28 = reg_0811;
    47: op1_07_in28 = reg_0444;
    48: op1_07_in28 = reg_0166;
    49: op1_07_in28 = reg_0496;
    51: op1_07_in28 = reg_0722;
    52: op1_07_in28 = reg_0488;
    53: op1_07_in28 = reg_0294;
    54: op1_07_in28 = reg_0718;
    57: op1_07_in28 = reg_0522;
    58: op1_07_in28 = reg_0837;
    59: op1_07_in28 = reg_0109;
    60: op1_07_in28 = reg_0980;
    61: op1_07_in28 = reg_0006;
    71: op1_07_in28 = reg_0006;
    62: op1_07_in28 = imem05_in[19:16];
    65: op1_07_in28 = reg_0354;
    66: op1_07_in28 = reg_0238;
    67: op1_07_in28 = reg_0114;
    68: op1_07_in28 = imem04_in[3:0];
    69: op1_07_in28 = reg_0630;
    70: op1_07_in28 = reg_0111;
    73: op1_07_in28 = reg_0916;
    74: op1_07_in28 = reg_0227;
    75: op1_07_in28 = reg_0581;
    76: op1_07_in28 = reg_0688;
    77: op1_07_in28 = reg_0143;
    78: op1_07_in28 = reg_0289;
    80: op1_07_in28 = reg_0877;
    81: op1_07_in28 = reg_0046;
    82: op1_07_in28 = imem02_in[35:32];
    84: op1_07_in28 = reg_0067;
    85: op1_07_in28 = reg_0616;
    87: op1_07_in28 = reg_0220;
    89: op1_07_in28 = reg_0895;
    90: op1_07_in28 = reg_0737;
    91: op1_07_in28 = reg_0122;
    92: op1_07_in28 = reg_0232;
    93: op1_07_in28 = imem05_in[71:68];
    94: op1_07_in28 = reg_0732;
    95: op1_07_in28 = reg_0507;
    96: op1_07_in28 = reg_0960;
    97: op1_07_in28 = reg_0779;
    default: op1_07_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv28 = 1;
    9: op1_07_inv28 = 1;
    14: op1_07_inv28 = 1;
    16: op1_07_inv28 = 1;
    17: op1_07_inv28 = 1;
    23: op1_07_inv28 = 1;
    24: op1_07_inv28 = 1;
    27: op1_07_inv28 = 1;
    28: op1_07_inv28 = 1;
    29: op1_07_inv28 = 1;
    32: op1_07_inv28 = 1;
    33: op1_07_inv28 = 1;
    35: op1_07_inv28 = 1;
    43: op1_07_inv28 = 1;
    44: op1_07_inv28 = 1;
    46: op1_07_inv28 = 1;
    48: op1_07_inv28 = 1;
    51: op1_07_inv28 = 1;
    52: op1_07_inv28 = 1;
    61: op1_07_inv28 = 1;
    62: op1_07_inv28 = 1;
    65: op1_07_inv28 = 1;
    70: op1_07_inv28 = 1;
    74: op1_07_inv28 = 1;
    76: op1_07_inv28 = 1;
    81: op1_07_inv28 = 1;
    85: op1_07_inv28 = 1;
    92: op1_07_inv28 = 1;
    95: op1_07_inv28 = 1;
    96: op1_07_inv28 = 1;
    default: op1_07_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in29 = reg_0070;
    6: op1_07_in29 = reg_0384;
    7: op1_07_in29 = imem07_in[19:16];
    8: op1_07_in29 = reg_0522;
    9: op1_07_in29 = reg_0041;
    10: op1_07_in29 = imem03_in[103:100];
    43: op1_07_in29 = imem03_in[103:100];
    11: op1_07_in29 = reg_0960;
    12: op1_07_in29 = reg_0342;
    13: op1_07_in29 = reg_0185;
    14: op1_07_in29 = reg_0220;
    15: op1_07_in29 = imem03_in[71:68];
    16: op1_07_in29 = reg_0386;
    17: op1_07_in29 = reg_0726;
    18: op1_07_in29 = reg_0827;
    20: op1_07_in29 = reg_0134;
    22: op1_07_in29 = reg_0946;
    23: op1_07_in29 = reg_0044;
    24: op1_07_in29 = reg_0288;
    25: op1_07_in29 = imem06_in[67:64];
    26: op1_07_in29 = reg_0227;
    27: op1_07_in29 = reg_0404;
    28: op1_07_in29 = reg_0179;
    29: op1_07_in29 = imem05_in[3:0];
    30: op1_07_in29 = reg_0752;
    32: op1_07_in29 = reg_0343;
    33: op1_07_in29 = reg_0985;
    34: op1_07_in29 = reg_0032;
    35: op1_07_in29 = imem02_in[123:120];
    36: op1_07_in29 = reg_0118;
    37: op1_07_in29 = imem03_in[99:96];
    86: op1_07_in29 = imem03_in[99:96];
    38: op1_07_in29 = reg_0658;
    39: op1_07_in29 = reg_0966;
    40: op1_07_in29 = reg_0605;
    41: op1_07_in29 = reg_0783;
    42: op1_07_in29 = reg_0500;
    44: op1_07_in29 = reg_0256;
    46: op1_07_in29 = reg_0238;
    47: op1_07_in29 = reg_0367;
    49: op1_07_in29 = reg_0869;
    51: op1_07_in29 = reg_0704;
    52: op1_07_in29 = reg_0757;
    53: op1_07_in29 = reg_0594;
    54: op1_07_in29 = reg_0744;
    57: op1_07_in29 = reg_1043;
    58: op1_07_in29 = reg_0423;
    59: op1_07_in29 = reg_0117;
    60: op1_07_in29 = reg_0990;
    61: op1_07_in29 = reg_0307;
    62: op1_07_in29 = imem05_in[31:28];
    65: op1_07_in29 = reg_0610;
    66: op1_07_in29 = reg_0501;
    67: op1_07_in29 = reg_0860;
    70: op1_07_in29 = reg_0860;
    68: op1_07_in29 = imem04_in[111:108];
    69: op1_07_in29 = reg_0371;
    71: op1_07_in29 = reg_0012;
    73: op1_07_in29 = reg_0885;
    74: op1_07_in29 = reg_1031;
    75: op1_07_in29 = reg_0385;
    76: op1_07_in29 = reg_0707;
    77: op1_07_in29 = reg_0235;
    78: op1_07_in29 = reg_0755;
    80: op1_07_in29 = imem02_in[75:72];
    81: op1_07_in29 = reg_0823;
    82: op1_07_in29 = imem02_in[51:48];
    84: op1_07_in29 = reg_0065;
    85: op1_07_in29 = reg_0832;
    87: op1_07_in29 = reg_0612;
    89: op1_07_in29 = reg_0595;
    90: op1_07_in29 = reg_0740;
    91: op1_07_in29 = reg_1032;
    92: op1_07_in29 = reg_0769;
    93: op1_07_in29 = imem05_in[103:100];
    94: op1_07_in29 = reg_0764;
    95: op1_07_in29 = reg_0848;
    96: op1_07_in29 = reg_0486;
    97: op1_07_in29 = reg_0767;
    default: op1_07_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_07_inv29 = 1;
    8: op1_07_inv29 = 1;
    9: op1_07_inv29 = 1;
    12: op1_07_inv29 = 1;
    14: op1_07_inv29 = 1;
    17: op1_07_inv29 = 1;
    23: op1_07_inv29 = 1;
    25: op1_07_inv29 = 1;
    26: op1_07_inv29 = 1;
    27: op1_07_inv29 = 1;
    28: op1_07_inv29 = 1;
    30: op1_07_inv29 = 1;
    33: op1_07_inv29 = 1;
    34: op1_07_inv29 = 1;
    36: op1_07_inv29 = 1;
    38: op1_07_inv29 = 1;
    41: op1_07_inv29 = 1;
    42: op1_07_inv29 = 1;
    43: op1_07_inv29 = 1;
    46: op1_07_inv29 = 1;
    54: op1_07_inv29 = 1;
    60: op1_07_inv29 = 1;
    61: op1_07_inv29 = 1;
    62: op1_07_inv29 = 1;
    65: op1_07_inv29 = 1;
    66: op1_07_inv29 = 1;
    67: op1_07_inv29 = 1;
    68: op1_07_inv29 = 1;
    69: op1_07_inv29 = 1;
    74: op1_07_inv29 = 1;
    76: op1_07_inv29 = 1;
    80: op1_07_inv29 = 1;
    81: op1_07_inv29 = 1;
    87: op1_07_inv29 = 1;
    89: op1_07_inv29 = 1;
    92: op1_07_inv29 = 1;
    95: op1_07_inv29 = 1;
    default: op1_07_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_07_in30 = imem05_in[23:20];
    6: op1_07_in30 = reg_0387;
    7: op1_07_in30 = imem07_in[27:24];
    8: op1_07_in30 = reg_0511;
    9: op1_07_in30 = reg_0057;
    47: op1_07_in30 = reg_0057;
    10: op1_07_in30 = imem03_in[111:108];
    11: op1_07_in30 = reg_0262;
    12: op1_07_in30 = reg_0045;
    13: op1_07_in30 = reg_0171;
    14: op1_07_in30 = reg_0234;
    15: op1_07_in30 = imem03_in[75:72];
    16: op1_07_in30 = reg_0409;
    17: op1_07_in30 = reg_0702;
    18: op1_07_in30 = reg_0828;
    20: op1_07_in30 = imem06_in[15:12];
    22: op1_07_in30 = reg_0960;
    23: op1_07_in30 = imem05_in[15:12];
    24: op1_07_in30 = reg_0556;
    25: op1_07_in30 = imem06_in[71:68];
    26: op1_07_in30 = reg_1017;
    90: op1_07_in30 = reg_1017;
    27: op1_07_in30 = reg_0401;
    28: op1_07_in30 = reg_0161;
    29: op1_07_in30 = imem05_in[83:80];
    30: op1_07_in30 = reg_1028;
    32: op1_07_in30 = reg_0346;
    33: op1_07_in30 = reg_0987;
    34: op1_07_in30 = reg_0780;
    35: op1_07_in30 = reg_0666;
    38: op1_07_in30 = reg_0666;
    36: op1_07_in30 = reg_0120;
    37: op1_07_in30 = imem03_in[107:104];
    39: op1_07_in30 = reg_0954;
    40: op1_07_in30 = reg_0017;
    87: op1_07_in30 = reg_0017;
    41: op1_07_in30 = reg_0595;
    42: op1_07_in30 = reg_1037;
    57: op1_07_in30 = reg_1037;
    43: op1_07_in30 = imem03_in[115:112];
    44: op1_07_in30 = reg_0827;
    67: op1_07_in30 = reg_0827;
    46: op1_07_in30 = reg_0249;
    49: op1_07_in30 = reg_0354;
    74: op1_07_in30 = reg_0354;
    51: op1_07_in30 = reg_0719;
    52: op1_07_in30 = reg_0150;
    53: op1_07_in30 = reg_0241;
    54: op1_07_in30 = reg_0029;
    58: op1_07_in30 = reg_0368;
    59: op1_07_in30 = reg_0110;
    60: op1_07_in30 = reg_0976;
    61: op1_07_in30 = reg_0322;
    62: op1_07_in30 = imem05_in[71:68];
    65: op1_07_in30 = reg_0610;
    66: op1_07_in30 = reg_0522;
    68: op1_07_in30 = reg_0536;
    69: op1_07_in30 = reg_0957;
    70: op1_07_in30 = imem02_in[27:24];
    71: op1_07_in30 = reg_0434;
    73: op1_07_in30 = reg_0907;
    75: op1_07_in30 = reg_0551;
    76: op1_07_in30 = reg_0970;
    77: op1_07_in30 = reg_0689;
    78: op1_07_in30 = reg_0566;
    80: op1_07_in30 = imem02_in[91:88];
    81: op1_07_in30 = reg_0397;
    82: op1_07_in30 = imem02_in[67:64];
    84: op1_07_in30 = reg_0627;
    85: op1_07_in30 = reg_0733;
    92: op1_07_in30 = reg_0733;
    86: op1_07_in30 = imem03_in[103:100];
    89: op1_07_in30 = reg_0606;
    91: op1_07_in30 = reg_0337;
    93: op1_07_in30 = imem05_in[107:104];
    94: op1_07_in30 = reg_0061;
    95: op1_07_in30 = reg_0850;
    96: op1_07_in30 = reg_0741;
    97: op1_07_in30 = reg_0597;
    default: op1_07_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv30 = 1;
    9: op1_07_inv30 = 1;
    11: op1_07_inv30 = 1;
    12: op1_07_inv30 = 1;
    17: op1_07_inv30 = 1;
    18: op1_07_inv30 = 1;
    20: op1_07_inv30 = 1;
    25: op1_07_inv30 = 1;
    26: op1_07_inv30 = 1;
    27: op1_07_inv30 = 1;
    28: op1_07_inv30 = 1;
    29: op1_07_inv30 = 1;
    30: op1_07_inv30 = 1;
    32: op1_07_inv30 = 1;
    35: op1_07_inv30 = 1;
    36: op1_07_inv30 = 1;
    37: op1_07_inv30 = 1;
    38: op1_07_inv30 = 1;
    39: op1_07_inv30 = 1;
    41: op1_07_inv30 = 1;
    52: op1_07_inv30 = 1;
    57: op1_07_inv30 = 1;
    60: op1_07_inv30 = 1;
    65: op1_07_inv30 = 1;
    75: op1_07_inv30 = 1;
    77: op1_07_inv30 = 1;
    82: op1_07_inv30 = 1;
    84: op1_07_inv30 = 1;
    85: op1_07_inv30 = 1;
    87: op1_07_inv30 = 1;
    90: op1_07_inv30 = 1;
    91: op1_07_inv30 = 1;
    92: op1_07_inv30 = 1;
    93: op1_07_inv30 = 1;
    default: op1_07_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_07_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_07_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in00 = imem05_in[31:28];
    84: op1_08_in00 = imem05_in[31:28];
    6: op1_08_in00 = reg_0391;
    7: op1_08_in00 = imem07_in[47:44];
    3: op1_08_in00 = imem07_in[47:44];
    8: op1_08_in00 = reg_0503;
    9: op1_08_in00 = imem05_in[39:36];
    10: op1_08_in00 = reg_0586;
    11: op1_08_in00 = reg_0259;
    24: op1_08_in00 = reg_0259;
    12: op1_08_in00 = reg_0052;
    13: op1_08_in00 = imem00_in[11:8];
    14: op1_08_in00 = reg_1050;
    15: op1_08_in00 = imem03_in[95:92];
    4: op1_08_in00 = imem07_in[15:12];
    16: op1_08_in00 = reg_0313;
    17: op1_08_in00 = imem00_in[59:56];
    64: op1_08_in00 = imem00_in[59:56];
    18: op1_08_in00 = reg_0254;
    19: op1_08_in00 = imem00_in[91:88];
    20: op1_08_in00 = imem06_in[43:40];
    21: op1_08_in00 = imem00_in[15:12];
    28: op1_08_in00 = imem00_in[15:12];
    83: op1_08_in00 = imem00_in[15:12];
    22: op1_08_in00 = reg_0256;
    23: op1_08_in00 = imem05_in[47:44];
    25: op1_08_in00 = imem06_in[123:120];
    26: op1_08_in00 = reg_0123;
    27: op1_08_in00 = reg_0799;
    2: op1_08_in00 = imem07_in[95:92];
    29: op1_08_in00 = imem05_in[99:96];
    30: op1_08_in00 = reg_0753;
    31: op1_08_in00 = imem00_in[43:40];
    32: op1_08_in00 = reg_0396;
    33: op1_08_in00 = reg_0981;
    34: op1_08_in00 = reg_0404;
    35: op1_08_in00 = reg_0647;
    36: op1_08_in00 = reg_0112;
    37: op1_08_in00 = reg_0938;
    38: op1_08_in00 = reg_0664;
    39: op1_08_in00 = reg_0968;
    40: op1_08_in00 = reg_0609;
    41: op1_08_in00 = reg_0344;
    42: op1_08_in00 = reg_0227;
    43: op1_08_in00 = reg_0006;
    86: op1_08_in00 = reg_0006;
    44: op1_08_in00 = reg_0896;
    45: op1_08_in00 = imem00_in[71:68];
    56: op1_08_in00 = imem00_in[71:68];
    46: op1_08_in00 = reg_0501;
    47: op1_08_in00 = reg_0864;
    48: op1_08_in00 = imem00_in[31:28];
    79: op1_08_in00 = imem00_in[31:28];
    49: op1_08_in00 = reg_0120;
    50: op1_08_in00 = imem00_in[19:16];
    51: op1_08_in00 = reg_0717;
    52: op1_08_in00 = reg_0138;
    53: op1_08_in00 = reg_0617;
    54: op1_08_in00 = reg_0420;
    55: op1_08_in00 = reg_0409;
    57: op1_08_in00 = reg_0354;
    58: op1_08_in00 = reg_0372;
    59: op1_08_in00 = imem02_in[19:16];
    60: op1_08_in00 = imem04_in[59:56];
    61: op1_08_in00 = reg_0661;
    62: op1_08_in00 = imem05_in[87:84];
    63: op1_08_in00 = imem00_in[55:52];
    65: op1_08_in00 = reg_0740;
    66: op1_08_in00 = reg_1017;
    67: op1_08_in00 = reg_0115;
    68: op1_08_in00 = reg_0265;
    69: op1_08_in00 = imem07_in[11:8];
    70: op1_08_in00 = imem02_in[51:48];
    71: op1_08_in00 = reg_0046;
    72: op1_08_in00 = imem00_in[63:60];
    73: op1_08_in00 = reg_0098;
    74: op1_08_in00 = reg_0304;
    90: op1_08_in00 = reg_0304;
    75: op1_08_in00 = reg_0985;
    76: op1_08_in00 = reg_0145;
    77: op1_08_in00 = reg_0226;
    78: op1_08_in00 = imem07_in[67:64];
    80: op1_08_in00 = imem02_in[99:96];
    81: op1_08_in00 = reg_0596;
    82: op1_08_in00 = imem02_in[115:112];
    85: op1_08_in00 = reg_0103;
    87: op1_08_in00 = reg_0403;
    88: op1_08_in00 = imem00_in[7:4];
    89: op1_08_in00 = imem06_in[3:0];
    91: op1_08_in00 = reg_1023;
    92: op1_08_in00 = reg_0860;
    93: op1_08_in00 = reg_0492;
    94: op1_08_in00 = reg_0243;
    95: op1_08_in00 = reg_0058;
    96: op1_08_in00 = imem06_in[15:12];
    97: op1_08_in00 = reg_0266;
    default: op1_08_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv00 = 1;
    7: op1_08_inv00 = 1;
    10: op1_08_inv00 = 1;
    11: op1_08_inv00 = 1;
    12: op1_08_inv00 = 1;
    13: op1_08_inv00 = 1;
    4: op1_08_inv00 = 1;
    18: op1_08_inv00 = 1;
    20: op1_08_inv00 = 1;
    22: op1_08_inv00 = 1;
    26: op1_08_inv00 = 1;
    27: op1_08_inv00 = 1;
    32: op1_08_inv00 = 1;
    33: op1_08_inv00 = 1;
    39: op1_08_inv00 = 1;
    40: op1_08_inv00 = 1;
    41: op1_08_inv00 = 1;
    43: op1_08_inv00 = 1;
    45: op1_08_inv00 = 1;
    47: op1_08_inv00 = 1;
    48: op1_08_inv00 = 1;
    49: op1_08_inv00 = 1;
    54: op1_08_inv00 = 1;
    55: op1_08_inv00 = 1;
    60: op1_08_inv00 = 1;
    64: op1_08_inv00 = 1;
    70: op1_08_inv00 = 1;
    71: op1_08_inv00 = 1;
    76: op1_08_inv00 = 1;
    77: op1_08_inv00 = 1;
    79: op1_08_inv00 = 1;
    82: op1_08_inv00 = 1;
    83: op1_08_inv00 = 1;
    84: op1_08_inv00 = 1;
    86: op1_08_inv00 = 1;
    87: op1_08_inv00 = 1;
    91: op1_08_inv00 = 1;
    92: op1_08_inv00 = 1;
    94: op1_08_inv00 = 1;
    95: op1_08_inv00 = 1;
    96: op1_08_inv00 = 1;
    97: op1_08_inv00 = 1;
    default: op1_08_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in01 = imem05_in[35:32];
    6: op1_08_in01 = reg_0321;
    7: op1_08_in01 = imem07_in[59:56];
    8: op1_08_in01 = reg_0235;
    9: op1_08_in01 = imem05_in[55:52];
    10: op1_08_in01 = reg_0587;
    11: op1_08_in01 = reg_0260;
    12: op1_08_in01 = reg_0098;
    13: op1_08_in01 = imem00_in[15:12];
    14: op1_08_in01 = reg_0249;
    15: op1_08_in01 = reg_0582;
    4: op1_08_in01 = imem07_in[47:44];
    16: op1_08_in01 = reg_0383;
    17: op1_08_in01 = imem00_in[75:72];
    18: op1_08_in01 = reg_0139;
    19: op1_08_in01 = imem00_in[123:120];
    31: op1_08_in01 = imem00_in[123:120];
    20: op1_08_in01 = imem06_in[63:60];
    21: op1_08_in01 = imem00_in[27:24];
    3: op1_08_in01 = imem07_in[99:96];
    2: op1_08_in01 = imem07_in[99:96];
    22: op1_08_in01 = reg_0491;
    23: op1_08_in01 = imem05_in[67:64];
    24: op1_08_in01 = reg_0755;
    25: op1_08_in01 = reg_0610;
    26: op1_08_in01 = reg_0122;
    27: op1_08_in01 = reg_0752;
    28: op1_08_in01 = imem00_in[59:56];
    29: op1_08_in01 = reg_0963;
    77: op1_08_in01 = reg_0963;
    30: op1_08_in01 = reg_1010;
    53: op1_08_in01 = reg_1010;
    32: op1_08_in01 = reg_0004;
    33: op1_08_in01 = reg_0988;
    34: op1_08_in01 = reg_0595;
    35: op1_08_in01 = reg_0095;
    36: op1_08_in01 = reg_0102;
    49: op1_08_in01 = reg_0102;
    37: op1_08_in01 = reg_0923;
    38: op1_08_in01 = reg_0657;
    39: op1_08_in01 = reg_0961;
    40: op1_08_in01 = reg_0008;
    41: op1_08_in01 = reg_0395;
    42: op1_08_in01 = reg_0216;
    43: op1_08_in01 = reg_0940;
    44: op1_08_in01 = reg_0132;
    45: op1_08_in01 = reg_0682;
    46: op1_08_in01 = reg_0500;
    47: op1_08_in01 = reg_0882;
    48: op1_08_in01 = imem00_in[55:52];
    50: op1_08_in01 = imem00_in[55:52];
    51: op1_08_in01 = reg_0705;
    52: op1_08_in01 = reg_0129;
    54: op1_08_in01 = reg_0868;
    55: op1_08_in01 = reg_0384;
    56: op1_08_in01 = imem00_in[127:124];
    57: op1_08_in01 = reg_0232;
    58: op1_08_in01 = reg_0007;
    59: op1_08_in01 = imem02_in[31:28];
    60: op1_08_in01 = imem04_in[71:68];
    61: op1_08_in01 = reg_0847;
    62: op1_08_in01 = reg_0935;
    63: op1_08_in01 = imem00_in[67:64];
    64: op1_08_in01 = imem00_in[71:68];
    72: op1_08_in01 = imem00_in[71:68];
    65: op1_08_in01 = reg_0304;
    66: op1_08_in01 = reg_0906;
    67: op1_08_in01 = reg_0109;
    68: op1_08_in01 = reg_0912;
    69: op1_08_in01 = imem07_in[23:20];
    70: op1_08_in01 = imem02_in[99:96];
    71: op1_08_in01 = reg_0240;
    73: op1_08_in01 = reg_0783;
    74: op1_08_in01 = reg_1051;
    75: op1_08_in01 = reg_0991;
    76: op1_08_in01 = reg_0965;
    78: op1_08_in01 = imem07_in[91:88];
    79: op1_08_in01 = imem00_in[47:44];
    80: op1_08_in01 = imem02_in[119:116];
    81: op1_08_in01 = reg_0239;
    82: op1_08_in01 = reg_0750;
    83: op1_08_in01 = imem00_in[23:20];
    84: op1_08_in01 = imem05_in[51:48];
    85: op1_08_in01 = reg_0821;
    86: op1_08_in01 = reg_0357;
    87: op1_08_in01 = reg_0369;
    88: op1_08_in01 = imem00_in[11:8];
    89: op1_08_in01 = imem06_in[23:20];
    90: op1_08_in01 = reg_0615;
    91: op1_08_in01 = reg_1056;
    92: op1_08_in01 = reg_0101;
    93: op1_08_in01 = reg_0944;
    94: op1_08_in01 = reg_0444;
    95: op1_08_in01 = reg_0015;
    96: op1_08_in01 = imem06_in[39:36];
    97: op1_08_in01 = reg_0060;
    default: op1_08_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_08_inv01 = 1;
    9: op1_08_inv01 = 1;
    10: op1_08_inv01 = 1;
    13: op1_08_inv01 = 1;
    15: op1_08_inv01 = 1;
    16: op1_08_inv01 = 1;
    3: op1_08_inv01 = 1;
    22: op1_08_inv01 = 1;
    25: op1_08_inv01 = 1;
    26: op1_08_inv01 = 1;
    2: op1_08_inv01 = 1;
    28: op1_08_inv01 = 1;
    30: op1_08_inv01 = 1;
    32: op1_08_inv01 = 1;
    36: op1_08_inv01 = 1;
    38: op1_08_inv01 = 1;
    40: op1_08_inv01 = 1;
    42: op1_08_inv01 = 1;
    45: op1_08_inv01 = 1;
    46: op1_08_inv01 = 1;
    47: op1_08_inv01 = 1;
    48: op1_08_inv01 = 1;
    51: op1_08_inv01 = 1;
    53: op1_08_inv01 = 1;
    54: op1_08_inv01 = 1;
    55: op1_08_inv01 = 1;
    57: op1_08_inv01 = 1;
    59: op1_08_inv01 = 1;
    61: op1_08_inv01 = 1;
    65: op1_08_inv01 = 1;
    66: op1_08_inv01 = 1;
    67: op1_08_inv01 = 1;
    68: op1_08_inv01 = 1;
    69: op1_08_inv01 = 1;
    73: op1_08_inv01 = 1;
    75: op1_08_inv01 = 1;
    77: op1_08_inv01 = 1;
    79: op1_08_inv01 = 1;
    81: op1_08_inv01 = 1;
    82: op1_08_inv01 = 1;
    83: op1_08_inv01 = 1;
    84: op1_08_inv01 = 1;
    86: op1_08_inv01 = 1;
    87: op1_08_inv01 = 1;
    89: op1_08_inv01 = 1;
    91: op1_08_inv01 = 1;
    95: op1_08_inv01 = 1;
    96: op1_08_inv01 = 1;
    97: op1_08_inv01 = 1;
    default: op1_08_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in02 = imem05_in[39:36];
    6: op1_08_in02 = reg_0370;
    7: op1_08_in02 = imem07_in[67:64];
    8: op1_08_in02 = reg_0242;
    9: op1_08_in02 = imem05_in[63:60];
    10: op1_08_in02 = reg_0597;
    11: op1_08_in02 = reg_0266;
    12: op1_08_in02 = reg_0060;
    13: op1_08_in02 = imem00_in[39:36];
    21: op1_08_in02 = imem00_in[39:36];
    14: op1_08_in02 = reg_0508;
    15: op1_08_in02 = reg_0573;
    4: op1_08_in02 = imem07_in[55:52];
    16: op1_08_in02 = reg_0337;
    17: op1_08_in02 = imem00_in[83:80];
    18: op1_08_in02 = reg_0138;
    19: op1_08_in02 = imem00_in[127:124];
    20: op1_08_in02 = imem06_in[83:80];
    3: op1_08_in02 = imem07_in[107:104];
    22: op1_08_in02 = reg_0275;
    23: op1_08_in02 = imem05_in[71:68];
    84: op1_08_in02 = imem05_in[71:68];
    24: op1_08_in02 = reg_0068;
    25: op1_08_in02 = reg_0604;
    26: op1_08_in02 = reg_0103;
    27: op1_08_in02 = reg_1028;
    28: op1_08_in02 = imem00_in[71:68];
    29: op1_08_in02 = reg_0959;
    30: op1_08_in02 = reg_0005;
    31: op1_08_in02 = reg_0686;
    32: op1_08_in02 = reg_0576;
    33: op1_08_in02 = reg_0976;
    34: op1_08_in02 = imem07_in[27:24];
    35: op1_08_in02 = reg_0318;
    36: op1_08_in02 = reg_0126;
    37: op1_08_in02 = reg_0793;
    38: op1_08_in02 = reg_0640;
    39: op1_08_in02 = reg_0834;
    40: op1_08_in02 = imem07_in[3:0];
    41: op1_08_in02 = reg_0295;
    42: op1_08_in02 = reg_0740;
    43: op1_08_in02 = reg_0327;
    86: op1_08_in02 = reg_0327;
    44: op1_08_in02 = reg_0148;
    45: op1_08_in02 = reg_0670;
    46: op1_08_in02 = reg_0354;
    47: op1_08_in02 = imem05_in[31:28];
    48: op1_08_in02 = imem00_in[119:116];
    49: op1_08_in02 = reg_0101;
    50: op1_08_in02 = imem00_in[99:96];
    51: op1_08_in02 = reg_0715;
    52: op1_08_in02 = reg_0130;
    53: op1_08_in02 = imem07_in[47:44];
    54: op1_08_in02 = reg_0162;
    55: op1_08_in02 = reg_0352;
    56: op1_08_in02 = reg_0841;
    64: op1_08_in02 = reg_0841;
    57: op1_08_in02 = reg_1055;
    65: op1_08_in02 = reg_1055;
    58: op1_08_in02 = reg_0482;
    59: op1_08_in02 = imem02_in[75:72];
    60: op1_08_in02 = imem04_in[119:116];
    61: op1_08_in02 = reg_0923;
    62: op1_08_in02 = reg_0237;
    63: op1_08_in02 = imem00_in[87:84];
    66: op1_08_in02 = reg_0232;
    67: op1_08_in02 = reg_0110;
    68: op1_08_in02 = reg_0306;
    69: op1_08_in02 = imem07_in[51:48];
    70: op1_08_in02 = reg_0666;
    71: op1_08_in02 = reg_0278;
    72: op1_08_in02 = reg_0682;
    73: op1_08_in02 = reg_0643;
    74: op1_08_in02 = reg_0769;
    75: op1_08_in02 = reg_1001;
    76: op1_08_in02 = imem06_in[15:12];
    77: op1_08_in02 = reg_0259;
    78: op1_08_in02 = imem07_in[95:92];
    79: op1_08_in02 = imem00_in[63:60];
    80: op1_08_in02 = imem02_in[127:124];
    81: op1_08_in02 = reg_0040;
    82: op1_08_in02 = reg_0844;
    83: op1_08_in02 = imem00_in[35:32];
    85: op1_08_in02 = reg_0745;
    87: op1_08_in02 = reg_0022;
    88: op1_08_in02 = imem00_in[31:28];
    89: op1_08_in02 = imem06_in[39:36];
    90: op1_08_in02 = reg_0512;
    91: op1_08_in02 = reg_0904;
    92: op1_08_in02 = reg_0109;
    93: op1_08_in02 = reg_0954;
    94: op1_08_in02 = reg_0027;
    95: op1_08_in02 = reg_0809;
    96: op1_08_in02 = imem06_in[67:64];
    97: op1_08_in02 = reg_0982;
    default: op1_08_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_08_inv02 = 1;
    9: op1_08_inv02 = 1;
    11: op1_08_inv02 = 1;
    12: op1_08_inv02 = 1;
    14: op1_08_inv02 = 1;
    4: op1_08_inv02 = 1;
    17: op1_08_inv02 = 1;
    18: op1_08_inv02 = 1;
    19: op1_08_inv02 = 1;
    3: op1_08_inv02 = 1;
    22: op1_08_inv02 = 1;
    25: op1_08_inv02 = 1;
    26: op1_08_inv02 = 1;
    28: op1_08_inv02 = 1;
    29: op1_08_inv02 = 1;
    30: op1_08_inv02 = 1;
    31: op1_08_inv02 = 1;
    34: op1_08_inv02 = 1;
    36: op1_08_inv02 = 1;
    37: op1_08_inv02 = 1;
    38: op1_08_inv02 = 1;
    42: op1_08_inv02 = 1;
    45: op1_08_inv02 = 1;
    47: op1_08_inv02 = 1;
    51: op1_08_inv02 = 1;
    52: op1_08_inv02 = 1;
    56: op1_08_inv02 = 1;
    58: op1_08_inv02 = 1;
    63: op1_08_inv02 = 1;
    64: op1_08_inv02 = 1;
    67: op1_08_inv02 = 1;
    70: op1_08_inv02 = 1;
    72: op1_08_inv02 = 1;
    73: op1_08_inv02 = 1;
    74: op1_08_inv02 = 1;
    75: op1_08_inv02 = 1;
    77: op1_08_inv02 = 1;
    78: op1_08_inv02 = 1;
    79: op1_08_inv02 = 1;
    81: op1_08_inv02 = 1;
    83: op1_08_inv02 = 1;
    84: op1_08_inv02 = 1;
    85: op1_08_inv02 = 1;
    88: op1_08_inv02 = 1;
    90: op1_08_inv02 = 1;
    94: op1_08_inv02 = 1;
    95: op1_08_inv02 = 1;
    default: op1_08_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in03 = imem05_in[75:72];
    6: op1_08_in03 = reg_0322;
    7: op1_08_in03 = imem07_in[83:80];
    8: op1_08_in03 = reg_0228;
    9: op1_08_in03 = reg_0959;
    10: op1_08_in03 = reg_0595;
    11: op1_08_in03 = reg_0152;
    12: op1_08_in03 = reg_0073;
    13: op1_08_in03 = imem00_in[43:40];
    14: op1_08_in03 = reg_1039;
    15: op1_08_in03 = reg_0583;
    4: op1_08_in03 = imem07_in[87:84];
    16: op1_08_in03 = reg_0368;
    17: op1_08_in03 = imem00_in[111:108];
    18: op1_08_in03 = reg_0130;
    19: op1_08_in03 = reg_0682;
    20: op1_08_in03 = reg_0625;
    21: op1_08_in03 = imem00_in[75:72];
    3: op1_08_in03 = imem07_in[127:124];
    22: op1_08_in03 = reg_0896;
    23: op1_08_in03 = imem05_in[119:116];
    24: op1_08_in03 = reg_0296;
    25: op1_08_in03 = reg_0630;
    26: op1_08_in03 = reg_0120;
    27: op1_08_in03 = reg_1010;
    28: op1_08_in03 = imem00_in[103:100];
    63: op1_08_in03 = imem00_in[103:100];
    29: op1_08_in03 = reg_0968;
    30: op1_08_in03 = imem07_in[19:16];
    31: op1_08_in03 = reg_0674;
    32: op1_08_in03 = reg_0793;
    33: op1_08_in03 = reg_0994;
    34: op1_08_in03 = imem07_in[35:32];
    35: op1_08_in03 = reg_0516;
    36: op1_08_in03 = imem02_in[3:0];
    37: op1_08_in03 = reg_0795;
    38: op1_08_in03 = reg_0648;
    39: op1_08_in03 = reg_0821;
    40: op1_08_in03 = imem07_in[23:20];
    41: op1_08_in03 = reg_0388;
    42: op1_08_in03 = reg_0925;
    43: op1_08_in03 = reg_0874;
    44: op1_08_in03 = reg_0142;
    45: op1_08_in03 = reg_0690;
    46: op1_08_in03 = reg_0740;
    47: op1_08_in03 = imem05_in[51:48];
    48: op1_08_in03 = reg_0685;
    56: op1_08_in03 = reg_0685;
    49: op1_08_in03 = reg_0115;
    50: op1_08_in03 = reg_0697;
    51: op1_08_in03 = reg_0707;
    52: op1_08_in03 = reg_0140;
    53: op1_08_in03 = imem07_in[107:104];
    54: op1_08_in03 = reg_0167;
    55: op1_08_in03 = reg_0679;
    57: op1_08_in03 = reg_0512;
    58: op1_08_in03 = reg_0085;
    59: op1_08_in03 = imem02_in[111:108];
    60: op1_08_in03 = reg_1006;
    61: op1_08_in03 = reg_0369;
    62: op1_08_in03 = reg_0949;
    64: op1_08_in03 = reg_0768;
    65: op1_08_in03 = reg_1033;
    66: op1_08_in03 = reg_0832;
    67: op1_08_in03 = imem02_in[11:8];
    68: op1_08_in03 = reg_0507;
    69: op1_08_in03 = imem07_in[67:64];
    70: op1_08_in03 = reg_0260;
    71: op1_08_in03 = reg_0571;
    86: op1_08_in03 = reg_0571;
    72: op1_08_in03 = reg_0841;
    73: op1_08_in03 = reg_0039;
    74: op1_08_in03 = reg_0555;
    75: op1_08_in03 = imem04_in[51:48];
    76: op1_08_in03 = imem06_in[27:24];
    77: op1_08_in03 = reg_0675;
    78: op1_08_in03 = reg_0716;
    79: op1_08_in03 = imem00_in[91:88];
    80: op1_08_in03 = reg_0750;
    81: op1_08_in03 = reg_0377;
    82: op1_08_in03 = reg_0700;
    83: op1_08_in03 = imem00_in[55:52];
    84: op1_08_in03 = reg_1021;
    85: op1_08_in03 = reg_0110;
    87: op1_08_in03 = imem07_in[3:0];
    88: op1_08_in03 = imem00_in[123:120];
    89: op1_08_in03 = imem06_in[51:48];
    90: op1_08_in03 = reg_0116;
    91: op1_08_in03 = reg_0501;
    92: op1_08_in03 = imem02_in[31:28];
    93: op1_08_in03 = reg_0319;
    94: op1_08_in03 = reg_0824;
    95: op1_08_in03 = reg_0432;
    96: op1_08_in03 = imem06_in[83:80];
    97: op1_08_in03 = reg_0613;
    default: op1_08_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv03 = 1;
    10: op1_08_inv03 = 1;
    11: op1_08_inv03 = 1;
    14: op1_08_inv03 = 1;
    15: op1_08_inv03 = 1;
    17: op1_08_inv03 = 1;
    21: op1_08_inv03 = 1;
    22: op1_08_inv03 = 1;
    23: op1_08_inv03 = 1;
    24: op1_08_inv03 = 1;
    25: op1_08_inv03 = 1;
    27: op1_08_inv03 = 1;
    28: op1_08_inv03 = 1;
    31: op1_08_inv03 = 1;
    32: op1_08_inv03 = 1;
    33: op1_08_inv03 = 1;
    37: op1_08_inv03 = 1;
    38: op1_08_inv03 = 1;
    39: op1_08_inv03 = 1;
    40: op1_08_inv03 = 1;
    42: op1_08_inv03 = 1;
    43: op1_08_inv03 = 1;
    44: op1_08_inv03 = 1;
    46: op1_08_inv03 = 1;
    49: op1_08_inv03 = 1;
    52: op1_08_inv03 = 1;
    53: op1_08_inv03 = 1;
    54: op1_08_inv03 = 1;
    55: op1_08_inv03 = 1;
    56: op1_08_inv03 = 1;
    58: op1_08_inv03 = 1;
    63: op1_08_inv03 = 1;
    66: op1_08_inv03 = 1;
    68: op1_08_inv03 = 1;
    70: op1_08_inv03 = 1;
    71: op1_08_inv03 = 1;
    76: op1_08_inv03 = 1;
    77: op1_08_inv03 = 1;
    78: op1_08_inv03 = 1;
    80: op1_08_inv03 = 1;
    83: op1_08_inv03 = 1;
    86: op1_08_inv03 = 1;
    87: op1_08_inv03 = 1;
    89: op1_08_inv03 = 1;
    91: op1_08_inv03 = 1;
    93: op1_08_inv03 = 1;
    94: op1_08_inv03 = 1;
    95: op1_08_inv03 = 1;
    96: op1_08_inv03 = 1;
    default: op1_08_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in04 = imem05_in[91:88];
    6: op1_08_in04 = imem03_in[95:92];
    7: op1_08_in04 = imem07_in[119:116];
    8: op1_08_in04 = reg_0102;
    9: op1_08_in04 = reg_0956;
    10: op1_08_in04 = reg_0388;
    11: op1_08_in04 = reg_0153;
    12: op1_08_in04 = imem03_in[59:56];
    13: op1_08_in04 = imem00_in[71:68];
    14: op1_08_in04 = reg_0869;
    15: op1_08_in04 = reg_0592;
    4: op1_08_in04 = imem07_in[127:124];
    16: op1_08_in04 = reg_1029;
    41: op1_08_in04 = reg_1029;
    17: op1_08_in04 = reg_0697;
    18: op1_08_in04 = imem06_in[7:4];
    19: op1_08_in04 = reg_0696;
    20: op1_08_in04 = reg_0626;
    21: op1_08_in04 = imem00_in[99:96];
    3: op1_08_in04 = reg_0174;
    22: op1_08_in04 = reg_0832;
    23: op1_08_in04 = reg_0962;
    24: op1_08_in04 = reg_0072;
    25: op1_08_in04 = reg_0618;
    26: op1_08_in04 = reg_0112;
    66: op1_08_in04 = reg_0112;
    27: op1_08_in04 = reg_0803;
    28: op1_08_in04 = reg_0686;
    64: op1_08_in04 = reg_0686;
    29: op1_08_in04 = reg_0946;
    30: op1_08_in04 = imem07_in[27:24];
    31: op1_08_in04 = reg_0678;
    32: op1_08_in04 = reg_0040;
    33: op1_08_in04 = imem04_in[15:12];
    34: op1_08_in04 = imem07_in[39:36];
    35: op1_08_in04 = reg_0772;
    36: op1_08_in04 = imem02_in[55:52];
    37: op1_08_in04 = reg_0051;
    38: op1_08_in04 = reg_0638;
    85: op1_08_in04 = reg_0638;
    39: op1_08_in04 = reg_0826;
    84: op1_08_in04 = reg_0826;
    40: op1_08_in04 = imem07_in[107:104];
    42: op1_08_in04 = reg_0106;
    43: op1_08_in04 = reg_0793;
    44: op1_08_in04 = reg_0134;
    45: op1_08_in04 = reg_0688;
    46: op1_08_in04 = imem02_in[35:32];
    47: op1_08_in04 = imem05_in[79:76];
    48: op1_08_in04 = reg_0676;
    50: op1_08_in04 = reg_0676;
    49: op1_08_in04 = reg_0127;
    51: op1_08_in04 = reg_0706;
    52: op1_08_in04 = imem06_in[63:60];
    53: op1_08_in04 = reg_0716;
    54: op1_08_in04 = reg_0166;
    55: op1_08_in04 = reg_0328;
    56: op1_08_in04 = reg_0748;
    57: op1_08_in04 = reg_0116;
    58: op1_08_in04 = reg_0090;
    59: op1_08_in04 = imem02_in[115:112];
    60: op1_08_in04 = reg_0912;
    61: op1_08_in04 = reg_0807;
    62: op1_08_in04 = reg_0063;
    63: op1_08_in04 = reg_0682;
    65: op1_08_in04 = reg_0273;
    67: op1_08_in04 = imem02_in[15:12];
    68: op1_08_in04 = reg_0524;
    69: op1_08_in04 = imem07_in[87:84];
    70: op1_08_in04 = reg_0098;
    71: op1_08_in04 = reg_1008;
    72: op1_08_in04 = reg_0825;
    79: op1_08_in04 = reg_0825;
    73: op1_08_in04 = reg_0394;
    74: op1_08_in04 = reg_0115;
    75: op1_08_in04 = imem04_in[71:68];
    76: op1_08_in04 = imem06_in[55:52];
    77: op1_08_in04 = reg_0947;
    78: op1_08_in04 = reg_0713;
    80: op1_08_in04 = reg_0886;
    81: op1_08_in04 = reg_0779;
    82: op1_08_in04 = reg_0441;
    83: op1_08_in04 = imem00_in[83:80];
    86: op1_08_in04 = reg_0038;
    87: op1_08_in04 = imem07_in[15:12];
    88: op1_08_in04 = reg_0683;
    89: op1_08_in04 = imem06_in[115:112];
    90: op1_08_in04 = reg_0101;
    91: op1_08_in04 = reg_0522;
    92: op1_08_in04 = imem02_in[39:36];
    93: op1_08_in04 = reg_0448;
    94: op1_08_in04 = reg_0332;
    95: op1_08_in04 = reg_0065;
    96: op1_08_in04 = imem06_in[103:100];
    97: op1_08_in04 = reg_0978;
    default: op1_08_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv04 = 1;
    6: op1_08_inv04 = 1;
    7: op1_08_inv04 = 1;
    9: op1_08_inv04 = 1;
    10: op1_08_inv04 = 1;
    11: op1_08_inv04 = 1;
    15: op1_08_inv04 = 1;
    4: op1_08_inv04 = 1;
    19: op1_08_inv04 = 1;
    21: op1_08_inv04 = 1;
    24: op1_08_inv04 = 1;
    26: op1_08_inv04 = 1;
    28: op1_08_inv04 = 1;
    29: op1_08_inv04 = 1;
    33: op1_08_inv04 = 1;
    34: op1_08_inv04 = 1;
    36: op1_08_inv04 = 1;
    42: op1_08_inv04 = 1;
    45: op1_08_inv04 = 1;
    47: op1_08_inv04 = 1;
    49: op1_08_inv04 = 1;
    53: op1_08_inv04 = 1;
    55: op1_08_inv04 = 1;
    56: op1_08_inv04 = 1;
    57: op1_08_inv04 = 1;
    60: op1_08_inv04 = 1;
    63: op1_08_inv04 = 1;
    66: op1_08_inv04 = 1;
    69: op1_08_inv04 = 1;
    73: op1_08_inv04 = 1;
    77: op1_08_inv04 = 1;
    83: op1_08_inv04 = 1;
    84: op1_08_inv04 = 1;
    85: op1_08_inv04 = 1;
    88: op1_08_inv04 = 1;
    89: op1_08_inv04 = 1;
    90: op1_08_inv04 = 1;
    91: op1_08_inv04 = 1;
    92: op1_08_inv04 = 1;
    95: op1_08_inv04 = 1;
    default: op1_08_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in05 = imem05_in[95:92];
    6: op1_08_in05 = imem04_in[23:20];
    7: op1_08_in05 = reg_0717;
    8: op1_08_in05 = reg_0107;
    9: op1_08_in05 = reg_0964;
    10: op1_08_in05 = reg_0377;
    11: op1_08_in05 = reg_0140;
    12: op1_08_in05 = imem03_in[63:60];
    13: op1_08_in05 = reg_0698;
    19: op1_08_in05 = reg_0698;
    14: op1_08_in05 = reg_0830;
    15: op1_08_in05 = reg_0600;
    4: op1_08_in05 = reg_0446;
    16: op1_08_in05 = reg_0027;
    17: op1_08_in05 = reg_0694;
    18: op1_08_in05 = imem06_in[27:24];
    20: op1_08_in05 = reg_0611;
    21: op1_08_in05 = reg_0695;
    3: op1_08_in05 = reg_0167;
    22: op1_08_in05 = reg_0819;
    23: op1_08_in05 = reg_0954;
    24: op1_08_in05 = reg_0738;
    25: op1_08_in05 = reg_0612;
    26: op1_08_in05 = reg_0320;
    27: op1_08_in05 = imem07_in[11:8];
    28: op1_08_in05 = reg_0688;
    29: op1_08_in05 = reg_0256;
    39: op1_08_in05 = reg_0256;
    30: op1_08_in05 = imem07_in[31:28];
    87: op1_08_in05 = imem07_in[31:28];
    31: op1_08_in05 = reg_0668;
    32: op1_08_in05 = reg_0509;
    33: op1_08_in05 = imem04_in[43:40];
    97: op1_08_in05 = imem04_in[43:40];
    34: op1_08_in05 = imem07_in[87:84];
    35: op1_08_in05 = reg_0814;
    36: op1_08_in05 = imem02_in[119:116];
    37: op1_08_in05 = reg_0767;
    38: op1_08_in05 = reg_0636;
    40: op1_08_in05 = reg_0722;
    41: op1_08_in05 = reg_0332;
    42: op1_08_in05 = imem02_in[43:40];
    43: op1_08_in05 = reg_0543;
    44: op1_08_in05 = imem06_in[15:12];
    45: op1_08_in05 = reg_0687;
    48: op1_08_in05 = reg_0687;
    46: op1_08_in05 = imem02_in[111:108];
    47: op1_08_in05 = imem05_in[103:100];
    49: op1_08_in05 = reg_0110;
    50: op1_08_in05 = reg_0689;
    51: op1_08_in05 = reg_0421;
    52: op1_08_in05 = reg_0624;
    53: op1_08_in05 = reg_0704;
    55: op1_08_in05 = reg_0383;
    56: op1_08_in05 = reg_0842;
    64: op1_08_in05 = reg_0842;
    57: op1_08_in05 = reg_0109;
    58: op1_08_in05 = reg_0084;
    59: op1_08_in05 = reg_0515;
    60: op1_08_in05 = reg_0048;
    61: op1_08_in05 = reg_0513;
    62: op1_08_in05 = reg_0032;
    63: op1_08_in05 = reg_0748;
    65: op1_08_in05 = reg_0860;
    66: op1_08_in05 = reg_0860;
    67: op1_08_in05 = imem02_in[87:84];
    68: op1_08_in05 = reg_0815;
    69: op1_08_in05 = imem07_in[99:96];
    70: op1_08_in05 = reg_0887;
    71: op1_08_in05 = reg_0609;
    72: op1_08_in05 = reg_0686;
    73: op1_08_in05 = reg_0644;
    74: op1_08_in05 = imem02_in[63:60];
    75: op1_08_in05 = imem04_in[79:76];
    76: op1_08_in05 = imem06_in[83:80];
    77: op1_08_in05 = reg_0707;
    78: op1_08_in05 = reg_0428;
    79: op1_08_in05 = reg_0670;
    88: op1_08_in05 = reg_0670;
    80: op1_08_in05 = reg_0762;
    81: op1_08_in05 = reg_0376;
    82: op1_08_in05 = reg_0424;
    83: op1_08_in05 = imem00_in[87:84];
    84: op1_08_in05 = reg_0647;
    85: op1_08_in05 = reg_0844;
    86: op1_08_in05 = reg_0996;
    89: op1_08_in05 = reg_0715;
    90: op1_08_in05 = reg_0113;
    91: op1_08_in05 = reg_0496;
    92: op1_08_in05 = imem02_in[67:64];
    93: op1_08_in05 = reg_0137;
    94: op1_08_in05 = imem05_in[11:8];
    95: op1_08_in05 = reg_0627;
    96: op1_08_in05 = reg_0660;
    default: op1_08_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv05 = 1;
    9: op1_08_inv05 = 1;
    11: op1_08_inv05 = 1;
    13: op1_08_inv05 = 1;
    14: op1_08_inv05 = 1;
    4: op1_08_inv05 = 1;
    17: op1_08_inv05 = 1;
    19: op1_08_inv05 = 1;
    22: op1_08_inv05 = 1;
    23: op1_08_inv05 = 1;
    25: op1_08_inv05 = 1;
    27: op1_08_inv05 = 1;
    28: op1_08_inv05 = 1;
    29: op1_08_inv05 = 1;
    32: op1_08_inv05 = 1;
    33: op1_08_inv05 = 1;
    35: op1_08_inv05 = 1;
    36: op1_08_inv05 = 1;
    38: op1_08_inv05 = 1;
    39: op1_08_inv05 = 1;
    43: op1_08_inv05 = 1;
    45: op1_08_inv05 = 1;
    46: op1_08_inv05 = 1;
    47: op1_08_inv05 = 1;
    49: op1_08_inv05 = 1;
    51: op1_08_inv05 = 1;
    52: op1_08_inv05 = 1;
    53: op1_08_inv05 = 1;
    55: op1_08_inv05 = 1;
    59: op1_08_inv05 = 1;
    60: op1_08_inv05 = 1;
    61: op1_08_inv05 = 1;
    68: op1_08_inv05 = 1;
    71: op1_08_inv05 = 1;
    75: op1_08_inv05 = 1;
    76: op1_08_inv05 = 1;
    77: op1_08_inv05 = 1;
    80: op1_08_inv05 = 1;
    81: op1_08_inv05 = 1;
    85: op1_08_inv05 = 1;
    86: op1_08_inv05 = 1;
    88: op1_08_inv05 = 1;
    92: op1_08_inv05 = 1;
    93: op1_08_inv05 = 1;
    94: op1_08_inv05 = 1;
    95: op1_08_inv05 = 1;
    96: op1_08_inv05 = 1;
    default: op1_08_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in06 = imem05_in[115:112];
    6: op1_08_in06 = imem04_in[27:24];
    7: op1_08_in06 = reg_0724;
    8: op1_08_in06 = imem02_in[11:8];
    9: op1_08_in06 = reg_0942;
    10: op1_08_in06 = reg_0322;
    11: op1_08_in06 = imem06_in[51:48];
    12: op1_08_in06 = imem03_in[79:76];
    13: op1_08_in06 = reg_0691;
    14: op1_08_in06 = reg_1015;
    15: op1_08_in06 = reg_0578;
    4: op1_08_in06 = reg_0161;
    16: op1_08_in06 = reg_0753;
    17: op1_08_in06 = reg_0698;
    18: op1_08_in06 = imem06_in[71:68];
    19: op1_08_in06 = reg_0688;
    20: op1_08_in06 = reg_0618;
    21: op1_08_in06 = reg_0696;
    3: op1_08_in06 = reg_0164;
    22: op1_08_in06 = reg_0831;
    23: op1_08_in06 = reg_0950;
    24: op1_08_in06 = reg_0855;
    25: op1_08_in06 = reg_0356;
    26: op1_08_in06 = reg_0052;
    27: op1_08_in06 = imem07_in[27:24];
    28: op1_08_in06 = reg_0457;
    29: op1_08_in06 = reg_0139;
    30: op1_08_in06 = imem07_in[51:48];
    31: op1_08_in06 = reg_0675;
    32: op1_08_in06 = reg_0836;
    33: op1_08_in06 = imem04_in[99:96];
    34: op1_08_in06 = reg_0731;
    35: op1_08_in06 = reg_0084;
    36: op1_08_in06 = reg_0655;
    37: op1_08_in06 = reg_0985;
    38: op1_08_in06 = reg_0080;
    39: op1_08_in06 = reg_0827;
    66: op1_08_in06 = reg_0827;
    40: op1_08_in06 = reg_0721;
    41: op1_08_in06 = reg_0241;
    42: op1_08_in06 = imem02_in[63:60];
    43: op1_08_in06 = reg_0377;
    44: op1_08_in06 = imem06_in[43:40];
    45: op1_08_in06 = reg_0692;
    46: op1_08_in06 = imem02_in[115:112];
    47: op1_08_in06 = imem05_in[123:120];
    48: op1_08_in06 = reg_0463;
    49: op1_08_in06 = imem02_in[35:32];
    50: op1_08_in06 = reg_0690;
    51: op1_08_in06 = reg_0868;
    52: op1_08_in06 = reg_0486;
    53: op1_08_in06 = reg_0719;
    55: op1_08_in06 = imem00_in[15:12];
    56: op1_08_in06 = reg_0883;
    64: op1_08_in06 = reg_0883;
    57: op1_08_in06 = reg_0113;
    58: op1_08_in06 = reg_0016;
    59: op1_08_in06 = reg_0649;
    60: op1_08_in06 = reg_1057;
    61: op1_08_in06 = reg_0844;
    62: op1_08_in06 = reg_0774;
    63: op1_08_in06 = reg_0686;
    65: op1_08_in06 = reg_0101;
    67: op1_08_in06 = imem02_in[103:100];
    68: op1_08_in06 = reg_0893;
    69: op1_08_in06 = imem07_in[103:100];
    70: op1_08_in06 = reg_0636;
    71: op1_08_in06 = reg_0820;
    81: op1_08_in06 = reg_0820;
    72: op1_08_in06 = reg_0842;
    88: op1_08_in06 = reg_0842;
    73: op1_08_in06 = reg_0037;
    74: op1_08_in06 = imem02_in[79:76];
    75: op1_08_in06 = imem04_in[87:84];
    76: op1_08_in06 = reg_0344;
    77: op1_08_in06 = reg_0019;
    78: op1_08_in06 = reg_0641;
    79: op1_08_in06 = reg_0738;
    80: op1_08_in06 = reg_0039;
    82: op1_08_in06 = reg_0359;
    83: op1_08_in06 = reg_0001;
    84: op1_08_in06 = reg_0966;
    85: op1_08_in06 = reg_0536;
    86: op1_08_in06 = reg_1001;
    87: op1_08_in06 = imem07_in[39:36];
    89: op1_08_in06 = reg_0903;
    90: op1_08_in06 = reg_0110;
    91: op1_08_in06 = reg_0829;
    92: op1_08_in06 = imem02_in[107:104];
    93: op1_08_in06 = reg_0813;
    94: op1_08_in06 = imem05_in[23:20];
    95: op1_08_in06 = reg_0332;
    96: op1_08_in06 = reg_0391;
    97: op1_08_in06 = imem04_in[47:44];
    default: op1_08_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv06 = 1;
    7: op1_08_inv06 = 1;
    8: op1_08_inv06 = 1;
    11: op1_08_inv06 = 1;
    12: op1_08_inv06 = 1;
    16: op1_08_inv06 = 1;
    20: op1_08_inv06 = 1;
    21: op1_08_inv06 = 1;
    3: op1_08_inv06 = 1;
    22: op1_08_inv06 = 1;
    25: op1_08_inv06 = 1;
    26: op1_08_inv06 = 1;
    27: op1_08_inv06 = 1;
    28: op1_08_inv06 = 1;
    29: op1_08_inv06 = 1;
    30: op1_08_inv06 = 1;
    32: op1_08_inv06 = 1;
    36: op1_08_inv06 = 1;
    39: op1_08_inv06 = 1;
    42: op1_08_inv06 = 1;
    46: op1_08_inv06 = 1;
    48: op1_08_inv06 = 1;
    49: op1_08_inv06 = 1;
    50: op1_08_inv06 = 1;
    51: op1_08_inv06 = 1;
    55: op1_08_inv06 = 1;
    58: op1_08_inv06 = 1;
    60: op1_08_inv06 = 1;
    61: op1_08_inv06 = 1;
    63: op1_08_inv06 = 1;
    64: op1_08_inv06 = 1;
    66: op1_08_inv06 = 1;
    67: op1_08_inv06 = 1;
    68: op1_08_inv06 = 1;
    71: op1_08_inv06 = 1;
    72: op1_08_inv06 = 1;
    73: op1_08_inv06 = 1;
    75: op1_08_inv06 = 1;
    76: op1_08_inv06 = 1;
    78: op1_08_inv06 = 1;
    79: op1_08_inv06 = 1;
    81: op1_08_inv06 = 1;
    83: op1_08_inv06 = 1;
    85: op1_08_inv06 = 1;
    86: op1_08_inv06 = 1;
    87: op1_08_inv06 = 1;
    89: op1_08_inv06 = 1;
    90: op1_08_inv06 = 1;
    91: op1_08_inv06 = 1;
    92: op1_08_inv06 = 1;
    93: op1_08_inv06 = 1;
    95: op1_08_inv06 = 1;
    96: op1_08_inv06 = 1;
    default: op1_08_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in07 = reg_0488;
    62: op1_08_in07 = reg_0488;
    6: op1_08_in07 = imem04_in[43:40];
    7: op1_08_in07 = reg_0711;
    8: op1_08_in07 = imem02_in[83:80];
    9: op1_08_in07 = reg_0953;
    10: op1_08_in07 = reg_0309;
    11: op1_08_in07 = imem06_in[59:56];
    12: op1_08_in07 = imem03_in[99:96];
    13: op1_08_in07 = reg_0675;
    14: op1_08_in07 = reg_0871;
    15: op1_08_in07 = reg_0590;
    4: op1_08_in07 = reg_0162;
    16: op1_08_in07 = reg_1011;
    17: op1_08_in07 = reg_0677;
    18: op1_08_in07 = imem06_in[79:76];
    19: op1_08_in07 = reg_0451;
    20: op1_08_in07 = reg_0615;
    21: op1_08_in07 = reg_0686;
    3: op1_08_in07 = reg_0185;
    22: op1_08_in07 = reg_0489;
    23: op1_08_in07 = reg_0965;
    24: op1_08_in07 = reg_0044;
    95: op1_08_in07 = reg_0044;
    25: op1_08_in07 = reg_0405;
    26: op1_08_in07 = reg_0529;
    27: op1_08_in07 = imem07_in[39:36];
    28: op1_08_in07 = reg_0469;
    29: op1_08_in07 = reg_0141;
    30: op1_08_in07 = imem07_in[111:108];
    31: op1_08_in07 = reg_0476;
    32: op1_08_in07 = reg_0767;
    33: op1_08_in07 = imem04_in[123:120];
    34: op1_08_in07 = reg_0726;
    35: op1_08_in07 = reg_0291;
    36: op1_08_in07 = reg_0638;
    37: op1_08_in07 = reg_0987;
    38: op1_08_in07 = reg_0330;
    39: op1_08_in07 = reg_1046;
    40: op1_08_in07 = reg_0725;
    41: op1_08_in07 = reg_0029;
    42: op1_08_in07 = reg_0654;
    43: op1_08_in07 = reg_0807;
    44: op1_08_in07 = reg_0614;
    45: op1_08_in07 = reg_0464;
    46: op1_08_in07 = reg_0363;
    47: op1_08_in07 = reg_0963;
    48: op1_08_in07 = reg_0465;
    49: op1_08_in07 = imem02_in[43:40];
    50: op1_08_in07 = reg_0688;
    51: op1_08_in07 = reg_0640;
    52: op1_08_in07 = reg_0371;
    53: op1_08_in07 = reg_0720;
    55: op1_08_in07 = imem00_in[79:76];
    56: op1_08_in07 = reg_0674;
    57: op1_08_in07 = reg_0821;
    58: op1_08_in07 = reg_0884;
    59: op1_08_in07 = reg_0558;
    60: op1_08_in07 = reg_1020;
    61: op1_08_in07 = reg_0374;
    63: op1_08_in07 = reg_0687;
    64: op1_08_in07 = reg_0102;
    65: op1_08_in07 = reg_0109;
    66: op1_08_in07 = reg_0103;
    67: op1_08_in07 = imem02_in[127:124];
    68: op1_08_in07 = reg_0108;
    69: op1_08_in07 = imem07_in[119:116];
    70: op1_08_in07 = reg_0081;
    71: op1_08_in07 = reg_0985;
    72: op1_08_in07 = reg_0883;
    73: op1_08_in07 = reg_0335;
    74: op1_08_in07 = imem02_in[111:108];
    75: op1_08_in07 = reg_0937;
    76: op1_08_in07 = reg_1018;
    77: op1_08_in07 = reg_0145;
    78: op1_08_in07 = reg_0353;
    79: op1_08_in07 = reg_0356;
    88: op1_08_in07 = reg_0356;
    80: op1_08_in07 = reg_0368;
    81: op1_08_in07 = reg_0233;
    82: op1_08_in07 = reg_0052;
    83: op1_08_in07 = reg_0825;
    84: op1_08_in07 = reg_0107;
    85: op1_08_in07 = reg_0543;
    86: op1_08_in07 = imem04_in[71:68];
    87: op1_08_in07 = imem07_in[83:80];
    89: op1_08_in07 = reg_0250;
    90: op1_08_in07 = imem02_in[3:0];
    91: op1_08_in07 = reg_0830;
    92: op1_08_in07 = reg_0285;
    93: op1_08_in07 = reg_0892;
    94: op1_08_in07 = imem05_in[43:40];
    96: op1_08_in07 = reg_0025;
    97: op1_08_in07 = imem04_in[67:64];
    default: op1_08_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv07 = 1;
    7: op1_08_inv07 = 1;
    12: op1_08_inv07 = 1;
    13: op1_08_inv07 = 1;
    14: op1_08_inv07 = 1;
    15: op1_08_inv07 = 1;
    4: op1_08_inv07 = 1;
    17: op1_08_inv07 = 1;
    19: op1_08_inv07 = 1;
    22: op1_08_inv07 = 1;
    23: op1_08_inv07 = 1;
    26: op1_08_inv07 = 1;
    31: op1_08_inv07 = 1;
    32: op1_08_inv07 = 1;
    35: op1_08_inv07 = 1;
    36: op1_08_inv07 = 1;
    37: op1_08_inv07 = 1;
    38: op1_08_inv07 = 1;
    39: op1_08_inv07 = 1;
    40: op1_08_inv07 = 1;
    43: op1_08_inv07 = 1;
    44: op1_08_inv07 = 1;
    49: op1_08_inv07 = 1;
    50: op1_08_inv07 = 1;
    51: op1_08_inv07 = 1;
    52: op1_08_inv07 = 1;
    53: op1_08_inv07 = 1;
    55: op1_08_inv07 = 1;
    59: op1_08_inv07 = 1;
    61: op1_08_inv07 = 1;
    62: op1_08_inv07 = 1;
    64: op1_08_inv07 = 1;
    65: op1_08_inv07 = 1;
    66: op1_08_inv07 = 1;
    67: op1_08_inv07 = 1;
    69: op1_08_inv07 = 1;
    70: op1_08_inv07 = 1;
    73: op1_08_inv07 = 1;
    74: op1_08_inv07 = 1;
    80: op1_08_inv07 = 1;
    81: op1_08_inv07 = 1;
    83: op1_08_inv07 = 1;
    84: op1_08_inv07 = 1;
    85: op1_08_inv07 = 1;
    86: op1_08_inv07 = 1;
    91: op1_08_inv07 = 1;
    92: op1_08_inv07 = 1;
    96: op1_08_inv07 = 1;
    97: op1_08_inv07 = 1;
    default: op1_08_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in08 = reg_0489;
    6: op1_08_in08 = imem04_in[79:76];
    7: op1_08_in08 = reg_0707;
    8: op1_08_in08 = imem02_in[91:88];
    9: op1_08_in08 = reg_0268;
    10: op1_08_in08 = reg_0993;
    11: op1_08_in08 = imem06_in[67:64];
    12: op1_08_in08 = reg_0586;
    13: op1_08_in08 = reg_0680;
    64: op1_08_in08 = reg_0680;
    14: op1_08_in08 = reg_1038;
    15: op1_08_in08 = reg_0576;
    4: op1_08_in08 = reg_0163;
    16: op1_08_in08 = imem07_in[31:28];
    17: op1_08_in08 = reg_0678;
    18: op1_08_in08 = imem06_in[83:80];
    19: op1_08_in08 = reg_0472;
    20: op1_08_in08 = reg_0612;
    21: op1_08_in08 = reg_0679;
    3: op1_08_in08 = reg_0170;
    22: op1_08_in08 = reg_0497;
    23: op1_08_in08 = reg_0946;
    24: op1_08_in08 = imem05_in[15:12];
    25: op1_08_in08 = reg_0383;
    26: op1_08_in08 = reg_0328;
    27: op1_08_in08 = imem07_in[47:44];
    28: op1_08_in08 = reg_0481;
    29: op1_08_in08 = reg_0372;
    82: op1_08_in08 = reg_0372;
    30: op1_08_in08 = reg_0725;
    31: op1_08_in08 = reg_0458;
    32: op1_08_in08 = reg_0844;
    33: op1_08_in08 = reg_0301;
    34: op1_08_in08 = reg_0703;
    35: op1_08_in08 = imem03_in[55:52];
    36: op1_08_in08 = reg_0225;
    37: op1_08_in08 = reg_0996;
    38: op1_08_in08 = reg_0335;
    39: op1_08_in08 = reg_0254;
    40: op1_08_in08 = reg_0724;
    41: op1_08_in08 = imem07_in[15:12];
    42: op1_08_in08 = reg_0656;
    43: op1_08_in08 = reg_0982;
    44: op1_08_in08 = reg_0613;
    45: op1_08_in08 = reg_0187;
    46: op1_08_in08 = reg_0653;
    67: op1_08_in08 = reg_0653;
    47: op1_08_in08 = reg_0955;
    48: op1_08_in08 = reg_0464;
    49: op1_08_in08 = imem02_in[71:68];
    50: op1_08_in08 = reg_0669;
    51: op1_08_in08 = reg_0838;
    52: op1_08_in08 = reg_0556;
    53: op1_08_in08 = reg_0726;
    55: op1_08_in08 = imem00_in[99:96];
    56: op1_08_in08 = reg_0663;
    57: op1_08_in08 = imem02_in[15:12];
    58: op1_08_in08 = imem03_in[3:0];
    59: op1_08_in08 = reg_0424;
    60: op1_08_in08 = reg_0888;
    61: op1_08_in08 = reg_0998;
    62: op1_08_in08 = reg_0757;
    63: op1_08_in08 = reg_0465;
    65: op1_08_in08 = imem02_in[35:32];
    66: op1_08_in08 = imem02_in[11:8];
    90: op1_08_in08 = imem02_in[11:8];
    68: op1_08_in08 = reg_0070;
    69: op1_08_in08 = reg_0716;
    70: op1_08_in08 = reg_0359;
    85: op1_08_in08 = reg_0359;
    71: op1_08_in08 = reg_0979;
    72: op1_08_in08 = reg_0356;
    73: op1_08_in08 = reg_0516;
    74: op1_08_in08 = reg_0666;
    75: op1_08_in08 = reg_0932;
    76: op1_08_in08 = reg_0384;
    77: op1_08_in08 = reg_0144;
    78: op1_08_in08 = reg_0175;
    79: op1_08_in08 = reg_0674;
    80: op1_08_in08 = reg_0818;
    81: op1_08_in08 = imem04_in[3:0];
    83: op1_08_in08 = reg_0900;
    84: op1_08_in08 = reg_1015;
    86: op1_08_in08 = imem04_in[87:84];
    87: op1_08_in08 = imem07_in[95:92];
    88: op1_08_in08 = reg_0450;
    89: op1_08_in08 = reg_0422;
    91: op1_08_in08 = reg_1040;
    92: op1_08_in08 = reg_0639;
    93: op1_08_in08 = reg_0964;
    94: op1_08_in08 = imem05_in[55:52];
    95: op1_08_in08 = imem05_in[7:4];
    96: op1_08_in08 = reg_0021;
    97: op1_08_in08 = imem04_in[111:108];
    default: op1_08_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv08 = 1;
    6: op1_08_inv08 = 1;
    7: op1_08_inv08 = 1;
    9: op1_08_inv08 = 1;
    11: op1_08_inv08 = 1;
    12: op1_08_inv08 = 1;
    15: op1_08_inv08 = 1;
    16: op1_08_inv08 = 1;
    17: op1_08_inv08 = 1;
    18: op1_08_inv08 = 1;
    19: op1_08_inv08 = 1;
    21: op1_08_inv08 = 1;
    3: op1_08_inv08 = 1;
    22: op1_08_inv08 = 1;
    26: op1_08_inv08 = 1;
    28: op1_08_inv08 = 1;
    29: op1_08_inv08 = 1;
    34: op1_08_inv08 = 1;
    36: op1_08_inv08 = 1;
    37: op1_08_inv08 = 1;
    38: op1_08_inv08 = 1;
    39: op1_08_inv08 = 1;
    40: op1_08_inv08 = 1;
    42: op1_08_inv08 = 1;
    43: op1_08_inv08 = 1;
    45: op1_08_inv08 = 1;
    46: op1_08_inv08 = 1;
    47: op1_08_inv08 = 1;
    49: op1_08_inv08 = 1;
    50: op1_08_inv08 = 1;
    51: op1_08_inv08 = 1;
    53: op1_08_inv08 = 1;
    55: op1_08_inv08 = 1;
    58: op1_08_inv08 = 1;
    60: op1_08_inv08 = 1;
    63: op1_08_inv08 = 1;
    66: op1_08_inv08 = 1;
    69: op1_08_inv08 = 1;
    71: op1_08_inv08 = 1;
    72: op1_08_inv08 = 1;
    74: op1_08_inv08 = 1;
    75: op1_08_inv08 = 1;
    76: op1_08_inv08 = 1;
    77: op1_08_inv08 = 1;
    80: op1_08_inv08 = 1;
    81: op1_08_inv08 = 1;
    83: op1_08_inv08 = 1;
    87: op1_08_inv08 = 1;
    91: op1_08_inv08 = 1;
    94: op1_08_inv08 = 1;
    95: op1_08_inv08 = 1;
    97: op1_08_inv08 = 1;
    default: op1_08_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in09 = reg_0215;
    6: op1_08_in09 = imem04_in[107:104];
    7: op1_08_in09 = reg_0700;
    8: op1_08_in09 = imem02_in[115:112];
    9: op1_08_in09 = reg_0269;
    10: op1_08_in09 = reg_0986;
    11: op1_08_in09 = imem06_in[107:104];
    18: op1_08_in09 = imem06_in[107:104];
    12: op1_08_in09 = reg_0572;
    13: op1_08_in09 = reg_0455;
    14: op1_08_in09 = reg_0105;
    15: op1_08_in09 = reg_0360;
    16: op1_08_in09 = reg_0722;
    17: op1_08_in09 = reg_0699;
    19: op1_08_in09 = reg_0480;
    28: op1_08_in09 = reg_0480;
    20: op1_08_in09 = reg_0349;
    21: op1_08_in09 = reg_0675;
    3: op1_08_in09 = reg_0173;
    22: op1_08_in09 = reg_0136;
    23: op1_08_in09 = reg_0953;
    24: op1_08_in09 = imem05_in[67:64];
    25: op1_08_in09 = reg_0404;
    26: op1_08_in09 = reg_0657;
    27: op1_08_in09 = imem07_in[71:68];
    29: op1_08_in09 = reg_0915;
    30: op1_08_in09 = reg_0701;
    31: op1_08_in09 = reg_0187;
    32: op1_08_in09 = reg_0374;
    33: op1_08_in09 = reg_0265;
    34: op1_08_in09 = reg_0712;
    35: op1_08_in09 = imem03_in[107:104];
    36: op1_08_in09 = reg_0886;
    37: op1_08_in09 = imem04_in[63:60];
    38: op1_08_in09 = reg_0083;
    39: op1_08_in09 = reg_0489;
    40: op1_08_in09 = reg_0708;
    41: op1_08_in09 = imem07_in[43:40];
    42: op1_08_in09 = reg_0643;
    43: op1_08_in09 = reg_0995;
    44: op1_08_in09 = reg_0883;
    45: op1_08_in09 = reg_0194;
    46: op1_08_in09 = reg_0341;
    47: op1_08_in09 = reg_0964;
    48: op1_08_in09 = reg_0473;
    49: op1_08_in09 = imem02_in[107:104];
    50: op1_08_in09 = reg_0450;
    63: op1_08_in09 = reg_0450;
    51: op1_08_in09 = reg_0180;
    52: op1_08_in09 = reg_0632;
    53: op1_08_in09 = reg_0714;
    55: op1_08_in09 = reg_0457;
    56: op1_08_in09 = reg_0469;
    57: op1_08_in09 = imem02_in[47:44];
    58: op1_08_in09 = imem03_in[51:48];
    59: op1_08_in09 = reg_0039;
    60: op1_08_in09 = reg_0050;
    61: op1_08_in09 = reg_0974;
    62: op1_08_in09 = reg_0023;
    64: op1_08_in09 = reg_0687;
    65: op1_08_in09 = imem02_in[59:56];
    66: op1_08_in09 = imem02_in[99:96];
    67: op1_08_in09 = reg_0290;
    68: op1_08_in09 = reg_0774;
    69: op1_08_in09 = reg_0717;
    70: op1_08_in09 = reg_0389;
    71: op1_08_in09 = reg_0984;
    72: op1_08_in09 = reg_0828;
    73: op1_08_in09 = reg_0772;
    74: op1_08_in09 = reg_0095;
    75: op1_08_in09 = reg_0313;
    76: op1_08_in09 = reg_0534;
    77: op1_08_in09 = imem06_in[47:44];
    78: op1_08_in09 = reg_0167;
    79: op1_08_in09 = reg_0668;
    80: op1_08_in09 = reg_0347;
    81: op1_08_in09 = imem04_in[47:44];
    82: op1_08_in09 = reg_0037;
    83: op1_08_in09 = reg_0356;
    84: op1_08_in09 = reg_0736;
    85: op1_08_in09 = reg_0052;
    86: op1_08_in09 = imem04_in[119:116];
    87: op1_08_in09 = imem07_in[111:108];
    88: op1_08_in09 = reg_0461;
    89: op1_08_in09 = reg_0744;
    90: op1_08_in09 = imem02_in[35:32];
    91: op1_08_in09 = reg_0737;
    92: op1_08_in09 = reg_0087;
    93: op1_08_in09 = reg_0257;
    94: op1_08_in09 = imem05_in[83:80];
    95: op1_08_in09 = imem05_in[51:48];
    96: op1_08_in09 = reg_0338;
    97: op1_08_in09 = reg_0147;
    default: op1_08_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_08_inv09 = 1;
    9: op1_08_inv09 = 1;
    10: op1_08_inv09 = 1;
    13: op1_08_inv09 = 1;
    14: op1_08_inv09 = 1;
    15: op1_08_inv09 = 1;
    17: op1_08_inv09 = 1;
    18: op1_08_inv09 = 1;
    19: op1_08_inv09 = 1;
    3: op1_08_inv09 = 1;
    23: op1_08_inv09 = 1;
    24: op1_08_inv09 = 1;
    25: op1_08_inv09 = 1;
    26: op1_08_inv09 = 1;
    29: op1_08_inv09 = 1;
    31: op1_08_inv09 = 1;
    33: op1_08_inv09 = 1;
    36: op1_08_inv09 = 1;
    37: op1_08_inv09 = 1;
    39: op1_08_inv09 = 1;
    40: op1_08_inv09 = 1;
    42: op1_08_inv09 = 1;
    43: op1_08_inv09 = 1;
    44: op1_08_inv09 = 1;
    45: op1_08_inv09 = 1;
    46: op1_08_inv09 = 1;
    48: op1_08_inv09 = 1;
    53: op1_08_inv09 = 1;
    57: op1_08_inv09 = 1;
    60: op1_08_inv09 = 1;
    61: op1_08_inv09 = 1;
    62: op1_08_inv09 = 1;
    66: op1_08_inv09 = 1;
    68: op1_08_inv09 = 1;
    69: op1_08_inv09 = 1;
    74: op1_08_inv09 = 1;
    75: op1_08_inv09 = 1;
    76: op1_08_inv09 = 1;
    77: op1_08_inv09 = 1;
    82: op1_08_inv09 = 1;
    83: op1_08_inv09 = 1;
    85: op1_08_inv09 = 1;
    88: op1_08_inv09 = 1;
    90: op1_08_inv09 = 1;
    91: op1_08_inv09 = 1;
    92: op1_08_inv09 = 1;
    97: op1_08_inv09 = 1;
    default: op1_08_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in10 = reg_0261;
    6: op1_08_in10 = imem04_in[127:124];
    7: op1_08_in10 = reg_0429;
    8: op1_08_in10 = reg_0642;
    9: op1_08_in10 = reg_0244;
    10: op1_08_in10 = reg_0980;
    11: op1_08_in10 = reg_0614;
    12: op1_08_in10 = reg_0594;
    13: op1_08_in10 = reg_0470;
    19: op1_08_in10 = reg_0470;
    14: op1_08_in10 = reg_0111;
    15: op1_08_in10 = reg_0362;
    16: op1_08_in10 = reg_0730;
    17: op1_08_in10 = reg_0463;
    18: op1_08_in10 = reg_0619;
    20: op1_08_in10 = reg_0392;
    21: op1_08_in10 = reg_0680;
    79: op1_08_in10 = reg_0680;
    22: op1_08_in10 = reg_0151;
    23: op1_08_in10 = reg_0826;
    24: op1_08_in10 = imem05_in[71:68];
    25: op1_08_in10 = reg_0026;
    26: op1_08_in10 = reg_0651;
    27: op1_08_in10 = imem07_in[115:112];
    28: op1_08_in10 = reg_0214;
    55: op1_08_in10 = reg_0214;
    29: op1_08_in10 = reg_0371;
    30: op1_08_in10 = reg_0424;
    31: op1_08_in10 = reg_0212;
    32: op1_08_in10 = reg_0234;
    33: op1_08_in10 = reg_1009;
    34: op1_08_in10 = reg_0709;
    35: op1_08_in10 = imem03_in[119:116];
    36: op1_08_in10 = reg_0482;
    37: op1_08_in10 = reg_1006;
    38: op1_08_in10 = reg_0761;
    39: op1_08_in10 = reg_0145;
    40: op1_08_in10 = reg_0425;
    41: op1_08_in10 = imem07_in[79:76];
    42: op1_08_in10 = reg_0039;
    43: op1_08_in10 = reg_1001;
    44: op1_08_in10 = reg_0020;
    45: op1_08_in10 = reg_0213;
    46: op1_08_in10 = reg_0515;
    47: op1_08_in10 = reg_0835;
    48: op1_08_in10 = reg_0458;
    49: op1_08_in10 = imem02_in[111:108];
    50: op1_08_in10 = reg_0451;
    51: op1_08_in10 = reg_0172;
    52: op1_08_in10 = reg_0612;
    53: op1_08_in10 = reg_0708;
    56: op1_08_in10 = reg_0475;
    57: op1_08_in10 = imem02_in[63:60];
    58: op1_08_in10 = imem03_in[59:56];
    59: op1_08_in10 = reg_0664;
    60: op1_08_in10 = reg_0537;
    61: op1_08_in10 = imem04_in[87:84];
    62: op1_08_in10 = reg_0819;
    63: op1_08_in10 = reg_0481;
    64: op1_08_in10 = reg_0749;
    65: op1_08_in10 = imem02_in[103:100];
    66: op1_08_in10 = reg_0759;
    67: op1_08_in10 = reg_0873;
    68: op1_08_in10 = reg_0435;
    69: op1_08_in10 = reg_0724;
    70: op1_08_in10 = reg_0335;
    82: op1_08_in10 = reg_0335;
    71: op1_08_in10 = imem04_in[31:28];
    72: op1_08_in10 = reg_0687;
    73: op1_08_in10 = reg_0083;
    74: op1_08_in10 = reg_0645;
    75: op1_08_in10 = reg_0524;
    76: op1_08_in10 = reg_0804;
    77: op1_08_in10 = imem06_in[79:76];
    78: op1_08_in10 = reg_0183;
    80: op1_08_in10 = reg_0776;
    81: op1_08_in10 = imem04_in[59:56];
    83: op1_08_in10 = reg_0674;
    84: op1_08_in10 = reg_0795;
    85: op1_08_in10 = reg_0331;
    86: op1_08_in10 = reg_0942;
    97: op1_08_in10 = reg_0942;
    87: op1_08_in10 = imem07_in[123:120];
    88: op1_08_in10 = reg_0469;
    89: op1_08_in10 = reg_0419;
    90: op1_08_in10 = imem02_in[39:36];
    91: op1_08_in10 = reg_0616;
    92: op1_08_in10 = reg_0650;
    93: op1_08_in10 = reg_0970;
    94: op1_08_in10 = imem05_in[103:100];
    95: op1_08_in10 = imem05_in[55:52];
    96: op1_08_in10 = reg_0735;
    default: op1_08_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_08_inv10 = 1;
    13: op1_08_inv10 = 1;
    14: op1_08_inv10 = 1;
    15: op1_08_inv10 = 1;
    17: op1_08_inv10 = 1;
    18: op1_08_inv10 = 1;
    20: op1_08_inv10 = 1;
    21: op1_08_inv10 = 1;
    22: op1_08_inv10 = 1;
    25: op1_08_inv10 = 1;
    26: op1_08_inv10 = 1;
    28: op1_08_inv10 = 1;
    29: op1_08_inv10 = 1;
    31: op1_08_inv10 = 1;
    32: op1_08_inv10 = 1;
    33: op1_08_inv10 = 1;
    34: op1_08_inv10 = 1;
    36: op1_08_inv10 = 1;
    37: op1_08_inv10 = 1;
    39: op1_08_inv10 = 1;
    41: op1_08_inv10 = 1;
    42: op1_08_inv10 = 1;
    43: op1_08_inv10 = 1;
    45: op1_08_inv10 = 1;
    47: op1_08_inv10 = 1;
    53: op1_08_inv10 = 1;
    55: op1_08_inv10 = 1;
    56: op1_08_inv10 = 1;
    60: op1_08_inv10 = 1;
    66: op1_08_inv10 = 1;
    67: op1_08_inv10 = 1;
    70: op1_08_inv10 = 1;
    71: op1_08_inv10 = 1;
    72: op1_08_inv10 = 1;
    74: op1_08_inv10 = 1;
    78: op1_08_inv10 = 1;
    80: op1_08_inv10 = 1;
    83: op1_08_inv10 = 1;
    86: op1_08_inv10 = 1;
    87: op1_08_inv10 = 1;
    90: op1_08_inv10 = 1;
    93: op1_08_inv10 = 1;
    96: op1_08_inv10 = 1;
    97: op1_08_inv10 = 1;
    default: op1_08_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in11 = reg_0147;
    6: op1_08_in11 = reg_0545;
    7: op1_08_in11 = reg_0426;
    8: op1_08_in11 = reg_0645;
    9: op1_08_in11 = reg_0272;
    10: op1_08_in11 = reg_0978;
    11: op1_08_in11 = reg_0624;
    12: op1_08_in11 = reg_0593;
    13: op1_08_in11 = reg_0474;
    14: op1_08_in11 = reg_0118;
    15: op1_08_in11 = reg_0373;
    16: op1_08_in11 = reg_0705;
    17: op1_08_in11 = reg_0455;
    50: op1_08_in11 = reg_0455;
    18: op1_08_in11 = reg_0633;
    19: op1_08_in11 = reg_0471;
    20: op1_08_in11 = reg_0405;
    86: op1_08_in11 = reg_0405;
    21: op1_08_in11 = reg_0687;
    22: op1_08_in11 = reg_0154;
    23: op1_08_in11 = reg_0900;
    24: op1_08_in11 = reg_0944;
    25: op1_08_in11 = reg_0808;
    26: op1_08_in11 = reg_0643;
    27: op1_08_in11 = reg_0716;
    28: op1_08_in11 = imem01_in[3:0];
    29: op1_08_in11 = reg_0554;
    30: op1_08_in11 = reg_0447;
    31: op1_08_in11 = imem01_in[15:12];
    32: op1_08_in11 = reg_0822;
    33: op1_08_in11 = reg_0306;
    34: op1_08_in11 = reg_0715;
    35: op1_08_in11 = imem03_in[123:120];
    36: op1_08_in11 = reg_0776;
    73: op1_08_in11 = reg_0776;
    37: op1_08_in11 = reg_0530;
    38: op1_08_in11 = reg_0872;
    39: op1_08_in11 = reg_0136;
    40: op1_08_in11 = reg_0424;
    41: op1_08_in11 = imem07_in[123:120];
    42: op1_08_in11 = reg_0096;
    43: op1_08_in11 = reg_0999;
    44: op1_08_in11 = reg_0754;
    45: op1_08_in11 = reg_0202;
    56: op1_08_in11 = reg_0202;
    46: op1_08_in11 = reg_0639;
    47: op1_08_in11 = reg_0256;
    48: op1_08_in11 = reg_0191;
    49: op1_08_in11 = reg_0355;
    92: op1_08_in11 = reg_0355;
    51: op1_08_in11 = reg_0159;
    52: op1_08_in11 = reg_0385;
    53: op1_08_in11 = reg_0707;
    55: op1_08_in11 = reg_0209;
    57: op1_08_in11 = imem02_in[67:64];
    58: op1_08_in11 = imem03_in[103:100];
    59: op1_08_in11 = reg_0368;
    60: op1_08_in11 = reg_0752;
    61: op1_08_in11 = reg_0912;
    62: op1_08_in11 = reg_0438;
    63: op1_08_in11 = reg_0470;
    64: op1_08_in11 = reg_0472;
    65: op1_08_in11 = reg_0341;
    66: op1_08_in11 = reg_0741;
    67: op1_08_in11 = reg_0914;
    68: op1_08_in11 = reg_0942;
    69: op1_08_in11 = reg_0709;
    70: op1_08_in11 = reg_0758;
    71: op1_08_in11 = imem04_in[39:36];
    72: op1_08_in11 = reg_0749;
    79: op1_08_in11 = reg_0749;
    74: op1_08_in11 = reg_0394;
    75: op1_08_in11 = reg_0076;
    76: op1_08_in11 = reg_0921;
    77: op1_08_in11 = imem06_in[115:112];
    78: op1_08_in11 = reg_0168;
    80: op1_08_in11 = reg_0090;
    81: op1_08_in11 = imem04_in[111:108];
    82: op1_08_in11 = reg_0077;
    83: op1_08_in11 = reg_0828;
    84: op1_08_in11 = reg_0951;
    85: op1_08_in11 = reg_0818;
    87: op1_08_in11 = reg_0567;
    88: op1_08_in11 = reg_0475;
    89: op1_08_in11 = reg_0181;
    90: op1_08_in11 = reg_0285;
    91: op1_08_in11 = reg_0615;
    93: op1_08_in11 = reg_0135;
    94: op1_08_in11 = imem05_in[107:104];
    95: op1_08_in11 = reg_0866;
    96: op1_08_in11 = reg_0384;
    97: op1_08_in11 = reg_0430;
    default: op1_08_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv11 = 1;
    10: op1_08_inv11 = 1;
    11: op1_08_inv11 = 1;
    12: op1_08_inv11 = 1;
    13: op1_08_inv11 = 1;
    14: op1_08_inv11 = 1;
    15: op1_08_inv11 = 1;
    16: op1_08_inv11 = 1;
    17: op1_08_inv11 = 1;
    20: op1_08_inv11 = 1;
    21: op1_08_inv11 = 1;
    22: op1_08_inv11 = 1;
    23: op1_08_inv11 = 1;
    24: op1_08_inv11 = 1;
    25: op1_08_inv11 = 1;
    28: op1_08_inv11 = 1;
    30: op1_08_inv11 = 1;
    31: op1_08_inv11 = 1;
    34: op1_08_inv11 = 1;
    36: op1_08_inv11 = 1;
    38: op1_08_inv11 = 1;
    45: op1_08_inv11 = 1;
    47: op1_08_inv11 = 1;
    48: op1_08_inv11 = 1;
    51: op1_08_inv11 = 1;
    52: op1_08_inv11 = 1;
    53: op1_08_inv11 = 1;
    55: op1_08_inv11 = 1;
    59: op1_08_inv11 = 1;
    61: op1_08_inv11 = 1;
    64: op1_08_inv11 = 1;
    66: op1_08_inv11 = 1;
    67: op1_08_inv11 = 1;
    70: op1_08_inv11 = 1;
    77: op1_08_inv11 = 1;
    79: op1_08_inv11 = 1;
    80: op1_08_inv11 = 1;
    81: op1_08_inv11 = 1;
    82: op1_08_inv11 = 1;
    83: op1_08_inv11 = 1;
    84: op1_08_inv11 = 1;
    85: op1_08_inv11 = 1;
    86: op1_08_inv11 = 1;
    90: op1_08_inv11 = 1;
    92: op1_08_inv11 = 1;
    95: op1_08_inv11 = 1;
    96: op1_08_inv11 = 1;
    97: op1_08_inv11 = 1;
    default: op1_08_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in12 = reg_0148;
    6: op1_08_in12 = reg_0536;
    7: op1_08_in12 = reg_0172;
    8: op1_08_in12 = reg_0665;
    9: op1_08_in12 = reg_0261;
    10: op1_08_in12 = reg_0981;
    43: op1_08_in12 = reg_0981;
    11: op1_08_in12 = reg_0577;
    12: op1_08_in12 = reg_0311;
    13: op1_08_in12 = reg_0187;
    14: op1_08_in12 = reg_0112;
    15: op1_08_in12 = reg_0396;
    16: op1_08_in12 = reg_0701;
    53: op1_08_in12 = reg_0701;
    17: op1_08_in12 = reg_0461;
    50: op1_08_in12 = reg_0461;
    18: op1_08_in12 = reg_0623;
    19: op1_08_in12 = reg_0191;
    20: op1_08_in12 = reg_0386;
    21: op1_08_in12 = reg_0454;
    22: op1_08_in12 = imem06_in[3:0];
    23: op1_08_in12 = reg_0256;
    24: op1_08_in12 = reg_0955;
    25: op1_08_in12 = reg_0752;
    26: op1_08_in12 = reg_0652;
    46: op1_08_in12 = reg_0652;
    27: op1_08_in12 = reg_0710;
    28: op1_08_in12 = imem01_in[27:24];
    29: op1_08_in12 = reg_0610;
    30: op1_08_in12 = reg_0434;
    31: op1_08_in12 = imem01_in[23:20];
    32: op1_08_in12 = reg_0996;
    33: op1_08_in12 = reg_0539;
    34: op1_08_in12 = reg_0436;
    35: op1_08_in12 = reg_0535;
    36: op1_08_in12 = imem03_in[23:20];
    37: op1_08_in12 = reg_0778;
    38: op1_08_in12 = reg_0079;
    39: op1_08_in12 = reg_0128;
    40: op1_08_in12 = reg_0445;
    41: op1_08_in12 = reg_0704;
    42: op1_08_in12 = reg_0886;
    44: op1_08_in12 = reg_0344;
    77: op1_08_in12 = reg_0344;
    45: op1_08_in12 = imem01_in[15:12];
    47: op1_08_in12 = reg_0257;
    48: op1_08_in12 = reg_0210;
    49: op1_08_in12 = reg_0657;
    52: op1_08_in12 = reg_0387;
    55: op1_08_in12 = reg_0186;
    56: op1_08_in12 = imem01_in[19:16];
    57: op1_08_in12 = imem02_in[87:84];
    58: op1_08_in12 = reg_0060;
    59: op1_08_in12 = reg_0087;
    60: op1_08_in12 = reg_0568;
    61: op1_08_in12 = reg_1057;
    62: op1_08_in12 = reg_0497;
    63: op1_08_in12 = reg_0474;
    64: op1_08_in12 = reg_0480;
    65: op1_08_in12 = reg_0873;
    66: op1_08_in12 = reg_0290;
    67: op1_08_in12 = reg_0643;
    68: op1_08_in12 = imem05_in[7:4];
    69: op1_08_in12 = reg_0706;
    70: op1_08_in12 = reg_0867;
    71: op1_08_in12 = imem04_in[59:56];
    72: op1_08_in12 = reg_0451;
    73: op1_08_in12 = reg_0077;
    90: op1_08_in12 = reg_0077;
    74: op1_08_in12 = reg_0368;
    75: op1_08_in12 = reg_0067;
    76: op1_08_in12 = reg_0807;
    78: op1_08_in12 = reg_0184;
    79: op1_08_in12 = reg_0453;
    83: op1_08_in12 = reg_0453;
    80: op1_08_in12 = reg_0840;
    81: op1_08_in12 = reg_1006;
    82: op1_08_in12 = reg_0291;
    84: op1_08_in12 = reg_0965;
    85: op1_08_in12 = reg_0772;
    86: op1_08_in12 = reg_0395;
    87: op1_08_in12 = reg_0165;
    88: op1_08_in12 = reg_0207;
    89: op1_08_in12 = reg_0703;
    91: op1_08_in12 = reg_0832;
    92: op1_08_in12 = reg_0624;
    93: op1_08_in12 = reg_0795;
    94: op1_08_in12 = reg_0141;
    95: op1_08_in12 = reg_0944;
    96: op1_08_in12 = reg_0792;
    97: op1_08_in12 = reg_1005;
    default: op1_08_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv12 = 1;
    6: op1_08_inv12 = 1;
    7: op1_08_inv12 = 1;
    8: op1_08_inv12 = 1;
    9: op1_08_inv12 = 1;
    10: op1_08_inv12 = 1;
    11: op1_08_inv12 = 1;
    12: op1_08_inv12 = 1;
    14: op1_08_inv12 = 1;
    16: op1_08_inv12 = 1;
    19: op1_08_inv12 = 1;
    20: op1_08_inv12 = 1;
    28: op1_08_inv12 = 1;
    29: op1_08_inv12 = 1;
    31: op1_08_inv12 = 1;
    32: op1_08_inv12 = 1;
    33: op1_08_inv12 = 1;
    34: op1_08_inv12 = 1;
    35: op1_08_inv12 = 1;
    37: op1_08_inv12 = 1;
    47: op1_08_inv12 = 1;
    48: op1_08_inv12 = 1;
    50: op1_08_inv12 = 1;
    52: op1_08_inv12 = 1;
    53: op1_08_inv12 = 1;
    56: op1_08_inv12 = 1;
    57: op1_08_inv12 = 1;
    59: op1_08_inv12 = 1;
    61: op1_08_inv12 = 1;
    66: op1_08_inv12 = 1;
    68: op1_08_inv12 = 1;
    69: op1_08_inv12 = 1;
    72: op1_08_inv12 = 1;
    73: op1_08_inv12 = 1;
    76: op1_08_inv12 = 1;
    78: op1_08_inv12 = 1;
    79: op1_08_inv12 = 1;
    80: op1_08_inv12 = 1;
    81: op1_08_inv12 = 1;
    82: op1_08_inv12 = 1;
    84: op1_08_inv12 = 1;
    85: op1_08_inv12 = 1;
    86: op1_08_inv12 = 1;
    87: op1_08_inv12 = 1;
    89: op1_08_inv12 = 1;
    90: op1_08_inv12 = 1;
    95: op1_08_inv12 = 1;
    96: op1_08_inv12 = 1;
    default: op1_08_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in13 = reg_0149;
    6: op1_08_in13 = reg_0553;
    7: op1_08_in13 = reg_0170;
    8: op1_08_in13 = reg_0659;
    9: op1_08_in13 = reg_0266;
    10: op1_08_in13 = reg_0976;
    11: op1_08_in13 = reg_0618;
    12: op1_08_in13 = reg_0319;
    13: op1_08_in13 = reg_0209;
    14: op1_08_in13 = reg_0121;
    15: op1_08_in13 = reg_0985;
    16: op1_08_in13 = reg_0700;
    17: op1_08_in13 = reg_0466;
    18: op1_08_in13 = reg_0612;
    19: op1_08_in13 = reg_0187;
    20: op1_08_in13 = reg_0390;
    21: op1_08_in13 = reg_0451;
    22: op1_08_in13 = imem06_in[27:24];
    23: op1_08_in13 = reg_0827;
    24: op1_08_in13 = reg_0942;
    25: op1_08_in13 = reg_0753;
    26: op1_08_in13 = imem02_in[3:0];
    85: op1_08_in13 = imem02_in[3:0];
    27: op1_08_in13 = reg_0723;
    89: op1_08_in13 = reg_0723;
    28: op1_08_in13 = imem01_in[31:28];
    29: op1_08_in13 = reg_0611;
    30: op1_08_in13 = reg_0444;
    31: op1_08_in13 = imem01_in[27:24];
    32: op1_08_in13 = reg_0986;
    33: op1_08_in13 = reg_1020;
    61: op1_08_in13 = reg_1020;
    34: op1_08_in13 = reg_0433;
    69: op1_08_in13 = reg_0433;
    35: op1_08_in13 = reg_1049;
    36: op1_08_in13 = reg_0006;
    37: op1_08_in13 = reg_1016;
    38: op1_08_in13 = imem03_in[31:28];
    39: op1_08_in13 = reg_0156;
    86: op1_08_in13 = reg_0156;
    40: op1_08_in13 = reg_0434;
    41: op1_08_in13 = reg_0726;
    42: op1_08_in13 = reg_0857;
    43: op1_08_in13 = imem04_in[27:24];
    44: op1_08_in13 = reg_0264;
    45: op1_08_in13 = imem01_in[35:32];
    46: op1_08_in13 = reg_0290;
    47: op1_08_in13 = reg_0785;
    48: op1_08_in13 = reg_0203;
    49: op1_08_in13 = reg_0326;
    50: op1_08_in13 = reg_0473;
    52: op1_08_in13 = reg_0804;
    53: op1_08_in13 = reg_0805;
    55: op1_08_in13 = imem01_in[15:12];
    56: op1_08_in13 = imem01_in[23:20];
    57: op1_08_in13 = imem02_in[119:116];
    58: op1_08_in13 = reg_0681;
    59: op1_08_in13 = reg_0037;
    60: op1_08_in13 = reg_0524;
    62: op1_08_in13 = reg_0132;
    63: op1_08_in13 = reg_0471;
    64: op1_08_in13 = reg_0467;
    65: op1_08_in13 = reg_0098;
    66: op1_08_in13 = reg_0233;
    67: op1_08_in13 = reg_0516;
    68: op1_08_in13 = imem05_in[51:48];
    70: op1_08_in13 = reg_0792;
    71: op1_08_in13 = imem04_in[67:64];
    72: op1_08_in13 = reg_0457;
    73: op1_08_in13 = reg_0884;
    82: op1_08_in13 = reg_0884;
    74: op1_08_in13 = reg_0372;
    75: op1_08_in13 = reg_0014;
    76: op1_08_in13 = reg_0782;
    77: op1_08_in13 = reg_0244;
    79: op1_08_in13 = reg_0477;
    80: op1_08_in13 = reg_0484;
    81: op1_08_in13 = reg_0511;
    83: op1_08_in13 = reg_0462;
    84: op1_08_in13 = imem06_in[59:56];
    87: op1_08_in13 = reg_0159;
    88: op1_08_in13 = reg_0211;
    90: op1_08_in13 = reg_0359;
    91: op1_08_in13 = reg_0116;
    92: op1_08_in13 = imem03_in[15:12];
    93: op1_08_in13 = reg_0949;
    94: op1_08_in13 = reg_0269;
    95: op1_08_in13 = reg_0217;
    96: op1_08_in13 = reg_0606;
    97: op1_08_in13 = reg_0292;
    default: op1_08_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv13 = 1;
    6: op1_08_inv13 = 1;
    7: op1_08_inv13 = 1;
    9: op1_08_inv13 = 1;
    11: op1_08_inv13 = 1;
    12: op1_08_inv13 = 1;
    13: op1_08_inv13 = 1;
    14: op1_08_inv13 = 1;
    17: op1_08_inv13 = 1;
    18: op1_08_inv13 = 1;
    19: op1_08_inv13 = 1;
    21: op1_08_inv13 = 1;
    23: op1_08_inv13 = 1;
    24: op1_08_inv13 = 1;
    25: op1_08_inv13 = 1;
    29: op1_08_inv13 = 1;
    31: op1_08_inv13 = 1;
    33: op1_08_inv13 = 1;
    35: op1_08_inv13 = 1;
    36: op1_08_inv13 = 1;
    42: op1_08_inv13 = 1;
    44: op1_08_inv13 = 1;
    45: op1_08_inv13 = 1;
    48: op1_08_inv13 = 1;
    55: op1_08_inv13 = 1;
    60: op1_08_inv13 = 1;
    61: op1_08_inv13 = 1;
    65: op1_08_inv13 = 1;
    66: op1_08_inv13 = 1;
    67: op1_08_inv13 = 1;
    69: op1_08_inv13 = 1;
    71: op1_08_inv13 = 1;
    73: op1_08_inv13 = 1;
    75: op1_08_inv13 = 1;
    76: op1_08_inv13 = 1;
    79: op1_08_inv13 = 1;
    81: op1_08_inv13 = 1;
    83: op1_08_inv13 = 1;
    85: op1_08_inv13 = 1;
    87: op1_08_inv13 = 1;
    88: op1_08_inv13 = 1;
    89: op1_08_inv13 = 1;
    91: op1_08_inv13 = 1;
    93: op1_08_inv13 = 1;
    94: op1_08_inv13 = 1;
    95: op1_08_inv13 = 1;
    default: op1_08_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in14 = reg_0150;
    6: op1_08_in14 = reg_0303;
    8: op1_08_in14 = reg_0325;
    9: op1_08_in14 = reg_0136;
    10: op1_08_in14 = reg_0994;
    11: op1_08_in14 = reg_0627;
    12: op1_08_in14 = reg_0369;
    13: op1_08_in14 = reg_0199;
    14: op1_08_in14 = imem02_in[23:20];
    15: op1_08_in14 = reg_0998;
    16: op1_08_in14 = reg_0424;
    17: op1_08_in14 = reg_0456;
    18: op1_08_in14 = reg_0402;
    19: op1_08_in14 = reg_0213;
    20: op1_08_in14 = reg_0401;
    21: op1_08_in14 = reg_0200;
    50: op1_08_in14 = reg_0200;
    22: op1_08_in14 = imem06_in[55:52];
    23: op1_08_in14 = reg_0251;
    24: op1_08_in14 = reg_0972;
    25: op1_08_in14 = reg_0805;
    26: op1_08_in14 = imem02_in[55:52];
    27: op1_08_in14 = reg_0717;
    41: op1_08_in14 = reg_0717;
    28: op1_08_in14 = imem01_in[119:116];
    29: op1_08_in14 = reg_0623;
    30: op1_08_in14 = reg_0420;
    31: op1_08_in14 = imem01_in[55:52];
    32: op1_08_in14 = reg_0980;
    33: op1_08_in14 = reg_1005;
    34: op1_08_in14 = reg_0428;
    35: op1_08_in14 = reg_0358;
    66: op1_08_in14 = reg_0358;
    36: op1_08_in14 = reg_1008;
    37: op1_08_in14 = reg_0932;
    61: op1_08_in14 = reg_0932;
    38: op1_08_in14 = imem03_in[59:56];
    39: op1_08_in14 = reg_0130;
    40: op1_08_in14 = reg_0443;
    42: op1_08_in14 = reg_0338;
    43: op1_08_in14 = imem04_in[35:32];
    44: op1_08_in14 = reg_0383;
    45: op1_08_in14 = imem01_in[115:112];
    46: op1_08_in14 = reg_0818;
    47: op1_08_in14 = reg_0147;
    48: op1_08_in14 = reg_0196;
    49: op1_08_in14 = reg_0656;
    52: op1_08_in14 = reg_0388;
    53: op1_08_in14 = reg_0002;
    55: op1_08_in14 = imem01_in[35:32];
    56: op1_08_in14 = imem01_in[39:36];
    57: op1_08_in14 = imem02_in[127:124];
    58: op1_08_in14 = reg_0099;
    59: op1_08_in14 = reg_0867;
    60: op1_08_in14 = reg_0014;
    62: op1_08_in14 = reg_0135;
    63: op1_08_in14 = reg_0479;
    64: op1_08_in14 = reg_0471;
    65: op1_08_in14 = reg_0887;
    67: op1_08_in14 = reg_0347;
    68: op1_08_in14 = imem05_in[79:76];
    69: op1_08_in14 = reg_0744;
    70: op1_08_in14 = reg_0261;
    71: op1_08_in14 = reg_1004;
    72: op1_08_in14 = reg_0476;
    73: op1_08_in14 = reg_0872;
    74: op1_08_in14 = reg_0608;
    75: op1_08_in14 = reg_0302;
    76: op1_08_in14 = reg_0022;
    77: op1_08_in14 = reg_0021;
    79: op1_08_in14 = reg_0473;
    80: op1_08_in14 = imem03_in[3:0];
    82: op1_08_in14 = imem03_in[3:0];
    81: op1_08_in14 = reg_1009;
    83: op1_08_in14 = reg_0191;
    84: op1_08_in14 = imem06_in[91:88];
    85: op1_08_in14 = imem02_in[11:8];
    86: op1_08_in14 = reg_0912;
    87: op1_08_in14 = reg_0726;
    88: op1_08_in14 = reg_0205;
    89: op1_08_in14 = reg_0449;
    90: op1_08_in14 = reg_0329;
    91: op1_08_in14 = reg_1033;
    92: op1_08_in14 = imem03_in[47:44];
    93: op1_08_in14 = imem06_in[23:20];
    94: op1_08_in14 = reg_0057;
    95: op1_08_in14 = reg_0954;
    96: op1_08_in14 = reg_0029;
    97: op1_08_in14 = reg_0909;
    default: op1_08_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv14 = 1;
    6: op1_08_inv14 = 1;
    9: op1_08_inv14 = 1;
    11: op1_08_inv14 = 1;
    12: op1_08_inv14 = 1;
    14: op1_08_inv14 = 1;
    16: op1_08_inv14 = 1;
    18: op1_08_inv14 = 1;
    23: op1_08_inv14 = 1;
    24: op1_08_inv14 = 1;
    26: op1_08_inv14 = 1;
    27: op1_08_inv14 = 1;
    33: op1_08_inv14 = 1;
    36: op1_08_inv14 = 1;
    37: op1_08_inv14 = 1;
    38: op1_08_inv14 = 1;
    39: op1_08_inv14 = 1;
    42: op1_08_inv14 = 1;
    44: op1_08_inv14 = 1;
    46: op1_08_inv14 = 1;
    50: op1_08_inv14 = 1;
    53: op1_08_inv14 = 1;
    56: op1_08_inv14 = 1;
    59: op1_08_inv14 = 1;
    61: op1_08_inv14 = 1;
    63: op1_08_inv14 = 1;
    65: op1_08_inv14 = 1;
    71: op1_08_inv14 = 1;
    73: op1_08_inv14 = 1;
    77: op1_08_inv14 = 1;
    80: op1_08_inv14 = 1;
    82: op1_08_inv14 = 1;
    83: op1_08_inv14 = 1;
    84: op1_08_inv14 = 1;
    86: op1_08_inv14 = 1;
    87: op1_08_inv14 = 1;
    92: op1_08_inv14 = 1;
    default: op1_08_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in15 = reg_0129;
    6: op1_08_in15 = reg_0289;
    8: op1_08_in15 = reg_0324;
    9: op1_08_in15 = reg_0142;
    10: op1_08_in15 = imem04_in[11:8];
    11: op1_08_in15 = reg_0622;
    12: op1_08_in15 = reg_0309;
    13: op1_08_in15 = imem01_in[7:4];
    14: op1_08_in15 = imem02_in[39:36];
    15: op1_08_in15 = reg_0995;
    16: op1_08_in15 = reg_0434;
    17: op1_08_in15 = reg_0207;
    83: op1_08_in15 = reg_0207;
    18: op1_08_in15 = reg_0344;
    19: op1_08_in15 = reg_0212;
    20: op1_08_in15 = reg_0800;
    21: op1_08_in15 = reg_0203;
    22: op1_08_in15 = imem06_in[59:56];
    23: op1_08_in15 = reg_0148;
    24: op1_08_in15 = reg_0256;
    25: op1_08_in15 = imem07_in[11:8];
    26: op1_08_in15 = imem02_in[63:60];
    27: op1_08_in15 = reg_0724;
    28: op1_08_in15 = imem01_in[123:120];
    29: op1_08_in15 = imem06_in[31:28];
    30: op1_08_in15 = reg_0180;
    31: op1_08_in15 = reg_0786;
    32: op1_08_in15 = reg_0978;
    33: op1_08_in15 = reg_0292;
    34: op1_08_in15 = reg_0438;
    35: op1_08_in15 = reg_0933;
    36: op1_08_in15 = reg_1049;
    37: op1_08_in15 = reg_0740;
    38: op1_08_in15 = imem03_in[63:60];
    39: op1_08_in15 = reg_0604;
    40: op1_08_in15 = reg_0437;
    41: op1_08_in15 = reg_0714;
    42: op1_08_in15 = reg_0516;
    43: op1_08_in15 = imem04_in[67:64];
    44: op1_08_in15 = reg_0617;
    45: op1_08_in15 = imem01_in[127:124];
    46: op1_08_in15 = reg_0817;
    47: op1_08_in15 = reg_0133;
    48: op1_08_in15 = reg_0037;
    49: op1_08_in15 = reg_0639;
    50: op1_08_in15 = imem01_in[43:40];
    52: op1_08_in15 = reg_0384;
    53: op1_08_in15 = reg_0744;
    55: op1_08_in15 = imem01_in[47:44];
    56: op1_08_in15 = imem01_in[47:44];
    57: op1_08_in15 = reg_0655;
    58: op1_08_in15 = reg_0445;
    59: op1_08_in15 = reg_0086;
    60: op1_08_in15 = reg_0552;
    61: op1_08_in15 = reg_0524;
    62: op1_08_in15 = reg_0139;
    63: op1_08_in15 = reg_0208;
    64: op1_08_in15 = reg_0479;
    65: op1_08_in15 = reg_0908;
    66: op1_08_in15 = reg_0739;
    67: op1_08_in15 = reg_0007;
    68: op1_08_in15 = imem05_in[119:116];
    69: op1_08_in15 = reg_0419;
    70: op1_08_in15 = reg_0765;
    71: op1_08_in15 = reg_1003;
    72: op1_08_in15 = reg_0462;
    73: op1_08_in15 = imem03_in[7:4];
    74: op1_08_in15 = reg_0083;
    75: op1_08_in15 = reg_0401;
    76: op1_08_in15 = reg_0545;
    77: op1_08_in15 = reg_0699;
    79: op1_08_in15 = reg_0456;
    80: op1_08_in15 = imem03_in[99:96];
    81: op1_08_in15 = reg_0912;
    82: op1_08_in15 = imem03_in[15:12];
    84: op1_08_in15 = imem06_in[103:100];
    85: op1_08_in15 = imem02_in[19:16];
    86: op1_08_in15 = reg_0048;
    87: op1_08_in15 = reg_0718;
    88: op1_08_in15 = reg_0192;
    89: op1_08_in15 = reg_0157;
    90: op1_08_in15 = reg_0389;
    91: op1_08_in15 = reg_0115;
    92: op1_08_in15 = imem03_in[59:56];
    93: op1_08_in15 = imem06_in[55:52];
    94: op1_08_in15 = reg_0958;
    95: op1_08_in15 = reg_0143;
    96: op1_08_in15 = reg_0811;
    97: op1_08_in15 = reg_0067;
    default: op1_08_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv15 = 1;
    6: op1_08_inv15 = 1;
    10: op1_08_inv15 = 1;
    12: op1_08_inv15 = 1;
    15: op1_08_inv15 = 1;
    16: op1_08_inv15 = 1;
    17: op1_08_inv15 = 1;
    18: op1_08_inv15 = 1;
    22: op1_08_inv15 = 1;
    23: op1_08_inv15 = 1;
    28: op1_08_inv15 = 1;
    29: op1_08_inv15 = 1;
    35: op1_08_inv15 = 1;
    37: op1_08_inv15 = 1;
    39: op1_08_inv15 = 1;
    46: op1_08_inv15 = 1;
    48: op1_08_inv15 = 1;
    55: op1_08_inv15 = 1;
    56: op1_08_inv15 = 1;
    59: op1_08_inv15 = 1;
    64: op1_08_inv15 = 1;
    67: op1_08_inv15 = 1;
    70: op1_08_inv15 = 1;
    71: op1_08_inv15 = 1;
    73: op1_08_inv15 = 1;
    74: op1_08_inv15 = 1;
    75: op1_08_inv15 = 1;
    76: op1_08_inv15 = 1;
    80: op1_08_inv15 = 1;
    81: op1_08_inv15 = 1;
    83: op1_08_inv15 = 1;
    84: op1_08_inv15 = 1;
    85: op1_08_inv15 = 1;
    86: op1_08_inv15 = 1;
    87: op1_08_inv15 = 1;
    88: op1_08_inv15 = 1;
    89: op1_08_inv15 = 1;
    90: op1_08_inv15 = 1;
    93: op1_08_inv15 = 1;
    94: op1_08_inv15 = 1;
    default: op1_08_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in16 = imem06_in[11:8];
    62: op1_08_in16 = imem06_in[11:8];
    6: op1_08_in16 = reg_0054;
    8: op1_08_in16 = reg_0353;
    9: op1_08_in16 = reg_0143;
    10: op1_08_in16 = imem04_in[15:12];
    11: op1_08_in16 = reg_0381;
    12: op1_08_in16 = reg_0987;
    13: op1_08_in16 = imem01_in[15:12];
    14: op1_08_in16 = imem02_in[103:100];
    15: op1_08_in16 = reg_0996;
    16: op1_08_in16 = reg_0440;
    17: op1_08_in16 = reg_0186;
    18: op1_08_in16 = reg_0372;
    90: op1_08_in16 = reg_0372;
    19: op1_08_in16 = reg_0199;
    20: op1_08_in16 = imem07_in[23:20];
    21: op1_08_in16 = reg_0194;
    22: op1_08_in16 = imem06_in[83:80];
    23: op1_08_in16 = reg_0133;
    24: op1_08_in16 = reg_0813;
    25: op1_08_in16 = imem07_in[19:16];
    26: op1_08_in16 = imem02_in[119:116];
    27: op1_08_in16 = reg_0705;
    28: op1_08_in16 = reg_0218;
    29: op1_08_in16 = imem06_in[47:44];
    30: op1_08_in16 = reg_0165;
    40: op1_08_in16 = reg_0165;
    31: op1_08_in16 = reg_0224;
    32: op1_08_in16 = reg_0997;
    33: op1_08_in16 = reg_0078;
    34: op1_08_in16 = reg_0180;
    35: op1_08_in16 = reg_0396;
    36: op1_08_in16 = reg_0245;
    37: op1_08_in16 = reg_0276;
    38: op1_08_in16 = imem03_in[71:68];
    39: op1_08_in16 = reg_0026;
    41: op1_08_in16 = reg_0703;
    42: op1_08_in16 = reg_0762;
    46: op1_08_in16 = reg_0762;
    43: op1_08_in16 = imem04_in[79:76];
    44: op1_08_in16 = reg_0633;
    45: op1_08_in16 = reg_0013;
    47: op1_08_in16 = reg_0156;
    48: op1_08_in16 = reg_1053;
    49: op1_08_in16 = reg_0334;
    50: op1_08_in16 = imem01_in[47:44];
    52: op1_08_in16 = reg_0629;
    53: op1_08_in16 = reg_0315;
    55: op1_08_in16 = imem01_in[119:116];
    56: op1_08_in16 = reg_0786;
    57: op1_08_in16 = reg_0649;
    58: op1_08_in16 = reg_0370;
    59: op1_08_in16 = imem03_in[7:4];
    60: op1_08_in16 = reg_0517;
    61: op1_08_in16 = reg_0014;
    63: op1_08_in16 = reg_0191;
    64: op1_08_in16 = reg_0209;
    65: op1_08_in16 = reg_0645;
    66: op1_08_in16 = reg_0368;
    67: op1_08_in16 = reg_0086;
    68: op1_08_in16 = imem05_in[127:124];
    69: op1_08_in16 = reg_0838;
    70: op1_08_in16 = reg_0961;
    71: op1_08_in16 = reg_0055;
    72: op1_08_in16 = reg_0471;
    73: op1_08_in16 = imem03_in[11:8];
    74: op1_08_in16 = reg_0867;
    75: op1_08_in16 = reg_0284;
    76: op1_08_in16 = imem07_in[79:76];
    77: op1_08_in16 = reg_0270;
    79: op1_08_in16 = reg_0478;
    80: op1_08_in16 = reg_0580;
    81: op1_08_in16 = reg_0888;
    82: op1_08_in16 = imem03_in[27:24];
    83: op1_08_in16 = reg_0198;
    84: op1_08_in16 = imem06_in[115:112];
    85: op1_08_in16 = imem02_in[27:24];
    86: op1_08_in16 = reg_1005;
    87: op1_08_in16 = reg_0805;
    88: op1_08_in16 = imem01_in[11:8];
    89: op1_08_in16 = reg_0184;
    91: op1_08_in16 = reg_0877;
    92: op1_08_in16 = imem03_in[119:116];
    93: op1_08_in16 = imem06_in[91:88];
    94: op1_08_in16 = reg_0675;
    95: op1_08_in16 = reg_0139;
    96: op1_08_in16 = reg_0177;
    97: op1_08_in16 = reg_0243;
    default: op1_08_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv16 = 1;
    8: op1_08_inv16 = 1;
    9: op1_08_inv16 = 1;
    10: op1_08_inv16 = 1;
    11: op1_08_inv16 = 1;
    15: op1_08_inv16 = 1;
    18: op1_08_inv16 = 1;
    19: op1_08_inv16 = 1;
    20: op1_08_inv16 = 1;
    22: op1_08_inv16 = 1;
    25: op1_08_inv16 = 1;
    29: op1_08_inv16 = 1;
    30: op1_08_inv16 = 1;
    31: op1_08_inv16 = 1;
    32: op1_08_inv16 = 1;
    34: op1_08_inv16 = 1;
    35: op1_08_inv16 = 1;
    36: op1_08_inv16 = 1;
    38: op1_08_inv16 = 1;
    41: op1_08_inv16 = 1;
    45: op1_08_inv16 = 1;
    46: op1_08_inv16 = 1;
    47: op1_08_inv16 = 1;
    50: op1_08_inv16 = 1;
    52: op1_08_inv16 = 1;
    56: op1_08_inv16 = 1;
    57: op1_08_inv16 = 1;
    58: op1_08_inv16 = 1;
    60: op1_08_inv16 = 1;
    61: op1_08_inv16 = 1;
    62: op1_08_inv16 = 1;
    63: op1_08_inv16 = 1;
    66: op1_08_inv16 = 1;
    67: op1_08_inv16 = 1;
    68: op1_08_inv16 = 1;
    69: op1_08_inv16 = 1;
    71: op1_08_inv16 = 1;
    75: op1_08_inv16 = 1;
    79: op1_08_inv16 = 1;
    80: op1_08_inv16 = 1;
    83: op1_08_inv16 = 1;
    87: op1_08_inv16 = 1;
    88: op1_08_inv16 = 1;
    89: op1_08_inv16 = 1;
    90: op1_08_inv16 = 1;
    91: op1_08_inv16 = 1;
    92: op1_08_inv16 = 1;
    93: op1_08_inv16 = 1;
    95: op1_08_inv16 = 1;
    default: op1_08_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in17 = reg_0607;
    6: op1_08_in17 = reg_0043;
    8: op1_08_in17 = reg_0310;
    9: op1_08_in17 = reg_0130;
    10: op1_08_in17 = imem04_in[71:68];
    11: op1_08_in17 = reg_0367;
    12: op1_08_in17 = reg_0984;
    13: op1_08_in17 = imem01_in[55:52];
    14: op1_08_in17 = imem02_in[107:104];
    15: op1_08_in17 = reg_1001;
    16: op1_08_in17 = reg_0427;
    17: op1_08_in17 = reg_0198;
    18: op1_08_in17 = reg_0407;
    19: op1_08_in17 = imem01_in[7:4];
    20: op1_08_in17 = imem07_in[75:72];
    21: op1_08_in17 = imem01_in[11:8];
    22: op1_08_in17 = imem06_in[95:92];
    23: op1_08_in17 = reg_0150;
    24: op1_08_in17 = reg_0785;
    25: op1_08_in17 = imem07_in[43:40];
    44: op1_08_in17 = imem07_in[43:40];
    26: op1_08_in17 = reg_0758;
    27: op1_08_in17 = reg_0711;
    28: op1_08_in17 = reg_0299;
    29: op1_08_in17 = imem06_in[51:48];
    30: op1_08_in17 = reg_0177;
    40: op1_08_in17 = reg_0177;
    31: op1_08_in17 = reg_0555;
    32: op1_08_in17 = imem04_in[31:28];
    33: op1_08_in17 = reg_0259;
    34: op1_08_in17 = reg_0172;
    35: op1_08_in17 = reg_0823;
    36: op1_08_in17 = reg_0322;
    37: op1_08_in17 = reg_0063;
    38: op1_08_in17 = imem03_in[87:84];
    39: op1_08_in17 = reg_1028;
    41: op1_08_in17 = reg_0708;
    42: op1_08_in17 = reg_0336;
    43: op1_08_in17 = imem04_in[127:124];
    45: op1_08_in17 = reg_0786;
    55: op1_08_in17 = reg_0786;
    46: op1_08_in17 = reg_0482;
    47: op1_08_in17 = reg_0143;
    48: op1_08_in17 = reg_0860;
    49: op1_08_in17 = reg_0290;
    50: op1_08_in17 = imem01_in[51:48];
    52: op1_08_in17 = reg_0017;
    53: op1_08_in17 = reg_0180;
    56: op1_08_in17 = reg_1056;
    57: op1_08_in17 = reg_0637;
    58: op1_08_in17 = reg_0807;
    59: op1_08_in17 = imem03_in[39:36];
    60: op1_08_in17 = reg_0542;
    61: op1_08_in17 = reg_0276;
    62: op1_08_in17 = reg_0391;
    63: op1_08_in17 = reg_0207;
    64: op1_08_in17 = reg_0190;
    65: op1_08_in17 = reg_0664;
    66: op1_08_in17 = reg_0089;
    67: op1_08_in17 = reg_0016;
    68: op1_08_in17 = reg_0940;
    69: op1_08_in17 = reg_0174;
    70: op1_08_in17 = reg_0743;
    71: op1_08_in17 = reg_1005;
    72: op1_08_in17 = reg_0479;
    73: op1_08_in17 = imem03_in[27:24];
    74: op1_08_in17 = reg_0814;
    75: op1_08_in17 = reg_0243;
    76: op1_08_in17 = imem07_in[91:88];
    77: op1_08_in17 = imem07_in[31:28];
    79: op1_08_in17 = reg_0458;
    80: op1_08_in17 = reg_0662;
    81: op1_08_in17 = reg_0568;
    82: op1_08_in17 = imem03_in[31:28];
    83: op1_08_in17 = reg_0201;
    84: op1_08_in17 = reg_0080;
    85: op1_08_in17 = imem02_in[103:100];
    86: op1_08_in17 = reg_0540;
    87: op1_08_in17 = reg_0303;
    88: op1_08_in17 = imem01_in[87:84];
    90: op1_08_in17 = reg_0608;
    91: op1_08_in17 = imem02_in[55:52];
    92: op1_08_in17 = imem03_in[123:120];
    93: op1_08_in17 = reg_0010;
    94: op1_08_in17 = reg_0437;
    95: op1_08_in17 = reg_0275;
    96: op1_08_in17 = imem07_in[51:48];
    97: op1_08_in17 = reg_0495;
    default: op1_08_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_08_inv17 = 1;
    10: op1_08_inv17 = 1;
    13: op1_08_inv17 = 1;
    15: op1_08_inv17 = 1;
    17: op1_08_inv17 = 1;
    19: op1_08_inv17 = 1;
    20: op1_08_inv17 = 1;
    21: op1_08_inv17 = 1;
    23: op1_08_inv17 = 1;
    24: op1_08_inv17 = 1;
    26: op1_08_inv17 = 1;
    29: op1_08_inv17 = 1;
    30: op1_08_inv17 = 1;
    32: op1_08_inv17 = 1;
    33: op1_08_inv17 = 1;
    35: op1_08_inv17 = 1;
    36: op1_08_inv17 = 1;
    38: op1_08_inv17 = 1;
    39: op1_08_inv17 = 1;
    41: op1_08_inv17 = 1;
    45: op1_08_inv17 = 1;
    46: op1_08_inv17 = 1;
    47: op1_08_inv17 = 1;
    48: op1_08_inv17 = 1;
    53: op1_08_inv17 = 1;
    55: op1_08_inv17 = 1;
    57: op1_08_inv17 = 1;
    59: op1_08_inv17 = 1;
    62: op1_08_inv17 = 1;
    63: op1_08_inv17 = 1;
    65: op1_08_inv17 = 1;
    70: op1_08_inv17 = 1;
    73: op1_08_inv17 = 1;
    74: op1_08_inv17 = 1;
    75: op1_08_inv17 = 1;
    80: op1_08_inv17 = 1;
    81: op1_08_inv17 = 1;
    85: op1_08_inv17 = 1;
    87: op1_08_inv17 = 1;
    88: op1_08_inv17 = 1;
    93: op1_08_inv17 = 1;
    94: op1_08_inv17 = 1;
    95: op1_08_inv17 = 1;
    default: op1_08_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in18 = reg_0616;
    39: op1_08_in18 = reg_0616;
    6: op1_08_in18 = reg_0063;
    8: op1_08_in18 = reg_0350;
    9: op1_08_in18 = reg_0155;
    10: op1_08_in18 = imem04_in[79:76];
    32: op1_08_in18 = imem04_in[79:76];
    11: op1_08_in18 = reg_0337;
    12: op1_08_in18 = reg_1001;
    13: op1_08_in18 = imem01_in[87:84];
    14: op1_08_in18 = imem02_in[123:120];
    15: op1_08_in18 = reg_0977;
    16: op1_08_in18 = reg_0435;
    17: op1_08_in18 = reg_0213;
    18: op1_08_in18 = reg_0383;
    19: op1_08_in18 = imem01_in[11:8];
    63: op1_08_in18 = imem01_in[11:8];
    20: op1_08_in18 = reg_0719;
    21: op1_08_in18 = imem01_in[43:40];
    22: op1_08_in18 = imem06_in[103:100];
    23: op1_08_in18 = reg_0144;
    24: op1_08_in18 = reg_0497;
    25: op1_08_in18 = imem07_in[51:48];
    44: op1_08_in18 = imem07_in[51:48];
    26: op1_08_in18 = reg_0261;
    27: op1_08_in18 = reg_0433;
    28: op1_08_in18 = reg_0555;
    29: op1_08_in18 = imem06_in[67:64];
    31: op1_08_in18 = reg_0905;
    33: op1_08_in18 = reg_0296;
    37: op1_08_in18 = reg_0296;
    34: op1_08_in18 = reg_0177;
    35: op1_08_in18 = reg_0784;
    36: op1_08_in18 = reg_0397;
    38: op1_08_in18 = imem03_in[91:88];
    40: op1_08_in18 = reg_0184;
    41: op1_08_in18 = reg_0727;
    42: op1_08_in18 = reg_0761;
    43: op1_08_in18 = reg_0265;
    45: op1_08_in18 = reg_0223;
    46: op1_08_in18 = reg_0089;
    47: op1_08_in18 = reg_0139;
    48: op1_08_in18 = imem01_in[27:24];
    49: op1_08_in18 = reg_0818;
    50: op1_08_in18 = imem01_in[91:88];
    52: op1_08_in18 = imem07_in[19:16];
    53: op1_08_in18 = reg_0181;
    55: op1_08_in18 = reg_0592;
    56: op1_08_in18 = reg_0829;
    57: op1_08_in18 = reg_0739;
    58: op1_08_in18 = reg_0376;
    59: op1_08_in18 = imem03_in[55:52];
    73: op1_08_in18 = imem03_in[55:52];
    60: op1_08_in18 = reg_0531;
    61: op1_08_in18 = reg_0284;
    62: op1_08_in18 = reg_0926;
    64: op1_08_in18 = reg_0199;
    65: op1_08_in18 = reg_0329;
    66: op1_08_in18 = reg_0090;
    67: op1_08_in18 = imem03_in[43:40];
    68: op1_08_in18 = reg_0274;
    69: op1_08_in18 = reg_0162;
    70: op1_08_in18 = reg_0060;
    71: op1_08_in18 = reg_0932;
    72: op1_08_in18 = reg_0191;
    74: op1_08_in18 = reg_0506;
    75: op1_08_in18 = reg_0854;
    76: op1_08_in18 = imem07_in[95:92];
    77: op1_08_in18 = imem07_in[47:44];
    79: op1_08_in18 = reg_0189;
    80: op1_08_in18 = reg_0590;
    81: op1_08_in18 = reg_0067;
    82: op1_08_in18 = imem03_in[51:48];
    83: op1_08_in18 = reg_0212;
    84: op1_08_in18 = reg_0625;
    85: op1_08_in18 = imem02_in[111:108];
    86: op1_08_in18 = reg_0909;
    87: op1_08_in18 = reg_0315;
    88: op1_08_in18 = reg_0106;
    90: op1_08_in18 = reg_0650;
    91: op1_08_in18 = reg_0285;
    92: op1_08_in18 = reg_0317;
    93: op1_08_in18 = reg_0694;
    94: op1_08_in18 = reg_0135;
    95: op1_08_in18 = reg_0013;
    96: op1_08_in18 = imem07_in[67:64];
    97: op1_08_in18 = reg_0627;
    default: op1_08_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv18 = 1;
    12: op1_08_inv18 = 1;
    16: op1_08_inv18 = 1;
    19: op1_08_inv18 = 1;
    24: op1_08_inv18 = 1;
    26: op1_08_inv18 = 1;
    27: op1_08_inv18 = 1;
    29: op1_08_inv18 = 1;
    31: op1_08_inv18 = 1;
    32: op1_08_inv18 = 1;
    34: op1_08_inv18 = 1;
    36: op1_08_inv18 = 1;
    43: op1_08_inv18 = 1;
    44: op1_08_inv18 = 1;
    50: op1_08_inv18 = 1;
    53: op1_08_inv18 = 1;
    55: op1_08_inv18 = 1;
    56: op1_08_inv18 = 1;
    58: op1_08_inv18 = 1;
    60: op1_08_inv18 = 1;
    61: op1_08_inv18 = 1;
    62: op1_08_inv18 = 1;
    64: op1_08_inv18 = 1;
    65: op1_08_inv18 = 1;
    67: op1_08_inv18 = 1;
    79: op1_08_inv18 = 1;
    81: op1_08_inv18 = 1;
    83: op1_08_inv18 = 1;
    84: op1_08_inv18 = 1;
    85: op1_08_inv18 = 1;
    86: op1_08_inv18 = 1;
    90: op1_08_inv18 = 1;
    92: op1_08_inv18 = 1;
    93: op1_08_inv18 = 1;
    94: op1_08_inv18 = 1;
    95: op1_08_inv18 = 1;
    default: op1_08_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in19 = reg_0609;
    6: op1_08_in19 = reg_0072;
    8: op1_08_in19 = reg_0080;
    9: op1_08_in19 = reg_0137;
    10: op1_08_in19 = imem04_in[87:84];
    11: op1_08_in19 = reg_1028;
    12: op1_08_in19 = reg_0978;
    13: op1_08_in19 = imem01_in[91:88];
    14: op1_08_in19 = reg_0666;
    15: op1_08_in19 = reg_0997;
    16: op1_08_in19 = reg_0159;
    17: op1_08_in19 = reg_0205;
    18: op1_08_in19 = reg_1029;
    19: op1_08_in19 = imem01_in[15:12];
    64: op1_08_in19 = imem01_in[15:12];
    20: op1_08_in19 = reg_0723;
    21: op1_08_in19 = imem01_in[51:48];
    22: op1_08_in19 = reg_0630;
    23: op1_08_in19 = imem06_in[19:16];
    24: op1_08_in19 = reg_0135;
    25: op1_08_in19 = imem07_in[63:60];
    44: op1_08_in19 = imem07_in[63:60];
    26: op1_08_in19 = reg_0484;
    27: op1_08_in19 = reg_0442;
    28: op1_08_in19 = reg_0248;
    29: op1_08_in19 = imem06_in[83:80];
    31: op1_08_in19 = reg_1042;
    32: op1_08_in19 = imem04_in[99:96];
    33: op1_08_in19 = reg_0009;
    34: op1_08_in19 = reg_0164;
    35: op1_08_in19 = reg_0377;
    36: op1_08_in19 = reg_0847;
    37: op1_08_in19 = reg_0075;
    38: op1_08_in19 = reg_1007;
    39: op1_08_in19 = reg_0877;
    41: op1_08_in19 = reg_0430;
    42: op1_08_in19 = reg_0876;
    43: op1_08_in19 = reg_0931;
    45: op1_08_in19 = reg_0560;
    46: op1_08_in19 = reg_0077;
    47: op1_08_in19 = reg_0140;
    48: op1_08_in19 = imem01_in[47:44];
    49: op1_08_in19 = reg_0083;
    50: op1_08_in19 = imem01_in[99:96];
    52: op1_08_in19 = imem07_in[47:44];
    53: op1_08_in19 = reg_0179;
    55: op1_08_in19 = reg_1036;
    56: op1_08_in19 = reg_0514;
    57: op1_08_in19 = reg_0372;
    58: op1_08_in19 = reg_0518;
    59: op1_08_in19 = imem03_in[79:76];
    60: op1_08_in19 = imem05_in[11:8];
    61: op1_08_in19 = reg_0243;
    62: op1_08_in19 = reg_0440;
    63: op1_08_in19 = imem01_in[19:16];
    65: op1_08_in19 = reg_0331;
    66: op1_08_in19 = reg_0091;
    67: op1_08_in19 = imem03_in[71:68];
    68: op1_08_in19 = reg_0688;
    69: op1_08_in19 = reg_0160;
    70: op1_08_in19 = reg_0620;
    71: op1_08_in19 = reg_0050;
    72: op1_08_in19 = reg_0189;
    73: op1_08_in19 = imem03_in[107:104];
    74: op1_08_in19 = reg_0084;
    75: op1_08_in19 = reg_0071;
    76: op1_08_in19 = reg_0429;
    77: op1_08_in19 = imem07_in[55:52];
    79: op1_08_in19 = reg_0188;
    80: op1_08_in19 = reg_0823;
    81: op1_08_in19 = reg_0276;
    82: op1_08_in19 = imem03_in[55:52];
    83: op1_08_in19 = imem01_in[7:4];
    84: op1_08_in19 = reg_0694;
    85: op1_08_in19 = imem03_in[3:0];
    86: op1_08_in19 = reg_0799;
    87: op1_08_in19 = reg_0024;
    88: op1_08_in19 = reg_0337;
    90: op1_08_in19 = reg_0776;
    91: op1_08_in19 = reg_0536;
    92: op1_08_in19 = reg_0578;
    93: op1_08_in19 = reg_0244;
    94: op1_08_in19 = reg_0528;
    95: op1_08_in19 = reg_0648;
    96: op1_08_in19 = reg_0720;
    97: op1_08_in19 = imem05_in[19:16];
    default: op1_08_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv19 = 1;
    8: op1_08_inv19 = 1;
    9: op1_08_inv19 = 1;
    13: op1_08_inv19 = 1;
    14: op1_08_inv19 = 1;
    15: op1_08_inv19 = 1;
    17: op1_08_inv19 = 1;
    20: op1_08_inv19 = 1;
    22: op1_08_inv19 = 1;
    23: op1_08_inv19 = 1;
    25: op1_08_inv19 = 1;
    26: op1_08_inv19 = 1;
    27: op1_08_inv19 = 1;
    31: op1_08_inv19 = 1;
    32: op1_08_inv19 = 1;
    33: op1_08_inv19 = 1;
    35: op1_08_inv19 = 1;
    36: op1_08_inv19 = 1;
    38: op1_08_inv19 = 1;
    39: op1_08_inv19 = 1;
    41: op1_08_inv19 = 1;
    42: op1_08_inv19 = 1;
    43: op1_08_inv19 = 1;
    44: op1_08_inv19 = 1;
    46: op1_08_inv19 = 1;
    47: op1_08_inv19 = 1;
    52: op1_08_inv19 = 1;
    53: op1_08_inv19 = 1;
    59: op1_08_inv19 = 1;
    60: op1_08_inv19 = 1;
    61: op1_08_inv19 = 1;
    63: op1_08_inv19 = 1;
    64: op1_08_inv19 = 1;
    67: op1_08_inv19 = 1;
    68: op1_08_inv19 = 1;
    69: op1_08_inv19 = 1;
    70: op1_08_inv19 = 1;
    71: op1_08_inv19 = 1;
    73: op1_08_inv19 = 1;
    74: op1_08_inv19 = 1;
    75: op1_08_inv19 = 1;
    76: op1_08_inv19 = 1;
    77: op1_08_inv19 = 1;
    79: op1_08_inv19 = 1;
    82: op1_08_inv19 = 1;
    83: op1_08_inv19 = 1;
    88: op1_08_inv19 = 1;
    90: op1_08_inv19 = 1;
    91: op1_08_inv19 = 1;
    92: op1_08_inv19 = 1;
    93: op1_08_inv19 = 1;
    94: op1_08_inv19 = 1;
    96: op1_08_inv19 = 1;
    default: op1_08_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in20 = reg_0402;
    6: op1_08_in20 = reg_0827;
    8: op1_08_in20 = reg_0090;
    9: op1_08_in20 = reg_0131;
    10: op1_08_in20 = imem04_in[91:88];
    11: op1_08_in20 = reg_0802;
    71: op1_08_in20 = reg_0802;
    12: op1_08_in20 = reg_0994;
    13: op1_08_in20 = reg_0246;
    14: op1_08_in20 = reg_0639;
    15: op1_08_in20 = imem04_in[35:32];
    16: op1_08_in20 = reg_0182;
    17: op1_08_in20 = reg_0197;
    18: op1_08_in20 = reg_0026;
    19: op1_08_in20 = imem01_in[23:20];
    20: op1_08_in20 = reg_0712;
    21: op1_08_in20 = imem01_in[55:52];
    48: op1_08_in20 = imem01_in[55:52];
    22: op1_08_in20 = reg_0605;
    23: op1_08_in20 = imem06_in[31:28];
    39: op1_08_in20 = imem06_in[31:28];
    24: op1_08_in20 = reg_0152;
    25: op1_08_in20 = imem07_in[67:64];
    77: op1_08_in20 = imem07_in[67:64];
    26: op1_08_in20 = imem03_in[15:12];
    27: op1_08_in20 = reg_0443;
    28: op1_08_in20 = reg_0544;
    29: op1_08_in20 = imem06_in[87:84];
    31: op1_08_in20 = reg_0869;
    32: op1_08_in20 = imem04_in[111:108];
    33: op1_08_in20 = reg_0059;
    34: op1_08_in20 = reg_0171;
    35: op1_08_in20 = reg_0767;
    36: op1_08_in20 = reg_0543;
    37: op1_08_in20 = reg_0074;
    38: op1_08_in20 = reg_0245;
    41: op1_08_in20 = reg_0433;
    42: op1_08_in20 = reg_0086;
    90: op1_08_in20 = reg_0086;
    43: op1_08_in20 = reg_0313;
    44: op1_08_in20 = imem07_in[87:84];
    45: op1_08_in20 = reg_0510;
    46: op1_08_in20 = imem03_in[63:60];
    47: op1_08_in20 = imem06_in[19:16];
    49: op1_08_in20 = reg_0482;
    50: op1_08_in20 = imem01_in[103:100];
    52: op1_08_in20 = imem07_in[51:48];
    53: op1_08_in20 = reg_0177;
    55: op1_08_in20 = reg_0253;
    56: op1_08_in20 = reg_1037;
    57: op1_08_in20 = reg_0818;
    58: op1_08_in20 = reg_0234;
    59: op1_08_in20 = imem03_in[91:88];
    60: op1_08_in20 = imem05_in[55:52];
    61: op1_08_in20 = reg_0658;
    62: op1_08_in20 = reg_0395;
    63: op1_08_in20 = imem01_in[39:36];
    64: op1_08_in20 = imem01_in[27:24];
    65: op1_08_in20 = reg_0335;
    66: op1_08_in20 = reg_0484;
    67: op1_08_in20 = imem03_in[87:84];
    68: op1_08_in20 = reg_0221;
    69: op1_08_in20 = reg_0166;
    70: op1_08_in20 = reg_1007;
    72: op1_08_in20 = reg_0187;
    73: op1_08_in20 = imem03_in[119:116];
    74: op1_08_in20 = imem03_in[27:24];
    75: op1_08_in20 = imem05_in[15:12];
    76: op1_08_in20 = reg_0646;
    79: op1_08_in20 = imem01_in[15:12];
    80: op1_08_in20 = reg_0278;
    81: op1_08_in20 = reg_0065;
    82: op1_08_in20 = imem03_in[71:68];
    83: op1_08_in20 = imem01_in[87:84];
    84: op1_08_in20 = reg_1019;
    85: op1_08_in20 = imem03_in[7:4];
    86: op1_08_in20 = reg_0058;
    87: op1_08_in20 = reg_0731;
    88: op1_08_in20 = reg_0503;
    91: op1_08_in20 = reg_0075;
    92: op1_08_in20 = reg_0007;
    93: op1_08_in20 = reg_0229;
    94: op1_08_in20 = reg_0490;
    95: op1_08_in20 = reg_0583;
    96: op1_08_in20 = reg_0923;
    97: op1_08_in20 = imem05_in[39:36];
    default: op1_08_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    11: op1_08_inv20 = 1;
    12: op1_08_inv20 = 1;
    13: op1_08_inv20 = 1;
    15: op1_08_inv20 = 1;
    18: op1_08_inv20 = 1;
    19: op1_08_inv20 = 1;
    25: op1_08_inv20 = 1;
    27: op1_08_inv20 = 1;
    28: op1_08_inv20 = 1;
    31: op1_08_inv20 = 1;
    32: op1_08_inv20 = 1;
    33: op1_08_inv20 = 1;
    34: op1_08_inv20 = 1;
    35: op1_08_inv20 = 1;
    38: op1_08_inv20 = 1;
    41: op1_08_inv20 = 1;
    43: op1_08_inv20 = 1;
    44: op1_08_inv20 = 1;
    45: op1_08_inv20 = 1;
    46: op1_08_inv20 = 1;
    50: op1_08_inv20 = 1;
    53: op1_08_inv20 = 1;
    55: op1_08_inv20 = 1;
    57: op1_08_inv20 = 1;
    58: op1_08_inv20 = 1;
    59: op1_08_inv20 = 1;
    60: op1_08_inv20 = 1;
    61: op1_08_inv20 = 1;
    62: op1_08_inv20 = 1;
    64: op1_08_inv20 = 1;
    65: op1_08_inv20 = 1;
    67: op1_08_inv20 = 1;
    71: op1_08_inv20 = 1;
    75: op1_08_inv20 = 1;
    77: op1_08_inv20 = 1;
    80: op1_08_inv20 = 1;
    81: op1_08_inv20 = 1;
    86: op1_08_inv20 = 1;
    87: op1_08_inv20 = 1;
    90: op1_08_inv20 = 1;
    91: op1_08_inv20 = 1;
    92: op1_08_inv20 = 1;
    93: op1_08_inv20 = 1;
    94: op1_08_inv20 = 1;
    95: op1_08_inv20 = 1;
    96: op1_08_inv20 = 1;
    97: op1_08_inv20 = 1;
    default: op1_08_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in21 = reg_0348;
    6: op1_08_in21 = reg_0822;
    8: op1_08_in21 = reg_0055;
    9: op1_08_in21 = reg_0134;
    10: op1_08_in21 = imem04_in[107:104];
    11: op1_08_in21 = reg_0803;
    12: op1_08_in21 = imem04_in[7:4];
    13: op1_08_in21 = reg_0735;
    14: op1_08_in21 = reg_0649;
    15: op1_08_in21 = imem04_in[55:52];
    16: op1_08_in21 = reg_0177;
    17: op1_08_in21 = imem01_in[83:80];
    63: op1_08_in21 = imem01_in[83:80];
    79: op1_08_in21 = imem01_in[83:80];
    18: op1_08_in21 = reg_1028;
    19: op1_08_in21 = imem01_in[31:28];
    20: op1_08_in21 = reg_0709;
    21: op1_08_in21 = imem01_in[67:64];
    22: op1_08_in21 = reg_0626;
    23: op1_08_in21 = imem06_in[35:32];
    94: op1_08_in21 = imem06_in[35:32];
    24: op1_08_in21 = reg_0156;
    25: op1_08_in21 = imem07_in[91:88];
    44: op1_08_in21 = imem07_in[91:88];
    26: op1_08_in21 = imem03_in[39:36];
    74: op1_08_in21 = imem03_in[39:36];
    27: op1_08_in21 = reg_0431;
    28: op1_08_in21 = reg_0249;
    29: op1_08_in21 = reg_0799;
    31: op1_08_in21 = reg_1031;
    55: op1_08_in21 = reg_1031;
    32: op1_08_in21 = reg_1004;
    33: op1_08_in21 = reg_0047;
    35: op1_08_in21 = reg_0820;
    36: op1_08_in21 = reg_0373;
    37: op1_08_in21 = reg_0072;
    38: op1_08_in21 = reg_0046;
    39: op1_08_in21 = imem06_in[39:36];
    41: op1_08_in21 = reg_0426;
    42: op1_08_in21 = reg_0049;
    43: op1_08_in21 = reg_0066;
    45: op1_08_in21 = reg_0224;
    46: op1_08_in21 = imem03_in[71:68];
    47: op1_08_in21 = imem06_in[83:80];
    48: op1_08_in21 = imem01_in[99:96];
    49: op1_08_in21 = reg_0867;
    50: op1_08_in21 = imem01_in[111:108];
    52: op1_08_in21 = imem07_in[63:60];
    53: op1_08_in21 = reg_0178;
    56: op1_08_in21 = reg_0902;
    57: op1_08_in21 = reg_0087;
    58: op1_08_in21 = reg_0985;
    59: op1_08_in21 = imem03_in[95:92];
    60: op1_08_in21 = imem05_in[59:56];
    75: op1_08_in21 = imem05_in[59:56];
    61: op1_08_in21 = reg_0854;
    62: op1_08_in21 = reg_0698;
    64: op1_08_in21 = imem01_in[39:36];
    65: op1_08_in21 = reg_0088;
    66: op1_08_in21 = imem03_in[127:124];
    67: op1_08_in21 = imem03_in[127:124];
    68: op1_08_in21 = reg_0786;
    69: op1_08_in21 = reg_0168;
    70: op1_08_in21 = reg_0547;
    71: op1_08_in21 = reg_0524;
    72: op1_08_in21 = reg_0202;
    73: op1_08_in21 = reg_0012;
    76: op1_08_in21 = reg_0653;
    77: op1_08_in21 = imem07_in[111:108];
    80: op1_08_in21 = reg_0239;
    81: op1_08_in21 = reg_0824;
    82: op1_08_in21 = imem03_in[75:72];
    83: op1_08_in21 = reg_0234;
    84: op1_08_in21 = reg_0351;
    85: op1_08_in21 = imem03_in[11:8];
    86: op1_08_in21 = reg_0432;
    87: op1_08_in21 = reg_0183;
    88: op1_08_in21 = reg_0869;
    90: op1_08_in21 = reg_0624;
    91: op1_08_in21 = reg_0543;
    92: op1_08_in21 = reg_0346;
    93: op1_08_in21 = reg_0889;
    95: op1_08_in21 = reg_0675;
    96: op1_08_in21 = reg_0002;
    97: op1_08_in21 = imem05_in[67:64];
    default: op1_08_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv21 = 1;
    8: op1_08_inv21 = 1;
    9: op1_08_inv21 = 1;
    11: op1_08_inv21 = 1;
    12: op1_08_inv21 = 1;
    13: op1_08_inv21 = 1;
    16: op1_08_inv21 = 1;
    17: op1_08_inv21 = 1;
    21: op1_08_inv21 = 1;
    22: op1_08_inv21 = 1;
    24: op1_08_inv21 = 1;
    25: op1_08_inv21 = 1;
    27: op1_08_inv21 = 1;
    28: op1_08_inv21 = 1;
    29: op1_08_inv21 = 1;
    31: op1_08_inv21 = 1;
    33: op1_08_inv21 = 1;
    35: op1_08_inv21 = 1;
    36: op1_08_inv21 = 1;
    37: op1_08_inv21 = 1;
    39: op1_08_inv21 = 1;
    44: op1_08_inv21 = 1;
    45: op1_08_inv21 = 1;
    47: op1_08_inv21 = 1;
    48: op1_08_inv21 = 1;
    49: op1_08_inv21 = 1;
    50: op1_08_inv21 = 1;
    52: op1_08_inv21 = 1;
    55: op1_08_inv21 = 1;
    57: op1_08_inv21 = 1;
    58: op1_08_inv21 = 1;
    60: op1_08_inv21 = 1;
    62: op1_08_inv21 = 1;
    63: op1_08_inv21 = 1;
    65: op1_08_inv21 = 1;
    66: op1_08_inv21 = 1;
    68: op1_08_inv21 = 1;
    69: op1_08_inv21 = 1;
    72: op1_08_inv21 = 1;
    77: op1_08_inv21 = 1;
    80: op1_08_inv21 = 1;
    81: op1_08_inv21 = 1;
    83: op1_08_inv21 = 1;
    87: op1_08_inv21 = 1;
    88: op1_08_inv21 = 1;
    93: op1_08_inv21 = 1;
    95: op1_08_inv21 = 1;
    default: op1_08_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in22 = reg_0379;
    93: op1_08_in22 = reg_0379;
    6: op1_08_in22 = reg_0828;
    45: op1_08_in22 = reg_0828;
    8: op1_08_in22 = reg_0060;
    59: op1_08_in22 = reg_0060;
    9: op1_08_in22 = reg_1020;
    10: op1_08_in22 = reg_0536;
    11: op1_08_in22 = reg_0805;
    18: op1_08_in22 = reg_0805;
    76: op1_08_in22 = reg_0805;
    12: op1_08_in22 = imem04_in[27:24];
    13: op1_08_in22 = reg_0248;
    14: op1_08_in22 = reg_0663;
    15: op1_08_in22 = imem04_in[59:56];
    16: op1_08_in22 = reg_0164;
    17: op1_08_in22 = imem01_in[87:84];
    19: op1_08_in22 = imem01_in[59:56];
    20: op1_08_in22 = reg_0706;
    21: op1_08_in22 = imem01_in[123:120];
    22: op1_08_in22 = reg_0611;
    23: op1_08_in22 = imem06_in[103:100];
    24: op1_08_in22 = reg_0143;
    25: op1_08_in22 = imem07_in[95:92];
    26: op1_08_in22 = imem03_in[99:96];
    46: op1_08_in22 = imem03_in[99:96];
    27: op1_08_in22 = reg_0172;
    28: op1_08_in22 = reg_0496;
    29: op1_08_in22 = reg_0798;
    31: op1_08_in22 = reg_1041;
    32: op1_08_in22 = reg_0265;
    33: op1_08_in22 = reg_0738;
    35: op1_08_in22 = reg_0844;
    36: op1_08_in22 = reg_0991;
    37: op1_08_in22 = reg_0748;
    38: op1_08_in22 = reg_0396;
    39: op1_08_in22 = imem06_in[55:52];
    41: op1_08_in22 = reg_0434;
    42: op1_08_in22 = imem03_in[71:68];
    43: op1_08_in22 = reg_0302;
    44: op1_08_in22 = reg_0728;
    47: op1_08_in22 = imem06_in[95:92];
    48: op1_08_in22 = reg_1039;
    49: op1_08_in22 = reg_0077;
    50: op1_08_in22 = reg_0918;
    52: op1_08_in22 = imem07_in[79:76];
    55: op1_08_in22 = reg_0521;
    56: op1_08_in22 = reg_0354;
    57: op1_08_in22 = reg_0644;
    58: op1_08_in22 = reg_0998;
    60: op1_08_in22 = imem05_in[63:60];
    61: op1_08_in22 = reg_0542;
    62: op1_08_in22 = reg_0222;
    63: op1_08_in22 = imem01_in[107:104];
    64: op1_08_in22 = imem01_in[43:40];
    65: op1_08_in22 = reg_0792;
    66: op1_08_in22 = reg_0012;
    67: op1_08_in22 = reg_0012;
    68: op1_08_in22 = reg_0145;
    70: op1_08_in22 = reg_0576;
    71: op1_08_in22 = reg_0296;
    72: op1_08_in22 = imem01_in[79:76];
    73: op1_08_in22 = reg_0307;
    74: op1_08_in22 = imem03_in[91:88];
    82: op1_08_in22 = imem03_in[91:88];
    75: op1_08_in22 = imem05_in[103:100];
    77: op1_08_in22 = imem07_in[123:120];
    79: op1_08_in22 = imem01_in[103:100];
    80: op1_08_in22 = reg_1008;
    81: op1_08_in22 = imem05_in[3:0];
    83: op1_08_in22 = reg_0869;
    84: op1_08_in22 = reg_0025;
    85: op1_08_in22 = imem03_in[35:32];
    86: op1_08_in22 = reg_0332;
    87: op1_08_in22 = reg_0449;
    88: op1_08_in22 = reg_0832;
    90: op1_08_in22 = reg_0367;
    91: op1_08_in22 = reg_0305;
    92: op1_08_in22 = reg_0823;
    94: op1_08_in22 = imem06_in[43:40];
    95: op1_08_in22 = reg_0152;
    96: op1_08_in22 = reg_0047;
    97: op1_08_in22 = imem05_in[79:76];
    default: op1_08_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv22 = 1;
    8: op1_08_inv22 = 1;
    9: op1_08_inv22 = 1;
    11: op1_08_inv22 = 1;
    12: op1_08_inv22 = 1;
    14: op1_08_inv22 = 1;
    15: op1_08_inv22 = 1;
    17: op1_08_inv22 = 1;
    18: op1_08_inv22 = 1;
    20: op1_08_inv22 = 1;
    22: op1_08_inv22 = 1;
    24: op1_08_inv22 = 1;
    28: op1_08_inv22 = 1;
    31: op1_08_inv22 = 1;
    39: op1_08_inv22 = 1;
    41: op1_08_inv22 = 1;
    43: op1_08_inv22 = 1;
    47: op1_08_inv22 = 1;
    58: op1_08_inv22 = 1;
    59: op1_08_inv22 = 1;
    60: op1_08_inv22 = 1;
    63: op1_08_inv22 = 1;
    64: op1_08_inv22 = 1;
    66: op1_08_inv22 = 1;
    68: op1_08_inv22 = 1;
    71: op1_08_inv22 = 1;
    80: op1_08_inv22 = 1;
    81: op1_08_inv22 = 1;
    86: op1_08_inv22 = 1;
    88: op1_08_inv22 = 1;
    90: op1_08_inv22 = 1;
    93: op1_08_inv22 = 1;
    94: op1_08_inv22 = 1;
    96: op1_08_inv22 = 1;
    default: op1_08_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in23 = reg_0349;
    6: op1_08_in23 = reg_0819;
    8: op1_08_in23 = imem03_in[19:16];
    9: op1_08_in23 = reg_0914;
    10: op1_08_in23 = reg_0557;
    11: op1_08_in23 = imem07_in[55:52];
    12: op1_08_in23 = imem04_in[75:72];
    13: op1_08_in23 = reg_0238;
    14: op1_08_in23 = reg_0325;
    76: op1_08_in23 = reg_0325;
    15: op1_08_in23 = reg_0544;
    16: op1_08_in23 = reg_0185;
    17: op1_08_in23 = imem01_in[119:116];
    18: op1_08_in23 = reg_0798;
    19: op1_08_in23 = imem01_in[63:60];
    20: op1_08_in23 = reg_0441;
    21: op1_08_in23 = reg_0239;
    22: op1_08_in23 = reg_0622;
    23: op1_08_in23 = imem06_in[127:124];
    24: op1_08_in23 = reg_0139;
    25: op1_08_in23 = imem07_in[103:100];
    26: op1_08_in23 = reg_0597;
    27: op1_08_in23 = reg_0166;
    28: op1_08_in23 = reg_0230;
    29: op1_08_in23 = imem07_in[19:16];
    31: op1_08_in23 = reg_1038;
    32: op1_08_in23 = reg_0937;
    33: op1_08_in23 = imem05_in[59:56];
    35: op1_08_in23 = reg_0980;
    58: op1_08_in23 = reg_0980;
    36: op1_08_in23 = reg_0999;
    37: op1_08_in23 = reg_0864;
    38: op1_08_in23 = reg_0824;
    39: op1_08_in23 = imem06_in[91:88];
    41: op1_08_in23 = reg_0427;
    42: op1_08_in23 = imem03_in[119:116];
    43: op1_08_in23 = reg_0068;
    44: op1_08_in23 = reg_0719;
    45: op1_08_in23 = reg_0236;
    46: op1_08_in23 = imem03_in[115:112];
    47: op1_08_in23 = imem06_in[99:96];
    48: op1_08_in23 = reg_0522;
    49: op1_08_in23 = reg_0884;
    50: op1_08_in23 = reg_0928;
    52: op1_08_in23 = imem07_in[83:80];
    55: op1_08_in23 = reg_0925;
    56: op1_08_in23 = reg_1017;
    57: op1_08_in23 = reg_0335;
    59: op1_08_in23 = reg_0760;
    60: op1_08_in23 = imem05_in[87:84];
    97: op1_08_in23 = imem05_in[87:84];
    61: op1_08_in23 = reg_0070;
    62: op1_08_in23 = reg_0241;
    63: op1_08_in23 = imem01_in[111:108];
    64: op1_08_in23 = imem01_in[67:64];
    65: op1_08_in23 = reg_0814;
    66: op1_08_in23 = reg_0357;
    67: op1_08_in23 = reg_0099;
    68: op1_08_in23 = reg_0142;
    70: op1_08_in23 = imem03_in[111:108];
    71: op1_08_in23 = reg_0074;
    72: op1_08_in23 = imem01_in[83:80];
    73: op1_08_in23 = reg_0590;
    74: op1_08_in23 = imem03_in[103:100];
    75: op1_08_in23 = imem05_in[127:124];
    77: op1_08_in23 = reg_0712;
    79: op1_08_in23 = imem01_in[115:112];
    80: op1_08_in23 = reg_0051;
    81: op1_08_in23 = imem05_in[7:4];
    82: op1_08_in23 = reg_0060;
    83: op1_08_in23 = reg_0604;
    84: op1_08_in23 = reg_0626;
    85: op1_08_in23 = imem03_in[87:84];
    86: op1_08_in23 = imem05_in[19:16];
    87: op1_08_in23 = reg_0690;
    88: op1_08_in23 = reg_0116;
    90: op1_08_in23 = reg_0000;
    91: op1_08_in23 = reg_0887;
    92: op1_08_in23 = reg_0596;
    93: op1_08_in23 = reg_1028;
    94: op1_08_in23 = imem06_in[47:44];
    95: op1_08_in23 = reg_0023;
    96: op1_08_in23 = reg_0599;
    default: op1_08_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    11: op1_08_inv23 = 1;
    12: op1_08_inv23 = 1;
    13: op1_08_inv23 = 1;
    16: op1_08_inv23 = 1;
    19: op1_08_inv23 = 1;
    20: op1_08_inv23 = 1;
    25: op1_08_inv23 = 1;
    27: op1_08_inv23 = 1;
    29: op1_08_inv23 = 1;
    33: op1_08_inv23 = 1;
    36: op1_08_inv23 = 1;
    38: op1_08_inv23 = 1;
    41: op1_08_inv23 = 1;
    42: op1_08_inv23 = 1;
    44: op1_08_inv23 = 1;
    52: op1_08_inv23 = 1;
    58: op1_08_inv23 = 1;
    59: op1_08_inv23 = 1;
    60: op1_08_inv23 = 1;
    62: op1_08_inv23 = 1;
    66: op1_08_inv23 = 1;
    67: op1_08_inv23 = 1;
    71: op1_08_inv23 = 1;
    72: op1_08_inv23 = 1;
    74: op1_08_inv23 = 1;
    76: op1_08_inv23 = 1;
    77: op1_08_inv23 = 1;
    79: op1_08_inv23 = 1;
    80: op1_08_inv23 = 1;
    81: op1_08_inv23 = 1;
    84: op1_08_inv23 = 1;
    85: op1_08_inv23 = 1;
    88: op1_08_inv23 = 1;
    91: op1_08_inv23 = 1;
    94: op1_08_inv23 = 1;
    96: op1_08_inv23 = 1;
    default: op1_08_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in24 = reg_0403;
    6: op1_08_in24 = reg_0832;
    8: op1_08_in24 = imem03_in[23:20];
    9: op1_08_in24 = reg_0020;
    10: op1_08_in24 = reg_0534;
    11: op1_08_in24 = imem07_in[95:92];
    12: op1_08_in24 = imem04_in[87:84];
    13: op1_08_in24 = reg_0508;
    14: op1_08_in24 = reg_0326;
    15: op1_08_in24 = reg_0530;
    16: op1_08_in24 = reg_0158;
    17: op1_08_in24 = reg_0240;
    59: op1_08_in24 = reg_0240;
    18: op1_08_in24 = imem07_in[19:16];
    19: op1_08_in24 = reg_1051;
    20: op1_08_in24 = reg_0429;
    21: op1_08_in24 = reg_1050;
    22: op1_08_in24 = reg_0402;
    23: op1_08_in24 = reg_0629;
    24: op1_08_in24 = reg_0129;
    25: op1_08_in24 = reg_0727;
    26: op1_08_in24 = reg_0581;
    27: op1_08_in24 = reg_0184;
    28: op1_08_in24 = reg_0830;
    29: op1_08_in24 = imem07_in[67:64];
    31: op1_08_in24 = reg_0111;
    56: op1_08_in24 = reg_0111;
    32: op1_08_in24 = reg_0282;
    33: op1_08_in24 = imem05_in[115:112];
    35: op1_08_in24 = imem04_in[35:32];
    36: op1_08_in24 = reg_0974;
    37: op1_08_in24 = reg_0021;
    38: op1_08_in24 = reg_0847;
    39: op1_08_in24 = imem06_in[107:104];
    41: op1_08_in24 = reg_0437;
    42: op1_08_in24 = reg_1008;
    43: op1_08_in24 = reg_0584;
    44: op1_08_in24 = reg_0710;
    45: op1_08_in24 = reg_0274;
    46: op1_08_in24 = reg_0535;
    47: op1_08_in24 = reg_0915;
    48: op1_08_in24 = reg_0869;
    49: op1_08_in24 = imem03_in[7:4];
    50: op1_08_in24 = reg_1044;
    52: op1_08_in24 = imem07_in[99:96];
    55: op1_08_in24 = reg_0232;
    57: op1_08_in24 = reg_0772;
    58: op1_08_in24 = reg_0978;
    60: op1_08_in24 = reg_1021;
    61: op1_08_in24 = reg_0970;
    62: op1_08_in24 = reg_0386;
    63: op1_08_in24 = reg_0786;
    64: op1_08_in24 = imem01_in[115:112];
    65: op1_08_in24 = reg_0049;
    66: op1_08_in24 = reg_0580;
    67: op1_08_in24 = reg_0357;
    68: op1_08_in24 = reg_0134;
    70: op1_08_in24 = imem03_in[115:112];
    85: op1_08_in24 = imem03_in[115:112];
    71: op1_08_in24 = reg_0243;
    72: op1_08_in24 = reg_1042;
    73: op1_08_in24 = reg_0576;
    74: op1_08_in24 = reg_0345;
    75: op1_08_in24 = reg_0142;
    76: op1_08_in24 = reg_0315;
    77: op1_08_in24 = reg_0265;
    79: op1_08_in24 = reg_0122;
    80: op1_08_in24 = reg_0377;
    81: op1_08_in24 = imem05_in[11:8];
    82: op1_08_in24 = reg_0620;
    83: op1_08_in24 = reg_0216;
    84: op1_08_in24 = reg_0817;
    86: op1_08_in24 = imem05_in[27:24];
    87: op1_08_in24 = reg_0371;
    88: op1_08_in24 = reg_1033;
    90: op1_08_in24 = reg_0681;
    91: op1_08_in24 = reg_0765;
    92: op1_08_in24 = reg_0773;
    93: op1_08_in24 = reg_0698;
    94: op1_08_in24 = imem06_in[55:52];
    95: op1_08_in24 = reg_0145;
    96: op1_08_in24 = reg_0838;
    97: op1_08_in24 = imem05_in[107:104];
    default: op1_08_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv24 = 1;
    9: op1_08_inv24 = 1;
    11: op1_08_inv24 = 1;
    12: op1_08_inv24 = 1;
    15: op1_08_inv24 = 1;
    16: op1_08_inv24 = 1;
    18: op1_08_inv24 = 1;
    23: op1_08_inv24 = 1;
    27: op1_08_inv24 = 1;
    29: op1_08_inv24 = 1;
    35: op1_08_inv24 = 1;
    37: op1_08_inv24 = 1;
    38: op1_08_inv24 = 1;
    39: op1_08_inv24 = 1;
    42: op1_08_inv24 = 1;
    47: op1_08_inv24 = 1;
    48: op1_08_inv24 = 1;
    49: op1_08_inv24 = 1;
    50: op1_08_inv24 = 1;
    52: op1_08_inv24 = 1;
    57: op1_08_inv24 = 1;
    59: op1_08_inv24 = 1;
    60: op1_08_inv24 = 1;
    61: op1_08_inv24 = 1;
    62: op1_08_inv24 = 1;
    63: op1_08_inv24 = 1;
    65: op1_08_inv24 = 1;
    66: op1_08_inv24 = 1;
    70: op1_08_inv24 = 1;
    71: op1_08_inv24 = 1;
    73: op1_08_inv24 = 1;
    76: op1_08_inv24 = 1;
    81: op1_08_inv24 = 1;
    82: op1_08_inv24 = 1;
    84: op1_08_inv24 = 1;
    85: op1_08_inv24 = 1;
    87: op1_08_inv24 = 1;
    88: op1_08_inv24 = 1;
    91: op1_08_inv24 = 1;
    92: op1_08_inv24 = 1;
    94: op1_08_inv24 = 1;
    default: op1_08_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in25 = reg_0367;
    6: op1_08_in25 = imem05_in[19:16];
    8: op1_08_in25 = imem03_in[51:48];
    9: op1_08_in25 = reg_0864;
    10: op1_08_in25 = reg_0555;
    11: op1_08_in25 = imem07_in[103:100];
    29: op1_08_in25 = imem07_in[103:100];
    12: op1_08_in25 = imem04_in[127:124];
    13: op1_08_in25 = reg_0905;
    14: op1_08_in25 = reg_0359;
    15: op1_08_in25 = reg_0553;
    17: op1_08_in25 = reg_0508;
    95: op1_08_in25 = reg_0508;
    18: op1_08_in25 = imem07_in[23:20];
    19: op1_08_in25 = reg_0511;
    20: op1_08_in25 = reg_0428;
    21: op1_08_in25 = reg_0226;
    22: op1_08_in25 = reg_0379;
    23: op1_08_in25 = reg_0616;
    24: op1_08_in25 = reg_0141;
    25: op1_08_in25 = reg_0175;
    26: op1_08_in25 = reg_0590;
    28: op1_08_in25 = reg_0216;
    31: op1_08_in25 = reg_0116;
    32: op1_08_in25 = reg_0912;
    33: op1_08_in25 = reg_0973;
    72: op1_08_in25 = reg_0973;
    35: op1_08_in25 = imem04_in[43:40];
    36: op1_08_in25 = reg_0977;
    37: op1_08_in25 = imem05_in[3:0];
    38: op1_08_in25 = reg_0923;
    39: op1_08_in25 = imem06_in[127:124];
    41: op1_08_in25 = reg_0438;
    42: op1_08_in25 = reg_1019;
    43: op1_08_in25 = reg_0072;
    44: op1_08_in25 = reg_0731;
    45: op1_08_in25 = reg_0238;
    46: op1_08_in25 = reg_0571;
    47: op1_08_in25 = reg_0781;
    48: op1_08_in25 = reg_1031;
    83: op1_08_in25 = reg_1031;
    49: op1_08_in25 = imem03_in[47:44];
    50: op1_08_in25 = reg_0503;
    52: op1_08_in25 = imem07_in[107:104];
    55: op1_08_in25 = reg_0109;
    56: op1_08_in25 = reg_0283;
    57: op1_08_in25 = reg_0482;
    58: op1_08_in25 = reg_0999;
    59: op1_08_in25 = reg_0765;
    60: op1_08_in25 = reg_0255;
    61: op1_08_in25 = reg_0966;
    62: op1_08_in25 = reg_0264;
    63: op1_08_in25 = reg_0779;
    64: op1_08_in25 = reg_0928;
    65: op1_08_in25 = reg_0840;
    66: op1_08_in25 = reg_0307;
    67: op1_08_in25 = reg_0547;
    68: op1_08_in25 = imem06_in[11:8];
    70: op1_08_in25 = reg_0982;
    71: op1_08_in25 = reg_0542;
    73: op1_08_in25 = reg_0239;
    74: op1_08_in25 = reg_0580;
    75: op1_08_in25 = reg_0319;
    76: op1_08_in25 = reg_0419;
    77: op1_08_in25 = reg_0628;
    79: op1_08_in25 = reg_1014;
    80: op1_08_in25 = reg_0767;
    81: op1_08_in25 = imem05_in[51:48];
    82: op1_08_in25 = reg_0345;
    84: op1_08_in25 = reg_0735;
    85: op1_08_in25 = reg_0012;
    86: op1_08_in25 = imem05_in[35:32];
    87: op1_08_in25 = reg_0184;
    88: op1_08_in25 = reg_0114;
    90: op1_08_in25 = reg_0984;
    91: op1_08_in25 = reg_0418;
    92: op1_08_in25 = reg_0051;
    93: op1_08_in25 = reg_0822;
    94: op1_08_in25 = imem06_in[83:80];
    96: op1_08_in25 = reg_0539;
    97: op1_08_in25 = imem05_in[123:120];
    default: op1_08_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv25 = 1;
    8: op1_08_inv25 = 1;
    9: op1_08_inv25 = 1;
    11: op1_08_inv25 = 1;
    12: op1_08_inv25 = 1;
    13: op1_08_inv25 = 1;
    14: op1_08_inv25 = 1;
    17: op1_08_inv25 = 1;
    19: op1_08_inv25 = 1;
    21: op1_08_inv25 = 1;
    23: op1_08_inv25 = 1;
    25: op1_08_inv25 = 1;
    29: op1_08_inv25 = 1;
    32: op1_08_inv25 = 1;
    37: op1_08_inv25 = 1;
    38: op1_08_inv25 = 1;
    39: op1_08_inv25 = 1;
    41: op1_08_inv25 = 1;
    44: op1_08_inv25 = 1;
    47: op1_08_inv25 = 1;
    55: op1_08_inv25 = 1;
    56: op1_08_inv25 = 1;
    57: op1_08_inv25 = 1;
    59: op1_08_inv25 = 1;
    60: op1_08_inv25 = 1;
    63: op1_08_inv25 = 1;
    67: op1_08_inv25 = 1;
    68: op1_08_inv25 = 1;
    72: op1_08_inv25 = 1;
    73: op1_08_inv25 = 1;
    74: op1_08_inv25 = 1;
    75: op1_08_inv25 = 1;
    79: op1_08_inv25 = 1;
    80: op1_08_inv25 = 1;
    84: op1_08_inv25 = 1;
    85: op1_08_inv25 = 1;
    86: op1_08_inv25 = 1;
    90: op1_08_inv25 = 1;
    94: op1_08_inv25 = 1;
    95: op1_08_inv25 = 1;
    96: op1_08_inv25 = 1;
    97: op1_08_inv25 = 1;
    default: op1_08_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in26 = reg_0380;
    6: op1_08_in26 = imem05_in[67:64];
    8: op1_08_in26 = imem03_in[63:60];
    9: op1_08_in26 = reg_0630;
    10: op1_08_in26 = reg_0558;
    11: op1_08_in26 = imem07_in[107:104];
    12: op1_08_in26 = reg_0540;
    13: op1_08_in26 = reg_1043;
    14: op1_08_in26 = reg_0339;
    15: op1_08_in26 = reg_0529;
    17: op1_08_in26 = reg_1042;
    21: op1_08_in26 = reg_1042;
    18: op1_08_in26 = imem07_in[27:24];
    19: op1_08_in26 = reg_1049;
    20: op1_08_in26 = reg_0446;
    22: op1_08_in26 = reg_0372;
    23: op1_08_in26 = reg_0618;
    24: op1_08_in26 = imem06_in[63:60];
    25: op1_08_in26 = reg_0165;
    26: op1_08_in26 = reg_0370;
    28: op1_08_in26 = reg_0871;
    29: op1_08_in26 = imem07_in[119:116];
    31: op1_08_in26 = imem02_in[79:76];
    32: op1_08_in26 = reg_0055;
    33: op1_08_in26 = reg_0954;
    35: op1_08_in26 = imem04_in[59:56];
    36: op1_08_in26 = reg_0975;
    37: op1_08_in26 = imem05_in[7:4];
    38: op1_08_in26 = reg_0833;
    39: op1_08_in26 = reg_0348;
    41: op1_08_in26 = reg_0435;
    42: op1_08_in26 = reg_0389;
    43: op1_08_in26 = reg_0054;
    44: op1_08_in26 = reg_0723;
    45: op1_08_in26 = reg_0520;
    46: op1_08_in26 = reg_0357;
    47: op1_08_in26 = reg_0403;
    48: op1_08_in26 = reg_0354;
    49: op1_08_in26 = imem03_in[51:48];
    50: op1_08_in26 = reg_0274;
    52: op1_08_in26 = reg_0728;
    55: op1_08_in26 = imem02_in[15:12];
    56: op1_08_in26 = imem02_in[3:0];
    57: op1_08_in26 = reg_0085;
    58: op1_08_in26 = reg_0988;
    59: op1_08_in26 = reg_0836;
    60: op1_08_in26 = reg_0866;
    61: op1_08_in26 = reg_0782;
    62: op1_08_in26 = reg_0633;
    63: op1_08_in26 = reg_0928;
    64: op1_08_in26 = reg_0236;
    65: op1_08_in26 = reg_0310;
    66: op1_08_in26 = reg_0322;
    67: op1_08_in26 = reg_0346;
    68: op1_08_in26 = imem06_in[15:12];
    70: op1_08_in26 = reg_0984;
    71: op1_08_in26 = reg_0070;
    72: op1_08_in26 = reg_0831;
    73: op1_08_in26 = reg_0230;
    74: op1_08_in26 = reg_0327;
    75: op1_08_in26 = reg_0448;
    76: op1_08_in26 = reg_0868;
    77: op1_08_in26 = reg_0250;
    79: op1_08_in26 = reg_1044;
    80: op1_08_in26 = reg_0981;
    81: op1_08_in26 = imem05_in[63:60];
    82: op1_08_in26 = reg_0099;
    83: op1_08_in26 = reg_0737;
    84: op1_08_in26 = reg_0384;
    85: op1_08_in26 = reg_1007;
    86: op1_08_in26 = imem05_in[87:84];
    88: op1_08_in26 = reg_0103;
    90: op1_08_in26 = reg_0635;
    91: op1_08_in26 = reg_0081;
    92: op1_08_in26 = reg_0385;
    93: op1_08_in26 = reg_0811;
    94: op1_08_in26 = imem06_in[103:100];
    95: op1_08_in26 = reg_0146;
    97: op1_08_in26 = reg_1021;
    default: op1_08_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv26 = 1;
    6: op1_08_inv26 = 1;
    8: op1_08_inv26 = 1;
    9: op1_08_inv26 = 1;
    10: op1_08_inv26 = 1;
    12: op1_08_inv26 = 1;
    15: op1_08_inv26 = 1;
    18: op1_08_inv26 = 1;
    19: op1_08_inv26 = 1;
    23: op1_08_inv26 = 1;
    24: op1_08_inv26 = 1;
    31: op1_08_inv26 = 1;
    32: op1_08_inv26 = 1;
    35: op1_08_inv26 = 1;
    37: op1_08_inv26 = 1;
    39: op1_08_inv26 = 1;
    41: op1_08_inv26 = 1;
    42: op1_08_inv26 = 1;
    46: op1_08_inv26 = 1;
    48: op1_08_inv26 = 1;
    50: op1_08_inv26 = 1;
    52: op1_08_inv26 = 1;
    55: op1_08_inv26 = 1;
    56: op1_08_inv26 = 1;
    62: op1_08_inv26 = 1;
    65: op1_08_inv26 = 1;
    66: op1_08_inv26 = 1;
    67: op1_08_inv26 = 1;
    68: op1_08_inv26 = 1;
    70: op1_08_inv26 = 1;
    72: op1_08_inv26 = 1;
    74: op1_08_inv26 = 1;
    77: op1_08_inv26 = 1;
    79: op1_08_inv26 = 1;
    82: op1_08_inv26 = 1;
    88: op1_08_inv26 = 1;
    90: op1_08_inv26 = 1;
    94: op1_08_inv26 = 1;
    95: op1_08_inv26 = 1;
    97: op1_08_inv26 = 1;
    default: op1_08_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in27 = reg_0026;
    6: op1_08_in27 = imem05_in[75:72];
    8: op1_08_in27 = reg_0579;
    9: op1_08_in27 = reg_0624;
    10: op1_08_in27 = reg_0559;
    11: op1_08_in27 = imem07_in[115:112];
    12: op1_08_in27 = reg_0304;
    13: op1_08_in27 = reg_1033;
    14: op1_08_in27 = reg_0346;
    46: op1_08_in27 = reg_0346;
    15: op1_08_in27 = reg_0537;
    17: op1_08_in27 = reg_1031;
    18: op1_08_in27 = imem07_in[31:28];
    19: op1_08_in27 = reg_1056;
    79: op1_08_in27 = reg_1056;
    20: op1_08_in27 = reg_0175;
    21: op1_08_in27 = reg_1043;
    22: op1_08_in27 = reg_0407;
    23: op1_08_in27 = reg_0402;
    24: op1_08_in27 = imem06_in[95:92];
    25: op1_08_in27 = reg_0179;
    26: op1_08_in27 = reg_0369;
    28: op1_08_in27 = reg_1017;
    29: op1_08_in27 = reg_0714;
    31: op1_08_in27 = imem02_in[83:80];
    32: op1_08_in27 = reg_0048;
    33: op1_08_in27 = reg_0950;
    35: op1_08_in27 = imem04_in[63:60];
    36: op1_08_in27 = imem04_in[43:40];
    37: op1_08_in27 = imem05_in[39:36];
    38: op1_08_in27 = reg_0807;
    39: op1_08_in27 = reg_0356;
    41: op1_08_in27 = reg_0431;
    42: op1_08_in27 = reg_0509;
    43: op1_08_in27 = reg_0738;
    44: op1_08_in27 = reg_0700;
    45: op1_08_in27 = reg_0737;
    47: op1_08_in27 = reg_0783;
    48: op1_08_in27 = reg_0906;
    49: op1_08_in27 = imem03_in[67:64];
    50: op1_08_in27 = reg_0238;
    52: op1_08_in27 = reg_0720;
    55: op1_08_in27 = imem02_in[31:28];
    56: op1_08_in27 = imem02_in[7:4];
    57: op1_08_in27 = reg_0086;
    58: op1_08_in27 = reg_0990;
    59: op1_08_in27 = reg_0246;
    60: op1_08_in27 = reg_0675;
    75: op1_08_in27 = reg_0675;
    61: op1_08_in27 = reg_0954;
    62: op1_08_in27 = reg_0349;
    63: op1_08_in27 = reg_0218;
    64: op1_08_in27 = reg_0871;
    65: op1_08_in27 = reg_0291;
    66: op1_08_in27 = reg_0434;
    67: op1_08_in27 = reg_0543;
    68: op1_08_in27 = imem06_in[39:36];
    70: op1_08_in27 = reg_0993;
    71: op1_08_in27 = reg_0332;
    72: op1_08_in27 = reg_0862;
    73: op1_08_in27 = reg_0982;
    74: op1_08_in27 = reg_0322;
    76: op1_08_in27 = reg_0640;
    77: op1_08_in27 = reg_0047;
    80: op1_08_in27 = reg_0977;
    81: op1_08_in27 = imem05_in[83:80];
    82: op1_08_in27 = reg_1007;
    83: op1_08_in27 = reg_0610;
    84: op1_08_in27 = reg_0895;
    85: op1_08_in27 = reg_0046;
    86: op1_08_in27 = reg_0636;
    88: op1_08_in27 = reg_0745;
    90: op1_08_in27 = reg_0245;
    91: op1_08_in27 = reg_0424;
    92: op1_08_in27 = reg_0233;
    93: op1_08_in27 = reg_0169;
    94: op1_08_in27 = imem06_in[115:112];
    95: op1_08_in27 = reg_0851;
    97: op1_08_in27 = reg_0136;
    default: op1_08_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv27 = 1;
    6: op1_08_inv27 = 1;
    8: op1_08_inv27 = 1;
    9: op1_08_inv27 = 1;
    11: op1_08_inv27 = 1;
    12: op1_08_inv27 = 1;
    13: op1_08_inv27 = 1;
    14: op1_08_inv27 = 1;
    15: op1_08_inv27 = 1;
    18: op1_08_inv27 = 1;
    19: op1_08_inv27 = 1;
    20: op1_08_inv27 = 1;
    21: op1_08_inv27 = 1;
    22: op1_08_inv27 = 1;
    23: op1_08_inv27 = 1;
    25: op1_08_inv27 = 1;
    26: op1_08_inv27 = 1;
    28: op1_08_inv27 = 1;
    32: op1_08_inv27 = 1;
    37: op1_08_inv27 = 1;
    42: op1_08_inv27 = 1;
    44: op1_08_inv27 = 1;
    46: op1_08_inv27 = 1;
    47: op1_08_inv27 = 1;
    49: op1_08_inv27 = 1;
    50: op1_08_inv27 = 1;
    55: op1_08_inv27 = 1;
    59: op1_08_inv27 = 1;
    60: op1_08_inv27 = 1;
    62: op1_08_inv27 = 1;
    64: op1_08_inv27 = 1;
    67: op1_08_inv27 = 1;
    68: op1_08_inv27 = 1;
    70: op1_08_inv27 = 1;
    72: op1_08_inv27 = 1;
    74: op1_08_inv27 = 1;
    76: op1_08_inv27 = 1;
    77: op1_08_inv27 = 1;
    79: op1_08_inv27 = 1;
    84: op1_08_inv27 = 1;
    86: op1_08_inv27 = 1;
    88: op1_08_inv27 = 1;
    92: op1_08_inv27 = 1;
    97: op1_08_inv27 = 1;
    default: op1_08_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in28 = reg_0020;
    6: op1_08_in28 = imem05_in[103:100];
    8: op1_08_in28 = reg_0569;
    9: op1_08_in28 = reg_0633;
    10: op1_08_in28 = reg_0531;
    11: op1_08_in28 = imem07_in[127:124];
    12: op1_08_in28 = reg_0279;
    13: op1_08_in28 = reg_0830;
    14: op1_08_in28 = reg_0353;
    15: op1_08_in28 = reg_0549;
    17: op1_08_in28 = reg_1036;
    18: op1_08_in28 = imem07_in[67:64];
    19: op1_08_in28 = reg_0220;
    20: op1_08_in28 = reg_0180;
    21: op1_08_in28 = reg_0216;
    22: op1_08_in28 = reg_0403;
    23: op1_08_in28 = reg_0344;
    24: op1_08_in28 = imem06_in[127:124];
    25: op1_08_in28 = reg_0161;
    26: op1_08_in28 = reg_0377;
    28: op1_08_in28 = reg_1038;
    29: op1_08_in28 = reg_0711;
    31: op1_08_in28 = imem02_in[87:84];
    32: op1_08_in28 = reg_0733;
    33: op1_08_in28 = reg_0951;
    35: op1_08_in28 = imem04_in[71:68];
    36: op1_08_in28 = imem04_in[55:52];
    37: op1_08_in28 = imem05_in[63:60];
    38: op1_08_in28 = reg_0513;
    39: op1_08_in28 = reg_0381;
    41: op1_08_in28 = reg_0166;
    42: op1_08_in28 = reg_0807;
    67: op1_08_in28 = reg_0807;
    43: op1_08_in28 = reg_0777;
    44: op1_08_in28 = reg_0727;
    45: op1_08_in28 = reg_1041;
    46: op1_08_in28 = reg_0396;
    47: op1_08_in28 = reg_0356;
    48: op1_08_in28 = reg_0123;
    49: op1_08_in28 = imem03_in[71:68];
    50: op1_08_in28 = reg_0285;
    52: op1_08_in28 = reg_0721;
    55: op1_08_in28 = imem02_in[79:76];
    56: op1_08_in28 = imem02_in[67:64];
    57: op1_08_in28 = reg_0084;
    58: op1_08_in28 = reg_0997;
    59: op1_08_in28 = reg_0991;
    60: op1_08_in28 = reg_0688;
    75: op1_08_in28 = reg_0688;
    61: op1_08_in28 = reg_0260;
    62: op1_08_in28 = imem07_in[3:0];
    63: op1_08_in28 = reg_1056;
    64: op1_08_in28 = reg_0496;
    65: op1_08_in28 = reg_0079;
    66: op1_08_in28 = reg_0346;
    68: op1_08_in28 = imem06_in[103:100];
    70: op1_08_in28 = reg_0999;
    71: op1_08_in28 = reg_0856;
    72: op1_08_in28 = reg_0869;
    73: op1_08_in28 = reg_0980;
    74: op1_08_in28 = reg_0585;
    76: op1_08_in28 = reg_0162;
    77: op1_08_in28 = reg_0175;
    79: op1_08_in28 = reg_0592;
    80: op1_08_in28 = imem04_in[31:28];
    81: op1_08_in28 = imem05_in[127:124];
    82: op1_08_in28 = reg_0307;
    83: op1_08_in28 = reg_0925;
    84: op1_08_in28 = reg_0392;
    85: op1_08_in28 = reg_0661;
    86: op1_08_in28 = reg_0866;
    88: op1_08_in28 = imem02_in[19:16];
    90: op1_08_in28 = reg_0974;
    91: op1_08_in28 = reg_0664;
    92: op1_08_in28 = reg_0266;
    93: op1_08_in28 = reg_0628;
    94: op1_08_in28 = reg_0660;
    95: op1_08_in28 = reg_0657;
    97: op1_08_in28 = reg_0954;
    default: op1_08_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv28 = 1;
    8: op1_08_inv28 = 1;
    13: op1_08_inv28 = 1;
    14: op1_08_inv28 = 1;
    18: op1_08_inv28 = 1;
    20: op1_08_inv28 = 1;
    21: op1_08_inv28 = 1;
    23: op1_08_inv28 = 1;
    26: op1_08_inv28 = 1;
    41: op1_08_inv28 = 1;
    45: op1_08_inv28 = 1;
    46: op1_08_inv28 = 1;
    47: op1_08_inv28 = 1;
    49: op1_08_inv28 = 1;
    52: op1_08_inv28 = 1;
    55: op1_08_inv28 = 1;
    56: op1_08_inv28 = 1;
    60: op1_08_inv28 = 1;
    62: op1_08_inv28 = 1;
    64: op1_08_inv28 = 1;
    65: op1_08_inv28 = 1;
    68: op1_08_inv28 = 1;
    70: op1_08_inv28 = 1;
    71: op1_08_inv28 = 1;
    72: op1_08_inv28 = 1;
    73: op1_08_inv28 = 1;
    75: op1_08_inv28 = 1;
    79: op1_08_inv28 = 1;
    82: op1_08_inv28 = 1;
    83: op1_08_inv28 = 1;
    84: op1_08_inv28 = 1;
    85: op1_08_inv28 = 1;
    88: op1_08_inv28 = 1;
    90: op1_08_inv28 = 1;
    91: op1_08_inv28 = 1;
    95: op1_08_inv28 = 1;
    97: op1_08_inv28 = 1;
    default: op1_08_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in29 = reg_0030;
    6: op1_08_in29 = imem05_in[107:104];
    8: op1_08_in29 = reg_0595;
    9: op1_08_in29 = reg_0608;
    10: op1_08_in29 = reg_0281;
    11: op1_08_in29 = reg_0719;
    12: op1_08_in29 = reg_0306;
    13: op1_08_in29 = reg_0216;
    14: op1_08_in29 = reg_0089;
    15: op1_08_in29 = reg_0558;
    17: op1_08_in29 = reg_1041;
    18: op1_08_in29 = imem07_in[79:76];
    19: op1_08_in29 = reg_0248;
    20: op1_08_in29 = reg_0159;
    21: op1_08_in29 = reg_1036;
    22: op1_08_in29 = reg_0390;
    23: op1_08_in29 = reg_0405;
    24: op1_08_in29 = reg_0628;
    25: op1_08_in29 = reg_0169;
    26: op1_08_in29 = reg_0398;
    28: op1_08_in29 = reg_0108;
    29: op1_08_in29 = reg_0706;
    31: op1_08_in29 = imem02_in[91:88];
    32: op1_08_in29 = reg_0763;
    33: op1_08_in29 = reg_0835;
    35: op1_08_in29 = imem04_in[83:80];
    36: op1_08_in29 = imem04_in[63:60];
    37: op1_08_in29 = imem05_in[91:88];
    38: op1_08_in29 = reg_0822;
    39: op1_08_in29 = reg_0395;
    47: op1_08_in29 = reg_0395;
    41: op1_08_in29 = reg_0157;
    42: op1_08_in29 = reg_0985;
    43: op1_08_in29 = reg_0285;
    44: op1_08_in29 = reg_0002;
    45: op1_08_in29 = reg_1017;
    46: op1_08_in29 = reg_0923;
    48: op1_08_in29 = reg_0122;
    49: op1_08_in29 = imem03_in[111:108];
    50: op1_08_in29 = reg_1039;
    52: op1_08_in29 = reg_0709;
    55: op1_08_in29 = imem02_in[123:120];
    56: op1_08_in29 = imem02_in[71:68];
    57: op1_08_in29 = reg_0291;
    58: op1_08_in29 = imem04_in[11:8];
    59: op1_08_in29 = reg_0978;
    60: op1_08_in29 = reg_0950;
    61: op1_08_in29 = reg_0968;
    62: op1_08_in29 = imem07_in[19:16];
    63: op1_08_in29 = reg_0592;
    64: op1_08_in29 = reg_0830;
    65: op1_08_in29 = imem03_in[43:40];
    66: op1_08_in29 = reg_0240;
    67: op1_08_in29 = reg_0836;
    68: op1_08_in29 = imem06_in[107:104];
    70: op1_08_in29 = reg_0981;
    71: op1_08_in29 = imem05_in[51:48];
    72: op1_08_in29 = reg_0514;
    73: op1_08_in29 = reg_0977;
    74: op1_08_in29 = reg_0396;
    82: op1_08_in29 = reg_0396;
    75: op1_08_in29 = reg_0707;
    76: op1_08_in29 = reg_0160;
    77: op1_08_in29 = reg_0172;
    79: op1_08_in29 = reg_0831;
    80: op1_08_in29 = imem04_in[35:32];
    81: op1_08_in29 = reg_0136;
    83: op1_08_in29 = reg_0615;
    84: op1_08_in29 = reg_0617;
    85: op1_08_in29 = reg_0823;
    86: op1_08_in29 = reg_0826;
    88: op1_08_in29 = imem02_in[51:48];
    90: op1_08_in29 = reg_0352;
    91: op1_08_in29 = reg_0359;
    92: op1_08_in29 = reg_0242;
    93: op1_08_in29 = reg_0611;
    94: op1_08_in29 = reg_0010;
    95: op1_08_in29 = reg_0144;
    97: op1_08_in29 = reg_0655;
    default: op1_08_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv29 = 1;
    6: op1_08_inv29 = 1;
    10: op1_08_inv29 = 1;
    12: op1_08_inv29 = 1;
    13: op1_08_inv29 = 1;
    15: op1_08_inv29 = 1;
    17: op1_08_inv29 = 1;
    18: op1_08_inv29 = 1;
    20: op1_08_inv29 = 1;
    22: op1_08_inv29 = 1;
    25: op1_08_inv29 = 1;
    26: op1_08_inv29 = 1;
    28: op1_08_inv29 = 1;
    29: op1_08_inv29 = 1;
    33: op1_08_inv29 = 1;
    39: op1_08_inv29 = 1;
    41: op1_08_inv29 = 1;
    42: op1_08_inv29 = 1;
    44: op1_08_inv29 = 1;
    45: op1_08_inv29 = 1;
    57: op1_08_inv29 = 1;
    61: op1_08_inv29 = 1;
    62: op1_08_inv29 = 1;
    66: op1_08_inv29 = 1;
    67: op1_08_inv29 = 1;
    68: op1_08_inv29 = 1;
    71: op1_08_inv29 = 1;
    72: op1_08_inv29 = 1;
    73: op1_08_inv29 = 1;
    80: op1_08_inv29 = 1;
    81: op1_08_inv29 = 1;
    82: op1_08_inv29 = 1;
    83: op1_08_inv29 = 1;
    85: op1_08_inv29 = 1;
    86: op1_08_inv29 = 1;
    91: op1_08_inv29 = 1;
    94: op1_08_inv29 = 1;
    95: op1_08_inv29 = 1;
    97: op1_08_inv29 = 1;
    default: op1_08_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_08_in30 = reg_0011;
    6: op1_08_in30 = imem05_in[119:116];
    8: op1_08_in30 = reg_0588;
    9: op1_08_in30 = reg_0632;
    10: op1_08_in30 = reg_0279;
    11: op1_08_in30 = reg_0731;
    12: op1_08_in30 = reg_0291;
    13: op1_08_in30 = reg_1036;
    14: op1_08_in30 = reg_0095;
    15: op1_08_in30 = reg_0282;
    17: op1_08_in30 = reg_0871;
    18: op1_08_in30 = imem07_in[99:96];
    19: op1_08_in30 = reg_0905;
    20: op1_08_in30 = reg_0182;
    21: op1_08_in30 = reg_1041;
    22: op1_08_in30 = reg_0380;
    23: op1_08_in30 = reg_0026;
    24: op1_08_in30 = reg_0620;
    25: op1_08_in30 = reg_0183;
    26: op1_08_in30 = reg_0376;
    28: op1_08_in30 = reg_0114;
    29: op1_08_in30 = reg_0430;
    31: op1_08_in30 = imem02_in[111:108];
    32: op1_08_in30 = reg_0062;
    33: op1_08_in30 = reg_0813;
    35: op1_08_in30 = imem04_in[95:92];
    36: op1_08_in30 = imem04_in[83:80];
    37: op1_08_in30 = reg_0970;
    38: op1_08_in30 = reg_0992;
    39: op1_08_in30 = reg_0042;
    42: op1_08_in30 = reg_0987;
    43: op1_08_in30 = imem05_in[27:24];
    44: op1_08_in30 = reg_0421;
    45: op1_08_in30 = reg_0111;
    46: op1_08_in30 = reg_0765;
    47: op1_08_in30 = reg_0386;
    48: op1_08_in30 = reg_0119;
    49: op1_08_in30 = imem03_in[119:116];
    50: op1_08_in30 = reg_0869;
    52: op1_08_in30 = reg_0715;
    55: op1_08_in30 = reg_0621;
    56: op1_08_in30 = imem02_in[75:72];
    57: op1_08_in30 = reg_0884;
    58: op1_08_in30 = imem04_in[19:16];
    59: op1_08_in30 = reg_0873;
    60: op1_08_in30 = reg_0221;
    61: op1_08_in30 = reg_0755;
    62: op1_08_in30 = imem07_in[23:20];
    63: op1_08_in30 = reg_0238;
    64: op1_08_in30 = reg_0500;
    65: op1_08_in30 = imem03_in[51:48];
    66: op1_08_in30 = reg_0833;
    67: op1_08_in30 = reg_0513;
    68: op1_08_in30 = imem06_in[119:116];
    70: op1_08_in30 = imem04_in[79:76];
    71: op1_08_in30 = imem05_in[87:84];
    72: op1_08_in30 = reg_0830;
    73: op1_08_in30 = reg_0990;
    74: op1_08_in30 = reg_0662;
    75: op1_08_in30 = reg_0019;
    76: op1_08_in30 = reg_0163;
    79: op1_08_in30 = reg_1043;
    80: op1_08_in30 = imem04_in[67:64];
    81: op1_08_in30 = reg_0139;
    82: op1_08_in30 = reg_0661;
    83: op1_08_in30 = reg_1053;
    84: op1_08_in30 = reg_0439;
    85: op1_08_in30 = reg_0038;
    86: op1_08_in30 = reg_0652;
    88: op1_08_in30 = imem02_in[79:76];
    90: op1_08_in30 = reg_0677;
    91: op1_08_in30 = reg_0423;
    92: op1_08_in30 = reg_0318;
    93: op1_08_in30 = imem07_in[27:24];
    94: op1_08_in30 = reg_0244;
    95: op1_08_in30 = imem06_in[27:24];
    97: op1_08_in30 = reg_0138;
    default: op1_08_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv30 = 1;
    11: op1_08_inv30 = 1;
    12: op1_08_inv30 = 1;
    13: op1_08_inv30 = 1;
    14: op1_08_inv30 = 1;
    15: op1_08_inv30 = 1;
    18: op1_08_inv30 = 1;
    19: op1_08_inv30 = 1;
    20: op1_08_inv30 = 1;
    21: op1_08_inv30 = 1;
    22: op1_08_inv30 = 1;
    24: op1_08_inv30 = 1;
    26: op1_08_inv30 = 1;
    28: op1_08_inv30 = 1;
    29: op1_08_inv30 = 1;
    33: op1_08_inv30 = 1;
    35: op1_08_inv30 = 1;
    37: op1_08_inv30 = 1;
    39: op1_08_inv30 = 1;
    47: op1_08_inv30 = 1;
    48: op1_08_inv30 = 1;
    50: op1_08_inv30 = 1;
    52: op1_08_inv30 = 1;
    55: op1_08_inv30 = 1;
    56: op1_08_inv30 = 1;
    58: op1_08_inv30 = 1;
    60: op1_08_inv30 = 1;
    64: op1_08_inv30 = 1;
    66: op1_08_inv30 = 1;
    70: op1_08_inv30 = 1;
    71: op1_08_inv30 = 1;
    72: op1_08_inv30 = 1;
    73: op1_08_inv30 = 1;
    74: op1_08_inv30 = 1;
    75: op1_08_inv30 = 1;
    79: op1_08_inv30 = 1;
    81: op1_08_inv30 = 1;
    83: op1_08_inv30 = 1;
    84: op1_08_inv30 = 1;
    88: op1_08_inv30 = 1;
    90: op1_08_inv30 = 1;
    94: op1_08_inv30 = 1;
    97: op1_08_inv30 = 1;
    default: op1_08_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_08_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_08_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in00 = imem07_in[43:40];
    6: op1_09_in00 = reg_0217;
    7: op1_09_in00 = imem00_in[79:76];
    8: op1_09_in00 = reg_0570;
    9: op1_09_in00 = reg_0623;
    10: op1_09_in00 = reg_0297;
    11: op1_09_in00 = imem00_in[35:32];
    54: op1_09_in00 = imem00_in[35:32];
    12: op1_09_in00 = reg_0292;
    13: op1_09_in00 = reg_1015;
    14: op1_09_in00 = reg_0085;
    15: op1_09_in00 = reg_0078;
    16: op1_09_in00 = imem00_in[31:28];
    41: op1_09_in00 = imem00_in[31:28];
    4: op1_09_in00 = imem07_in[79:76];
    17: op1_09_in00 = reg_1038;
    18: op1_09_in00 = imem00_in[15:12];
    87: op1_09_in00 = imem00_in[15:12];
    89: op1_09_in00 = imem00_in[15:12];
    19: op1_09_in00 = reg_1039;
    20: op1_09_in00 = imem00_in[19:16];
    21: op1_09_in00 = reg_1017;
    22: op1_09_in00 = reg_0799;
    23: op1_09_in00 = reg_0800;
    24: op1_09_in00 = reg_0631;
    3: op1_09_in00 = imem07_in[123:120];
    25: op1_09_in00 = imem00_in[39:36];
    26: op1_09_in00 = reg_0998;
    27: op1_09_in00 = imem00_in[59:56];
    28: op1_09_in00 = reg_0106;
    2: op1_09_in00 = imem07_in[51:48];
    29: op1_09_in00 = imem00_in[7:4];
    69: op1_09_in00 = imem00_in[7:4];
    96: op1_09_in00 = imem00_in[7:4];
    30: op1_09_in00 = imem00_in[75:72];
    31: op1_09_in00 = reg_0642;
    32: op1_09_in00 = reg_0755;
    33: op1_09_in00 = reg_0832;
    34: op1_09_in00 = imem00_in[11:8];
    53: op1_09_in00 = imem00_in[11:8];
    35: op1_09_in00 = imem04_in[119:116];
    36: op1_09_in00 = imem04_in[87:84];
    37: op1_09_in00 = reg_0956;
    38: op1_09_in00 = reg_0979;
    39: op1_09_in00 = reg_0388;
    40: op1_09_in00 = imem00_in[47:44];
    78: op1_09_in00 = imem00_in[47:44];
    42: op1_09_in00 = reg_0990;
    43: op1_09_in00 = imem05_in[39:36];
    44: op1_09_in00 = reg_0321;
    45: op1_09_in00 = reg_0104;
    46: op1_09_in00 = reg_0038;
    47: op1_09_in00 = reg_0349;
    48: op1_09_in00 = reg_0102;
    49: op1_09_in00 = imem03_in[127:124];
    50: op1_09_in00 = reg_0520;
    51: op1_09_in00 = imem00_in[3:0];
    77: op1_09_in00 = imem00_in[3:0];
    52: op1_09_in00 = reg_0599;
    55: op1_09_in00 = reg_0300;
    56: op1_09_in00 = reg_0326;
    57: op1_09_in00 = imem03_in[11:8];
    58: op1_09_in00 = imem04_in[35:32];
    59: op1_09_in00 = reg_0122;
    60: op1_09_in00 = reg_0035;
    61: op1_09_in00 = imem05_in[31:28];
    62: op1_09_in00 = imem07_in[27:24];
    63: op1_09_in00 = reg_0604;
    64: op1_09_in00 = reg_0216;
    65: op1_09_in00 = imem03_in[59:56];
    66: op1_09_in00 = reg_0051;
    67: op1_09_in00 = reg_0844;
    68: op1_09_in00 = imem06_in[127:124];
    70: op1_09_in00 = reg_1009;
    71: op1_09_in00 = imem05_in[115:112];
    72: op1_09_in00 = reg_0616;
    73: op1_09_in00 = imem04_in[15:12];
    92: op1_09_in00 = imem04_in[15:12];
    74: op1_09_in00 = reg_0238;
    75: op1_09_in00 = reg_0806;
    76: op1_09_in00 = reg_0164;
    79: op1_09_in00 = reg_0830;
    80: op1_09_in00 = reg_0301;
    81: op1_09_in00 = reg_0138;
    82: op1_09_in00 = reg_0576;
    83: op1_09_in00 = reg_1033;
    84: op1_09_in00 = reg_0382;
    85: op1_09_in00 = reg_0609;
    86: op1_09_in00 = reg_0128;
    88: op1_09_in00 = imem02_in[87:84];
    90: op1_09_in00 = reg_0004;
    91: op1_09_in00 = reg_0394;
    93: op1_09_in00 = imem07_in[31:28];
    94: op1_09_in00 = reg_0267;
    95: op1_09_in00 = imem06_in[91:88];
    97: op1_09_in00 = reg_0448;
    default: op1_09_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv00 = 1;
    7: op1_09_inv00 = 1;
    12: op1_09_inv00 = 1;
    14: op1_09_inv00 = 1;
    16: op1_09_inv00 = 1;
    19: op1_09_inv00 = 1;
    20: op1_09_inv00 = 1;
    25: op1_09_inv00 = 1;
    29: op1_09_inv00 = 1;
    31: op1_09_inv00 = 1;
    36: op1_09_inv00 = 1;
    38: op1_09_inv00 = 1;
    39: op1_09_inv00 = 1;
    41: op1_09_inv00 = 1;
    42: op1_09_inv00 = 1;
    43: op1_09_inv00 = 1;
    45: op1_09_inv00 = 1;
    50: op1_09_inv00 = 1;
    51: op1_09_inv00 = 1;
    52: op1_09_inv00 = 1;
    55: op1_09_inv00 = 1;
    56: op1_09_inv00 = 1;
    57: op1_09_inv00 = 1;
    59: op1_09_inv00 = 1;
    60: op1_09_inv00 = 1;
    62: op1_09_inv00 = 1;
    63: op1_09_inv00 = 1;
    64: op1_09_inv00 = 1;
    66: op1_09_inv00 = 1;
    74: op1_09_inv00 = 1;
    75: op1_09_inv00 = 1;
    76: op1_09_inv00 = 1;
    77: op1_09_inv00 = 1;
    79: op1_09_inv00 = 1;
    80: op1_09_inv00 = 1;
    81: op1_09_inv00 = 1;
    83: op1_09_inv00 = 1;
    86: op1_09_inv00 = 1;
    92: op1_09_inv00 = 1;
    94: op1_09_inv00 = 1;
    95: op1_09_inv00 = 1;
    96: op1_09_inv00 = 1;
    97: op1_09_inv00 = 1;
    default: op1_09_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in01 = imem07_in[115:112];
    6: op1_09_in01 = reg_0269;
    7: op1_09_in01 = imem00_in[87:84];
    8: op1_09_in01 = reg_0311;
    9: op1_09_in01 = reg_0348;
    10: op1_09_in01 = reg_0275;
    12: op1_09_in01 = reg_0275;
    11: op1_09_in01 = imem00_in[75:72];
    27: op1_09_in01 = imem00_in[75:72];
    13: op1_09_in01 = reg_1017;
    14: op1_09_in01 = reg_0096;
    15: op1_09_in01 = reg_0065;
    16: op1_09_in01 = imem00_in[39:36];
    18: op1_09_in01 = imem00_in[39:36];
    20: op1_09_in01 = imem00_in[39:36];
    54: op1_09_in01 = imem00_in[39:36];
    89: op1_09_in01 = imem00_in[39:36];
    4: op1_09_in01 = imem07_in[91:88];
    17: op1_09_in01 = reg_0122;
    19: op1_09_in01 = reg_0869;
    21: op1_09_in01 = reg_0114;
    22: op1_09_in01 = reg_1028;
    23: op1_09_in01 = reg_0808;
    24: op1_09_in01 = reg_0608;
    3: op1_09_in01 = reg_0174;
    25: op1_09_in01 = imem00_in[71:68];
    26: op1_09_in01 = reg_0986;
    28: op1_09_in01 = reg_0110;
    2: op1_09_in01 = imem07_in[99:96];
    29: op1_09_in01 = imem00_in[27:24];
    77: op1_09_in01 = imem00_in[27:24];
    30: op1_09_in01 = imem00_in[99:96];
    31: op1_09_in01 = reg_0661;
    32: op1_09_in01 = reg_0071;
    33: op1_09_in01 = reg_0135;
    34: op1_09_in01 = reg_0693;
    35: op1_09_in01 = reg_0277;
    36: op1_09_in01 = imem04_in[107:104];
    37: op1_09_in01 = reg_0957;
    38: op1_09_in01 = reg_0978;
    39: op1_09_in01 = reg_0628;
    40: op1_09_in01 = imem00_in[51:48];
    41: op1_09_in01 = imem00_in[47:44];
    42: op1_09_in01 = reg_0305;
    43: op1_09_in01 = imem05_in[51:48];
    44: op1_09_in01 = reg_0353;
    45: op1_09_in01 = reg_0119;
    46: op1_09_in01 = reg_0985;
    47: op1_09_in01 = reg_0222;
    48: op1_09_in01 = reg_0107;
    49: op1_09_in01 = reg_0004;
    50: op1_09_in01 = reg_1043;
    51: op1_09_in01 = imem00_in[11:8];
    52: op1_09_in01 = reg_0024;
    53: op1_09_in01 = imem00_in[31:28];
    55: op1_09_in01 = reg_0648;
    86: op1_09_in01 = reg_0648;
    56: op1_09_in01 = reg_0636;
    57: op1_09_in01 = imem03_in[23:20];
    58: op1_09_in01 = imem04_in[43:40];
    59: op1_09_in01 = reg_0367;
    60: op1_09_in01 = reg_0952;
    61: op1_09_in01 = imem05_in[115:112];
    62: op1_09_in01 = imem07_in[39:36];
    63: op1_09_in01 = reg_0829;
    64: op1_09_in01 = reg_0354;
    65: op1_09_in01 = imem03_in[83:80];
    66: op1_09_in01 = reg_0981;
    67: op1_09_in01 = reg_0822;
    68: op1_09_in01 = reg_0338;
    69: op1_09_in01 = imem00_in[35:32];
    70: op1_09_in01 = reg_0282;
    71: op1_09_in01 = reg_0030;
    72: op1_09_in01 = reg_0610;
    73: op1_09_in01 = imem04_in[23:20];
    74: op1_09_in01 = reg_0756;
    75: op1_09_in01 = reg_0706;
    76: op1_09_in01 = reg_0185;
    78: op1_09_in01 = imem00_in[67:64];
    79: op1_09_in01 = reg_0902;
    80: op1_09_in01 = reg_1003;
    81: op1_09_in01 = reg_0137;
    82: op1_09_in01 = reg_0397;
    83: op1_09_in01 = reg_0112;
    84: op1_09_in01 = reg_0591;
    85: op1_09_in01 = reg_0051;
    87: op1_09_in01 = imem00_in[43:40];
    88: op1_09_in01 = imem02_in[123:120];
    90: op1_09_in01 = reg_0570;
    91: op1_09_in01 = reg_0087;
    92: op1_09_in01 = imem04_in[35:32];
    93: op1_09_in01 = imem07_in[51:48];
    94: op1_09_in01 = reg_0393;
    95: op1_09_in01 = imem06_in[107:104];
    96: op1_09_in01 = imem00_in[19:16];
    97: op1_09_in01 = reg_0689;
    default: op1_09_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv01 = 1;
    6: op1_09_inv01 = 1;
    8: op1_09_inv01 = 1;
    15: op1_09_inv01 = 1;
    4: op1_09_inv01 = 1;
    17: op1_09_inv01 = 1;
    18: op1_09_inv01 = 1;
    20: op1_09_inv01 = 1;
    3: op1_09_inv01 = 1;
    25: op1_09_inv01 = 1;
    27: op1_09_inv01 = 1;
    28: op1_09_inv01 = 1;
    30: op1_09_inv01 = 1;
    33: op1_09_inv01 = 1;
    35: op1_09_inv01 = 1;
    37: op1_09_inv01 = 1;
    38: op1_09_inv01 = 1;
    40: op1_09_inv01 = 1;
    41: op1_09_inv01 = 1;
    42: op1_09_inv01 = 1;
    44: op1_09_inv01 = 1;
    45: op1_09_inv01 = 1;
    48: op1_09_inv01 = 1;
    49: op1_09_inv01 = 1;
    50: op1_09_inv01 = 1;
    52: op1_09_inv01 = 1;
    53: op1_09_inv01 = 1;
    54: op1_09_inv01 = 1;
    56: op1_09_inv01 = 1;
    57: op1_09_inv01 = 1;
    58: op1_09_inv01 = 1;
    59: op1_09_inv01 = 1;
    61: op1_09_inv01 = 1;
    62: op1_09_inv01 = 1;
    63: op1_09_inv01 = 1;
    65: op1_09_inv01 = 1;
    69: op1_09_inv01 = 1;
    70: op1_09_inv01 = 1;
    71: op1_09_inv01 = 1;
    72: op1_09_inv01 = 1;
    73: op1_09_inv01 = 1;
    75: op1_09_inv01 = 1;
    76: op1_09_inv01 = 1;
    81: op1_09_inv01 = 1;
    85: op1_09_inv01 = 1;
    87: op1_09_inv01 = 1;
    88: op1_09_inv01 = 1;
    91: op1_09_inv01 = 1;
    92: op1_09_inv01 = 1;
    94: op1_09_inv01 = 1;
    95: op1_09_inv01 = 1;
    97: op1_09_inv01 = 1;
    default: op1_09_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in02 = imem07_in[127:124];
    6: op1_09_in02 = reg_0263;
    7: op1_09_in02 = imem00_in[91:88];
    8: op1_09_in02 = reg_0376;
    9: op1_09_in02 = reg_0313;
    10: op1_09_in02 = reg_0065;
    11: op1_09_in02 = imem00_in[83:80];
    12: op1_09_in02 = reg_0054;
    13: op1_09_in02 = reg_0111;
    14: op1_09_in02 = reg_0097;
    15: op1_09_in02 = reg_0048;
    16: op1_09_in02 = imem00_in[47:44];
    18: op1_09_in02 = imem00_in[47:44];
    87: op1_09_in02 = imem00_in[47:44];
    4: op1_09_in02 = imem07_in[99:96];
    17: op1_09_in02 = reg_0116;
    79: op1_09_in02 = reg_0116;
    19: op1_09_in02 = reg_1033;
    20: op1_09_in02 = imem00_in[55:52];
    41: op1_09_in02 = imem00_in[55:52];
    54: op1_09_in02 = imem00_in[55:52];
    21: op1_09_in02 = reg_0109;
    22: op1_09_in02 = reg_0801;
    23: op1_09_in02 = reg_0486;
    24: op1_09_in02 = reg_0632;
    3: op1_09_in02 = reg_0161;
    25: op1_09_in02 = imem00_in[99:96];
    26: op1_09_in02 = reg_0980;
    27: op1_09_in02 = imem00_in[115:112];
    28: op1_09_in02 = imem02_in[19:16];
    29: op1_09_in02 = imem00_in[35:32];
    96: op1_09_in02 = imem00_in[35:32];
    30: op1_09_in02 = reg_0682;
    31: op1_09_in02 = reg_0656;
    32: op1_09_in02 = reg_0069;
    33: op1_09_in02 = reg_0139;
    34: op1_09_in02 = reg_0694;
    35: op1_09_in02 = reg_0055;
    36: op1_09_in02 = reg_0265;
    37: op1_09_in02 = reg_0942;
    38: op1_09_in02 = reg_0990;
    39: op1_09_in02 = reg_0625;
    40: op1_09_in02 = imem00_in[71:68];
    42: op1_09_in02 = reg_0750;
    43: op1_09_in02 = imem05_in[71:68];
    44: op1_09_in02 = reg_0599;
    45: op1_09_in02 = reg_0100;
    46: op1_09_in02 = reg_0982;
    47: op1_09_in02 = reg_0628;
    48: op1_09_in02 = imem02_in[43:40];
    49: op1_09_in02 = reg_0576;
    50: op1_09_in02 = reg_0830;
    51: op1_09_in02 = imem00_in[19:16];
    52: op1_09_in02 = reg_0431;
    53: op1_09_in02 = imem00_in[59:56];
    55: op1_09_in02 = reg_0854;
    56: op1_09_in02 = reg_0739;
    57: op1_09_in02 = imem03_in[51:48];
    58: op1_09_in02 = imem04_in[59:56];
    59: op1_09_in02 = reg_0773;
    60: op1_09_in02 = reg_0953;
    61: op1_09_in02 = imem05_in[127:124];
    62: op1_09_in02 = imem07_in[107:104];
    63: op1_09_in02 = reg_1041;
    64: op1_09_in02 = reg_0832;
    65: op1_09_in02 = reg_0006;
    66: op1_09_in02 = reg_0983;
    67: op1_09_in02 = reg_0996;
    68: op1_09_in02 = reg_0614;
    69: op1_09_in02 = imem00_in[51:48];
    70: op1_09_in02 = reg_0912;
    71: op1_09_in02 = reg_0326;
    72: op1_09_in02 = reg_1017;
    73: op1_09_in02 = imem04_in[27:24];
    74: op1_09_in02 = reg_0596;
    75: op1_09_in02 = reg_0795;
    77: op1_09_in02 = imem00_in[43:40];
    78: op1_09_in02 = imem00_in[119:116];
    89: op1_09_in02 = imem00_in[119:116];
    80: op1_09_in02 = reg_0277;
    81: op1_09_in02 = reg_0648;
    82: op1_09_in02 = reg_0579;
    83: op1_09_in02 = reg_0860;
    84: op1_09_in02 = reg_0699;
    85: op1_09_in02 = reg_0820;
    86: op1_09_in02 = reg_0057;
    88: op1_09_in02 = reg_0255;
    90: op1_09_in02 = reg_0785;
    91: op1_09_in02 = reg_0608;
    92: op1_09_in02 = imem04_in[55:52];
    93: op1_09_in02 = imem07_in[63:60];
    94: op1_09_in02 = reg_0440;
    95: op1_09_in02 = reg_0660;
    97: op1_09_in02 = reg_0269;
    default: op1_09_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv02 = 1;
    11: op1_09_inv02 = 1;
    12: op1_09_inv02 = 1;
    13: op1_09_inv02 = 1;
    4: op1_09_inv02 = 1;
    17: op1_09_inv02 = 1;
    24: op1_09_inv02 = 1;
    3: op1_09_inv02 = 1;
    26: op1_09_inv02 = 1;
    28: op1_09_inv02 = 1;
    30: op1_09_inv02 = 1;
    32: op1_09_inv02 = 1;
    35: op1_09_inv02 = 1;
    36: op1_09_inv02 = 1;
    40: op1_09_inv02 = 1;
    41: op1_09_inv02 = 1;
    42: op1_09_inv02 = 1;
    43: op1_09_inv02 = 1;
    45: op1_09_inv02 = 1;
    47: op1_09_inv02 = 1;
    51: op1_09_inv02 = 1;
    53: op1_09_inv02 = 1;
    55: op1_09_inv02 = 1;
    56: op1_09_inv02 = 1;
    57: op1_09_inv02 = 1;
    59: op1_09_inv02 = 1;
    60: op1_09_inv02 = 1;
    61: op1_09_inv02 = 1;
    66: op1_09_inv02 = 1;
    68: op1_09_inv02 = 1;
    71: op1_09_inv02 = 1;
    73: op1_09_inv02 = 1;
    74: op1_09_inv02 = 1;
    75: op1_09_inv02 = 1;
    80: op1_09_inv02 = 1;
    81: op1_09_inv02 = 1;
    82: op1_09_inv02 = 1;
    83: op1_09_inv02 = 1;
    87: op1_09_inv02 = 1;
    88: op1_09_inv02 = 1;
    94: op1_09_inv02 = 1;
    95: op1_09_inv02 = 1;
    default: op1_09_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in03 = reg_0719;
    6: op1_09_in03 = reg_0149;
    7: op1_09_in03 = imem00_in[103:100];
    8: op1_09_in03 = reg_0996;
    9: op1_09_in03 = imem06_in[27:24];
    10: op1_09_in03 = reg_0058;
    11: op1_09_in03 = imem00_in[111:108];
    69: op1_09_in03 = imem00_in[111:108];
    12: op1_09_in03 = reg_0065;
    13: op1_09_in03 = reg_0116;
    63: op1_09_in03 = reg_0116;
    14: op1_09_in03 = reg_0087;
    15: op1_09_in03 = reg_0050;
    16: op1_09_in03 = imem00_in[79:76];
    18: op1_09_in03 = imem00_in[79:76];
    4: op1_09_in03 = imem07_in[115:112];
    17: op1_09_in03 = reg_0120;
    19: op1_09_in03 = reg_0227;
    20: op1_09_in03 = imem00_in[91:88];
    21: op1_09_in03 = reg_0535;
    22: op1_09_in03 = imem07_in[19:16];
    23: op1_09_in03 = reg_0801;
    24: op1_09_in03 = reg_0332;
    3: op1_09_in03 = reg_0162;
    25: op1_09_in03 = imem00_in[123:120];
    26: op1_09_in03 = reg_0975;
    27: op1_09_in03 = imem00_in[127:124];
    40: op1_09_in03 = imem00_in[127:124];
    28: op1_09_in03 = imem02_in[47:44];
    48: op1_09_in03 = imem02_in[47:44];
    29: op1_09_in03 = imem00_in[67:64];
    54: op1_09_in03 = imem00_in[67:64];
    30: op1_09_in03 = reg_0693;
    31: op1_09_in03 = reg_0641;
    32: op1_09_in03 = reg_0064;
    33: op1_09_in03 = imem06_in[3:0];
    34: op1_09_in03 = reg_0689;
    35: op1_09_in03 = reg_0048;
    36: op1_09_in03 = reg_1057;
    37: op1_09_in03 = reg_0961;
    38: op1_09_in03 = reg_0976;
    39: op1_09_in03 = reg_0617;
    68: op1_09_in03 = reg_0617;
    41: op1_09_in03 = imem00_in[83:80];
    53: op1_09_in03 = imem00_in[83:80];
    42: op1_09_in03 = reg_0588;
    43: op1_09_in03 = imem05_in[79:76];
    44: op1_09_in03 = reg_0589;
    45: op1_09_in03 = reg_0113;
    46: op1_09_in03 = reg_1001;
    47: op1_09_in03 = reg_0894;
    49: op1_09_in03 = reg_0373;
    50: op1_09_in03 = reg_0500;
    51: op1_09_in03 = imem00_in[35:32];
    52: op1_09_in03 = reg_0174;
    55: op1_09_in03 = reg_0652;
    56: op1_09_in03 = reg_0441;
    57: op1_09_in03 = imem03_in[71:68];
    58: op1_09_in03 = imem04_in[79:76];
    59: op1_09_in03 = reg_0539;
    80: op1_09_in03 = reg_0539;
    60: op1_09_in03 = reg_0019;
    61: op1_09_in03 = reg_0019;
    62: op1_09_in03 = reg_0726;
    64: op1_09_in03 = reg_0273;
    65: op1_09_in03 = reg_0760;
    66: op1_09_in03 = reg_0994;
    67: op1_09_in03 = reg_0993;
    70: op1_09_in03 = reg_0778;
    71: op1_09_in03 = reg_0667;
    72: op1_09_in03 = reg_0615;
    73: op1_09_in03 = imem04_in[59:56];
    74: op1_09_in03 = reg_0820;
    75: op1_09_in03 = reg_0950;
    77: op1_09_in03 = imem00_in[87:84];
    78: op1_09_in03 = reg_0768;
    79: op1_09_in03 = reg_1033;
    81: op1_09_in03 = reg_0966;
    82: op1_09_in03 = reg_1008;
    83: op1_09_in03 = reg_0101;
    84: op1_09_in03 = reg_0289;
    85: op1_09_in03 = reg_0233;
    86: op1_09_in03 = reg_0953;
    87: op1_09_in03 = imem00_in[99:96];
    88: op1_09_in03 = reg_0091;
    89: op1_09_in03 = reg_0519;
    90: op1_09_in03 = reg_0317;
    91: op1_09_in03 = reg_0650;
    92: op1_09_in03 = imem04_in[63:60];
    93: op1_09_in03 = imem07_in[71:68];
    94: op1_09_in03 = reg_0895;
    95: op1_09_in03 = reg_0267;
    96: op1_09_in03 = imem00_in[43:40];
    97: op1_09_in03 = reg_0057;
    default: op1_09_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv03 = 1;
    7: op1_09_inv03 = 1;
    9: op1_09_inv03 = 1;
    11: op1_09_inv03 = 1;
    13: op1_09_inv03 = 1;
    14: op1_09_inv03 = 1;
    15: op1_09_inv03 = 1;
    16: op1_09_inv03 = 1;
    22: op1_09_inv03 = 1;
    3: op1_09_inv03 = 1;
    25: op1_09_inv03 = 1;
    29: op1_09_inv03 = 1;
    32: op1_09_inv03 = 1;
    34: op1_09_inv03 = 1;
    35: op1_09_inv03 = 1;
    38: op1_09_inv03 = 1;
    39: op1_09_inv03 = 1;
    40: op1_09_inv03 = 1;
    42: op1_09_inv03 = 1;
    43: op1_09_inv03 = 1;
    44: op1_09_inv03 = 1;
    46: op1_09_inv03 = 1;
    47: op1_09_inv03 = 1;
    49: op1_09_inv03 = 1;
    50: op1_09_inv03 = 1;
    51: op1_09_inv03 = 1;
    54: op1_09_inv03 = 1;
    55: op1_09_inv03 = 1;
    58: op1_09_inv03 = 1;
    59: op1_09_inv03 = 1;
    60: op1_09_inv03 = 1;
    62: op1_09_inv03 = 1;
    63: op1_09_inv03 = 1;
    64: op1_09_inv03 = 1;
    71: op1_09_inv03 = 1;
    74: op1_09_inv03 = 1;
    78: op1_09_inv03 = 1;
    79: op1_09_inv03 = 1;
    83: op1_09_inv03 = 1;
    85: op1_09_inv03 = 1;
    87: op1_09_inv03 = 1;
    88: op1_09_inv03 = 1;
    90: op1_09_inv03 = 1;
    92: op1_09_inv03 = 1;
    93: op1_09_inv03 = 1;
    94: op1_09_inv03 = 1;
    97: op1_09_inv03 = 1;
    default: op1_09_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in04 = reg_0720;
    6: op1_09_in04 = reg_0150;
    7: op1_09_in04 = reg_0682;
    87: op1_09_in04 = reg_0682;
    8: op1_09_in04 = reg_0978;
    9: op1_09_in04 = imem07_in[39:36];
    10: op1_09_in04 = reg_0068;
    11: op1_09_in04 = reg_0685;
    12: op1_09_in04 = reg_0048;
    13: op1_09_in04 = reg_0113;
    14: op1_09_in04 = reg_0094;
    15: op1_09_in04 = imem05_in[39:36];
    16: op1_09_in04 = imem00_in[87:84];
    4: op1_09_in04 = reg_0422;
    17: op1_09_in04 = reg_0114;
    18: op1_09_in04 = imem00_in[95:92];
    41: op1_09_in04 = imem00_in[95:92];
    19: op1_09_in04 = reg_0228;
    20: op1_09_in04 = imem00_in[99:96];
    53: op1_09_in04 = imem00_in[99:96];
    21: op1_09_in04 = reg_0793;
    22: op1_09_in04 = imem07_in[59:56];
    23: op1_09_in04 = reg_0802;
    24: op1_09_in04 = reg_0381;
    3: op1_09_in04 = reg_0184;
    25: op1_09_in04 = reg_0693;
    26: op1_09_in04 = reg_0988;
    46: op1_09_in04 = reg_0988;
    27: op1_09_in04 = reg_0672;
    28: op1_09_in04 = imem02_in[51:48];
    29: op1_09_in04 = imem00_in[75:72];
    30: op1_09_in04 = reg_0697;
    40: op1_09_in04 = reg_0697;
    31: op1_09_in04 = reg_0636;
    32: op1_09_in04 = reg_0732;
    33: op1_09_in04 = imem06_in[87:84];
    34: op1_09_in04 = reg_0677;
    35: op1_09_in04 = reg_0292;
    59: op1_09_in04 = reg_0292;
    36: op1_09_in04 = reg_1016;
    37: op1_09_in04 = reg_0806;
    38: op1_09_in04 = imem04_in[11:8];
    39: op1_09_in04 = reg_0626;
    42: op1_09_in04 = reg_0265;
    43: op1_09_in04 = imem05_in[87:84];
    44: op1_09_in04 = reg_0502;
    45: op1_09_in04 = reg_0645;
    47: op1_09_in04 = reg_0241;
    48: op1_09_in04 = imem02_in[55:52];
    49: op1_09_in04 = reg_0836;
    50: op1_09_in04 = reg_1040;
    51: op1_09_in04 = imem00_in[43:40];
    52: op1_09_in04 = reg_0175;
    54: op1_09_in04 = imem00_in[83:80];
    55: op1_09_in04 = reg_0424;
    56: op1_09_in04 = reg_0424;
    57: op1_09_in04 = imem03_in[95:92];
    58: op1_09_in04 = imem04_in[91:88];
    60: op1_09_in04 = reg_0022;
    61: op1_09_in04 = reg_0493;
    62: op1_09_in04 = reg_0725;
    63: op1_09_in04 = reg_0283;
    64: op1_09_in04 = reg_0745;
    65: op1_09_in04 = reg_0580;
    66: op1_09_in04 = imem04_in[7:4];
    67: op1_09_in04 = reg_0980;
    68: op1_09_in04 = reg_0533;
    69: op1_09_in04 = reg_0900;
    70: op1_09_in04 = reg_0537;
    71: op1_09_in04 = reg_0255;
    72: op1_09_in04 = reg_0832;
    73: op1_09_in04 = imem04_in[95:92];
    74: op1_09_in04 = reg_0581;
    75: op1_09_in04 = reg_0741;
    77: op1_09_in04 = imem00_in[127:124];
    78: op1_09_in04 = reg_0686;
    79: op1_09_in04 = reg_0273;
    80: op1_09_in04 = reg_0752;
    81: op1_09_in04 = reg_0948;
    82: op1_09_in04 = reg_1049;
    83: op1_09_in04 = reg_0115;
    84: op1_09_in04 = reg_1010;
    85: op1_09_in04 = reg_0266;
    86: op1_09_in04 = reg_0314;
    88: op1_09_in04 = reg_0279;
    89: op1_09_in04 = reg_0768;
    90: op1_09_in04 = reg_0743;
    91: op1_09_in04 = reg_0045;
    92: op1_09_in04 = reg_0511;
    93: op1_09_in04 = imem07_in[83:80];
    94: op1_09_in04 = reg_0792;
    95: op1_09_in04 = reg_0229;
    96: op1_09_in04 = imem00_in[47:44];
    97: op1_09_in04 = reg_0935;
    default: op1_09_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv04 = 1;
    12: op1_09_inv04 = 1;
    16: op1_09_inv04 = 1;
    17: op1_09_inv04 = 1;
    20: op1_09_inv04 = 1;
    24: op1_09_inv04 = 1;
    3: op1_09_inv04 = 1;
    25: op1_09_inv04 = 1;
    28: op1_09_inv04 = 1;
    31: op1_09_inv04 = 1;
    34: op1_09_inv04 = 1;
    35: op1_09_inv04 = 1;
    36: op1_09_inv04 = 1;
    39: op1_09_inv04 = 1;
    40: op1_09_inv04 = 1;
    42: op1_09_inv04 = 1;
    43: op1_09_inv04 = 1;
    47: op1_09_inv04 = 1;
    51: op1_09_inv04 = 1;
    52: op1_09_inv04 = 1;
    53: op1_09_inv04 = 1;
    54: op1_09_inv04 = 1;
    55: op1_09_inv04 = 1;
    56: op1_09_inv04 = 1;
    57: op1_09_inv04 = 1;
    60: op1_09_inv04 = 1;
    65: op1_09_inv04 = 1;
    68: op1_09_inv04 = 1;
    69: op1_09_inv04 = 1;
    70: op1_09_inv04 = 1;
    71: op1_09_inv04 = 1;
    72: op1_09_inv04 = 1;
    73: op1_09_inv04 = 1;
    74: op1_09_inv04 = 1;
    77: op1_09_inv04 = 1;
    78: op1_09_inv04 = 1;
    79: op1_09_inv04 = 1;
    81: op1_09_inv04 = 1;
    84: op1_09_inv04 = 1;
    85: op1_09_inv04 = 1;
    88: op1_09_inv04 = 1;
    91: op1_09_inv04 = 1;
    92: op1_09_inv04 = 1;
    94: op1_09_inv04 = 1;
    96: op1_09_inv04 = 1;
    default: op1_09_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in05 = reg_0721;
    6: op1_09_in05 = reg_0152;
    7: op1_09_in05 = reg_0684;
    89: op1_09_in05 = reg_0684;
    8: op1_09_in05 = reg_0989;
    9: op1_09_in05 = imem07_in[123:120];
    10: op1_09_in05 = reg_0048;
    11: op1_09_in05 = reg_0688;
    12: op1_09_in05 = reg_1021;
    13: op1_09_in05 = imem02_in[3:0];
    14: op1_09_in05 = imem03_in[7:4];
    15: op1_09_in05 = imem05_in[75:72];
    16: op1_09_in05 = imem00_in[107:104];
    4: op1_09_in05 = reg_0423;
    17: op1_09_in05 = reg_0127;
    18: op1_09_in05 = reg_0693;
    20: op1_09_in05 = reg_0693;
    19: op1_09_in05 = reg_1017;
    21: op1_09_in05 = reg_0666;
    22: op1_09_in05 = imem07_in[67:64];
    23: op1_09_in05 = reg_0753;
    24: op1_09_in05 = reg_0390;
    25: op1_09_in05 = reg_0689;
    26: op1_09_in05 = reg_0990;
    27: op1_09_in05 = reg_0670;
    28: op1_09_in05 = imem02_in[55:52];
    29: op1_09_in05 = imem00_in[99:96];
    51: op1_09_in05 = imem00_in[99:96];
    54: op1_09_in05 = imem00_in[99:96];
    30: op1_09_in05 = reg_0683;
    40: op1_09_in05 = reg_0683;
    31: op1_09_in05 = reg_0096;
    32: op1_09_in05 = reg_0059;
    33: op1_09_in05 = imem06_in[95:92];
    34: op1_09_in05 = reg_0678;
    35: op1_09_in05 = reg_0074;
    36: op1_09_in05 = reg_0065;
    37: op1_09_in05 = reg_0149;
    38: op1_09_in05 = imem04_in[15:12];
    39: op1_09_in05 = reg_0926;
    41: op1_09_in05 = reg_0697;
    42: op1_09_in05 = imem04_in[7:4];
    43: op1_09_in05 = reg_0963;
    44: op1_09_in05 = reg_0024;
    45: op1_09_in05 = imem02_in[11:8];
    46: op1_09_in05 = reg_0352;
    47: op1_09_in05 = reg_0631;
    48: op1_09_in05 = reg_0650;
    49: op1_09_in05 = reg_1002;
    50: op1_09_in05 = reg_0616;
    52: op1_09_in05 = reg_0165;
    53: op1_09_in05 = reg_0695;
    55: op1_09_in05 = reg_0331;
    56: op1_09_in05 = reg_0425;
    57: op1_09_in05 = imem03_in[111:108];
    58: op1_09_in05 = imem04_in[127:124];
    59: op1_09_in05 = reg_0931;
    60: op1_09_in05 = reg_0032;
    61: op1_09_in05 = reg_0819;
    62: op1_09_in05 = reg_0729;
    94: op1_09_in05 = reg_0729;
    63: op1_09_in05 = reg_0860;
    64: op1_09_in05 = imem02_in[27:24];
    65: op1_09_in05 = reg_0585;
    66: op1_09_in05 = imem04_in[43:40];
    67: op1_09_in05 = reg_0999;
    74: op1_09_in05 = reg_0999;
    68: op1_09_in05 = reg_0011;
    69: op1_09_in05 = reg_0356;
    70: op1_09_in05 = reg_0802;
    71: op1_09_in05 = reg_0259;
    72: op1_09_in05 = reg_1055;
    73: op1_09_in05 = reg_1003;
    75: op1_09_in05 = imem06_in[63:60];
    77: op1_09_in05 = reg_0768;
    78: op1_09_in05 = reg_0451;
    79: op1_09_in05 = reg_0109;
    80: op1_09_in05 = reg_0288;
    81: op1_09_in05 = reg_1046;
    82: op1_09_in05 = reg_0376;
    83: op1_09_in05 = reg_0110;
    84: op1_09_in05 = reg_0403;
    85: op1_09_in05 = reg_0982;
    86: op1_09_in05 = reg_0957;
    87: op1_09_in05 = reg_0671;
    88: op1_09_in05 = reg_0359;
    90: op1_09_in05 = reg_0049;
    91: op1_09_in05 = reg_0776;
    92: op1_09_in05 = reg_1009;
    93: op1_09_in05 = imem07_in[95:92];
    95: op1_09_in05 = reg_0735;
    96: op1_09_in05 = imem00_in[63:60];
    97: op1_09_in05 = reg_0146;
    default: op1_09_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv05 = 1;
    7: op1_09_inv05 = 1;
    9: op1_09_inv05 = 1;
    10: op1_09_inv05 = 1;
    12: op1_09_inv05 = 1;
    13: op1_09_inv05 = 1;
    14: op1_09_inv05 = 1;
    16: op1_09_inv05 = 1;
    17: op1_09_inv05 = 1;
    18: op1_09_inv05 = 1;
    20: op1_09_inv05 = 1;
    21: op1_09_inv05 = 1;
    22: op1_09_inv05 = 1;
    23: op1_09_inv05 = 1;
    24: op1_09_inv05 = 1;
    25: op1_09_inv05 = 1;
    26: op1_09_inv05 = 1;
    27: op1_09_inv05 = 1;
    29: op1_09_inv05 = 1;
    31: op1_09_inv05 = 1;
    33: op1_09_inv05 = 1;
    35: op1_09_inv05 = 1;
    37: op1_09_inv05 = 1;
    40: op1_09_inv05 = 1;
    43: op1_09_inv05 = 1;
    47: op1_09_inv05 = 1;
    50: op1_09_inv05 = 1;
    52: op1_09_inv05 = 1;
    55: op1_09_inv05 = 1;
    56: op1_09_inv05 = 1;
    58: op1_09_inv05 = 1;
    59: op1_09_inv05 = 1;
    60: op1_09_inv05 = 1;
    61: op1_09_inv05 = 1;
    64: op1_09_inv05 = 1;
    65: op1_09_inv05 = 1;
    66: op1_09_inv05 = 1;
    69: op1_09_inv05 = 1;
    70: op1_09_inv05 = 1;
    72: op1_09_inv05 = 1;
    74: op1_09_inv05 = 1;
    77: op1_09_inv05 = 1;
    78: op1_09_inv05 = 1;
    79: op1_09_inv05 = 1;
    81: op1_09_inv05 = 1;
    83: op1_09_inv05 = 1;
    84: op1_09_inv05 = 1;
    85: op1_09_inv05 = 1;
    89: op1_09_inv05 = 1;
    90: op1_09_inv05 = 1;
    93: op1_09_inv05 = 1;
    94: op1_09_inv05 = 1;
    97: op1_09_inv05 = 1;
    default: op1_09_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in06 = reg_0702;
    6: op1_09_in06 = reg_0141;
    7: op1_09_in06 = reg_0450;
    8: op1_09_in06 = reg_0974;
    9: op1_09_in06 = reg_0710;
    10: op1_09_in06 = imem05_in[55:52];
    11: op1_09_in06 = reg_0463;
    12: op1_09_in06 = reg_0491;
    13: op1_09_in06 = imem02_in[43:40];
    14: op1_09_in06 = imem03_in[11:8];
    15: op1_09_in06 = imem05_in[87:84];
    16: op1_09_in06 = reg_0685;
    77: op1_09_in06 = reg_0685;
    4: op1_09_in06 = reg_0445;
    17: op1_09_in06 = reg_0113;
    18: op1_09_in06 = reg_0697;
    19: op1_09_in06 = reg_1034;
    20: op1_09_in06 = reg_0694;
    21: op1_09_in06 = reg_0639;
    22: op1_09_in06 = imem07_in[111:108];
    23: op1_09_in06 = reg_0781;
    24: op1_09_in06 = reg_0752;
    25: op1_09_in06 = reg_0686;
    30: op1_09_in06 = reg_0686;
    26: op1_09_in06 = reg_0994;
    27: op1_09_in06 = reg_0688;
    28: op1_09_in06 = imem02_in[59:56];
    29: op1_09_in06 = imem00_in[115:112];
    31: op1_09_in06 = reg_0290;
    32: op1_09_in06 = reg_0283;
    33: op1_09_in06 = reg_0614;
    95: op1_09_in06 = reg_0614;
    34: op1_09_in06 = reg_0687;
    35: op1_09_in06 = reg_0525;
    36: op1_09_in06 = reg_0063;
    37: op1_09_in06 = reg_0145;
    38: op1_09_in06 = imem04_in[27:24];
    39: op1_09_in06 = imem07_in[31:28];
    40: op1_09_in06 = reg_0696;
    41: op1_09_in06 = reg_0672;
    42: op1_09_in06 = imem04_in[11:8];
    82: op1_09_in06 = imem04_in[11:8];
    43: op1_09_in06 = reg_0971;
    44: op1_09_in06 = reg_0838;
    45: op1_09_in06 = imem02_in[35:32];
    46: op1_09_in06 = reg_0062;
    47: op1_09_in06 = reg_0029;
    48: op1_09_in06 = reg_0657;
    49: op1_09_in06 = reg_1001;
    50: op1_09_in06 = reg_1041;
    51: op1_09_in06 = imem00_in[127:124];
    52: op1_09_in06 = reg_0161;
    53: op1_09_in06 = reg_0683;
    54: op1_09_in06 = imem00_in[107:104];
    55: op1_09_in06 = reg_0818;
    56: op1_09_in06 = reg_0083;
    57: op1_09_in06 = reg_0012;
    58: op1_09_in06 = reg_0265;
    73: op1_09_in06 = reg_0265;
    59: op1_09_in06 = reg_0313;
    60: op1_09_in06 = reg_0757;
    61: op1_09_in06 = reg_0136;
    62: op1_09_in06 = reg_0708;
    63: op1_09_in06 = reg_0117;
    64: op1_09_in06 = imem02_in[39:36];
    65: op1_09_in06 = reg_0547;
    66: op1_09_in06 = imem04_in[87:84];
    67: op1_09_in06 = reg_0990;
    68: op1_09_in06 = reg_0222;
    69: op1_09_in06 = reg_0472;
    70: op1_09_in06 = reg_0568;
    71: op1_09_in06 = reg_1046;
    72: op1_09_in06 = reg_0827;
    74: op1_09_in06 = reg_0988;
    75: op1_09_in06 = imem06_in[67:64];
    78: op1_09_in06 = reg_0457;
    79: op1_09_in06 = reg_0103;
    80: op1_09_in06 = reg_0732;
    81: op1_09_in06 = reg_0736;
    83: op1_09_in06 = imem02_in[11:8];
    84: op1_09_in06 = imem07_in[19:16];
    85: op1_09_in06 = reg_0991;
    86: op1_09_in06 = reg_0970;
    87: op1_09_in06 = reg_0883;
    88: op1_09_in06 = reg_0372;
    89: op1_09_in06 = reg_0842;
    90: op1_09_in06 = reg_0007;
    91: op1_09_in06 = reg_0086;
    92: op1_09_in06 = reg_0224;
    93: op1_09_in06 = imem07_in[103:100];
    94: op1_09_in06 = reg_0382;
    96: op1_09_in06 = imem00_in[95:92];
    97: op1_09_in06 = reg_0795;
    default: op1_09_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv06 = 1;
    7: op1_09_inv06 = 1;
    8: op1_09_inv06 = 1;
    9: op1_09_inv06 = 1;
    10: op1_09_inv06 = 1;
    11: op1_09_inv06 = 1;
    13: op1_09_inv06 = 1;
    4: op1_09_inv06 = 1;
    18: op1_09_inv06 = 1;
    19: op1_09_inv06 = 1;
    21: op1_09_inv06 = 1;
    23: op1_09_inv06 = 1;
    24: op1_09_inv06 = 1;
    25: op1_09_inv06 = 1;
    26: op1_09_inv06 = 1;
    28: op1_09_inv06 = 1;
    29: op1_09_inv06 = 1;
    33: op1_09_inv06 = 1;
    37: op1_09_inv06 = 1;
    40: op1_09_inv06 = 1;
    42: op1_09_inv06 = 1;
    45: op1_09_inv06 = 1;
    47: op1_09_inv06 = 1;
    50: op1_09_inv06 = 1;
    52: op1_09_inv06 = 1;
    58: op1_09_inv06 = 1;
    60: op1_09_inv06 = 1;
    62: op1_09_inv06 = 1;
    63: op1_09_inv06 = 1;
    64: op1_09_inv06 = 1;
    65: op1_09_inv06 = 1;
    67: op1_09_inv06 = 1;
    68: op1_09_inv06 = 1;
    69: op1_09_inv06 = 1;
    71: op1_09_inv06 = 1;
    72: op1_09_inv06 = 1;
    77: op1_09_inv06 = 1;
    78: op1_09_inv06 = 1;
    79: op1_09_inv06 = 1;
    80: op1_09_inv06 = 1;
    82: op1_09_inv06 = 1;
    85: op1_09_inv06 = 1;
    86: op1_09_inv06 = 1;
    87: op1_09_inv06 = 1;
    88: op1_09_inv06 = 1;
    89: op1_09_inv06 = 1;
    92: op1_09_inv06 = 1;
    94: op1_09_inv06 = 1;
    95: op1_09_inv06 = 1;
    96: op1_09_inv06 = 1;
    default: op1_09_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in07 = reg_0426;
    6: op1_09_in07 = reg_0130;
    7: op1_09_in07 = reg_0457;
    8: op1_09_in07 = reg_0977;
    9: op1_09_in07 = reg_0725;
    10: op1_09_in07 = imem05_in[75:72];
    11: op1_09_in07 = reg_0451;
    12: op1_09_in07 = reg_0244;
    13: op1_09_in07 = imem02_in[91:88];
    14: op1_09_in07 = imem03_in[39:36];
    15: op1_09_in07 = reg_0944;
    16: op1_09_in07 = reg_0680;
    4: op1_09_in07 = reg_0434;
    17: op1_09_in07 = imem02_in[35:32];
    18: op1_09_in07 = reg_0676;
    19: op1_09_in07 = reg_0111;
    20: op1_09_in07 = reg_0686;
    21: op1_09_in07 = reg_0643;
    22: op1_09_in07 = reg_0702;
    23: op1_09_in07 = reg_0782;
    24: op1_09_in07 = reg_0780;
    25: op1_09_in07 = reg_0691;
    26: op1_09_in07 = imem04_in[27:24];
    42: op1_09_in07 = imem04_in[27:24];
    27: op1_09_in07 = reg_0455;
    28: op1_09_in07 = reg_0658;
    80: op1_09_in07 = reg_0658;
    29: op1_09_in07 = reg_0682;
    30: op1_09_in07 = reg_0679;
    31: op1_09_in07 = reg_0818;
    32: op1_09_in07 = reg_0043;
    33: op1_09_in07 = reg_0611;
    34: op1_09_in07 = reg_0453;
    35: op1_09_in07 = reg_0748;
    36: op1_09_in07 = reg_0070;
    37: op1_09_in07 = reg_0152;
    38: op1_09_in07 = imem04_in[39:36];
    39: op1_09_in07 = imem07_in[39:36];
    40: op1_09_in07 = reg_0672;
    41: op1_09_in07 = reg_0694;
    43: op1_09_in07 = reg_0964;
    44: op1_09_in07 = reg_0175;
    45: op1_09_in07 = imem02_in[63:60];
    46: op1_09_in07 = reg_0259;
    47: op1_09_in07 = imem07_in[19:16];
    48: op1_09_in07 = reg_0653;
    49: op1_09_in07 = reg_0978;
    50: op1_09_in07 = reg_0304;
    51: op1_09_in07 = reg_0693;
    52: op1_09_in07 = reg_0169;
    53: op1_09_in07 = reg_0685;
    54: op1_09_in07 = imem00_in[115:112];
    55: op1_09_in07 = reg_0037;
    56: op1_09_in07 = reg_0792;
    57: op1_09_in07 = reg_0345;
    58: op1_09_in07 = reg_0306;
    59: op1_09_in07 = reg_0568;
    60: op1_09_in07 = reg_0252;
    61: op1_09_in07 = reg_0133;
    62: op1_09_in07 = reg_0713;
    63: op1_09_in07 = reg_0363;
    64: op1_09_in07 = imem02_in[47:44];
    83: op1_09_in07 = imem02_in[47:44];
    65: op1_09_in07 = reg_0240;
    66: op1_09_in07 = reg_0483;
    67: op1_09_in07 = reg_0976;
    68: op1_09_in07 = reg_0348;
    69: op1_09_in07 = reg_0480;
    70: op1_09_in07 = reg_0850;
    71: op1_09_in07 = reg_0333;
    72: op1_09_in07 = reg_0877;
    73: op1_09_in07 = reg_0937;
    74: op1_09_in07 = imem04_in[3:0];
    75: op1_09_in07 = reg_1019;
    77: op1_09_in07 = reg_0670;
    78: op1_09_in07 = reg_0464;
    79: op1_09_in07 = reg_0110;
    81: op1_09_in07 = reg_0970;
    82: op1_09_in07 = imem04_in[15:12];
    84: op1_09_in07 = imem07_in[23:20];
    85: op1_09_in07 = reg_0979;
    86: op1_09_in07 = reg_0486;
    87: op1_09_in07 = reg_0674;
    88: op1_09_in07 = reg_0054;
    89: op1_09_in07 = reg_0356;
    90: op1_09_in07 = reg_0346;
    91: op1_09_in07 = reg_0367;
    92: op1_09_in07 = reg_0586;
    93: op1_09_in07 = reg_0567;
    94: op1_09_in07 = reg_0029;
    95: op1_09_in07 = reg_0729;
    96: op1_09_in07 = reg_0857;
    97: op1_09_in07 = reg_0950;
    default: op1_09_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv07 = 1;
    6: op1_09_inv07 = 1;
    7: op1_09_inv07 = 1;
    8: op1_09_inv07 = 1;
    9: op1_09_inv07 = 1;
    11: op1_09_inv07 = 1;
    12: op1_09_inv07 = 1;
    13: op1_09_inv07 = 1;
    15: op1_09_inv07 = 1;
    19: op1_09_inv07 = 1;
    20: op1_09_inv07 = 1;
    24: op1_09_inv07 = 1;
    25: op1_09_inv07 = 1;
    26: op1_09_inv07 = 1;
    28: op1_09_inv07 = 1;
    32: op1_09_inv07 = 1;
    35: op1_09_inv07 = 1;
    37: op1_09_inv07 = 1;
    40: op1_09_inv07 = 1;
    44: op1_09_inv07 = 1;
    45: op1_09_inv07 = 1;
    46: op1_09_inv07 = 1;
    51: op1_09_inv07 = 1;
    59: op1_09_inv07 = 1;
    61: op1_09_inv07 = 1;
    62: op1_09_inv07 = 1;
    63: op1_09_inv07 = 1;
    64: op1_09_inv07 = 1;
    66: op1_09_inv07 = 1;
    67: op1_09_inv07 = 1;
    68: op1_09_inv07 = 1;
    72: op1_09_inv07 = 1;
    75: op1_09_inv07 = 1;
    78: op1_09_inv07 = 1;
    80: op1_09_inv07 = 1;
    81: op1_09_inv07 = 1;
    82: op1_09_inv07 = 1;
    85: op1_09_inv07 = 1;
    86: op1_09_inv07 = 1;
    87: op1_09_inv07 = 1;
    88: op1_09_inv07 = 1;
    89: op1_09_inv07 = 1;
    90: op1_09_inv07 = 1;
    91: op1_09_inv07 = 1;
    92: op1_09_inv07 = 1;
    93: op1_09_inv07 = 1;
    default: op1_09_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in08 = reg_0181;
    6: op1_09_in08 = imem06_in[3:0];
    97: op1_09_in08 = imem06_in[3:0];
    7: op1_09_in08 = reg_0469;
    11: op1_09_in08 = reg_0469;
    8: op1_09_in08 = reg_0983;
    9: op1_09_in08 = reg_0714;
    10: op1_09_in08 = imem05_in[99:96];
    12: op1_09_in08 = reg_1046;
    13: op1_09_in08 = imem02_in[95:92];
    14: op1_09_in08 = imem03_in[63:60];
    15: op1_09_in08 = reg_0959;
    16: op1_09_in08 = reg_0688;
    40: op1_09_in08 = reg_0688;
    4: op1_09_in08 = reg_0427;
    17: op1_09_in08 = imem02_in[59:56];
    18: op1_09_in08 = reg_0674;
    25: op1_09_in08 = reg_0674;
    89: op1_09_in08 = reg_0674;
    19: op1_09_in08 = reg_0118;
    96: op1_09_in08 = reg_0118;
    20: op1_09_in08 = reg_0690;
    21: op1_09_in08 = reg_0328;
    22: op1_09_in08 = reg_0708;
    23: op1_09_in08 = reg_0754;
    24: op1_09_in08 = reg_0802;
    26: op1_09_in08 = reg_0301;
    66: op1_09_in08 = reg_0301;
    27: op1_09_in08 = reg_0457;
    28: op1_09_in08 = reg_0653;
    29: op1_09_in08 = reg_0681;
    30: op1_09_in08 = reg_0677;
    31: op1_09_in08 = reg_0338;
    32: op1_09_in08 = reg_0856;
    33: op1_09_in08 = reg_0618;
    34: op1_09_in08 = reg_0481;
    35: op1_09_in08 = reg_0736;
    36: op1_09_in08 = reg_0882;
    37: op1_09_in08 = reg_0143;
    38: op1_09_in08 = imem04_in[79:76];
    39: op1_09_in08 = imem07_in[59:56];
    41: op1_09_in08 = reg_0689;
    42: op1_09_in08 = imem04_in[71:68];
    43: op1_09_in08 = reg_0953;
    44: op1_09_in08 = reg_0180;
    45: op1_09_in08 = reg_0916;
    46: op1_09_in08 = reg_0364;
    47: op1_09_in08 = imem07_in[35:32];
    48: op1_09_in08 = reg_0651;
    49: op1_09_in08 = reg_0989;
    50: op1_09_in08 = reg_0105;
    51: op1_09_in08 = reg_0676;
    52: op1_09_in08 = reg_0160;
    53: op1_09_in08 = reg_0698;
    54: op1_09_in08 = imem00_in[119:116];
    55: op1_09_in08 = reg_0085;
    56: op1_09_in08 = reg_0506;
    57: op1_09_in08 = reg_0245;
    58: op1_09_in08 = reg_0055;
    59: op1_09_in08 = reg_0058;
    60: op1_09_in08 = reg_0094;
    61: op1_09_in08 = reg_0134;
    62: op1_09_in08 = reg_0707;
    63: op1_09_in08 = reg_0035;
    64: op1_09_in08 = imem02_in[67:64];
    65: op1_09_in08 = reg_0823;
    90: op1_09_in08 = reg_0823;
    67: op1_09_in08 = imem04_in[7:4];
    68: op1_09_in08 = reg_0780;
    69: op1_09_in08 = reg_0452;
    70: op1_09_in08 = reg_0076;
    71: op1_09_in08 = reg_0136;
    72: op1_09_in08 = reg_0745;
    73: op1_09_in08 = reg_0050;
    74: op1_09_in08 = imem04_in[39:36];
    75: op1_09_in08 = reg_0696;
    77: op1_09_in08 = reg_0668;
    78: op1_09_in08 = reg_0477;
    79: op1_09_in08 = imem02_in[19:16];
    80: op1_09_in08 = reg_0517;
    81: op1_09_in08 = reg_0135;
    82: op1_09_in08 = imem04_in[27:24];
    83: op1_09_in08 = imem02_in[55:52];
    84: op1_09_in08 = imem07_in[83:80];
    85: op1_09_in08 = reg_0977;
    86: op1_09_in08 = reg_0950;
    87: op1_09_in08 = reg_0102;
    88: op1_09_in08 = reg_0086;
    91: op1_09_in08 = imem03_in[23:20];
    92: op1_09_in08 = reg_0850;
    93: op1_09_in08 = reg_0710;
    94: op1_09_in08 = reg_0011;
    95: op1_09_in08 = reg_0510;
    default: op1_09_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv08 = 1;
    12: op1_09_inv08 = 1;
    15: op1_09_inv08 = 1;
    16: op1_09_inv08 = 1;
    17: op1_09_inv08 = 1;
    19: op1_09_inv08 = 1;
    20: op1_09_inv08 = 1;
    22: op1_09_inv08 = 1;
    24: op1_09_inv08 = 1;
    29: op1_09_inv08 = 1;
    33: op1_09_inv08 = 1;
    36: op1_09_inv08 = 1;
    39: op1_09_inv08 = 1;
    40: op1_09_inv08 = 1;
    41: op1_09_inv08 = 1;
    45: op1_09_inv08 = 1;
    47: op1_09_inv08 = 1;
    51: op1_09_inv08 = 1;
    53: op1_09_inv08 = 1;
    54: op1_09_inv08 = 1;
    60: op1_09_inv08 = 1;
    63: op1_09_inv08 = 1;
    64: op1_09_inv08 = 1;
    67: op1_09_inv08 = 1;
    69: op1_09_inv08 = 1;
    70: op1_09_inv08 = 1;
    73: op1_09_inv08 = 1;
    74: op1_09_inv08 = 1;
    77: op1_09_inv08 = 1;
    80: op1_09_inv08 = 1;
    81: op1_09_inv08 = 1;
    82: op1_09_inv08 = 1;
    84: op1_09_inv08 = 1;
    90: op1_09_inv08 = 1;
    93: op1_09_inv08 = 1;
    95: op1_09_inv08 = 1;
    97: op1_09_inv08 = 1;
    default: op1_09_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in09 = reg_0182;
    6: op1_09_in09 = imem06_in[19:16];
    7: op1_09_in09 = reg_0471;
    8: op1_09_in09 = reg_0994;
    9: op1_09_in09 = reg_0712;
    10: op1_09_in09 = imem05_in[111:108];
    11: op1_09_in09 = reg_0474;
    12: op1_09_in09 = reg_0958;
    13: op1_09_in09 = imem02_in[107:104];
    14: op1_09_in09 = imem03_in[95:92];
    15: op1_09_in09 = reg_0954;
    16: op1_09_in09 = reg_0673;
    4: op1_09_in09 = reg_0435;
    17: op1_09_in09 = imem02_in[91:88];
    18: op1_09_in09 = reg_0671;
    19: op1_09_in09 = reg_0099;
    20: op1_09_in09 = reg_0691;
    30: op1_09_in09 = reg_0691;
    21: op1_09_in09 = imem02_in[7:4];
    22: op1_09_in09 = reg_0709;
    23: op1_09_in09 = reg_0798;
    24: op1_09_in09 = reg_0025;
    25: op1_09_in09 = reg_0675;
    26: op1_09_in09 = reg_0530;
    27: op1_09_in09 = reg_0452;
    28: op1_09_in09 = reg_0664;
    29: op1_09_in09 = reg_0685;
    31: op1_09_in09 = reg_0336;
    32: op1_09_in09 = imem05_in[15:12];
    33: op1_09_in09 = reg_0622;
    34: op1_09_in09 = reg_0473;
    35: op1_09_in09 = reg_0517;
    36: op1_09_in09 = reg_0732;
    37: op1_09_in09 = reg_0138;
    38: op1_09_in09 = imem04_in[103:100];
    39: op1_09_in09 = imem07_in[67:64];
    40: op1_09_in09 = reg_0469;
    41: op1_09_in09 = reg_0668;
    42: op1_09_in09 = imem04_in[83:80];
    43: op1_09_in09 = reg_0826;
    44: op1_09_in09 = reg_0162;
    45: op1_09_in09 = reg_0863;
    46: op1_09_in09 = reg_0585;
    47: op1_09_in09 = imem07_in[47:44];
    48: op1_09_in09 = reg_0636;
    49: op1_09_in09 = reg_0997;
    50: op1_09_in09 = reg_0111;
    51: op1_09_in09 = reg_0677;
    52: op1_09_in09 = reg_0163;
    53: op1_09_in09 = reg_0686;
    54: op1_09_in09 = reg_0693;
    55: op1_09_in09 = reg_0792;
    56: op1_09_in09 = reg_0310;
    57: op1_09_in09 = reg_0577;
    58: op1_09_in09 = reg_0292;
    59: op1_09_in09 = reg_0056;
    60: op1_09_in09 = reg_0819;
    61: op1_09_in09 = reg_0593;
    62: op1_09_in09 = reg_0727;
    63: op1_09_in09 = reg_0634;
    64: op1_09_in09 = imem02_in[123:120];
    65: op1_09_in09 = reg_0051;
    66: op1_09_in09 = reg_0265;
    67: op1_09_in09 = imem04_in[51:48];
    74: op1_09_in09 = imem04_in[51:48];
    68: op1_09_in09 = reg_1028;
    69: op1_09_in09 = reg_0189;
    78: op1_09_in09 = reg_0189;
    70: op1_09_in09 = reg_0068;
    71: op1_09_in09 = reg_0156;
    72: op1_09_in09 = reg_0110;
    73: op1_09_in09 = reg_0313;
    75: op1_09_in09 = reg_1018;
    77: op1_09_in09 = reg_0461;
    79: op1_09_in09 = imem02_in[55:52];
    80: op1_09_in09 = imem05_in[19:16];
    81: op1_09_in09 = reg_0706;
    82: op1_09_in09 = imem04_in[43:40];
    83: op1_09_in09 = imem02_in[63:60];
    84: op1_09_in09 = imem07_in[91:88];
    85: op1_09_in09 = reg_0990;
    86: op1_09_in09 = reg_0151;
    87: op1_09_in09 = reg_0669;
    88: op1_09_in09 = reg_0885;
    89: op1_09_in09 = reg_0453;
    90: op1_09_in09 = reg_0238;
    91: op1_09_in09 = imem03_in[67:64];
    92: op1_09_in09 = reg_0764;
    93: op1_09_in09 = reg_0721;
    94: op1_09_in09 = reg_0289;
    95: op1_09_in09 = reg_0380;
    96: op1_09_in09 = reg_0899;
    97: op1_09_in09 = imem06_in[7:4];
    default: op1_09_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_09_inv09 = 1;
    9: op1_09_inv09 = 1;
    10: op1_09_inv09 = 1;
    11: op1_09_inv09 = 1;
    13: op1_09_inv09 = 1;
    14: op1_09_inv09 = 1;
    15: op1_09_inv09 = 1;
    16: op1_09_inv09 = 1;
    4: op1_09_inv09 = 1;
    17: op1_09_inv09 = 1;
    18: op1_09_inv09 = 1;
    19: op1_09_inv09 = 1;
    21: op1_09_inv09 = 1;
    22: op1_09_inv09 = 1;
    23: op1_09_inv09 = 1;
    24: op1_09_inv09 = 1;
    29: op1_09_inv09 = 1;
    32: op1_09_inv09 = 1;
    35: op1_09_inv09 = 1;
    36: op1_09_inv09 = 1;
    42: op1_09_inv09 = 1;
    43: op1_09_inv09 = 1;
    45: op1_09_inv09 = 1;
    46: op1_09_inv09 = 1;
    47: op1_09_inv09 = 1;
    49: op1_09_inv09 = 1;
    51: op1_09_inv09 = 1;
    55: op1_09_inv09 = 1;
    56: op1_09_inv09 = 1;
    57: op1_09_inv09 = 1;
    60: op1_09_inv09 = 1;
    61: op1_09_inv09 = 1;
    64: op1_09_inv09 = 1;
    66: op1_09_inv09 = 1;
    67: op1_09_inv09 = 1;
    68: op1_09_inv09 = 1;
    70: op1_09_inv09 = 1;
    73: op1_09_inv09 = 1;
    79: op1_09_inv09 = 1;
    80: op1_09_inv09 = 1;
    81: op1_09_inv09 = 1;
    82: op1_09_inv09 = 1;
    83: op1_09_inv09 = 1;
    86: op1_09_inv09 = 1;
    87: op1_09_inv09 = 1;
    90: op1_09_inv09 = 1;
    93: op1_09_inv09 = 1;
    94: op1_09_inv09 = 1;
    95: op1_09_inv09 = 1;
    97: op1_09_inv09 = 1;
    default: op1_09_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in10 = reg_0166;
    6: op1_09_in10 = imem06_in[67:64];
    7: op1_09_in10 = reg_0191;
    8: op1_09_in10 = imem04_in[11:8];
    9: op1_09_in10 = reg_0709;
    10: op1_09_in10 = reg_0271;
    11: op1_09_in10 = reg_0193;
    69: op1_09_in10 = reg_0193;
    78: op1_09_in10 = reg_0193;
    12: op1_09_in10 = reg_0959;
    13: op1_09_in10 = imem02_in[127:124];
    14: op1_09_in10 = reg_0599;
    15: op1_09_in10 = reg_0964;
    16: op1_09_in10 = reg_0455;
    4: op1_09_in10 = reg_0183;
    17: op1_09_in10 = imem02_in[115:112];
    18: op1_09_in10 = reg_0465;
    41: op1_09_in10 = reg_0465;
    19: op1_09_in10 = reg_0114;
    20: op1_09_in10 = reg_0680;
    21: op1_09_in10 = imem02_in[31:28];
    22: op1_09_in10 = reg_0713;
    23: op1_09_in10 = imem07_in[7:4];
    24: op1_09_in10 = reg_0018;
    25: op1_09_in10 = reg_0463;
    26: op1_09_in10 = reg_0539;
    27: op1_09_in10 = reg_0458;
    28: op1_09_in10 = reg_0656;
    29: op1_09_in10 = reg_0684;
    30: op1_09_in10 = reg_0453;
    31: op1_09_in10 = reg_0758;
    32: op1_09_in10 = imem05_in[35:32];
    33: op1_09_in10 = reg_0356;
    34: op1_09_in10 = reg_0214;
    35: op1_09_in10 = reg_0777;
    92: op1_09_in10 = reg_0777;
    36: op1_09_in10 = reg_0054;
    37: op1_09_in10 = reg_0141;
    38: op1_09_in10 = imem04_in[115:112];
    39: op1_09_in10 = imem07_in[83:80];
    40: op1_09_in10 = reg_0460;
    42: op1_09_in10 = reg_0525;
    43: op1_09_in10 = reg_0022;
    44: op1_09_in10 = reg_0170;
    45: op1_09_in10 = reg_0290;
    46: op1_09_in10 = reg_0579;
    47: op1_09_in10 = reg_0704;
    48: op1_09_in10 = reg_0045;
    49: op1_09_in10 = reg_0555;
    50: op1_09_in10 = reg_0104;
    51: op1_09_in10 = reg_0674;
    53: op1_09_in10 = reg_0688;
    54: op1_09_in10 = reg_0696;
    55: op1_09_in10 = reg_0405;
    68: op1_09_in10 = reg_0405;
    56: op1_09_in10 = imem03_in[31:28];
    57: op1_09_in10 = reg_0661;
    58: op1_09_in10 = reg_0540;
    59: op1_09_in10 = reg_0584;
    70: op1_09_in10 = reg_0584;
    60: op1_09_in10 = reg_0438;
    61: op1_09_in10 = reg_0759;
    62: op1_09_in10 = reg_0325;
    63: op1_09_in10 = reg_0857;
    64: op1_09_in10 = reg_0810;
    65: op1_09_in10 = reg_0376;
    66: op1_09_in10 = reg_0937;
    67: op1_09_in10 = imem04_in[67:64];
    71: op1_09_in10 = reg_0138;
    72: op1_09_in10 = reg_0657;
    73: op1_09_in10 = reg_0058;
    74: op1_09_in10 = imem04_in[63:60];
    75: op1_09_in10 = reg_0267;
    77: op1_09_in10 = reg_0211;
    79: op1_09_in10 = imem02_in[63:60];
    80: op1_09_in10 = imem05_in[43:40];
    81: op1_09_in10 = reg_0258;
    82: op1_09_in10 = imem04_in[79:76];
    83: op1_09_in10 = imem02_in[107:104];
    84: op1_09_in10 = imem07_in[103:100];
    85: op1_09_in10 = imem04_in[23:20];
    86: op1_09_in10 = reg_0631;
    87: op1_09_in10 = reg_0461;
    88: op1_09_in10 = reg_0082;
    89: op1_09_in10 = reg_0207;
    90: op1_09_in10 = reg_0596;
    91: op1_09_in10 = imem03_in[87:84];
    93: op1_09_in10 = reg_0164;
    94: op1_09_in10 = reg_0370;
    95: op1_09_in10 = reg_0811;
    96: op1_09_in10 = reg_0310;
    97: op1_09_in10 = imem06_in[31:28];
    default: op1_09_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv10 = 1;
    6: op1_09_inv10 = 1;
    8: op1_09_inv10 = 1;
    9: op1_09_inv10 = 1;
    10: op1_09_inv10 = 1;
    11: op1_09_inv10 = 1;
    12: op1_09_inv10 = 1;
    13: op1_09_inv10 = 1;
    15: op1_09_inv10 = 1;
    4: op1_09_inv10 = 1;
    17: op1_09_inv10 = 1;
    18: op1_09_inv10 = 1;
    20: op1_09_inv10 = 1;
    21: op1_09_inv10 = 1;
    23: op1_09_inv10 = 1;
    24: op1_09_inv10 = 1;
    26: op1_09_inv10 = 1;
    27: op1_09_inv10 = 1;
    28: op1_09_inv10 = 1;
    29: op1_09_inv10 = 1;
    30: op1_09_inv10 = 1;
    32: op1_09_inv10 = 1;
    33: op1_09_inv10 = 1;
    40: op1_09_inv10 = 1;
    44: op1_09_inv10 = 1;
    46: op1_09_inv10 = 1;
    47: op1_09_inv10 = 1;
    49: op1_09_inv10 = 1;
    50: op1_09_inv10 = 1;
    56: op1_09_inv10 = 1;
    58: op1_09_inv10 = 1;
    60: op1_09_inv10 = 1;
    61: op1_09_inv10 = 1;
    63: op1_09_inv10 = 1;
    65: op1_09_inv10 = 1;
    66: op1_09_inv10 = 1;
    68: op1_09_inv10 = 1;
    70: op1_09_inv10 = 1;
    74: op1_09_inv10 = 1;
    77: op1_09_inv10 = 1;
    78: op1_09_inv10 = 1;
    79: op1_09_inv10 = 1;
    80: op1_09_inv10 = 1;
    82: op1_09_inv10 = 1;
    87: op1_09_inv10 = 1;
    89: op1_09_inv10 = 1;
    90: op1_09_inv10 = 1;
    92: op1_09_inv10 = 1;
    94: op1_09_inv10 = 1;
    default: op1_09_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の11番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in11 = reg_0628;
    7: op1_09_in11 = reg_0212;
    11: op1_09_in11 = reg_0212;
    8: op1_09_in11 = imem04_in[15:12];
    9: op1_09_in11 = reg_0701;
    10: op1_09_in11 = reg_0259;
    12: op1_09_in11 = reg_0956;
    13: op1_09_in11 = reg_0648;
    14: op1_09_in11 = reg_0583;
    15: op1_09_in11 = reg_0949;
    16: op1_09_in11 = reg_0476;
    87: op1_09_in11 = reg_0476;
    4: op1_09_in11 = reg_0168;
    17: op1_09_in11 = reg_0647;
    18: op1_09_in11 = reg_0469;
    19: op1_09_in11 = reg_0113;
    20: op1_09_in11 = reg_0459;
    21: op1_09_in11 = imem03_in[7:4];
    22: op1_09_in11 = reg_0441;
    23: op1_09_in11 = imem07_in[23:20];
    24: op1_09_in11 = reg_0805;
    25: op1_09_in11 = reg_0457;
    26: op1_09_in11 = reg_0292;
    27: op1_09_in11 = reg_0188;
    28: op1_09_in11 = reg_0644;
    29: op1_09_in11 = reg_0690;
    30: op1_09_in11 = reg_0481;
    31: op1_09_in11 = reg_0261;
    32: op1_09_in11 = imem05_in[55:52];
    33: op1_09_in11 = reg_0914;
    34: op1_09_in11 = reg_0208;
    35: op1_09_in11 = reg_0286;
    36: op1_09_in11 = reg_0736;
    37: op1_09_in11 = reg_0130;
    38: op1_09_in11 = reg_0483;
    82: op1_09_in11 = reg_0483;
    39: op1_09_in11 = imem07_in[99:96];
    40: op1_09_in11 = reg_0473;
    41: op1_09_in11 = reg_0450;
    42: op1_09_in11 = reg_0528;
    43: op1_09_in11 = reg_0260;
    45: op1_09_in11 = reg_0886;
    46: op1_09_in11 = reg_0301;
    47: op1_09_in11 = reg_0719;
    48: op1_09_in11 = reg_0818;
    49: op1_09_in11 = reg_0499;
    50: op1_09_in11 = reg_0112;
    51: op1_09_in11 = reg_0678;
    53: op1_09_in11 = reg_0464;
    54: op1_09_in11 = reg_0698;
    55: op1_09_in11 = reg_0677;
    56: op1_09_in11 = imem03_in[43:40];
    57: op1_09_in11 = reg_0767;
    58: op1_09_in11 = reg_0524;
    59: op1_09_in11 = reg_0401;
    60: op1_09_in11 = reg_0497;
    61: op1_09_in11 = reg_0845;
    62: op1_09_in11 = reg_0426;
    63: op1_09_in11 = reg_0642;
    64: op1_09_in11 = reg_0741;
    65: op1_09_in11 = reg_0312;
    66: op1_09_in11 = reg_0277;
    67: op1_09_in11 = imem04_in[71:68];
    68: op1_09_in11 = reg_0449;
    69: op1_09_in11 = reg_0207;
    70: op1_09_in11 = reg_0808;
    73: op1_09_in11 = reg_0808;
    71: op1_09_in11 = reg_0594;
    72: op1_09_in11 = reg_0621;
    74: op1_09_in11 = imem04_in[75:72];
    75: op1_09_in11 = reg_0817;
    77: op1_09_in11 = imem01_in[67:64];
    78: op1_09_in11 = reg_0198;
    79: op1_09_in11 = imem02_in[107:104];
    80: op1_09_in11 = imem05_in[47:44];
    92: op1_09_in11 = imem05_in[47:44];
    81: op1_09_in11 = reg_0326;
    83: op1_09_in11 = imem02_in[123:120];
    84: op1_09_in11 = imem07_in[115:112];
    85: op1_09_in11 = imem04_in[43:40];
    86: op1_09_in11 = reg_0053;
    88: op1_09_in11 = reg_0643;
    89: op1_09_in11 = reg_0206;
    90: op1_09_in11 = reg_0579;
    91: op1_09_in11 = reg_0317;
    93: op1_09_in11 = reg_0708;
    94: op1_09_in11 = reg_0392;
    95: op1_09_in11 = reg_0133;
    96: op1_09_in11 = reg_0760;
    97: op1_09_in11 = imem06_in[47:44];
    default: op1_09_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_09_inv11 = 1;
    10: op1_09_inv11 = 1;
    11: op1_09_inv11 = 1;
    15: op1_09_inv11 = 1;
    19: op1_09_inv11 = 1;
    20: op1_09_inv11 = 1;
    21: op1_09_inv11 = 1;
    23: op1_09_inv11 = 1;
    24: op1_09_inv11 = 1;
    25: op1_09_inv11 = 1;
    26: op1_09_inv11 = 1;
    28: op1_09_inv11 = 1;
    29: op1_09_inv11 = 1;
    30: op1_09_inv11 = 1;
    37: op1_09_inv11 = 1;
    42: op1_09_inv11 = 1;
    43: op1_09_inv11 = 1;
    45: op1_09_inv11 = 1;
    47: op1_09_inv11 = 1;
    48: op1_09_inv11 = 1;
    49: op1_09_inv11 = 1;
    51: op1_09_inv11 = 1;
    53: op1_09_inv11 = 1;
    55: op1_09_inv11 = 1;
    56: op1_09_inv11 = 1;
    61: op1_09_inv11 = 1;
    62: op1_09_inv11 = 1;
    63: op1_09_inv11 = 1;
    64: op1_09_inv11 = 1;
    69: op1_09_inv11 = 1;
    72: op1_09_inv11 = 1;
    74: op1_09_inv11 = 1;
    75: op1_09_inv11 = 1;
    77: op1_09_inv11 = 1;
    80: op1_09_inv11 = 1;
    81: op1_09_inv11 = 1;
    82: op1_09_inv11 = 1;
    90: op1_09_inv11 = 1;
    94: op1_09_inv11 = 1;
    95: op1_09_inv11 = 1;
    default: op1_09_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の12番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in12 = reg_0610;
    7: op1_09_in12 = imem01_in[23:20];
    8: op1_09_in12 = imem04_in[23:20];
    9: op1_09_in12 = reg_0700;
    10: op1_09_in12 = reg_0252;
    11: op1_09_in12 = reg_0190;
    12: op1_09_in12 = reg_0951;
    13: op1_09_in12 = reg_0652;
    14: op1_09_in12 = reg_0591;
    15: op1_09_in12 = reg_0965;
    16: op1_09_in12 = reg_0479;
    17: op1_09_in12 = reg_0640;
    18: op1_09_in12 = reg_0476;
    19: op1_09_in12 = imem02_in[51:48];
    20: op1_09_in12 = reg_0191;
    21: op1_09_in12 = imem03_in[23:20];
    22: op1_09_in12 = reg_0430;
    23: op1_09_in12 = imem07_in[103:100];
    39: op1_09_in12 = imem07_in[103:100];
    24: op1_09_in12 = reg_1011;
    25: op1_09_in12 = reg_0475;
    26: op1_09_in12 = reg_1016;
    27: op1_09_in12 = reg_0203;
    28: op1_09_in12 = reg_0636;
    29: op1_09_in12 = reg_0668;
    30: op1_09_in12 = reg_0472;
    31: op1_09_in12 = reg_0049;
    32: op1_09_in12 = imem05_in[71:68];
    33: op1_09_in12 = reg_0388;
    34: op1_09_in12 = reg_0207;
    35: op1_09_in12 = reg_0044;
    36: op1_09_in12 = reg_0056;
    37: op1_09_in12 = reg_0144;
    38: op1_09_in12 = reg_1009;
    40: op1_09_in12 = reg_0470;
    41: op1_09_in12 = reg_0469;
    42: op1_09_in12 = reg_0854;
    43: op1_09_in12 = reg_0785;
    45: op1_09_in12 = reg_0772;
    46: op1_09_in12 = reg_0530;
    47: op1_09_in12 = reg_0710;
    48: op1_09_in12 = reg_0817;
    49: op1_09_in12 = reg_0301;
    50: op1_09_in12 = reg_0106;
    51: op1_09_in12 = reg_0675;
    53: op1_09_in12 = reg_0478;
    54: op1_09_in12 = reg_0689;
    55: op1_09_in12 = reg_0570;
    56: op1_09_in12 = imem03_in[95:92];
    57: op1_09_in12 = reg_0246;
    65: op1_09_in12 = reg_0246;
    58: op1_09_in12 = reg_0276;
    59: op1_09_in12 = imem04_in[31:28];
    60: op1_09_in12 = reg_0147;
    61: op1_09_in12 = reg_0690;
    62: op1_09_in12 = reg_0589;
    63: op1_09_in12 = imem02_in[31:28];
    64: op1_09_in12 = reg_0666;
    66: op1_09_in12 = reg_0912;
    67: op1_09_in12 = imem04_in[87:84];
    68: op1_09_in12 = reg_0371;
    69: op1_09_in12 = reg_0194;
    70: op1_09_in12 = reg_0809;
    71: op1_09_in12 = reg_0349;
    72: op1_09_in12 = imem02_in[23:20];
    73: op1_09_in12 = reg_0495;
    74: op1_09_in12 = imem04_in[79:76];
    75: op1_09_in12 = reg_0735;
    77: op1_09_in12 = imem01_in[83:80];
    78: op1_09_in12 = reg_0199;
    79: op1_09_in12 = imem02_in[115:112];
    80: op1_09_in12 = imem05_in[55:52];
    81: op1_09_in12 = reg_0851;
    82: op1_09_in12 = reg_0282;
    83: op1_09_in12 = reg_0813;
    84: op1_09_in12 = reg_0165;
    85: op1_09_in12 = imem04_in[103:100];
    86: op1_09_in12 = reg_0005;
    87: op1_09_in12 = reg_0471;
    88: op1_09_in12 = reg_0341;
    89: op1_09_in12 = reg_0197;
    90: op1_09_in12 = reg_0038;
    91: op1_09_in12 = reg_0761;
    92: op1_09_in12 = imem05_in[59:56];
    93: op1_09_in12 = reg_0247;
    94: op1_09_in12 = reg_0040;
    95: op1_09_in12 = reg_0084;
    96: op1_09_in12 = reg_0680;
    97: op1_09_in12 = reg_0696;
    default: op1_09_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv12 = 1;
    9: op1_09_inv12 = 1;
    12: op1_09_inv12 = 1;
    16: op1_09_inv12 = 1;
    17: op1_09_inv12 = 1;
    18: op1_09_inv12 = 1;
    19: op1_09_inv12 = 1;
    22: op1_09_inv12 = 1;
    24: op1_09_inv12 = 1;
    25: op1_09_inv12 = 1;
    27: op1_09_inv12 = 1;
    31: op1_09_inv12 = 1;
    34: op1_09_inv12 = 1;
    41: op1_09_inv12 = 1;
    42: op1_09_inv12 = 1;
    43: op1_09_inv12 = 1;
    45: op1_09_inv12 = 1;
    48: op1_09_inv12 = 1;
    51: op1_09_inv12 = 1;
    53: op1_09_inv12 = 1;
    56: op1_09_inv12 = 1;
    59: op1_09_inv12 = 1;
    60: op1_09_inv12 = 1;
    61: op1_09_inv12 = 1;
    62: op1_09_inv12 = 1;
    64: op1_09_inv12 = 1;
    65: op1_09_inv12 = 1;
    67: op1_09_inv12 = 1;
    69: op1_09_inv12 = 1;
    72: op1_09_inv12 = 1;
    75: op1_09_inv12 = 1;
    78: op1_09_inv12 = 1;
    79: op1_09_inv12 = 1;
    81: op1_09_inv12 = 1;
    82: op1_09_inv12 = 1;
    84: op1_09_inv12 = 1;
    87: op1_09_inv12 = 1;
    88: op1_09_inv12 = 1;
    90: op1_09_inv12 = 1;
    91: op1_09_inv12 = 1;
    default: op1_09_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の13番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in13 = reg_0629;
    7: op1_09_in13 = imem01_in[27:24];
    8: op1_09_in13 = imem04_in[55:52];
    9: op1_09_in13 = reg_0421;
    10: op1_09_in13 = reg_0258;
    11: op1_09_in13 = reg_0202;
    12: op1_09_in13 = reg_0946;
    13: op1_09_in13 = reg_0352;
    14: op1_09_in13 = reg_0563;
    15: op1_09_in13 = reg_0947;
    16: op1_09_in13 = reg_0214;
    17: op1_09_in13 = reg_0648;
    18: op1_09_in13 = reg_0481;
    19: op1_09_in13 = imem02_in[63:60];
    20: op1_09_in13 = reg_0209;
    21: op1_09_in13 = reg_0584;
    22: op1_09_in13 = reg_0447;
    23: op1_09_in13 = reg_0704;
    24: op1_09_in13 = imem07_in[23:20];
    25: op1_09_in13 = reg_0480;
    51: op1_09_in13 = reg_0480;
    26: op1_09_in13 = reg_0764;
    27: op1_09_in13 = imem01_in[3:0];
    78: op1_09_in13 = imem01_in[3:0];
    28: op1_09_in13 = reg_0045;
    29: op1_09_in13 = reg_0675;
    30: op1_09_in13 = reg_0470;
    31: op1_09_in13 = reg_0084;
    32: op1_09_in13 = reg_0962;
    33: op1_09_in13 = reg_0222;
    34: op1_09_in13 = reg_0213;
    35: op1_09_in13 = imem05_in[3:0];
    36: op1_09_in13 = reg_0053;
    37: op1_09_in13 = reg_0915;
    38: op1_09_in13 = reg_0277;
    39: op1_09_in13 = reg_0716;
    40: op1_09_in13 = reg_0193;
    41: op1_09_in13 = reg_0476;
    42: op1_09_in13 = reg_0777;
    43: op1_09_in13 = reg_0819;
    45: op1_09_in13 = reg_0761;
    46: op1_09_in13 = reg_0539;
    47: op1_09_in13 = reg_0723;
    48: op1_09_in13 = reg_0772;
    49: op1_09_in13 = reg_0055;
    66: op1_09_in13 = reg_0055;
    82: op1_09_in13 = reg_0055;
    50: op1_09_in13 = reg_0115;
    53: op1_09_in13 = reg_0208;
    54: op1_09_in13 = reg_0690;
    55: op1_09_in13 = imem03_in[15:12];
    56: op1_09_in13 = imem03_in[115:112];
    57: op1_09_in13 = reg_0992;
    58: op1_09_in13 = reg_0899;
    59: op1_09_in13 = imem04_in[47:44];
    60: op1_09_in13 = reg_0128;
    61: op1_09_in13 = reg_0693;
    62: op1_09_in13 = reg_0420;
    63: op1_09_in13 = imem02_in[55:52];
    64: op1_09_in13 = reg_0654;
    65: op1_09_in13 = reg_0374;
    67: op1_09_in13 = imem04_in[95:92];
    68: op1_09_in13 = reg_0264;
    69: op1_09_in13 = reg_0196;
    70: op1_09_in13 = reg_0284;
    71: op1_09_in13 = reg_0093;
    72: op1_09_in13 = imem02_in[51:48];
    73: op1_09_in13 = reg_0953;
    74: op1_09_in13 = imem04_in[119:116];
    75: op1_09_in13 = reg_0440;
    77: op1_09_in13 = imem01_in[87:84];
    79: op1_09_in13 = imem02_in[123:120];
    80: op1_09_in13 = imem05_in[71:68];
    81: op1_09_in13 = reg_0490;
    83: op1_09_in13 = reg_0896;
    84: op1_09_in13 = reg_0717;
    85: op1_09_in13 = reg_0577;
    86: op1_09_in13 = reg_0263;
    87: op1_09_in13 = reg_0468;
    88: op1_09_in13 = reg_0367;
    89: op1_09_in13 = imem01_in[19:16];
    90: op1_09_in13 = reg_0672;
    91: op1_09_in13 = reg_0836;
    92: op1_09_in13 = imem05_in[95:92];
    93: op1_09_in13 = reg_0805;
    94: op1_09_in13 = reg_0403;
    95: op1_09_in13 = imem07_in[15:12];
    96: op1_09_in13 = reg_0030;
    97: op1_09_in13 = reg_0351;
    default: op1_09_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv13 = 1;
    8: op1_09_inv13 = 1;
    11: op1_09_inv13 = 1;
    12: op1_09_inv13 = 1;
    14: op1_09_inv13 = 1;
    15: op1_09_inv13 = 1;
    18: op1_09_inv13 = 1;
    19: op1_09_inv13 = 1;
    21: op1_09_inv13 = 1;
    22: op1_09_inv13 = 1;
    23: op1_09_inv13 = 1;
    24: op1_09_inv13 = 1;
    30: op1_09_inv13 = 1;
    32: op1_09_inv13 = 1;
    34: op1_09_inv13 = 1;
    36: op1_09_inv13 = 1;
    39: op1_09_inv13 = 1;
    41: op1_09_inv13 = 1;
    42: op1_09_inv13 = 1;
    43: op1_09_inv13 = 1;
    45: op1_09_inv13 = 1;
    46: op1_09_inv13 = 1;
    47: op1_09_inv13 = 1;
    48: op1_09_inv13 = 1;
    53: op1_09_inv13 = 1;
    54: op1_09_inv13 = 1;
    55: op1_09_inv13 = 1;
    57: op1_09_inv13 = 1;
    58: op1_09_inv13 = 1;
    60: op1_09_inv13 = 1;
    61: op1_09_inv13 = 1;
    62: op1_09_inv13 = 1;
    67: op1_09_inv13 = 1;
    68: op1_09_inv13 = 1;
    69: op1_09_inv13 = 1;
    70: op1_09_inv13 = 1;
    71: op1_09_inv13 = 1;
    72: op1_09_inv13 = 1;
    73: op1_09_inv13 = 1;
    75: op1_09_inv13 = 1;
    77: op1_09_inv13 = 1;
    80: op1_09_inv13 = 1;
    82: op1_09_inv13 = 1;
    84: op1_09_inv13 = 1;
    87: op1_09_inv13 = 1;
    91: op1_09_inv13 = 1;
    94: op1_09_inv13 = 1;
    97: op1_09_inv13 = 1;
    default: op1_09_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の14番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in14 = reg_0630;
    7: op1_09_in14 = imem01_in[87:84];
    8: op1_09_in14 = imem04_in[95:92];
    9: op1_09_in14 = reg_0447;
    10: op1_09_in14 = reg_0265;
    11: op1_09_in14 = reg_0788;
    12: op1_09_in14 = reg_0953;
    13: op1_09_in14 = reg_0333;
    17: op1_09_in14 = reg_0333;
    14: op1_09_in14 = reg_0594;
    15: op1_09_in14 = reg_0960;
    16: op1_09_in14 = reg_0200;
    18: op1_09_in14 = reg_0470;
    19: op1_09_in14 = imem02_in[99:96];
    20: op1_09_in14 = reg_0207;
    21: op1_09_in14 = reg_0585;
    22: op1_09_in14 = reg_0418;
    23: op1_09_in14 = reg_0720;
    24: op1_09_in14 = imem07_in[55:52];
    25: op1_09_in14 = reg_0473;
    51: op1_09_in14 = reg_0473;
    26: op1_09_in14 = reg_0733;
    27: op1_09_in14 = imem01_in[67:64];
    28: op1_09_in14 = reg_0916;
    29: op1_09_in14 = reg_0673;
    30: op1_09_in14 = reg_0198;
    40: op1_09_in14 = reg_0198;
    31: op1_09_in14 = reg_0016;
    32: op1_09_in14 = reg_0973;
    33: op1_09_in14 = reg_0917;
    34: op1_09_in14 = reg_0195;
    35: op1_09_in14 = imem05_in[7:4];
    36: op1_09_in14 = reg_0044;
    37: op1_09_in14 = reg_0534;
    38: op1_09_in14 = reg_0540;
    39: op1_09_in14 = reg_0726;
    47: op1_09_in14 = reg_0726;
    41: op1_09_in14 = reg_0456;
    42: op1_09_in14 = imem05_in[11:8];
    43: op1_09_in14 = reg_0489;
    45: op1_09_in14 = imem03_in[7:4];
    46: op1_09_in14 = reg_0048;
    48: op1_09_in14 = reg_0758;
    49: op1_09_in14 = reg_0292;
    50: op1_09_in14 = reg_0127;
    53: op1_09_in14 = reg_0204;
    54: op1_09_in14 = reg_0688;
    55: op1_09_in14 = imem03_in[87:84];
    56: op1_09_in14 = imem03_in[119:116];
    57: op1_09_in14 = reg_0990;
    58: op1_09_in14 = reg_0554;
    59: op1_09_in14 = imem04_in[63:60];
    60: op1_09_in14 = reg_0142;
    61: op1_09_in14 = reg_0787;
    62: op1_09_in14 = reg_0640;
    63: op1_09_in14 = imem02_in[71:68];
    64: op1_09_in14 = reg_0865;
    65: op1_09_in14 = reg_0979;
    66: op1_09_in14 = reg_0050;
    67: op1_09_in14 = imem04_in[99:96];
    68: op1_09_in14 = reg_0633;
    69: op1_09_in14 = reg_0885;
    83: op1_09_in14 = reg_0885;
    70: op1_09_in14 = reg_0627;
    71: op1_09_in14 = reg_0119;
    72: op1_09_in14 = imem02_in[63:60];
    73: op1_09_in14 = imem05_in[67:64];
    74: op1_09_in14 = reg_0937;
    75: op1_09_in14 = reg_0698;
    77: op1_09_in14 = reg_0968;
    78: op1_09_in14 = imem01_in[11:8];
    79: op1_09_in14 = reg_0803;
    80: op1_09_in14 = imem05_in[83:80];
    81: op1_09_in14 = imem06_in[7:4];
    82: op1_09_in14 = reg_1016;
    84: op1_09_in14 = reg_0923;
    85: op1_09_in14 = reg_0942;
    86: op1_09_in14 = reg_0010;
    87: op1_09_in14 = reg_0479;
    88: op1_09_in14 = reg_0678;
    89: op1_09_in14 = imem01_in[47:44];
    90: op1_09_in14 = reg_0767;
    91: op1_09_in14 = reg_0049;
    92: op1_09_in14 = reg_0319;
    93: op1_09_in14 = reg_0047;
    94: op1_09_in14 = reg_0632;
    95: op1_09_in14 = imem07_in[23:20];
    96: op1_09_in14 = reg_0469;
    97: op1_09_in14 = reg_0267;
    default: op1_09_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    11: op1_09_inv14 = 1;
    17: op1_09_inv14 = 1;
    19: op1_09_inv14 = 1;
    21: op1_09_inv14 = 1;
    24: op1_09_inv14 = 1;
    32: op1_09_inv14 = 1;
    33: op1_09_inv14 = 1;
    35: op1_09_inv14 = 1;
    38: op1_09_inv14 = 1;
    39: op1_09_inv14 = 1;
    40: op1_09_inv14 = 1;
    41: op1_09_inv14 = 1;
    43: op1_09_inv14 = 1;
    47: op1_09_inv14 = 1;
    50: op1_09_inv14 = 1;
    54: op1_09_inv14 = 1;
    55: op1_09_inv14 = 1;
    57: op1_09_inv14 = 1;
    60: op1_09_inv14 = 1;
    62: op1_09_inv14 = 1;
    67: op1_09_inv14 = 1;
    85: op1_09_inv14 = 1;
    86: op1_09_inv14 = 1;
    87: op1_09_inv14 = 1;
    89: op1_09_inv14 = 1;
    90: op1_09_inv14 = 1;
    96: op1_09_inv14 = 1;
    97: op1_09_inv14 = 1;
    default: op1_09_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の15番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in15 = reg_0631;
    7: op1_09_in15 = imem01_in[111:108];
    8: op1_09_in15 = imem04_in[119:116];
    9: op1_09_in15 = reg_0419;
    10: op1_09_in15 = reg_0272;
    11: op1_09_in15 = reg_0786;
    12: op1_09_in15 = imem05_in[63:60];
    36: op1_09_in15 = imem05_in[63:60];
    13: op1_09_in15 = reg_0320;
    14: op1_09_in15 = reg_0395;
    15: op1_09_in15 = reg_0217;
    16: op1_09_in15 = reg_0186;
    20: op1_09_in15 = reg_0186;
    17: op1_09_in15 = reg_0329;
    18: op1_09_in15 = reg_0456;
    19: op1_09_in15 = imem02_in[103:100];
    21: op1_09_in15 = reg_0578;
    22: op1_09_in15 = reg_0434;
    23: op1_09_in15 = reg_0721;
    24: op1_09_in15 = imem07_in[71:68];
    25: op1_09_in15 = reg_0452;
    87: op1_09_in15 = reg_0452;
    26: op1_09_in15 = reg_0763;
    27: op1_09_in15 = imem01_in[123:120];
    28: op1_09_in15 = reg_0081;
    29: op1_09_in15 = reg_0692;
    54: op1_09_in15 = reg_0692;
    30: op1_09_in15 = reg_0212;
    31: op1_09_in15 = reg_0077;
    32: op1_09_in15 = reg_0966;
    33: op1_09_in15 = reg_0486;
    34: op1_09_in15 = reg_0199;
    35: op1_09_in15 = imem05_in[23:20];
    37: op1_09_in15 = reg_0027;
    38: op1_09_in15 = reg_0931;
    39: op1_09_in15 = reg_0717;
    40: op1_09_in15 = reg_0197;
    41: op1_09_in15 = reg_0188;
    42: op1_09_in15 = imem05_in[55:52];
    43: op1_09_in15 = reg_0128;
    45: op1_09_in15 = imem03_in[15:12];
    46: op1_09_in15 = reg_0848;
    82: op1_09_in15 = reg_0848;
    47: op1_09_in15 = reg_0361;
    48: op1_09_in15 = reg_0867;
    49: op1_09_in15 = reg_1016;
    50: op1_09_in15 = reg_0110;
    51: op1_09_in15 = reg_0470;
    53: op1_09_in15 = reg_0194;
    55: op1_09_in15 = imem03_in[111:108];
    56: op1_09_in15 = reg_0012;
    57: op1_09_in15 = imem04_in[11:8];
    58: op1_09_in15 = reg_0075;
    59: op1_09_in15 = imem04_in[75:72];
    60: op1_09_in15 = reg_0146;
    61: op1_09_in15 = reg_0573;
    62: op1_09_in15 = reg_0161;
    63: op1_09_in15 = imem02_in[87:84];
    64: op1_09_in15 = reg_0894;
    65: op1_09_in15 = reg_0980;
    66: op1_09_in15 = reg_0537;
    67: op1_09_in15 = imem04_in[103:100];
    68: op1_09_in15 = reg_0955;
    69: op1_09_in15 = reg_0100;
    70: op1_09_in15 = reg_0854;
    71: op1_09_in15 = reg_0696;
    72: op1_09_in15 = imem02_in[71:68];
    73: op1_09_in15 = imem05_in[103:100];
    74: op1_09_in15 = reg_0282;
    75: op1_09_in15 = reg_0807;
    77: op1_09_in15 = reg_0592;
    78: op1_09_in15 = imem01_in[79:76];
    79: op1_09_in15 = reg_0637;
    80: op1_09_in15 = imem05_in[95:92];
    81: op1_09_in15 = imem06_in[15:12];
    83: op1_09_in15 = reg_0260;
    84: op1_09_in15 = reg_0353;
    85: op1_09_in15 = reg_0306;
    86: op1_09_in15 = reg_1018;
    88: op1_09_in15 = reg_0396;
    89: op1_09_in15 = reg_0122;
    90: op1_09_in15 = reg_0581;
    91: op1_09_in15 = reg_0609;
    92: op1_09_in15 = reg_0013;
    93: op1_09_in15 = reg_0744;
    94: op1_09_in15 = reg_0084;
    95: op1_09_in15 = imem07_in[31:28];
    96: op1_09_in15 = reg_0472;
    97: op1_09_in15 = reg_0025;
    default: op1_09_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv15 = 1;
    9: op1_09_inv15 = 1;
    13: op1_09_inv15 = 1;
    14: op1_09_inv15 = 1;
    15: op1_09_inv15 = 1;
    18: op1_09_inv15 = 1;
    20: op1_09_inv15 = 1;
    21: op1_09_inv15 = 1;
    23: op1_09_inv15 = 1;
    25: op1_09_inv15 = 1;
    26: op1_09_inv15 = 1;
    29: op1_09_inv15 = 1;
    33: op1_09_inv15 = 1;
    35: op1_09_inv15 = 1;
    36: op1_09_inv15 = 1;
    39: op1_09_inv15 = 1;
    41: op1_09_inv15 = 1;
    42: op1_09_inv15 = 1;
    43: op1_09_inv15 = 1;
    47: op1_09_inv15 = 1;
    48: op1_09_inv15 = 1;
    49: op1_09_inv15 = 1;
    50: op1_09_inv15 = 1;
    57: op1_09_inv15 = 1;
    59: op1_09_inv15 = 1;
    60: op1_09_inv15 = 1;
    61: op1_09_inv15 = 1;
    63: op1_09_inv15 = 1;
    64: op1_09_inv15 = 1;
    65: op1_09_inv15 = 1;
    70: op1_09_inv15 = 1;
    72: op1_09_inv15 = 1;
    73: op1_09_inv15 = 1;
    74: op1_09_inv15 = 1;
    75: op1_09_inv15 = 1;
    77: op1_09_inv15 = 1;
    78: op1_09_inv15 = 1;
    79: op1_09_inv15 = 1;
    80: op1_09_inv15 = 1;
    81: op1_09_inv15 = 1;
    85: op1_09_inv15 = 1;
    87: op1_09_inv15 = 1;
    88: op1_09_inv15 = 1;
    89: op1_09_inv15 = 1;
    90: op1_09_inv15 = 1;
    95: op1_09_inv15 = 1;
    97: op1_09_inv15 = 1;
    default: op1_09_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の16番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in16 = reg_0626;
    7: op1_09_in16 = imem01_in[127:124];
    8: op1_09_in16 = reg_0548;
    9: op1_09_in16 = reg_0434;
    10: op1_09_in16 = reg_0254;
    11: op1_09_in16 = reg_0218;
    12: op1_09_in16 = imem05_in[71:68];
    13: op1_09_in16 = reg_0359;
    14: op1_09_in16 = reg_0360;
    15: op1_09_in16 = reg_0835;
    75: op1_09_in16 = reg_0835;
    16: op1_09_in16 = reg_0194;
    20: op1_09_in16 = reg_0194;
    17: op1_09_in16 = reg_0346;
    18: op1_09_in16 = reg_0196;
    53: op1_09_in16 = reg_0196;
    19: op1_09_in16 = imem02_in[115:112];
    21: op1_09_in16 = reg_0597;
    33: op1_09_in16 = reg_0597;
    22: op1_09_in16 = reg_0443;
    23: op1_09_in16 = reg_0725;
    24: op1_09_in16 = imem07_in[79:76];
    25: op1_09_in16 = reg_0188;
    26: op1_09_in16 = reg_0015;
    27: op1_09_in16 = reg_0510;
    28: op1_09_in16 = reg_0817;
    29: op1_09_in16 = reg_0463;
    30: op1_09_in16 = imem01_in[47:44];
    31: op1_09_in16 = reg_0502;
    32: op1_09_in16 = reg_0955;
    34: op1_09_in16 = imem01_in[51:48];
    35: op1_09_in16 = imem05_in[31:28];
    36: op1_09_in16 = imem05_in[87:84];
    37: op1_09_in16 = reg_0897;
    38: op1_09_in16 = reg_0074;
    39: op1_09_in16 = reg_0703;
    40: op1_09_in16 = reg_0735;
    41: op1_09_in16 = reg_0190;
    42: op1_09_in16 = imem05_in[63:60];
    43: op1_09_in16 = reg_0139;
    45: op1_09_in16 = imem03_in[27:24];
    46: op1_09_in16 = reg_0752;
    47: op1_09_in16 = reg_0744;
    48: op1_09_in16 = reg_0310;
    49: op1_09_in16 = reg_0066;
    50: op1_09_in16 = imem02_in[3:0];
    51: op1_09_in16 = reg_0456;
    54: op1_09_in16 = reg_0454;
    55: op1_09_in16 = imem03_in[119:116];
    56: op1_09_in16 = reg_0580;
    57: op1_09_in16 = imem04_in[23:20];
    58: op1_09_in16 = imem05_in[3:0];
    59: op1_09_in16 = imem05_in[59:56];
    60: op1_09_in16 = reg_0153;
    61: op1_09_in16 = reg_0660;
    62: op1_09_in16 = reg_0185;
    63: op1_09_in16 = imem02_in[91:88];
    64: op1_09_in16 = reg_0441;
    65: op1_09_in16 = reg_0976;
    66: op1_09_in16 = reg_0507;
    67: op1_09_in16 = reg_1004;
    68: op1_09_in16 = imem07_in[23:20];
    69: op1_09_in16 = reg_0646;
    92: op1_09_in16 = reg_0646;
    70: op1_09_in16 = reg_0071;
    71: op1_09_in16 = reg_0025;
    72: op1_09_in16 = imem02_in[79:76];
    73: op1_09_in16 = imem05_in[123:120];
    74: op1_09_in16 = reg_0067;
    77: op1_09_in16 = reg_1035;
    78: op1_09_in16 = imem01_in[99:96];
    79: op1_09_in16 = reg_0833;
    80: op1_09_in16 = imem05_in[115:112];
    81: op1_09_in16 = imem06_in[71:68];
    82: op1_09_in16 = reg_0568;
    83: op1_09_in16 = reg_0082;
    84: op1_09_in16 = reg_0174;
    85: op1_09_in16 = reg_0882;
    86: op1_09_in16 = reg_0393;
    87: op1_09_in16 = reg_0204;
    88: op1_09_in16 = reg_0661;
    89: op1_09_in16 = reg_1014;
    90: op1_09_in16 = reg_0385;
    91: op1_09_in16 = reg_0672;
    93: op1_09_in16 = reg_0428;
    94: op1_09_in16 = imem07_in[43:40];
    95: op1_09_in16 = imem07_in[83:80];
    96: op1_09_in16 = reg_0480;
    97: op1_09_in16 = reg_0822;
    default: op1_09_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_09_inv16 = 1;
    10: op1_09_inv16 = 1;
    11: op1_09_inv16 = 1;
    12: op1_09_inv16 = 1;
    13: op1_09_inv16 = 1;
    16: op1_09_inv16 = 1;
    21: op1_09_inv16 = 1;
    23: op1_09_inv16 = 1;
    25: op1_09_inv16 = 1;
    26: op1_09_inv16 = 1;
    29: op1_09_inv16 = 1;
    31: op1_09_inv16 = 1;
    33: op1_09_inv16 = 1;
    35: op1_09_inv16 = 1;
    36: op1_09_inv16 = 1;
    37: op1_09_inv16 = 1;
    39: op1_09_inv16 = 1;
    40: op1_09_inv16 = 1;
    41: op1_09_inv16 = 1;
    53: op1_09_inv16 = 1;
    54: op1_09_inv16 = 1;
    55: op1_09_inv16 = 1;
    58: op1_09_inv16 = 1;
    60: op1_09_inv16 = 1;
    61: op1_09_inv16 = 1;
    62: op1_09_inv16 = 1;
    64: op1_09_inv16 = 1;
    68: op1_09_inv16 = 1;
    70: op1_09_inv16 = 1;
    71: op1_09_inv16 = 1;
    73: op1_09_inv16 = 1;
    74: op1_09_inv16 = 1;
    75: op1_09_inv16 = 1;
    79: op1_09_inv16 = 1;
    80: op1_09_inv16 = 1;
    81: op1_09_inv16 = 1;
    83: op1_09_inv16 = 1;
    84: op1_09_inv16 = 1;
    86: op1_09_inv16 = 1;
    91: op1_09_inv16 = 1;
    92: op1_09_inv16 = 1;
    96: op1_09_inv16 = 1;
    default: op1_09_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の17番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in17 = reg_0379;
    7: op1_09_in17 = reg_0509;
    8: op1_09_in17 = reg_0537;
    9: op1_09_in17 = reg_0444;
    10: op1_09_in17 = reg_0255;
    73: op1_09_in17 = reg_0255;
    11: op1_09_in17 = reg_0224;
    12: op1_09_in17 = imem05_in[79:76];
    13: op1_09_in17 = reg_0355;
    14: op1_09_in17 = reg_0343;
    15: op1_09_in17 = reg_0251;
    70: op1_09_in17 = reg_0251;
    16: op1_09_in17 = reg_0198;
    17: op1_09_in17 = reg_0097;
    18: op1_09_in17 = reg_0202;
    19: op1_09_in17 = reg_0650;
    20: op1_09_in17 = imem01_in[27:24];
    21: op1_09_in17 = reg_0588;
    37: op1_09_in17 = reg_0588;
    22: op1_09_in17 = reg_0172;
    23: op1_09_in17 = reg_0707;
    24: op1_09_in17 = imem07_in[111:108];
    25: op1_09_in17 = reg_0205;
    26: op1_09_in17 = reg_0854;
    27: op1_09_in17 = reg_1032;
    28: op1_09_in17 = reg_0037;
    29: op1_09_in17 = reg_0450;
    30: op1_09_in17 = imem01_in[75:72];
    31: op1_09_in17 = reg_0561;
    32: op1_09_in17 = reg_0967;
    33: op1_09_in17 = imem07_in[23:20];
    34: op1_09_in17 = imem01_in[67:64];
    35: op1_09_in17 = imem05_in[87:84];
    36: op1_09_in17 = imem05_in[95:92];
    38: op1_09_in17 = reg_0072;
    39: op1_09_in17 = reg_0709;
    40: op1_09_in17 = reg_0870;
    41: op1_09_in17 = reg_0849;
    42: op1_09_in17 = imem05_in[115:112];
    43: op1_09_in17 = imem06_in[15:12];
    45: op1_09_in17 = imem03_in[67:64];
    46: op1_09_in17 = reg_0524;
    47: op1_09_in17 = reg_0419;
    48: op1_09_in17 = reg_0077;
    49: op1_09_in17 = reg_0014;
    82: op1_09_in17 = reg_0014;
    50: op1_09_in17 = imem02_in[23:20];
    51: op1_09_in17 = reg_0209;
    53: op1_09_in17 = reg_0212;
    54: op1_09_in17 = reg_0451;
    55: op1_09_in17 = imem03_in[123:120];
    56: op1_09_in17 = reg_0662;
    57: op1_09_in17 = imem04_in[75:72];
    58: op1_09_in17 = imem05_in[27:24];
    59: op1_09_in17 = imem05_in[91:88];
    60: op1_09_in17 = reg_0134;
    61: op1_09_in17 = reg_0625;
    62: op1_09_in17 = reg_0157;
    63: op1_09_in17 = imem02_in[115:112];
    64: op1_09_in17 = reg_0372;
    65: op1_09_in17 = imem04_in[7:4];
    66: op1_09_in17 = reg_0848;
    67: op1_09_in17 = reg_0937;
    68: op1_09_in17 = imem07_in[71:68];
    69: op1_09_in17 = reg_0544;
    71: op1_09_in17 = reg_0817;
    72: op1_09_in17 = imem02_in[99:96];
    74: op1_09_in17 = reg_0056;
    75: op1_09_in17 = reg_1010;
    77: op1_09_in17 = reg_0488;
    78: op1_09_in17 = reg_0122;
    79: op1_09_in17 = reg_0763;
    80: op1_09_in17 = reg_0215;
    81: op1_09_in17 = imem06_in[83:80];
    83: op1_09_in17 = reg_0886;
    84: op1_09_in17 = reg_0175;
    85: op1_09_in17 = reg_0123;
    86: op1_09_in17 = reg_0926;
    87: op1_09_in17 = reg_0186;
    88: op1_09_in17 = imem03_in[7:4];
    89: op1_09_in17 = reg_0971;
    90: op1_09_in17 = imem03_in[51:48];
    91: op1_09_in17 = reg_0820;
    92: op1_09_in17 = reg_0695;
    93: op1_09_in17 = reg_0599;
    94: op1_09_in17 = imem07_in[47:44];
    95: op1_09_in17 = reg_0710;
    96: op1_09_in17 = reg_0473;
    97: op1_09_in17 = reg_0370;
    default: op1_09_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv17 = 1;
    8: op1_09_inv17 = 1;
    9: op1_09_inv17 = 1;
    12: op1_09_inv17 = 1;
    13: op1_09_inv17 = 1;
    15: op1_09_inv17 = 1;
    16: op1_09_inv17 = 1;
    17: op1_09_inv17 = 1;
    18: op1_09_inv17 = 1;
    19: op1_09_inv17 = 1;
    20: op1_09_inv17 = 1;
    21: op1_09_inv17 = 1;
    23: op1_09_inv17 = 1;
    24: op1_09_inv17 = 1;
    25: op1_09_inv17 = 1;
    26: op1_09_inv17 = 1;
    27: op1_09_inv17 = 1;
    28: op1_09_inv17 = 1;
    29: op1_09_inv17 = 1;
    35: op1_09_inv17 = 1;
    36: op1_09_inv17 = 1;
    38: op1_09_inv17 = 1;
    41: op1_09_inv17 = 1;
    43: op1_09_inv17 = 1;
    46: op1_09_inv17 = 1;
    47: op1_09_inv17 = 1;
    48: op1_09_inv17 = 1;
    50: op1_09_inv17 = 1;
    53: op1_09_inv17 = 1;
    55: op1_09_inv17 = 1;
    56: op1_09_inv17 = 1;
    57: op1_09_inv17 = 1;
    58: op1_09_inv17 = 1;
    60: op1_09_inv17 = 1;
    62: op1_09_inv17 = 1;
    66: op1_09_inv17 = 1;
    68: op1_09_inv17 = 1;
    71: op1_09_inv17 = 1;
    72: op1_09_inv17 = 1;
    73: op1_09_inv17 = 1;
    77: op1_09_inv17 = 1;
    78: op1_09_inv17 = 1;
    79: op1_09_inv17 = 1;
    82: op1_09_inv17 = 1;
    88: op1_09_inv17 = 1;
    90: op1_09_inv17 = 1;
    93: op1_09_inv17 = 1;
    94: op1_09_inv17 = 1;
    96: op1_09_inv17 = 1;
    97: op1_09_inv17 = 1;
    default: op1_09_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の18番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in18 = reg_0381;
    7: op1_09_in18 = reg_0503;
    8: op1_09_in18 = reg_0555;
    9: op1_09_in18 = reg_0442;
    10: op1_09_in18 = reg_0142;
    11: op1_09_in18 = reg_0737;
    12: op1_09_in18 = imem05_in[87:84];
    13: op1_09_in18 = reg_0350;
    14: op1_09_in18 = reg_0396;
    15: op1_09_in18 = reg_0898;
    16: op1_09_in18 = imem01_in[7:4];
    17: op1_09_in18 = reg_0082;
    18: op1_09_in18 = imem01_in[67:64];
    19: op1_09_in18 = reg_0658;
    20: op1_09_in18 = imem01_in[47:44];
    21: op1_09_in18 = reg_0388;
    22: op1_09_in18 = reg_0179;
    23: op1_09_in18 = reg_0426;
    24: op1_09_in18 = reg_0720;
    25: op1_09_in18 = reg_0199;
    26: op1_09_in18 = reg_0856;
    27: op1_09_in18 = reg_0869;
    28: op1_09_in18 = reg_0091;
    29: op1_09_in18 = reg_0464;
    30: op1_09_in18 = imem01_in[87:84];
    31: op1_09_in18 = reg_0515;
    32: op1_09_in18 = reg_0954;
    33: op1_09_in18 = imem07_in[39:36];
    34: op1_09_in18 = imem01_in[79:76];
    35: op1_09_in18 = imem05_in[99:96];
    36: op1_09_in18 = reg_0966;
    37: op1_09_in18 = reg_0385;
    38: op1_09_in18 = reg_0882;
    39: op1_09_in18 = reg_0701;
    40: op1_09_in18 = reg_0560;
    41: op1_09_in18 = reg_1056;
    89: op1_09_in18 = reg_1056;
    42: op1_09_in18 = reg_0958;
    43: op1_09_in18 = imem06_in[19:16];
    45: op1_09_in18 = imem03_in[79:76];
    46: op1_09_in18 = reg_0076;
    47: op1_09_in18 = reg_0532;
    48: op1_09_in18 = reg_0884;
    49: op1_09_in18 = reg_0276;
    50: op1_09_in18 = imem02_in[95:92];
    51: op1_09_in18 = reg_0188;
    53: op1_09_in18 = reg_0197;
    54: op1_09_in18 = reg_0469;
    55: op1_09_in18 = imem03_in[127:124];
    56: op1_09_in18 = reg_0576;
    57: op1_09_in18 = imem04_in[79:76];
    58: op1_09_in18 = imem05_in[47:44];
    59: op1_09_in18 = imem05_in[111:108];
    60: op1_09_in18 = reg_0144;
    61: op1_09_in18 = reg_0926;
    63: op1_09_in18 = imem02_in[127:124];
    64: op1_09_in18 = reg_0347;
    65: op1_09_in18 = imem04_in[43:40];
    66: op1_09_in18 = reg_0752;
    67: op1_09_in18 = reg_0055;
    68: op1_09_in18 = imem07_in[87:84];
    69: op1_09_in18 = reg_0360;
    70: op1_09_in18 = reg_0332;
    71: op1_09_in18 = reg_0392;
    72: op1_09_in18 = reg_0739;
    73: op1_09_in18 = reg_0940;
    74: op1_09_in18 = reg_0401;
    75: op1_09_in18 = reg_0403;
    77: op1_09_in18 = reg_1022;
    78: op1_09_in18 = reg_1032;
    79: op1_09_in18 = reg_0762;
    80: op1_09_in18 = reg_0826;
    81: op1_09_in18 = imem06_in[87:84];
    82: op1_09_in18 = reg_0809;
    83: op1_09_in18 = reg_0279;
    84: op1_09_in18 = reg_0731;
    85: op1_09_in18 = reg_0848;
    86: op1_09_in18 = reg_0229;
    87: op1_09_in18 = reg_0198;
    88: op1_09_in18 = reg_0278;
    90: op1_09_in18 = imem03_in[59:56];
    91: op1_09_in18 = reg_0581;
    92: op1_09_in18 = reg_0956;
    93: op1_09_in18 = reg_0868;
    94: op1_09_in18 = imem07_in[51:48];
    95: op1_09_in18 = reg_0923;
    96: op1_09_in18 = reg_0470;
    97: op1_09_in18 = reg_0628;
    default: op1_09_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_09_inv18 = 1;
    9: op1_09_inv18 = 1;
    13: op1_09_inv18 = 1;
    14: op1_09_inv18 = 1;
    17: op1_09_inv18 = 1;
    18: op1_09_inv18 = 1;
    24: op1_09_inv18 = 1;
    25: op1_09_inv18 = 1;
    27: op1_09_inv18 = 1;
    28: op1_09_inv18 = 1;
    29: op1_09_inv18 = 1;
    30: op1_09_inv18 = 1;
    31: op1_09_inv18 = 1;
    32: op1_09_inv18 = 1;
    36: op1_09_inv18 = 1;
    37: op1_09_inv18 = 1;
    38: op1_09_inv18 = 1;
    39: op1_09_inv18 = 1;
    40: op1_09_inv18 = 1;
    43: op1_09_inv18 = 1;
    45: op1_09_inv18 = 1;
    48: op1_09_inv18 = 1;
    49: op1_09_inv18 = 1;
    53: op1_09_inv18 = 1;
    54: op1_09_inv18 = 1;
    55: op1_09_inv18 = 1;
    57: op1_09_inv18 = 1;
    58: op1_09_inv18 = 1;
    59: op1_09_inv18 = 1;
    60: op1_09_inv18 = 1;
    61: op1_09_inv18 = 1;
    64: op1_09_inv18 = 1;
    65: op1_09_inv18 = 1;
    67: op1_09_inv18 = 1;
    70: op1_09_inv18 = 1;
    72: op1_09_inv18 = 1;
    73: op1_09_inv18 = 1;
    74: op1_09_inv18 = 1;
    78: op1_09_inv18 = 1;
    81: op1_09_inv18 = 1;
    84: op1_09_inv18 = 1;
    86: op1_09_inv18 = 1;
    88: op1_09_inv18 = 1;
    91: op1_09_inv18 = 1;
    93: op1_09_inv18 = 1;
    96: op1_09_inv18 = 1;
    97: op1_09_inv18 = 1;
    default: op1_09_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の19番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in19 = reg_0392;
    7: op1_09_in19 = reg_0506;
    8: op1_09_in19 = reg_0540;
    9: op1_09_in19 = reg_0443;
    10: op1_09_in19 = reg_0143;
    11: op1_09_in19 = reg_0740;
    12: op1_09_in19 = imem05_in[107:104];
    13: op1_09_in19 = reg_0347;
    72: op1_09_in19 = reg_0347;
    14: op1_09_in19 = reg_0985;
    15: op1_09_in19 = reg_0254;
    16: op1_09_in19 = imem01_in[11:8];
    17: op1_09_in19 = reg_0084;
    18: op1_09_in19 = imem01_in[71:68];
    20: op1_09_in19 = imem01_in[71:68];
    19: op1_09_in19 = reg_0653;
    21: op1_09_in19 = reg_0369;
    22: op1_09_in19 = reg_0161;
    23: op1_09_in19 = reg_0419;
    24: op1_09_in19 = reg_0710;
    25: op1_09_in19 = reg_0197;
    26: op1_09_in19 = reg_0044;
    70: op1_09_in19 = reg_0044;
    27: op1_09_in19 = reg_0105;
    28: op1_09_in19 = reg_0049;
    29: op1_09_in19 = reg_0480;
    30: op1_09_in19 = imem01_in[91:88];
    31: op1_09_in19 = reg_0503;
    32: op1_09_in19 = reg_0961;
    33: op1_09_in19 = imem07_in[75:72];
    34: op1_09_in19 = reg_0860;
    35: op1_09_in19 = imem05_in[123:120];
    36: op1_09_in19 = reg_0954;
    37: op1_09_in19 = reg_0294;
    38: op1_09_in19 = reg_0278;
    39: op1_09_in19 = reg_0727;
    40: op1_09_in19 = reg_0003;
    41: op1_09_in19 = reg_0250;
    42: op1_09_in19 = reg_0971;
    78: op1_09_in19 = reg_0971;
    43: op1_09_in19 = imem06_in[39:36];
    45: op1_09_in19 = imem03_in[91:88];
    46: op1_09_in19 = reg_0067;
    47: op1_09_in19 = reg_0427;
    48: op1_09_in19 = imem03_in[19:16];
    49: op1_09_in19 = reg_0284;
    66: op1_09_in19 = reg_0284;
    50: op1_09_in19 = imem02_in[123:120];
    51: op1_09_in19 = reg_0193;
    53: op1_09_in19 = reg_0560;
    54: op1_09_in19 = reg_0472;
    55: op1_09_in19 = reg_0823;
    56: op1_09_in19 = reg_0795;
    57: op1_09_in19 = imem04_in[91:88];
    58: op1_09_in19 = imem05_in[67:64];
    59: op1_09_in19 = reg_0944;
    60: op1_09_in19 = imem06_in[7:4];
    61: op1_09_in19 = reg_1030;
    63: op1_09_in19 = reg_0323;
    64: op1_09_in19 = reg_0482;
    65: op1_09_in19 = imem04_in[51:48];
    67: op1_09_in19 = reg_1020;
    68: op1_09_in19 = imem07_in[107:104];
    69: op1_09_in19 = reg_1052;
    71: op1_09_in19 = reg_0617;
    73: op1_09_in19 = reg_0020;
    74: op1_09_in19 = reg_0815;
    75: op1_09_in19 = reg_0567;
    77: op1_09_in19 = reg_0518;
    79: op1_09_in19 = reg_0837;
    80: op1_09_in19 = reg_0492;
    81: op1_09_in19 = imem06_in[107:104];
    82: op1_09_in19 = reg_0732;
    83: op1_09_in19 = reg_0441;
    84: op1_09_in19 = reg_0339;
    85: op1_09_in19 = reg_0058;
    86: op1_09_in19 = reg_0889;
    87: op1_09_in19 = reg_0212;
    88: op1_09_in19 = reg_0756;
    89: op1_09_in19 = reg_0488;
    90: op1_09_in19 = imem03_in[75:72];
    91: op1_09_in19 = reg_0445;
    92: op1_09_in19 = reg_0129;
    93: op1_09_in19 = reg_0024;
    94: op1_09_in19 = imem07_in[111:108];
    95: op1_09_in19 = reg_0442;
    96: op1_09_in19 = reg_0471;
    97: op1_09_in19 = reg_0804;
    default: op1_09_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv19 = 1;
    10: op1_09_inv19 = 1;
    11: op1_09_inv19 = 1;
    12: op1_09_inv19 = 1;
    13: op1_09_inv19 = 1;
    14: op1_09_inv19 = 1;
    15: op1_09_inv19 = 1;
    19: op1_09_inv19 = 1;
    21: op1_09_inv19 = 1;
    22: op1_09_inv19 = 1;
    26: op1_09_inv19 = 1;
    27: op1_09_inv19 = 1;
    28: op1_09_inv19 = 1;
    29: op1_09_inv19 = 1;
    30: op1_09_inv19 = 1;
    31: op1_09_inv19 = 1;
    32: op1_09_inv19 = 1;
    33: op1_09_inv19 = 1;
    35: op1_09_inv19 = 1;
    36: op1_09_inv19 = 1;
    39: op1_09_inv19 = 1;
    40: op1_09_inv19 = 1;
    41: op1_09_inv19 = 1;
    42: op1_09_inv19 = 1;
    45: op1_09_inv19 = 1;
    46: op1_09_inv19 = 1;
    47: op1_09_inv19 = 1;
    49: op1_09_inv19 = 1;
    54: op1_09_inv19 = 1;
    56: op1_09_inv19 = 1;
    59: op1_09_inv19 = 1;
    60: op1_09_inv19 = 1;
    61: op1_09_inv19 = 1;
    63: op1_09_inv19 = 1;
    64: op1_09_inv19 = 1;
    70: op1_09_inv19 = 1;
    72: op1_09_inv19 = 1;
    77: op1_09_inv19 = 1;
    78: op1_09_inv19 = 1;
    79: op1_09_inv19 = 1;
    80: op1_09_inv19 = 1;
    81: op1_09_inv19 = 1;
    86: op1_09_inv19 = 1;
    87: op1_09_inv19 = 1;
    88: op1_09_inv19 = 1;
    93: op1_09_inv19 = 1;
    95: op1_09_inv19 = 1;
    default: op1_09_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の20番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in20 = reg_0371;
    7: op1_09_in20 = reg_0233;
    8: op1_09_in20 = reg_0532;
    25: op1_09_in20 = reg_0532;
    9: op1_09_in20 = reg_0435;
    10: op1_09_in20 = reg_0134;
    11: op1_09_in20 = reg_0793;
    12: op1_09_in20 = reg_0147;
    13: op1_09_in20 = reg_0083;
    14: op1_09_in20 = reg_0980;
    15: op1_09_in20 = reg_0255;
    16: op1_09_in20 = imem01_in[39:36];
    17: op1_09_in20 = reg_0079;
    18: op1_09_in20 = imem01_in[87:84];
    19: op1_09_in20 = reg_0637;
    20: op1_09_in20 = imem01_in[107:104];
    21: op1_09_in20 = reg_0377;
    22: op1_09_in20 = reg_0182;
    23: op1_09_in20 = reg_0439;
    24: op1_09_in20 = reg_0706;
    26: op1_09_in20 = imem05_in[59:56];
    27: op1_09_in20 = reg_0107;
    28: op1_09_in20 = reg_0016;
    29: op1_09_in20 = reg_0470;
    30: op1_09_in20 = imem01_in[111:108];
    31: op1_09_in20 = imem03_in[3:0];
    64: op1_09_in20 = imem03_in[3:0];
    32: op1_09_in20 = reg_0022;
    33: op1_09_in20 = imem07_in[87:84];
    34: op1_09_in20 = reg_0544;
    35: op1_09_in20 = reg_0959;
    36: op1_09_in20 = reg_0949;
    37: op1_09_in20 = reg_0383;
    38: op1_09_in20 = reg_0777;
    39: op1_09_in20 = reg_0441;
    40: op1_09_in20 = reg_0299;
    41: op1_09_in20 = reg_0013;
    42: op1_09_in20 = reg_0955;
    43: op1_09_in20 = imem06_in[43:40];
    45: op1_09_in20 = imem03_in[123:120];
    46: op1_09_in20 = reg_0584;
    47: op1_09_in20 = reg_0175;
    48: op1_09_in20 = imem03_in[67:64];
    49: op1_09_in20 = imem04_in[3:0];
    50: op1_09_in20 = reg_0656;
    51: op1_09_in20 = reg_0207;
    53: op1_09_in20 = reg_0099;
    54: op1_09_in20 = reg_0480;
    55: op1_09_in20 = reg_0874;
    56: op1_09_in20 = reg_0246;
    57: op1_09_in20 = imem04_in[111:108];
    58: op1_09_in20 = imem05_in[83:80];
    59: op1_09_in20 = reg_0675;
    60: op1_09_in20 = imem06_in[31:28];
    61: op1_09_in20 = reg_0011;
    63: op1_09_in20 = reg_0358;
    79: op1_09_in20 = reg_0358;
    65: op1_09_in20 = imem04_in[55:52];
    66: op1_09_in20 = reg_0764;
    82: op1_09_in20 = reg_0764;
    67: op1_09_in20 = reg_0292;
    68: op1_09_in20 = reg_0719;
    69: op1_09_in20 = imem01_in[15:12];
    70: op1_09_in20 = imem05_in[7:4];
    71: op1_09_in20 = reg_0863;
    72: op1_09_in20 = reg_0089;
    73: op1_09_in20 = reg_0688;
    74: op1_09_in20 = reg_0809;
    75: op1_09_in20 = reg_0704;
    77: op1_09_in20 = reg_0234;
    78: op1_09_in20 = reg_1024;
    80: op1_09_in20 = reg_0235;
    81: op1_09_in20 = imem06_in[115:112];
    83: op1_09_in20 = reg_0039;
    84: op1_09_in20 = reg_0183;
    85: op1_09_in20 = reg_0401;
    86: op1_09_in20 = reg_0384;
    87: op1_09_in20 = imem01_in[47:44];
    88: op1_09_in20 = reg_0551;
    89: op1_09_in20 = reg_1022;
    90: op1_09_in20 = imem03_in[99:96];
    91: op1_09_in20 = reg_0978;
    92: op1_09_in20 = reg_0437;
    93: op1_09_in20 = reg_0429;
    94: op1_09_in20 = imem07_in[119:116];
    95: op1_09_in20 = reg_0759;
    96: op1_09_in20 = reg_0208;
    97: op1_09_in20 = imem07_in[43:40];
    default: op1_09_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv20 = 1;
    9: op1_09_inv20 = 1;
    12: op1_09_inv20 = 1;
    13: op1_09_inv20 = 1;
    14: op1_09_inv20 = 1;
    15: op1_09_inv20 = 1;
    16: op1_09_inv20 = 1;
    17: op1_09_inv20 = 1;
    19: op1_09_inv20 = 1;
    20: op1_09_inv20 = 1;
    21: op1_09_inv20 = 1;
    25: op1_09_inv20 = 1;
    27: op1_09_inv20 = 1;
    29: op1_09_inv20 = 1;
    34: op1_09_inv20 = 1;
    36: op1_09_inv20 = 1;
    39: op1_09_inv20 = 1;
    46: op1_09_inv20 = 1;
    49: op1_09_inv20 = 1;
    50: op1_09_inv20 = 1;
    51: op1_09_inv20 = 1;
    53: op1_09_inv20 = 1;
    57: op1_09_inv20 = 1;
    58: op1_09_inv20 = 1;
    63: op1_09_inv20 = 1;
    64: op1_09_inv20 = 1;
    65: op1_09_inv20 = 1;
    66: op1_09_inv20 = 1;
    67: op1_09_inv20 = 1;
    70: op1_09_inv20 = 1;
    72: op1_09_inv20 = 1;
    73: op1_09_inv20 = 1;
    78: op1_09_inv20 = 1;
    82: op1_09_inv20 = 1;
    83: op1_09_inv20 = 1;
    84: op1_09_inv20 = 1;
    86: op1_09_inv20 = 1;
    87: op1_09_inv20 = 1;
    90: op1_09_inv20 = 1;
    93: op1_09_inv20 = 1;
    94: op1_09_inv20 = 1;
    95: op1_09_inv20 = 1;
    default: op1_09_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の21番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in21 = reg_0390;
    7: op1_09_in21 = reg_0218;
    8: op1_09_in21 = reg_0301;
    57: op1_09_in21 = reg_0301;
    9: op1_09_in21 = reg_0181;
    93: op1_09_in21 = reg_0181;
    10: op1_09_in21 = imem06_in[7:4];
    11: op1_09_in21 = reg_0221;
    12: op1_09_in21 = reg_0151;
    13: op1_09_in21 = reg_0092;
    14: op1_09_in21 = imem04_in[95:92];
    15: op1_09_in21 = reg_0253;
    16: op1_09_in21 = imem01_in[47:44];
    69: op1_09_in21 = imem01_in[47:44];
    17: op1_09_in21 = imem03_in[39:36];
    18: op1_09_in21 = imem01_in[95:92];
    19: op1_09_in21 = reg_0648;
    20: op1_09_in21 = reg_0013;
    21: op1_09_in21 = reg_0984;
    22: op1_09_in21 = reg_0163;
    23: op1_09_in21 = reg_0428;
    24: op1_09_in21 = reg_0429;
    25: op1_09_in21 = reg_0926;
    26: op1_09_in21 = reg_0967;
    27: op1_09_in21 = reg_0113;
    28: op1_09_in21 = reg_0872;
    29: op1_09_in21 = reg_0459;
    30: op1_09_in21 = reg_0779;
    31: op1_09_in21 = imem03_in[47:44];
    32: op1_09_in21 = reg_0835;
    33: op1_09_in21 = imem07_in[111:108];
    34: op1_09_in21 = reg_0087;
    35: op1_09_in21 = reg_0948;
    36: op1_09_in21 = reg_0947;
    37: op1_09_in21 = reg_0399;
    38: op1_09_in21 = imem05_in[11:8];
    39: op1_09_in21 = reg_0445;
    40: op1_09_in21 = reg_0240;
    41: op1_09_in21 = reg_0299;
    42: op1_09_in21 = reg_0957;
    43: op1_09_in21 = imem06_in[67:64];
    45: op1_09_in21 = reg_1050;
    46: op1_09_in21 = reg_0815;
    85: op1_09_in21 = reg_0815;
    47: op1_09_in21 = reg_0179;
    48: op1_09_in21 = imem03_in[87:84];
    49: op1_09_in21 = imem04_in[11:8];
    50: op1_09_in21 = reg_0082;
    51: op1_09_in21 = reg_0196;
    53: op1_09_in21 = reg_0107;
    54: op1_09_in21 = reg_0471;
    55: op1_09_in21 = reg_0833;
    56: op1_09_in21 = reg_0998;
    58: op1_09_in21 = imem05_in[103:100];
    59: op1_09_in21 = reg_0955;
    60: op1_09_in21 = imem06_in[59:56];
    61: op1_09_in21 = imem06_in[3:0];
    63: op1_09_in21 = reg_0248;
    64: op1_09_in21 = imem03_in[19:16];
    65: op1_09_in21 = imem04_in[87:84];
    66: op1_09_in21 = reg_0432;
    67: op1_09_in21 = reg_0540;
    68: op1_09_in21 = reg_0726;
    70: op1_09_in21 = imem05_in[91:88];
    71: op1_09_in21 = imem06_in[19:16];
    72: op1_09_in21 = reg_0086;
    73: op1_09_in21 = reg_0125;
    74: op1_09_in21 = reg_0764;
    75: op1_09_in21 = reg_0308;
    77: op1_09_in21 = reg_0225;
    78: op1_09_in21 = reg_0522;
    79: op1_09_in21 = reg_0441;
    80: op1_09_in21 = reg_0137;
    81: op1_09_in21 = reg_0010;
    82: op1_09_in21 = reg_0494;
    83: op1_09_in21 = reg_0664;
    84: op1_09_in21 = reg_0565;
    86: op1_09_in21 = imem06_in[23:20];
    87: op1_09_in21 = imem01_in[91:88];
    88: op1_09_in21 = reg_0987;
    89: op1_09_in21 = reg_0234;
    90: op1_09_in21 = imem04_in[3:0];
    91: op1_09_in21 = reg_0396;
    92: op1_09_in21 = reg_0651;
    94: op1_09_in21 = reg_0567;
    95: op1_09_in21 = reg_0002;
    96: op1_09_in21 = reg_0204;
    97: op1_09_in21 = imem07_in[87:84];
    default: op1_09_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    11: op1_09_inv21 = 1;
    15: op1_09_inv21 = 1;
    17: op1_09_inv21 = 1;
    21: op1_09_inv21 = 1;
    22: op1_09_inv21 = 1;
    25: op1_09_inv21 = 1;
    26: op1_09_inv21 = 1;
    33: op1_09_inv21 = 1;
    35: op1_09_inv21 = 1;
    36: op1_09_inv21 = 1;
    39: op1_09_inv21 = 1;
    40: op1_09_inv21 = 1;
    41: op1_09_inv21 = 1;
    42: op1_09_inv21 = 1;
    45: op1_09_inv21 = 1;
    46: op1_09_inv21 = 1;
    47: op1_09_inv21 = 1;
    48: op1_09_inv21 = 1;
    50: op1_09_inv21 = 1;
    58: op1_09_inv21 = 1;
    59: op1_09_inv21 = 1;
    60: op1_09_inv21 = 1;
    61: op1_09_inv21 = 1;
    63: op1_09_inv21 = 1;
    66: op1_09_inv21 = 1;
    67: op1_09_inv21 = 1;
    68: op1_09_inv21 = 1;
    69: op1_09_inv21 = 1;
    70: op1_09_inv21 = 1;
    71: op1_09_inv21 = 1;
    73: op1_09_inv21 = 1;
    74: op1_09_inv21 = 1;
    78: op1_09_inv21 = 1;
    80: op1_09_inv21 = 1;
    81: op1_09_inv21 = 1;
    87: op1_09_inv21 = 1;
    89: op1_09_inv21 = 1;
    90: op1_09_inv21 = 1;
    91: op1_09_inv21 = 1;
    93: op1_09_inv21 = 1;
    95: op1_09_inv21 = 1;
    96: op1_09_inv21 = 1;
    97: op1_09_inv21 = 1;
    default: op1_09_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の22番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in22 = reg_0367;
    7: op1_09_in22 = reg_0245;
    8: op1_09_in22 = reg_0279;
    9: op1_09_in22 = reg_0162;
    10: op1_09_in22 = imem06_in[23:20];
    11: op1_09_in22 = reg_0812;
    12: op1_09_in22 = reg_0153;
    13: op1_09_in22 = reg_0049;
    14: op1_09_in22 = imem04_in[107:104];
    15: op1_09_in22 = reg_0148;
    16: op1_09_in22 = imem01_in[51:48];
    69: op1_09_in22 = imem01_in[51:48];
    17: op1_09_in22 = imem03_in[63:60];
    18: op1_09_in22 = imem01_in[99:96];
    19: op1_09_in22 = reg_0638;
    20: op1_09_in22 = reg_0762;
    21: op1_09_in22 = reg_0974;
    22: op1_09_in22 = reg_0178;
    23: op1_09_in22 = reg_0431;
    24: op1_09_in22 = reg_0418;
    25: op1_09_in22 = reg_0220;
    26: op1_09_in22 = reg_0956;
    27: op1_09_in22 = imem02_in[31:28];
    28: op1_09_in22 = reg_0012;
    29: op1_09_in22 = reg_0208;
    30: op1_09_in22 = reg_0510;
    31: op1_09_in22 = imem03_in[55:52];
    32: op1_09_in22 = reg_0900;
    33: op1_09_in22 = imem07_in[119:116];
    34: op1_09_in22 = reg_0221;
    35: op1_09_in22 = reg_0964;
    36: op1_09_in22 = reg_0943;
    37: op1_09_in22 = reg_0390;
    38: op1_09_in22 = imem05_in[15:12];
    39: op1_09_in22 = reg_0438;
    40: op1_09_in22 = reg_0544;
    41: op1_09_in22 = reg_0224;
    42: op1_09_in22 = reg_0948;
    43: op1_09_in22 = imem06_in[103:100];
    45: op1_09_in22 = reg_0317;
    46: op1_09_in22 = reg_0064;
    47: op1_09_in22 = reg_0168;
    48: op1_09_in22 = imem03_in[115:112];
    49: op1_09_in22 = imem04_in[27:24];
    50: op1_09_in22 = reg_0643;
    51: op1_09_in22 = imem01_in[27:24];
    53: op1_09_in22 = reg_0523;
    54: op1_09_in22 = reg_0209;
    55: op1_09_in22 = reg_0376;
    56: op1_09_in22 = reg_0982;
    57: op1_09_in22 = reg_0511;
    58: op1_09_in22 = imem05_in[107:104];
    70: op1_09_in22 = imem05_in[107:104];
    59: op1_09_in22 = reg_0022;
    60: op1_09_in22 = imem06_in[71:68];
    61: op1_09_in22 = imem06_in[19:16];
    63: op1_09_in22 = reg_0818;
    64: op1_09_in22 = imem03_in[39:36];
    65: op1_09_in22 = imem04_in[103:100];
    66: op1_09_in22 = reg_0243;
    67: op1_09_in22 = reg_0050;
    68: op1_09_in22 = reg_0727;
    71: op1_09_in22 = imem06_in[27:24];
    72: op1_09_in22 = reg_0506;
    73: op1_09_in22 = reg_0447;
    74: op1_09_in22 = reg_0494;
    75: op1_09_in22 = reg_0092;
    77: op1_09_in22 = reg_0500;
    78: op1_09_in22 = reg_0798;
    79: op1_09_in22 = reg_0389;
    80: op1_09_in22 = reg_0256;
    81: op1_09_in22 = reg_0244;
    82: op1_09_in22 = reg_0627;
    83: op1_09_in22 = reg_0248;
    84: op1_09_in22 = reg_0724;
    85: op1_09_in22 = reg_0072;
    86: op1_09_in22 = imem06_in[43:40];
    87: op1_09_in22 = reg_0973;
    88: op1_09_in22 = reg_0989;
    89: op1_09_in22 = reg_0962;
    90: op1_09_in22 = imem04_in[31:28];
    91: op1_09_in22 = imem04_in[3:0];
    92: op1_09_in22 = reg_0146;
    93: op1_09_in22 = reg_0183;
    94: op1_09_in22 = reg_0563;
    95: op1_09_in22 = reg_0433;
    96: op1_09_in22 = reg_0203;
    97: op1_09_in22 = imem07_in[99:96];
    default: op1_09_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv22 = 1;
    9: op1_09_inv22 = 1;
    11: op1_09_inv22 = 1;
    13: op1_09_inv22 = 1;
    16: op1_09_inv22 = 1;
    17: op1_09_inv22 = 1;
    19: op1_09_inv22 = 1;
    25: op1_09_inv22 = 1;
    27: op1_09_inv22 = 1;
    29: op1_09_inv22 = 1;
    31: op1_09_inv22 = 1;
    32: op1_09_inv22 = 1;
    34: op1_09_inv22 = 1;
    35: op1_09_inv22 = 1;
    36: op1_09_inv22 = 1;
    39: op1_09_inv22 = 1;
    40: op1_09_inv22 = 1;
    41: op1_09_inv22 = 1;
    42: op1_09_inv22 = 1;
    45: op1_09_inv22 = 1;
    48: op1_09_inv22 = 1;
    49: op1_09_inv22 = 1;
    56: op1_09_inv22 = 1;
    57: op1_09_inv22 = 1;
    59: op1_09_inv22 = 1;
    60: op1_09_inv22 = 1;
    61: op1_09_inv22 = 1;
    63: op1_09_inv22 = 1;
    64: op1_09_inv22 = 1;
    65: op1_09_inv22 = 1;
    67: op1_09_inv22 = 1;
    69: op1_09_inv22 = 1;
    70: op1_09_inv22 = 1;
    73: op1_09_inv22 = 1;
    85: op1_09_inv22 = 1;
    86: op1_09_inv22 = 1;
    87: op1_09_inv22 = 1;
    90: op1_09_inv22 = 1;
    92: op1_09_inv22 = 1;
    94: op1_09_inv22 = 1;
    97: op1_09_inv22 = 1;
    default: op1_09_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の23番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in23 = reg_0035;
    7: op1_09_in23 = reg_0219;
    8: op1_09_in23 = reg_0293;
    9: op1_09_in23 = reg_0182;
    10: op1_09_in23 = imem06_in[55:52];
    11: op1_09_in23 = reg_1042;
    12: op1_09_in23 = imem06_in[43:40];
    13: op1_09_in23 = reg_0087;
    14: op1_09_in23 = reg_0560;
    15: op1_09_in23 = reg_0128;
    16: op1_09_in23 = imem01_in[63:60];
    17: op1_09_in23 = imem03_in[79:76];
    18: op1_09_in23 = imem01_in[111:108];
    19: op1_09_in23 = reg_0659;
    20: op1_09_in23 = reg_0242;
    21: op1_09_in23 = reg_0990;
    22: op1_09_in23 = reg_0157;
    23: op1_09_in23 = reg_0165;
    24: op1_09_in23 = reg_0442;
    25: op1_09_in23 = imem01_in[35:32];
    26: op1_09_in23 = reg_0942;
    42: op1_09_in23 = reg_0942;
    27: op1_09_in23 = imem02_in[107:104];
    28: op1_09_in23 = reg_0360;
    29: op1_09_in23 = reg_0201;
    30: op1_09_in23 = reg_0299;
    75: op1_09_in23 = reg_0299;
    31: op1_09_in23 = imem03_in[99:96];
    32: op1_09_in23 = reg_0275;
    33: op1_09_in23 = imem07_in[123:120];
    34: op1_09_in23 = reg_1039;
    35: op1_09_in23 = reg_0951;
    36: op1_09_in23 = reg_0960;
    37: op1_09_in23 = reg_0380;
    38: op1_09_in23 = imem05_in[19:16];
    39: op1_09_in23 = reg_0175;
    40: op1_09_in23 = imem01_in[75:72];
    41: op1_09_in23 = reg_0810;
    43: op1_09_in23 = imem06_in[119:116];
    45: op1_09_in23 = reg_1019;
    46: op1_09_in23 = imem04_in[7:4];
    47: op1_09_in23 = reg_0170;
    48: op1_09_in23 = reg_0394;
    49: op1_09_in23 = imem04_in[67:64];
    50: op1_09_in23 = reg_0648;
    51: op1_09_in23 = imem01_in[79:76];
    53: op1_09_in23 = reg_1018;
    54: op1_09_in23 = reg_0196;
    55: op1_09_in23 = reg_0513;
    56: op1_09_in23 = reg_0977;
    57: op1_09_in23 = reg_0277;
    58: op1_09_in23 = reg_0255;
    59: op1_09_in23 = reg_0237;
    60: op1_09_in23 = imem06_in[83:80];
    61: op1_09_in23 = imem06_in[47:44];
    63: op1_09_in23 = reg_0608;
    64: op1_09_in23 = imem03_in[95:92];
    65: op1_09_in23 = reg_1006;
    66: op1_09_in23 = reg_0027;
    67: op1_09_in23 = reg_0537;
    68: op1_09_in23 = reg_0303;
    69: op1_09_in23 = imem01_in[95:92];
    70: op1_09_in23 = imem05_in[119:116];
    71: op1_09_in23 = imem06_in[31:28];
    72: op1_09_in23 = reg_0091;
    73: op1_09_in23 = reg_0156;
    74: op1_09_in23 = reg_0409;
    77: op1_09_in23 = reg_1037;
    78: op1_09_in23 = reg_0604;
    79: op1_09_in23 = reg_0037;
    80: op1_09_in23 = reg_0963;
    81: op1_09_in23 = reg_0262;
    82: op1_09_in23 = reg_0777;
    83: op1_09_in23 = reg_0818;
    85: op1_09_in23 = reg_0243;
    86: op1_09_in23 = imem06_in[95:92];
    87: op1_09_in23 = reg_0337;
    88: op1_09_in23 = imem04_in[15:12];
    89: op1_09_in23 = reg_0798;
    90: op1_09_in23 = imem04_in[43:40];
    91: op1_09_in23 = imem04_in[55:52];
    92: op1_09_in23 = reg_0949;
    93: op1_09_in23 = reg_0690;
    94: op1_09_in23 = reg_0420;
    95: op1_09_in23 = reg_0321;
    96: op1_09_in23 = reg_0205;
    97: op1_09_in23 = imem07_in[103:100];
    default: op1_09_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv23 = 1;
    8: op1_09_inv23 = 1;
    11: op1_09_inv23 = 1;
    12: op1_09_inv23 = 1;
    15: op1_09_inv23 = 1;
    16: op1_09_inv23 = 1;
    17: op1_09_inv23 = 1;
    18: op1_09_inv23 = 1;
    19: op1_09_inv23 = 1;
    20: op1_09_inv23 = 1;
    22: op1_09_inv23 = 1;
    23: op1_09_inv23 = 1;
    24: op1_09_inv23 = 1;
    27: op1_09_inv23 = 1;
    30: op1_09_inv23 = 1;
    31: op1_09_inv23 = 1;
    32: op1_09_inv23 = 1;
    33: op1_09_inv23 = 1;
    38: op1_09_inv23 = 1;
    39: op1_09_inv23 = 1;
    41: op1_09_inv23 = 1;
    43: op1_09_inv23 = 1;
    45: op1_09_inv23 = 1;
    46: op1_09_inv23 = 1;
    47: op1_09_inv23 = 1;
    50: op1_09_inv23 = 1;
    54: op1_09_inv23 = 1;
    56: op1_09_inv23 = 1;
    59: op1_09_inv23 = 1;
    61: op1_09_inv23 = 1;
    65: op1_09_inv23 = 1;
    66: op1_09_inv23 = 1;
    67: op1_09_inv23 = 1;
    68: op1_09_inv23 = 1;
    69: op1_09_inv23 = 1;
    72: op1_09_inv23 = 1;
    77: op1_09_inv23 = 1;
    79: op1_09_inv23 = 1;
    80: op1_09_inv23 = 1;
    82: op1_09_inv23 = 1;
    91: op1_09_inv23 = 1;
    96: op1_09_inv23 = 1;
    default: op1_09_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の24番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in24 = reg_0020;
    7: op1_09_in24 = reg_0118;
    8: op1_09_in24 = reg_0307;
    9: op1_09_in24 = reg_0183;
    10: op1_09_in24 = imem06_in[75:72];
    11: op1_09_in24 = reg_1032;
    12: op1_09_in24 = imem06_in[51:48];
    13: op1_09_in24 = reg_0073;
    14: op1_09_in24 = reg_0554;
    15: op1_09_in24 = reg_0139;
    16: op1_09_in24 = reg_0235;
    17: op1_09_in24 = reg_0602;
    18: op1_09_in24 = reg_0735;
    19: op1_09_in24 = reg_0329;
    20: op1_09_in24 = reg_0502;
    21: op1_09_in24 = imem04_in[23:20];
    23: op1_09_in24 = reg_0168;
    24: op1_09_in24 = reg_0165;
    25: op1_09_in24 = imem01_in[95:92];
    26: op1_09_in24 = reg_0949;
    27: op1_09_in24 = imem02_in[119:116];
    28: op1_09_in24 = reg_0302;
    29: op1_09_in24 = reg_0212;
    30: op1_09_in24 = reg_0224;
    31: op1_09_in24 = imem03_in[115:112];
    32: op1_09_in24 = reg_0896;
    33: op1_09_in24 = imem07_in[127:124];
    34: op1_09_in24 = reg_0226;
    35: op1_09_in24 = reg_0942;
    36: op1_09_in24 = reg_0215;
    37: op1_09_in24 = imem06_in[67:64];
    38: op1_09_in24 = imem05_in[27:24];
    39: op1_09_in24 = reg_0166;
    40: op1_09_in24 = imem01_in[83:80];
    41: op1_09_in24 = reg_0248;
    42: op1_09_in24 = reg_1021;
    43: op1_09_in24 = reg_0883;
    45: op1_09_in24 = reg_0397;
    46: op1_09_in24 = imem04_in[19:16];
    48: op1_09_in24 = reg_1007;
    49: op1_09_in24 = imem04_in[83:80];
    50: op1_09_in24 = reg_0045;
    51: op1_09_in24 = imem01_in[91:88];
    53: op1_09_in24 = reg_0905;
    54: op1_09_in24 = reg_0205;
    55: op1_09_in24 = reg_0246;
    56: op1_09_in24 = reg_0983;
    57: op1_09_in24 = reg_0912;
    58: op1_09_in24 = reg_0866;
    59: op1_09_in24 = reg_0497;
    60: op1_09_in24 = imem06_in[99:96];
    61: op1_09_in24 = imem06_in[91:88];
    63: op1_09_in24 = reg_0772;
    64: op1_09_in24 = reg_0345;
    65: op1_09_in24 = reg_0530;
    66: op1_09_in24 = reg_0627;
    67: op1_09_in24 = reg_0313;
    68: op1_09_in24 = reg_0325;
    69: op1_09_in24 = imem01_in[99:96];
    70: op1_09_in24 = reg_1015;
    71: op1_09_in24 = imem06_in[43:40];
    72: op1_09_in24 = reg_0077;
    73: op1_09_in24 = reg_0155;
    74: op1_09_in24 = reg_0495;
    75: op1_09_in24 = reg_0708;
    77: op1_09_in24 = reg_0906;
    78: op1_09_in24 = reg_1040;
    79: op1_09_in24 = reg_0347;
    83: op1_09_in24 = reg_0347;
    80: op1_09_in24 = reg_0525;
    81: op1_09_in24 = reg_0679;
    82: op1_09_in24 = reg_0542;
    85: op1_09_in24 = reg_0552;
    86: op1_09_in24 = imem06_in[127:124];
    87: op1_09_in24 = reg_0546;
    88: op1_09_in24 = imem04_in[47:44];
    89: op1_09_in24 = reg_0830;
    90: op1_09_in24 = imem04_in[79:76];
    91: op1_09_in24 = imem04_in[59:56];
    92: op1_09_in24 = reg_0965;
    94: op1_09_in24 = reg_0427;
    95: op1_09_in24 = reg_0406;
    96: op1_09_in24 = reg_0202;
    97: op1_09_in24 = reg_0162;
    default: op1_09_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv24 = 1;
    7: op1_09_inv24 = 1;
    8: op1_09_inv24 = 1;
    9: op1_09_inv24 = 1;
    10: op1_09_inv24 = 1;
    11: op1_09_inv24 = 1;
    12: op1_09_inv24 = 1;
    13: op1_09_inv24 = 1;
    14: op1_09_inv24 = 1;
    15: op1_09_inv24 = 1;
    17: op1_09_inv24 = 1;
    19: op1_09_inv24 = 1;
    20: op1_09_inv24 = 1;
    21: op1_09_inv24 = 1;
    23: op1_09_inv24 = 1;
    25: op1_09_inv24 = 1;
    26: op1_09_inv24 = 1;
    27: op1_09_inv24 = 1;
    28: op1_09_inv24 = 1;
    29: op1_09_inv24 = 1;
    30: op1_09_inv24 = 1;
    31: op1_09_inv24 = 1;
    33: op1_09_inv24 = 1;
    38: op1_09_inv24 = 1;
    39: op1_09_inv24 = 1;
    41: op1_09_inv24 = 1;
    42: op1_09_inv24 = 1;
    43: op1_09_inv24 = 1;
    48: op1_09_inv24 = 1;
    50: op1_09_inv24 = 1;
    51: op1_09_inv24 = 1;
    53: op1_09_inv24 = 1;
    54: op1_09_inv24 = 1;
    55: op1_09_inv24 = 1;
    56: op1_09_inv24 = 1;
    58: op1_09_inv24 = 1;
    60: op1_09_inv24 = 1;
    63: op1_09_inv24 = 1;
    66: op1_09_inv24 = 1;
    67: op1_09_inv24 = 1;
    68: op1_09_inv24 = 1;
    70: op1_09_inv24 = 1;
    73: op1_09_inv24 = 1;
    77: op1_09_inv24 = 1;
    78: op1_09_inv24 = 1;
    79: op1_09_inv24 = 1;
    80: op1_09_inv24 = 1;
    82: op1_09_inv24 = 1;
    85: op1_09_inv24 = 1;
    86: op1_09_inv24 = 1;
    87: op1_09_inv24 = 1;
    88: op1_09_inv24 = 1;
    90: op1_09_inv24 = 1;
    94: op1_09_inv24 = 1;
    96: op1_09_inv24 = 1;
    default: op1_09_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の25番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in25 = reg_0023;
    7: op1_09_in25 = reg_0125;
    8: op1_09_in25 = reg_0059;
    9: op1_09_in25 = reg_0166;
    10: op1_09_in25 = imem06_in[95:92];
    61: op1_09_in25 = imem06_in[95:92];
    11: op1_09_in25 = reg_1041;
    12: op1_09_in25 = imem06_in[63:60];
    13: op1_09_in25 = imem03_in[43:40];
    14: op1_09_in25 = reg_0558;
    15: op1_09_in25 = reg_0140;
    16: op1_09_in25 = reg_0246;
    17: op1_09_in25 = reg_0579;
    18: op1_09_in25 = reg_0766;
    19: op1_09_in25 = reg_0365;
    75: op1_09_in25 = reg_0365;
    20: op1_09_in25 = reg_0220;
    43: op1_09_in25 = reg_0220;
    21: op1_09_in25 = imem04_in[75:72];
    23: op1_09_in25 = reg_0170;
    24: op1_09_in25 = reg_0179;
    25: op1_09_in25 = imem01_in[103:100];
    26: op1_09_in25 = reg_0945;
    27: op1_09_in25 = reg_0655;
    28: op1_09_in25 = reg_0217;
    29: op1_09_in25 = imem01_in[11:8];
    30: op1_09_in25 = reg_0555;
    31: op1_09_in25 = reg_0793;
    32: op1_09_in25 = reg_0149;
    33: op1_09_in25 = reg_0722;
    34: op1_09_in25 = reg_0885;
    35: op1_09_in25 = reg_0229;
    36: op1_09_in25 = reg_0022;
    37: op1_09_in25 = imem06_in[87:84];
    38: op1_09_in25 = reg_0954;
    39: op1_09_in25 = reg_0177;
    40: op1_09_in25 = imem01_in[91:88];
    41: op1_09_in25 = imem01_in[15:12];
    42: op1_09_in25 = reg_0489;
    45: op1_09_in25 = reg_0004;
    46: op1_09_in25 = imem04_in[47:44];
    48: op1_09_in25 = reg_0245;
    49: op1_09_in25 = imem04_in[111:108];
    50: op1_09_in25 = reg_0863;
    51: op1_09_in25 = imem01_in[95:92];
    53: op1_09_in25 = reg_0918;
    54: op1_09_in25 = reg_0190;
    55: op1_09_in25 = reg_1002;
    56: op1_09_in25 = imem04_in[15:12];
    57: op1_09_in25 = reg_1057;
    58: op1_09_in25 = reg_0581;
    59: op1_09_in25 = reg_0132;
    60: op1_09_in25 = imem06_in[103:100];
    63: op1_09_in25 = reg_0085;
    64: op1_09_in25 = reg_0099;
    65: op1_09_in25 = reg_1003;
    66: op1_09_in25 = reg_0854;
    67: op1_09_in25 = reg_0799;
    68: op1_09_in25 = reg_0433;
    69: op1_09_in25 = imem01_in[115:112];
    70: op1_09_in25 = reg_0030;
    71: op1_09_in25 = imem06_in[51:48];
    72: op1_09_in25 = imem03_in[59:56];
    73: op1_09_in25 = imem06_in[3:0];
    74: op1_09_in25 = reg_0531;
    77: op1_09_in25 = reg_0832;
    78: op1_09_in25 = reg_0902;
    79: op1_09_in25 = reg_0049;
    80: op1_09_in25 = reg_0150;
    81: op1_09_in25 = reg_0392;
    82: op1_09_in25 = imem05_in[47:44];
    83: op1_09_in25 = reg_0772;
    85: op1_09_in25 = reg_0542;
    86: op1_09_in25 = reg_0270;
    87: op1_09_in25 = reg_0798;
    88: op1_09_in25 = imem04_in[79:76];
    89: op1_09_in25 = reg_0216;
    90: op1_09_in25 = imem04_in[83:80];
    91: op1_09_in25 = imem04_in[83:80];
    92: op1_09_in25 = imem06_in[23:20];
    94: op1_09_in25 = reg_0429;
    95: op1_09_in25 = reg_0714;
    96: op1_09_in25 = reg_0541;
    97: op1_09_in25 = reg_0726;
    default: op1_09_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv25 = 1;
    8: op1_09_inv25 = 1;
    10: op1_09_inv25 = 1;
    11: op1_09_inv25 = 1;
    16: op1_09_inv25 = 1;
    17: op1_09_inv25 = 1;
    20: op1_09_inv25 = 1;
    21: op1_09_inv25 = 1;
    27: op1_09_inv25 = 1;
    28: op1_09_inv25 = 1;
    29: op1_09_inv25 = 1;
    30: op1_09_inv25 = 1;
    33: op1_09_inv25 = 1;
    36: op1_09_inv25 = 1;
    37: op1_09_inv25 = 1;
    39: op1_09_inv25 = 1;
    40: op1_09_inv25 = 1;
    41: op1_09_inv25 = 1;
    42: op1_09_inv25 = 1;
    46: op1_09_inv25 = 1;
    57: op1_09_inv25 = 1;
    59: op1_09_inv25 = 1;
    61: op1_09_inv25 = 1;
    65: op1_09_inv25 = 1;
    66: op1_09_inv25 = 1;
    69: op1_09_inv25 = 1;
    70: op1_09_inv25 = 1;
    77: op1_09_inv25 = 1;
    79: op1_09_inv25 = 1;
    81: op1_09_inv25 = 1;
    83: op1_09_inv25 = 1;
    85: op1_09_inv25 = 1;
    86: op1_09_inv25 = 1;
    90: op1_09_inv25 = 1;
    91: op1_09_inv25 = 1;
    92: op1_09_inv25 = 1;
    94: op1_09_inv25 = 1;
    95: op1_09_inv25 = 1;
    97: op1_09_inv25 = 1;
    default: op1_09_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の26番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in26 = imem07_in[15:12];
    7: op1_09_in26 = reg_0107;
    8: op1_09_in26 = reg_0076;
    9: op1_09_in26 = reg_0178;
    10: op1_09_in26 = imem06_in[99:96];
    11: op1_09_in26 = reg_0109;
    12: op1_09_in26 = reg_0610;
    13: op1_09_in26 = imem03_in[59:56];
    14: op1_09_in26 = reg_0531;
    15: op1_09_in26 = imem06_in[3:0];
    16: op1_09_in26 = reg_0242;
    17: op1_09_in26 = reg_0572;
    18: op1_09_in26 = reg_0234;
    19: op1_09_in26 = reg_0342;
    20: op1_09_in26 = reg_0237;
    21: op1_09_in26 = imem04_in[103:100];
    24: op1_09_in26 = reg_0162;
    25: op1_09_in26 = reg_0226;
    26: op1_09_in26 = reg_0489;
    27: op1_09_in26 = reg_0640;
    28: op1_09_in26 = reg_0925;
    29: op1_09_in26 = imem01_in[35:32];
    30: op1_09_in26 = reg_0236;
    31: op1_09_in26 = reg_0767;
    32: op1_09_in26 = reg_0133;
    33: op1_09_in26 = reg_0710;
    34: op1_09_in26 = reg_0500;
    35: op1_09_in26 = reg_0257;
    36: op1_09_in26 = reg_0827;
    37: op1_09_in26 = imem06_in[107:104];
    60: op1_09_in26 = imem06_in[107:104];
    38: op1_09_in26 = reg_0946;
    39: op1_09_in26 = reg_0158;
    40: op1_09_in26 = imem01_in[95:92];
    41: op1_09_in26 = imem01_in[107:104];
    51: op1_09_in26 = imem01_in[107:104];
    42: op1_09_in26 = reg_0132;
    43: op1_09_in26 = reg_0856;
    45: op1_09_in26 = reg_0543;
    46: op1_09_in26 = imem04_in[51:48];
    48: op1_09_in26 = reg_0327;
    49: op1_09_in26 = imem05_in[19:16];
    50: op1_09_in26 = reg_0081;
    53: op1_09_in26 = reg_0779;
    54: op1_09_in26 = imem01_in[11:8];
    55: op1_09_in26 = reg_0974;
    56: op1_09_in26 = imem04_in[27:24];
    57: op1_09_in26 = reg_1020;
    58: op1_09_in26 = reg_0675;
    59: op1_09_in26 = reg_0135;
    61: op1_09_in26 = imem07_in[51:48];
    63: op1_09_in26 = reg_0049;
    64: op1_09_in26 = reg_0760;
    65: op1_09_in26 = reg_0511;
    66: op1_09_in26 = reg_0824;
    67: op1_09_in26 = reg_0848;
    68: op1_09_in26 = reg_0024;
    69: op1_09_in26 = reg_0522;
    70: op1_09_in26 = reg_0949;
    71: op1_09_in26 = imem06_in[95:92];
    72: op1_09_in26 = imem03_in[75:72];
    73: op1_09_in26 = imem06_in[47:44];
    74: op1_09_in26 = reg_0958;
    75: op1_09_in26 = imem07_in[11:8];
    77: op1_09_in26 = reg_0111;
    78: op1_09_in26 = reg_0521;
    79: op1_09_in26 = imem03_in[11:8];
    80: op1_09_in26 = reg_0947;
    81: op1_09_in26 = reg_0632;
    82: op1_09_in26 = imem05_in[107:104];
    83: op1_09_in26 = reg_0007;
    85: op1_09_in26 = reg_0295;
    86: op1_09_in26 = reg_0022;
    87: op1_09_in26 = reg_0869;
    88: op1_09_in26 = imem04_in[95:92];
    89: op1_09_in26 = reg_0737;
    90: op1_09_in26 = reg_0942;
    91: op1_09_in26 = imem04_in[107:104];
    92: op1_09_in26 = imem06_in[43:40];
    94: op1_09_in26 = reg_0714;
    95: op1_09_in26 = reg_0701;
    96: op1_09_in26 = reg_0789;
    97: op1_09_in26 = reg_0247;
    default: op1_09_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv26 = 1;
    8: op1_09_inv26 = 1;
    11: op1_09_inv26 = 1;
    13: op1_09_inv26 = 1;
    14: op1_09_inv26 = 1;
    15: op1_09_inv26 = 1;
    18: op1_09_inv26 = 1;
    20: op1_09_inv26 = 1;
    24: op1_09_inv26 = 1;
    25: op1_09_inv26 = 1;
    26: op1_09_inv26 = 1;
    30: op1_09_inv26 = 1;
    31: op1_09_inv26 = 1;
    34: op1_09_inv26 = 1;
    37: op1_09_inv26 = 1;
    40: op1_09_inv26 = 1;
    42: op1_09_inv26 = 1;
    43: op1_09_inv26 = 1;
    45: op1_09_inv26 = 1;
    46: op1_09_inv26 = 1;
    48: op1_09_inv26 = 1;
    49: op1_09_inv26 = 1;
    50: op1_09_inv26 = 1;
    54: op1_09_inv26 = 1;
    57: op1_09_inv26 = 1;
    60: op1_09_inv26 = 1;
    61: op1_09_inv26 = 1;
    65: op1_09_inv26 = 1;
    71: op1_09_inv26 = 1;
    72: op1_09_inv26 = 1;
    73: op1_09_inv26 = 1;
    74: op1_09_inv26 = 1;
    75: op1_09_inv26 = 1;
    79: op1_09_inv26 = 1;
    80: op1_09_inv26 = 1;
    83: op1_09_inv26 = 1;
    88: op1_09_inv26 = 1;
    92: op1_09_inv26 = 1;
    95: op1_09_inv26 = 1;
    96: op1_09_inv26 = 1;
    97: op1_09_inv26 = 1;
    default: op1_09_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の27番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in27 = imem07_in[51:48];
    75: op1_09_in27 = imem07_in[51:48];
    7: op1_09_in27 = imem02_in[31:28];
    8: op1_09_in27 = reg_0048;
    9: op1_09_in27 = reg_0157;
    10: op1_09_in27 = reg_0625;
    11: op1_09_in27 = reg_0107;
    12: op1_09_in27 = reg_0626;
    13: op1_09_in27 = imem03_in[67:64];
    14: op1_09_in27 = reg_0541;
    15: op1_09_in27 = imem06_in[39:36];
    16: op1_09_in27 = reg_0503;
    17: op1_09_in27 = reg_0576;
    18: op1_09_in27 = reg_0508;
    19: op1_09_in27 = reg_0314;
    20: op1_09_in27 = reg_0245;
    21: op1_09_in27 = reg_0543;
    24: op1_09_in27 = reg_0166;
    25: op1_09_in27 = reg_0496;
    26: op1_09_in27 = reg_0497;
    27: op1_09_in27 = reg_0863;
    28: op1_09_in27 = reg_0589;
    29: op1_09_in27 = imem01_in[39:36];
    30: op1_09_in27 = reg_0274;
    31: op1_09_in27 = reg_0822;
    32: op1_09_in27 = reg_0151;
    33: op1_09_in27 = reg_0717;
    34: op1_09_in27 = reg_1045;
    35: op1_09_in27 = reg_0819;
    36: op1_09_in27 = reg_0816;
    37: op1_09_in27 = imem07_in[19:16];
    38: op1_09_in27 = reg_0834;
    40: op1_09_in27 = imem01_in[103:100];
    41: op1_09_in27 = imem01_in[111:108];
    42: op1_09_in27 = reg_0145;
    43: op1_09_in27 = reg_0892;
    45: op1_09_in27 = reg_0795;
    46: op1_09_in27 = imem04_in[111:108];
    48: op1_09_in27 = reg_0346;
    49: op1_09_in27 = imem05_in[35:32];
    50: op1_09_in27 = reg_0225;
    51: op1_09_in27 = reg_0918;
    53: op1_09_in27 = reg_0223;
    54: op1_09_in27 = imem01_in[31:28];
    55: op1_09_in27 = reg_0990;
    56: op1_09_in27 = reg_0483;
    57: op1_09_in27 = reg_0292;
    58: op1_09_in27 = reg_0221;
    59: op1_09_in27 = reg_0133;
    60: op1_09_in27 = imem06_in[111:108];
    61: op1_09_in27 = imem07_in[63:60];
    63: op1_09_in27 = reg_0840;
    64: op1_09_in27 = reg_0445;
    65: op1_09_in27 = reg_0282;
    66: op1_09_in27 = reg_0650;
    67: op1_09_in27 = reg_0068;
    68: op1_09_in27 = reg_0176;
    69: op1_09_in27 = reg_0514;
    70: op1_09_in27 = reg_0953;
    71: op1_09_in27 = imem06_in[99:96];
    72: op1_09_in27 = imem03_in[79:76];
    73: op1_09_in27 = imem06_in[71:68];
    92: op1_09_in27 = imem06_in[71:68];
    74: op1_09_in27 = reg_0509;
    77: op1_09_in27 = reg_1053;
    78: op1_09_in27 = reg_0906;
    79: op1_09_in27 = imem03_in[15:12];
    80: op1_09_in27 = reg_1015;
    81: op1_09_in27 = reg_0380;
    82: op1_09_in27 = reg_0636;
    83: op1_09_in27 = reg_0482;
    85: op1_09_in27 = imem05_in[39:36];
    86: op1_09_in27 = imem07_in[43:40];
    87: op1_09_in27 = reg_0216;
    88: op1_09_in27 = imem04_in[127:124];
    89: op1_09_in27 = reg_0610;
    90: op1_09_in27 = reg_0446;
    91: op1_09_in27 = reg_0942;
    94: op1_09_in27 = reg_0701;
    95: op1_09_in27 = reg_0449;
    96: op1_09_in27 = reg_0968;
    97: op1_09_in27 = reg_0715;
    default: op1_09_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_09_inv27 = 1;
    10: op1_09_inv27 = 1;
    12: op1_09_inv27 = 1;
    13: op1_09_inv27 = 1;
    14: op1_09_inv27 = 1;
    15: op1_09_inv27 = 1;
    16: op1_09_inv27 = 1;
    17: op1_09_inv27 = 1;
    19: op1_09_inv27 = 1;
    24: op1_09_inv27 = 1;
    25: op1_09_inv27 = 1;
    26: op1_09_inv27 = 1;
    27: op1_09_inv27 = 1;
    31: op1_09_inv27 = 1;
    33: op1_09_inv27 = 1;
    35: op1_09_inv27 = 1;
    36: op1_09_inv27 = 1;
    38: op1_09_inv27 = 1;
    42: op1_09_inv27 = 1;
    43: op1_09_inv27 = 1;
    45: op1_09_inv27 = 1;
    46: op1_09_inv27 = 1;
    50: op1_09_inv27 = 1;
    51: op1_09_inv27 = 1;
    54: op1_09_inv27 = 1;
    55: op1_09_inv27 = 1;
    61: op1_09_inv27 = 1;
    63: op1_09_inv27 = 1;
    67: op1_09_inv27 = 1;
    70: op1_09_inv27 = 1;
    77: op1_09_inv27 = 1;
    78: op1_09_inv27 = 1;
    79: op1_09_inv27 = 1;
    80: op1_09_inv27 = 1;
    82: op1_09_inv27 = 1;
    83: op1_09_inv27 = 1;
    85: op1_09_inv27 = 1;
    90: op1_09_inv27 = 1;
    91: op1_09_inv27 = 1;
    92: op1_09_inv27 = 1;
    94: op1_09_inv27 = 1;
    95: op1_09_inv27 = 1;
    default: op1_09_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の28番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in28 = imem07_in[115:112];
    7: op1_09_in28 = imem02_in[123:120];
    8: op1_09_in28 = imem05_in[7:4];
    10: op1_09_in28 = reg_0607;
    11: op1_09_in28 = reg_0117;
    12: op1_09_in28 = reg_0608;
    13: op1_09_in28 = reg_0596;
    14: op1_09_in28 = reg_0547;
    15: op1_09_in28 = imem06_in[43:40];
    16: op1_09_in28 = reg_0905;
    17: op1_09_in28 = reg_0394;
    18: op1_09_in28 = reg_1035;
    19: op1_09_in28 = reg_0092;
    20: op1_09_in28 = reg_0226;
    21: op1_09_in28 = reg_0557;
    24: op1_09_in28 = reg_0176;
    25: op1_09_in28 = reg_1033;
    26: op1_09_in28 = reg_0147;
    88: op1_09_in28 = reg_0147;
    27: op1_09_in28 = reg_0080;
    28: op1_09_in28 = reg_0585;
    29: op1_09_in28 = imem01_in[51:48];
    30: op1_09_in28 = reg_0221;
    31: op1_09_in28 = reg_1002;
    32: op1_09_in28 = reg_0134;
    33: op1_09_in28 = reg_0708;
    34: op1_09_in28 = reg_0104;
    35: op1_09_in28 = reg_0489;
    36: op1_09_in28 = reg_0489;
    37: op1_09_in28 = imem07_in[31:28];
    38: op1_09_in28 = reg_0757;
    40: op1_09_in28 = imem01_in[111:108];
    41: op1_09_in28 = imem01_in[115:112];
    42: op1_09_in28 = reg_0133;
    43: op1_09_in28 = reg_0627;
    45: op1_09_in28 = reg_0311;
    46: op1_09_in28 = imem05_in[3:0];
    48: op1_09_in28 = reg_0004;
    49: op1_09_in28 = imem05_in[39:36];
    50: op1_09_in28 = reg_0085;
    51: op1_09_in28 = reg_0586;
    53: op1_09_in28 = reg_1044;
    54: op1_09_in28 = imem01_in[79:76];
    55: op1_09_in28 = imem04_in[35:32];
    56: op1_09_in28 = reg_0306;
    57: op1_09_in28 = reg_0541;
    58: op1_09_in28 = reg_0785;
    59: op1_09_in28 = reg_0151;
    60: op1_09_in28 = imem06_in[119:116];
    61: op1_09_in28 = imem07_in[95:92];
    63: op1_09_in28 = reg_0310;
    64: op1_09_in28 = reg_0577;
    65: op1_09_in28 = reg_0055;
    66: op1_09_in28 = reg_0951;
    67: op1_09_in28 = reg_0015;
    69: op1_09_in28 = reg_0830;
    70: op1_09_in28 = reg_0675;
    71: op1_09_in28 = imem07_in[15:12];
    72: op1_09_in28 = imem03_in[119:116];
    73: op1_09_in28 = imem06_in[95:92];
    74: op1_09_in28 = reg_0129;
    75: op1_09_in28 = imem07_in[59:56];
    77: op1_09_in28 = reg_0555;
    78: op1_09_in28 = reg_0232;
    79: op1_09_in28 = imem03_in[31:28];
    80: op1_09_in28 = reg_1046;
    81: op1_09_in28 = reg_0695;
    82: op1_09_in28 = reg_0128;
    83: op1_09_in28 = reg_0776;
    85: op1_09_in28 = imem05_in[63:60];
    86: op1_09_in28 = imem07_in[91:88];
    87: op1_09_in28 = reg_0512;
    89: op1_09_in28 = reg_0769;
    90: op1_09_in28 = reg_0511;
    91: op1_09_in28 = reg_0048;
    92: op1_09_in28 = imem06_in[111:108];
    94: op1_09_in28 = reg_0697;
    95: op1_09_in28 = reg_0724;
    96: op1_09_in28 = reg_0592;
    97: op1_09_in28 = reg_0321;
    default: op1_09_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv28 = 1;
    11: op1_09_inv28 = 1;
    12: op1_09_inv28 = 1;
    15: op1_09_inv28 = 1;
    19: op1_09_inv28 = 1;
    20: op1_09_inv28 = 1;
    21: op1_09_inv28 = 1;
    24: op1_09_inv28 = 1;
    26: op1_09_inv28 = 1;
    27: op1_09_inv28 = 1;
    29: op1_09_inv28 = 1;
    35: op1_09_inv28 = 1;
    36: op1_09_inv28 = 1;
    38: op1_09_inv28 = 1;
    40: op1_09_inv28 = 1;
    41: op1_09_inv28 = 1;
    45: op1_09_inv28 = 1;
    48: op1_09_inv28 = 1;
    50: op1_09_inv28 = 1;
    55: op1_09_inv28 = 1;
    56: op1_09_inv28 = 1;
    59: op1_09_inv28 = 1;
    61: op1_09_inv28 = 1;
    63: op1_09_inv28 = 1;
    64: op1_09_inv28 = 1;
    66: op1_09_inv28 = 1;
    67: op1_09_inv28 = 1;
    70: op1_09_inv28 = 1;
    75: op1_09_inv28 = 1;
    77: op1_09_inv28 = 1;
    79: op1_09_inv28 = 1;
    82: op1_09_inv28 = 1;
    83: op1_09_inv28 = 1;
    86: op1_09_inv28 = 1;
    87: op1_09_inv28 = 1;
    88: op1_09_inv28 = 1;
    92: op1_09_inv28 = 1;
    94: op1_09_inv28 = 1;
    95: op1_09_inv28 = 1;
    default: op1_09_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の29番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in29 = reg_0728;
    7: op1_09_in29 = reg_0642;
    8: op1_09_in29 = imem05_in[39:36];
    10: op1_09_in29 = reg_0631;
    11: op1_09_in29 = imem02_in[3:0];
    12: op1_09_in29 = reg_0349;
    13: op1_09_in29 = reg_0587;
    14: op1_09_in29 = reg_0301;
    15: op1_09_in29 = imem06_in[47:44];
    16: op1_09_in29 = reg_1039;
    17: op1_09_in29 = reg_0373;
    18: op1_09_in29 = reg_1031;
    19: op1_09_in29 = reg_0085;
    20: op1_09_in29 = reg_0496;
    21: op1_09_in29 = reg_0552;
    25: op1_09_in29 = reg_0871;
    26: op1_09_in29 = reg_0145;
    27: op1_09_in29 = reg_0095;
    28: op1_09_in29 = reg_0588;
    29: op1_09_in29 = imem01_in[67:64];
    30: op1_09_in29 = reg_0249;
    31: op1_09_in29 = reg_0995;
    32: op1_09_in29 = reg_0921;
    33: op1_09_in29 = reg_0713;
    34: op1_09_in29 = reg_0108;
    35: op1_09_in29 = reg_0132;
    36: op1_09_in29 = reg_0132;
    37: op1_09_in29 = imem07_in[63:60];
    38: op1_09_in29 = reg_0275;
    40: op1_09_in29 = imem01_in[119:116];
    41: op1_09_in29 = reg_0111;
    42: op1_09_in29 = reg_0129;
    43: op1_09_in29 = reg_0042;
    45: op1_09_in29 = reg_0369;
    46: op1_09_in29 = imem05_in[7:4];
    48: op1_09_in29 = reg_0833;
    49: op1_09_in29 = imem05_in[43:40];
    50: op1_09_in29 = reg_0792;
    51: op1_09_in29 = reg_0223;
    53: op1_09_in29 = reg_1056;
    54: op1_09_in29 = imem01_in[99:96];
    55: op1_09_in29 = imem04_in[63:60];
    56: op1_09_in29 = reg_0909;
    57: op1_09_in29 = reg_0850;
    58: op1_09_in29 = reg_0032;
    59: op1_09_in29 = reg_0152;
    60: op1_09_in29 = reg_0010;
    61: op1_09_in29 = imem07_in[115:112];
    63: op1_09_in29 = reg_0872;
    64: op1_09_in29 = reg_0661;
    65: op1_09_in29 = reg_0888;
    66: op1_09_in29 = reg_0667;
    67: op1_09_in29 = reg_0072;
    69: op1_09_in29 = reg_0610;
    70: op1_09_in29 = reg_0508;
    71: op1_09_in29 = imem07_in[31:28];
    72: op1_09_in29 = reg_0445;
    73: op1_09_in29 = imem06_in[119:116];
    92: op1_09_in29 = imem06_in[119:116];
    74: op1_09_in29 = reg_0946;
    75: op1_09_in29 = imem07_in[75:72];
    77: op1_09_in29 = reg_0114;
    78: op1_09_in29 = reg_0114;
    89: op1_09_in29 = reg_0114;
    79: op1_09_in29 = imem03_in[39:36];
    80: op1_09_in29 = reg_0957;
    81: op1_09_in29 = reg_0834;
    82: op1_09_in29 = reg_0319;
    83: op1_09_in29 = reg_0867;
    85: op1_09_in29 = imem05_in[83:80];
    86: op1_09_in29 = imem07_in[95:92];
    87: op1_09_in29 = reg_1053;
    88: op1_09_in29 = reg_1009;
    90: op1_09_in29 = reg_0550;
    91: op1_09_in29 = reg_0430;
    96: op1_09_in29 = reg_0237;
    97: op1_09_in29 = reg_0589;
    default: op1_09_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv29 = 1;
    7: op1_09_inv29 = 1;
    8: op1_09_inv29 = 1;
    10: op1_09_inv29 = 1;
    12: op1_09_inv29 = 1;
    13: op1_09_inv29 = 1;
    14: op1_09_inv29 = 1;
    15: op1_09_inv29 = 1;
    18: op1_09_inv29 = 1;
    19: op1_09_inv29 = 1;
    20: op1_09_inv29 = 1;
    21: op1_09_inv29 = 1;
    26: op1_09_inv29 = 1;
    28: op1_09_inv29 = 1;
    30: op1_09_inv29 = 1;
    31: op1_09_inv29 = 1;
    32: op1_09_inv29 = 1;
    33: op1_09_inv29 = 1;
    34: op1_09_inv29 = 1;
    35: op1_09_inv29 = 1;
    40: op1_09_inv29 = 1;
    41: op1_09_inv29 = 1;
    42: op1_09_inv29 = 1;
    43: op1_09_inv29 = 1;
    46: op1_09_inv29 = 1;
    51: op1_09_inv29 = 1;
    53: op1_09_inv29 = 1;
    57: op1_09_inv29 = 1;
    63: op1_09_inv29 = 1;
    71: op1_09_inv29 = 1;
    74: op1_09_inv29 = 1;
    81: op1_09_inv29 = 1;
    82: op1_09_inv29 = 1;
    83: op1_09_inv29 = 1;
    85: op1_09_inv29 = 1;
    86: op1_09_inv29 = 1;
    87: op1_09_inv29 = 1;
    88: op1_09_inv29 = 1;
    89: op1_09_inv29 = 1;
    91: op1_09_inv29 = 1;
    default: op1_09_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の30番目の入力
  always @ ( * ) begin
    case ( state )
    6: op1_09_in30 = reg_0702;
    7: op1_09_in30 = reg_0646;
    8: op1_09_in30 = imem05_in[79:76];
    10: op1_09_in30 = reg_0626;
    11: op1_09_in30 = imem02_in[31:28];
    12: op1_09_in30 = reg_0404;
    13: op1_09_in30 = reg_0592;
    53: op1_09_in30 = reg_0592;
    14: op1_09_in30 = reg_0306;
    15: op1_09_in30 = reg_0835;
    16: op1_09_in30 = reg_1042;
    17: op1_09_in30 = reg_0322;
    18: op1_09_in30 = reg_0913;
    19: op1_09_in30 = imem03_in[59:56];
    20: op1_09_in30 = reg_1032;
    21: op1_09_in30 = reg_0555;
    25: op1_09_in30 = reg_1017;
    69: op1_09_in30 = reg_1017;
    26: op1_09_in30 = reg_0128;
    27: op1_09_in30 = reg_0865;
    28: op1_09_in30 = imem03_in[3:0];
    29: op1_09_in30 = imem01_in[79:76];
    30: op1_09_in30 = reg_0769;
    31: op1_09_in30 = reg_0984;
    32: op1_09_in30 = reg_0894;
    33: op1_09_in30 = reg_0701;
    34: op1_09_in30 = reg_0114;
    35: op1_09_in30 = reg_0135;
    36: op1_09_in30 = reg_0135;
    37: op1_09_in30 = imem07_in[75:72];
    38: op1_09_in30 = reg_1046;
    40: op1_09_in30 = reg_0123;
    41: op1_09_in30 = reg_0100;
    86: op1_09_in30 = reg_0100;
    42: op1_09_in30 = reg_0140;
    43: op1_09_in30 = reg_0295;
    45: op1_09_in30 = reg_0807;
    46: op1_09_in30 = imem05_in[123:120];
    48: op1_09_in30 = reg_0373;
    49: op1_09_in30 = imem05_in[91:88];
    50: op1_09_in30 = reg_0814;
    51: op1_09_in30 = reg_0218;
    54: op1_09_in30 = imem01_in[123:120];
    55: op1_09_in30 = imem04_in[103:100];
    56: op1_09_in30 = reg_0802;
    57: op1_09_in30 = reg_0076;
    58: op1_09_in30 = reg_0508;
    59: op1_09_in30 = reg_0154;
    60: op1_09_in30 = reg_0625;
    61: op1_09_in30 = reg_0722;
    63: op1_09_in30 = reg_0079;
    64: op1_09_in30 = reg_0040;
    65: op1_09_in30 = reg_0931;
    66: op1_09_in30 = reg_0490;
    67: op1_09_in30 = reg_0764;
    70: op1_09_in30 = reg_0786;
    71: op1_09_in30 = imem07_in[59:56];
    72: op1_09_in30 = reg_0434;
    73: op1_09_in30 = reg_0391;
    74: op1_09_in30 = reg_0134;
    75: op1_09_in30 = imem07_in[83:80];
    77: op1_09_in30 = reg_0860;
    78: op1_09_in30 = reg_0860;
    79: op1_09_in30 = imem03_in[47:44];
    80: op1_09_in30 = reg_0145;
    81: op1_09_in30 = reg_0017;
    82: op1_09_in30 = reg_0448;
    83: op1_09_in30 = reg_0086;
    85: op1_09_in30 = imem05_in[87:84];
    87: op1_09_in30 = reg_1033;
    88: op1_09_in30 = reg_0014;
    89: op1_09_in30 = reg_0109;
    90: op1_09_in30 = reg_0016;
    91: op1_09_in30 = reg_0008;
    92: op1_09_in30 = reg_0021;
    96: op1_09_in30 = reg_0544;
    97: op1_09_in30 = reg_0024;
    default: op1_09_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv30 = 1;
    7: op1_09_inv30 = 1;
    10: op1_09_inv30 = 1;
    11: op1_09_inv30 = 1;
    14: op1_09_inv30 = 1;
    17: op1_09_inv30 = 1;
    25: op1_09_inv30 = 1;
    26: op1_09_inv30 = 1;
    27: op1_09_inv30 = 1;
    28: op1_09_inv30 = 1;
    29: op1_09_inv30 = 1;
    31: op1_09_inv30 = 1;
    32: op1_09_inv30 = 1;
    34: op1_09_inv30 = 1;
    37: op1_09_inv30 = 1;
    38: op1_09_inv30 = 1;
    40: op1_09_inv30 = 1;
    42: op1_09_inv30 = 1;
    46: op1_09_inv30 = 1;
    49: op1_09_inv30 = 1;
    53: op1_09_inv30 = 1;
    63: op1_09_inv30 = 1;
    64: op1_09_inv30 = 1;
    65: op1_09_inv30 = 1;
    69: op1_09_inv30 = 1;
    80: op1_09_inv30 = 1;
    81: op1_09_inv30 = 1;
    83: op1_09_inv30 = 1;
    96: op1_09_inv30 = 1;
    97: op1_09_inv30 = 1;
    default: op1_09_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_09_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_09_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in00 = imem00_in[103:100];
    6: op1_10_in00 = imem00_in[31:28];
    93: op1_10_in00 = imem00_in[31:28];
    7: op1_10_in00 = reg_0664;
    8: op1_10_in00 = imem05_in[107:104];
    9: op1_10_in00 = imem00_in[47:44];
    10: op1_10_in00 = reg_0601;
    11: op1_10_in00 = imem02_in[83:80];
    12: op1_10_in00 = reg_0367;
    13: op1_10_in00 = reg_0589;
    14: op1_10_in00 = reg_0302;
    57: op1_10_in00 = reg_0302;
    15: op1_10_in00 = imem06_in[59:56];
    16: op1_10_in00 = reg_0885;
    17: op1_10_in00 = reg_0331;
    4: op1_10_in00 = imem07_in[31:28];
    18: op1_10_in00 = reg_0904;
    19: op1_10_in00 = imem03_in[79:76];
    20: op1_10_in00 = reg_1040;
    21: op1_10_in00 = reg_0551;
    22: op1_10_in00 = reg_0685;
    23: op1_10_in00 = imem00_in[59:56];
    24: op1_10_in00 = imem00_in[3:0];
    47: op1_10_in00 = imem00_in[3:0];
    25: op1_10_in00 = reg_0105;
    3: op1_10_in00 = imem07_in[107:104];
    71: op1_10_in00 = imem07_in[107:104];
    26: op1_10_in00 = reg_0156;
    27: op1_10_in00 = reg_0083;
    28: op1_10_in00 = imem03_in[27:24];
    29: op1_10_in00 = imem01_in[95:92];
    30: op1_10_in00 = reg_1042;
    31: op1_10_in00 = reg_0990;
    2: op1_10_in00 = imem07_in[67:64];
    32: op1_10_in00 = reg_0925;
    69: op1_10_in00 = reg_0925;
    33: op1_10_in00 = reg_0706;
    34: op1_10_in00 = reg_0100;
    35: op1_10_in00 = reg_0150;
    36: op1_10_in00 = reg_0154;
    37: op1_10_in00 = imem07_in[79:76];
    38: op1_10_in00 = reg_0254;
    39: op1_10_in00 = imem00_in[15:12];
    68: op1_10_in00 = imem00_in[15:12];
    76: op1_10_in00 = imem00_in[15:12];
    94: op1_10_in00 = imem00_in[15:12];
    40: op1_10_in00 = reg_0111;
    41: op1_10_in00 = reg_0106;
    42: op1_10_in00 = reg_0131;
    43: op1_10_in00 = reg_0383;
    44: op1_10_in00 = imem00_in[19:16];
    45: op1_10_in00 = reg_0376;
    46: op1_10_in00 = reg_0958;
    48: op1_10_in00 = reg_0051;
    49: op1_10_in00 = reg_0962;
    50: op1_10_in00 = reg_0506;
    51: op1_10_in00 = reg_0871;
    52: op1_10_in00 = imem00_in[7:4];
    84: op1_10_in00 = imem00_in[7:4];
    53: op1_10_in00 = reg_1035;
    54: op1_10_in00 = reg_1056;
    55: op1_10_in00 = imem04_in[111:108];
    56: op1_10_in00 = reg_0068;
    58: op1_10_in00 = reg_0813;
    59: op1_10_in00 = reg_0129;
    60: op1_10_in00 = reg_0694;
    61: op1_10_in00 = reg_0704;
    62: op1_10_in00 = imem00_in[67:64];
    63: op1_10_in00 = imem03_in[11:8];
    64: op1_10_in00 = reg_0509;
    65: op1_10_in00 = reg_0932;
    66: op1_10_in00 = reg_0950;
    67: op1_10_in00 = reg_0065;
    70: op1_10_in00 = reg_0972;
    72: op1_10_in00 = reg_0298;
    73: op1_10_in00 = reg_0626;
    74: op1_10_in00 = reg_0943;
    75: op1_10_in00 = imem07_in[87:84];
    77: op1_10_in00 = reg_0115;
    78: op1_10_in00 = reg_0113;
    79: op1_10_in00 = imem03_in[71:68];
    80: op1_10_in00 = reg_0135;
    81: op1_10_in00 = reg_0755;
    82: op1_10_in00 = reg_0137;
    83: op1_10_in00 = imem03_in[7:4];
    85: op1_10_in00 = imem05_in[111:108];
    86: op1_10_in00 = reg_0653;
    87: op1_10_in00 = reg_0555;
    88: op1_10_in00 = reg_0809;
    89: op1_10_in00 = imem02_in[39:36];
    90: op1_10_in00 = reg_0537;
    91: op1_10_in00 = reg_0537;
    92: op1_10_in00 = reg_0692;
    95: op1_10_in00 = imem00_in[71:68];
    96: op1_10_in00 = imem01_in[11:8];
    97: op1_10_in00 = reg_0640;
    default: op1_10_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv00 = 1;
    6: op1_10_inv00 = 1;
    11: op1_10_inv00 = 1;
    13: op1_10_inv00 = 1;
    14: op1_10_inv00 = 1;
    15: op1_10_inv00 = 1;
    17: op1_10_inv00 = 1;
    18: op1_10_inv00 = 1;
    19: op1_10_inv00 = 1;
    20: op1_10_inv00 = 1;
    21: op1_10_inv00 = 1;
    22: op1_10_inv00 = 1;
    24: op1_10_inv00 = 1;
    3: op1_10_inv00 = 1;
    27: op1_10_inv00 = 1;
    28: op1_10_inv00 = 1;
    29: op1_10_inv00 = 1;
    2: op1_10_inv00 = 1;
    33: op1_10_inv00 = 1;
    36: op1_10_inv00 = 1;
    37: op1_10_inv00 = 1;
    38: op1_10_inv00 = 1;
    41: op1_10_inv00 = 1;
    43: op1_10_inv00 = 1;
    45: op1_10_inv00 = 1;
    46: op1_10_inv00 = 1;
    47: op1_10_inv00 = 1;
    52: op1_10_inv00 = 1;
    57: op1_10_inv00 = 1;
    58: op1_10_inv00 = 1;
    60: op1_10_inv00 = 1;
    62: op1_10_inv00 = 1;
    63: op1_10_inv00 = 1;
    67: op1_10_inv00 = 1;
    69: op1_10_inv00 = 1;
    70: op1_10_inv00 = 1;
    71: op1_10_inv00 = 1;
    72: op1_10_inv00 = 1;
    76: op1_10_inv00 = 1;
    78: op1_10_inv00 = 1;
    83: op1_10_inv00 = 1;
    87: op1_10_inv00 = 1;
    88: op1_10_inv00 = 1;
    89: op1_10_inv00 = 1;
    90: op1_10_inv00 = 1;
    93: op1_10_inv00 = 1;
    94: op1_10_inv00 = 1;
    default: op1_10_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in01 = imem00_in[115:112];
    6: op1_10_in01 = imem00_in[35:32];
    7: op1_10_in01 = reg_0663;
    8: op1_10_in01 = reg_0970;
    9: op1_10_in01 = imem00_in[51:48];
    44: op1_10_in01 = imem00_in[51:48];
    10: op1_10_in01 = reg_0356;
    11: op1_10_in01 = reg_0650;
    12: op1_10_in01 = reg_0780;
    13: op1_10_in01 = reg_0580;
    14: op1_10_in01 = reg_0293;
    15: op1_10_in01 = reg_0614;
    92: op1_10_in01 = reg_0614;
    16: op1_10_in01 = reg_1044;
    17: op1_10_in01 = reg_0992;
    4: op1_10_in01 = imem07_in[39:36];
    18: op1_10_in01 = reg_0118;
    19: op1_10_in01 = imem03_in[91:88];
    20: op1_10_in01 = reg_0111;
    21: op1_10_in01 = reg_0061;
    22: op1_10_in01 = reg_0686;
    23: op1_10_in01 = imem00_in[103:100];
    24: op1_10_in01 = imem00_in[11:8];
    84: op1_10_in01 = imem00_in[11:8];
    25: op1_10_in01 = reg_0122;
    3: op1_10_in01 = imem07_in[111:108];
    75: op1_10_in01 = imem07_in[111:108];
    26: op1_10_in01 = reg_0154;
    27: op1_10_in01 = reg_0086;
    28: op1_10_in01 = imem03_in[31:28];
    83: op1_10_in01 = imem03_in[31:28];
    29: op1_10_in01 = reg_0003;
    30: op1_10_in01 = reg_0230;
    31: op1_10_in01 = reg_1000;
    2: op1_10_in01 = imem07_in[103:100];
    32: op1_10_in01 = reg_0926;
    33: op1_10_in01 = reg_0436;
    34: op1_10_in01 = reg_0127;
    35: op1_10_in01 = reg_0156;
    36: op1_10_in01 = reg_0129;
    37: op1_10_in01 = imem07_in[91:88];
    38: op1_10_in01 = reg_0128;
    39: op1_10_in01 = imem00_in[47:44];
    40: op1_10_in01 = reg_0116;
    41: op1_10_in01 = reg_0115;
    42: op1_10_in01 = imem06_in[11:8];
    43: op1_10_in01 = reg_0380;
    45: op1_10_in01 = reg_0844;
    46: op1_10_in01 = reg_0971;
    47: op1_10_in01 = imem00_in[31:28];
    48: op1_10_in01 = reg_0822;
    49: op1_10_in01 = reg_0963;
    50: op1_10_in01 = reg_0091;
    51: op1_10_in01 = reg_1031;
    52: op1_10_in01 = imem00_in[15:12];
    53: op1_10_in01 = reg_0236;
    54: op1_10_in01 = reg_0285;
    55: op1_10_in01 = reg_0048;
    56: op1_10_in01 = reg_0809;
    57: op1_10_in01 = reg_0296;
    58: op1_10_in01 = reg_0336;
    59: op1_10_in01 = imem06_in[35:32];
    60: op1_10_in01 = reg_0393;
    61: op1_10_in01 = reg_0712;
    62: op1_10_in01 = imem00_in[83:80];
    63: op1_10_in01 = imem03_in[63:60];
    64: op1_10_in01 = reg_0836;
    65: op1_10_in01 = reg_0568;
    66: op1_10_in01 = reg_0968;
    67: op1_10_in01 = reg_0108;
    68: op1_10_in01 = imem00_in[59:56];
    69: op1_10_in01 = reg_1055;
    70: op1_10_in01 = reg_0136;
    71: op1_10_in01 = reg_0719;
    72: op1_10_in01 = reg_0239;
    73: op1_10_in01 = reg_0338;
    74: op1_10_in01 = reg_0866;
    76: op1_10_in01 = imem00_in[23:20];
    77: op1_10_in01 = reg_0113;
    78: op1_10_in01 = imem02_in[15:12];
    79: op1_10_in01 = imem03_in[107:104];
    80: op1_10_in01 = reg_0146;
    81: op1_10_in01 = reg_1010;
    82: op1_10_in01 = reg_0689;
    85: op1_10_in01 = reg_1021;
    86: op1_10_in01 = reg_0589;
    87: op1_10_in01 = imem02_in[35:32];
    88: op1_10_in01 = reg_0407;
    89: op1_10_in01 = imem02_in[47:44];
    90: op1_10_in01 = reg_0848;
    91: op1_10_in01 = reg_0123;
    93: op1_10_in01 = imem00_in[55:52];
    94: op1_10_in01 = imem00_in[19:16];
    95: op1_10_in01 = reg_0899;
    96: op1_10_in01 = imem01_in[27:24];
    97: op1_10_in01 = reg_0180;
    default: op1_10_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv01 = 1;
    7: op1_10_inv01 = 1;
    8: op1_10_inv01 = 1;
    10: op1_10_inv01 = 1;
    16: op1_10_inv01 = 1;
    17: op1_10_inv01 = 1;
    18: op1_10_inv01 = 1;
    20: op1_10_inv01 = 1;
    21: op1_10_inv01 = 1;
    22: op1_10_inv01 = 1;
    24: op1_10_inv01 = 1;
    3: op1_10_inv01 = 1;
    26: op1_10_inv01 = 1;
    28: op1_10_inv01 = 1;
    29: op1_10_inv01 = 1;
    30: op1_10_inv01 = 1;
    31: op1_10_inv01 = 1;
    34: op1_10_inv01 = 1;
    35: op1_10_inv01 = 1;
    37: op1_10_inv01 = 1;
    38: op1_10_inv01 = 1;
    41: op1_10_inv01 = 1;
    42: op1_10_inv01 = 1;
    43: op1_10_inv01 = 1;
    48: op1_10_inv01 = 1;
    49: op1_10_inv01 = 1;
    52: op1_10_inv01 = 1;
    53: op1_10_inv01 = 1;
    54: op1_10_inv01 = 1;
    56: op1_10_inv01 = 1;
    58: op1_10_inv01 = 1;
    59: op1_10_inv01 = 1;
    62: op1_10_inv01 = 1;
    63: op1_10_inv01 = 1;
    64: op1_10_inv01 = 1;
    65: op1_10_inv01 = 1;
    66: op1_10_inv01 = 1;
    68: op1_10_inv01 = 1;
    71: op1_10_inv01 = 1;
    74: op1_10_inv01 = 1;
    75: op1_10_inv01 = 1;
    76: op1_10_inv01 = 1;
    77: op1_10_inv01 = 1;
    78: op1_10_inv01 = 1;
    81: op1_10_inv01 = 1;
    87: op1_10_inv01 = 1;
    92: op1_10_inv01 = 1;
    93: op1_10_inv01 = 1;
    97: op1_10_inv01 = 1;
    default: op1_10_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in02 = reg_0685;
    6: op1_10_in02 = imem00_in[47:44];
    7: op1_10_in02 = reg_0358;
    8: op1_10_in02 = reg_0966;
    9: op1_10_in02 = imem00_in[71:68];
    10: op1_10_in02 = reg_0344;
    11: op1_10_in02 = reg_0647;
    12: op1_10_in02 = reg_1028;
    13: op1_10_in02 = reg_0588;
    14: op1_10_in02 = reg_0048;
    15: op1_10_in02 = reg_0625;
    16: op1_10_in02 = reg_1033;
    17: op1_10_in02 = reg_0977;
    4: op1_10_in02 = imem07_in[71:68];
    18: op1_10_in02 = reg_0116;
    19: op1_10_in02 = imem03_in[107:104];
    63: op1_10_in02 = imem03_in[107:104];
    20: op1_10_in02 = reg_0125;
    21: op1_10_in02 = reg_0067;
    22: op1_10_in02 = reg_0679;
    23: op1_10_in02 = reg_0679;
    24: op1_10_in02 = imem00_in[35:32];
    25: op1_10_in02 = reg_0104;
    3: op1_10_in02 = reg_0175;
    26: op1_10_in02 = imem06_in[115:112];
    27: op1_10_in02 = reg_0090;
    28: op1_10_in02 = imem03_in[79:76];
    29: op1_10_in02 = reg_0299;
    30: op1_10_in02 = reg_0830;
    31: op1_10_in02 = reg_0997;
    2: op1_10_in02 = imem07_in[111:108];
    32: op1_10_in02 = reg_0614;
    33: op1_10_in02 = reg_0434;
    34: op1_10_in02 = imem02_in[7:4];
    77: op1_10_in02 = imem02_in[7:4];
    35: op1_10_in02 = reg_0130;
    36: op1_10_in02 = reg_0141;
    37: op1_10_in02 = imem07_in[119:116];
    38: op1_10_in02 = reg_0154;
    70: op1_10_in02 = reg_0154;
    39: op1_10_in02 = imem00_in[59:56];
    40: op1_10_in02 = reg_0108;
    41: op1_10_in02 = reg_0126;
    42: op1_10_in02 = imem06_in[31:28];
    43: op1_10_in02 = reg_0309;
    44: op1_10_in02 = imem00_in[83:80];
    45: op1_10_in02 = reg_0991;
    46: op1_10_in02 = reg_0957;
    47: op1_10_in02 = imem00_in[39:36];
    76: op1_10_in02 = imem00_in[39:36];
    48: op1_10_in02 = reg_0998;
    49: op1_10_in02 = reg_0950;
    50: op1_10_in02 = reg_0049;
    51: op1_10_in02 = reg_0610;
    52: op1_10_in02 = imem00_in[51:48];
    53: op1_10_in02 = reg_0520;
    54: op1_10_in02 = reg_0514;
    55: op1_10_in02 = reg_0888;
    56: op1_10_in02 = reg_0288;
    57: op1_10_in02 = reg_0078;
    58: op1_10_in02 = reg_0436;
    59: op1_10_in02 = imem06_in[111:108];
    60: op1_10_in02 = reg_0626;
    61: op1_10_in02 = reg_0709;
    62: op1_10_in02 = imem00_in[115:112];
    93: op1_10_in02 = imem00_in[115:112];
    64: op1_10_in02 = reg_0374;
    65: op1_10_in02 = reg_0276;
    66: op1_10_in02 = reg_0945;
    67: op1_10_in02 = reg_0531;
    68: op1_10_in02 = imem00_in[67:64];
    69: op1_10_in02 = reg_0111;
    71: op1_10_in02 = reg_0721;
    72: op1_10_in02 = reg_0233;
    73: op1_10_in02 = reg_0926;
    74: op1_10_in02 = reg_0217;
    85: op1_10_in02 = reg_0217;
    75: op1_10_in02 = reg_0575;
    78: op1_10_in02 = imem02_in[31:28];
    79: op1_10_in02 = imem03_in[115:112];
    80: op1_10_in02 = imem06_in[19:16];
    81: op1_10_in02 = reg_0782;
    82: op1_10_in02 = reg_0269;
    83: op1_10_in02 = imem03_in[39:36];
    84: op1_10_in02 = imem00_in[27:24];
    86: op1_10_in02 = reg_0724;
    87: op1_10_in02 = imem02_in[43:40];
    88: op1_10_in02 = imem05_in[47:44];
    89: op1_10_in02 = imem02_in[59:56];
    90: op1_10_in02 = reg_0058;
    91: op1_10_in02 = reg_0802;
    92: op1_10_in02 = reg_0787;
    94: op1_10_in02 = imem00_in[79:76];
    95: op1_10_in02 = reg_0738;
    96: op1_10_in02 = imem01_in[31:28];
    97: op1_10_in02 = reg_0731;
    default: op1_10_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv02 = 1;
    9: op1_10_inv02 = 1;
    11: op1_10_inv02 = 1;
    12: op1_10_inv02 = 1;
    14: op1_10_inv02 = 1;
    16: op1_10_inv02 = 1;
    4: op1_10_inv02 = 1;
    20: op1_10_inv02 = 1;
    21: op1_10_inv02 = 1;
    22: op1_10_inv02 = 1;
    23: op1_10_inv02 = 1;
    24: op1_10_inv02 = 1;
    3: op1_10_inv02 = 1;
    28: op1_10_inv02 = 1;
    29: op1_10_inv02 = 1;
    30: op1_10_inv02 = 1;
    31: op1_10_inv02 = 1;
    33: op1_10_inv02 = 1;
    34: op1_10_inv02 = 1;
    37: op1_10_inv02 = 1;
    39: op1_10_inv02 = 1;
    40: op1_10_inv02 = 1;
    42: op1_10_inv02 = 1;
    43: op1_10_inv02 = 1;
    45: op1_10_inv02 = 1;
    46: op1_10_inv02 = 1;
    47: op1_10_inv02 = 1;
    55: op1_10_inv02 = 1;
    56: op1_10_inv02 = 1;
    57: op1_10_inv02 = 1;
    58: op1_10_inv02 = 1;
    60: op1_10_inv02 = 1;
    62: op1_10_inv02 = 1;
    63: op1_10_inv02 = 1;
    64: op1_10_inv02 = 1;
    66: op1_10_inv02 = 1;
    68: op1_10_inv02 = 1;
    70: op1_10_inv02 = 1;
    71: op1_10_inv02 = 1;
    73: op1_10_inv02 = 1;
    74: op1_10_inv02 = 1;
    78: op1_10_inv02 = 1;
    80: op1_10_inv02 = 1;
    83: op1_10_inv02 = 1;
    84: op1_10_inv02 = 1;
    85: op1_10_inv02 = 1;
    86: op1_10_inv02 = 1;
    87: op1_10_inv02 = 1;
    88: op1_10_inv02 = 1;
    89: op1_10_inv02 = 1;
    91: op1_10_inv02 = 1;
    92: op1_10_inv02 = 1;
    93: op1_10_inv02 = 1;
    94: op1_10_inv02 = 1;
    96: op1_10_inv02 = 1;
    default: op1_10_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in03 = reg_0689;
    6: op1_10_in03 = imem00_in[51:48];
    47: op1_10_in03 = imem00_in[51:48];
    7: op1_10_in03 = reg_0325;
    8: op1_10_in03 = reg_0972;
    9: op1_10_in03 = imem00_in[75:72];
    10: op1_10_in03 = reg_0381;
    11: op1_10_in03 = reg_0648;
    12: op1_10_in03 = reg_1010;
    13: op1_10_in03 = reg_0590;
    14: op1_10_in03 = imem05_in[11:8];
    15: op1_10_in03 = reg_0630;
    16: op1_10_in03 = reg_1017;
    17: op1_10_in03 = reg_1000;
    4: op1_10_in03 = imem07_in[75:72];
    18: op1_10_in03 = reg_0119;
    19: op1_10_in03 = reg_0569;
    20: op1_10_in03 = reg_0106;
    21: op1_10_in03 = reg_0259;
    22: op1_10_in03 = reg_0691;
    23: op1_10_in03 = reg_0690;
    24: op1_10_in03 = imem00_in[43:40];
    25: op1_10_in03 = reg_0120;
    3: op1_10_in03 = reg_0181;
    26: op1_10_in03 = reg_0614;
    27: op1_10_in03 = imem03_in[47:44];
    28: op1_10_in03 = imem03_in[111:108];
    29: op1_10_in03 = reg_0224;
    30: op1_10_in03 = reg_0500;
    31: op1_10_in03 = imem04_in[15:12];
    32: op1_10_in03 = reg_0607;
    33: op1_10_in03 = reg_0446;
    34: op1_10_in03 = imem02_in[27:24];
    35: op1_10_in03 = imem06_in[11:8];
    36: op1_10_in03 = reg_0137;
    37: op1_10_in03 = reg_0713;
    38: op1_10_in03 = reg_0134;
    39: op1_10_in03 = imem00_in[83:80];
    40: op1_10_in03 = reg_0100;
    41: op1_10_in03 = imem02_in[7:4];
    42: op1_10_in03 = reg_0534;
    43: op1_10_in03 = reg_0626;
    44: op1_10_in03 = imem00_in[103:100];
    45: op1_10_in03 = reg_0978;
    46: op1_10_in03 = reg_0948;
    48: op1_10_in03 = reg_0984;
    49: op1_10_in03 = reg_0964;
    50: op1_10_in03 = reg_0016;
    51: op1_10_in03 = reg_0925;
    52: op1_10_in03 = reg_0695;
    53: op1_10_in03 = reg_1043;
    54: op1_10_in03 = reg_0830;
    55: op1_10_in03 = reg_0931;
    56: op1_10_in03 = reg_0281;
    57: op1_10_in03 = reg_0027;
    58: op1_10_in03 = reg_0094;
    59: op1_10_in03 = reg_0660;
    60: op1_10_in03 = reg_0735;
    61: op1_10_in03 = reg_0718;
    62: op1_10_in03 = imem00_in[119:116];
    63: op1_10_in03 = reg_0681;
    64: op1_10_in03 = reg_0234;
    65: op1_10_in03 = reg_0074;
    66: op1_10_in03 = reg_0896;
    67: op1_10_in03 = imem05_in[31:28];
    68: op1_10_in03 = imem00_in[95:92];
    94: op1_10_in03 = imem00_in[95:92];
    69: op1_10_in03 = reg_0003;
    70: op1_10_in03 = imem06_in[47:44];
    71: op1_10_in03 = reg_0723;
    97: op1_10_in03 = reg_0723;
    72: op1_10_in03 = reg_0551;
    73: op1_10_in03 = reg_0692;
    74: op1_10_in03 = reg_0652;
    75: op1_10_in03 = reg_0303;
    76: op1_10_in03 = reg_0768;
    77: op1_10_in03 = imem02_in[15:12];
    78: op1_10_in03 = imem02_in[35:32];
    79: op1_10_in03 = reg_0620;
    80: op1_10_in03 = imem06_in[39:36];
    81: op1_10_in03 = reg_0566;
    82: op1_10_in03 = reg_0947;
    83: op1_10_in03 = imem03_in[75:72];
    84: op1_10_in03 = imem00_in[35:32];
    85: op1_10_in03 = reg_0141;
    87: op1_10_in03 = imem02_in[75:72];
    88: op1_10_in03 = imem05_in[51:48];
    89: op1_10_in03 = imem02_in[71:68];
    90: op1_10_in03 = reg_0076;
    91: op1_10_in03 = reg_0068;
    92: op1_10_in03 = reg_0440;
    93: op1_10_in03 = reg_0683;
    95: op1_10_in03 = reg_0078;
    96: op1_10_in03 = imem01_in[35:32];
    default: op1_10_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv03 = 1;
    9: op1_10_inv03 = 1;
    10: op1_10_inv03 = 1;
    12: op1_10_inv03 = 1;
    15: op1_10_inv03 = 1;
    17: op1_10_inv03 = 1;
    4: op1_10_inv03 = 1;
    18: op1_10_inv03 = 1;
    19: op1_10_inv03 = 1;
    20: op1_10_inv03 = 1;
    22: op1_10_inv03 = 1;
    24: op1_10_inv03 = 1;
    25: op1_10_inv03 = 1;
    26: op1_10_inv03 = 1;
    27: op1_10_inv03 = 1;
    29: op1_10_inv03 = 1;
    32: op1_10_inv03 = 1;
    37: op1_10_inv03 = 1;
    39: op1_10_inv03 = 1;
    40: op1_10_inv03 = 1;
    41: op1_10_inv03 = 1;
    44: op1_10_inv03 = 1;
    46: op1_10_inv03 = 1;
    48: op1_10_inv03 = 1;
    49: op1_10_inv03 = 1;
    51: op1_10_inv03 = 1;
    53: op1_10_inv03 = 1;
    55: op1_10_inv03 = 1;
    57: op1_10_inv03 = 1;
    66: op1_10_inv03 = 1;
    67: op1_10_inv03 = 1;
    68: op1_10_inv03 = 1;
    71: op1_10_inv03 = 1;
    72: op1_10_inv03 = 1;
    73: op1_10_inv03 = 1;
    74: op1_10_inv03 = 1;
    75: op1_10_inv03 = 1;
    76: op1_10_inv03 = 1;
    77: op1_10_inv03 = 1;
    78: op1_10_inv03 = 1;
    79: op1_10_inv03 = 1;
    80: op1_10_inv03 = 1;
    81: op1_10_inv03 = 1;
    82: op1_10_inv03 = 1;
    87: op1_10_inv03 = 1;
    90: op1_10_inv03 = 1;
    92: op1_10_inv03 = 1;
    96: op1_10_inv03 = 1;
    97: op1_10_inv03 = 1;
    default: op1_10_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in04 = reg_0679;
    6: op1_10_in04 = imem00_in[99:96];
    7: op1_10_in04 = reg_0341;
    8: op1_10_in04 = reg_0960;
    9: op1_10_in04 = imem00_in[123:120];
    10: op1_10_in04 = reg_0372;
    11: op1_10_in04 = reg_0665;
    12: op1_10_in04 = reg_0782;
    13: op1_10_in04 = reg_0391;
    14: op1_10_in04 = imem05_in[15:12];
    15: op1_10_in04 = reg_0618;
    16: op1_10_in04 = reg_0122;
    17: op1_10_in04 = reg_0994;
    4: op1_10_in04 = imem07_in[111:108];
    18: op1_10_in04 = reg_0114;
    19: op1_10_in04 = reg_0369;
    20: op1_10_in04 = reg_0109;
    21: op1_10_in04 = reg_0069;
    22: op1_10_in04 = reg_0680;
    23: op1_10_in04 = reg_0677;
    24: op1_10_in04 = imem00_in[47:44];
    84: op1_10_in04 = imem00_in[47:44];
    25: op1_10_in04 = reg_0106;
    40: op1_10_in04 = reg_0106;
    3: op1_10_in04 = reg_0162;
    26: op1_10_in04 = reg_0625;
    59: op1_10_in04 = reg_0625;
    27: op1_10_in04 = imem03_in[103:100];
    28: op1_10_in04 = imem03_in[123:120];
    29: op1_10_in04 = reg_0555;
    30: op1_10_in04 = reg_0216;
    31: op1_10_in04 = imem04_in[23:20];
    32: op1_10_in04 = reg_0620;
    33: op1_10_in04 = reg_0449;
    34: op1_10_in04 = imem02_in[63:60];
    35: op1_10_in04 = imem06_in[15:12];
    36: op1_10_in04 = reg_0144;
    38: op1_10_in04 = reg_0144;
    37: op1_10_in04 = reg_0711;
    39: op1_10_in04 = imem00_in[87:84];
    41: op1_10_in04 = imem02_in[11:8];
    42: op1_10_in04 = reg_0624;
    43: op1_10_in04 = reg_0531;
    44: op1_10_in04 = imem00_in[127:124];
    45: op1_10_in04 = imem04_in[39:36];
    46: op1_10_in04 = reg_0964;
    47: op1_10_in04 = imem00_in[75:72];
    48: op1_10_in04 = imem04_in[15:12];
    49: op1_10_in04 = reg_0949;
    50: op1_10_in04 = imem03_in[43:40];
    51: op1_10_in04 = reg_0113;
    52: op1_10_in04 = reg_0681;
    53: op1_10_in04 = reg_0227;
    54: op1_10_in04 = reg_0227;
    55: op1_10_in04 = reg_0541;
    56: op1_10_in04 = reg_0078;
    57: op1_10_in04 = reg_0517;
    58: op1_10_in04 = reg_1046;
    60: op1_10_in04 = reg_0692;
    61: op1_10_in04 = reg_0361;
    62: op1_10_in04 = reg_0841;
    63: op1_10_in04 = reg_1007;
    64: op1_10_in04 = reg_0984;
    65: op1_10_in04 = reg_0732;
    66: op1_10_in04 = imem05_in[23:20];
    67: op1_10_in04 = imem05_in[51:48];
    68: op1_10_in04 = reg_0519;
    69: op1_10_in04 = reg_0283;
    70: op1_10_in04 = imem06_in[95:92];
    71: op1_10_in04 = reg_0715;
    72: op1_10_in04 = reg_0998;
    73: op1_10_in04 = reg_0895;
    74: op1_10_in04 = reg_0142;
    75: op1_10_in04 = reg_0744;
    76: op1_10_in04 = reg_0748;
    77: op1_10_in04 = imem02_in[19:16];
    78: op1_10_in04 = imem02_in[87:84];
    79: op1_10_in04 = reg_0756;
    80: op1_10_in04 = imem06_in[51:48];
    81: op1_10_in04 = reg_0716;
    82: op1_10_in04 = reg_0943;
    83: op1_10_in04 = imem03_in[91:88];
    85: op1_10_in04 = reg_0269;
    87: op1_10_in04 = imem02_in[83:80];
    89: op1_10_in04 = imem02_in[83:80];
    88: op1_10_in04 = imem05_in[67:64];
    90: op1_10_in04 = reg_0056;
    91: op1_10_in04 = reg_0015;
    92: op1_10_in04 = reg_0698;
    93: op1_10_in04 = reg_0762;
    94: op1_10_in04 = reg_0684;
    95: op1_10_in04 = reg_0521;
    96: op1_10_in04 = imem01_in[63:60];
    97: op1_10_in04 = reg_0182;
    default: op1_10_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv04 = 1;
    8: op1_10_inv04 = 1;
    9: op1_10_inv04 = 1;
    11: op1_10_inv04 = 1;
    16: op1_10_inv04 = 1;
    17: op1_10_inv04 = 1;
    20: op1_10_inv04 = 1;
    22: op1_10_inv04 = 1;
    23: op1_10_inv04 = 1;
    28: op1_10_inv04 = 1;
    29: op1_10_inv04 = 1;
    30: op1_10_inv04 = 1;
    31: op1_10_inv04 = 1;
    33: op1_10_inv04 = 1;
    36: op1_10_inv04 = 1;
    37: op1_10_inv04 = 1;
    38: op1_10_inv04 = 1;
    41: op1_10_inv04 = 1;
    42: op1_10_inv04 = 1;
    43: op1_10_inv04 = 1;
    44: op1_10_inv04 = 1;
    45: op1_10_inv04 = 1;
    46: op1_10_inv04 = 1;
    50: op1_10_inv04 = 1;
    52: op1_10_inv04 = 1;
    53: op1_10_inv04 = 1;
    55: op1_10_inv04 = 1;
    57: op1_10_inv04 = 1;
    59: op1_10_inv04 = 1;
    60: op1_10_inv04 = 1;
    62: op1_10_inv04 = 1;
    64: op1_10_inv04 = 1;
    68: op1_10_inv04 = 1;
    71: op1_10_inv04 = 1;
    72: op1_10_inv04 = 1;
    73: op1_10_inv04 = 1;
    75: op1_10_inv04 = 1;
    76: op1_10_inv04 = 1;
    77: op1_10_inv04 = 1;
    79: op1_10_inv04 = 1;
    80: op1_10_inv04 = 1;
    81: op1_10_inv04 = 1;
    84: op1_10_inv04 = 1;
    85: op1_10_inv04 = 1;
    88: op1_10_inv04 = 1;
    89: op1_10_inv04 = 1;
    90: op1_10_inv04 = 1;
    91: op1_10_inv04 = 1;
    93: op1_10_inv04 = 1;
    94: op1_10_inv04 = 1;
    96: op1_10_inv04 = 1;
    97: op1_10_inv04 = 1;
    default: op1_10_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in05 = reg_0690;
    52: op1_10_in05 = reg_0690;
    6: op1_10_in05 = reg_0693;
    7: op1_10_in05 = reg_0346;
    8: op1_10_in05 = reg_0256;
    9: op1_10_in05 = reg_0688;
    10: op1_10_in05 = reg_0408;
    11: op1_10_in05 = reg_0341;
    12: op1_10_in05 = imem07_in[15:12];
    13: op1_10_in05 = reg_0360;
    14: op1_10_in05 = imem05_in[51:48];
    15: op1_10_in05 = reg_0632;
    16: op1_10_in05 = reg_0124;
    17: op1_10_in05 = imem04_in[115:112];
    4: op1_10_in05 = imem07_in[119:116];
    18: op1_10_in05 = reg_0106;
    19: op1_10_in05 = reg_0396;
    20: op1_10_in05 = reg_0107;
    25: op1_10_in05 = reg_0107;
    85: op1_10_in05 = reg_0107;
    21: op1_10_in05 = reg_0296;
    91: op1_10_in05 = reg_0296;
    22: op1_10_in05 = reg_0687;
    23: op1_10_in05 = reg_0675;
    24: op1_10_in05 = imem00_in[71:68];
    3: op1_10_in05 = reg_0183;
    26: op1_10_in05 = reg_0613;
    73: op1_10_in05 = reg_0613;
    27: op1_10_in05 = imem03_in[107:104];
    83: op1_10_in05 = imem03_in[107:104];
    28: op1_10_in05 = reg_0984;
    29: op1_10_in05 = reg_0810;
    30: op1_10_in05 = reg_0871;
    31: op1_10_in05 = imem04_in[51:48];
    45: op1_10_in05 = imem04_in[51:48];
    32: op1_10_in05 = reg_0608;
    33: op1_10_in05 = reg_0442;
    34: op1_10_in05 = imem02_in[87:84];
    35: op1_10_in05 = imem06_in[19:16];
    36: op1_10_in05 = reg_0604;
    37: op1_10_in05 = reg_0707;
    38: op1_10_in05 = imem06_in[15:12];
    39: op1_10_in05 = reg_0695;
    47: op1_10_in05 = reg_0695;
    40: op1_10_in05 = reg_0115;
    41: op1_10_in05 = imem02_in[63:60];
    42: op1_10_in05 = reg_0556;
    43: op1_10_in05 = reg_0633;
    44: op1_10_in05 = reg_0682;
    46: op1_10_in05 = reg_0945;
    48: op1_10_in05 = imem04_in[31:28];
    49: op1_10_in05 = reg_0961;
    50: op1_10_in05 = imem03_in[87:84];
    51: op1_10_in05 = reg_0126;
    53: op1_10_in05 = imem01_in[15:12];
    54: op1_10_in05 = reg_0521;
    55: op1_10_in05 = reg_0276;
    56: op1_10_in05 = reg_0485;
    57: op1_10_in05 = reg_0529;
    58: op1_10_in05 = reg_0333;
    59: op1_10_in05 = reg_0262;
    60: op1_10_in05 = reg_0439;
    61: op1_10_in05 = reg_0002;
    62: op1_10_in05 = reg_0768;
    63: op1_10_in05 = reg_0765;
    64: op1_10_in05 = reg_0993;
    65: op1_10_in05 = reg_0065;
    66: op1_10_in05 = imem05_in[43:40];
    67: op1_10_in05 = imem05_in[59:56];
    68: op1_10_in05 = reg_0683;
    69: op1_10_in05 = reg_1033;
    70: op1_10_in05 = reg_1018;
    71: op1_10_in05 = reg_0718;
    72: op1_10_in05 = reg_0991;
    74: op1_10_in05 = reg_0140;
    75: op1_10_in05 = reg_0350;
    76: op1_10_in05 = reg_0684;
    77: op1_10_in05 = imem02_in[79:76];
    78: op1_10_in05 = imem02_in[103:100];
    87: op1_10_in05 = imem02_in[103:100];
    79: op1_10_in05 = reg_0596;
    80: op1_10_in05 = imem06_in[75:72];
    81: op1_10_in05 = reg_0497;
    82: op1_10_in05 = reg_0972;
    84: op1_10_in05 = imem00_in[55:52];
    88: op1_10_in05 = imem05_in[99:96];
    89: op1_10_in05 = imem02_in[111:108];
    90: op1_10_in05 = reg_0068;
    92: op1_10_in05 = reg_0928;
    93: op1_10_in05 = reg_0344;
    94: op1_10_in05 = reg_0760;
    95: op1_10_in05 = reg_0132;
    96: op1_10_in05 = imem01_in[67:64];
    97: op1_10_in05 = reg_0565;
    default: op1_10_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_10_inv05 = 1;
    9: op1_10_inv05 = 1;
    10: op1_10_inv05 = 1;
    14: op1_10_inv05 = 1;
    17: op1_10_inv05 = 1;
    19: op1_10_inv05 = 1;
    22: op1_10_inv05 = 1;
    23: op1_10_inv05 = 1;
    25: op1_10_inv05 = 1;
    26: op1_10_inv05 = 1;
    27: op1_10_inv05 = 1;
    28: op1_10_inv05 = 1;
    29: op1_10_inv05 = 1;
    30: op1_10_inv05 = 1;
    31: op1_10_inv05 = 1;
    32: op1_10_inv05 = 1;
    33: op1_10_inv05 = 1;
    34: op1_10_inv05 = 1;
    35: op1_10_inv05 = 1;
    37: op1_10_inv05 = 1;
    39: op1_10_inv05 = 1;
    41: op1_10_inv05 = 1;
    49: op1_10_inv05 = 1;
    50: op1_10_inv05 = 1;
    51: op1_10_inv05 = 1;
    53: op1_10_inv05 = 1;
    54: op1_10_inv05 = 1;
    55: op1_10_inv05 = 1;
    58: op1_10_inv05 = 1;
    62: op1_10_inv05 = 1;
    69: op1_10_inv05 = 1;
    70: op1_10_inv05 = 1;
    71: op1_10_inv05 = 1;
    73: op1_10_inv05 = 1;
    74: op1_10_inv05 = 1;
    76: op1_10_inv05 = 1;
    77: op1_10_inv05 = 1;
    78: op1_10_inv05 = 1;
    83: op1_10_inv05 = 1;
    90: op1_10_inv05 = 1;
    95: op1_10_inv05 = 1;
    96: op1_10_inv05 = 1;
    97: op1_10_inv05 = 1;
    default: op1_10_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in06 = reg_0691;
    52: op1_10_in06 = reg_0691;
    6: op1_10_in06 = reg_0694;
    7: op1_10_in06 = reg_0324;
    8: op1_10_in06 = reg_0252;
    9: op1_10_in06 = reg_0465;
    23: op1_10_in06 = reg_0465;
    10: op1_10_in06 = reg_0313;
    11: op1_10_in06 = reg_0353;
    12: op1_10_in06 = imem07_in[19:16];
    13: op1_10_in06 = reg_0317;
    14: op1_10_in06 = imem05_in[55:52];
    15: op1_10_in06 = reg_0623;
    16: op1_10_in06 = reg_0125;
    17: op1_10_in06 = imem04_in[119:116];
    4: op1_10_in06 = reg_0447;
    18: op1_10_in06 = reg_0110;
    19: op1_10_in06 = reg_0331;
    20: op1_10_in06 = reg_0127;
    21: op1_10_in06 = reg_0075;
    22: op1_10_in06 = reg_0699;
    24: op1_10_in06 = imem00_in[87:84];
    25: op1_10_in06 = imem02_in[19:16];
    3: op1_10_in06 = reg_0166;
    26: op1_10_in06 = reg_0606;
    27: op1_10_in06 = imem03_in[111:108];
    28: op1_10_in06 = reg_0993;
    29: op1_10_in06 = reg_0274;
    30: op1_10_in06 = reg_0119;
    31: op1_10_in06 = imem04_in[59:56];
    32: op1_10_in06 = reg_0622;
    33: op1_10_in06 = reg_0443;
    34: op1_10_in06 = imem02_in[103:100];
    35: op1_10_in06 = imem06_in[87:84];
    36: op1_10_in06 = reg_0026;
    37: op1_10_in06 = reg_0701;
    38: op1_10_in06 = imem06_in[27:24];
    39: op1_10_in06 = reg_0670;
    40: op1_10_in06 = reg_0107;
    41: op1_10_in06 = imem02_in[107:104];
    87: op1_10_in06 = imem02_in[107:104];
    42: op1_10_in06 = reg_0889;
    43: op1_10_in06 = reg_0008;
    44: op1_10_in06 = reg_0457;
    45: op1_10_in06 = imem04_in[91:88];
    46: op1_10_in06 = reg_0806;
    47: op1_10_in06 = reg_0683;
    48: op1_10_in06 = imem04_in[63:60];
    49: op1_10_in06 = reg_0943;
    50: op1_10_in06 = imem03_in[95:92];
    51: op1_10_in06 = imem02_in[7:4];
    53: op1_10_in06 = imem01_in[27:24];
    54: op1_10_in06 = reg_0354;
    55: op1_10_in06 = reg_0584;
    56: op1_10_in06 = reg_0942;
    57: op1_10_in06 = reg_0756;
    58: op1_10_in06 = reg_0438;
    59: op1_10_in06 = reg_0926;
    60: op1_10_in06 = reg_0781;
    61: op1_10_in06 = reg_0303;
    62: op1_10_in06 = reg_0523;
    63: op1_10_in06 = reg_0833;
    64: op1_10_in06 = reg_0981;
    65: op1_10_in06 = reg_0251;
    66: op1_10_in06 = imem05_in[59:56];
    67: op1_10_in06 = reg_0962;
    68: op1_10_in06 = reg_0668;
    69: op1_10_in06 = reg_0273;
    70: op1_10_in06 = reg_0021;
    71: op1_10_in06 = reg_0805;
    72: op1_10_in06 = reg_0980;
    73: op1_10_in06 = reg_0533;
    74: op1_10_in06 = reg_0057;
    75: op1_10_in06 = reg_0024;
    76: op1_10_in06 = reg_0356;
    77: op1_10_in06 = imem02_in[87:84];
    78: op1_10_in06 = reg_0666;
    79: op1_10_in06 = reg_0991;
    80: op1_10_in06 = reg_0010;
    81: op1_10_in06 = reg_0167;
    82: op1_10_in06 = reg_0707;
    83: op1_10_in06 = reg_0006;
    84: op1_10_in06 = imem00_in[63:60];
    85: op1_10_in06 = reg_0947;
    88: op1_10_in06 = imem05_in[107:104];
    89: op1_10_in06 = reg_0285;
    90: op1_10_in06 = reg_0276;
    91: op1_10_in06 = reg_0809;
    92: op1_10_in06 = reg_0783;
    93: op1_10_in06 = reg_0760;
    94: op1_10_in06 = reg_0030;
    95: op1_10_in06 = reg_0580;
    96: op1_10_in06 = imem01_in[91:88];
    97: op1_10_in06 = reg_0157;
    default: op1_10_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_10_inv06 = 1;
    9: op1_10_inv06 = 1;
    12: op1_10_inv06 = 1;
    13: op1_10_inv06 = 1;
    14: op1_10_inv06 = 1;
    16: op1_10_inv06 = 1;
    18: op1_10_inv06 = 1;
    21: op1_10_inv06 = 1;
    22: op1_10_inv06 = 1;
    24: op1_10_inv06 = 1;
    25: op1_10_inv06 = 1;
    26: op1_10_inv06 = 1;
    27: op1_10_inv06 = 1;
    29: op1_10_inv06 = 1;
    31: op1_10_inv06 = 1;
    32: op1_10_inv06 = 1;
    33: op1_10_inv06 = 1;
    34: op1_10_inv06 = 1;
    36: op1_10_inv06 = 1;
    37: op1_10_inv06 = 1;
    44: op1_10_inv06 = 1;
    45: op1_10_inv06 = 1;
    46: op1_10_inv06 = 1;
    48: op1_10_inv06 = 1;
    49: op1_10_inv06 = 1;
    50: op1_10_inv06 = 1;
    53: op1_10_inv06 = 1;
    56: op1_10_inv06 = 1;
    60: op1_10_inv06 = 1;
    61: op1_10_inv06 = 1;
    63: op1_10_inv06 = 1;
    64: op1_10_inv06 = 1;
    66: op1_10_inv06 = 1;
    67: op1_10_inv06 = 1;
    68: op1_10_inv06 = 1;
    69: op1_10_inv06 = 1;
    72: op1_10_inv06 = 1;
    73: op1_10_inv06 = 1;
    74: op1_10_inv06 = 1;
    75: op1_10_inv06 = 1;
    78: op1_10_inv06 = 1;
    80: op1_10_inv06 = 1;
    82: op1_10_inv06 = 1;
    83: op1_10_inv06 = 1;
    85: op1_10_inv06 = 1;
    89: op1_10_inv06 = 1;
    91: op1_10_inv06 = 1;
    92: op1_10_inv06 = 1;
    default: op1_10_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in07 = reg_0675;
    6: op1_10_in07 = reg_0676;
    7: op1_10_in07 = reg_0335;
    11: op1_10_in07 = reg_0335;
    8: op1_10_in07 = reg_0254;
    9: op1_10_in07 = reg_0453;
    22: op1_10_in07 = reg_0453;
    23: op1_10_in07 = reg_0453;
    10: op1_10_in07 = reg_0375;
    12: op1_10_in07 = imem07_in[31:28];
    13: op1_10_in07 = reg_0361;
    71: op1_10_in07 = reg_0361;
    14: op1_10_in07 = imem05_in[59:56];
    15: op1_10_in07 = reg_0615;
    16: op1_10_in07 = reg_0114;
    17: op1_10_in07 = reg_0530;
    4: op1_10_in07 = reg_0419;
    61: op1_10_in07 = reg_0419;
    18: op1_10_in07 = imem02_in[51:48];
    19: op1_10_in07 = reg_0996;
    20: op1_10_in07 = imem02_in[23:20];
    25: op1_10_in07 = imem02_in[23:20];
    21: op1_10_in07 = reg_0064;
    55: op1_10_in07 = reg_0064;
    24: op1_10_in07 = imem00_in[103:100];
    26: op1_10_in07 = reg_0609;
    27: op1_10_in07 = imem03_in[123:120];
    28: op1_10_in07 = reg_0981;
    29: op1_10_in07 = reg_0544;
    30: op1_10_in07 = reg_0112;
    31: op1_10_in07 = imem04_in[75:72];
    32: op1_10_in07 = reg_0392;
    33: op1_10_in07 = reg_0169;
    34: op1_10_in07 = imem02_in[123:120];
    35: op1_10_in07 = reg_0625;
    36: op1_10_in07 = reg_0612;
    37: op1_10_in07 = reg_0425;
    38: op1_10_in07 = imem06_in[47:44];
    39: op1_10_in07 = reg_0687;
    40: op1_10_in07 = imem02_in[19:16];
    41: op1_10_in07 = imem02_in[127:124];
    42: op1_10_in07 = reg_0344;
    43: op1_10_in07 = reg_0005;
    44: op1_10_in07 = reg_0466;
    45: op1_10_in07 = reg_0277;
    46: op1_10_in07 = reg_0827;
    69: op1_10_in07 = reg_0827;
    47: op1_10_in07 = reg_0696;
    48: op1_10_in07 = imem04_in[71:68];
    49: op1_10_in07 = reg_0256;
    50: op1_10_in07 = imem03_in[103:100];
    51: op1_10_in07 = imem02_in[99:96];
    52: op1_10_in07 = reg_0680;
    93: op1_10_in07 = reg_0680;
    53: op1_10_in07 = imem01_in[83:80];
    54: op1_10_in07 = reg_1051;
    56: op1_10_in07 = imem05_in[15:12];
    57: op1_10_in07 = reg_0864;
    58: op1_10_in07 = reg_0489;
    59: op1_10_in07 = reg_0632;
    60: op1_10_in07 = reg_0008;
    62: op1_10_in07 = reg_0748;
    63: op1_10_in07 = reg_0795;
    64: op1_10_in07 = imem04_in[7:4];
    65: op1_10_in07 = reg_0650;
    66: op1_10_in07 = imem05_in[87:84];
    67: op1_10_in07 = reg_0834;
    68: op1_10_in07 = reg_0454;
    70: op1_10_in07 = reg_0328;
    72: op1_10_in07 = reg_0974;
    73: op1_10_in07 = reg_0439;
    74: op1_10_in07 = reg_0583;
    75: op1_10_in07 = reg_0838;
    76: op1_10_in07 = reg_0469;
    77: op1_10_in07 = imem02_in[119:116];
    78: op1_10_in07 = reg_0637;
    79: op1_10_in07 = reg_0990;
    80: op1_10_in07 = reg_0393;
    81: op1_10_in07 = reg_0822;
    82: op1_10_in07 = reg_0970;
    83: op1_10_in07 = reg_0012;
    84: op1_10_in07 = imem00_in[119:116];
    85: op1_10_in07 = reg_0967;
    87: op1_10_in07 = imem02_in[111:108];
    88: op1_10_in07 = imem05_in[123:120];
    89: op1_10_in07 = reg_0090;
    90: op1_10_in07 = reg_0296;
    91: op1_10_in07 = reg_0444;
    92: op1_10_in07 = reg_0011;
    94: op1_10_in07 = reg_0580;
    95: op1_10_in07 = reg_0699;
    96: op1_10_in07 = imem01_in[95:92];
    default: op1_10_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv07 = 1;
    6: op1_10_inv07 = 1;
    10: op1_10_inv07 = 1;
    12: op1_10_inv07 = 1;
    13: op1_10_inv07 = 1;
    14: op1_10_inv07 = 1;
    16: op1_10_inv07 = 1;
    17: op1_10_inv07 = 1;
    4: op1_10_inv07 = 1;
    18: op1_10_inv07 = 1;
    20: op1_10_inv07 = 1;
    21: op1_10_inv07 = 1;
    26: op1_10_inv07 = 1;
    27: op1_10_inv07 = 1;
    30: op1_10_inv07 = 1;
    31: op1_10_inv07 = 1;
    32: op1_10_inv07 = 1;
    34: op1_10_inv07 = 1;
    36: op1_10_inv07 = 1;
    38: op1_10_inv07 = 1;
    40: op1_10_inv07 = 1;
    41: op1_10_inv07 = 1;
    45: op1_10_inv07 = 1;
    46: op1_10_inv07 = 1;
    48: op1_10_inv07 = 1;
    50: op1_10_inv07 = 1;
    51: op1_10_inv07 = 1;
    52: op1_10_inv07 = 1;
    53: op1_10_inv07 = 1;
    54: op1_10_inv07 = 1;
    55: op1_10_inv07 = 1;
    59: op1_10_inv07 = 1;
    60: op1_10_inv07 = 1;
    61: op1_10_inv07 = 1;
    62: op1_10_inv07 = 1;
    64: op1_10_inv07 = 1;
    68: op1_10_inv07 = 1;
    71: op1_10_inv07 = 1;
    74: op1_10_inv07 = 1;
    76: op1_10_inv07 = 1;
    77: op1_10_inv07 = 1;
    78: op1_10_inv07 = 1;
    80: op1_10_inv07 = 1;
    82: op1_10_inv07 = 1;
    84: op1_10_inv07 = 1;
    85: op1_10_inv07 = 1;
    88: op1_10_inv07 = 1;
    89: op1_10_inv07 = 1;
    90: op1_10_inv07 = 1;
    91: op1_10_inv07 = 1;
    92: op1_10_inv07 = 1;
    93: op1_10_inv07 = 1;
    default: op1_10_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in08 = reg_0680;
    6: op1_10_in08 = reg_0671;
    7: op1_10_in08 = reg_0347;
    8: op1_10_in08 = reg_0255;
    9: op1_10_in08 = reg_0460;
    10: op1_10_in08 = reg_0382;
    11: op1_10_in08 = reg_0328;
    12: op1_10_in08 = imem07_in[43:40];
    13: op1_10_in08 = reg_0396;
    14: op1_10_in08 = imem05_in[103:100];
    15: op1_10_in08 = reg_0405;
    16: op1_10_in08 = imem02_in[15:12];
    17: op1_10_in08 = reg_0534;
    4: op1_10_in08 = reg_0443;
    18: op1_10_in08 = imem02_in[71:68];
    19: op1_10_in08 = reg_0978;
    20: op1_10_in08 = imem02_in[47:44];
    21: op1_10_in08 = reg_0278;
    22: op1_10_in08 = reg_0454;
    23: op1_10_in08 = reg_0457;
    94: op1_10_in08 = reg_0457;
    24: op1_10_in08 = reg_0672;
    25: op1_10_in08 = imem02_in[115:112];
    26: op1_10_in08 = reg_0611;
    27: op1_10_in08 = reg_0572;
    28: op1_10_in08 = reg_0977;
    29: op1_10_in08 = reg_0905;
    30: op1_10_in08 = reg_0106;
    31: op1_10_in08 = reg_0536;
    32: op1_10_in08 = reg_0390;
    33: op1_10_in08 = reg_0177;
    34: op1_10_in08 = reg_0645;
    35: op1_10_in08 = reg_0629;
    36: op1_10_in08 = reg_0521;
    37: op1_10_in08 = reg_0433;
    38: op1_10_in08 = imem06_in[67:64];
    39: op1_10_in08 = reg_0450;
    68: op1_10_in08 = reg_0450;
    40: op1_10_in08 = imem02_in[51:48];
    41: op1_10_in08 = reg_0664;
    42: op1_10_in08 = reg_0392;
    43: op1_10_in08 = reg_0425;
    44: op1_10_in08 = reg_0472;
    45: op1_10_in08 = reg_1020;
    46: op1_10_in08 = reg_0254;
    47: op1_10_in08 = reg_0676;
    48: op1_10_in08 = imem04_in[79:76];
    49: op1_10_in08 = reg_0825;
    50: op1_10_in08 = imem03_in[111:108];
    51: op1_10_in08 = reg_0642;
    52: op1_10_in08 = reg_0453;
    93: op1_10_in08 = reg_0453;
    53: op1_10_in08 = imem02_in[19:16];
    54: op1_10_in08 = reg_0116;
    55: op1_10_in08 = reg_0284;
    56: op1_10_in08 = imem05_in[31:28];
    57: op1_10_in08 = reg_0031;
    58: op1_10_in08 = reg_0497;
    59: op1_10_in08 = reg_0222;
    60: op1_10_in08 = reg_0380;
    61: op1_10_in08 = reg_0502;
    62: op1_10_in08 = reg_0684;
    63: op1_10_in08 = reg_0373;
    64: op1_10_in08 = imem04_in[11:8];
    65: op1_10_in08 = reg_0971;
    66: op1_10_in08 = reg_0132;
    67: op1_10_in08 = reg_0022;
    69: op1_10_in08 = reg_0115;
    70: op1_10_in08 = reg_0889;
    71: op1_10_in08 = reg_0422;
    72: op1_10_in08 = reg_0988;
    73: op1_10_in08 = reg_0695;
    74: op1_10_in08 = reg_0020;
    75: op1_10_in08 = reg_0174;
    76: op1_10_in08 = reg_0481;
    77: op1_10_in08 = imem02_in[123:120];
    87: op1_10_in08 = imem02_in[123:120];
    78: op1_10_in08 = reg_0765;
    79: op1_10_in08 = imem04_in[23:20];
    80: op1_10_in08 = reg_0262;
    81: op1_10_in08 = reg_0705;
    82: op1_10_in08 = reg_0145;
    83: op1_10_in08 = reg_0760;
    84: op1_10_in08 = reg_0682;
    85: op1_10_in08 = reg_0153;
    88: op1_10_in08 = reg_0136;
    89: op1_10_in08 = reg_0091;
    90: op1_10_in08 = reg_0732;
    91: op1_10_in08 = reg_0065;
    92: op1_10_in08 = reg_0169;
    95: op1_10_in08 = reg_0464;
    96: op1_10_in08 = imem01_in[111:108];
    default: op1_10_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_10_inv08 = 1;
    9: op1_10_inv08 = 1;
    10: op1_10_inv08 = 1;
    12: op1_10_inv08 = 1;
    13: op1_10_inv08 = 1;
    14: op1_10_inv08 = 1;
    17: op1_10_inv08 = 1;
    4: op1_10_inv08 = 1;
    19: op1_10_inv08 = 1;
    22: op1_10_inv08 = 1;
    24: op1_10_inv08 = 1;
    30: op1_10_inv08 = 1;
    31: op1_10_inv08 = 1;
    32: op1_10_inv08 = 1;
    35: op1_10_inv08 = 1;
    37: op1_10_inv08 = 1;
    40: op1_10_inv08 = 1;
    42: op1_10_inv08 = 1;
    45: op1_10_inv08 = 1;
    48: op1_10_inv08 = 1;
    49: op1_10_inv08 = 1;
    50: op1_10_inv08 = 1;
    57: op1_10_inv08 = 1;
    59: op1_10_inv08 = 1;
    60: op1_10_inv08 = 1;
    61: op1_10_inv08 = 1;
    62: op1_10_inv08 = 1;
    64: op1_10_inv08 = 1;
    65: op1_10_inv08 = 1;
    70: op1_10_inv08 = 1;
    71: op1_10_inv08 = 1;
    73: op1_10_inv08 = 1;
    78: op1_10_inv08 = 1;
    79: op1_10_inv08 = 1;
    80: op1_10_inv08 = 1;
    82: op1_10_inv08 = 1;
    83: op1_10_inv08 = 1;
    85: op1_10_inv08 = 1;
    88: op1_10_inv08 = 1;
    89: op1_10_inv08 = 1;
    90: op1_10_inv08 = 1;
    93: op1_10_inv08 = 1;
    95: op1_10_inv08 = 1;
    default: op1_10_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in09 = reg_0451;
    6: op1_10_in09 = reg_0465;
    7: op1_10_in09 = imem03_in[35:32];
    8: op1_10_in09 = reg_0263;
    9: op1_10_in09 = reg_0480;
    10: op1_10_in09 = reg_0404;
    11: op1_10_in09 = reg_0097;
    12: op1_10_in09 = imem07_in[91:88];
    13: op1_10_in09 = reg_0985;
    14: op1_10_in09 = imem05_in[107:104];
    15: op1_10_in09 = reg_1011;
    16: op1_10_in09 = imem02_in[87:84];
    17: op1_10_in09 = reg_0537;
    4: op1_10_in09 = reg_0437;
    18: op1_10_in09 = imem02_in[115:112];
    20: op1_10_in09 = imem02_in[115:112];
    19: op1_10_in09 = reg_0999;
    21: op1_10_in09 = reg_0059;
    22: op1_10_in09 = reg_0469;
    23: op1_10_in09 = reg_0476;
    24: op1_10_in09 = reg_0670;
    84: op1_10_in09 = reg_0670;
    25: op1_10_in09 = reg_0664;
    26: op1_10_in09 = reg_0577;
    27: op1_10_in09 = reg_0594;
    60: op1_10_in09 = reg_0594;
    28: op1_10_in09 = reg_0983;
    29: op1_10_in09 = reg_0226;
    30: op1_10_in09 = reg_0115;
    31: op1_10_in09 = reg_0301;
    32: op1_10_in09 = imem06_in[27:24];
    33: op1_10_in09 = reg_0157;
    34: op1_10_in09 = reg_0654;
    35: op1_10_in09 = reg_0624;
    70: op1_10_in09 = reg_0624;
    36: op1_10_in09 = reg_0915;
    37: op1_10_in09 = reg_0439;
    38: op1_10_in09 = imem06_in[87:84];
    39: op1_10_in09 = reg_0455;
    68: op1_10_in09 = reg_0455;
    40: op1_10_in09 = imem02_in[63:60];
    41: op1_10_in09 = reg_0661;
    42: op1_10_in09 = reg_0383;
    43: op1_10_in09 = reg_0289;
    44: op1_10_in09 = reg_0468;
    45: op1_10_in09 = reg_0932;
    46: op1_10_in09 = reg_0831;
    47: op1_10_in09 = reg_0688;
    48: op1_10_in09 = imem04_in[83:80];
    49: op1_10_in09 = reg_0254;
    50: op1_10_in09 = imem03_in[127:124];
    51: op1_10_in09 = reg_0643;
    52: op1_10_in09 = reg_0470;
    53: op1_10_in09 = imem02_in[55:52];
    54: op1_10_in09 = imem02_in[3:0];
    55: op1_10_in09 = reg_0816;
    56: op1_10_in09 = imem05_in[123:120];
    57: op1_10_in09 = reg_0882;
    58: op1_10_in09 = reg_0148;
    66: op1_10_in09 = reg_0148;
    59: op1_10_in09 = reg_0630;
    61: op1_10_in09 = reg_0431;
    62: op1_10_in09 = reg_0499;
    63: op1_10_in09 = reg_0509;
    64: op1_10_in09 = imem04_in[15:12];
    65: op1_10_in09 = reg_0689;
    67: op1_10_in09 = reg_0835;
    69: op1_10_in09 = reg_0110;
    71: op1_10_in09 = reg_0744;
    72: op1_10_in09 = imem04_in[3:0];
    73: op1_10_in09 = reg_0370;
    74: op1_10_in09 = reg_0603;
    75: op1_10_in09 = reg_0182;
    76: op1_10_in09 = reg_0473;
    77: op1_10_in09 = reg_0750;
    78: op1_10_in09 = reg_0418;
    79: op1_10_in09 = imem04_in[67:64];
    80: op1_10_in09 = reg_0817;
    81: op1_10_in09 = reg_0123;
    82: op1_10_in09 = reg_0508;
    83: op1_10_in09 = reg_0346;
    85: op1_10_in09 = reg_1046;
    87: op1_10_in09 = reg_0334;
    88: op1_10_in09 = reg_0652;
    89: op1_10_in09 = reg_0765;
    90: op1_10_in09 = reg_0517;
    91: op1_10_in09 = reg_0517;
    92: op1_10_in09 = reg_0124;
    93: op1_10_in09 = reg_0454;
    94: op1_10_in09 = reg_0466;
    95: op1_10_in09 = reg_0461;
    96: op1_10_in09 = imem01_in[119:116];
    default: op1_10_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv09 = 1;
    13: op1_10_inv09 = 1;
    16: op1_10_inv09 = 1;
    18: op1_10_inv09 = 1;
    21: op1_10_inv09 = 1;
    25: op1_10_inv09 = 1;
    27: op1_10_inv09 = 1;
    28: op1_10_inv09 = 1;
    29: op1_10_inv09 = 1;
    30: op1_10_inv09 = 1;
    31: op1_10_inv09 = 1;
    33: op1_10_inv09 = 1;
    34: op1_10_inv09 = 1;
    35: op1_10_inv09 = 1;
    36: op1_10_inv09 = 1;
    39: op1_10_inv09 = 1;
    40: op1_10_inv09 = 1;
    43: op1_10_inv09 = 1;
    44: op1_10_inv09 = 1;
    45: op1_10_inv09 = 1;
    47: op1_10_inv09 = 1;
    48: op1_10_inv09 = 1;
    49: op1_10_inv09 = 1;
    50: op1_10_inv09 = 1;
    53: op1_10_inv09 = 1;
    54: op1_10_inv09 = 1;
    56: op1_10_inv09 = 1;
    57: op1_10_inv09 = 1;
    58: op1_10_inv09 = 1;
    59: op1_10_inv09 = 1;
    60: op1_10_inv09 = 1;
    62: op1_10_inv09 = 1;
    63: op1_10_inv09 = 1;
    66: op1_10_inv09 = 1;
    67: op1_10_inv09 = 1;
    68: op1_10_inv09 = 1;
    69: op1_10_inv09 = 1;
    70: op1_10_inv09 = 1;
    73: op1_10_inv09 = 1;
    76: op1_10_inv09 = 1;
    77: op1_10_inv09 = 1;
    81: op1_10_inv09 = 1;
    83: op1_10_inv09 = 1;
    85: op1_10_inv09 = 1;
    88: op1_10_inv09 = 1;
    90: op1_10_inv09 = 1;
    92: op1_10_inv09 = 1;
    93: op1_10_inv09 = 1;
    94: op1_10_inv09 = 1;
    96: op1_10_inv09 = 1;
    default: op1_10_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in10 = reg_0473;
    6: op1_10_in10 = reg_0457;
    7: op1_10_in10 = imem03_in[47:44];
    8: op1_10_in10 = reg_0154;
    9: op1_10_in10 = reg_0456;
    52: op1_10_in10 = reg_0456;
    10: op1_10_in10 = reg_0406;
    11: op1_10_in10 = reg_0051;
    12: op1_10_in10 = imem07_in[95:92];
    13: op1_10_in10 = reg_0995;
    14: op1_10_in10 = imem05_in[123:120];
    15: op1_10_in10 = imem07_in[3:0];
    16: op1_10_in10 = reg_0642;
    17: op1_10_in10 = reg_0541;
    4: op1_10_in10 = reg_0435;
    18: op1_10_in10 = imem02_in[127:124];
    20: op1_10_in10 = imem02_in[127:124];
    19: op1_10_in10 = reg_0974;
    21: op1_10_in10 = reg_0525;
    22: op1_10_in10 = reg_0480;
    23: op1_10_in10 = reg_0466;
    24: op1_10_in10 = reg_0679;
    25: op1_10_in10 = reg_0647;
    88: op1_10_in10 = reg_0647;
    26: op1_10_in10 = reg_0618;
    27: op1_10_in10 = reg_0578;
    28: op1_10_in10 = reg_0997;
    29: op1_10_in10 = reg_0230;
    30: op1_10_in10 = reg_0110;
    31: op1_10_in10 = reg_0912;
    32: op1_10_in10 = imem06_in[35:32];
    33: op1_10_in10 = reg_0158;
    34: op1_10_in10 = reg_0660;
    35: op1_10_in10 = reg_0620;
    36: op1_10_in10 = reg_0036;
    37: op1_10_in10 = reg_0449;
    38: op1_10_in10 = imem06_in[107:104];
    39: op1_10_in10 = reg_0469;
    40: op1_10_in10 = imem02_in[79:76];
    41: op1_10_in10 = reg_0639;
    42: op1_10_in10 = reg_0399;
    43: op1_10_in10 = reg_0866;
    44: op1_10_in10 = reg_0214;
    45: op1_10_in10 = reg_0050;
    46: op1_10_in10 = reg_0489;
    47: op1_10_in10 = reg_0673;
    48: op1_10_in10 = imem04_in[107:104];
    49: op1_10_in10 = reg_0831;
    50: op1_10_in10 = reg_0535;
    51: op1_10_in10 = reg_0636;
    53: op1_10_in10 = imem02_in[67:64];
    54: op1_10_in10 = imem02_in[111:108];
    55: op1_10_in10 = reg_0864;
    56: op1_10_in10 = reg_0032;
    57: op1_10_in10 = imem05_in[31:28];
    58: op1_10_in10 = reg_0149;
    59: op1_10_in10 = reg_0241;
    60: op1_10_in10 = reg_0596;
    61: op1_10_in10 = reg_0159;
    62: op1_10_in10 = reg_0069;
    63: op1_10_in10 = reg_0377;
    64: op1_10_in10 = imem04_in[23:20];
    65: op1_10_in10 = reg_0497;
    66: op1_10_in10 = reg_0133;
    67: op1_10_in10 = reg_0800;
    68: op1_10_in10 = reg_0467;
    69: op1_10_in10 = imem02_in[43:40];
    70: op1_10_in10 = reg_0617;
    71: op1_10_in10 = reg_0641;
    72: op1_10_in10 = imem04_in[7:4];
    73: op1_10_in10 = reg_0612;
    74: op1_10_in10 = reg_0436;
    75: op1_10_in10 = reg_0177;
    76: op1_10_in10 = reg_0471;
    77: op1_10_in10 = reg_0666;
    78: op1_10_in10 = reg_0358;
    79: op1_10_in10 = imem04_in[71:68];
    80: op1_10_in10 = reg_1011;
    81: op1_10_in10 = reg_0728;
    82: op1_10_in10 = imem06_in[55:52];
    83: op1_10_in10 = reg_0240;
    84: op1_10_in10 = reg_0883;
    85: op1_10_in10 = reg_0736;
    87: op1_10_in10 = reg_0543;
    89: op1_10_in10 = reg_0394;
    90: op1_10_in10 = reg_0495;
    91: op1_10_in10 = reg_0108;
    92: op1_10_in10 = imem07_in[75:72];
    93: op1_10_in10 = reg_0461;
    94: op1_10_in10 = reg_0472;
    95: op1_10_in10 = reg_0460;
    96: op1_10_in10 = reg_0235;
    default: op1_10_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_10_inv10 = 1;
    13: op1_10_inv10 = 1;
    17: op1_10_inv10 = 1;
    4: op1_10_inv10 = 1;
    21: op1_10_inv10 = 1;
    24: op1_10_inv10 = 1;
    26: op1_10_inv10 = 1;
    28: op1_10_inv10 = 1;
    32: op1_10_inv10 = 1;
    33: op1_10_inv10 = 1;
    35: op1_10_inv10 = 1;
    37: op1_10_inv10 = 1;
    44: op1_10_inv10 = 1;
    45: op1_10_inv10 = 1;
    46: op1_10_inv10 = 1;
    50: op1_10_inv10 = 1;
    51: op1_10_inv10 = 1;
    53: op1_10_inv10 = 1;
    54: op1_10_inv10 = 1;
    55: op1_10_inv10 = 1;
    56: op1_10_inv10 = 1;
    58: op1_10_inv10 = 1;
    59: op1_10_inv10 = 1;
    61: op1_10_inv10 = 1;
    65: op1_10_inv10 = 1;
    68: op1_10_inv10 = 1;
    69: op1_10_inv10 = 1;
    70: op1_10_inv10 = 1;
    74: op1_10_inv10 = 1;
    75: op1_10_inv10 = 1;
    79: op1_10_inv10 = 1;
    80: op1_10_inv10 = 1;
    81: op1_10_inv10 = 1;
    82: op1_10_inv10 = 1;
    83: op1_10_inv10 = 1;
    90: op1_10_inv10 = 1;
    93: op1_10_inv10 = 1;
    94: op1_10_inv10 = 1;
    95: op1_10_inv10 = 1;
    default: op1_10_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in11 = reg_0459;
    76: op1_10_in11 = reg_0459;
    6: op1_10_in11 = reg_0469;
    7: op1_10_in11 = imem03_in[79:76];
    8: op1_10_in11 = reg_0140;
    9: op1_10_in11 = reg_0209;
    10: op1_10_in11 = reg_0367;
    11: op1_10_in11 = reg_0094;
    12: op1_10_in11 = imem07_in[103:100];
    13: op1_10_in11 = reg_0996;
    14: op1_10_in11 = reg_0954;
    67: op1_10_in11 = reg_0954;
    15: op1_10_in11 = imem07_in[7:4];
    16: op1_10_in11 = reg_0650;
    17: op1_10_in11 = reg_0300;
    4: op1_10_in11 = reg_0174;
    18: op1_10_in11 = reg_0658;
    19: op1_10_in11 = reg_0997;
    20: op1_10_in11 = reg_0645;
    21: op1_10_in11 = reg_0054;
    22: op1_10_in11 = reg_0473;
    39: op1_10_in11 = reg_0473;
    95: op1_10_in11 = reg_0473;
    23: op1_10_in11 = reg_0187;
    24: op1_10_in11 = reg_0673;
    25: op1_10_in11 = reg_0352;
    26: op1_10_in11 = reg_0408;
    27: op1_10_in11 = reg_0393;
    28: op1_10_in11 = imem04_in[87:84];
    29: op1_10_in11 = reg_1033;
    30: op1_10_in11 = imem02_in[3:0];
    31: op1_10_in11 = reg_1005;
    32: op1_10_in11 = imem06_in[67:64];
    34: op1_10_in11 = reg_0640;
    35: op1_10_in11 = reg_0632;
    36: op1_10_in11 = reg_0782;
    37: op1_10_in11 = reg_0427;
    38: op1_10_in11 = reg_0372;
    40: op1_10_in11 = imem02_in[111:108];
    41: op1_10_in11 = reg_0649;
    42: op1_10_in11 = reg_0222;
    96: op1_10_in11 = reg_0222;
    43: op1_10_in11 = reg_0636;
    44: op1_10_in11 = reg_0198;
    45: op1_10_in11 = reg_0524;
    46: op1_10_in11 = reg_0497;
    47: op1_10_in11 = reg_0699;
    48: op1_10_in11 = imem04_in[111:108];
    49: op1_10_in11 = reg_0148;
    50: op1_10_in11 = reg_1049;
    51: op1_10_in11 = reg_0863;
    70: op1_10_in11 = reg_0863;
    52: op1_10_in11 = reg_0478;
    53: op1_10_in11 = imem02_in[71:68];
    54: op1_10_in11 = reg_0642;
    55: op1_10_in11 = reg_0882;
    56: op1_10_in11 = reg_0488;
    57: op1_10_in11 = imem05_in[83:80];
    58: op1_10_in11 = reg_0135;
    59: op1_10_in11 = reg_0596;
    60: op1_10_in11 = reg_0609;
    62: op1_10_in11 = reg_0687;
    63: op1_10_in11 = reg_0985;
    64: op1_10_in11 = imem04_in[39:36];
    65: op1_10_in11 = imem05_in[15:12];
    66: op1_10_in11 = reg_0142;
    68: op1_10_in11 = reg_0468;
    94: op1_10_in11 = reg_0468;
    69: op1_10_in11 = imem02_in[47:44];
    71: op1_10_in11 = reg_0532;
    72: op1_10_in11 = imem04_in[23:20];
    73: op1_10_in11 = reg_0383;
    74: op1_10_in11 = reg_0947;
    75: op1_10_in11 = reg_0173;
    77: op1_10_in11 = reg_0803;
    78: op1_10_in11 = reg_0329;
    79: op1_10_in11 = imem04_in[103:100];
    80: op1_10_in11 = reg_0613;
    81: op1_10_in11 = reg_0569;
    82: op1_10_in11 = imem06_in[59:56];
    83: op1_10_in11 = reg_0312;
    84: op1_10_in11 = reg_0356;
    85: op1_10_in11 = reg_0780;
    87: op1_10_in11 = reg_0483;
    88: op1_10_in11 = reg_0448;
    89: op1_10_in11 = reg_0248;
    90: op1_10_in11 = reg_0108;
    91: op1_10_in11 = imem05_in[19:16];
    92: op1_10_in11 = imem07_in[87:84];
    93: op1_10_in11 = reg_0477;
    default: op1_10_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv11 = 1;
    8: op1_10_inv11 = 1;
    13: op1_10_inv11 = 1;
    15: op1_10_inv11 = 1;
    16: op1_10_inv11 = 1;
    17: op1_10_inv11 = 1;
    4: op1_10_inv11 = 1;
    18: op1_10_inv11 = 1;
    20: op1_10_inv11 = 1;
    26: op1_10_inv11 = 1;
    27: op1_10_inv11 = 1;
    28: op1_10_inv11 = 1;
    29: op1_10_inv11 = 1;
    30: op1_10_inv11 = 1;
    31: op1_10_inv11 = 1;
    32: op1_10_inv11 = 1;
    35: op1_10_inv11 = 1;
    37: op1_10_inv11 = 1;
    38: op1_10_inv11 = 1;
    39: op1_10_inv11 = 1;
    45: op1_10_inv11 = 1;
    46: op1_10_inv11 = 1;
    47: op1_10_inv11 = 1;
    50: op1_10_inv11 = 1;
    51: op1_10_inv11 = 1;
    56: op1_10_inv11 = 1;
    60: op1_10_inv11 = 1;
    62: op1_10_inv11 = 1;
    64: op1_10_inv11 = 1;
    65: op1_10_inv11 = 1;
    67: op1_10_inv11 = 1;
    68: op1_10_inv11 = 1;
    71: op1_10_inv11 = 1;
    75: op1_10_inv11 = 1;
    76: op1_10_inv11 = 1;
    77: op1_10_inv11 = 1;
    78: op1_10_inv11 = 1;
    81: op1_10_inv11 = 1;
    83: op1_10_inv11 = 1;
    85: op1_10_inv11 = 1;
    88: op1_10_inv11 = 1;
    89: op1_10_inv11 = 1;
    93: op1_10_inv11 = 1;
    95: op1_10_inv11 = 1;
    default: op1_10_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in12 = reg_0452;
    6: op1_10_in12 = reg_0476;
    7: op1_10_in12 = reg_0572;
    8: op1_10_in12 = reg_0134;
    9: op1_10_in12 = reg_0205;
    10: op1_10_in12 = reg_0380;
    11: op1_10_in12 = reg_0093;
    12: op1_10_in12 = imem07_in[123:120];
    13: op1_10_in12 = reg_0993;
    14: op1_10_in12 = reg_0947;
    15: op1_10_in12 = imem07_in[15:12];
    16: op1_10_in12 = reg_0643;
    17: op1_10_in12 = reg_0299;
    4: op1_10_in12 = reg_0179;
    18: op1_10_in12 = reg_0653;
    19: op1_10_in12 = reg_0994;
    20: op1_10_in12 = reg_0661;
    21: op1_10_in12 = reg_0736;
    22: op1_10_in12 = reg_0470;
    23: op1_10_in12 = reg_0194;
    24: op1_10_in12 = reg_0669;
    25: op1_10_in12 = reg_0341;
    26: op1_10_in12 = reg_0386;
    27: op1_10_in12 = imem04_in[3:0];
    28: op1_10_in12 = imem04_in[103:100];
    29: op1_10_in12 = reg_0830;
    30: op1_10_in12 = imem02_in[23:20];
    31: op1_10_in12 = reg_0537;
    32: op1_10_in12 = imem06_in[71:68];
    34: op1_10_in12 = reg_0638;
    35: op1_10_in12 = reg_0627;
    36: op1_10_in12 = reg_0745;
    37: op1_10_in12 = reg_0438;
    38: op1_10_in12 = reg_0593;
    39: op1_10_in12 = reg_0474;
    95: op1_10_in12 = reg_0474;
    40: op1_10_in12 = imem02_in[119:116];
    41: op1_10_in12 = reg_0916;
    42: op1_10_in12 = reg_0917;
    43: op1_10_in12 = reg_0709;
    44: op1_10_in12 = reg_0197;
    45: op1_10_in12 = reg_0067;
    46: op1_10_in12 = reg_0136;
    47: op1_10_in12 = reg_0475;
    48: op1_10_in12 = reg_0301;
    49: op1_10_in12 = reg_0145;
    50: op1_10_in12 = reg_0358;
    51: op1_10_in12 = reg_0318;
    52: op1_10_in12 = reg_0208;
    53: op1_10_in12 = imem02_in[91:88];
    54: op1_10_in12 = reg_0650;
    55: op1_10_in12 = imem05_in[3:0];
    56: op1_10_in12 = reg_0435;
    57: op1_10_in12 = imem05_in[115:112];
    58: op1_10_in12 = reg_0152;
    59: op1_10_in12 = reg_0633;
    60: op1_10_in12 = reg_0029;
    62: op1_10_in12 = reg_0749;
    63: op1_10_in12 = reg_0997;
    64: op1_10_in12 = imem04_in[71:68];
    65: op1_10_in12 = imem05_in[39:36];
    66: op1_10_in12 = imem06_in[3:0];
    67: op1_10_in12 = reg_0969;
    68: op1_10_in12 = reg_0210;
    76: op1_10_in12 = reg_0210;
    69: op1_10_in12 = imem02_in[79:76];
    70: op1_10_in12 = reg_0804;
    71: op1_10_in12 = reg_0350;
    72: op1_10_in12 = imem04_in[31:28];
    73: op1_10_in12 = reg_0403;
    74: op1_10_in12 = imem05_in[19:16];
    77: op1_10_in12 = reg_0096;
    78: op1_10_in12 = reg_0423;
    79: op1_10_in12 = imem04_in[107:104];
    80: op1_10_in12 = reg_0439;
    81: op1_10_in12 = reg_0923;
    82: op1_10_in12 = imem06_in[83:80];
    83: op1_10_in12 = reg_0385;
    84: op1_10_in12 = reg_0668;
    85: op1_10_in12 = reg_0486;
    87: op1_10_in12 = reg_0887;
    88: op1_10_in12 = reg_0675;
    89: op1_10_in12 = reg_0608;
    90: op1_10_in12 = reg_0251;
    91: op1_10_in12 = imem05_in[35:32];
    92: op1_10_in12 = imem07_in[115:112];
    93: op1_10_in12 = reg_0462;
    94: op1_10_in12 = reg_0479;
    96: op1_10_in12 = reg_0120;
    default: op1_10_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv12 = 1;
    7: op1_10_inv12 = 1;
    8: op1_10_inv12 = 1;
    12: op1_10_inv12 = 1;
    13: op1_10_inv12 = 1;
    15: op1_10_inv12 = 1;
    16: op1_10_inv12 = 1;
    21: op1_10_inv12 = 1;
    23: op1_10_inv12 = 1;
    26: op1_10_inv12 = 1;
    27: op1_10_inv12 = 1;
    29: op1_10_inv12 = 1;
    32: op1_10_inv12 = 1;
    37: op1_10_inv12 = 1;
    41: op1_10_inv12 = 1;
    42: op1_10_inv12 = 1;
    43: op1_10_inv12 = 1;
    44: op1_10_inv12 = 1;
    51: op1_10_inv12 = 1;
    54: op1_10_inv12 = 1;
    58: op1_10_inv12 = 1;
    65: op1_10_inv12 = 1;
    67: op1_10_inv12 = 1;
    69: op1_10_inv12 = 1;
    72: op1_10_inv12 = 1;
    74: op1_10_inv12 = 1;
    78: op1_10_inv12 = 1;
    81: op1_10_inv12 = 1;
    85: op1_10_inv12 = 1;
    88: op1_10_inv12 = 1;
    90: op1_10_inv12 = 1;
    94: op1_10_inv12 = 1;
    96: op1_10_inv12 = 1;
    default: op1_10_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in13 = reg_0456;
    94: op1_10_in13 = reg_0456;
    6: op1_10_in13 = reg_0466;
    7: op1_10_in13 = reg_0593;
    8: op1_10_in13 = imem06_in[3:0];
    9: op1_10_in13 = reg_0195;
    10: op1_10_in13 = reg_0787;
    11: op1_10_in13 = imem03_in[15:12];
    12: op1_10_in13 = imem07_in[127:124];
    13: op1_10_in13 = reg_0976;
    14: op1_10_in13 = reg_0217;
    15: op1_10_in13 = imem07_in[39:36];
    16: op1_10_in13 = reg_0659;
    17: op1_10_in13 = reg_0289;
    4: op1_10_in13 = reg_0170;
    18: op1_10_in13 = reg_0661;
    19: op1_10_in13 = reg_0277;
    20: op1_10_in13 = reg_0647;
    21: op1_10_in13 = reg_0864;
    22: op1_10_in13 = reg_0459;
    23: op1_10_in13 = imem01_in[15:12];
    24: op1_10_in13 = reg_0453;
    25: op1_10_in13 = reg_0359;
    26: op1_10_in13 = reg_0375;
    27: op1_10_in13 = imem04_in[19:16];
    28: op1_10_in13 = imem04_in[107:104];
    29: op1_10_in13 = reg_0227;
    30: op1_10_in13 = imem02_in[27:24];
    31: op1_10_in13 = reg_0259;
    32: op1_10_in13 = imem06_in[79:76];
    34: op1_10_in13 = reg_0665;
    35: op1_10_in13 = reg_0622;
    36: op1_10_in13 = imem06_in[35:32];
    37: op1_10_in13 = reg_0167;
    38: op1_10_in13 = reg_0925;
    39: op1_10_in13 = reg_0478;
    40: op1_10_in13 = imem02_in[123:120];
    41: op1_10_in13 = reg_0097;
    42: op1_10_in13 = reg_0894;
    43: op1_10_in13 = imem07_in[71:68];
    44: op1_10_in13 = imem01_in[19:16];
    45: op1_10_in13 = reg_0284;
    46: op1_10_in13 = reg_0152;
    47: op1_10_in13 = reg_0452;
    48: op1_10_in13 = reg_0055;
    49: op1_10_in13 = reg_0128;
    50: op1_10_in13 = reg_0923;
    51: op1_10_in13 = reg_0886;
    52: op1_10_in13 = reg_0191;
    53: op1_10_in13 = reg_0649;
    54: op1_10_in13 = reg_0655;
    55: op1_10_in13 = imem05_in[55:52];
    56: op1_10_in13 = reg_0336;
    57: op1_10_in13 = reg_0569;
    58: op1_10_in13 = reg_0142;
    59: op1_10_in13 = reg_0005;
    60: op1_10_in13 = reg_0005;
    62: op1_10_in13 = reg_0669;
    63: op1_10_in13 = imem04_in[15:12];
    64: op1_10_in13 = reg_1004;
    65: op1_10_in13 = imem05_in[63:60];
    66: op1_10_in13 = imem06_in[31:28];
    67: op1_10_in13 = reg_0964;
    68: op1_10_in13 = reg_0209;
    69: op1_10_in13 = imem02_in[87:84];
    70: op1_10_in13 = reg_0386;
    71: op1_10_in13 = reg_0838;
    72: op1_10_in13 = imem04_in[43:40];
    73: op1_10_in13 = imem07_in[3:0];
    74: op1_10_in13 = imem06_in[11:8];
    76: op1_10_in13 = reg_0186;
    77: op1_10_in13 = reg_0762;
    78: op1_10_in13 = reg_0368;
    79: op1_10_in13 = imem04_in[123:120];
    80: op1_10_in13 = reg_0382;
    81: op1_10_in13 = reg_0718;
    82: op1_10_in13 = imem06_in[95:92];
    83: op1_10_in13 = reg_0979;
    84: op1_10_in13 = reg_0680;
    85: op1_10_in13 = reg_0651;
    87: op1_10_in13 = reg_0052;
    88: op1_10_in13 = reg_0947;
    89: op1_10_in13 = reg_0335;
    90: op1_10_in13 = reg_0295;
    91: op1_10_in13 = imem05_in[59:56];
    92: op1_10_in13 = reg_0567;
    93: op1_10_in13 = reg_0205;
    95: op1_10_in13 = reg_0471;
    96: op1_10_in13 = reg_0216;
    default: op1_10_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv13 = 1;
    6: op1_10_inv13 = 1;
    7: op1_10_inv13 = 1;
    11: op1_10_inv13 = 1;
    17: op1_10_inv13 = 1;
    19: op1_10_inv13 = 1;
    20: op1_10_inv13 = 1;
    21: op1_10_inv13 = 1;
    22: op1_10_inv13 = 1;
    23: op1_10_inv13 = 1;
    28: op1_10_inv13 = 1;
    35: op1_10_inv13 = 1;
    36: op1_10_inv13 = 1;
    37: op1_10_inv13 = 1;
    38: op1_10_inv13 = 1;
    41: op1_10_inv13 = 1;
    43: op1_10_inv13 = 1;
    46: op1_10_inv13 = 1;
    47: op1_10_inv13 = 1;
    49: op1_10_inv13 = 1;
    52: op1_10_inv13 = 1;
    54: op1_10_inv13 = 1;
    55: op1_10_inv13 = 1;
    57: op1_10_inv13 = 1;
    59: op1_10_inv13 = 1;
    60: op1_10_inv13 = 1;
    62: op1_10_inv13 = 1;
    63: op1_10_inv13 = 1;
    66: op1_10_inv13 = 1;
    67: op1_10_inv13 = 1;
    68: op1_10_inv13 = 1;
    71: op1_10_inv13 = 1;
    72: op1_10_inv13 = 1;
    74: op1_10_inv13 = 1;
    77: op1_10_inv13 = 1;
    78: op1_10_inv13 = 1;
    81: op1_10_inv13 = 1;
    83: op1_10_inv13 = 1;
    85: op1_10_inv13 = 1;
    87: op1_10_inv13 = 1;
    89: op1_10_inv13 = 1;
    91: op1_10_inv13 = 1;
    92: op1_10_inv13 = 1;
    96: op1_10_inv13 = 1;
    default: op1_10_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in14 = reg_0191;
    6: op1_10_in14 = reg_0470;
    7: op1_10_in14 = reg_0395;
    8: op1_10_in14 = imem06_in[15:12];
    9: op1_10_in14 = imem01_in[35:32];
    76: op1_10_in14 = imem01_in[35:32];
    10: op1_10_in14 = reg_0025;
    11: op1_10_in14 = imem03_in[19:16];
    12: op1_10_in14 = reg_0731;
    13: op1_10_in14 = imem04_in[11:8];
    14: op1_10_in14 = reg_0836;
    15: op1_10_in14 = imem07_in[95:92];
    16: op1_10_in14 = reg_0352;
    17: op1_10_in14 = reg_0306;
    4: op1_10_in14 = reg_0176;
    96: op1_10_in14 = reg_0176;
    18: op1_10_in14 = reg_0641;
    19: op1_10_in14 = reg_0048;
    20: op1_10_in14 = reg_0640;
    21: op1_10_in14 = reg_0856;
    22: op1_10_in14 = reg_0209;
    23: op1_10_in14 = imem01_in[59:56];
    24: op1_10_in14 = reg_0450;
    25: op1_10_in14 = reg_0345;
    26: op1_10_in14 = reg_0404;
    27: op1_10_in14 = imem04_in[27:24];
    28: op1_10_in14 = reg_1004;
    79: op1_10_in14 = reg_1004;
    29: op1_10_in14 = reg_1031;
    30: op1_10_in14 = imem02_in[47:44];
    31: op1_10_in14 = reg_0071;
    32: op1_10_in14 = imem06_in[103:100];
    34: op1_10_in14 = reg_0652;
    35: op1_10_in14 = reg_0385;
    36: op1_10_in14 = imem06_in[51:48];
    37: op1_10_in14 = reg_0169;
    38: op1_10_in14 = reg_0618;
    39: op1_10_in14 = reg_0198;
    40: op1_10_in14 = imem02_in[127:124];
    41: op1_10_in14 = reg_0225;
    42: op1_10_in14 = reg_0241;
    43: op1_10_in14 = imem07_in[107:104];
    44: op1_10_in14 = imem01_in[23:20];
    45: op1_10_in14 = reg_0748;
    46: op1_10_in14 = reg_0130;
    47: op1_10_in14 = reg_0456;
    48: op1_10_in14 = reg_0507;
    49: op1_10_in14 = reg_0154;
    50: op1_10_in14 = reg_0370;
    51: op1_10_in14 = reg_0865;
    52: op1_10_in14 = reg_0186;
    53: op1_10_in14 = reg_0651;
    54: op1_10_in14 = reg_0854;
    55: op1_10_in14 = imem05_in[79:76];
    56: op1_10_in14 = reg_0132;
    57: op1_10_in14 = reg_0835;
    58: op1_10_in14 = reg_0137;
    59: op1_10_in14 = reg_0545;
    60: op1_10_in14 = imem07_in[39:36];
    62: op1_10_in14 = reg_0473;
    63: op1_10_in14 = imem04_in[51:48];
    64: op1_10_in14 = reg_0055;
    65: op1_10_in14 = imem05_in[67:64];
    66: op1_10_in14 = imem06_in[43:40];
    67: op1_10_in14 = reg_0782;
    68: op1_10_in14 = imem01_in[7:4];
    69: op1_10_in14 = imem02_in[103:100];
    70: op1_10_in14 = reg_0633;
    71: op1_10_in14 = reg_0161;
    72: op1_10_in14 = imem04_in[47:44];
    73: op1_10_in14 = imem07_in[7:4];
    74: op1_10_in14 = imem06_in[63:60];
    77: op1_10_in14 = reg_0323;
    78: op1_10_in14 = reg_0425;
    80: op1_10_in14 = reg_0632;
    81: op1_10_in14 = reg_0002;
    82: op1_10_in14 = imem06_in[99:96];
    83: op1_10_in14 = reg_0980;
    84: op1_10_in14 = reg_0454;
    85: op1_10_in14 = reg_0146;
    87: op1_10_in14 = reg_0368;
    88: op1_10_in14 = reg_0152;
    89: op1_10_in14 = reg_0347;
    90: op1_10_in14 = imem05_in[27:24];
    91: op1_10_in14 = imem05_in[71:68];
    92: op1_10_in14 = reg_0710;
    93: op1_10_in14 = reg_0364;
    94: op1_10_in14 = reg_0458;
    95: op1_10_in14 = reg_0200;
    default: op1_10_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv14 = 1;
    6: op1_10_inv14 = 1;
    8: op1_10_inv14 = 1;
    9: op1_10_inv14 = 1;
    12: op1_10_inv14 = 1;
    13: op1_10_inv14 = 1;
    14: op1_10_inv14 = 1;
    15: op1_10_inv14 = 1;
    17: op1_10_inv14 = 1;
    24: op1_10_inv14 = 1;
    25: op1_10_inv14 = 1;
    27: op1_10_inv14 = 1;
    29: op1_10_inv14 = 1;
    30: op1_10_inv14 = 1;
    37: op1_10_inv14 = 1;
    40: op1_10_inv14 = 1;
    41: op1_10_inv14 = 1;
    42: op1_10_inv14 = 1;
    44: op1_10_inv14 = 1;
    45: op1_10_inv14 = 1;
    46: op1_10_inv14 = 1;
    47: op1_10_inv14 = 1;
    49: op1_10_inv14 = 1;
    53: op1_10_inv14 = 1;
    54: op1_10_inv14 = 1;
    55: op1_10_inv14 = 1;
    56: op1_10_inv14 = 1;
    62: op1_10_inv14 = 1;
    65: op1_10_inv14 = 1;
    67: op1_10_inv14 = 1;
    68: op1_10_inv14 = 1;
    71: op1_10_inv14 = 1;
    72: op1_10_inv14 = 1;
    73: op1_10_inv14 = 1;
    74: op1_10_inv14 = 1;
    78: op1_10_inv14 = 1;
    79: op1_10_inv14 = 1;
    82: op1_10_inv14 = 1;
    84: op1_10_inv14 = 1;
    85: op1_10_inv14 = 1;
    88: op1_10_inv14 = 1;
    91: op1_10_inv14 = 1;
    92: op1_10_inv14 = 1;
    93: op1_10_inv14 = 1;
    94: op1_10_inv14 = 1;
    95: op1_10_inv14 = 1;
    default: op1_10_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in15 = reg_0210;
    6: op1_10_in15 = reg_0203;
    22: op1_10_in15 = reg_0203;
    95: op1_10_in15 = reg_0203;
    7: op1_10_in15 = reg_0391;
    8: op1_10_in15 = imem06_in[47:44];
    9: op1_10_in15 = imem01_in[55:52];
    68: op1_10_in15 = imem01_in[55:52];
    10: op1_10_in15 = reg_0781;
    11: op1_10_in15 = imem03_in[47:44];
    12: op1_10_in15 = reg_0702;
    13: op1_10_in15 = imem04_in[59:56];
    14: op1_10_in15 = reg_0258;
    15: op1_10_in15 = imem07_in[103:100];
    16: op1_10_in15 = reg_0364;
    17: op1_10_in15 = reg_0302;
    4: op1_10_in15 = reg_0158;
    18: op1_10_in15 = reg_0325;
    19: op1_10_in15 = reg_0756;
    20: op1_10_in15 = reg_0649;
    21: op1_10_in15 = imem05_in[11:8];
    23: op1_10_in15 = imem01_in[79:76];
    24: op1_10_in15 = reg_0464;
    25: op1_10_in15 = reg_0363;
    26: op1_10_in15 = reg_0027;
    27: op1_10_in15 = imem04_in[43:40];
    28: op1_10_in15 = reg_0483;
    29: op1_10_in15 = reg_1015;
    30: op1_10_in15 = imem02_in[123:120];
    31: op1_10_in15 = reg_0063;
    32: op1_10_in15 = imem07_in[3:0];
    34: op1_10_in15 = reg_0097;
    35: op1_10_in15 = reg_0356;
    36: op1_10_in15 = imem06_in[71:68];
    37: op1_10_in15 = reg_0170;
    38: op1_10_in15 = reg_0406;
    39: op1_10_in15 = reg_0196;
    40: op1_10_in15 = reg_0666;
    41: op1_10_in15 = reg_0098;
    42: op1_10_in15 = reg_0596;
    43: op1_10_in15 = imem07_in[115:112];
    44: op1_10_in15 = imem01_in[27:24];
    45: op1_10_in15 = reg_0773;
    46: op1_10_in15 = reg_0155;
    47: op1_10_in15 = reg_0209;
    48: op1_10_in15 = reg_0014;
    49: op1_10_in15 = reg_0139;
    50: op1_10_in15 = reg_0246;
    51: op1_10_in15 = reg_0482;
    52: op1_10_in15 = reg_0194;
    94: op1_10_in15 = reg_0194;
    53: op1_10_in15 = reg_0621;
    54: op1_10_in15 = reg_0664;
    55: op1_10_in15 = imem05_in[103:100];
    56: op1_10_in15 = reg_0154;
    57: op1_10_in15 = reg_0233;
    58: op1_10_in15 = reg_0486;
    59: op1_10_in15 = reg_0263;
    60: op1_10_in15 = imem07_in[67:64];
    62: op1_10_in15 = reg_0467;
    63: op1_10_in15 = imem04_in[67:64];
    64: op1_10_in15 = reg_0292;
    65: op1_10_in15 = imem05_in[87:84];
    66: op1_10_in15 = imem06_in[55:52];
    67: op1_10_in15 = reg_0968;
    69: op1_10_in15 = imem02_in[107:104];
    70: op1_10_in15 = reg_0399;
    71: op1_10_in15 = reg_0169;
    72: op1_10_in15 = imem04_in[75:72];
    73: op1_10_in15 = imem07_in[35:32];
    74: op1_10_in15 = imem06_in[91:88];
    76: op1_10_in15 = imem01_in[63:60];
    77: op1_10_in15 = reg_0358;
    78: op1_10_in15 = reg_0248;
    79: op1_10_in15 = reg_1003;
    80: op1_10_in15 = reg_0026;
    81: op1_10_in15 = reg_0422;
    82: op1_10_in15 = imem06_in[111:108];
    83: op1_10_in15 = reg_0977;
    84: op1_10_in15 = reg_0450;
    85: op1_10_in15 = reg_0795;
    87: op1_10_in15 = reg_0335;
    88: op1_10_in15 = reg_0956;
    89: op1_10_in15 = reg_0341;
    90: op1_10_in15 = reg_0492;
    91: op1_10_in15 = imem05_in[91:88];
    92: op1_10_in15 = reg_0721;
    93: op1_10_in15 = reg_0369;
    96: op1_10_in15 = reg_0737;
    default: op1_10_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv15 = 1;
    8: op1_10_inv15 = 1;
    15: op1_10_inv15 = 1;
    16: op1_10_inv15 = 1;
    17: op1_10_inv15 = 1;
    4: op1_10_inv15 = 1;
    18: op1_10_inv15 = 1;
    20: op1_10_inv15 = 1;
    21: op1_10_inv15 = 1;
    22: op1_10_inv15 = 1;
    25: op1_10_inv15 = 1;
    26: op1_10_inv15 = 1;
    27: op1_10_inv15 = 1;
    28: op1_10_inv15 = 1;
    29: op1_10_inv15 = 1;
    30: op1_10_inv15 = 1;
    34: op1_10_inv15 = 1;
    35: op1_10_inv15 = 1;
    37: op1_10_inv15 = 1;
    39: op1_10_inv15 = 1;
    40: op1_10_inv15 = 1;
    42: op1_10_inv15 = 1;
    44: op1_10_inv15 = 1;
    45: op1_10_inv15 = 1;
    48: op1_10_inv15 = 1;
    51: op1_10_inv15 = 1;
    52: op1_10_inv15 = 1;
    55: op1_10_inv15 = 1;
    56: op1_10_inv15 = 1;
    57: op1_10_inv15 = 1;
    59: op1_10_inv15 = 1;
    60: op1_10_inv15 = 1;
    62: op1_10_inv15 = 1;
    64: op1_10_inv15 = 1;
    67: op1_10_inv15 = 1;
    71: op1_10_inv15 = 1;
    72: op1_10_inv15 = 1;
    74: op1_10_inv15 = 1;
    76: op1_10_inv15 = 1;
    81: op1_10_inv15 = 1;
    82: op1_10_inv15 = 1;
    84: op1_10_inv15 = 1;
    88: op1_10_inv15 = 1;
    89: op1_10_inv15 = 1;
    92: op1_10_inv15 = 1;
    94: op1_10_inv15 = 1;
    95: op1_10_inv15 = 1;
    96: op1_10_inv15 = 1;
    default: op1_10_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in16 = reg_0204;
    6: op1_10_in16 = reg_0193;
    7: op1_10_in16 = reg_0362;
    8: op1_10_in16 = imem06_in[71:68];
    9: op1_10_in16 = imem01_in[111:108];
    10: op1_10_in16 = reg_1010;
    11: op1_10_in16 = imem03_in[55:52];
    12: op1_10_in16 = reg_0718;
    13: op1_10_in16 = imem04_in[87:84];
    14: op1_10_in16 = reg_0898;
    15: op1_10_in16 = imem07_in[107:104];
    16: op1_10_in16 = reg_0310;
    17: op1_10_in16 = reg_0291;
    4: op1_10_in16 = reg_0171;
    18: op1_10_in16 = reg_0359;
    19: op1_10_in16 = reg_0857;
    20: op1_10_in16 = reg_0644;
    78: op1_10_in16 = reg_0644;
    21: op1_10_in16 = imem05_in[55:52];
    22: op1_10_in16 = reg_0207;
    23: op1_10_in16 = reg_0013;
    90: op1_10_in16 = reg_0013;
    24: op1_10_in16 = reg_0459;
    25: op1_10_in16 = reg_0365;
    26: op1_10_in16 = reg_0752;
    27: op1_10_in16 = imem04_in[103:100];
    28: op1_10_in16 = reg_1006;
    29: op1_10_in16 = reg_1045;
    30: op1_10_in16 = reg_0658;
    31: op1_10_in16 = reg_0882;
    32: op1_10_in16 = imem07_in[15:12];
    34: op1_10_in16 = reg_0338;
    35: op1_10_in16 = reg_0395;
    36: op1_10_in16 = imem06_in[95:92];
    37: op1_10_in16 = reg_0184;
    38: op1_10_in16 = reg_0588;
    39: op1_10_in16 = reg_0206;
    40: op1_10_in16 = reg_0637;
    41: op1_10_in16 = reg_0762;
    42: op1_10_in16 = reg_0631;
    43: op1_10_in16 = imem07_in[123:120];
    44: op1_10_in16 = imem01_in[35:32];
    45: op1_10_in16 = reg_0970;
    46: op1_10_in16 = reg_0131;
    47: op1_10_in16 = reg_0186;
    48: op1_10_in16 = reg_0015;
    49: op1_10_in16 = reg_0130;
    50: op1_10_in16 = reg_0987;
    51: op1_10_in16 = reg_0876;
    52: op1_10_in16 = reg_0190;
    53: op1_10_in16 = reg_0300;
    54: op1_10_in16 = reg_0394;
    55: op1_10_in16 = imem05_in[111:108];
    56: op1_10_in16 = reg_0139;
    57: op1_10_in16 = reg_0215;
    58: op1_10_in16 = reg_0317;
    59: op1_10_in16 = imem07_in[31:28];
    60: op1_10_in16 = imem07_in[87:84];
    62: op1_10_in16 = reg_0470;
    63: op1_10_in16 = imem04_in[95:92];
    64: op1_10_in16 = reg_0888;
    65: op1_10_in16 = imem05_in[91:88];
    66: op1_10_in16 = imem06_in[87:84];
    67: op1_10_in16 = reg_0896;
    68: op1_10_in16 = imem01_in[71:68];
    69: op1_10_in16 = reg_0355;
    70: op1_10_in16 = reg_0219;
    71: op1_10_in16 = reg_0182;
    72: op1_10_in16 = imem04_in[107:104];
    73: op1_10_in16 = imem07_in[43:40];
    74: op1_10_in16 = reg_0696;
    76: op1_10_in16 = imem01_in[99:96];
    77: op1_10_in16 = reg_0441;
    79: op1_10_in16 = reg_0937;
    80: op1_10_in16 = reg_0017;
    81: op1_10_in16 = reg_0421;
    82: op1_10_in16 = imem06_in[115:112];
    83: op1_10_in16 = reg_0990;
    84: op1_10_in16 = reg_0464;
    85: op1_10_in16 = reg_0950;
    87: op1_10_in16 = reg_0734;
    88: op1_10_in16 = reg_0260;
    89: op1_10_in16 = imem03_in[39:36];
    91: op1_10_in16 = reg_0652;
    92: op1_10_in16 = reg_0299;
    93: op1_10_in16 = reg_0849;
    94: op1_10_in16 = reg_0198;
    95: op1_10_in16 = reg_0236;
    96: op1_10_in16 = reg_0877;
    default: op1_10_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv16 = 1;
    9: op1_10_inv16 = 1;
    10: op1_10_inv16 = 1;
    16: op1_10_inv16 = 1;
    17: op1_10_inv16 = 1;
    22: op1_10_inv16 = 1;
    23: op1_10_inv16 = 1;
    26: op1_10_inv16 = 1;
    27: op1_10_inv16 = 1;
    29: op1_10_inv16 = 1;
    30: op1_10_inv16 = 1;
    34: op1_10_inv16 = 1;
    35: op1_10_inv16 = 1;
    36: op1_10_inv16 = 1;
    37: op1_10_inv16 = 1;
    38: op1_10_inv16 = 1;
    39: op1_10_inv16 = 1;
    40: op1_10_inv16 = 1;
    41: op1_10_inv16 = 1;
    43: op1_10_inv16 = 1;
    45: op1_10_inv16 = 1;
    48: op1_10_inv16 = 1;
    49: op1_10_inv16 = 1;
    51: op1_10_inv16 = 1;
    55: op1_10_inv16 = 1;
    57: op1_10_inv16 = 1;
    59: op1_10_inv16 = 1;
    60: op1_10_inv16 = 1;
    62: op1_10_inv16 = 1;
    65: op1_10_inv16 = 1;
    67: op1_10_inv16 = 1;
    69: op1_10_inv16 = 1;
    79: op1_10_inv16 = 1;
    83: op1_10_inv16 = 1;
    85: op1_10_inv16 = 1;
    89: op1_10_inv16 = 1;
    90: op1_10_inv16 = 1;
    91: op1_10_inv16 = 1;
    92: op1_10_inv16 = 1;
    94: op1_10_inv16 = 1;
    95: op1_10_inv16 = 1;
    default: op1_10_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in17 = reg_0211;
    6: op1_10_in17 = reg_0207;
    7: op1_10_in17 = reg_0373;
    8: op1_10_in17 = imem06_in[111:108];
    9: op1_10_in17 = reg_0514;
    10: op1_10_in17 = reg_1011;
    11: op1_10_in17 = imem03_in[95:92];
    12: op1_10_in17 = reg_0711;
    13: op1_10_in17 = reg_0549;
    14: op1_10_in17 = reg_0132;
    15: op1_10_in17 = reg_0722;
    16: op1_10_in17 = reg_0365;
    17: op1_10_in17 = reg_0297;
    18: op1_10_in17 = reg_0083;
    19: op1_10_in17 = reg_0484;
    20: op1_10_in17 = reg_0663;
    21: op1_10_in17 = reg_0959;
    22: op1_10_in17 = reg_0206;
    23: op1_10_in17 = reg_0242;
    24: op1_10_in17 = reg_0214;
    25: op1_10_in17 = reg_0342;
    26: op1_10_in17 = imem07_in[35:32];
    27: op1_10_in17 = reg_1016;
    28: op1_10_in17 = reg_0301;
    29: op1_10_in17 = reg_0871;
    30: op1_10_in17 = reg_0656;
    31: op1_10_in17 = reg_0009;
    32: op1_10_in17 = imem07_in[39:36];
    34: op1_10_in17 = reg_0007;
    35: op1_10_in17 = reg_0914;
    36: op1_10_in17 = imem06_in[115:112];
    66: op1_10_in17 = imem06_in[115:112];
    38: op1_10_in17 = reg_0042;
    39: op1_10_in17 = imem01_in[7:4];
    52: op1_10_in17 = imem01_in[7:4];
    40: op1_10_in17 = reg_0640;
    41: op1_10_in17 = reg_0772;
    42: op1_10_in17 = reg_0029;
    43: op1_10_in17 = reg_0181;
    44: op1_10_in17 = imem01_in[43:40];
    45: op1_10_in17 = reg_0969;
    46: op1_10_in17 = imem06_in[27:24];
    47: op1_10_in17 = imem01_in[3:0];
    48: op1_10_in17 = reg_0074;
    49: op1_10_in17 = reg_0140;
    50: op1_10_in17 = reg_0979;
    51: op1_10_in17 = reg_0090;
    53: op1_10_in17 = reg_0652;
    54: op1_10_in17 = reg_0368;
    55: op1_10_in17 = reg_0970;
    56: op1_10_in17 = reg_0138;
    57: op1_10_in17 = reg_0488;
    58: op1_10_in17 = reg_0093;
    59: op1_10_in17 = imem07_in[83:80];
    60: op1_10_in17 = imem07_in[91:88];
    62: op1_10_in17 = reg_0479;
    63: op1_10_in17 = imem04_in[119:116];
    64: op1_10_in17 = reg_0313;
    65: op1_10_in17 = imem05_in[107:104];
    67: op1_10_in17 = reg_0256;
    68: op1_10_in17 = imem01_in[115:112];
    69: op1_10_in17 = reg_0666;
    70: op1_10_in17 = imem07_in[43:40];
    71: op1_10_in17 = reg_0158;
    72: op1_10_in17 = reg_0483;
    73: op1_10_in17 = imem07_in[47:44];
    74: op1_10_in17 = reg_0691;
    76: op1_10_in17 = imem01_in[127:124];
    77: op1_10_in17 = reg_0424;
    78: op1_10_in17 = reg_0037;
    79: op1_10_in17 = reg_0912;
    80: op1_10_in17 = reg_0915;
    81: op1_10_in17 = reg_0350;
    82: op1_10_in17 = reg_1019;
    83: op1_10_in17 = reg_0997;
    84: op1_10_in17 = reg_0469;
    85: op1_10_in17 = imem06_in[7:4];
    87: op1_10_in17 = reg_0381;
    88: op1_10_in17 = reg_0587;
    89: op1_10_in17 = imem03_in[91:88];
    90: op1_10_in17 = reg_0226;
    91: op1_10_in17 = reg_0954;
    92: op1_10_in17 = reg_0250;
    93: op1_10_in17 = reg_0120;
    94: op1_10_in17 = reg_0196;
    95: op1_10_in17 = reg_0399;
    96: op1_10_in17 = reg_0096;
    default: op1_10_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_10_inv17 = 1;
    8: op1_10_inv17 = 1;
    10: op1_10_inv17 = 1;
    12: op1_10_inv17 = 1;
    13: op1_10_inv17 = 1;
    16: op1_10_inv17 = 1;
    20: op1_10_inv17 = 1;
    21: op1_10_inv17 = 1;
    22: op1_10_inv17 = 1;
    24: op1_10_inv17 = 1;
    26: op1_10_inv17 = 1;
    28: op1_10_inv17 = 1;
    29: op1_10_inv17 = 1;
    35: op1_10_inv17 = 1;
    39: op1_10_inv17 = 1;
    40: op1_10_inv17 = 1;
    41: op1_10_inv17 = 1;
    43: op1_10_inv17 = 1;
    45: op1_10_inv17 = 1;
    47: op1_10_inv17 = 1;
    49: op1_10_inv17 = 1;
    50: op1_10_inv17 = 1;
    51: op1_10_inv17 = 1;
    53: op1_10_inv17 = 1;
    54: op1_10_inv17 = 1;
    56: op1_10_inv17 = 1;
    58: op1_10_inv17 = 1;
    59: op1_10_inv17 = 1;
    60: op1_10_inv17 = 1;
    63: op1_10_inv17 = 1;
    66: op1_10_inv17 = 1;
    67: op1_10_inv17 = 1;
    68: op1_10_inv17 = 1;
    69: op1_10_inv17 = 1;
    72: op1_10_inv17 = 1;
    76: op1_10_inv17 = 1;
    77: op1_10_inv17 = 1;
    78: op1_10_inv17 = 1;
    83: op1_10_inv17 = 1;
    88: op1_10_inv17 = 1;
    89: op1_10_inv17 = 1;
    90: op1_10_inv17 = 1;
    92: op1_10_inv17 = 1;
    93: op1_10_inv17 = 1;
    95: op1_10_inv17 = 1;
    default: op1_10_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in18 = reg_0196;
    6: op1_10_in18 = reg_0211;
    24: op1_10_in18 = reg_0211;
    7: op1_10_in18 = reg_0369;
    8: op1_10_in18 = reg_0628;
    9: op1_10_in18 = reg_0517;
    10: op1_10_in18 = reg_0798;
    11: op1_10_in18 = imem03_in[99:96];
    12: op1_10_in18 = reg_0706;
    13: op1_10_in18 = reg_0533;
    14: op1_10_in18 = reg_0129;
    15: op1_10_in18 = reg_0717;
    16: op1_10_in18 = reg_0342;
    17: op1_10_in18 = reg_0069;
    18: op1_10_in18 = reg_0088;
    19: op1_10_in18 = reg_0742;
    20: op1_10_in18 = reg_0334;
    21: op1_10_in18 = reg_0956;
    22: op1_10_in18 = reg_0192;
    23: op1_10_in18 = reg_0248;
    25: op1_10_in18 = reg_0355;
    26: op1_10_in18 = imem07_in[55:52];
    27: op1_10_in18 = reg_0541;
    28: op1_10_in18 = reg_0530;
    83: op1_10_in18 = reg_0530;
    29: op1_10_in18 = reg_0123;
    30: op1_10_in18 = reg_0639;
    31: op1_10_in18 = reg_0047;
    32: op1_10_in18 = reg_0726;
    34: op1_10_in18 = reg_0084;
    35: op1_10_in18 = reg_0392;
    36: op1_10_in18 = reg_0914;
    38: op1_10_in18 = reg_0386;
    39: op1_10_in18 = imem01_in[11:8];
    40: op1_10_in18 = reg_0638;
    41: op1_10_in18 = reg_0007;
    42: op1_10_in18 = imem07_in[15:12];
    43: op1_10_in18 = reg_0161;
    44: op1_10_in18 = imem01_in[67:64];
    45: op1_10_in18 = reg_0950;
    46: op1_10_in18 = imem06_in[43:40];
    47: op1_10_in18 = imem01_in[47:44];
    48: op1_10_in18 = reg_0893;
    49: op1_10_in18 = imem06_in[7:4];
    50: op1_10_in18 = reg_0984;
    51: op1_10_in18 = imem03_in[43:40];
    52: op1_10_in18 = imem01_in[19:16];
    53: op1_10_in18 = reg_0418;
    54: op1_10_in18 = reg_0037;
    55: op1_10_in18 = reg_0967;
    56: op1_10_in18 = reg_0614;
    57: op1_10_in18 = reg_0508;
    58: op1_10_in18 = reg_0673;
    59: op1_10_in18 = imem07_in[103:100];
    60: op1_10_in18 = imem07_in[119:116];
    62: op1_10_in18 = imem01_in[3:0];
    63: op1_10_in18 = reg_1004;
    64: op1_10_in18 = reg_0802;
    65: op1_10_in18 = imem05_in[111:108];
    66: op1_10_in18 = reg_0694;
    67: op1_10_in18 = reg_0603;
    68: op1_10_in18 = imem01_in[119:116];
    69: op1_10_in18 = reg_0654;
    70: op1_10_in18 = imem07_in[67:64];
    81: op1_10_in18 = imem07_in[67:64];
    72: op1_10_in18 = reg_0277;
    73: op1_10_in18 = imem07_in[79:76];
    74: op1_10_in18 = reg_1018;
    76: op1_10_in18 = reg_0973;
    77: op1_10_in18 = reg_0644;
    78: op1_10_in18 = reg_0335;
    79: op1_10_in18 = reg_0539;
    80: op1_10_in18 = reg_0383;
    82: op1_10_in18 = reg_0025;
    84: op1_10_in18 = reg_0474;
    85: op1_10_in18 = imem06_in[23:20];
    87: op1_10_in18 = reg_0700;
    88: op1_10_in18 = reg_0951;
    89: op1_10_in18 = imem03_in[127:124];
    90: op1_10_in18 = reg_0152;
    91: op1_10_in18 = reg_0319;
    92: op1_10_in18 = reg_0422;
    93: op1_10_in18 = reg_0237;
    94: op1_10_in18 = reg_0197;
    95: op1_10_in18 = reg_1039;
    96: op1_10_in18 = reg_0845;
    default: op1_10_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv18 = 1;
    6: op1_10_inv18 = 1;
    7: op1_10_inv18 = 1;
    8: op1_10_inv18 = 1;
    12: op1_10_inv18 = 1;
    16: op1_10_inv18 = 1;
    17: op1_10_inv18 = 1;
    18: op1_10_inv18 = 1;
    19: op1_10_inv18 = 1;
    21: op1_10_inv18 = 1;
    22: op1_10_inv18 = 1;
    23: op1_10_inv18 = 1;
    24: op1_10_inv18 = 1;
    25: op1_10_inv18 = 1;
    28: op1_10_inv18 = 1;
    35: op1_10_inv18 = 1;
    43: op1_10_inv18 = 1;
    44: op1_10_inv18 = 1;
    45: op1_10_inv18 = 1;
    46: op1_10_inv18 = 1;
    50: op1_10_inv18 = 1;
    51: op1_10_inv18 = 1;
    52: op1_10_inv18 = 1;
    55: op1_10_inv18 = 1;
    56: op1_10_inv18 = 1;
    57: op1_10_inv18 = 1;
    58: op1_10_inv18 = 1;
    59: op1_10_inv18 = 1;
    60: op1_10_inv18 = 1;
    62: op1_10_inv18 = 1;
    63: op1_10_inv18 = 1;
    65: op1_10_inv18 = 1;
    67: op1_10_inv18 = 1;
    68: op1_10_inv18 = 1;
    76: op1_10_inv18 = 1;
    77: op1_10_inv18 = 1;
    78: op1_10_inv18 = 1;
    80: op1_10_inv18 = 1;
    82: op1_10_inv18 = 1;
    83: op1_10_inv18 = 1;
    85: op1_10_inv18 = 1;
    87: op1_10_inv18 = 1;
    88: op1_10_inv18 = 1;
    89: op1_10_inv18 = 1;
    90: op1_10_inv18 = 1;
    94: op1_10_inv18 = 1;
    96: op1_10_inv18 = 1;
    default: op1_10_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in19 = reg_0195;
    6: op1_10_in19 = reg_0201;
    7: op1_10_in19 = reg_0322;
    8: op1_10_in19 = reg_0621;
    9: op1_10_in19 = reg_0506;
    10: op1_10_in19 = imem07_in[7:4];
    11: op1_10_in19 = imem03_in[119:116];
    12: op1_10_in19 = reg_0429;
    13: op1_10_in19 = reg_0531;
    14: op1_10_in19 = reg_0131;
    15: op1_10_in19 = reg_0712;
    32: op1_10_in19 = reg_0712;
    16: op1_10_in19 = reg_0086;
    17: op1_10_in19 = reg_0074;
    18: op1_10_in19 = reg_0080;
    19: op1_10_in19 = reg_0485;
    20: op1_10_in19 = reg_0359;
    21: op1_10_in19 = reg_0951;
    22: op1_10_in19 = reg_0197;
    23: op1_10_in19 = reg_0487;
    93: op1_10_in19 = reg_0487;
    24: op1_10_in19 = reg_0186;
    25: op1_10_in19 = reg_0007;
    26: op1_10_in19 = imem07_in[63:60];
    27: op1_10_in19 = reg_0537;
    28: op1_10_in19 = reg_0937;
    29: op1_10_in19 = reg_0105;
    30: op1_10_in19 = reg_0647;
    31: op1_10_in19 = reg_0855;
    34: op1_10_in19 = reg_0840;
    35: op1_10_in19 = reg_0741;
    38: op1_10_in19 = reg_0741;
    36: op1_10_in19 = reg_0351;
    39: op1_10_in19 = imem01_in[35:32];
    40: op1_10_in19 = reg_0644;
    41: op1_10_in19 = reg_0758;
    42: op1_10_in19 = imem07_in[31:28];
    43: op1_10_in19 = reg_0159;
    44: op1_10_in19 = imem01_in[127:124];
    45: op1_10_in19 = reg_0942;
    46: op1_10_in19 = imem06_in[95:92];
    47: op1_10_in19 = imem01_in[83:80];
    48: op1_10_in19 = reg_0279;
    49: op1_10_in19 = imem06_in[23:20];
    50: op1_10_in19 = imem04_in[39:36];
    51: op1_10_in19 = imem03_in[47:44];
    52: op1_10_in19 = imem01_in[87:84];
    53: op1_10_in19 = reg_0664;
    54: op1_10_in19 = reg_0088;
    55: op1_10_in19 = reg_0968;
    56: op1_10_in19 = reg_0073;
    57: op1_10_in19 = reg_0252;
    58: op1_10_in19 = reg_0573;
    59: op1_10_in19 = imem07_in[119:116];
    60: op1_10_in19 = reg_0723;
    62: op1_10_in19 = imem01_in[15:12];
    63: op1_10_in19 = reg_0483;
    64: op1_10_in19 = reg_0568;
    65: op1_10_in19 = reg_0774;
    66: op1_10_in19 = reg_0624;
    87: op1_10_in19 = reg_0624;
    67: op1_10_in19 = reg_0948;
    68: op1_10_in19 = imem01_in[123:120];
    69: op1_10_in19 = reg_0290;
    70: op1_10_in19 = reg_0716;
    72: op1_10_in19 = reg_0282;
    73: op1_10_in19 = imem07_in[83:80];
    74: op1_10_in19 = reg_0391;
    76: op1_10_in19 = reg_1023;
    77: op1_10_in19 = reg_0876;
    78: op1_10_in19 = reg_0516;
    79: op1_10_in19 = reg_0055;
    80: op1_10_in19 = reg_0022;
    81: op1_10_in19 = imem07_in[71:68];
    82: op1_10_in19 = reg_0229;
    83: op1_10_in19 = reg_0268;
    84: op1_10_in19 = reg_0459;
    85: op1_10_in19 = imem06_in[63:60];
    88: op1_10_in19 = reg_0945;
    89: op1_10_in19 = reg_0859;
    90: op1_10_in19 = reg_0129;
    91: op1_10_in19 = reg_0143;
    92: op1_10_in19 = reg_0426;
    94: op1_10_in19 = reg_0369;
    95: op1_10_in19 = reg_1014;
    96: op1_10_in19 = reg_0232;
    default: op1_10_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv19 = 1;
    6: op1_10_inv19 = 1;
    7: op1_10_inv19 = 1;
    8: op1_10_inv19 = 1;
    10: op1_10_inv19 = 1;
    11: op1_10_inv19 = 1;
    14: op1_10_inv19 = 1;
    17: op1_10_inv19 = 1;
    19: op1_10_inv19 = 1;
    20: op1_10_inv19 = 1;
    24: op1_10_inv19 = 1;
    25: op1_10_inv19 = 1;
    29: op1_10_inv19 = 1;
    31: op1_10_inv19 = 1;
    34: op1_10_inv19 = 1;
    35: op1_10_inv19 = 1;
    38: op1_10_inv19 = 1;
    40: op1_10_inv19 = 1;
    44: op1_10_inv19 = 1;
    45: op1_10_inv19 = 1;
    46: op1_10_inv19 = 1;
    49: op1_10_inv19 = 1;
    50: op1_10_inv19 = 1;
    51: op1_10_inv19 = 1;
    52: op1_10_inv19 = 1;
    53: op1_10_inv19 = 1;
    54: op1_10_inv19 = 1;
    56: op1_10_inv19 = 1;
    63: op1_10_inv19 = 1;
    64: op1_10_inv19 = 1;
    68: op1_10_inv19 = 1;
    70: op1_10_inv19 = 1;
    73: op1_10_inv19 = 1;
    74: op1_10_inv19 = 1;
    82: op1_10_inv19 = 1;
    83: op1_10_inv19 = 1;
    90: op1_10_inv19 = 1;
    92: op1_10_inv19 = 1;
    93: op1_10_inv19 = 1;
    94: op1_10_inv19 = 1;
    default: op1_10_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in20 = imem01_in[51:48];
    6: op1_10_in20 = reg_0197;
    7: op1_10_in20 = reg_0374;
    8: op1_10_in20 = reg_0616;
    9: op1_10_in20 = reg_0508;
    10: op1_10_in20 = imem07_in[43:40];
    11: op1_10_in20 = reg_0569;
    12: op1_10_in20 = reg_0419;
    13: op1_10_in20 = reg_0303;
    14: op1_10_in20 = reg_0144;
    15: op1_10_in20 = reg_0708;
    16: op1_10_in20 = reg_0084;
    17: op1_10_in20 = imem05_in[19:16];
    18: op1_10_in20 = reg_0085;
    19: op1_10_in20 = reg_0552;
    20: op1_10_in20 = reg_0330;
    21: op1_10_in20 = reg_0960;
    22: op1_10_in20 = imem01_in[55:52];
    23: op1_10_in20 = reg_0226;
    24: op1_10_in20 = reg_0196;
    25: op1_10_in20 = reg_0086;
    26: op1_10_in20 = reg_0723;
    27: op1_10_in20 = reg_0268;
    28: op1_10_in20 = reg_1009;
    29: op1_10_in20 = reg_0103;
    30: op1_10_in20 = reg_0648;
    31: op1_10_in20 = imem05_in[7:4];
    32: op1_10_in20 = reg_0707;
    34: op1_10_in20 = reg_0310;
    35: op1_10_in20 = reg_0388;
    36: op1_10_in20 = reg_0390;
    38: op1_10_in20 = reg_0383;
    39: op1_10_in20 = reg_0235;
    40: op1_10_in20 = reg_0667;
    41: op1_10_in20 = reg_0077;
    42: op1_10_in20 = imem07_in[119:116];
    43: op1_10_in20 = reg_0182;
    44: op1_10_in20 = reg_0786;
    45: op1_10_in20 = reg_0965;
    46: op1_10_in20 = imem06_in[103:100];
    47: op1_10_in20 = reg_0223;
    48: op1_10_in20 = reg_0525;
    49: op1_10_in20 = imem06_in[43:40];
    50: op1_10_in20 = imem04_in[55:52];
    51: op1_10_in20 = imem03_in[67:64];
    52: op1_10_in20 = imem01_in[91:88];
    53: op1_10_in20 = reg_0389;
    54: op1_10_in20 = reg_0872;
    55: op1_10_in20 = reg_0961;
    56: op1_10_in20 = reg_0611;
    82: op1_10_in20 = reg_0611;
    57: op1_10_in20 = reg_0446;
    58: op1_10_in20 = reg_0000;
    59: op1_10_in20 = reg_0728;
    60: op1_10_in20 = reg_0726;
    70: op1_10_in20 = reg_0726;
    62: op1_10_in20 = imem01_in[35:32];
    63: op1_10_in20 = reg_0536;
    64: op1_10_in20 = reg_0066;
    65: op1_10_in20 = reg_0493;
    66: op1_10_in20 = reg_1029;
    67: op1_10_in20 = reg_0865;
    68: op1_10_in20 = reg_0928;
    69: op1_10_in20 = reg_0873;
    72: op1_10_in20 = reg_0932;
    73: op1_10_in20 = imem07_in[87:84];
    81: op1_10_in20 = imem07_in[87:84];
    74: op1_10_in20 = reg_0021;
    76: op1_10_in20 = reg_0592;
    77: op1_10_in20 = reg_0049;
    89: op1_10_in20 = reg_0049;
    78: op1_10_in20 = reg_0054;
    79: op1_10_in20 = reg_0778;
    80: op1_10_in20 = imem07_in[35:32];
    83: op1_10_in20 = reg_0078;
    84: op1_10_in20 = reg_0191;
    85: op1_10_in20 = imem06_in[91:88];
    87: op1_10_in20 = imem03_in[15:12];
    88: op1_10_in20 = reg_0741;
    90: op1_10_in20 = reg_0130;
    91: op1_10_in20 = reg_0139;
    92: op1_10_in20 = reg_0161;
    93: op1_10_in20 = reg_0368;
    94: op1_10_in20 = imem01_in[27:24];
    95: op1_10_in20 = reg_0829;
    96: op1_10_in20 = reg_0111;
    default: op1_10_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv20 = 1;
    6: op1_10_inv20 = 1;
    14: op1_10_inv20 = 1;
    19: op1_10_inv20 = 1;
    20: op1_10_inv20 = 1;
    23: op1_10_inv20 = 1;
    25: op1_10_inv20 = 1;
    26: op1_10_inv20 = 1;
    27: op1_10_inv20 = 1;
    28: op1_10_inv20 = 1;
    29: op1_10_inv20 = 1;
    30: op1_10_inv20 = 1;
    31: op1_10_inv20 = 1;
    34: op1_10_inv20 = 1;
    35: op1_10_inv20 = 1;
    36: op1_10_inv20 = 1;
    38: op1_10_inv20 = 1;
    39: op1_10_inv20 = 1;
    42: op1_10_inv20 = 1;
    45: op1_10_inv20 = 1;
    46: op1_10_inv20 = 1;
    47: op1_10_inv20 = 1;
    52: op1_10_inv20 = 1;
    53: op1_10_inv20 = 1;
    54: op1_10_inv20 = 1;
    58: op1_10_inv20 = 1;
    63: op1_10_inv20 = 1;
    65: op1_10_inv20 = 1;
    67: op1_10_inv20 = 1;
    68: op1_10_inv20 = 1;
    69: op1_10_inv20 = 1;
    73: op1_10_inv20 = 1;
    74: op1_10_inv20 = 1;
    77: op1_10_inv20 = 1;
    78: op1_10_inv20 = 1;
    79: op1_10_inv20 = 1;
    81: op1_10_inv20 = 1;
    82: op1_10_inv20 = 1;
    83: op1_10_inv20 = 1;
    84: op1_10_inv20 = 1;
    85: op1_10_inv20 = 1;
    87: op1_10_inv20 = 1;
    88: op1_10_inv20 = 1;
    89: op1_10_inv20 = 1;
    90: op1_10_inv20 = 1;
    92: op1_10_inv20 = 1;
    93: op1_10_inv20 = 1;
    95: op1_10_inv20 = 1;
    96: op1_10_inv20 = 1;
    default: op1_10_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in21 = imem01_in[91:88];
    6: op1_10_in21 = imem01_in[75:72];
    22: op1_10_in21 = imem01_in[75:72];
    7: op1_10_in21 = reg_0986;
    8: op1_10_in21 = reg_0626;
    9: op1_10_in21 = reg_0233;
    10: op1_10_in21 = imem07_in[51:48];
    11: op1_10_in21 = reg_0591;
    12: op1_10_in21 = reg_0437;
    13: op1_10_in21 = reg_0281;
    14: op1_10_in21 = imem06_in[19:16];
    15: op1_10_in21 = reg_0715;
    16: op1_10_in21 = reg_0087;
    17: op1_10_in21 = imem05_in[23:20];
    18: op1_10_in21 = reg_0086;
    53: op1_10_in21 = reg_0086;
    19: op1_10_in21 = reg_0537;
    20: op1_10_in21 = reg_0346;
    21: op1_10_in21 = reg_0813;
    23: op1_10_in21 = reg_0885;
    24: op1_10_in21 = reg_0192;
    25: op1_10_in21 = imem03_in[27:24];
    26: op1_10_in21 = reg_0703;
    27: op1_10_in21 = reg_0071;
    28: op1_10_in21 = reg_0539;
    92: op1_10_in21 = reg_0539;
    29: op1_10_in21 = reg_0111;
    30: op1_10_in21 = reg_0644;
    31: op1_10_in21 = imem05_in[43:40];
    32: op1_10_in21 = reg_0700;
    34: op1_10_in21 = reg_0884;
    35: op1_10_in21 = reg_0025;
    36: op1_10_in21 = reg_0753;
    38: op1_10_in21 = reg_0630;
    39: op1_10_in21 = reg_0218;
    44: op1_10_in21 = reg_0218;
    40: op1_10_in21 = reg_0096;
    41: op1_10_in21 = imem03_in[3:0];
    42: op1_10_in21 = reg_0723;
    43: op1_10_in21 = reg_0164;
    45: op1_10_in21 = reg_0827;
    46: op1_10_in21 = imem06_in[115:112];
    47: op1_10_in21 = reg_0242;
    48: op1_10_in21 = reg_0269;
    49: op1_10_in21 = imem06_in[83:80];
    50: op1_10_in21 = imem04_in[87:84];
    51: op1_10_in21 = imem03_in[79:76];
    52: op1_10_in21 = reg_0586;
    54: op1_10_in21 = reg_0009;
    55: op1_10_in21 = reg_0960;
    56: op1_10_in21 = reg_0782;
    57: op1_10_in21 = reg_0148;
    58: op1_10_in21 = reg_0660;
    85: op1_10_in21 = reg_0660;
    59: op1_10_in21 = reg_0702;
    60: op1_10_in21 = reg_0714;
    62: op1_10_in21 = imem01_in[39:36];
    63: op1_10_in21 = reg_0277;
    64: op1_10_in21 = reg_0064;
    65: op1_10_in21 = reg_0128;
    66: op1_10_in21 = reg_0348;
    67: op1_10_in21 = reg_1046;
    68: op1_10_in21 = reg_0936;
    69: op1_10_in21 = reg_0036;
    70: op1_10_in21 = reg_0725;
    72: op1_10_in21 = reg_0799;
    73: op1_10_in21 = reg_0716;
    74: op1_10_in21 = reg_1030;
    76: op1_10_in21 = reg_1035;
    77: op1_10_in21 = reg_0016;
    78: op1_10_in21 = reg_0007;
    79: op1_10_in21 = reg_0932;
    80: op1_10_in21 = imem07_in[39:36];
    81: op1_10_in21 = imem07_in[99:96];
    82: op1_10_in21 = reg_0619;
    83: op1_10_in21 = reg_0166;
    84: op1_10_in21 = reg_0187;
    87: op1_10_in21 = imem03_in[55:52];
    88: op1_10_in21 = reg_0144;
    89: op1_10_in21 = reg_0620;
    90: op1_10_in21 = reg_0831;
    91: op1_10_in21 = reg_0235;
    93: op1_10_in21 = reg_0225;
    94: op1_10_in21 = imem01_in[31:28];
    95: op1_10_in21 = reg_0875;
    96: op1_10_in21 = reg_0003;
    default: op1_10_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv21 = 1;
    7: op1_10_inv21 = 1;
    9: op1_10_inv21 = 1;
    13: op1_10_inv21 = 1;
    14: op1_10_inv21 = 1;
    15: op1_10_inv21 = 1;
    16: op1_10_inv21 = 1;
    18: op1_10_inv21 = 1;
    19: op1_10_inv21 = 1;
    20: op1_10_inv21 = 1;
    21: op1_10_inv21 = 1;
    22: op1_10_inv21 = 1;
    23: op1_10_inv21 = 1;
    27: op1_10_inv21 = 1;
    29: op1_10_inv21 = 1;
    31: op1_10_inv21 = 1;
    32: op1_10_inv21 = 1;
    34: op1_10_inv21 = 1;
    35: op1_10_inv21 = 1;
    39: op1_10_inv21 = 1;
    41: op1_10_inv21 = 1;
    42: op1_10_inv21 = 1;
    44: op1_10_inv21 = 1;
    45: op1_10_inv21 = 1;
    47: op1_10_inv21 = 1;
    49: op1_10_inv21 = 1;
    50: op1_10_inv21 = 1;
    51: op1_10_inv21 = 1;
    56: op1_10_inv21 = 1;
    57: op1_10_inv21 = 1;
    58: op1_10_inv21 = 1;
    59: op1_10_inv21 = 1;
    63: op1_10_inv21 = 1;
    65: op1_10_inv21 = 1;
    67: op1_10_inv21 = 1;
    68: op1_10_inv21 = 1;
    69: op1_10_inv21 = 1;
    70: op1_10_inv21 = 1;
    72: op1_10_inv21 = 1;
    73: op1_10_inv21 = 1;
    79: op1_10_inv21 = 1;
    81: op1_10_inv21 = 1;
    84: op1_10_inv21 = 1;
    88: op1_10_inv21 = 1;
    90: op1_10_inv21 = 1;
    93: op1_10_inv21 = 1;
    96: op1_10_inv21 = 1;
    default: op1_10_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in22 = imem01_in[95:92];
    6: op1_10_in22 = imem01_in[87:84];
    7: op1_10_in22 = reg_0981;
    8: op1_10_in22 = reg_0618;
    9: op1_10_in22 = reg_0242;
    10: op1_10_in22 = imem07_in[75:72];
    11: op1_10_in22 = reg_0584;
    12: op1_10_in22 = reg_0158;
    13: op1_10_in22 = reg_0305;
    14: op1_10_in22 = imem06_in[47:44];
    15: op1_10_in22 = reg_0706;
    16: op1_10_in22 = reg_0094;
    17: op1_10_in22 = imem05_in[59:56];
    18: op1_10_in22 = imem03_in[31:28];
    19: op1_10_in22 = imem04_in[19:16];
    20: op1_10_in22 = reg_0324;
    21: op1_10_in22 = reg_0147;
    22: op1_10_in22 = imem01_in[91:88];
    23: op1_10_in22 = reg_0904;
    24: op1_10_in22 = imem01_in[47:44];
    94: op1_10_in22 = imem01_in[47:44];
    25: op1_10_in22 = imem03_in[43:40];
    26: op1_10_in22 = reg_0712;
    59: op1_10_in22 = reg_0712;
    27: op1_10_in22 = reg_0063;
    83: op1_10_in22 = reg_0063;
    28: op1_10_in22 = reg_0932;
    29: op1_10_in22 = reg_0112;
    30: op1_10_in22 = reg_0039;
    31: op1_10_in22 = imem05_in[63:60];
    32: op1_10_in22 = reg_0429;
    34: op1_10_in22 = imem03_in[35:32];
    35: op1_10_in22 = reg_0404;
    36: op1_10_in22 = reg_0404;
    38: op1_10_in22 = reg_0631;
    39: op1_10_in22 = reg_0224;
    40: op1_10_in22 = reg_0037;
    41: op1_10_in22 = imem03_in[23:20];
    77: op1_10_in22 = imem03_in[23:20];
    42: op1_10_in22 = reg_0708;
    43: op1_10_in22 = reg_0170;
    44: op1_10_in22 = reg_0510;
    45: op1_10_in22 = reg_0229;
    46: op1_10_in22 = reg_0915;
    66: op1_10_in22 = reg_0915;
    47: op1_10_in22 = reg_0828;
    48: op1_10_in22 = reg_0873;
    49: op1_10_in22 = reg_0486;
    50: op1_10_in22 = imem04_in[95:92];
    51: op1_10_in22 = imem03_in[83:80];
    52: op1_10_in22 = reg_0786;
    53: op1_10_in22 = reg_0484;
    54: op1_10_in22 = reg_0676;
    55: op1_10_in22 = reg_0032;
    56: op1_10_in22 = reg_0632;
    57: op1_10_in22 = reg_0151;
    58: op1_10_in22 = reg_1019;
    60: op1_10_in22 = reg_0703;
    62: op1_10_in22 = imem01_in[55:52];
    63: op1_10_in22 = reg_0888;
    64: op1_10_in22 = reg_0809;
    72: op1_10_in22 = reg_0809;
    65: op1_10_in22 = reg_0129;
    67: op1_10_in22 = reg_0333;
    68: op1_10_in22 = reg_0870;
    69: op1_10_in22 = reg_0098;
    70: op1_10_in22 = reg_0702;
    73: op1_10_in22 = reg_0729;
    74: op1_10_in22 = reg_0611;
    76: op1_10_in22 = reg_0488;
    78: op1_10_in22 = reg_0086;
    79: op1_10_in22 = reg_0799;
    80: op1_10_in22 = imem07_in[47:44];
    81: op1_10_in22 = imem07_in[107:104];
    82: op1_10_in22 = reg_0857;
    84: op1_10_in22 = reg_0204;
    85: op1_10_in22 = reg_0691;
    87: op1_10_in22 = imem03_in[67:64];
    88: op1_10_in22 = imem06_in[19:16];
    89: op1_10_in22 = reg_0763;
    90: op1_10_in22 = reg_0970;
    91: op1_10_in22 = reg_0140;
    92: op1_10_in22 = reg_0185;
    93: op1_10_in22 = reg_1042;
    95: op1_10_in22 = reg_0616;
    96: op1_10_in22 = reg_0116;
    default: op1_10_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv22 = 1;
    7: op1_10_inv22 = 1;
    8: op1_10_inv22 = 1;
    10: op1_10_inv22 = 1;
    13: op1_10_inv22 = 1;
    14: op1_10_inv22 = 1;
    16: op1_10_inv22 = 1;
    18: op1_10_inv22 = 1;
    19: op1_10_inv22 = 1;
    20: op1_10_inv22 = 1;
    22: op1_10_inv22 = 1;
    24: op1_10_inv22 = 1;
    25: op1_10_inv22 = 1;
    29: op1_10_inv22 = 1;
    30: op1_10_inv22 = 1;
    31: op1_10_inv22 = 1;
    34: op1_10_inv22 = 1;
    35: op1_10_inv22 = 1;
    38: op1_10_inv22 = 1;
    39: op1_10_inv22 = 1;
    40: op1_10_inv22 = 1;
    42: op1_10_inv22 = 1;
    44: op1_10_inv22 = 1;
    45: op1_10_inv22 = 1;
    46: op1_10_inv22 = 1;
    50: op1_10_inv22 = 1;
    59: op1_10_inv22 = 1;
    60: op1_10_inv22 = 1;
    65: op1_10_inv22 = 1;
    66: op1_10_inv22 = 1;
    68: op1_10_inv22 = 1;
    70: op1_10_inv22 = 1;
    72: op1_10_inv22 = 1;
    73: op1_10_inv22 = 1;
    76: op1_10_inv22 = 1;
    78: op1_10_inv22 = 1;
    79: op1_10_inv22 = 1;
    81: op1_10_inv22 = 1;
    82: op1_10_inv22 = 1;
    83: op1_10_inv22 = 1;
    85: op1_10_inv22 = 1;
    89: op1_10_inv22 = 1;
    90: op1_10_inv22 = 1;
    91: op1_10_inv22 = 1;
    96: op1_10_inv22 = 1;
    default: op1_10_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in23 = imem01_in[111:108];
    6: op1_10_in23 = imem01_in[123:120];
    7: op1_10_in23 = reg_0975;
    8: op1_10_in23 = reg_0402;
    9: op1_10_in23 = reg_0247;
    39: op1_10_in23 = reg_0247;
    10: op1_10_in23 = imem07_in[119:116];
    11: op1_10_in23 = reg_0580;
    13: op1_10_in23 = reg_0277;
    14: op1_10_in23 = imem06_in[67:64];
    15: op1_10_in23 = reg_0422;
    16: op1_10_in23 = reg_0079;
    17: op1_10_in23 = imem05_in[107:104];
    18: op1_10_in23 = imem03_in[35:32];
    41: op1_10_in23 = imem03_in[35:32];
    19: op1_10_in23 = imem04_in[87:84];
    20: op1_10_in23 = reg_0365;
    21: op1_10_in23 = reg_0148;
    22: op1_10_in23 = imem01_in[95:92];
    23: op1_10_in23 = reg_0104;
    24: op1_10_in23 = imem01_in[99:96];
    25: op1_10_in23 = imem03_in[75:72];
    26: op1_10_in23 = reg_0729;
    27: op1_10_in23 = reg_0074;
    28: op1_10_in23 = reg_0050;
    29: op1_10_in23 = reg_0114;
    30: op1_10_in23 = reg_0096;
    31: op1_10_in23 = imem05_in[75:72];
    32: op1_10_in23 = reg_0432;
    72: op1_10_in23 = reg_0432;
    34: op1_10_in23 = imem03_in[39:36];
    35: op1_10_in23 = reg_0591;
    36: op1_10_in23 = reg_0018;
    38: op1_10_in23 = imem07_in[3:0];
    40: op1_10_in23 = reg_0772;
    42: op1_10_in23 = reg_0709;
    43: op1_10_in23 = reg_0157;
    44: op1_10_in23 = reg_0239;
    45: op1_10_in23 = reg_0825;
    46: op1_10_in23 = reg_0783;
    47: op1_10_in23 = reg_0249;
    48: op1_10_in23 = imem05_in[59:56];
    49: op1_10_in23 = reg_0781;
    50: op1_10_in23 = imem04_in[119:116];
    51: op1_10_in23 = imem03_in[103:100];
    52: op1_10_in23 = reg_0928;
    53: op1_10_in23 = imem03_in[3:0];
    54: op1_10_in23 = reg_0570;
    55: op1_10_in23 = reg_0023;
    56: op1_10_in23 = reg_0382;
    57: op1_10_in23 = reg_0142;
    58: op1_10_in23 = reg_0696;
    59: op1_10_in23 = reg_0724;
    60: op1_10_in23 = reg_0724;
    62: op1_10_in23 = reg_0933;
    63: op1_10_in23 = reg_0313;
    64: op1_10_in23 = reg_0243;
    65: op1_10_in23 = reg_0130;
    66: op1_10_in23 = reg_1028;
    67: op1_10_in23 = reg_0819;
    68: op1_10_in23 = reg_1036;
    69: op1_10_in23 = reg_0224;
    70: op1_10_in23 = reg_0703;
    73: op1_10_in23 = reg_0715;
    74: op1_10_in23 = reg_0699;
    76: op1_10_in23 = reg_0234;
    77: op1_10_in23 = imem03_in[31:28];
    78: op1_10_in23 = reg_0049;
    79: op1_10_in23 = reg_0067;
    80: op1_10_in23 = imem07_in[71:68];
    81: op1_10_in23 = imem07_in[115:112];
    82: op1_10_in23 = reg_0289;
    83: op1_10_in23 = reg_0654;
    84: op1_10_in23 = reg_0194;
    85: op1_10_in23 = reg_1018;
    87: op1_10_in23 = imem03_in[99:96];
    88: op1_10_in23 = imem06_in[35:32];
    89: op1_10_in23 = reg_0976;
    90: op1_10_in23 = reg_0145;
    91: op1_10_in23 = reg_0226;
    93: op1_10_in23 = reg_0488;
    94: op1_10_in23 = imem01_in[79:76];
    95: op1_10_in23 = reg_0962;
    96: op1_10_in23 = reg_0860;
    default: op1_10_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv23 = 1;
    6: op1_10_inv23 = 1;
    8: op1_10_inv23 = 1;
    9: op1_10_inv23 = 1;
    13: op1_10_inv23 = 1;
    14: op1_10_inv23 = 1;
    15: op1_10_inv23 = 1;
    19: op1_10_inv23 = 1;
    23: op1_10_inv23 = 1;
    26: op1_10_inv23 = 1;
    27: op1_10_inv23 = 1;
    28: op1_10_inv23 = 1;
    30: op1_10_inv23 = 1;
    31: op1_10_inv23 = 1;
    32: op1_10_inv23 = 1;
    35: op1_10_inv23 = 1;
    41: op1_10_inv23 = 1;
    43: op1_10_inv23 = 1;
    46: op1_10_inv23 = 1;
    47: op1_10_inv23 = 1;
    51: op1_10_inv23 = 1;
    53: op1_10_inv23 = 1;
    54: op1_10_inv23 = 1;
    56: op1_10_inv23 = 1;
    59: op1_10_inv23 = 1;
    60: op1_10_inv23 = 1;
    63: op1_10_inv23 = 1;
    64: op1_10_inv23 = 1;
    67: op1_10_inv23 = 1;
    70: op1_10_inv23 = 1;
    72: op1_10_inv23 = 1;
    73: op1_10_inv23 = 1;
    74: op1_10_inv23 = 1;
    80: op1_10_inv23 = 1;
    83: op1_10_inv23 = 1;
    84: op1_10_inv23 = 1;
    85: op1_10_inv23 = 1;
    87: op1_10_inv23 = 1;
    88: op1_10_inv23 = 1;
    89: op1_10_inv23 = 1;
    90: op1_10_inv23 = 1;
    93: op1_10_inv23 = 1;
    94: op1_10_inv23 = 1;
    95: op1_10_inv23 = 1;
    default: op1_10_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in24 = reg_0503;
    6: op1_10_in24 = imem01_in[127:124];
    7: op1_10_in24 = imem04_in[3:0];
    8: op1_10_in24 = reg_0356;
    9: op1_10_in24 = reg_0236;
    10: op1_10_in24 = reg_0704;
    11: op1_10_in24 = reg_0576;
    13: op1_10_in24 = reg_0276;
    14: op1_10_in24 = reg_0611;
    15: op1_10_in24 = reg_0433;
    16: op1_10_in24 = imem03_in[11:8];
    17: op1_10_in24 = imem05_in[111:108];
    18: op1_10_in24 = imem03_in[83:80];
    19: op1_10_in24 = imem04_in[99:96];
    20: op1_10_in24 = reg_0355;
    21: op1_10_in24 = reg_0136;
    22: op1_10_in24 = imem01_in[111:108];
    23: op1_10_in24 = reg_0120;
    24: op1_10_in24 = imem01_in[107:104];
    25: op1_10_in24 = imem03_in[99:96];
    26: op1_10_in24 = reg_0713;
    59: op1_10_in24 = reg_0713;
    27: op1_10_in24 = reg_0072;
    28: op1_10_in24 = reg_0537;
    29: op1_10_in24 = reg_0100;
    30: op1_10_in24 = reg_0318;
    31: op1_10_in24 = imem05_in[119:116];
    32: op1_10_in24 = reg_0436;
    34: op1_10_in24 = imem03_in[59:56];
    35: op1_10_in24 = reg_0029;
    36: op1_10_in24 = imem07_in[11:8];
    38: op1_10_in24 = imem07_in[71:68];
    39: op1_10_in24 = reg_0487;
    40: op1_10_in24 = reg_0007;
    41: op1_10_in24 = imem03_in[51:48];
    42: op1_10_in24 = reg_0441;
    44: op1_10_in24 = reg_0810;
    45: op1_10_in24 = reg_0896;
    46: op1_10_in24 = reg_0391;
    47: op1_10_in24 = reg_0501;
    48: op1_10_in24 = imem05_in[63:60];
    49: op1_10_in24 = reg_0595;
    50: op1_10_in24 = reg_0483;
    51: op1_10_in24 = imem03_in[107:104];
    52: op1_10_in24 = reg_0904;
    53: op1_10_in24 = imem03_in[47:44];
    54: op1_10_in24 = reg_0734;
    55: op1_10_in24 = reg_0448;
    56: op1_10_in24 = reg_0399;
    57: op1_10_in24 = reg_0146;
    58: op1_10_in24 = reg_0393;
    60: op1_10_in24 = reg_0708;
    62: op1_10_in24 = reg_0919;
    63: op1_10_in24 = reg_0799;
    64: op1_10_in24 = reg_0542;
    65: op1_10_in24 = reg_0140;
    66: op1_10_in24 = reg_0633;
    67: op1_10_in24 = reg_0142;
    68: op1_10_in24 = reg_0238;
    69: op1_10_in24 = reg_0643;
    70: op1_10_in24 = reg_0724;
    72: op1_10_in24 = reg_0444;
    73: op1_10_in24 = reg_0711;
    74: op1_10_in24 = reg_0289;
    76: op1_10_in24 = reg_0225;
    77: op1_10_in24 = imem03_in[55:52];
    78: op1_10_in24 = reg_0084;
    79: op1_10_in24 = reg_0064;
    80: op1_10_in24 = imem07_in[99:96];
    82: op1_10_in24 = reg_0381;
    83: op1_10_in24 = reg_0656;
    84: op1_10_in24 = reg_0196;
    85: op1_10_in24 = reg_1011;
    87: op1_10_in24 = reg_0345;
    88: op1_10_in24 = imem06_in[71:68];
    89: op1_10_in24 = reg_0558;
    90: op1_10_in24 = reg_0706;
    91: op1_10_in24 = reg_0259;
    93: op1_10_in24 = reg_1024;
    94: op1_10_in24 = imem01_in[103:100];
    95: op1_10_in24 = imem01_in[19:16];
    96: op1_10_in24 = reg_0109;
    default: op1_10_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv24 = 1;
    6: op1_10_inv24 = 1;
    7: op1_10_inv24 = 1;
    8: op1_10_inv24 = 1;
    10: op1_10_inv24 = 1;
    11: op1_10_inv24 = 1;
    14: op1_10_inv24 = 1;
    15: op1_10_inv24 = 1;
    16: op1_10_inv24 = 1;
    18: op1_10_inv24 = 1;
    21: op1_10_inv24 = 1;
    22: op1_10_inv24 = 1;
    23: op1_10_inv24 = 1;
    24: op1_10_inv24 = 1;
    27: op1_10_inv24 = 1;
    28: op1_10_inv24 = 1;
    31: op1_10_inv24 = 1;
    32: op1_10_inv24 = 1;
    36: op1_10_inv24 = 1;
    40: op1_10_inv24 = 1;
    42: op1_10_inv24 = 1;
    46: op1_10_inv24 = 1;
    47: op1_10_inv24 = 1;
    50: op1_10_inv24 = 1;
    53: op1_10_inv24 = 1;
    55: op1_10_inv24 = 1;
    56: op1_10_inv24 = 1;
    57: op1_10_inv24 = 1;
    58: op1_10_inv24 = 1;
    60: op1_10_inv24 = 1;
    62: op1_10_inv24 = 1;
    63: op1_10_inv24 = 1;
    65: op1_10_inv24 = 1;
    66: op1_10_inv24 = 1;
    67: op1_10_inv24 = 1;
    68: op1_10_inv24 = 1;
    72: op1_10_inv24 = 1;
    78: op1_10_inv24 = 1;
    80: op1_10_inv24 = 1;
    83: op1_10_inv24 = 1;
    84: op1_10_inv24 = 1;
    85: op1_10_inv24 = 1;
    87: op1_10_inv24 = 1;
    91: op1_10_inv24 = 1;
    94: op1_10_inv24 = 1;
    95: op1_10_inv24 = 1;
    default: op1_10_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in25 = reg_0517;
    6: op1_10_in25 = reg_0520;
    7: op1_10_in25 = imem04_in[71:68];
    8: op1_10_in25 = reg_0407;
    9: op1_10_in25 = reg_0248;
    10: op1_10_in25 = reg_0712;
    80: op1_10_in25 = reg_0712;
    11: op1_10_in25 = reg_0394;
    13: op1_10_in25 = reg_0291;
    14: op1_10_in25 = reg_0577;
    15: op1_10_in25 = reg_0423;
    32: op1_10_in25 = reg_0423;
    16: op1_10_in25 = imem03_in[31:28];
    17: op1_10_in25 = reg_0973;
    18: op1_10_in25 = imem03_in[103:100];
    41: op1_10_in25 = imem03_in[103:100];
    19: op1_10_in25 = reg_0059;
    20: op1_10_in25 = reg_0314;
    21: op1_10_in25 = reg_0152;
    91: op1_10_in25 = reg_0152;
    22: op1_10_in25 = imem01_in[127:124];
    23: op1_10_in25 = reg_0126;
    24: op1_10_in25 = imem01_in[123:120];
    25: op1_10_in25 = imem03_in[115:112];
    26: op1_10_in25 = reg_0425;
    27: op1_10_in25 = reg_0279;
    28: op1_10_in25 = reg_0763;
    29: op1_10_in25 = reg_0106;
    30: op1_10_in25 = reg_0886;
    31: op1_10_in25 = reg_0968;
    34: op1_10_in25 = imem03_in[91:88];
    35: op1_10_in25 = reg_0005;
    36: op1_10_in25 = imem07_in[31:28];
    38: op1_10_in25 = imem07_in[99:96];
    39: op1_10_in25 = reg_1039;
    44: op1_10_in25 = reg_1039;
    40: op1_10_in25 = reg_0814;
    42: op1_10_in25 = reg_0447;
    45: op1_10_in25 = reg_0819;
    46: op1_10_in25 = reg_0386;
    47: op1_10_in25 = reg_1041;
    48: op1_10_in25 = imem05_in[75:72];
    49: op1_10_in25 = reg_0889;
    50: op1_10_in25 = reg_0536;
    51: op1_10_in25 = reg_0571;
    52: op1_10_in25 = reg_0242;
    53: op1_10_in25 = reg_0357;
    54: op1_10_in25 = imem03_in[3:0];
    55: op1_10_in25 = reg_0136;
    56: op1_10_in25 = reg_0804;
    57: op1_10_in25 = reg_0156;
    58: op1_10_in25 = reg_0817;
    59: op1_10_in25 = reg_0002;
    60: op1_10_in25 = reg_0718;
    62: op1_10_in25 = reg_0274;
    63: op1_10_in25 = reg_0584;
    64: op1_10_in25 = reg_0295;
    65: op1_10_in25 = reg_0134;
    66: op1_10_in25 = reg_0955;
    67: op1_10_in25 = reg_0146;
    68: op1_10_in25 = reg_1037;
    69: op1_10_in25 = reg_0908;
    70: op1_10_in25 = reg_0708;
    72: op1_10_in25 = reg_0856;
    73: op1_10_in25 = reg_0727;
    74: op1_10_in25 = reg_0921;
    76: op1_10_in25 = reg_1043;
    77: op1_10_in25 = reg_0006;
    78: op1_10_in25 = reg_0310;
    79: op1_10_in25 = reg_0288;
    82: op1_10_in25 = reg_0220;
    83: op1_10_in25 = reg_0931;
    84: op1_10_in25 = reg_0205;
    85: op1_10_in25 = reg_0926;
    87: op1_10_in25 = reg_0760;
    88: op1_10_in25 = imem06_in[75:72];
    89: op1_10_in25 = reg_0662;
    90: op1_10_in25 = reg_0951;
    93: op1_10_in25 = imem01_in[51:48];
    94: op1_10_in25 = reg_0501;
    95: op1_10_in25 = imem01_in[63:60];
    96: op1_10_in25 = reg_0113;
    default: op1_10_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv25 = 1;
    9: op1_10_inv25 = 1;
    10: op1_10_inv25 = 1;
    11: op1_10_inv25 = 1;
    13: op1_10_inv25 = 1;
    14: op1_10_inv25 = 1;
    15: op1_10_inv25 = 1;
    16: op1_10_inv25 = 1;
    17: op1_10_inv25 = 1;
    18: op1_10_inv25 = 1;
    20: op1_10_inv25 = 1;
    23: op1_10_inv25 = 1;
    24: op1_10_inv25 = 1;
    27: op1_10_inv25 = 1;
    29: op1_10_inv25 = 1;
    31: op1_10_inv25 = 1;
    34: op1_10_inv25 = 1;
    36: op1_10_inv25 = 1;
    38: op1_10_inv25 = 1;
    40: op1_10_inv25 = 1;
    42: op1_10_inv25 = 1;
    45: op1_10_inv25 = 1;
    46: op1_10_inv25 = 1;
    47: op1_10_inv25 = 1;
    55: op1_10_inv25 = 1;
    56: op1_10_inv25 = 1;
    59: op1_10_inv25 = 1;
    62: op1_10_inv25 = 1;
    63: op1_10_inv25 = 1;
    64: op1_10_inv25 = 1;
    66: op1_10_inv25 = 1;
    67: op1_10_inv25 = 1;
    68: op1_10_inv25 = 1;
    70: op1_10_inv25 = 1;
    72: op1_10_inv25 = 1;
    73: op1_10_inv25 = 1;
    77: op1_10_inv25 = 1;
    79: op1_10_inv25 = 1;
    83: op1_10_inv25 = 1;
    84: op1_10_inv25 = 1;
    90: op1_10_inv25 = 1;
    93: op1_10_inv25 = 1;
    94: op1_10_inv25 = 1;
    95: op1_10_inv25 = 1;
    default: op1_10_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in26 = reg_0518;
    6: op1_10_in26 = reg_0521;
    7: op1_10_in26 = imem04_in[75:72];
    8: op1_10_in26 = reg_0405;
    9: op1_10_in26 = reg_0234;
    10: op1_10_in26 = reg_0729;
    11: op1_10_in26 = reg_0360;
    13: op1_10_in26 = reg_0297;
    14: op1_10_in26 = reg_0615;
    15: op1_10_in26 = reg_0439;
    16: op1_10_in26 = imem03_in[43:40];
    17: op1_10_in26 = reg_0944;
    18: op1_10_in26 = reg_0602;
    19: op1_10_in26 = reg_0283;
    20: op1_10_in26 = reg_0092;
    21: op1_10_in26 = imem06_in[79:76];
    22: op1_10_in26 = reg_1055;
    23: op1_10_in26 = imem02_in[27:24];
    24: op1_10_in26 = reg_0246;
    25: op1_10_in26 = reg_0598;
    26: op1_10_in26 = reg_0441;
    27: op1_10_in26 = reg_0058;
    28: op1_10_in26 = reg_0065;
    29: op1_10_in26 = reg_0101;
    30: op1_10_in26 = reg_0082;
    31: op1_10_in26 = reg_0961;
    32: op1_10_in26 = reg_0448;
    34: op1_10_in26 = imem03_in[107:104];
    35: op1_10_in26 = imem07_in[11:8];
    36: op1_10_in26 = imem07_in[43:40];
    38: op1_10_in26 = imem07_in[111:108];
    39: op1_10_in26 = reg_0500;
    40: op1_10_in26 = reg_0090;
    41: op1_10_in26 = reg_0394;
    69: op1_10_in26 = reg_0394;
    42: op1_10_in26 = reg_0434;
    44: op1_10_in26 = reg_1043;
    45: op1_10_in26 = reg_0147;
    46: op1_10_in26 = reg_0382;
    47: op1_10_in26 = reg_0116;
    48: op1_10_in26 = imem05_in[95:92];
    49: op1_10_in26 = reg_0348;
    50: op1_10_in26 = reg_0937;
    51: op1_10_in26 = reg_1050;
    52: op1_10_in26 = reg_1056;
    53: op1_10_in26 = reg_0327;
    54: op1_10_in26 = imem03_in[7:4];
    55: op1_10_in26 = reg_0144;
    56: op1_10_in26 = reg_0222;
    57: op1_10_in26 = reg_0387;
    58: op1_10_in26 = reg_1011;
    59: op1_10_in26 = reg_0303;
    60: op1_10_in26 = reg_0706;
    62: op1_10_in26 = reg_0249;
    63: op1_10_in26 = reg_0296;
    64: op1_10_in26 = imem05_in[7:4];
    65: op1_10_in26 = imem06_in[15:12];
    66: op1_10_in26 = imem07_in[3:0];
    67: op1_10_in26 = reg_0138;
    68: op1_10_in26 = reg_0216;
    70: op1_10_in26 = reg_0321;
    72: op1_10_in26 = reg_0531;
    73: op1_10_in26 = reg_0433;
    74: op1_10_in26 = reg_0612;
    76: op1_10_in26 = reg_1040;
    77: op1_10_in26 = reg_0099;
    78: op1_10_in26 = imem03_in[11:8];
    79: op1_10_in26 = reg_0432;
    80: op1_10_in26 = reg_0100;
    82: op1_10_in26 = reg_0383;
    83: op1_10_in26 = reg_0313;
    84: op1_10_in26 = reg_0197;
    85: op1_10_in26 = reg_0692;
    87: op1_10_in26 = reg_1007;
    88: op1_10_in26 = reg_0660;
    89: op1_10_in26 = reg_0823;
    90: op1_10_in26 = reg_0258;
    91: op1_10_in26 = reg_0956;
    93: op1_10_in26 = imem01_in[95:92];
    95: op1_10_in26 = imem01_in[95:92];
    94: op1_10_in26 = reg_0227;
    96: op1_10_in26 = reg_0821;
    default: op1_10_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv26 = 1;
    8: op1_10_inv26 = 1;
    9: op1_10_inv26 = 1;
    13: op1_10_inv26 = 1;
    14: op1_10_inv26 = 1;
    16: op1_10_inv26 = 1;
    18: op1_10_inv26 = 1;
    19: op1_10_inv26 = 1;
    22: op1_10_inv26 = 1;
    23: op1_10_inv26 = 1;
    24: op1_10_inv26 = 1;
    25: op1_10_inv26 = 1;
    27: op1_10_inv26 = 1;
    32: op1_10_inv26 = 1;
    34: op1_10_inv26 = 1;
    35: op1_10_inv26 = 1;
    38: op1_10_inv26 = 1;
    40: op1_10_inv26 = 1;
    44: op1_10_inv26 = 1;
    45: op1_10_inv26 = 1;
    46: op1_10_inv26 = 1;
    51: op1_10_inv26 = 1;
    52: op1_10_inv26 = 1;
    53: op1_10_inv26 = 1;
    54: op1_10_inv26 = 1;
    55: op1_10_inv26 = 1;
    57: op1_10_inv26 = 1;
    62: op1_10_inv26 = 1;
    65: op1_10_inv26 = 1;
    66: op1_10_inv26 = 1;
    67: op1_10_inv26 = 1;
    70: op1_10_inv26 = 1;
    72: op1_10_inv26 = 1;
    73: op1_10_inv26 = 1;
    76: op1_10_inv26 = 1;
    77: op1_10_inv26 = 1;
    82: op1_10_inv26 = 1;
    84: op1_10_inv26 = 1;
    88: op1_10_inv26 = 1;
    91: op1_10_inv26 = 1;
    93: op1_10_inv26 = 1;
    94: op1_10_inv26 = 1;
    default: op1_10_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in27 = reg_0506;
    6: op1_10_in27 = reg_0499;
    7: op1_10_in27 = imem04_in[79:76];
    8: op1_10_in27 = reg_0406;
    9: op1_10_in27 = reg_0245;
    10: op1_10_in27 = reg_0709;
    11: op1_10_in27 = reg_0343;
    13: op1_10_in27 = reg_0298;
    14: op1_10_in27 = reg_0348;
    15: op1_10_in27 = reg_0446;
    16: op1_10_in27 = imem03_in[51:48];
    17: op1_10_in27 = reg_0959;
    18: op1_10_in27 = reg_0572;
    19: op1_10_in27 = reg_0058;
    20: op1_10_in27 = reg_0095;
    21: op1_10_in27 = imem06_in[127:124];
    22: op1_10_in27 = reg_0766;
    23: op1_10_in27 = imem02_in[91:88];
    24: op1_10_in27 = reg_0735;
    25: op1_10_in27 = reg_0571;
    41: op1_10_in27 = reg_0571;
    26: op1_10_in27 = reg_0422;
    27: op1_10_in27 = reg_0056;
    28: op1_10_in27 = reg_0076;
    29: op1_10_in27 = reg_0115;
    30: op1_10_in27 = reg_0516;
    31: op1_10_in27 = reg_0972;
    32: op1_10_in27 = reg_0431;
    34: op1_10_in27 = reg_0940;
    35: op1_10_in27 = imem07_in[63:60];
    36: op1_10_in27 = imem07_in[59:56];
    38: op1_10_in27 = imem07_in[115:112];
    39: op1_10_in27 = reg_1041;
    40: op1_10_in27 = reg_0291;
    42: op1_10_in27 = reg_0440;
    44: op1_10_in27 = reg_0616;
    45: op1_10_in27 = reg_0136;
    46: op1_10_in27 = reg_0243;
    47: op1_10_in27 = reg_0104;
    48: op1_10_in27 = reg_0957;
    49: op1_10_in27 = reg_0344;
    50: op1_10_in27 = reg_0277;
    51: op1_10_in27 = reg_0357;
    77: op1_10_in27 = reg_0357;
    52: op1_10_in27 = reg_1045;
    53: op1_10_in27 = reg_0874;
    54: op1_10_in27 = imem03_in[23:20];
    55: op1_10_in27 = imem06_in[7:4];
    56: op1_10_in27 = reg_0609;
    57: op1_10_in27 = reg_0915;
    58: op1_10_in27 = reg_0229;
    59: op1_10_in27 = reg_0325;
    60: op1_10_in27 = reg_0700;
    62: op1_10_in27 = reg_0607;
    63: op1_10_in27 = reg_0288;
    64: op1_10_in27 = imem05_in[39:36];
    65: op1_10_in27 = imem06_in[47:44];
    66: op1_10_in27 = imem07_in[7:4];
    67: op1_10_in27 = reg_0153;
    68: op1_10_in27 = reg_0902;
    69: op1_10_in27 = reg_0368;
    70: op1_10_in27 = reg_0419;
    72: op1_10_in27 = imem05_in[7:4];
    73: op1_10_in27 = reg_0428;
    74: op1_10_in27 = reg_0017;
    76: op1_10_in27 = reg_0925;
    78: op1_10_in27 = imem03_in[19:16];
    79: op1_10_in27 = reg_0444;
    80: op1_10_in27 = reg_0563;
    82: op1_10_in27 = reg_0403;
    83: op1_10_in27 = imem04_in[3:0];
    84: op1_10_in27 = imem01_in[7:4];
    85: op1_10_in27 = reg_0028;
    87: op1_10_in27 = reg_0327;
    88: op1_10_in27 = reg_0696;
    89: op1_10_in27 = reg_0597;
    90: op1_10_in27 = reg_0490;
    91: op1_10_in27 = reg_0129;
    93: op1_10_in27 = imem01_in[107:104];
    94: op1_10_in27 = reg_0622;
    95: op1_10_in27 = reg_0003;
    96: op1_10_in27 = reg_0110;
    default: op1_10_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_10_inv27 = 1;
    17: op1_10_inv27 = 1;
    18: op1_10_inv27 = 1;
    20: op1_10_inv27 = 1;
    23: op1_10_inv27 = 1;
    26: op1_10_inv27 = 1;
    29: op1_10_inv27 = 1;
    30: op1_10_inv27 = 1;
    31: op1_10_inv27 = 1;
    34: op1_10_inv27 = 1;
    35: op1_10_inv27 = 1;
    38: op1_10_inv27 = 1;
    39: op1_10_inv27 = 1;
    40: op1_10_inv27 = 1;
    41: op1_10_inv27 = 1;
    44: op1_10_inv27 = 1;
    47: op1_10_inv27 = 1;
    48: op1_10_inv27 = 1;
    49: op1_10_inv27 = 1;
    50: op1_10_inv27 = 1;
    51: op1_10_inv27 = 1;
    54: op1_10_inv27 = 1;
    55: op1_10_inv27 = 1;
    57: op1_10_inv27 = 1;
    58: op1_10_inv27 = 1;
    60: op1_10_inv27 = 1;
    62: op1_10_inv27 = 1;
    66: op1_10_inv27 = 1;
    67: op1_10_inv27 = 1;
    69: op1_10_inv27 = 1;
    73: op1_10_inv27 = 1;
    77: op1_10_inv27 = 1;
    78: op1_10_inv27 = 1;
    79: op1_10_inv27 = 1;
    88: op1_10_inv27 = 1;
    89: op1_10_inv27 = 1;
    90: op1_10_inv27 = 1;
    94: op1_10_inv27 = 1;
    95: op1_10_inv27 = 1;
    default: op1_10_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in28 = reg_0507;
    6: op1_10_in28 = reg_0518;
    7: op1_10_in28 = imem04_in[107:104];
    8: op1_10_in28 = reg_0032;
    9: op1_10_in28 = reg_0238;
    10: op1_10_in28 = reg_0701;
    11: op1_10_in28 = reg_0319;
    13: op1_10_in28 = reg_0288;
    14: op1_10_in28 = reg_0332;
    15: op1_10_in28 = reg_0449;
    16: op1_10_in28 = imem03_in[91:88];
    17: op1_10_in28 = reg_0967;
    18: op1_10_in28 = reg_0592;
    19: op1_10_in28 = reg_0528;
    20: op1_10_in28 = reg_0098;
    21: op1_10_in28 = reg_0610;
    22: op1_10_in28 = reg_1056;
    23: op1_10_in28 = reg_0642;
    24: op1_10_in28 = reg_0766;
    25: op1_10_in28 = reg_0596;
    46: op1_10_in28 = reg_0596;
    26: op1_10_in28 = reg_0421;
    27: op1_10_in28 = reg_0043;
    28: op1_10_in28 = reg_0074;
    29: op1_10_in28 = reg_0121;
    30: op1_10_in28 = reg_0007;
    31: op1_10_in28 = reg_1021;
    32: op1_10_in28 = reg_0165;
    34: op1_10_in28 = reg_0535;
    35: op1_10_in28 = imem07_in[111:108];
    36: op1_10_in28 = imem07_in[71:68];
    38: op1_10_in28 = reg_0717;
    39: op1_10_in28 = reg_0124;
    44: op1_10_in28 = reg_0124;
    40: op1_10_in28 = imem03_in[3:0];
    41: op1_10_in28 = reg_0245;
    42: op1_10_in28 = reg_0442;
    45: op1_10_in28 = reg_0138;
    47: op1_10_in28 = reg_0114;
    48: op1_10_in28 = reg_0969;
    49: op1_10_in28 = reg_0042;
    50: op1_10_in28 = reg_0055;
    51: op1_10_in28 = reg_0398;
    52: op1_10_in28 = reg_0869;
    53: op1_10_in28 = reg_0923;
    54: op1_10_in28 = imem03_in[51:48];
    55: op1_10_in28 = imem06_in[19:16];
    56: op1_10_in28 = reg_1010;
    57: op1_10_in28 = reg_0856;
    63: op1_10_in28 = reg_0856;
    58: op1_10_in28 = reg_0735;
    59: op1_10_in28 = reg_0047;
    60: op1_10_in28 = reg_0361;
    62: op1_10_in28 = reg_0496;
    64: op1_10_in28 = imem05_in[51:48];
    65: op1_10_in28 = imem06_in[71:68];
    66: op1_10_in28 = imem07_in[23:20];
    67: op1_10_in28 = reg_0141;
    68: op1_10_in28 = reg_0737;
    69: op1_10_in28 = reg_0331;
    70: op1_10_in28 = reg_0353;
    72: op1_10_in28 = imem05_in[11:8];
    73: op1_10_in28 = reg_0174;
    74: op1_10_in28 = reg_0403;
    76: op1_10_in28 = reg_0832;
    77: op1_10_in28 = reg_0396;
    78: op1_10_in28 = imem03_in[71:68];
    79: op1_10_in28 = reg_0360;
    80: op1_10_in28 = reg_0727;
    82: op1_10_in28 = reg_0095;
    83: op1_10_in28 = imem04_in[15:12];
    84: op1_10_in28 = imem01_in[11:8];
    85: op1_10_in28 = reg_0534;
    87: op1_10_in28 = reg_0322;
    88: op1_10_in28 = reg_0244;
    89: op1_10_in28 = reg_0385;
    90: op1_10_in28 = imem06_in[39:36];
    91: op1_10_in28 = reg_0437;
    93: op1_10_in28 = imem01_in[119:116];
    94: op1_10_in28 = reg_1038;
    95: op1_10_in28 = reg_1053;
    96: op1_10_in28 = imem02_in[3:0];
    default: op1_10_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_10_inv28 = 1;
    9: op1_10_inv28 = 1;
    13: op1_10_inv28 = 1;
    14: op1_10_inv28 = 1;
    16: op1_10_inv28 = 1;
    18: op1_10_inv28 = 1;
    19: op1_10_inv28 = 1;
    20: op1_10_inv28 = 1;
    25: op1_10_inv28 = 1;
    28: op1_10_inv28 = 1;
    29: op1_10_inv28 = 1;
    32: op1_10_inv28 = 1;
    34: op1_10_inv28 = 1;
    35: op1_10_inv28 = 1;
    41: op1_10_inv28 = 1;
    46: op1_10_inv28 = 1;
    48: op1_10_inv28 = 1;
    49: op1_10_inv28 = 1;
    51: op1_10_inv28 = 1;
    52: op1_10_inv28 = 1;
    53: op1_10_inv28 = 1;
    55: op1_10_inv28 = 1;
    57: op1_10_inv28 = 1;
    58: op1_10_inv28 = 1;
    62: op1_10_inv28 = 1;
    63: op1_10_inv28 = 1;
    67: op1_10_inv28 = 1;
    68: op1_10_inv28 = 1;
    70: op1_10_inv28 = 1;
    78: op1_10_inv28 = 1;
    79: op1_10_inv28 = 1;
    82: op1_10_inv28 = 1;
    83: op1_10_inv28 = 1;
    85: op1_10_inv28 = 1;
    87: op1_10_inv28 = 1;
    95: op1_10_inv28 = 1;
    96: op1_10_inv28 = 1;
    default: op1_10_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in29 = reg_0235;
    6: op1_10_in29 = reg_0515;
    7: op1_10_in29 = reg_0555;
    8: op1_10_in29 = reg_0029;
    9: op1_10_in29 = reg_0119;
    10: op1_10_in29 = reg_0706;
    11: op1_10_in29 = reg_0987;
    13: op1_10_in29 = reg_0059;
    14: op1_10_in29 = reg_0344;
    15: op1_10_in29 = reg_0431;
    16: op1_10_in29 = imem03_in[95:92];
    78: op1_10_in29 = imem03_in[95:92];
    17: op1_10_in29 = reg_0965;
    18: op1_10_in29 = reg_0597;
    19: op1_10_in29 = reg_0056;
    20: op1_10_in29 = reg_0094;
    21: op1_10_in29 = reg_0621;
    22: op1_10_in29 = reg_0220;
    23: op1_10_in29 = reg_0650;
    24: op1_10_in29 = reg_1056;
    25: op1_10_in29 = reg_0568;
    26: op1_10_in29 = reg_0449;
    27: op1_10_in29 = reg_0855;
    28: op1_10_in29 = reg_0738;
    29: op1_10_in29 = imem02_in[107:104];
    30: op1_10_in29 = reg_0758;
    31: op1_10_in29 = reg_0827;
    32: op1_10_in29 = reg_0162;
    34: op1_10_in29 = reg_0847;
    35: op1_10_in29 = reg_0721;
    36: op1_10_in29 = imem07_in[87:84];
    38: op1_10_in29 = reg_0725;
    39: op1_10_in29 = reg_0100;
    40: op1_10_in29 = imem03_in[35:32];
    41: op1_10_in29 = reg_0389;
    42: op1_10_in29 = reg_0435;
    44: op1_10_in29 = reg_0104;
    45: op1_10_in29 = reg_0155;
    46: op1_10_in29 = reg_0626;
    47: op1_10_in29 = imem02_in[7:4];
    96: op1_10_in29 = imem02_in[7:4];
    48: op1_10_in29 = reg_0960;
    49: op1_10_in29 = reg_0392;
    50: op1_10_in29 = reg_0050;
    51: op1_10_in29 = reg_0793;
    52: op1_10_in29 = reg_0604;
    53: op1_10_in29 = reg_0311;
    54: op1_10_in29 = imem03_in[67:64];
    55: op1_10_in29 = imem06_in[35:32];
    56: op1_10_in29 = imem07_in[83:80];
    57: op1_10_in29 = reg_0571;
    58: op1_10_in29 = imem06_in[19:16];
    59: op1_10_in29 = reg_0641;
    60: op1_10_in29 = reg_0419;
    62: op1_10_in29 = reg_0869;
    63: op1_10_in29 = imem05_in[15:12];
    64: op1_10_in29 = imem05_in[63:60];
    65: op1_10_in29 = reg_1019;
    66: op1_10_in29 = imem07_in[31:28];
    67: op1_10_in29 = reg_0140;
    68: op1_10_in29 = reg_1033;
    76: op1_10_in29 = reg_1033;
    69: op1_10_in29 = reg_0772;
    70: op1_10_in29 = reg_0024;
    72: op1_10_in29 = imem05_in[23:20];
    73: op1_10_in29 = reg_0179;
    74: op1_10_in29 = reg_0573;
    77: op1_10_in29 = reg_0661;
    79: op1_10_in29 = reg_0676;
    80: op1_10_in29 = reg_0002;
    82: op1_10_in29 = reg_0497;
    83: op1_10_in29 = imem04_in[23:20];
    84: op1_10_in29 = reg_0546;
    85: op1_10_in29 = reg_0591;
    87: op1_10_in29 = reg_0230;
    88: op1_10_in29 = reg_0391;
    89: op1_10_in29 = reg_1002;
    90: op1_10_in29 = imem06_in[47:44];
    91: op1_10_in29 = reg_0272;
    93: op1_10_in29 = reg_0232;
    94: op1_10_in29 = reg_0769;
    95: op1_10_in29 = reg_0733;
    default: op1_10_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv29 = 1;
    8: op1_10_inv29 = 1;
    9: op1_10_inv29 = 1;
    10: op1_10_inv29 = 1;
    13: op1_10_inv29 = 1;
    14: op1_10_inv29 = 1;
    17: op1_10_inv29 = 1;
    18: op1_10_inv29 = 1;
    21: op1_10_inv29 = 1;
    23: op1_10_inv29 = 1;
    24: op1_10_inv29 = 1;
    26: op1_10_inv29 = 1;
    28: op1_10_inv29 = 1;
    30: op1_10_inv29 = 1;
    34: op1_10_inv29 = 1;
    38: op1_10_inv29 = 1;
    41: op1_10_inv29 = 1;
    45: op1_10_inv29 = 1;
    46: op1_10_inv29 = 1;
    48: op1_10_inv29 = 1;
    50: op1_10_inv29 = 1;
    51: op1_10_inv29 = 1;
    57: op1_10_inv29 = 1;
    58: op1_10_inv29 = 1;
    59: op1_10_inv29 = 1;
    60: op1_10_inv29 = 1;
    63: op1_10_inv29 = 1;
    64: op1_10_inv29 = 1;
    66: op1_10_inv29 = 1;
    72: op1_10_inv29 = 1;
    74: op1_10_inv29 = 1;
    77: op1_10_inv29 = 1;
    79: op1_10_inv29 = 1;
    80: op1_10_inv29 = 1;
    83: op1_10_inv29 = 1;
    84: op1_10_inv29 = 1;
    85: op1_10_inv29 = 1;
    89: op1_10_inv29 = 1;
    90: op1_10_inv29 = 1;
    91: op1_10_inv29 = 1;
    default: op1_10_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_10_in30 = reg_0239;
    6: op1_10_in30 = reg_0233;
    7: op1_10_in30 = reg_0281;
    8: op1_10_in30 = imem07_in[3:0];
    9: op1_10_in30 = reg_0108;
    10: op1_10_in30 = reg_0425;
    11: op1_10_in30 = reg_0979;
    13: op1_10_in30 = reg_0046;
    14: op1_10_in30 = reg_0383;
    15: op1_10_in30 = reg_0180;
    16: op1_10_in30 = imem03_in[115:112];
    17: op1_10_in30 = reg_0215;
    48: op1_10_in30 = reg_0215;
    18: op1_10_in30 = reg_0395;
    19: op1_10_in30 = reg_0875;
    20: op1_10_in30 = reg_0093;
    21: op1_10_in30 = reg_0626;
    22: op1_10_in30 = reg_0234;
    23: op1_10_in30 = reg_0666;
    24: op1_10_in30 = reg_0507;
    25: op1_10_in30 = reg_0587;
    26: op1_10_in30 = reg_0444;
    27: op1_10_in30 = reg_0773;
    87: op1_10_in30 = reg_0773;
    28: op1_10_in30 = reg_0056;
    29: op1_10_in30 = imem02_in[111:108];
    30: op1_10_in30 = reg_0085;
    31: op1_10_in30 = reg_0252;
    32: op1_10_in30 = imem06_in[71:68];
    34: op1_10_in30 = reg_0311;
    35: op1_10_in30 = reg_0703;
    36: op1_10_in30 = reg_0728;
    38: op1_10_in30 = reg_0709;
    39: op1_10_in30 = reg_0110;
    40: op1_10_in30 = imem03_in[55:52];
    41: op1_10_in30 = reg_0765;
    51: op1_10_in30 = reg_0765;
    42: op1_10_in30 = reg_0175;
    60: op1_10_in30 = reg_0175;
    44: op1_10_in30 = reg_0126;
    45: op1_10_in30 = imem06_in[7:4];
    46: op1_10_in30 = reg_1010;
    47: op1_10_in30 = imem02_in[15:12];
    49: op1_10_in30 = reg_0017;
    50: op1_10_in30 = reg_0909;
    52: op1_10_in30 = reg_0830;
    53: op1_10_in30 = reg_0987;
    54: op1_10_in30 = imem03_in[87:84];
    55: op1_10_in30 = reg_0895;
    56: op1_10_in30 = reg_0730;
    57: op1_10_in30 = reg_0390;
    58: op1_10_in30 = imem06_in[63:60];
    59: op1_10_in30 = reg_0161;
    62: op1_10_in30 = reg_1037;
    63: op1_10_in30 = imem05_in[35:32];
    64: op1_10_in30 = imem05_in[67:64];
    65: op1_10_in30 = reg_0691;
    66: op1_10_in30 = imem07_in[43:40];
    67: op1_10_in30 = imem06_in[15:12];
    68: op1_10_in30 = reg_0112;
    69: op1_10_in30 = reg_0089;
    70: op1_10_in30 = reg_0172;
    72: op1_10_in30 = imem05_in[31:28];
    73: op1_10_in30 = reg_0162;
    74: op1_10_in30 = imem07_in[51:48];
    76: op1_10_in30 = reg_0273;
    77: op1_10_in30 = reg_0571;
    78: op1_10_in30 = reg_0345;
    79: op1_10_in30 = reg_0330;
    80: op1_10_in30 = reg_0406;
    82: op1_10_in30 = reg_0713;
    83: op1_10_in30 = imem04_in[79:76];
    84: op1_10_in30 = reg_1035;
    85: op1_10_in30 = reg_0270;
    88: op1_10_in30 = reg_0267;
    89: op1_10_in30 = reg_0996;
    90: op1_10_in30 = imem06_in[91:88];
    91: op1_10_in30 = reg_0706;
    93: op1_10_in30 = reg_1055;
    94: op1_10_in30 = reg_0283;
    95: op1_10_in30 = reg_0860;
    96: op1_10_in30 = imem02_in[79:76];
    default: op1_10_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv30 = 1;
    8: op1_10_inv30 = 1;
    9: op1_10_inv30 = 1;
    13: op1_10_inv30 = 1;
    15: op1_10_inv30 = 1;
    16: op1_10_inv30 = 1;
    17: op1_10_inv30 = 1;
    18: op1_10_inv30 = 1;
    19: op1_10_inv30 = 1;
    21: op1_10_inv30 = 1;
    22: op1_10_inv30 = 1;
    27: op1_10_inv30 = 1;
    28: op1_10_inv30 = 1;
    31: op1_10_inv30 = 1;
    32: op1_10_inv30 = 1;
    34: op1_10_inv30 = 1;
    35: op1_10_inv30 = 1;
    38: op1_10_inv30 = 1;
    39: op1_10_inv30 = 1;
    41: op1_10_inv30 = 1;
    44: op1_10_inv30 = 1;
    45: op1_10_inv30 = 1;
    46: op1_10_inv30 = 1;
    47: op1_10_inv30 = 1;
    48: op1_10_inv30 = 1;
    54: op1_10_inv30 = 1;
    57: op1_10_inv30 = 1;
    60: op1_10_inv30 = 1;
    62: op1_10_inv30 = 1;
    63: op1_10_inv30 = 1;
    64: op1_10_inv30 = 1;
    67: op1_10_inv30 = 1;
    68: op1_10_inv30 = 1;
    69: op1_10_inv30 = 1;
    73: op1_10_inv30 = 1;
    78: op1_10_inv30 = 1;
    79: op1_10_inv30 = 1;
    82: op1_10_inv30 = 1;
    89: op1_10_inv30 = 1;
    93: op1_10_inv30 = 1;
    95: op1_10_inv30 = 1;
    default: op1_10_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_10_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_10_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in00 = reg_0240;
    6: op1_11_in00 = reg_0236;
    7: op1_11_in00 = reg_0301;
    8: op1_11_in00 = imem07_in[7:4];
    9: op1_11_in00 = reg_0100;
    10: op1_11_in00 = imem00_in[59:56];
    11: op1_11_in00 = reg_0986;
    12: op1_11_in00 = imem00_in[19:16];
    13: op1_11_in00 = reg_0058;
    14: op1_11_in00 = reg_0367;
    15: op1_11_in00 = imem00_in[15:12];
    16: op1_11_in00 = imem03_in[119:116];
    17: op1_11_in00 = reg_0826;
    48: op1_11_in00 = reg_0826;
    18: op1_11_in00 = reg_0384;
    19: op1_11_in00 = reg_0855;
    20: op1_11_in00 = imem03_in[15:12];
    4: op1_11_in00 = imem07_in[55:52];
    21: op1_11_in00 = reg_0632;
    22: op1_11_in00 = reg_0245;
    23: op1_11_in00 = reg_0637;
    24: op1_11_in00 = reg_1042;
    25: op1_11_in00 = reg_0592;
    3: op1_11_in00 = imem07_in[99:96];
    26: op1_11_in00 = imem00_in[3:0];
    27: op1_11_in00 = imem05_in[63:60];
    28: op1_11_in00 = reg_0875;
    29: op1_11_in00 = imem02_in[115:112];
    30: op1_11_in00 = reg_0086;
    31: op1_11_in00 = reg_0229;
    2: op1_11_in00 = imem07_in[31:28];
    32: op1_11_in00 = imem00_in[7:4];
    33: op1_11_in00 = imem00_in[7:4];
    61: op1_11_in00 = imem00_in[7:4];
    86: op1_11_in00 = imem00_in[7:4];
    34: op1_11_in00 = reg_0807;
    35: op1_11_in00 = reg_0432;
    36: op1_11_in00 = reg_0430;
    37: op1_11_in00 = imem00_in[123:120];
    38: op1_11_in00 = reg_0707;
    39: op1_11_in00 = imem02_in[15:12];
    40: op1_11_in00 = imem03_in[59:56];
    41: op1_11_in00 = reg_0784;
    42: op1_11_in00 = reg_0181;
    70: op1_11_in00 = reg_0181;
    43: op1_11_in00 = imem00_in[39:36];
    92: op1_11_in00 = imem00_in[39:36];
    44: op1_11_in00 = imem02_in[7:4];
    45: op1_11_in00 = imem06_in[19:16];
    46: op1_11_in00 = imem07_in[103:100];
    47: op1_11_in00 = imem02_in[55:52];
    49: op1_11_in00 = reg_0626;
    50: op1_11_in00 = reg_0524;
    51: op1_11_in00 = reg_0370;
    52: op1_11_in00 = reg_0216;
    53: op1_11_in00 = reg_0991;
    54: op1_11_in00 = imem03_in[99:96];
    55: op1_11_in00 = reg_0220;
    56: op1_11_in00 = reg_0703;
    57: op1_11_in00 = imem06_in[55:52];
    58: op1_11_in00 = imem06_in[91:88];
    59: op1_11_in00 = reg_0162;
    60: op1_11_in00 = reg_0180;
    62: op1_11_in00 = reg_0616;
    63: op1_11_in00 = imem05_in[67:64];
    64: op1_11_in00 = imem05_in[71:68];
    65: op1_11_in00 = reg_1018;
    66: op1_11_in00 = imem07_in[51:48];
    67: op1_11_in00 = imem06_in[47:44];
    68: op1_11_in00 = reg_0103;
    69: op1_11_in00 = reg_0876;
    71: op1_11_in00 = imem00_in[51:48];
    72: op1_11_in00 = imem05_in[43:40];
    73: op1_11_in00 = reg_0166;
    74: op1_11_in00 = imem07_in[63:60];
    75: op1_11_in00 = imem00_in[75:72];
    76: op1_11_in00 = imem02_in[31:28];
    77: op1_11_in00 = reg_0397;
    78: op1_11_in00 = reg_0585;
    79: op1_11_in00 = reg_0530;
    80: op1_11_in00 = reg_0641;
    81: op1_11_in00 = imem00_in[23:20];
    82: op1_11_in00 = reg_0167;
    83: op1_11_in00 = imem04_in[87:84];
    84: op1_11_in00 = reg_0488;
    85: op1_11_in00 = reg_0485;
    87: op1_11_in00 = reg_0979;
    88: op1_11_in00 = reg_0692;
    89: op1_11_in00 = reg_1001;
    90: op1_11_in00 = reg_0660;
    91: op1_11_in00 = imem06_in[15:12];
    93: op1_11_in00 = reg_0003;
    94: op1_11_in00 = reg_0733;
    95: op1_11_in00 = reg_0113;
    96: op1_11_in00 = imem02_in[87:84];
    default: op1_11_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv00 = 1;
    9: op1_11_inv00 = 1;
    11: op1_11_inv00 = 1;
    12: op1_11_inv00 = 1;
    13: op1_11_inv00 = 1;
    15: op1_11_inv00 = 1;
    20: op1_11_inv00 = 1;
    4: op1_11_inv00 = 1;
    21: op1_11_inv00 = 1;
    24: op1_11_inv00 = 1;
    25: op1_11_inv00 = 1;
    26: op1_11_inv00 = 1;
    2: op1_11_inv00 = 1;
    36: op1_11_inv00 = 1;
    39: op1_11_inv00 = 1;
    40: op1_11_inv00 = 1;
    42: op1_11_inv00 = 1;
    47: op1_11_inv00 = 1;
    48: op1_11_inv00 = 1;
    50: op1_11_inv00 = 1;
    51: op1_11_inv00 = 1;
    52: op1_11_inv00 = 1;
    57: op1_11_inv00 = 1;
    59: op1_11_inv00 = 1;
    60: op1_11_inv00 = 1;
    61: op1_11_inv00 = 1;
    62: op1_11_inv00 = 1;
    64: op1_11_inv00 = 1;
    65: op1_11_inv00 = 1;
    66: op1_11_inv00 = 1;
    67: op1_11_inv00 = 1;
    68: op1_11_inv00 = 1;
    69: op1_11_inv00 = 1;
    72: op1_11_inv00 = 1;
    73: op1_11_inv00 = 1;
    74: op1_11_inv00 = 1;
    75: op1_11_inv00 = 1;
    76: op1_11_inv00 = 1;
    77: op1_11_inv00 = 1;
    78: op1_11_inv00 = 1;
    79: op1_11_inv00 = 1;
    80: op1_11_inv00 = 1;
    81: op1_11_inv00 = 1;
    84: op1_11_inv00 = 1;
    85: op1_11_inv00 = 1;
    88: op1_11_inv00 = 1;
    89: op1_11_inv00 = 1;
    92: op1_11_inv00 = 1;
    94: op1_11_inv00 = 1;
    96: op1_11_inv00 = 1;
    default: op1_11_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in01 = reg_0234;
    84: op1_11_in01 = reg_0234;
    6: op1_11_in01 = reg_0245;
    7: op1_11_in01 = reg_0294;
    8: op1_11_in01 = imem07_in[43:40];
    9: op1_11_in01 = reg_0101;
    10: op1_11_in01 = imem00_in[63:60];
    92: op1_11_in01 = imem00_in[63:60];
    11: op1_11_in01 = reg_0990;
    12: op1_11_in01 = imem00_in[27:24];
    61: op1_11_in01 = imem00_in[27:24];
    81: op1_11_in01 = imem00_in[27:24];
    86: op1_11_in01 = imem00_in[27:24];
    13: op1_11_in01 = imem05_in[7:4];
    28: op1_11_in01 = imem05_in[7:4];
    14: op1_11_in01 = reg_0026;
    15: op1_11_in01 = imem00_in[31:28];
    32: op1_11_in01 = imem00_in[31:28];
    16: op1_11_in01 = imem03_in[123:120];
    17: op1_11_in01 = reg_0835;
    18: op1_11_in01 = reg_0317;
    19: op1_11_in01 = imem05_in[55:52];
    72: op1_11_in01 = imem05_in[55:52];
    20: op1_11_in01 = imem03_in[39:36];
    4: op1_11_in01 = reg_0441;
    38: op1_11_in01 = reg_0441;
    21: op1_11_in01 = reg_0601;
    22: op1_11_in01 = reg_1042;
    23: op1_11_in01 = reg_0639;
    24: op1_11_in01 = reg_1043;
    25: op1_11_in01 = reg_0589;
    3: op1_11_in01 = imem07_in[111:108];
    26: op1_11_in01 = imem00_in[15:12];
    27: op1_11_in01 = imem05_in[75:72];
    29: op1_11_in01 = imem02_in[123:120];
    30: op1_11_in01 = reg_0310;
    69: op1_11_in01 = reg_0310;
    31: op1_11_in01 = reg_0785;
    2: op1_11_in01 = imem07_in[35:32];
    33: op1_11_in01 = imem00_in[71:68];
    43: op1_11_in01 = imem00_in[71:68];
    34: op1_11_in01 = reg_0312;
    35: op1_11_in01 = reg_0421;
    36: op1_11_in01 = reg_0433;
    37: op1_11_in01 = reg_0693;
    82: op1_11_in01 = reg_0693;
    39: op1_11_in01 = imem02_in[43:40];
    40: op1_11_in01 = imem03_in[83:80];
    41: op1_11_in01 = reg_0509;
    42: op1_11_in01 = reg_0160;
    44: op1_11_in01 = imem02_in[39:36];
    45: op1_11_in01 = imem06_in[39:36];
    46: op1_11_in01 = reg_0716;
    47: op1_11_in01 = imem02_in[59:56];
    48: op1_11_in01 = reg_0251;
    49: op1_11_in01 = reg_0622;
    50: op1_11_in01 = reg_0056;
    51: op1_11_in01 = reg_0373;
    52: op1_11_in01 = reg_0902;
    53: op1_11_in01 = reg_0996;
    54: op1_11_in01 = imem03_in[107:104];
    55: op1_11_in01 = reg_0371;
    56: op1_11_in01 = reg_0707;
    57: op1_11_in01 = imem06_in[83:80];
    58: op1_11_in01 = imem06_in[127:124];
    59: op1_11_in01 = reg_0177;
    60: op1_11_in01 = reg_0169;
    62: op1_11_in01 = reg_0925;
    63: op1_11_in01 = imem05_in[71:68];
    64: op1_11_in01 = imem05_in[103:100];
    65: op1_11_in01 = reg_0626;
    66: op1_11_in01 = imem07_in[71:68];
    74: op1_11_in01 = imem07_in[71:68];
    67: op1_11_in01 = reg_1019;
    68: op1_11_in01 = reg_0117;
    70: op1_11_in01 = reg_0162;
    71: op1_11_in01 = imem00_in[59:56];
    73: op1_11_in01 = reg_0168;
    75: op1_11_in01 = imem00_in[79:76];
    76: op1_11_in01 = imem02_in[35:32];
    77: op1_11_in01 = reg_0040;
    78: op1_11_in01 = reg_0046;
    79: op1_11_in01 = reg_0652;
    80: op1_11_in01 = reg_0502;
    83: op1_11_in01 = imem04_in[115:112];
    85: op1_11_in01 = reg_0018;
    87: op1_11_in01 = reg_0984;
    88: op1_11_in01 = reg_0814;
    89: op1_11_in01 = reg_0993;
    90: op1_11_in01 = reg_0694;
    91: op1_11_in01 = imem06_in[19:16];
    93: op1_11_in01 = reg_0555;
    94: op1_11_in01 = imem02_in[3:0];
    95: op1_11_in01 = imem02_in[23:20];
    96: op1_11_in01 = reg_0334;
    default: op1_11_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv01 = 1;
    6: op1_11_inv01 = 1;
    7: op1_11_inv01 = 1;
    8: op1_11_inv01 = 1;
    9: op1_11_inv01 = 1;
    12: op1_11_inv01 = 1;
    14: op1_11_inv01 = 1;
    15: op1_11_inv01 = 1;
    18: op1_11_inv01 = 1;
    19: op1_11_inv01 = 1;
    21: op1_11_inv01 = 1;
    22: op1_11_inv01 = 1;
    24: op1_11_inv01 = 1;
    27: op1_11_inv01 = 1;
    28: op1_11_inv01 = 1;
    30: op1_11_inv01 = 1;
    31: op1_11_inv01 = 1;
    2: op1_11_inv01 = 1;
    32: op1_11_inv01 = 1;
    33: op1_11_inv01 = 1;
    37: op1_11_inv01 = 1;
    38: op1_11_inv01 = 1;
    39: op1_11_inv01 = 1;
    42: op1_11_inv01 = 1;
    45: op1_11_inv01 = 1;
    49: op1_11_inv01 = 1;
    50: op1_11_inv01 = 1;
    56: op1_11_inv01 = 1;
    57: op1_11_inv01 = 1;
    59: op1_11_inv01 = 1;
    60: op1_11_inv01 = 1;
    61: op1_11_inv01 = 1;
    62: op1_11_inv01 = 1;
    64: op1_11_inv01 = 1;
    65: op1_11_inv01 = 1;
    66: op1_11_inv01 = 1;
    67: op1_11_inv01 = 1;
    69: op1_11_inv01 = 1;
    72: op1_11_inv01 = 1;
    74: op1_11_inv01 = 1;
    79: op1_11_inv01 = 1;
    81: op1_11_inv01 = 1;
    83: op1_11_inv01 = 1;
    86: op1_11_inv01 = 1;
    87: op1_11_inv01 = 1;
    90: op1_11_inv01 = 1;
    91: op1_11_inv01 = 1;
    93: op1_11_inv01 = 1;
    94: op1_11_inv01 = 1;
    95: op1_11_inv01 = 1;
    default: op1_11_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in02 = reg_0101;
    6: op1_11_in02 = reg_0221;
    7: op1_11_in02 = reg_0276;
    8: op1_11_in02 = imem07_in[51:48];
    9: op1_11_in02 = reg_0121;
    10: op1_11_in02 = imem00_in[71:68];
    11: op1_11_in02 = reg_1000;
    89: op1_11_in02 = reg_1000;
    12: op1_11_in02 = imem00_in[67:64];
    26: op1_11_in02 = imem00_in[67:64];
    13: op1_11_in02 = imem05_in[15:12];
    14: op1_11_in02 = reg_0800;
    15: op1_11_in02 = imem00_in[35:32];
    81: op1_11_in02 = imem00_in[35:32];
    16: op1_11_in02 = reg_0579;
    17: op1_11_in02 = reg_0827;
    18: op1_11_in02 = reg_0343;
    19: op1_11_in02 = imem05_in[103:100];
    20: op1_11_in02 = imem03_in[95:92];
    4: op1_11_in02 = reg_0432;
    21: op1_11_in02 = reg_0349;
    22: op1_11_in02 = reg_0230;
    23: op1_11_in02 = reg_0665;
    24: op1_11_in02 = reg_0216;
    25: op1_11_in02 = reg_0593;
    3: op1_11_in02 = imem07_in[115:112];
    27: op1_11_in02 = imem05_in[99:96];
    28: op1_11_in02 = imem05_in[19:16];
    29: op1_11_in02 = reg_0658;
    30: op1_11_in02 = imem03_in[27:24];
    31: op1_11_in02 = reg_0132;
    2: op1_11_in02 = imem07_in[43:40];
    32: op1_11_in02 = imem00_in[59:56];
    33: op1_11_in02 = imem00_in[75:72];
    34: op1_11_in02 = reg_0822;
    51: op1_11_in02 = reg_0822;
    35: op1_11_in02 = reg_0426;
    36: op1_11_in02 = reg_0440;
    37: op1_11_in02 = reg_0674;
    38: op1_11_in02 = reg_0429;
    39: op1_11_in02 = reg_0645;
    40: op1_11_in02 = imem03_in[103:100];
    41: op1_11_in02 = reg_0807;
    42: op1_11_in02 = reg_0158;
    43: op1_11_in02 = imem00_in[123:120];
    44: op1_11_in02 = imem02_in[51:48];
    45: op1_11_in02 = imem06_in[43:40];
    46: op1_11_in02 = reg_0725;
    47: op1_11_in02 = imem02_in[87:84];
    48: op1_11_in02 = reg_0825;
    49: op1_11_in02 = imem07_in[39:36];
    50: op1_11_in02 = reg_0014;
    52: op1_11_in02 = reg_0119;
    53: op1_11_in02 = reg_1001;
    87: op1_11_in02 = reg_1001;
    54: op1_11_in02 = reg_0847;
    55: op1_11_in02 = reg_0611;
    56: op1_11_in02 = reg_0427;
    57: op1_11_in02 = imem06_in[123:120];
    58: op1_11_in02 = reg_0628;
    59: op1_11_in02 = reg_0170;
    60: op1_11_in02 = reg_0168;
    61: op1_11_in02 = imem00_in[111:108];
    62: op1_11_in02 = reg_1033;
    63: op1_11_in02 = imem05_in[123:120];
    64: op1_11_in02 = reg_0042;
    65: op1_11_in02 = reg_0021;
    66: op1_11_in02 = imem07_in[79:76];
    67: op1_11_in02 = reg_0244;
    68: op1_11_in02 = reg_0821;
    69: op1_11_in02 = imem03_in[3:0];
    70: op1_11_in02 = reg_0159;
    71: op1_11_in02 = imem00_in[127:124];
    72: op1_11_in02 = imem05_in[71:68];
    73: op1_11_in02 = reg_0173;
    74: op1_11_in02 = imem07_in[103:100];
    75: op1_11_in02 = imem00_in[83:80];
    76: op1_11_in02 = imem02_in[39:36];
    77: op1_11_in02 = reg_0672;
    78: op1_11_in02 = reg_0396;
    79: op1_11_in02 = reg_0648;
    80: op1_11_in02 = reg_0868;
    82: op1_11_in02 = reg_0342;
    83: op1_11_in02 = imem04_in[127:124];
    84: op1_11_in02 = reg_0798;
    85: op1_11_in02 = reg_0403;
    86: op1_11_in02 = imem00_in[31:28];
    88: op1_11_in02 = reg_0630;
    90: op1_11_in02 = reg_0926;
    91: op1_11_in02 = imem06_in[27:24];
    92: op1_11_in02 = imem00_in[79:76];
    93: op1_11_in02 = reg_0115;
    94: op1_11_in02 = imem02_in[11:8];
    95: op1_11_in02 = reg_0255;
    96: op1_11_in02 = reg_0536;
    default: op1_11_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv02 = 1;
    7: op1_11_inv02 = 1;
    9: op1_11_inv02 = 1;
    12: op1_11_inv02 = 1;
    14: op1_11_inv02 = 1;
    16: op1_11_inv02 = 1;
    17: op1_11_inv02 = 1;
    18: op1_11_inv02 = 1;
    19: op1_11_inv02 = 1;
    20: op1_11_inv02 = 1;
    23: op1_11_inv02 = 1;
    25: op1_11_inv02 = 1;
    3: op1_11_inv02 = 1;
    26: op1_11_inv02 = 1;
    28: op1_11_inv02 = 1;
    32: op1_11_inv02 = 1;
    33: op1_11_inv02 = 1;
    34: op1_11_inv02 = 1;
    38: op1_11_inv02 = 1;
    39: op1_11_inv02 = 1;
    43: op1_11_inv02 = 1;
    44: op1_11_inv02 = 1;
    49: op1_11_inv02 = 1;
    55: op1_11_inv02 = 1;
    56: op1_11_inv02 = 1;
    57: op1_11_inv02 = 1;
    58: op1_11_inv02 = 1;
    60: op1_11_inv02 = 1;
    61: op1_11_inv02 = 1;
    62: op1_11_inv02 = 1;
    68: op1_11_inv02 = 1;
    70: op1_11_inv02 = 1;
    72: op1_11_inv02 = 1;
    77: op1_11_inv02 = 1;
    80: op1_11_inv02 = 1;
    81: op1_11_inv02 = 1;
    82: op1_11_inv02 = 1;
    83: op1_11_inv02 = 1;
    85: op1_11_inv02 = 1;
    88: op1_11_inv02 = 1;
    89: op1_11_inv02 = 1;
    92: op1_11_inv02 = 1;
    93: op1_11_inv02 = 1;
    95: op1_11_inv02 = 1;
    96: op1_11_inv02 = 1;
    default: op1_11_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in03 = reg_0659;
    6: op1_11_in03 = reg_0105;
    7: op1_11_in03 = reg_0295;
    8: op1_11_in03 = imem07_in[55:52];
    9: op1_11_in03 = reg_0650;
    10: op1_11_in03 = imem00_in[87:84];
    11: op1_11_in03 = imem04_in[11:8];
    12: op1_11_in03 = imem00_in[75:72];
    13: op1_11_in03 = imem05_in[35:32];
    14: op1_11_in03 = reg_0801;
    15: op1_11_in03 = imem00_in[83:80];
    33: op1_11_in03 = imem00_in[83:80];
    86: op1_11_in03 = imem00_in[83:80];
    16: op1_11_in03 = reg_0580;
    17: op1_11_in03 = reg_0258;
    18: op1_11_in03 = reg_0388;
    19: op1_11_in03 = reg_0963;
    20: op1_11_in03 = imem03_in[99:96];
    4: op1_11_in03 = reg_0445;
    21: op1_11_in03 = reg_0403;
    22: op1_11_in03 = reg_1033;
    23: op1_11_in03 = reg_0667;
    24: op1_11_in03 = reg_1035;
    25: op1_11_in03 = reg_0576;
    3: op1_11_in03 = imem07_in[127:124];
    26: op1_11_in03 = reg_0694;
    27: op1_11_in03 = reg_0966;
    28: op1_11_in03 = imem05_in[31:28];
    29: op1_11_in03 = reg_0664;
    39: op1_11_in03 = reg_0664;
    30: op1_11_in03 = imem03_in[51:48];
    31: op1_11_in03 = reg_0133;
    2: op1_11_in03 = imem07_in[87:84];
    32: op1_11_in03 = reg_0681;
    43: op1_11_in03 = reg_0681;
    34: op1_11_in03 = reg_0979;
    35: op1_11_in03 = reg_0423;
    36: op1_11_in03 = reg_0444;
    37: op1_11_in03 = reg_0680;
    38: op1_11_in03 = reg_0440;
    40: op1_11_in03 = imem03_in[127:124];
    41: op1_11_in03 = reg_0820;
    44: op1_11_in03 = imem02_in[75:72];
    45: op1_11_in03 = imem06_in[75:72];
    46: op1_11_in03 = reg_0724;
    47: op1_11_in03 = imem02_in[107:104];
    48: op1_11_in03 = reg_1046;
    49: op1_11_in03 = imem07_in[67:64];
    50: op1_11_in03 = reg_0276;
    51: op1_11_in03 = reg_0982;
    52: op1_11_in03 = reg_0120;
    53: op1_11_in03 = reg_0993;
    54: op1_11_in03 = reg_0874;
    55: op1_11_in03 = reg_0627;
    56: op1_11_in03 = reg_0431;
    57: op1_11_in03 = reg_0348;
    58: op1_11_in03 = reg_0780;
    59: op1_11_in03 = reg_0157;
    60: op1_11_in03 = reg_0157;
    61: op1_11_in03 = imem00_in[119:116];
    62: op1_11_in03 = reg_0273;
    63: op1_11_in03 = reg_0437;
    64: op1_11_in03 = reg_0967;
    65: op1_11_in03 = reg_0692;
    66: op1_11_in03 = reg_0728;
    67: op1_11_in03 = reg_0393;
    68: op1_11_in03 = reg_0110;
    93: op1_11_in03 = reg_0110;
    69: op1_11_in03 = imem03_in[11:8];
    70: op1_11_in03 = reg_0169;
    71: op1_11_in03 = reg_0519;
    72: op1_11_in03 = imem05_in[103:100];
    74: op1_11_in03 = reg_0719;
    75: op1_11_in03 = imem00_in[123:120];
    76: op1_11_in03 = imem02_in[55:52];
    77: op1_11_in03 = reg_0597;
    78: op1_11_in03 = reg_0662;
    79: op1_11_in03 = imem05_in[11:8];
    80: op1_11_in03 = reg_0024;
    81: op1_11_in03 = imem00_in[47:44];
    82: op1_11_in03 = reg_0711;
    83: op1_11_in03 = reg_0799;
    84: op1_11_in03 = reg_1037;
    85: op1_11_in03 = imem07_in[7:4];
    87: op1_11_in03 = reg_0980;
    88: op1_11_in03 = reg_0343;
    89: op1_11_in03 = imem04_in[15:12];
    90: op1_11_in03 = reg_0229;
    91: op1_11_in03 = imem06_in[35:32];
    92: op1_11_in03 = imem00_in[99:96];
    94: op1_11_in03 = imem02_in[15:12];
    95: op1_11_in03 = reg_0090;
    96: op1_11_in03 = reg_0075;
    default: op1_11_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv03 = 1;
    8: op1_11_inv03 = 1;
    9: op1_11_inv03 = 1;
    10: op1_11_inv03 = 1;
    14: op1_11_inv03 = 1;
    17: op1_11_inv03 = 1;
    19: op1_11_inv03 = 1;
    4: op1_11_inv03 = 1;
    21: op1_11_inv03 = 1;
    25: op1_11_inv03 = 1;
    31: op1_11_inv03 = 1;
    33: op1_11_inv03 = 1;
    35: op1_11_inv03 = 1;
    36: op1_11_inv03 = 1;
    38: op1_11_inv03 = 1;
    40: op1_11_inv03 = 1;
    41: op1_11_inv03 = 1;
    43: op1_11_inv03 = 1;
    44: op1_11_inv03 = 1;
    45: op1_11_inv03 = 1;
    46: op1_11_inv03 = 1;
    48: op1_11_inv03 = 1;
    57: op1_11_inv03 = 1;
    63: op1_11_inv03 = 1;
    69: op1_11_inv03 = 1;
    70: op1_11_inv03 = 1;
    74: op1_11_inv03 = 1;
    75: op1_11_inv03 = 1;
    76: op1_11_inv03 = 1;
    77: op1_11_inv03 = 1;
    78: op1_11_inv03 = 1;
    79: op1_11_inv03 = 1;
    82: op1_11_inv03 = 1;
    83: op1_11_inv03 = 1;
    85: op1_11_inv03 = 1;
    86: op1_11_inv03 = 1;
    87: op1_11_inv03 = 1;
    88: op1_11_inv03 = 1;
    95: op1_11_inv03 = 1;
    96: op1_11_inv03 = 1;
    default: op1_11_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in04 = reg_0334;
    6: op1_11_in04 = reg_0116;
    7: op1_11_in04 = reg_0307;
    8: op1_11_in04 = imem07_in[83:80];
    49: op1_11_in04 = imem07_in[83:80];
    9: op1_11_in04 = reg_0653;
    10: op1_11_in04 = reg_0679;
    11: op1_11_in04 = imem04_in[15:12];
    12: op1_11_in04 = imem00_in[95:92];
    33: op1_11_in04 = imem00_in[95:92];
    13: op1_11_in04 = imem05_in[67:64];
    14: op1_11_in04 = reg_1011;
    15: op1_11_in04 = reg_0682;
    16: op1_11_in04 = reg_0578;
    17: op1_11_in04 = reg_0147;
    18: op1_11_in04 = reg_0362;
    19: op1_11_in04 = reg_0970;
    20: op1_11_in04 = imem03_in[107:104];
    4: op1_11_in04 = reg_0437;
    35: op1_11_in04 = reg_0437;
    21: op1_11_in04 = reg_0406;
    22: op1_11_in04 = reg_1031;
    23: op1_11_in04 = reg_0325;
    24: op1_11_in04 = reg_0913;
    25: op1_11_in04 = reg_0391;
    3: op1_11_in04 = reg_0159;
    26: op1_11_in04 = reg_0688;
    27: op1_11_in04 = reg_0971;
    28: op1_11_in04 = imem05_in[59:56];
    29: op1_11_in04 = reg_0639;
    30: op1_11_in04 = imem03_in[71:68];
    31: op1_11_in04 = reg_0156;
    32: op1_11_in04 = reg_0676;
    34: op1_11_in04 = reg_0984;
    36: op1_11_in04 = reg_0442;
    37: op1_11_in04 = reg_0699;
    38: op1_11_in04 = reg_0169;
    39: op1_11_in04 = reg_0661;
    40: op1_11_in04 = reg_0317;
    41: op1_11_in04 = reg_0844;
    43: op1_11_in04 = reg_0696;
    44: op1_11_in04 = imem02_in[87:84];
    45: op1_11_in04 = imem06_in[83:80];
    46: op1_11_in04 = reg_0361;
    47: op1_11_in04 = reg_0654;
    48: op1_11_in04 = reg_0149;
    50: op1_11_in04 = reg_0401;
    51: op1_11_in04 = reg_0991;
    52: op1_11_in04 = reg_0121;
    53: op1_11_in04 = reg_0978;
    54: op1_11_in04 = reg_0370;
    55: op1_11_in04 = reg_0754;
    57: op1_11_in04 = reg_0914;
    58: op1_11_in04 = reg_0605;
    59: op1_11_in04 = reg_0158;
    60: op1_11_in04 = reg_0184;
    61: op1_11_in04 = reg_0001;
    75: op1_11_in04 = reg_0001;
    62: op1_11_in04 = reg_0113;
    63: op1_11_in04 = reg_0941;
    64: op1_11_in04 = reg_0972;
    65: op1_11_in04 = reg_0534;
    66: op1_11_in04 = reg_0704;
    67: op1_11_in04 = reg_0262;
    68: op1_11_in04 = imem02_in[7:4];
    69: op1_11_in04 = imem03_in[63:60];
    70: op1_11_in04 = reg_0182;
    71: op1_11_in04 = reg_0738;
    72: op1_11_in04 = imem05_in[119:116];
    74: op1_11_in04 = reg_0724;
    76: op1_11_in04 = imem02_in[67:64];
    77: op1_11_in04 = reg_0233;
    78: op1_11_in04 = reg_0038;
    79: op1_11_in04 = imem05_in[51:48];
    80: op1_11_in04 = reg_0183;
    81: op1_11_in04 = imem00_in[51:48];
    82: op1_11_in04 = reg_0705;
    83: op1_11_in04 = reg_0056;
    84: op1_11_in04 = reg_1053;
    85: op1_11_in04 = imem07_in[11:8];
    86: op1_11_in04 = imem00_in[107:104];
    87: op1_11_in04 = reg_0999;
    88: op1_11_in04 = reg_0822;
    89: op1_11_in04 = imem04_in[23:20];
    90: op1_11_in04 = reg_0889;
    91: op1_11_in04 = imem06_in[87:84];
    92: op1_11_in04 = imem00_in[115:112];
    93: op1_11_in04 = imem02_in[11:8];
    94: op1_11_in04 = imem02_in[39:36];
    95: op1_11_in04 = reg_0621;
    96: op1_11_in04 = reg_0543;
    default: op1_11_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv04 = 1;
    6: op1_11_inv04 = 1;
    8: op1_11_inv04 = 1;
    10: op1_11_inv04 = 1;
    12: op1_11_inv04 = 1;
    14: op1_11_inv04 = 1;
    15: op1_11_inv04 = 1;
    16: op1_11_inv04 = 1;
    17: op1_11_inv04 = 1;
    20: op1_11_inv04 = 1;
    21: op1_11_inv04 = 1;
    23: op1_11_inv04 = 1;
    26: op1_11_inv04 = 1;
    31: op1_11_inv04 = 1;
    32: op1_11_inv04 = 1;
    34: op1_11_inv04 = 1;
    35: op1_11_inv04 = 1;
    38: op1_11_inv04 = 1;
    40: op1_11_inv04 = 1;
    41: op1_11_inv04 = 1;
    47: op1_11_inv04 = 1;
    48: op1_11_inv04 = 1;
    49: op1_11_inv04 = 1;
    50: op1_11_inv04 = 1;
    51: op1_11_inv04 = 1;
    53: op1_11_inv04 = 1;
    54: op1_11_inv04 = 1;
    55: op1_11_inv04 = 1;
    57: op1_11_inv04 = 1;
    58: op1_11_inv04 = 1;
    59: op1_11_inv04 = 1;
    61: op1_11_inv04 = 1;
    62: op1_11_inv04 = 1;
    64: op1_11_inv04 = 1;
    66: op1_11_inv04 = 1;
    67: op1_11_inv04 = 1;
    69: op1_11_inv04 = 1;
    78: op1_11_inv04 = 1;
    79: op1_11_inv04 = 1;
    80: op1_11_inv04 = 1;
    82: op1_11_inv04 = 1;
    83: op1_11_inv04 = 1;
    84: op1_11_inv04 = 1;
    85: op1_11_inv04 = 1;
    86: op1_11_inv04 = 1;
    89: op1_11_inv04 = 1;
    91: op1_11_inv04 = 1;
    92: op1_11_inv04 = 1;
    93: op1_11_inv04 = 1;
    default: op1_11_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in05 = reg_0350;
    6: op1_11_in05 = reg_0119;
    7: op1_11_in05 = reg_0054;
    8: op1_11_in05 = imem07_in[119:116];
    9: op1_11_in05 = reg_0656;
    10: op1_11_in05 = reg_0688;
    11: op1_11_in05 = imem04_in[51:48];
    12: op1_11_in05 = reg_0693;
    13: op1_11_in05 = imem05_in[75:72];
    28: op1_11_in05 = imem05_in[75:72];
    14: op1_11_in05 = imem07_in[11:8];
    15: op1_11_in05 = reg_0681;
    16: op1_11_in05 = reg_0576;
    17: op1_11_in05 = reg_0149;
    18: op1_11_in05 = reg_0385;
    19: op1_11_in05 = reg_0950;
    20: op1_11_in05 = reg_0585;
    4: op1_11_in05 = reg_0420;
    21: op1_11_in05 = reg_0337;
    22: op1_11_in05 = reg_0913;
    23: op1_11_in05 = reg_0345;
    24: op1_11_in05 = reg_1017;
    25: op1_11_in05 = reg_0360;
    26: op1_11_in05 = reg_0465;
    27: op1_11_in05 = reg_0967;
    29: op1_11_in05 = reg_0651;
    30: op1_11_in05 = imem03_in[87:84];
    31: op1_11_in05 = imem06_in[11:8];
    32: op1_11_in05 = reg_0671;
    33: op1_11_in05 = reg_0697;
    34: op1_11_in05 = reg_0993;
    35: op1_11_in05 = reg_0431;
    36: op1_11_in05 = reg_0160;
    37: op1_11_in05 = reg_0470;
    38: op1_11_in05 = reg_0178;
    39: op1_11_in05 = reg_0842;
    40: op1_11_in05 = reg_0358;
    41: op1_11_in05 = reg_0985;
    43: op1_11_in05 = reg_0676;
    44: op1_11_in05 = imem02_in[111:108];
    45: op1_11_in05 = imem06_in[87:84];
    46: op1_11_in05 = reg_0744;
    47: op1_11_in05 = reg_0515;
    48: op1_11_in05 = reg_0135;
    49: op1_11_in05 = reg_0722;
    50: op1_11_in05 = reg_0815;
    51: op1_11_in05 = reg_0984;
    52: op1_11_in05 = reg_0768;
    53: op1_11_in05 = imem04_in[7:4];
    54: op1_11_in05 = reg_0833;
    55: op1_11_in05 = reg_0391;
    57: op1_11_in05 = reg_0741;
    58: op1_11_in05 = reg_0017;
    61: op1_11_in05 = reg_0683;
    62: op1_11_in05 = imem02_in[23:20];
    63: op1_11_in05 = reg_0835;
    64: op1_11_in05 = reg_0215;
    65: op1_11_in05 = reg_0297;
    66: op1_11_in05 = reg_0720;
    67: op1_11_in05 = reg_0817;
    68: op1_11_in05 = imem02_in[15:12];
    69: op1_11_in05 = imem03_in[67:64];
    70: op1_11_in05 = reg_0183;
    71: op1_11_in05 = reg_0663;
    72: op1_11_in05 = imem05_in[127:124];
    74: op1_11_in05 = reg_0422;
    75: op1_11_in05 = reg_0843;
    76: op1_11_in05 = imem02_in[87:84];
    77: op1_11_in05 = reg_0998;
    78: op1_11_in05 = reg_0239;
    79: op1_11_in05 = imem05_in[111:108];
    80: op1_11_in05 = reg_0185;
    81: op1_11_in05 = imem00_in[55:52];
    82: op1_11_in05 = reg_0438;
    83: op1_11_in05 = reg_0809;
    84: op1_11_in05 = reg_0860;
    85: op1_11_in05 = imem07_in[43:40];
    86: op1_11_in05 = imem00_in[111:108];
    87: op1_11_in05 = reg_0981;
    88: op1_11_in05 = reg_0121;
    89: op1_11_in05 = imem04_in[43:40];
    90: op1_11_in05 = reg_0692;
    91: op1_11_in05 = imem06_in[119:116];
    92: op1_11_in05 = reg_0386;
    93: op1_11_in05 = imem02_in[39:36];
    94: op1_11_in05 = imem02_in[43:40];
    95: op1_11_in05 = reg_0073;
    96: op1_11_in05 = reg_0090;
    default: op1_11_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_11_inv05 = 1;
    9: op1_11_inv05 = 1;
    10: op1_11_inv05 = 1;
    12: op1_11_inv05 = 1;
    13: op1_11_inv05 = 1;
    14: op1_11_inv05 = 1;
    15: op1_11_inv05 = 1;
    17: op1_11_inv05 = 1;
    18: op1_11_inv05 = 1;
    19: op1_11_inv05 = 1;
    24: op1_11_inv05 = 1;
    25: op1_11_inv05 = 1;
    27: op1_11_inv05 = 1;
    29: op1_11_inv05 = 1;
    34: op1_11_inv05 = 1;
    36: op1_11_inv05 = 1;
    37: op1_11_inv05 = 1;
    38: op1_11_inv05 = 1;
    40: op1_11_inv05 = 1;
    41: op1_11_inv05 = 1;
    45: op1_11_inv05 = 1;
    46: op1_11_inv05 = 1;
    47: op1_11_inv05 = 1;
    48: op1_11_inv05 = 1;
    49: op1_11_inv05 = 1;
    50: op1_11_inv05 = 1;
    51: op1_11_inv05 = 1;
    52: op1_11_inv05 = 1;
    58: op1_11_inv05 = 1;
    62: op1_11_inv05 = 1;
    64: op1_11_inv05 = 1;
    66: op1_11_inv05 = 1;
    67: op1_11_inv05 = 1;
    68: op1_11_inv05 = 1;
    69: op1_11_inv05 = 1;
    71: op1_11_inv05 = 1;
    72: op1_11_inv05 = 1;
    74: op1_11_inv05 = 1;
    76: op1_11_inv05 = 1;
    78: op1_11_inv05 = 1;
    79: op1_11_inv05 = 1;
    80: op1_11_inv05 = 1;
    81: op1_11_inv05 = 1;
    83: op1_11_inv05 = 1;
    84: op1_11_inv05 = 1;
    86: op1_11_inv05 = 1;
    88: op1_11_inv05 = 1;
    90: op1_11_inv05 = 1;
    95: op1_11_inv05 = 1;
    default: op1_11_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in06 = reg_0085;
    6: op1_11_in06 = reg_0106;
    7: op1_11_in06 = reg_0041;
    8: op1_11_in06 = reg_0719;
    49: op1_11_in06 = reg_0719;
    9: op1_11_in06 = reg_0639;
    47: op1_11_in06 = reg_0639;
    10: op1_11_in06 = reg_0699;
    11: op1_11_in06 = imem04_in[87:84];
    12: op1_11_in06 = reg_0694;
    91: op1_11_in06 = reg_0694;
    13: op1_11_in06 = imem05_in[115:112];
    28: op1_11_in06 = imem05_in[115:112];
    14: op1_11_in06 = imem07_in[75:72];
    15: op1_11_in06 = reg_0685;
    16: op1_11_in06 = reg_0388;
    17: op1_11_in06 = reg_0133;
    18: op1_11_in06 = reg_0396;
    19: op1_11_in06 = reg_0964;
    20: op1_11_in06 = reg_0362;
    4: op1_11_in06 = reg_0179;
    21: op1_11_in06 = reg_0800;
    22: op1_11_in06 = reg_1045;
    23: op1_11_in06 = reg_0339;
    24: op1_11_in06 = reg_0125;
    25: op1_11_in06 = reg_0361;
    26: op1_11_in06 = reg_0476;
    27: op1_11_in06 = reg_0957;
    29: op1_11_in06 = reg_0643;
    30: op1_11_in06 = imem03_in[95:92];
    31: op1_11_in06 = imem06_in[15:12];
    32: op1_11_in06 = reg_0668;
    33: op1_11_in06 = reg_0683;
    34: op1_11_in06 = reg_0980;
    35: op1_11_in06 = reg_0175;
    36: op1_11_in06 = reg_0163;
    37: op1_11_in06 = reg_0471;
    39: op1_11_in06 = reg_0039;
    40: op1_11_in06 = reg_0765;
    95: op1_11_in06 = reg_0765;
    41: op1_11_in06 = reg_0996;
    43: op1_11_in06 = reg_0689;
    44: op1_11_in06 = reg_0664;
    45: op1_11_in06 = imem06_in[115:112];
    46: op1_11_in06 = reg_0589;
    48: op1_11_in06 = reg_0139;
    50: op1_11_in06 = reg_0281;
    51: op1_11_in06 = reg_0989;
    52: op1_11_in06 = reg_0916;
    53: op1_11_in06 = imem04_in[27:24];
    54: op1_11_in06 = reg_0040;
    55: op1_11_in06 = reg_0264;
    57: op1_11_in06 = reg_0780;
    58: op1_11_in06 = reg_0633;
    61: op1_11_in06 = reg_0768;
    62: op1_11_in06 = imem02_in[55:52];
    63: op1_11_in06 = reg_0967;
    64: op1_11_in06 = reg_0259;
    65: op1_11_in06 = reg_0595;
    66: op1_11_in06 = reg_0702;
    67: op1_11_in06 = reg_0889;
    68: op1_11_in06 = imem02_in[23:20];
    69: op1_11_in06 = reg_0547;
    70: op1_11_in06 = reg_0173;
    71: op1_11_in06 = reg_0454;
    72: op1_11_in06 = reg_0970;
    74: op1_11_in06 = reg_0641;
    75: op1_11_in06 = reg_0738;
    76: op1_11_in06 = imem02_in[95:92];
    77: op1_11_in06 = reg_0979;
    78: op1_11_in06 = reg_0051;
    79: op1_11_in06 = reg_0707;
    81: op1_11_in06 = imem00_in[71:68];
    82: op1_11_in06 = reg_0725;
    83: op1_11_in06 = reg_0764;
    84: op1_11_in06 = reg_0877;
    85: op1_11_in06 = imem07_in[51:48];
    86: op1_11_in06 = reg_0001;
    87: op1_11_in06 = reg_0983;
    88: op1_11_in06 = reg_0220;
    89: op1_11_in06 = imem04_in[47:44];
    90: op1_11_in06 = reg_0630;
    92: op1_11_in06 = reg_0867;
    93: op1_11_in06 = imem02_in[43:40];
    94: op1_11_in06 = imem02_in[51:48];
    96: op1_11_in06 = reg_0642;
    default: op1_11_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv06 = 1;
    6: op1_11_inv06 = 1;
    8: op1_11_inv06 = 1;
    9: op1_11_inv06 = 1;
    10: op1_11_inv06 = 1;
    12: op1_11_inv06 = 1;
    14: op1_11_inv06 = 1;
    15: op1_11_inv06 = 1;
    16: op1_11_inv06 = 1;
    4: op1_11_inv06 = 1;
    21: op1_11_inv06 = 1;
    22: op1_11_inv06 = 1;
    24: op1_11_inv06 = 1;
    25: op1_11_inv06 = 1;
    26: op1_11_inv06 = 1;
    27: op1_11_inv06 = 1;
    28: op1_11_inv06 = 1;
    32: op1_11_inv06 = 1;
    34: op1_11_inv06 = 1;
    35: op1_11_inv06 = 1;
    36: op1_11_inv06 = 1;
    37: op1_11_inv06 = 1;
    44: op1_11_inv06 = 1;
    49: op1_11_inv06 = 1;
    50: op1_11_inv06 = 1;
    51: op1_11_inv06 = 1;
    52: op1_11_inv06 = 1;
    54: op1_11_inv06 = 1;
    58: op1_11_inv06 = 1;
    62: op1_11_inv06 = 1;
    65: op1_11_inv06 = 1;
    66: op1_11_inv06 = 1;
    72: op1_11_inv06 = 1;
    75: op1_11_inv06 = 1;
    78: op1_11_inv06 = 1;
    81: op1_11_inv06 = 1;
    82: op1_11_inv06 = 1;
    84: op1_11_inv06 = 1;
    86: op1_11_inv06 = 1;
    88: op1_11_inv06 = 1;
    89: op1_11_inv06 = 1;
    90: op1_11_inv06 = 1;
    92: op1_11_inv06 = 1;
    93: op1_11_inv06 = 1;
    94: op1_11_inv06 = 1;
    default: op1_11_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in07 = reg_0052;
    6: op1_11_in07 = reg_0101;
    7: op1_11_in07 = reg_0053;
    8: op1_11_in07 = reg_0713;
    9: op1_11_in07 = reg_0357;
    10: op1_11_in07 = reg_0476;
    11: op1_11_in07 = reg_0535;
    12: op1_11_in07 = reg_0676;
    13: op1_11_in07 = reg_0966;
    14: op1_11_in07 = imem07_in[103:100];
    15: op1_11_in07 = reg_0689;
    16: op1_11_in07 = reg_0369;
    17: op1_11_in07 = reg_0152;
    18: op1_11_in07 = reg_0374;
    25: op1_11_in07 = reg_0374;
    19: op1_11_in07 = reg_0961;
    20: op1_11_in07 = reg_0312;
    21: op1_11_in07 = reg_0753;
    22: op1_11_in07 = reg_1017;
    23: op1_11_in07 = reg_0355;
    24: op1_11_in07 = reg_0104;
    26: op1_11_in07 = reg_0480;
    27: op1_11_in07 = reg_0942;
    28: op1_11_in07 = reg_0962;
    29: op1_11_in07 = reg_0652;
    30: op1_11_in07 = imem03_in[123:120];
    31: op1_11_in07 = imem06_in[51:48];
    32: op1_11_in07 = reg_0687;
    33: op1_11_in07 = reg_0672;
    34: op1_11_in07 = reg_0978;
    35: op1_11_in07 = reg_0162;
    36: op1_11_in07 = reg_0183;
    37: op1_11_in07 = reg_0468;
    39: op1_11_in07 = reg_0330;
    40: op1_11_in07 = reg_0833;
    41: op1_11_in07 = reg_0980;
    43: op1_11_in07 = reg_0684;
    44: op1_11_in07 = reg_0661;
    69: op1_11_in07 = reg_0661;
    45: op1_11_in07 = reg_0624;
    46: op1_11_in07 = reg_0174;
    74: op1_11_in07 = reg_0174;
    47: op1_11_in07 = reg_0300;
    48: op1_11_in07 = reg_0140;
    49: op1_11_in07 = reg_0710;
    50: op1_11_in07 = reg_0899;
    51: op1_11_in07 = reg_0990;
    52: op1_11_in07 = reg_0095;
    53: op1_11_in07 = imem04_in[35:32];
    54: op1_11_in07 = reg_0784;
    55: op1_11_in07 = reg_0295;
    57: op1_11_in07 = reg_0241;
    58: op1_11_in07 = imem07_in[7:4];
    61: op1_11_in07 = reg_0900;
    62: op1_11_in07 = reg_0650;
    63: op1_11_in07 = reg_0254;
    64: op1_11_in07 = reg_0446;
    65: op1_11_in07 = reg_0781;
    66: op1_11_in07 = reg_0709;
    67: op1_11_in07 = reg_0297;
    68: op1_11_in07 = imem02_in[35:32];
    70: op1_11_in07 = reg_0184;
    71: op1_11_in07 = reg_0452;
    72: op1_11_in07 = reg_0693;
    75: op1_11_in07 = reg_0356;
    76: op1_11_in07 = reg_0750;
    77: op1_11_in07 = reg_0977;
    78: op1_11_in07 = reg_0376;
    79: op1_11_in07 = reg_0019;
    81: op1_11_in07 = reg_0843;
    82: op1_11_in07 = reg_0712;
    83: op1_11_in07 = reg_0061;
    84: op1_11_in07 = reg_0117;
    85: op1_11_in07 = imem07_in[59:56];
    86: op1_11_in07 = reg_0841;
    87: op1_11_in07 = imem04_in[83:80];
    88: op1_11_in07 = reg_0755;
    89: op1_11_in07 = imem04_in[51:48];
    90: op1_11_in07 = reg_0729;
    91: op1_11_in07 = reg_1019;
    92: op1_11_in07 = reg_0028;
    93: op1_11_in07 = imem02_in[83:80];
    94: op1_11_in07 = imem02_in[99:96];
    95: op1_11_in07 = reg_0423;
    96: op1_11_in07 = reg_0765;
    default: op1_11_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_11_inv07 = 1;
    9: op1_11_inv07 = 1;
    11: op1_11_inv07 = 1;
    14: op1_11_inv07 = 1;
    17: op1_11_inv07 = 1;
    18: op1_11_inv07 = 1;
    22: op1_11_inv07 = 1;
    25: op1_11_inv07 = 1;
    27: op1_11_inv07 = 1;
    28: op1_11_inv07 = 1;
    29: op1_11_inv07 = 1;
    31: op1_11_inv07 = 1;
    33: op1_11_inv07 = 1;
    36: op1_11_inv07 = 1;
    37: op1_11_inv07 = 1;
    39: op1_11_inv07 = 1;
    40: op1_11_inv07 = 1;
    41: op1_11_inv07 = 1;
    45: op1_11_inv07 = 1;
    46: op1_11_inv07 = 1;
    52: op1_11_inv07 = 1;
    53: op1_11_inv07 = 1;
    54: op1_11_inv07 = 1;
    57: op1_11_inv07 = 1;
    63: op1_11_inv07 = 1;
    65: op1_11_inv07 = 1;
    66: op1_11_inv07 = 1;
    68: op1_11_inv07 = 1;
    69: op1_11_inv07 = 1;
    72: op1_11_inv07 = 1;
    82: op1_11_inv07 = 1;
    83: op1_11_inv07 = 1;
    84: op1_11_inv07 = 1;
    86: op1_11_inv07 = 1;
    88: op1_11_inv07 = 1;
    89: op1_11_inv07 = 1;
    93: op1_11_inv07 = 1;
    94: op1_11_inv07 = 1;
    95: op1_11_inv07 = 1;
    96: op1_11_inv07 = 1;
    default: op1_11_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in08 = reg_0084;
    6: op1_11_in08 = reg_0121;
    7: op1_11_in08 = reg_0048;
    8: op1_11_in08 = reg_0423;
    9: op1_11_in08 = reg_0318;
    10: op1_11_in08 = reg_0473;
    11: op1_11_in08 = reg_0540;
    12: op1_11_in08 = reg_0689;
    13: op1_11_in08 = reg_0944;
    14: op1_11_in08 = reg_0716;
    15: op1_11_in08 = reg_0692;
    32: op1_11_in08 = reg_0692;
    16: op1_11_in08 = reg_0322;
    17: op1_11_in08 = reg_0142;
    18: op1_11_in08 = reg_0993;
    19: op1_11_in08 = reg_0250;
    20: op1_11_in08 = reg_0374;
    21: op1_11_in08 = reg_0805;
    22: op1_11_in08 = reg_1038;
    23: op1_11_in08 = reg_0291;
    24: op1_11_in08 = reg_0114;
    25: op1_11_in08 = reg_0991;
    26: op1_11_in08 = reg_0203;
    27: op1_11_in08 = reg_0968;
    28: op1_11_in08 = reg_0966;
    29: op1_11_in08 = reg_0334;
    30: op1_11_in08 = imem03_in[127:124];
    31: op1_11_in08 = imem06_in[91:88];
    33: op1_11_in08 = reg_0694;
    34: op1_11_in08 = reg_0981;
    35: op1_11_in08 = reg_0160;
    36: op1_11_in08 = reg_0168;
    37: op1_11_in08 = reg_0189;
    39: op1_11_in08 = reg_0082;
    40: op1_11_in08 = reg_0795;
    41: op1_11_in08 = reg_0989;
    43: op1_11_in08 = reg_0690;
    44: op1_11_in08 = reg_0665;
    45: op1_11_in08 = reg_0407;
    83: op1_11_in08 = reg_0407;
    46: op1_11_in08 = reg_0180;
    47: op1_11_in08 = reg_0418;
    48: op1_11_in08 = reg_0131;
    49: op1_11_in08 = reg_0712;
    50: op1_11_in08 = reg_0529;
    51: op1_11_in08 = reg_0994;
    52: op1_11_in08 = reg_0661;
    53: op1_11_in08 = imem04_in[55:52];
    54: op1_11_in08 = reg_0820;
    55: op1_11_in08 = reg_0243;
    57: op1_11_in08 = reg_0596;
    58: op1_11_in08 = imem07_in[19:16];
    61: op1_11_in08 = reg_0477;
    62: op1_11_in08 = reg_0646;
    63: op1_11_in08 = reg_0972;
    64: op1_11_in08 = reg_0493;
    65: op1_11_in08 = reg_0804;
    66: op1_11_in08 = reg_0325;
    67: op1_11_in08 = reg_0613;
    68: op1_11_in08 = imem02_in[47:44];
    69: op1_11_in08 = reg_0590;
    71: op1_11_in08 = reg_0478;
    72: op1_11_in08 = reg_0967;
    74: op1_11_in08 = reg_0181;
    75: op1_11_in08 = reg_0828;
    76: op1_11_in08 = reg_0096;
    77: op1_11_in08 = imem04_in[31:28];
    78: op1_11_in08 = reg_0581;
    79: op1_11_in08 = reg_0780;
    81: op1_11_in08 = reg_0674;
    82: op1_11_in08 = reg_0721;
    84: op1_11_in08 = reg_0745;
    85: op1_11_in08 = imem07_in[71:68];
    86: op1_11_in08 = reg_0825;
    87: op1_11_in08 = reg_0870;
    88: op1_11_in08 = imem07_in[7:4];
    89: op1_11_in08 = imem04_in[59:56];
    90: op1_11_in08 = reg_1028;
    91: op1_11_in08 = reg_0338;
    92: op1_11_in08 = reg_0451;
    93: op1_11_in08 = imem02_in[91:88];
    94: op1_11_in08 = imem02_in[103:100];
    95: op1_11_in08 = reg_0394;
    96: op1_11_in08 = reg_0323;
    default: op1_11_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv08 = 1;
    7: op1_11_inv08 = 1;
    9: op1_11_inv08 = 1;
    11: op1_11_inv08 = 1;
    13: op1_11_inv08 = 1;
    16: op1_11_inv08 = 1;
    17: op1_11_inv08 = 1;
    18: op1_11_inv08 = 1;
    19: op1_11_inv08 = 1;
    20: op1_11_inv08 = 1;
    23: op1_11_inv08 = 1;
    25: op1_11_inv08 = 1;
    26: op1_11_inv08 = 1;
    29: op1_11_inv08 = 1;
    34: op1_11_inv08 = 1;
    35: op1_11_inv08 = 1;
    36: op1_11_inv08 = 1;
    40: op1_11_inv08 = 1;
    43: op1_11_inv08 = 1;
    45: op1_11_inv08 = 1;
    47: op1_11_inv08 = 1;
    49: op1_11_inv08 = 1;
    50: op1_11_inv08 = 1;
    53: op1_11_inv08 = 1;
    54: op1_11_inv08 = 1;
    61: op1_11_inv08 = 1;
    67: op1_11_inv08 = 1;
    68: op1_11_inv08 = 1;
    69: op1_11_inv08 = 1;
    72: op1_11_inv08 = 1;
    74: op1_11_inv08 = 1;
    77: op1_11_inv08 = 1;
    82: op1_11_inv08 = 1;
    85: op1_11_inv08 = 1;
    86: op1_11_inv08 = 1;
    88: op1_11_inv08 = 1;
    89: op1_11_inv08 = 1;
    90: op1_11_inv08 = 1;
    96: op1_11_inv08 = 1;
    default: op1_11_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in09 = reg_0094;
    6: op1_11_in09 = reg_0110;
    84: op1_11_in09 = reg_0110;
    7: op1_11_in09 = reg_0074;
    8: op1_11_in09 = reg_0175;
    9: op1_11_in09 = reg_0330;
    10: op1_11_in09 = reg_0467;
    11: op1_11_in09 = reg_0301;
    12: op1_11_in09 = reg_0686;
    13: op1_11_in09 = reg_0955;
    14: op1_11_in09 = reg_0731;
    15: op1_11_in09 = reg_0463;
    32: op1_11_in09 = reg_0463;
    16: op1_11_in09 = reg_0323;
    17: op1_11_in09 = reg_0154;
    18: op1_11_in09 = reg_0986;
    19: op1_11_in09 = reg_0908;
    20: op1_11_in09 = reg_0991;
    21: op1_11_in09 = imem07_in[11:8];
    22: op1_11_in09 = reg_1034;
    23: op1_11_in09 = imem03_in[7:4];
    24: op1_11_in09 = reg_0101;
    25: op1_11_in09 = reg_0980;
    26: op1_11_in09 = reg_0193;
    27: op1_11_in09 = reg_0946;
    28: op1_11_in09 = reg_0954;
    29: op1_11_in09 = reg_0045;
    30: op1_11_in09 = reg_0589;
    31: op1_11_in09 = imem06_in[107:104];
    33: op1_11_in09 = reg_0676;
    34: op1_11_in09 = reg_0988;
    35: op1_11_in09 = reg_0183;
    37: op1_11_in09 = imem01_in[3:0];
    39: op1_11_in09 = reg_0007;
    40: op1_11_in09 = reg_0311;
    41: op1_11_in09 = imem04_in[27:24];
    43: op1_11_in09 = reg_0465;
    44: op1_11_in09 = reg_0667;
    45: op1_11_in09 = reg_0611;
    46: op1_11_in09 = reg_0161;
    74: op1_11_in09 = reg_0161;
    47: op1_11_in09 = reg_0081;
    48: op1_11_in09 = imem06_in[7:4];
    49: op1_11_in09 = reg_0708;
    50: op1_11_in09 = reg_0777;
    51: op1_11_in09 = imem04_in[39:36];
    78: op1_11_in09 = imem04_in[39:36];
    52: op1_11_in09 = reg_0035;
    53: op1_11_in09 = imem04_in[127:124];
    54: op1_11_in09 = reg_0844;
    69: op1_11_in09 = reg_0844;
    55: op1_11_in09 = reg_0804;
    57: op1_11_in09 = reg_0005;
    58: op1_11_in09 = imem07_in[39:36];
    61: op1_11_in09 = reg_0469;
    62: op1_11_in09 = reg_0639;
    63: op1_11_in09 = reg_0337;
    64: op1_11_in09 = reg_0448;
    65: op1_11_in09 = reg_0695;
    66: op1_11_in09 = reg_0047;
    67: op1_11_in09 = reg_0617;
    68: op1_11_in09 = imem02_in[79:76];
    71: op1_11_in09 = reg_0208;
    72: op1_11_in09 = reg_0949;
    75: op1_11_in09 = reg_0462;
    76: op1_11_in09 = reg_0649;
    77: op1_11_in09 = imem04_in[51:48];
    79: op1_11_in09 = reg_0970;
    81: op1_11_in09 = reg_0680;
    82: op1_11_in09 = reg_0560;
    83: op1_11_in09 = reg_0444;
    85: op1_11_in09 = imem07_in[91:88];
    86: op1_11_in09 = reg_0883;
    87: op1_11_in09 = reg_0156;
    88: op1_11_in09 = imem07_in[15:12];
    89: op1_11_in09 = imem04_in[63:60];
    90: op1_11_in09 = reg_0380;
    91: op1_11_in09 = reg_1011;
    92: op1_11_in09 = reg_0464;
    93: op1_11_in09 = imem02_in[99:96];
    94: op1_11_in09 = imem02_in[115:112];
    95: op1_11_in09 = reg_0389;
    96: op1_11_in09 = reg_0739;
    default: op1_11_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv09 = 1;
    11: op1_11_inv09 = 1;
    12: op1_11_inv09 = 1;
    13: op1_11_inv09 = 1;
    14: op1_11_inv09 = 1;
    15: op1_11_inv09 = 1;
    16: op1_11_inv09 = 1;
    19: op1_11_inv09 = 1;
    20: op1_11_inv09 = 1;
    21: op1_11_inv09 = 1;
    24: op1_11_inv09 = 1;
    28: op1_11_inv09 = 1;
    30: op1_11_inv09 = 1;
    37: op1_11_inv09 = 1;
    39: op1_11_inv09 = 1;
    40: op1_11_inv09 = 1;
    43: op1_11_inv09 = 1;
    44: op1_11_inv09 = 1;
    46: op1_11_inv09 = 1;
    49: op1_11_inv09 = 1;
    52: op1_11_inv09 = 1;
    53: op1_11_inv09 = 1;
    55: op1_11_inv09 = 1;
    57: op1_11_inv09 = 1;
    58: op1_11_inv09 = 1;
    61: op1_11_inv09 = 1;
    63: op1_11_inv09 = 1;
    64: op1_11_inv09 = 1;
    66: op1_11_inv09 = 1;
    67: op1_11_inv09 = 1;
    75: op1_11_inv09 = 1;
    76: op1_11_inv09 = 1;
    77: op1_11_inv09 = 1;
    81: op1_11_inv09 = 1;
    82: op1_11_inv09 = 1;
    84: op1_11_inv09 = 1;
    85: op1_11_inv09 = 1;
    86: op1_11_inv09 = 1;
    87: op1_11_inv09 = 1;
    88: op1_11_inv09 = 1;
    90: op1_11_inv09 = 1;
    93: op1_11_inv09 = 1;
    94: op1_11_inv09 = 1;
    default: op1_11_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in10 = imem03_in[27:24];
    6: op1_11_in10 = imem02_in[39:36];
    7: op1_11_in10 = imem05_in[67:64];
    8: op1_11_in10 = reg_0180;
    9: op1_11_in10 = reg_0314;
    10: op1_11_in10 = reg_0470;
    75: op1_11_in10 = reg_0470;
    11: op1_11_in10 = reg_0300;
    62: op1_11_in10 = reg_0300;
    12: op1_11_in10 = reg_0679;
    13: op1_11_in10 = reg_0957;
    28: op1_11_in10 = reg_0957;
    14: op1_11_in10 = reg_0702;
    15: op1_11_in10 = reg_0450;
    16: op1_11_in10 = reg_0992;
    20: op1_11_in10 = reg_0992;
    17: op1_11_in10 = reg_0143;
    18: op1_11_in10 = reg_0978;
    25: op1_11_in10 = reg_0978;
    19: op1_11_in10 = reg_0836;
    21: op1_11_in10 = imem07_in[19:16];
    22: op1_11_in10 = reg_0111;
    23: op1_11_in10 = imem03_in[15:12];
    24: op1_11_in10 = reg_0121;
    26: op1_11_in10 = reg_0201;
    27: op1_11_in10 = reg_0961;
    29: op1_11_in10 = reg_0290;
    30: op1_11_in10 = reg_0600;
    31: op1_11_in10 = reg_0605;
    32: op1_11_in10 = reg_0465;
    33: op1_11_in10 = reg_0670;
    34: op1_11_in10 = imem04_in[59:56];
    35: op1_11_in10 = reg_0177;
    74: op1_11_in10 = reg_0177;
    37: op1_11_in10 = imem01_in[11:8];
    39: op1_11_in10 = reg_0761;
    40: op1_11_in10 = reg_0979;
    41: op1_11_in10 = imem04_in[39:36];
    43: op1_11_in10 = reg_0457;
    44: op1_11_in10 = reg_0663;
    45: op1_11_in10 = reg_0595;
    46: op1_11_in10 = reg_0167;
    47: op1_11_in10 = reg_0039;
    48: op1_11_in10 = imem06_in[11:8];
    49: op1_11_in10 = reg_0705;
    50: op1_11_in10 = reg_0750;
    51: op1_11_in10 = imem04_in[63:60];
    52: op1_11_in10 = reg_0360;
    53: op1_11_in10 = reg_1003;
    54: op1_11_in10 = reg_0986;
    55: op1_11_in10 = reg_1029;
    57: op1_11_in10 = imem07_in[7:4];
    58: op1_11_in10 = imem07_in[47:44];
    61: op1_11_in10 = reg_0456;
    63: op1_11_in10 = reg_0404;
    64: op1_11_in10 = reg_0333;
    65: op1_11_in10 = reg_0946;
    66: op1_11_in10 = reg_0427;
    67: op1_11_in10 = reg_0533;
    68: op1_11_in10 = imem02_in[87:84];
    69: op1_11_in10 = reg_1002;
    71: op1_11_in10 = reg_0187;
    72: op1_11_in10 = reg_0326;
    76: op1_11_in10 = reg_0260;
    77: op1_11_in10 = imem04_in[55:52];
    78: op1_11_in10 = imem04_in[43:40];
    79: op1_11_in10 = reg_0135;
    81: op1_11_in10 = reg_0453;
    82: op1_11_in10 = reg_0708;
    83: op1_11_in10 = reg_0041;
    84: op1_11_in10 = reg_0079;
    85: op1_11_in10 = imem07_in[111:108];
    86: op1_11_in10 = reg_0674;
    87: op1_11_in10 = reg_0540;
    88: op1_11_in10 = imem07_in[23:20];
    89: op1_11_in10 = imem04_in[71:68];
    90: op1_11_in10 = reg_0918;
    91: op1_11_in10 = reg_0735;
    92: op1_11_in10 = reg_0191;
    93: op1_11_in10 = imem02_in[119:116];
    94: op1_11_in10 = reg_0536;
    95: op1_11_in10 = reg_0248;
    96: op1_11_in10 = reg_0664;
    default: op1_11_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv10 = 1;
    9: op1_11_inv10 = 1;
    14: op1_11_inv10 = 1;
    16: op1_11_inv10 = 1;
    18: op1_11_inv10 = 1;
    19: op1_11_inv10 = 1;
    20: op1_11_inv10 = 1;
    26: op1_11_inv10 = 1;
    28: op1_11_inv10 = 1;
    29: op1_11_inv10 = 1;
    30: op1_11_inv10 = 1;
    33: op1_11_inv10 = 1;
    34: op1_11_inv10 = 1;
    37: op1_11_inv10 = 1;
    40: op1_11_inv10 = 1;
    43: op1_11_inv10 = 1;
    44: op1_11_inv10 = 1;
    45: op1_11_inv10 = 1;
    46: op1_11_inv10 = 1;
    48: op1_11_inv10 = 1;
    50: op1_11_inv10 = 1;
    51: op1_11_inv10 = 1;
    52: op1_11_inv10 = 1;
    57: op1_11_inv10 = 1;
    58: op1_11_inv10 = 1;
    63: op1_11_inv10 = 1;
    64: op1_11_inv10 = 1;
    68: op1_11_inv10 = 1;
    71: op1_11_inv10 = 1;
    72: op1_11_inv10 = 1;
    74: op1_11_inv10 = 1;
    75: op1_11_inv10 = 1;
    83: op1_11_inv10 = 1;
    86: op1_11_inv10 = 1;
    87: op1_11_inv10 = 1;
    88: op1_11_inv10 = 1;
    93: op1_11_inv10 = 1;
    96: op1_11_inv10 = 1;
    default: op1_11_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in11 = imem03_in[47:44];
    6: op1_11_in11 = imem02_in[71:68];
    7: op1_11_in11 = imem05_in[79:76];
    8: op1_11_in11 = reg_0161;
    9: op1_11_in11 = reg_0347;
    10: op1_11_in11 = reg_0479;
    11: op1_11_in11 = reg_0302;
    12: op1_11_in11 = reg_0453;
    13: op1_11_in11 = reg_0964;
    14: op1_11_in11 = reg_0729;
    15: op1_11_in11 = reg_0451;
    16: op1_11_in11 = reg_0977;
    18: op1_11_in11 = reg_0977;
    17: op1_11_in11 = reg_0144;
    19: op1_11_in11 = reg_0902;
    20: op1_11_in11 = reg_0974;
    21: op1_11_in11 = imem07_in[35:32];
    22: op1_11_in11 = reg_0119;
    23: op1_11_in11 = imem03_in[19:16];
    24: op1_11_in11 = reg_0110;
    25: op1_11_in11 = reg_0988;
    26: op1_11_in11 = reg_0190;
    27: op1_11_in11 = reg_0943;
    28: op1_11_in11 = reg_0969;
    29: op1_11_in11 = reg_0225;
    30: op1_11_in11 = reg_0597;
    31: op1_11_in11 = reg_0626;
    32: op1_11_in11 = reg_0457;
    33: op1_11_in11 = reg_0687;
    34: op1_11_in11 = imem04_in[79:76];
    37: op1_11_in11 = imem01_in[79:76];
    39: op1_11_in11 = reg_0814;
    40: op1_11_in11 = reg_0980;
    69: op1_11_in11 = reg_0980;
    41: op1_11_in11 = imem04_in[51:48];
    43: op1_11_in11 = reg_0481;
    44: op1_11_in11 = reg_0080;
    45: op1_11_in11 = reg_0612;
    47: op1_11_in11 = reg_0097;
    48: op1_11_in11 = imem06_in[23:20];
    49: op1_11_in11 = reg_0718;
    50: op1_11_in11 = reg_0973;
    51: op1_11_in11 = imem04_in[87:84];
    52: op1_11_in11 = reg_0082;
    53: op1_11_in11 = reg_0937;
    54: op1_11_in11 = reg_0978;
    55: op1_11_in11 = reg_0625;
    57: op1_11_in11 = imem07_in[31:28];
    58: op1_11_in11 = imem07_in[63:60];
    61: op1_11_in11 = reg_0191;
    62: op1_11_in11 = reg_0279;
    76: op1_11_in11 = reg_0279;
    63: op1_11_in11 = reg_1046;
    64: op1_11_in11 = reg_0145;
    65: op1_11_in11 = reg_0816;
    66: op1_11_in11 = reg_0431;
    67: op1_11_in11 = reg_0439;
    68: op1_11_in11 = imem02_in[91:88];
    71: op1_11_in11 = reg_0203;
    72: op1_11_in11 = reg_0343;
    74: op1_11_in11 = reg_0178;
    75: op1_11_in11 = reg_0468;
    77: op1_11_in11 = reg_0483;
    78: op1_11_in11 = imem04_in[47:44];
    79: op1_11_in11 = reg_0486;
    81: op1_11_in11 = reg_0454;
    82: op1_11_in11 = reg_0442;
    83: op1_11_in11 = reg_0065;
    84: op1_11_in11 = imem02_in[19:16];
    85: op1_11_in11 = reg_0712;
    86: op1_11_in11 = reg_0102;
    87: op1_11_in11 = reg_0586;
    88: op1_11_in11 = imem07_in[27:24];
    89: op1_11_in11 = imem04_in[75:72];
    90: op1_11_in11 = reg_0293;
    91: op1_11_in11 = reg_0787;
    92: op1_11_in11 = reg_0194;
    93: op1_11_in11 = reg_0334;
    94: op1_11_in11 = reg_0255;
    95: op1_11_in11 = reg_0516;
    96: op1_11_in11 = reg_0329;
    default: op1_11_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv11 = 1;
    6: op1_11_inv11 = 1;
    7: op1_11_inv11 = 1;
    8: op1_11_inv11 = 1;
    10: op1_11_inv11 = 1;
    16: op1_11_inv11 = 1;
    18: op1_11_inv11 = 1;
    20: op1_11_inv11 = 1;
    22: op1_11_inv11 = 1;
    24: op1_11_inv11 = 1;
    25: op1_11_inv11 = 1;
    26: op1_11_inv11 = 1;
    28: op1_11_inv11 = 1;
    29: op1_11_inv11 = 1;
    31: op1_11_inv11 = 1;
    34: op1_11_inv11 = 1;
    37: op1_11_inv11 = 1;
    43: op1_11_inv11 = 1;
    45: op1_11_inv11 = 1;
    47: op1_11_inv11 = 1;
    48: op1_11_inv11 = 1;
    49: op1_11_inv11 = 1;
    50: op1_11_inv11 = 1;
    53: op1_11_inv11 = 1;
    63: op1_11_inv11 = 1;
    64: op1_11_inv11 = 1;
    65: op1_11_inv11 = 1;
    66: op1_11_inv11 = 1;
    71: op1_11_inv11 = 1;
    74: op1_11_inv11 = 1;
    76: op1_11_inv11 = 1;
    78: op1_11_inv11 = 1;
    81: op1_11_inv11 = 1;
    82: op1_11_inv11 = 1;
    83: op1_11_inv11 = 1;
    86: op1_11_inv11 = 1;
    88: op1_11_inv11 = 1;
    92: op1_11_inv11 = 1;
    95: op1_11_inv11 = 1;
    default: op1_11_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in12 = imem03_in[111:108];
    6: op1_11_in12 = imem02_in[111:108];
    68: op1_11_in12 = imem02_in[111:108];
    7: op1_11_in12 = imem05_in[87:84];
    8: op1_11_in12 = reg_0167;
    9: op1_11_in12 = reg_0092;
    10: op1_11_in12 = reg_0459;
    11: op1_11_in12 = reg_0293;
    12: op1_11_in12 = reg_0469;
    13: op1_11_in12 = reg_0968;
    14: op1_11_in12 = reg_0707;
    15: op1_11_in12 = reg_0455;
    16: op1_11_in12 = reg_0976;
    17: op1_11_in12 = imem06_in[19:16];
    18: op1_11_in12 = reg_0997;
    25: op1_11_in12 = reg_0997;
    19: op1_11_in12 = reg_0255;
    20: op1_11_in12 = imem04_in[15:12];
    21: op1_11_in12 = imem07_in[51:48];
    22: op1_11_in12 = reg_0102;
    23: op1_11_in12 = imem03_in[71:68];
    24: op1_11_in12 = imem02_in[11:8];
    26: op1_11_in12 = reg_0195;
    27: op1_11_in12 = reg_0215;
    28: op1_11_in12 = reg_0964;
    29: op1_11_in12 = reg_0886;
    30: op1_11_in12 = reg_0590;
    31: op1_11_in12 = reg_0632;
    32: op1_11_in12 = reg_0461;
    33: op1_11_in12 = reg_0463;
    34: op1_11_in12 = imem04_in[115:112];
    37: op1_11_in12 = imem01_in[127:124];
    39: op1_11_in12 = reg_0086;
    40: op1_11_in12 = reg_0994;
    41: op1_11_in12 = imem04_in[79:76];
    43: op1_11_in12 = reg_0201;
    44: op1_11_in12 = reg_0098;
    45: op1_11_in12 = reg_0387;
    47: op1_11_in12 = reg_0225;
    48: op1_11_in12 = imem06_in[55:52];
    49: op1_11_in12 = reg_0701;
    50: op1_11_in12 = reg_0959;
    51: op1_11_in12 = reg_0507;
    52: op1_11_in12 = reg_0300;
    53: op1_11_in12 = reg_1005;
    54: op1_11_in12 = reg_0977;
    55: op1_11_in12 = reg_1010;
    57: op1_11_in12 = imem07_in[67:64];
    58: op1_11_in12 = imem07_in[103:100];
    61: op1_11_in12 = reg_0210;
    62: op1_11_in12 = reg_0358;
    76: op1_11_in12 = reg_0358;
    63: op1_11_in12 = reg_0819;
    64: op1_11_in12 = reg_0136;
    65: op1_11_in12 = reg_0605;
    66: op1_11_in12 = reg_0174;
    67: op1_11_in12 = reg_0595;
    69: op1_11_in12 = reg_0988;
    71: op1_11_in12 = reg_0194;
    72: op1_11_in12 = reg_0963;
    74: op1_11_in12 = reg_0158;
    75: op1_11_in12 = reg_0478;
    77: op1_11_in12 = reg_0301;
    78: op1_11_in12 = reg_0937;
    79: op1_11_in12 = reg_0806;
    81: op1_11_in12 = reg_0450;
    82: op1_11_in12 = reg_0563;
    83: op1_11_in12 = reg_0517;
    84: op1_11_in12 = imem02_in[43:40];
    85: op1_11_in12 = reg_0374;
    86: op1_11_in12 = reg_0663;
    87: op1_11_in12 = reg_0066;
    88: op1_11_in12 = imem07_in[87:84];
    89: op1_11_in12 = imem04_in[87:84];
    90: op1_11_in12 = reg_0807;
    91: op1_11_in12 = reg_0895;
    92: op1_11_in12 = reg_0212;
    93: op1_11_in12 = reg_0844;
    94: op1_11_in12 = reg_0055;
    95: op1_11_in12 = reg_0083;
    96: op1_11_in12 = reg_0423;
    default: op1_11_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_11_inv12 = 1;
    8: op1_11_inv12 = 1;
    9: op1_11_inv12 = 1;
    10: op1_11_inv12 = 1;
    11: op1_11_inv12 = 1;
    17: op1_11_inv12 = 1;
    18: op1_11_inv12 = 1;
    25: op1_11_inv12 = 1;
    27: op1_11_inv12 = 1;
    28: op1_11_inv12 = 1;
    29: op1_11_inv12 = 1;
    31: op1_11_inv12 = 1;
    32: op1_11_inv12 = 1;
    39: op1_11_inv12 = 1;
    43: op1_11_inv12 = 1;
    47: op1_11_inv12 = 1;
    48: op1_11_inv12 = 1;
    50: op1_11_inv12 = 1;
    51: op1_11_inv12 = 1;
    52: op1_11_inv12 = 1;
    53: op1_11_inv12 = 1;
    63: op1_11_inv12 = 1;
    64: op1_11_inv12 = 1;
    65: op1_11_inv12 = 1;
    66: op1_11_inv12 = 1;
    67: op1_11_inv12 = 1;
    69: op1_11_inv12 = 1;
    71: op1_11_inv12 = 1;
    74: op1_11_inv12 = 1;
    75: op1_11_inv12 = 1;
    76: op1_11_inv12 = 1;
    77: op1_11_inv12 = 1;
    79: op1_11_inv12 = 1;
    82: op1_11_inv12 = 1;
    83: op1_11_inv12 = 1;
    84: op1_11_inv12 = 1;
    93: op1_11_inv12 = 1;
    95: op1_11_inv12 = 1;
    default: op1_11_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in13 = reg_0586;
    6: op1_11_in13 = reg_0655;
    7: op1_11_in13 = imem05_in[107:104];
    8: op1_11_in13 = reg_0163;
    9: op1_11_in13 = reg_0090;
    10: op1_11_in13 = reg_0210;
    11: op1_11_in13 = reg_0296;
    12: op1_11_in13 = reg_0473;
    13: op1_11_in13 = reg_0953;
    14: op1_11_in13 = reg_0430;
    15: op1_11_in13 = reg_0457;
    16: op1_11_in13 = imem04_in[15:12];
    17: op1_11_in13 = imem06_in[63:60];
    18: op1_11_in13 = reg_0265;
    19: op1_11_in13 = reg_0253;
    20: op1_11_in13 = imem04_in[19:16];
    21: op1_11_in13 = imem07_in[107:104];
    22: op1_11_in13 = reg_0126;
    23: op1_11_in13 = imem03_in[119:116];
    24: op1_11_in13 = imem02_in[27:24];
    25: op1_11_in13 = imem04_in[39:36];
    26: op1_11_in13 = reg_0199;
    27: op1_11_in13 = reg_0757;
    28: op1_11_in13 = reg_0968;
    29: op1_11_in13 = reg_0865;
    72: op1_11_in13 = reg_0865;
    30: op1_11_in13 = reg_0765;
    31: op1_11_in13 = reg_0627;
    32: op1_11_in13 = reg_0472;
    33: op1_11_in13 = reg_0477;
    86: op1_11_in13 = reg_0477;
    34: op1_11_in13 = imem04_in[119:116];
    37: op1_11_in13 = reg_0299;
    39: op1_11_in13 = reg_0310;
    40: op1_11_in13 = imem04_in[27:24];
    41: op1_11_in13 = imem04_in[83:80];
    43: op1_11_in13 = imem01_in[83:80];
    44: op1_11_in13 = reg_0817;
    45: op1_11_in13 = reg_0351;
    47: op1_11_in13 = reg_0818;
    48: op1_11_in13 = reg_0614;
    49: op1_11_in13 = reg_0706;
    50: op1_11_in13 = reg_0956;
    51: op1_11_in13 = reg_0067;
    52: op1_11_in13 = imem02_in[7:4];
    53: op1_11_in13 = reg_0888;
    54: op1_11_in13 = reg_0997;
    55: op1_11_in13 = reg_0531;
    57: op1_11_in13 = imem07_in[75:72];
    58: op1_11_in13 = reg_0730;
    61: op1_11_in13 = reg_0187;
    62: op1_11_in13 = reg_0739;
    63: op1_11_in13 = reg_0148;
    64: op1_11_in13 = reg_0133;
    65: op1_11_in13 = reg_0264;
    66: op1_11_in13 = reg_0175;
    67: op1_11_in13 = reg_0241;
    68: op1_11_in13 = reg_0653;
    69: op1_11_in13 = reg_1000;
    71: op1_11_in13 = reg_0202;
    75: op1_11_in13 = reg_0200;
    76: op1_11_in13 = reg_0329;
    77: op1_11_in13 = reg_0282;
    78: op1_11_in13 = reg_1009;
    79: op1_11_in13 = reg_0945;
    81: op1_11_in13 = reg_0455;
    82: op1_11_in13 = reg_0759;
    83: op1_11_in13 = reg_0854;
    84: op1_11_in13 = imem02_in[51:48];
    85: op1_11_in13 = reg_0923;
    87: op1_11_in13 = reg_0015;
    88: op1_11_in13 = reg_0728;
    89: op1_11_in13 = imem04_in[95:92];
    90: op1_11_in13 = reg_0392;
    91: op1_11_in13 = reg_0792;
    92: op1_11_in13 = reg_0205;
    93: op1_11_in13 = reg_0285;
    94: op1_11_in13 = reg_0323;
    95: op1_11_in13 = reg_0045;
    96: op1_11_in13 = reg_0037;
    default: op1_11_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv13 = 1;
    7: op1_11_inv13 = 1;
    9: op1_11_inv13 = 1;
    10: op1_11_inv13 = 1;
    14: op1_11_inv13 = 1;
    15: op1_11_inv13 = 1;
    18: op1_11_inv13 = 1;
    21: op1_11_inv13 = 1;
    22: op1_11_inv13 = 1;
    23: op1_11_inv13 = 1;
    24: op1_11_inv13 = 1;
    25: op1_11_inv13 = 1;
    27: op1_11_inv13 = 1;
    29: op1_11_inv13 = 1;
    32: op1_11_inv13 = 1;
    34: op1_11_inv13 = 1;
    40: op1_11_inv13 = 1;
    41: op1_11_inv13 = 1;
    43: op1_11_inv13 = 1;
    49: op1_11_inv13 = 1;
    51: op1_11_inv13 = 1;
    52: op1_11_inv13 = 1;
    53: op1_11_inv13 = 1;
    54: op1_11_inv13 = 1;
    57: op1_11_inv13 = 1;
    58: op1_11_inv13 = 1;
    62: op1_11_inv13 = 1;
    68: op1_11_inv13 = 1;
    69: op1_11_inv13 = 1;
    71: op1_11_inv13 = 1;
    77: op1_11_inv13 = 1;
    78: op1_11_inv13 = 1;
    81: op1_11_inv13 = 1;
    82: op1_11_inv13 = 1;
    83: op1_11_inv13 = 1;
    84: op1_11_inv13 = 1;
    85: op1_11_inv13 = 1;
    86: op1_11_inv13 = 1;
    92: op1_11_inv13 = 1;
    93: op1_11_inv13 = 1;
    94: op1_11_inv13 = 1;
    default: op1_11_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in14 = reg_0587;
    6: op1_11_in14 = reg_0654;
    7: op1_11_in14 = imem05_in[111:108];
    9: op1_11_in14 = imem03_in[39:36];
    10: op1_11_in14 = reg_0189;
    11: op1_11_in14 = reg_0278;
    12: op1_11_in14 = reg_0459;
    13: op1_11_in14 = reg_0835;
    14: op1_11_in14 = reg_0429;
    15: op1_11_in14 = reg_0480;
    33: op1_11_in14 = reg_0480;
    16: op1_11_in14 = imem04_in[23:20];
    69: op1_11_in14 = imem04_in[23:20];
    17: op1_11_in14 = reg_0613;
    18: op1_11_in14 = reg_0260;
    19: op1_11_in14 = reg_0135;
    20: op1_11_in14 = imem04_in[43:40];
    21: op1_11_in14 = reg_0730;
    22: op1_11_in14 = reg_0110;
    23: op1_11_in14 = reg_0598;
    24: op1_11_in14 = imem02_in[123:120];
    25: op1_11_in14 = imem04_in[83:80];
    26: op1_11_in14 = reg_0197;
    27: op1_11_in14 = reg_0251;
    83: op1_11_in14 = reg_0251;
    28: op1_11_in14 = reg_0945;
    29: op1_11_in14 = reg_0516;
    30: op1_11_in14 = reg_0543;
    31: op1_11_in14 = reg_0344;
    32: op1_11_in14 = reg_0473;
    34: op1_11_in14 = imem04_in[127:124];
    37: op1_11_in14 = reg_0811;
    39: op1_11_in14 = reg_0484;
    40: op1_11_in14 = imem04_in[31:28];
    41: op1_11_in14 = reg_1004;
    43: op1_11_in14 = imem01_in[95:92];
    44: op1_11_in14 = reg_0338;
    47: op1_11_in14 = reg_0338;
    45: op1_11_in14 = reg_0393;
    48: op1_11_in14 = reg_0407;
    49: op1_11_in14 = reg_0575;
    50: op1_11_in14 = reg_0957;
    51: op1_11_in14 = reg_0056;
    52: op1_11_in14 = imem02_in[11:8];
    53: op1_11_in14 = reg_1016;
    54: op1_11_in14 = imem04_in[3:0];
    55: op1_11_in14 = reg_0005;
    57: op1_11_in14 = imem07_in[83:80];
    58: op1_11_in14 = reg_0721;
    61: op1_11_in14 = reg_0209;
    62: op1_11_in14 = reg_0424;
    63: op1_11_in14 = reg_0151;
    64: op1_11_in14 = reg_0151;
    65: op1_11_in14 = reg_0633;
    66: op1_11_in14 = reg_0159;
    67: op1_11_in14 = reg_1028;
    68: op1_11_in14 = reg_0845;
    71: op1_11_in14 = imem01_in[19:16];
    72: op1_11_in14 = reg_0153;
    75: op1_11_in14 = reg_0210;
    76: op1_11_in14 = reg_0425;
    77: op1_11_in14 = reg_0306;
    78: op1_11_in14 = reg_0401;
    79: op1_11_in14 = reg_0741;
    81: op1_11_in14 = reg_0475;
    82: op1_11_in14 = reg_0727;
    84: op1_11_in14 = imem02_in[55:52];
    85: op1_11_in14 = reg_0759;
    86: op1_11_in14 = reg_0469;
    87: op1_11_in14 = reg_0893;
    88: op1_11_in14 = reg_0165;
    89: op1_11_in14 = reg_0126;
    90: op1_11_in14 = reg_0040;
    91: op1_11_in14 = reg_0533;
    92: op1_11_in14 = reg_0199;
    93: op1_11_in14 = reg_0075;
    94: op1_11_in14 = reg_0441;
    95: op1_11_in14 = reg_0778;
    96: op1_11_in14 = reg_0335;
    default: op1_11_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv14 = 1;
    7: op1_11_inv14 = 1;
    9: op1_11_inv14 = 1;
    10: op1_11_inv14 = 1;
    12: op1_11_inv14 = 1;
    13: op1_11_inv14 = 1;
    14: op1_11_inv14 = 1;
    15: op1_11_inv14 = 1;
    17: op1_11_inv14 = 1;
    18: op1_11_inv14 = 1;
    20: op1_11_inv14 = 1;
    22: op1_11_inv14 = 1;
    24: op1_11_inv14 = 1;
    25: op1_11_inv14 = 1;
    27: op1_11_inv14 = 1;
    31: op1_11_inv14 = 1;
    34: op1_11_inv14 = 1;
    39: op1_11_inv14 = 1;
    41: op1_11_inv14 = 1;
    43: op1_11_inv14 = 1;
    48: op1_11_inv14 = 1;
    51: op1_11_inv14 = 1;
    53: op1_11_inv14 = 1;
    58: op1_11_inv14 = 1;
    61: op1_11_inv14 = 1;
    62: op1_11_inv14 = 1;
    65: op1_11_inv14 = 1;
    68: op1_11_inv14 = 1;
    69: op1_11_inv14 = 1;
    71: op1_11_inv14 = 1;
    77: op1_11_inv14 = 1;
    79: op1_11_inv14 = 1;
    81: op1_11_inv14 = 1;
    82: op1_11_inv14 = 1;
    83: op1_11_inv14 = 1;
    84: op1_11_inv14 = 1;
    88: op1_11_inv14 = 1;
    89: op1_11_inv14 = 1;
    91: op1_11_inv14 = 1;
    92: op1_11_inv14 = 1;
    93: op1_11_inv14 = 1;
    94: op1_11_inv14 = 1;
    default: op1_11_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in15 = reg_0588;
    6: op1_11_in15 = reg_0656;
    95: op1_11_in15 = reg_0656;
    7: op1_11_in15 = imem05_in[115:112];
    9: op1_11_in15 = imem03_in[43:40];
    10: op1_11_in15 = reg_0186;
    11: op1_11_in15 = reg_0046;
    12: op1_11_in15 = reg_0452;
    13: op1_11_in15 = reg_0900;
    14: op1_11_in15 = reg_0432;
    15: op1_11_in15 = reg_0473;
    16: op1_11_in15 = imem04_in[27:24];
    17: op1_11_in15 = reg_0617;
    18: op1_11_in15 = reg_0776;
    19: op1_11_in15 = reg_0156;
    20: op1_11_in15 = imem04_in[67:64];
    21: op1_11_in15 = reg_0731;
    22: op1_11_in15 = imem02_in[11:8];
    23: op1_11_in15 = reg_0582;
    24: op1_11_in15 = reg_0650;
    25: op1_11_in15 = imem04_in[91:88];
    26: op1_11_in15 = imem01_in[19:16];
    27: op1_11_in15 = reg_0260;
    28: op1_11_in15 = reg_0946;
    29: op1_11_in15 = reg_0792;
    30: op1_11_in15 = reg_0795;
    31: op1_11_in15 = reg_0914;
    32: op1_11_in15 = reg_0467;
    33: op1_11_in15 = reg_0468;
    34: op1_11_in15 = reg_0277;
    37: op1_11_in15 = reg_0249;
    39: op1_11_in15 = imem03_in[39:36];
    40: op1_11_in15 = imem04_in[51:48];
    41: op1_11_in15 = reg_0912;
    43: op1_11_in15 = imem01_in[111:108];
    44: op1_11_in15 = reg_0516;
    45: op1_11_in15 = reg_0388;
    47: op1_11_in15 = reg_0083;
    48: op1_11_in15 = reg_0020;
    49: op1_11_in15 = reg_0419;
    50: op1_11_in15 = reg_0964;
    51: op1_11_in15 = reg_0068;
    52: op1_11_in15 = imem02_in[15:12];
    53: op1_11_in15 = reg_0537;
    54: op1_11_in15 = imem04_in[7:4];
    55: op1_11_in15 = reg_0263;
    57: op1_11_in15 = reg_0720;
    58: op1_11_in15 = reg_0717;
    61: op1_11_in15 = reg_0194;
    62: op1_11_in15 = reg_0372;
    63: op1_11_in15 = reg_0128;
    64: op1_11_in15 = reg_0142;
    65: op1_11_in15 = reg_0957;
    66: op1_11_in15 = reg_0169;
    67: op1_11_in15 = reg_0605;
    68: op1_11_in15 = reg_0290;
    69: op1_11_in15 = imem04_in[75:72];
    71: op1_11_in15 = imem01_in[47:44];
    72: op1_11_in15 = reg_0144;
    75: op1_11_in15 = reg_0189;
    76: op1_11_in15 = reg_0087;
    77: op1_11_in15 = reg_0539;
    78: op1_11_in15 = reg_0764;
    87: op1_11_in15 = reg_0764;
    79: op1_11_in15 = imem06_in[7:4];
    81: op1_11_in15 = reg_0462;
    82: op1_11_in15 = reg_0805;
    83: op1_11_in15 = reg_0070;
    84: op1_11_in15 = imem02_in[67:64];
    85: op1_11_in15 = reg_0653;
    86: op1_11_in15 = reg_0476;
    88: op1_11_in15 = reg_0710;
    89: op1_11_in15 = reg_0405;
    90: op1_11_in15 = reg_0177;
    91: op1_11_in15 = reg_0928;
    92: op1_11_in15 = reg_0192;
    93: op1_11_in15 = reg_0664;
    94: op1_11_in15 = reg_0423;
    96: op1_11_in15 = reg_0347;
    default: op1_11_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_11_inv15 = 1;
    9: op1_11_inv15 = 1;
    11: op1_11_inv15 = 1;
    12: op1_11_inv15 = 1;
    15: op1_11_inv15 = 1;
    16: op1_11_inv15 = 1;
    17: op1_11_inv15 = 1;
    19: op1_11_inv15 = 1;
    24: op1_11_inv15 = 1;
    25: op1_11_inv15 = 1;
    28: op1_11_inv15 = 1;
    31: op1_11_inv15 = 1;
    33: op1_11_inv15 = 1;
    37: op1_11_inv15 = 1;
    39: op1_11_inv15 = 1;
    44: op1_11_inv15 = 1;
    45: op1_11_inv15 = 1;
    47: op1_11_inv15 = 1;
    48: op1_11_inv15 = 1;
    49: op1_11_inv15 = 1;
    50: op1_11_inv15 = 1;
    51: op1_11_inv15 = 1;
    55: op1_11_inv15 = 1;
    58: op1_11_inv15 = 1;
    62: op1_11_inv15 = 1;
    68: op1_11_inv15 = 1;
    71: op1_11_inv15 = 1;
    75: op1_11_inv15 = 1;
    78: op1_11_inv15 = 1;
    83: op1_11_inv15 = 1;
    85: op1_11_inv15 = 1;
    86: op1_11_inv15 = 1;
    87: op1_11_inv15 = 1;
    89: op1_11_inv15 = 1;
    90: op1_11_inv15 = 1;
    93: op1_11_inv15 = 1;
    94: op1_11_inv15 = 1;
    95: op1_11_inv15 = 1;
    96: op1_11_inv15 = 1;
    default: op1_11_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in16 = reg_0311;
    6: op1_11_in16 = reg_0640;
    7: op1_11_in16 = reg_0963;
    9: op1_11_in16 = imem03_in[83:80];
    10: op1_11_in16 = reg_0790;
    11: op1_11_in16 = reg_0047;
    85: op1_11_in16 = reg_0047;
    12: op1_11_in16 = reg_0189;
    13: op1_11_in16 = reg_0252;
    14: op1_11_in16 = reg_0433;
    15: op1_11_in16 = reg_0474;
    16: op1_11_in16 = imem04_in[51:48];
    17: op1_11_in16 = reg_0616;
    18: op1_11_in16 = reg_0553;
    19: op1_11_in16 = reg_0131;
    20: op1_11_in16 = imem04_in[99:96];
    21: op1_11_in16 = reg_0721;
    22: op1_11_in16 = imem02_in[31:28];
    23: op1_11_in16 = reg_0596;
    24: op1_11_in16 = reg_0645;
    25: op1_11_in16 = reg_1006;
    26: op1_11_in16 = imem01_in[47:44];
    27: op1_11_in16 = reg_0254;
    28: op1_11_in16 = reg_0952;
    29: op1_11_in16 = reg_0484;
    30: op1_11_in16 = reg_0377;
    31: op1_11_in16 = reg_0294;
    32: op1_11_in16 = reg_0479;
    33: op1_11_in16 = reg_0458;
    34: op1_11_in16 = reg_0048;
    37: op1_11_in16 = reg_1033;
    39: op1_11_in16 = imem03_in[47:44];
    40: op1_11_in16 = imem04_in[71:68];
    41: op1_11_in16 = reg_1057;
    43: op1_11_in16 = reg_0779;
    44: op1_11_in16 = reg_0876;
    45: op1_11_in16 = reg_0349;
    65: op1_11_in16 = reg_0349;
    47: op1_11_in16 = reg_0776;
    48: op1_11_in16 = reg_0627;
    49: op1_11_in16 = reg_0181;
    50: op1_11_in16 = imem05_in[67:64];
    51: op1_11_in16 = reg_0276;
    52: op1_11_in16 = imem02_in[43:40];
    53: op1_11_in16 = reg_0313;
    54: op1_11_in16 = imem04_in[15:12];
    55: op1_11_in16 = imem07_in[7:4];
    57: op1_11_in16 = reg_0700;
    58: op1_11_in16 = reg_0709;
    61: op1_11_in16 = reg_0202;
    62: op1_11_in16 = reg_0792;
    63: op1_11_in16 = reg_0141;
    64: op1_11_in16 = reg_0153;
    66: op1_11_in16 = reg_0182;
    67: op1_11_in16 = reg_0405;
    68: op1_11_in16 = reg_0914;
    69: op1_11_in16 = imem04_in[87:84];
    71: op1_11_in16 = imem01_in[51:48];
    72: op1_11_in16 = imem06_in[15:12];
    75: op1_11_in16 = reg_0204;
    76: op1_11_in16 = reg_0054;
    77: op1_11_in16 = reg_0055;
    78: op1_11_in16 = reg_0027;
    79: op1_11_in16 = imem06_in[51:48];
    81: op1_11_in16 = reg_0472;
    82: op1_11_in16 = reg_0002;
    83: op1_11_in16 = reg_0295;
    84: op1_11_in16 = imem02_in[87:84];
    86: op1_11_in16 = reg_0475;
    87: op1_11_in16 = reg_0658;
    88: op1_11_in16 = reg_0247;
    89: op1_11_in16 = reg_0395;
    90: op1_11_in16 = reg_0036;
    91: op1_11_in16 = reg_0719;
    92: op1_11_in16 = imem01_in[59:56];
    93: op1_11_in16 = reg_0359;
    94: op1_11_in16 = reg_0394;
    95: op1_11_in16 = reg_0886;
    96: op1_11_in16 = reg_0650;
    default: op1_11_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv16 = 1;
    7: op1_11_inv16 = 1;
    12: op1_11_inv16 = 1;
    17: op1_11_inv16 = 1;
    18: op1_11_inv16 = 1;
    19: op1_11_inv16 = 1;
    20: op1_11_inv16 = 1;
    24: op1_11_inv16 = 1;
    26: op1_11_inv16 = 1;
    28: op1_11_inv16 = 1;
    31: op1_11_inv16 = 1;
    32: op1_11_inv16 = 1;
    33: op1_11_inv16 = 1;
    45: op1_11_inv16 = 1;
    47: op1_11_inv16 = 1;
    48: op1_11_inv16 = 1;
    49: op1_11_inv16 = 1;
    50: op1_11_inv16 = 1;
    51: op1_11_inv16 = 1;
    52: op1_11_inv16 = 1;
    54: op1_11_inv16 = 1;
    61: op1_11_inv16 = 1;
    63: op1_11_inv16 = 1;
    65: op1_11_inv16 = 1;
    68: op1_11_inv16 = 1;
    69: op1_11_inv16 = 1;
    75: op1_11_inv16 = 1;
    77: op1_11_inv16 = 1;
    78: op1_11_inv16 = 1;
    79: op1_11_inv16 = 1;
    85: op1_11_inv16 = 1;
    86: op1_11_inv16 = 1;
    89: op1_11_inv16 = 1;
    90: op1_11_inv16 = 1;
    92: op1_11_inv16 = 1;
    94: op1_11_inv16 = 1;
    95: op1_11_inv16 = 1;
    default: op1_11_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in17 = reg_0317;
    6: op1_11_in17 = reg_0648;
    7: op1_11_in17 = reg_0970;
    9: op1_11_in17 = reg_0583;
    10: op1_11_in17 = reg_0777;
    11: op1_11_in17 = imem05_in[35:32];
    12: op1_11_in17 = reg_0203;
    13: op1_11_in17 = reg_0251;
    14: op1_11_in17 = reg_0440;
    15: op1_11_in17 = reg_0478;
    16: op1_11_in17 = imem04_in[63:60];
    17: op1_11_in17 = reg_0611;
    18: op1_11_in17 = reg_0542;
    19: op1_11_in17 = reg_0134;
    63: op1_11_in17 = reg_0134;
    20: op1_11_in17 = imem04_in[111:108];
    21: op1_11_in17 = reg_0723;
    22: op1_11_in17 = imem02_in[79:76];
    23: op1_11_in17 = reg_0591;
    24: op1_11_in17 = reg_0666;
    25: op1_11_in17 = reg_0530;
    26: op1_11_in17 = imem01_in[63:60];
    92: op1_11_in17 = imem01_in[63:60];
    27: op1_11_in17 = reg_0819;
    28: op1_11_in17 = reg_0947;
    29: op1_11_in17 = imem03_in[3:0];
    30: op1_11_in17 = reg_0312;
    31: op1_11_in17 = reg_0295;
    32: op1_11_in17 = reg_0452;
    33: op1_11_in17 = reg_0191;
    34: op1_11_in17 = reg_1057;
    37: op1_11_in17 = reg_1031;
    39: op1_11_in17 = imem03_in[67:64];
    40: op1_11_in17 = imem04_in[91:88];
    69: op1_11_in17 = imem04_in[91:88];
    41: op1_11_in17 = reg_0313;
    43: op1_11_in17 = reg_0242;
    44: op1_11_in17 = reg_0086;
    62: op1_11_in17 = reg_0086;
    45: op1_11_in17 = reg_0222;
    47: op1_11_in17 = imem03_in[11:8];
    48: op1_11_in17 = reg_0381;
    49: op1_11_in17 = reg_0179;
    50: op1_11_in17 = imem05_in[87:84];
    51: op1_11_in17 = reg_0584;
    52: op1_11_in17 = reg_0506;
    53: op1_11_in17 = reg_0507;
    54: op1_11_in17 = imem04_in[51:48];
    55: op1_11_in17 = imem07_in[15:12];
    57: op1_11_in17 = reg_0421;
    58: op1_11_in17 = reg_0705;
    61: op1_11_in17 = imem01_in[7:4];
    64: op1_11_in17 = imem06_in[11:8];
    65: op1_11_in17 = imem07_in[51:48];
    66: op1_11_in17 = reg_0170;
    67: op1_11_in17 = reg_0264;
    68: op1_11_in17 = reg_0323;
    71: op1_11_in17 = reg_0105;
    72: op1_11_in17 = imem06_in[59:56];
    79: op1_11_in17 = imem06_in[59:56];
    75: op1_11_in17 = reg_0211;
    76: op1_11_in17 = reg_0347;
    77: op1_11_in17 = reg_0050;
    78: op1_11_in17 = imem05_in[23:20];
    81: op1_11_in17 = reg_0459;
    82: op1_11_in17 = reg_0047;
    83: op1_11_in17 = reg_0856;
    84: op1_11_in17 = imem02_in[103:100];
    85: op1_11_in17 = reg_0640;
    86: op1_11_in17 = reg_0480;
    87: op1_11_in17 = reg_0065;
    88: op1_11_in17 = reg_0718;
    89: op1_11_in17 = reg_0292;
    90: op1_11_in17 = reg_0403;
    91: op1_11_in17 = reg_0084;
    93: op1_11_in17 = reg_0329;
    94: op1_11_in17 = reg_0389;
    95: op1_11_in17 = reg_0218;
    96: op1_11_in17 = reg_0365;
    default: op1_11_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv17 = 1;
    7: op1_11_inv17 = 1;
    9: op1_11_inv17 = 1;
    10: op1_11_inv17 = 1;
    11: op1_11_inv17 = 1;
    13: op1_11_inv17 = 1;
    15: op1_11_inv17 = 1;
    16: op1_11_inv17 = 1;
    17: op1_11_inv17 = 1;
    18: op1_11_inv17 = 1;
    21: op1_11_inv17 = 1;
    22: op1_11_inv17 = 1;
    23: op1_11_inv17 = 1;
    24: op1_11_inv17 = 1;
    25: op1_11_inv17 = 1;
    27: op1_11_inv17 = 1;
    29: op1_11_inv17 = 1;
    34: op1_11_inv17 = 1;
    37: op1_11_inv17 = 1;
    40: op1_11_inv17 = 1;
    44: op1_11_inv17 = 1;
    45: op1_11_inv17 = 1;
    47: op1_11_inv17 = 1;
    50: op1_11_inv17 = 1;
    55: op1_11_inv17 = 1;
    61: op1_11_inv17 = 1;
    62: op1_11_inv17 = 1;
    64: op1_11_inv17 = 1;
    66: op1_11_inv17 = 1;
    67: op1_11_inv17 = 1;
    69: op1_11_inv17 = 1;
    75: op1_11_inv17 = 1;
    76: op1_11_inv17 = 1;
    77: op1_11_inv17 = 1;
    78: op1_11_inv17 = 1;
    81: op1_11_inv17 = 1;
    84: op1_11_inv17 = 1;
    87: op1_11_inv17 = 1;
    88: op1_11_inv17 = 1;
    89: op1_11_inv17 = 1;
    91: op1_11_inv17 = 1;
    92: op1_11_inv17 = 1;
    94: op1_11_inv17 = 1;
    95: op1_11_inv17 = 1;
    default: op1_11_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in18 = reg_0012;
    6: op1_11_in18 = reg_0662;
    7: op1_11_in18 = reg_0971;
    9: op1_11_in18 = reg_0587;
    10: op1_11_in18 = reg_0775;
    11: op1_11_in18 = imem05_in[39:36];
    12: op1_11_in18 = reg_0193;
    13: op1_11_in18 = reg_0836;
    14: op1_11_in18 = reg_0442;
    15: op1_11_in18 = reg_0214;
    16: op1_11_in18 = imem04_in[95:92];
    17: op1_11_in18 = reg_0577;
    18: op1_11_in18 = reg_0540;
    19: op1_11_in18 = imem06_in[7:4];
    20: op1_11_in18 = imem04_in[123:120];
    21: op1_11_in18 = reg_0702;
    22: op1_11_in18 = imem02_in[115:112];
    23: op1_11_in18 = reg_0563;
    24: op1_11_in18 = reg_0654;
    25: op1_11_in18 = reg_0277;
    26: op1_11_in18 = imem01_in[67:64];
    27: op1_11_in18 = reg_0831;
    28: op1_11_in18 = reg_0972;
    29: op1_11_in18 = imem03_in[35:32];
    30: op1_11_in18 = reg_0844;
    31: op1_11_in18 = imem07_in[7:4];
    32: op1_11_in18 = reg_0188;
    33: op1_11_in18 = reg_0188;
    34: op1_11_in18 = reg_0050;
    37: op1_11_in18 = reg_0228;
    39: op1_11_in18 = imem03_in[83:80];
    40: op1_11_in18 = imem04_in[107:104];
    41: op1_11_in18 = reg_0764;
    43: op1_11_in18 = reg_0274;
    44: op1_11_in18 = reg_0016;
    45: op1_11_in18 = reg_0780;
    47: op1_11_in18 = imem03_in[91:88];
    48: op1_11_in18 = reg_0264;
    49: op1_11_in18 = reg_0169;
    50: op1_11_in18 = imem05_in[91:88];
    51: op1_11_in18 = reg_0064;
    52: op1_11_in18 = reg_0261;
    53: op1_11_in18 = reg_0276;
    54: op1_11_in18 = imem04_in[59:56];
    55: op1_11_in18 = imem07_in[47:44];
    57: op1_11_in18 = reg_0321;
    58: op1_11_in18 = reg_0707;
    61: op1_11_in18 = imem01_in[75:72];
    62: op1_11_in18 = reg_0484;
    63: op1_11_in18 = imem06_in[43:40];
    64: op1_11_in18 = imem06_in[35:32];
    65: op1_11_in18 = imem07_in[63:60];
    67: op1_11_in18 = reg_0916;
    68: op1_11_in18 = reg_0358;
    69: op1_11_in18 = reg_1004;
    71: op1_11_in18 = reg_1032;
    72: op1_11_in18 = imem06_in[67:64];
    75: op1_11_in18 = reg_0186;
    76: op1_11_in18 = reg_0761;
    77: op1_11_in18 = reg_0067;
    78: op1_11_in18 = imem05_in[55:52];
    79: op1_11_in18 = imem06_in[87:84];
    81: op1_11_in18 = reg_0478;
    82: op1_11_in18 = imem07_in[19:16];
    83: op1_11_in18 = imem05_in[3:0];
    84: op1_11_in18 = reg_0645;
    85: op1_11_in18 = reg_0703;
    86: op1_11_in18 = reg_0473;
    87: op1_11_in18 = reg_0552;
    88: op1_11_in18 = reg_0805;
    89: op1_11_in18 = reg_0888;
    90: op1_11_in18 = reg_0804;
    91: op1_11_in18 = reg_0222;
    92: op1_11_in18 = imem01_in[91:88];
    93: op1_11_in18 = reg_0394;
    94: op1_11_in18 = reg_0425;
    95: op1_11_in18 = imem03_in[7:4];
    96: op1_11_in18 = imem03_in[47:44];
    default: op1_11_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv18 = 1;
    10: op1_11_inv18 = 1;
    11: op1_11_inv18 = 1;
    13: op1_11_inv18 = 1;
    14: op1_11_inv18 = 1;
    18: op1_11_inv18 = 1;
    21: op1_11_inv18 = 1;
    25: op1_11_inv18 = 1;
    26: op1_11_inv18 = 1;
    28: op1_11_inv18 = 1;
    30: op1_11_inv18 = 1;
    33: op1_11_inv18 = 1;
    34: op1_11_inv18 = 1;
    40: op1_11_inv18 = 1;
    43: op1_11_inv18 = 1;
    47: op1_11_inv18 = 1;
    48: op1_11_inv18 = 1;
    52: op1_11_inv18 = 1;
    53: op1_11_inv18 = 1;
    57: op1_11_inv18 = 1;
    58: op1_11_inv18 = 1;
    61: op1_11_inv18 = 1;
    63: op1_11_inv18 = 1;
    71: op1_11_inv18 = 1;
    72: op1_11_inv18 = 1;
    76: op1_11_inv18 = 1;
    78: op1_11_inv18 = 1;
    81: op1_11_inv18 = 1;
    82: op1_11_inv18 = 1;
    83: op1_11_inv18 = 1;
    85: op1_11_inv18 = 1;
    86: op1_11_inv18 = 1;
    88: op1_11_inv18 = 1;
    89: op1_11_inv18 = 1;
    91: op1_11_inv18 = 1;
    93: op1_11_inv18 = 1;
    default: op1_11_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in19 = reg_0002;
    6: op1_11_in19 = reg_0644;
    94: op1_11_in19 = reg_0644;
    7: op1_11_in19 = reg_0946;
    9: op1_11_in19 = reg_0388;
    10: op1_11_in19 = reg_0792;
    11: op1_11_in19 = imem05_in[123:120];
    12: op1_11_in19 = reg_0207;
    13: op1_11_in19 = reg_0152;
    14: op1_11_in19 = reg_0437;
    15: op1_11_in19 = reg_0191;
    16: op1_11_in19 = imem04_in[115:112];
    17: op1_11_in19 = reg_0408;
    18: op1_11_in19 = reg_0558;
    19: op1_11_in19 = imem06_in[47:44];
    20: op1_11_in19 = reg_0553;
    21: op1_11_in19 = reg_0709;
    22: op1_11_in19 = imem02_in[123:120];
    23: op1_11_in19 = reg_0595;
    24: op1_11_in19 = reg_0646;
    25: op1_11_in19 = reg_0306;
    26: op1_11_in19 = reg_0299;
    27: op1_11_in19 = reg_0140;
    28: op1_11_in19 = reg_0900;
    29: op1_11_in19 = imem03_in[63:60];
    30: op1_11_in19 = reg_0996;
    31: op1_11_in19 = imem07_in[43:40];
    32: op1_11_in19 = reg_0211;
    33: op1_11_in19 = imem01_in[23:20];
    34: op1_11_in19 = reg_0268;
    37: op1_11_in19 = reg_1018;
    39: op1_11_in19 = reg_0938;
    40: op1_11_in19 = reg_1004;
    41: op1_11_in19 = reg_0061;
    43: op1_11_in19 = reg_0487;
    44: op1_11_in19 = imem03_in[27:24];
    95: op1_11_in19 = imem03_in[27:24];
    45: op1_11_in19 = reg_0609;
    47: op1_11_in19 = imem03_in[127:124];
    48: op1_11_in19 = reg_0383;
    49: op1_11_in19 = reg_0170;
    50: op1_11_in19 = reg_0150;
    51: op1_11_in19 = reg_0281;
    52: op1_11_in19 = imem03_in[11:8];
    53: op1_11_in19 = reg_0401;
    54: op1_11_in19 = imem04_in[91:88];
    55: op1_11_in19 = imem07_in[83:80];
    57: op1_11_in19 = reg_0599;
    58: op1_11_in19 = reg_0706;
    61: op1_11_in19 = imem01_in[79:76];
    62: op1_11_in19 = imem03_in[59:56];
    63: op1_11_in19 = imem06_in[67:64];
    64: op1_11_in19 = imem06_in[39:36];
    65: op1_11_in19 = imem07_in[67:64];
    67: op1_11_in19 = reg_0955;
    68: op1_11_in19 = reg_0081;
    69: op1_11_in19 = reg_0912;
    71: op1_11_in19 = reg_1035;
    72: op1_11_in19 = imem06_in[71:68];
    75: op1_11_in19 = reg_0196;
    76: op1_11_in19 = reg_0085;
    77: op1_11_in19 = reg_0056;
    78: op1_11_in19 = imem05_in[83:80];
    79: op1_11_in19 = imem06_in[107:104];
    81: op1_11_in19 = reg_0203;
    82: op1_11_in19 = imem07_in[27:24];
    83: op1_11_in19 = imem05_in[59:56];
    84: op1_11_in19 = reg_0323;
    85: op1_11_in19 = reg_0339;
    86: op1_11_in19 = reg_0470;
    87: op1_11_in19 = reg_0027;
    88: op1_11_in19 = reg_0433;
    89: op1_11_in19 = reg_0850;
    90: op1_11_in19 = reg_0222;
    91: op1_11_in19 = imem07_in[19:16];
    92: op1_11_in19 = imem01_in[119:116];
    93: op1_11_in19 = reg_0372;
    96: op1_11_in19 = imem03_in[75:72];
    default: op1_11_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv19 = 1;
    7: op1_11_inv19 = 1;
    11: op1_11_inv19 = 1;
    12: op1_11_inv19 = 1;
    13: op1_11_inv19 = 1;
    16: op1_11_inv19 = 1;
    17: op1_11_inv19 = 1;
    18: op1_11_inv19 = 1;
    21: op1_11_inv19 = 1;
    23: op1_11_inv19 = 1;
    27: op1_11_inv19 = 1;
    28: op1_11_inv19 = 1;
    34: op1_11_inv19 = 1;
    39: op1_11_inv19 = 1;
    44: op1_11_inv19 = 1;
    45: op1_11_inv19 = 1;
    48: op1_11_inv19 = 1;
    49: op1_11_inv19 = 1;
    50: op1_11_inv19 = 1;
    51: op1_11_inv19 = 1;
    52: op1_11_inv19 = 1;
    53: op1_11_inv19 = 1;
    55: op1_11_inv19 = 1;
    57: op1_11_inv19 = 1;
    58: op1_11_inv19 = 1;
    62: op1_11_inv19 = 1;
    69: op1_11_inv19 = 1;
    71: op1_11_inv19 = 1;
    75: op1_11_inv19 = 1;
    76: op1_11_inv19 = 1;
    77: op1_11_inv19 = 1;
    78: op1_11_inv19 = 1;
    81: op1_11_inv19 = 1;
    82: op1_11_inv19 = 1;
    85: op1_11_inv19 = 1;
    88: op1_11_inv19 = 1;
    89: op1_11_inv19 = 1;
    93: op1_11_inv19 = 1;
    95: op1_11_inv19 = 1;
    96: op1_11_inv19 = 1;
    default: op1_11_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in20 = reg_0013;
    6: op1_11_in20 = reg_0643;
    7: op1_11_in20 = reg_0961;
    9: op1_11_in20 = reg_0327;
    10: op1_11_in20 = reg_0519;
    11: op1_11_in20 = reg_0973;
    12: op1_11_in20 = reg_0198;
    32: op1_11_in20 = reg_0198;
    13: op1_11_in20 = reg_0142;
    14: op1_11_in20 = reg_0179;
    15: op1_11_in20 = reg_0204;
    16: op1_11_in20 = imem04_in[119:116];
    54: op1_11_in20 = imem04_in[119:116];
    17: op1_11_in20 = reg_0349;
    18: op1_11_in20 = reg_0556;
    19: op1_11_in20 = imem06_in[63:60];
    20: op1_11_in20 = reg_0546;
    21: op1_11_in20 = reg_0713;
    22: op1_11_in20 = reg_0655;
    23: op1_11_in20 = reg_0384;
    24: op1_11_in20 = reg_0657;
    25: op1_11_in20 = reg_1020;
    26: op1_11_in20 = reg_0810;
    27: op1_11_in20 = imem06_in[15:12];
    28: op1_11_in20 = reg_0757;
    29: op1_11_in20 = imem03_in[67:64];
    30: op1_11_in20 = reg_1001;
    31: op1_11_in20 = imem07_in[63:60];
    33: op1_11_in20 = imem01_in[31:28];
    34: op1_11_in20 = reg_0068;
    37: op1_11_in20 = reg_1034;
    39: op1_11_in20 = reg_0824;
    40: op1_11_in20 = reg_0483;
    41: op1_11_in20 = reg_0755;
    43: op1_11_in20 = reg_0249;
    44: op1_11_in20 = imem03_in[71:68];
    45: op1_11_in20 = reg_0622;
    47: op1_11_in20 = reg_0940;
    48: op1_11_in20 = reg_0629;
    49: op1_11_in20 = reg_0158;
    50: op1_11_in20 = reg_0154;
    51: op1_11_in20 = reg_0834;
    52: op1_11_in20 = imem03_in[23:20];
    53: op1_11_in20 = reg_0288;
    55: op1_11_in20 = reg_0719;
    57: op1_11_in20 = reg_0420;
    58: op1_11_in20 = reg_0700;
    61: op1_11_in20 = imem01_in[107:104];
    62: op1_11_in20 = imem03_in[123:120];
    63: op1_11_in20 = imem06_in[123:120];
    64: op1_11_in20 = imem06_in[43:40];
    65: op1_11_in20 = imem07_in[71:68];
    67: op1_11_in20 = imem07_in[23:20];
    68: op1_11_in20 = reg_0052;
    84: op1_11_in20 = reg_0052;
    69: op1_11_in20 = reg_0537;
    71: op1_11_in20 = reg_0793;
    72: op1_11_in20 = imem06_in[75:72];
    75: op1_11_in20 = imem01_in[7:4];
    76: op1_11_in20 = reg_0291;
    77: op1_11_in20 = reg_0764;
    78: op1_11_in20 = reg_0826;
    79: op1_11_in20 = imem06_in[111:108];
    81: op1_11_in20 = reg_0212;
    82: op1_11_in20 = imem07_in[79:76];
    83: op1_11_in20 = imem05_in[71:68];
    86: op1_11_in20 = reg_0459;
    87: op1_11_in20 = reg_0854;
    88: op1_11_in20 = reg_0426;
    89: op1_11_in20 = reg_0067;
    90: op1_11_in20 = imem07_in[3:0];
    91: op1_11_in20 = imem07_in[75:72];
    92: op1_11_in20 = reg_0246;
    93: op1_11_in20 = reg_0248;
    94: op1_11_in20 = reg_0347;
    95: op1_11_in20 = imem03_in[63:60];
    96: op1_11_in20 = imem03_in[103:100];
    default: op1_11_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv20 = 1;
    6: op1_11_inv20 = 1;
    9: op1_11_inv20 = 1;
    12: op1_11_inv20 = 1;
    14: op1_11_inv20 = 1;
    15: op1_11_inv20 = 1;
    16: op1_11_inv20 = 1;
    17: op1_11_inv20 = 1;
    18: op1_11_inv20 = 1;
    19: op1_11_inv20 = 1;
    21: op1_11_inv20 = 1;
    22: op1_11_inv20 = 1;
    23: op1_11_inv20 = 1;
    27: op1_11_inv20 = 1;
    28: op1_11_inv20 = 1;
    29: op1_11_inv20 = 1;
    31: op1_11_inv20 = 1;
    32: op1_11_inv20 = 1;
    33: op1_11_inv20 = 1;
    34: op1_11_inv20 = 1;
    37: op1_11_inv20 = 1;
    39: op1_11_inv20 = 1;
    40: op1_11_inv20 = 1;
    44: op1_11_inv20 = 1;
    51: op1_11_inv20 = 1;
    52: op1_11_inv20 = 1;
    53: op1_11_inv20 = 1;
    62: op1_11_inv20 = 1;
    64: op1_11_inv20 = 1;
    67: op1_11_inv20 = 1;
    68: op1_11_inv20 = 1;
    69: op1_11_inv20 = 1;
    77: op1_11_inv20 = 1;
    81: op1_11_inv20 = 1;
    86: op1_11_inv20 = 1;
    87: op1_11_inv20 = 1;
    88: op1_11_inv20 = 1;
    91: op1_11_inv20 = 1;
    92: op1_11_inv20 = 1;
    93: op1_11_inv20 = 1;
    94: op1_11_inv20 = 1;
    default: op1_11_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in21 = reg_0014;
    6: op1_11_in21 = reg_0663;
    7: op1_11_in21 = reg_0250;
    9: op1_11_in21 = reg_0396;
    10: op1_11_in21 = reg_0517;
    11: op1_11_in21 = reg_0948;
    12: op1_11_in21 = reg_0201;
    32: op1_11_in21 = reg_0201;
    13: op1_11_in21 = reg_0146;
    14: op1_11_in21 = reg_0161;
    15: op1_11_in21 = reg_0188;
    16: op1_11_in21 = imem04_in[127:124];
    17: op1_11_in21 = reg_0409;
    18: op1_11_in21 = reg_0308;
    19: op1_11_in21 = imem06_in[91:88];
    20: op1_11_in21 = reg_0540;
    21: op1_11_in21 = reg_0430;
    22: op1_11_in21 = reg_0654;
    23: op1_11_in21 = reg_0373;
    24: op1_11_in21 = reg_0656;
    25: op1_11_in21 = reg_0050;
    26: op1_11_in21 = reg_0828;
    27: op1_11_in21 = imem06_in[75:72];
    28: op1_11_in21 = reg_0260;
    29: op1_11_in21 = imem03_in[75:72];
    44: op1_11_in21 = imem03_in[75:72];
    30: op1_11_in21 = reg_0974;
    31: op1_11_in21 = imem07_in[107:104];
    33: op1_11_in21 = imem01_in[59:56];
    34: op1_11_in21 = reg_0047;
    37: op1_11_in21 = reg_0105;
    39: op1_11_in21 = reg_0389;
    40: op1_11_in21 = reg_1006;
    41: op1_11_in21 = reg_0009;
    43: op1_11_in21 = reg_0501;
    45: op1_11_in21 = imem07_in[3:0];
    47: op1_11_in21 = reg_0535;
    48: op1_11_in21 = reg_0309;
    50: op1_11_in21 = reg_0143;
    51: op1_11_in21 = reg_0899;
    52: op1_11_in21 = imem03_in[47:44];
    53: op1_11_in21 = reg_0732;
    54: op1_11_in21 = reg_1004;
    55: op1_11_in21 = reg_0714;
    57: op1_11_in21 = reg_0502;
    58: op1_11_in21 = reg_0303;
    61: op1_11_in21 = imem01_in[111:108];
    62: op1_11_in21 = reg_0357;
    63: op1_11_in21 = reg_1019;
    64: op1_11_in21 = imem06_in[71:68];
    65: op1_11_in21 = imem07_in[75:72];
    67: op1_11_in21 = imem07_in[87:84];
    68: op1_11_in21 = reg_0423;
    84: op1_11_in21 = reg_0423;
    69: op1_11_in21 = reg_0909;
    71: op1_11_in21 = reg_0862;
    72: op1_11_in21 = imem06_in[79:76];
    75: op1_11_in21 = imem01_in[43:40];
    76: op1_11_in21 = imem03_in[19:16];
    77: op1_11_in21 = reg_0432;
    78: op1_11_in21 = reg_0226;
    79: op1_11_in21 = imem06_in[123:120];
    81: op1_11_in21 = reg_0202;
    82: op1_11_in21 = imem07_in[111:108];
    83: op1_11_in21 = imem05_in[79:76];
    86: op1_11_in21 = reg_0209;
    87: op1_11_in21 = reg_0295;
    88: op1_11_in21 = reg_0419;
    89: op1_11_in21 = reg_0401;
    90: op1_11_in21 = imem07_in[7:4];
    91: op1_11_in21 = imem07_in[103:100];
    92: op1_11_in21 = reg_1014;
    93: op1_11_in21 = reg_0516;
    94: op1_11_in21 = reg_0650;
    95: op1_11_in21 = imem03_in[67:64];
    96: op1_11_in21 = imem03_in[127:124];
    default: op1_11_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_11_inv21 = 1;
    14: op1_11_inv21 = 1;
    15: op1_11_inv21 = 1;
    16: op1_11_inv21 = 1;
    18: op1_11_inv21 = 1;
    19: op1_11_inv21 = 1;
    20: op1_11_inv21 = 1;
    21: op1_11_inv21 = 1;
    24: op1_11_inv21 = 1;
    25: op1_11_inv21 = 1;
    27: op1_11_inv21 = 1;
    28: op1_11_inv21 = 1;
    29: op1_11_inv21 = 1;
    33: op1_11_inv21 = 1;
    37: op1_11_inv21 = 1;
    41: op1_11_inv21 = 1;
    43: op1_11_inv21 = 1;
    47: op1_11_inv21 = 1;
    48: op1_11_inv21 = 1;
    52: op1_11_inv21 = 1;
    57: op1_11_inv21 = 1;
    58: op1_11_inv21 = 1;
    61: op1_11_inv21 = 1;
    62: op1_11_inv21 = 1;
    63: op1_11_inv21 = 1;
    65: op1_11_inv21 = 1;
    67: op1_11_inv21 = 1;
    68: op1_11_inv21 = 1;
    69: op1_11_inv21 = 1;
    72: op1_11_inv21 = 1;
    75: op1_11_inv21 = 1;
    78: op1_11_inv21 = 1;
    82: op1_11_inv21 = 1;
    88: op1_11_inv21 = 1;
    89: op1_11_inv21 = 1;
    90: op1_11_inv21 = 1;
    92: op1_11_inv21 = 1;
    93: op1_11_inv21 = 1;
    94: op1_11_inv21 = 1;
    96: op1_11_inv21 = 1;
    default: op1_11_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in22 = reg_0015;
    6: op1_11_in22 = reg_0359;
    7: op1_11_in22 = reg_0152;
    9: op1_11_in22 = reg_0389;
    10: op1_11_in22 = reg_0515;
    11: op1_11_in22 = reg_0942;
    12: op1_11_in22 = reg_0197;
    81: op1_11_in22 = reg_0197;
    13: op1_11_in22 = reg_0137;
    14: op1_11_in22 = reg_0160;
    15: op1_11_in22 = reg_0212;
    16: op1_11_in22 = reg_0543;
    17: op1_11_in22 = reg_0375;
    18: op1_11_in22 = reg_0301;
    19: op1_11_in22 = imem06_in[99:96];
    20: op1_11_in22 = reg_0558;
    21: op1_11_in22 = reg_0426;
    22: op1_11_in22 = reg_0637;
    23: op1_11_in22 = reg_0396;
    24: op1_11_in22 = reg_0649;
    25: op1_11_in22 = reg_0313;
    26: op1_11_in22 = reg_0236;
    27: op1_11_in22 = imem06_in[107:104];
    28: op1_11_in22 = reg_0825;
    29: op1_11_in22 = imem03_in[99:96];
    44: op1_11_in22 = imem03_in[99:96];
    30: op1_11_in22 = reg_0981;
    31: op1_11_in22 = reg_0721;
    32: op1_11_in22 = reg_0213;
    33: op1_11_in22 = imem01_in[83:80];
    34: op1_11_in22 = reg_0043;
    37: op1_11_in22 = reg_0124;
    39: op1_11_in22 = reg_1001;
    40: op1_11_in22 = reg_0937;
    41: op1_11_in22 = reg_0059;
    43: op1_11_in22 = reg_0798;
    45: op1_11_in22 = imem07_in[103:100];
    47: op1_11_in22 = reg_1050;
    48: op1_11_in22 = imem07_in[47:44];
    50: op1_11_in22 = reg_0153;
    51: op1_11_in22 = reg_0593;
    52: op1_11_in22 = imem03_in[55:52];
    53: op1_11_in22 = reg_0078;
    54: op1_11_in22 = reg_0931;
    55: op1_11_in22 = reg_0729;
    57: op1_11_in22 = reg_0180;
    58: op1_11_in22 = reg_0315;
    61: op1_11_in22 = reg_0242;
    62: op1_11_in22 = reg_1007;
    63: op1_11_in22 = reg_0696;
    64: op1_11_in22 = imem06_in[83:80];
    65: op1_11_in22 = imem07_in[83:80];
    67: op1_11_in22 = imem07_in[111:108];
    68: op1_11_in22 = reg_0394;
    69: op1_11_in22 = reg_0752;
    71: op1_11_in22 = reg_0604;
    72: op1_11_in22 = reg_0010;
    75: op1_11_in22 = reg_1032;
    76: op1_11_in22 = imem03_in[35:32];
    77: op1_11_in22 = reg_0856;
    78: op1_11_in22 = reg_0256;
    79: op1_11_in22 = reg_0691;
    83: op1_11_in22 = imem05_in[95:92];
    84: op1_11_in22 = reg_0372;
    86: op1_11_in22 = reg_0207;
    87: op1_11_in22 = reg_0966;
    88: op1_11_in22 = reg_0174;
    89: op1_11_in22 = reg_0815;
    90: op1_11_in22 = imem07_in[23:20];
    91: op1_11_in22 = imem07_in[107:104];
    92: op1_11_in22 = reg_1035;
    93: op1_11_in22 = reg_0347;
    94: op1_11_in22 = reg_0734;
    95: op1_11_in22 = imem03_in[79:76];
    96: op1_11_in22 = reg_0819;
    default: op1_11_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv22 = 1;
    6: op1_11_inv22 = 1;
    10: op1_11_inv22 = 1;
    17: op1_11_inv22 = 1;
    19: op1_11_inv22 = 1;
    20: op1_11_inv22 = 1;
    21: op1_11_inv22 = 1;
    23: op1_11_inv22 = 1;
    24: op1_11_inv22 = 1;
    25: op1_11_inv22 = 1;
    28: op1_11_inv22 = 1;
    29: op1_11_inv22 = 1;
    30: op1_11_inv22 = 1;
    32: op1_11_inv22 = 1;
    33: op1_11_inv22 = 1;
    34: op1_11_inv22 = 1;
    40: op1_11_inv22 = 1;
    41: op1_11_inv22 = 1;
    47: op1_11_inv22 = 1;
    48: op1_11_inv22 = 1;
    50: op1_11_inv22 = 1;
    51: op1_11_inv22 = 1;
    52: op1_11_inv22 = 1;
    53: op1_11_inv22 = 1;
    55: op1_11_inv22 = 1;
    57: op1_11_inv22 = 1;
    61: op1_11_inv22 = 1;
    64: op1_11_inv22 = 1;
    67: op1_11_inv22 = 1;
    69: op1_11_inv22 = 1;
    71: op1_11_inv22 = 1;
    76: op1_11_inv22 = 1;
    78: op1_11_inv22 = 1;
    86: op1_11_inv22 = 1;
    87: op1_11_inv22 = 1;
    90: op1_11_inv22 = 1;
    91: op1_11_inv22 = 1;
    92: op1_11_inv22 = 1;
    93: op1_11_inv22 = 1;
    96: op1_11_inv22 = 1;
    default: op1_11_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in23 = reg_0016;
    6: op1_11_in23 = reg_0083;
    7: op1_11_in23 = reg_0130;
    9: op1_11_in23 = reg_0982;
    10: op1_11_in23 = imem01_in[7:4];
    32: op1_11_in23 = imem01_in[7:4];
    81: op1_11_in23 = imem01_in[7:4];
    11: op1_11_in23 = reg_0968;
    12: op1_11_in23 = imem01_in[27:24];
    13: op1_11_in23 = reg_0134;
    14: op1_11_in23 = reg_0164;
    15: op1_11_in23 = reg_0195;
    16: op1_11_in23 = reg_0529;
    17: op1_11_in23 = reg_0404;
    18: op1_11_in23 = reg_0305;
    19: op1_11_in23 = imem06_in[127:124];
    20: op1_11_in23 = reg_0541;
    21: op1_11_in23 = reg_0423;
    22: op1_11_in23 = reg_0656;
    94: op1_11_in23 = reg_0656;
    23: op1_11_in23 = reg_1002;
    24: op1_11_in23 = reg_0641;
    25: op1_11_in23 = reg_0764;
    26: op1_11_in23 = reg_0248;
    27: op1_11_in23 = imem06_in[111:108];
    28: op1_11_in23 = reg_0142;
    29: op1_11_in23 = reg_0602;
    30: op1_11_in23 = reg_1000;
    39: op1_11_in23 = reg_1000;
    31: op1_11_in23 = reg_0718;
    33: op1_11_in23 = reg_0786;
    34: op1_11_in23 = reg_0855;
    37: op1_11_in23 = reg_0116;
    40: op1_11_in23 = reg_0539;
    41: op1_11_in23 = reg_0854;
    43: op1_11_in23 = reg_0604;
    44: op1_11_in23 = imem03_in[127:124];
    45: op1_11_in23 = imem07_in[111:108];
    47: op1_11_in23 = reg_0357;
    48: op1_11_in23 = imem07_in[51:48];
    50: op1_11_in23 = reg_0140;
    51: op1_11_in23 = reg_0031;
    52: op1_11_in23 = imem03_in[63:60];
    53: op1_11_in23 = reg_0578;
    54: op1_11_in23 = reg_0752;
    55: op1_11_in23 = reg_0713;
    57: op1_11_in23 = reg_0178;
    58: op1_11_in23 = reg_0353;
    61: op1_11_in23 = reg_0870;
    62: op1_11_in23 = reg_0576;
    63: op1_11_in23 = reg_0889;
    64: op1_11_in23 = imem06_in[87:84];
    65: op1_11_in23 = imem07_in[123:120];
    67: op1_11_in23 = reg_0719;
    68: op1_11_in23 = reg_0037;
    69: op1_11_in23 = reg_0076;
    71: op1_11_in23 = reg_0902;
    72: op1_11_in23 = reg_1019;
    75: op1_11_in23 = reg_1023;
    76: op1_11_in23 = imem03_in[59:56];
    77: op1_11_in23 = reg_0044;
    78: op1_11_in23 = reg_0941;
    79: op1_11_in23 = reg_1018;
    83: op1_11_in23 = imem05_in[107:104];
    84: op1_11_in23 = reg_0347;
    86: op1_11_in23 = reg_0194;
    87: op1_11_in23 = reg_0611;
    88: op1_11_in23 = reg_0172;
    89: op1_11_in23 = reg_0072;
    90: op1_11_in23 = imem07_in[27:24];
    91: op1_11_in23 = imem07_in[115:112];
    92: op1_11_in23 = reg_0503;
    93: op1_11_in23 = reg_0734;
    95: op1_11_in23 = imem03_in[95:92];
    96: op1_11_in23 = reg_0784;
    default: op1_11_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv23 = 1;
    6: op1_11_inv23 = 1;
    9: op1_11_inv23 = 1;
    16: op1_11_inv23 = 1;
    17: op1_11_inv23 = 1;
    19: op1_11_inv23 = 1;
    21: op1_11_inv23 = 1;
    22: op1_11_inv23 = 1;
    23: op1_11_inv23 = 1;
    24: op1_11_inv23 = 1;
    25: op1_11_inv23 = 1;
    28: op1_11_inv23 = 1;
    29: op1_11_inv23 = 1;
    31: op1_11_inv23 = 1;
    33: op1_11_inv23 = 1;
    39: op1_11_inv23 = 1;
    40: op1_11_inv23 = 1;
    43: op1_11_inv23 = 1;
    52: op1_11_inv23 = 1;
    53: op1_11_inv23 = 1;
    54: op1_11_inv23 = 1;
    57: op1_11_inv23 = 1;
    61: op1_11_inv23 = 1;
    63: op1_11_inv23 = 1;
    64: op1_11_inv23 = 1;
    65: op1_11_inv23 = 1;
    68: op1_11_inv23 = 1;
    69: op1_11_inv23 = 1;
    71: op1_11_inv23 = 1;
    75: op1_11_inv23 = 1;
    78: op1_11_inv23 = 1;
    81: op1_11_inv23 = 1;
    92: op1_11_inv23 = 1;
    93: op1_11_inv23 = 1;
    96: op1_11_inv23 = 1;
    default: op1_11_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in24 = imem04_in[23:20];
    6: op1_11_in24 = reg_0095;
    7: op1_11_in24 = imem06_in[27:24];
    9: op1_11_in24 = reg_0984;
    23: op1_11_in24 = reg_0984;
    10: op1_11_in24 = imem01_in[27:24];
    11: op1_11_in24 = reg_0952;
    12: op1_11_in24 = imem01_in[39:36];
    13: op1_11_in24 = imem06_in[3:0];
    15: op1_11_in24 = imem01_in[35:32];
    16: op1_11_in24 = reg_0555;
    17: op1_11_in24 = reg_0406;
    18: op1_11_in24 = reg_0306;
    19: op1_11_in24 = reg_0624;
    20: op1_11_in24 = reg_0740;
    21: op1_11_in24 = reg_0446;
    22: op1_11_in24 = reg_0636;
    24: op1_11_in24 = reg_0341;
    25: op1_11_in24 = reg_0733;
    26: op1_11_in24 = reg_0544;
    27: op1_11_in24 = imem06_in[127:124];
    28: op1_11_in24 = reg_0139;
    29: op1_11_in24 = reg_0586;
    30: op1_11_in24 = reg_0983;
    31: op1_11_in24 = reg_0424;
    32: op1_11_in24 = imem01_in[11:8];
    33: op1_11_in24 = reg_0810;
    34: op1_11_in24 = reg_0044;
    37: op1_11_in24 = reg_0104;
    39: op1_11_in24 = imem04_in[11:8];
    40: op1_11_in24 = reg_1020;
    41: op1_11_in24 = reg_0875;
    43: op1_11_in24 = reg_0829;
    44: op1_11_in24 = reg_0492;
    45: op1_11_in24 = reg_0716;
    47: op1_11_in24 = reg_0327;
    48: op1_11_in24 = imem07_in[127:124];
    50: op1_11_in24 = reg_0137;
    51: op1_11_in24 = imem05_in[51:48];
    52: op1_11_in24 = imem03_in[87:84];
    53: op1_11_in24 = reg_0864;
    54: op1_11_in24 = reg_0067;
    55: op1_11_in24 = reg_0718;
    58: op1_11_in24 = reg_0175;
    61: op1_11_in24 = reg_1056;
    62: op1_11_in24 = reg_0543;
    63: op1_11_in24 = reg_0692;
    64: op1_11_in24 = imem06_in[99:96];
    65: op1_11_in24 = reg_0719;
    67: op1_11_in24 = reg_0726;
    68: op1_11_in24 = reg_0608;
    69: op1_11_in24 = reg_0808;
    71: op1_11_in24 = reg_0521;
    72: op1_11_in24 = reg_0351;
    75: op1_11_in24 = reg_0488;
    76: op1_11_in24 = imem03_in[115:112];
    77: op1_11_in24 = imem05_in[71:68];
    78: op1_11_in24 = reg_0956;
    79: op1_11_in24 = reg_0338;
    81: op1_11_in24 = reg_1032;
    83: op1_11_in24 = imem05_in[119:116];
    84: op1_11_in24 = reg_0088;
    86: op1_11_in24 = reg_0198;
    87: op1_11_in24 = reg_0241;
    88: op1_11_in24 = reg_0181;
    89: op1_11_in24 = reg_0444;
    90: op1_11_in24 = imem07_in[35:32];
    91: op1_11_in24 = reg_0722;
    92: op1_11_in24 = reg_1022;
    93: op1_11_in24 = reg_0408;
    94: op1_11_in24 = reg_0788;
    95: op1_11_in24 = imem03_in[119:116];
    96: op1_11_in24 = reg_0049;
    default: op1_11_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv24 = 1;
    9: op1_11_inv24 = 1;
    10: op1_11_inv24 = 1;
    12: op1_11_inv24 = 1;
    15: op1_11_inv24 = 1;
    16: op1_11_inv24 = 1;
    17: op1_11_inv24 = 1;
    18: op1_11_inv24 = 1;
    23: op1_11_inv24 = 1;
    26: op1_11_inv24 = 1;
    28: op1_11_inv24 = 1;
    31: op1_11_inv24 = 1;
    34: op1_11_inv24 = 1;
    37: op1_11_inv24 = 1;
    41: op1_11_inv24 = 1;
    43: op1_11_inv24 = 1;
    44: op1_11_inv24 = 1;
    45: op1_11_inv24 = 1;
    47: op1_11_inv24 = 1;
    50: op1_11_inv24 = 1;
    52: op1_11_inv24 = 1;
    53: op1_11_inv24 = 1;
    54: op1_11_inv24 = 1;
    62: op1_11_inv24 = 1;
    65: op1_11_inv24 = 1;
    69: op1_11_inv24 = 1;
    75: op1_11_inv24 = 1;
    78: op1_11_inv24 = 1;
    81: op1_11_inv24 = 1;
    83: op1_11_inv24 = 1;
    84: op1_11_inv24 = 1;
    86: op1_11_inv24 = 1;
    87: op1_11_inv24 = 1;
    93: op1_11_inv24 = 1;
    95: op1_11_inv24 = 1;
    default: op1_11_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in25 = reg_0543;
    6: op1_11_in25 = reg_0090;
    7: op1_11_in25 = imem06_in[39:36];
    9: op1_11_in25 = reg_0996;
    10: op1_11_in25 = imem01_in[35:32];
    11: op1_11_in25 = reg_0268;
    12: op1_11_in25 = imem01_in[47:44];
    13: op1_11_in25 = imem06_in[43:40];
    15: op1_11_in25 = imem01_in[43:40];
    16: op1_11_in25 = reg_0551;
    17: op1_11_in25 = reg_0367;
    18: op1_11_in25 = reg_0302;
    19: op1_11_in25 = reg_0613;
    20: op1_11_in25 = reg_0062;
    25: op1_11_in25 = reg_0062;
    21: op1_11_in25 = reg_0438;
    22: op1_11_in25 = reg_0352;
    23: op1_11_in25 = reg_0990;
    24: op1_11_in25 = reg_0329;
    26: op1_11_in25 = reg_0905;
    27: op1_11_in25 = reg_0610;
    28: op1_11_in25 = reg_0129;
    29: op1_11_in25 = reg_0579;
    30: op1_11_in25 = reg_0994;
    31: op1_11_in25 = reg_0421;
    32: op1_11_in25 = imem01_in[51:48];
    33: op1_11_in25 = reg_0885;
    34: op1_11_in25 = imem05_in[23:20];
    53: op1_11_in25 = imem05_in[23:20];
    37: op1_11_in25 = reg_0119;
    39: op1_11_in25 = imem04_in[19:16];
    40: op1_11_in25 = reg_0292;
    41: op1_11_in25 = reg_0774;
    43: op1_11_in25 = reg_0925;
    44: op1_11_in25 = reg_1049;
    45: op1_11_in25 = reg_0719;
    47: op1_11_in25 = reg_0046;
    48: op1_11_in25 = reg_0723;
    50: op1_11_in25 = reg_0131;
    51: op1_11_in25 = imem05_in[103:100];
    52: op1_11_in25 = imem03_in[119:116];
    54: op1_11_in25 = reg_0078;
    55: op1_11_in25 = reg_0701;
    58: op1_11_in25 = reg_0161;
    61: op1_11_in25 = reg_1052;
    62: op1_11_in25 = reg_0370;
    63: op1_11_in25 = reg_0439;
    64: op1_11_in25 = imem06_in[127:124];
    65: op1_11_in25 = reg_0730;
    67: op1_11_in25 = reg_0717;
    68: op1_11_in25 = reg_0758;
    69: op1_11_in25 = reg_0288;
    71: op1_11_in25 = reg_0304;
    72: op1_11_in25 = reg_0262;
    75: op1_11_in25 = reg_0793;
    76: op1_11_in25 = imem03_in[123:120];
    95: op1_11_in25 = imem03_in[123:120];
    77: op1_11_in25 = reg_0866;
    78: op1_11_in25 = reg_0274;
    79: op1_11_in25 = reg_0735;
    81: op1_11_in25 = reg_0337;
    83: op1_11_in25 = imem05_in[127:124];
    84: op1_11_in25 = reg_0814;
    86: op1_11_in25 = reg_0196;
    87: op1_11_in25 = reg_0711;
    88: op1_11_in25 = reg_0157;
    89: op1_11_in25 = reg_0494;
    90: op1_11_in25 = imem07_in[43:40];
    91: op1_11_in25 = reg_0567;
    92: op1_11_in25 = reg_0604;
    93: op1_11_in25 = reg_0082;
    94: op1_11_in25 = imem03_in[43:40];
    96: op1_11_in25 = reg_0033;
    default: op1_11_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_11_inv25 = 1;
    9: op1_11_inv25 = 1;
    11: op1_11_inv25 = 1;
    12: op1_11_inv25 = 1;
    16: op1_11_inv25 = 1;
    17: op1_11_inv25 = 1;
    18: op1_11_inv25 = 1;
    20: op1_11_inv25 = 1;
    22: op1_11_inv25 = 1;
    23: op1_11_inv25 = 1;
    24: op1_11_inv25 = 1;
    29: op1_11_inv25 = 1;
    30: op1_11_inv25 = 1;
    31: op1_11_inv25 = 1;
    32: op1_11_inv25 = 1;
    37: op1_11_inv25 = 1;
    39: op1_11_inv25 = 1;
    40: op1_11_inv25 = 1;
    41: op1_11_inv25 = 1;
    51: op1_11_inv25 = 1;
    52: op1_11_inv25 = 1;
    54: op1_11_inv25 = 1;
    58: op1_11_inv25 = 1;
    65: op1_11_inv25 = 1;
    84: op1_11_inv25 = 1;
    87: op1_11_inv25 = 1;
    88: op1_11_inv25 = 1;
    89: op1_11_inv25 = 1;
    91: op1_11_inv25 = 1;
    93: op1_11_inv25 = 1;
    94: op1_11_inv25 = 1;
    default: op1_11_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in26 = reg_0545;
    6: op1_11_in26 = reg_0051;
    7: op1_11_in26 = imem06_in[55:52];
    9: op1_11_in26 = reg_0976;
    10: op1_11_in26 = imem01_in[87:84];
    11: op1_11_in26 = reg_0271;
    12: op1_11_in26 = imem01_in[67:64];
    13: op1_11_in26 = imem06_in[51:48];
    15: op1_11_in26 = imem01_in[51:48];
    16: op1_11_in26 = reg_0559;
    17: op1_11_in26 = reg_0401;
    18: op1_11_in26 = reg_0307;
    19: op1_11_in26 = reg_0633;
    20: op1_11_in26 = reg_0268;
    21: op1_11_in26 = reg_0181;
    22: op1_11_in26 = reg_0358;
    23: op1_11_in26 = imem04_in[11:8];
    24: op1_11_in26 = reg_0339;
    25: op1_11_in26 = reg_0076;
    26: op1_11_in26 = reg_1039;
    75: op1_11_in26 = reg_1039;
    27: op1_11_in26 = reg_0620;
    28: op1_11_in26 = reg_0153;
    29: op1_11_in26 = reg_0583;
    30: op1_11_in26 = imem04_in[51:48];
    31: op1_11_in26 = reg_0447;
    32: op1_11_in26 = imem01_in[59:56];
    33: op1_11_in26 = reg_1043;
    34: op1_11_in26 = reg_0971;
    37: op1_11_in26 = reg_0114;
    39: op1_11_in26 = imem04_in[47:44];
    40: op1_11_in26 = reg_0050;
    41: op1_11_in26 = reg_0864;
    43: op1_11_in26 = reg_0615;
    44: op1_11_in26 = reg_0397;
    45: op1_11_in26 = reg_0730;
    47: op1_11_in26 = reg_0396;
    48: op1_11_in26 = reg_0702;
    50: op1_11_in26 = reg_0134;
    87: op1_11_in26 = reg_0134;
    51: op1_11_in26 = reg_0973;
    52: op1_11_in26 = reg_0571;
    53: op1_11_in26 = imem05_in[55:52];
    54: op1_11_in26 = reg_0816;
    55: op1_11_in26 = reg_0700;
    58: op1_11_in26 = reg_0162;
    61: op1_11_in26 = reg_0238;
    62: op1_11_in26 = reg_0311;
    63: op1_11_in26 = reg_0804;
    64: op1_11_in26 = reg_0660;
    65: op1_11_in26 = reg_0726;
    67: op1_11_in26 = reg_0712;
    91: op1_11_in26 = reg_0712;
    68: op1_11_in26 = reg_0876;
    69: op1_11_in26 = reg_0432;
    71: op1_11_in26 = reg_0733;
    72: op1_11_in26 = reg_0817;
    76: op1_11_in26 = reg_0228;
    77: op1_11_in26 = reg_0057;
    78: op1_11_in26 = reg_0237;
    79: op1_11_in26 = reg_0533;
    81: op1_11_in26 = reg_0488;
    83: op1_11_in26 = reg_0319;
    84: op1_11_in26 = reg_0049;
    86: op1_11_in26 = reg_0212;
    89: op1_11_in26 = reg_0517;
    90: op1_11_in26 = imem07_in[83:80];
    92: op1_11_in26 = reg_1037;
    93: op1_11_in26 = reg_0367;
    94: op1_11_in26 = imem03_in[71:68];
    95: op1_11_in26 = reg_0819;
    96: op1_11_in26 = reg_0342;
    default: op1_11_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv26 = 1;
    9: op1_11_inv26 = 1;
    10: op1_11_inv26 = 1;
    12: op1_11_inv26 = 1;
    13: op1_11_inv26 = 1;
    15: op1_11_inv26 = 1;
    18: op1_11_inv26 = 1;
    20: op1_11_inv26 = 1;
    21: op1_11_inv26 = 1;
    23: op1_11_inv26 = 1;
    24: op1_11_inv26 = 1;
    26: op1_11_inv26 = 1;
    27: op1_11_inv26 = 1;
    28: op1_11_inv26 = 1;
    37: op1_11_inv26 = 1;
    40: op1_11_inv26 = 1;
    41: op1_11_inv26 = 1;
    43: op1_11_inv26 = 1;
    48: op1_11_inv26 = 1;
    53: op1_11_inv26 = 1;
    55: op1_11_inv26 = 1;
    58: op1_11_inv26 = 1;
    61: op1_11_inv26 = 1;
    63: op1_11_inv26 = 1;
    65: op1_11_inv26 = 1;
    67: op1_11_inv26 = 1;
    68: op1_11_inv26 = 1;
    76: op1_11_inv26 = 1;
    78: op1_11_inv26 = 1;
    79: op1_11_inv26 = 1;
    83: op1_11_inv26 = 1;
    86: op1_11_inv26 = 1;
    89: op1_11_inv26 = 1;
    90: op1_11_inv26 = 1;
    91: op1_11_inv26 = 1;
    93: op1_11_inv26 = 1;
    96: op1_11_inv26 = 1;
    default: op1_11_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in27 = reg_0550;
    6: op1_11_in27 = reg_0055;
    7: op1_11_in27 = imem06_in[71:68];
    9: op1_11_in27 = reg_0994;
    10: op1_11_in27 = imem01_in[119:116];
    11: op1_11_in27 = reg_0260;
    12: op1_11_in27 = reg_1051;
    13: op1_11_in27 = imem06_in[95:92];
    15: op1_11_in27 = imem01_in[71:68];
    16: op1_11_in27 = reg_0308;
    17: op1_11_in27 = reg_0799;
    18: op1_11_in27 = imem04_in[55:52];
    30: op1_11_in27 = imem04_in[55:52];
    19: op1_11_in27 = reg_0608;
    20: op1_11_in27 = reg_0259;
    21: op1_11_in27 = reg_0166;
    22: op1_11_in27 = reg_0354;
    23: op1_11_in27 = imem04_in[19:16];
    24: op1_11_in27 = reg_0346;
    25: op1_11_in27 = reg_0064;
    26: op1_11_in27 = reg_1043;
    27: op1_11_in27 = reg_0402;
    28: op1_11_in27 = reg_0140;
    29: op1_11_in27 = reg_0587;
    31: op1_11_in27 = reg_0419;
    32: op1_11_in27 = imem01_in[127:124];
    33: op1_11_in27 = reg_1044;
    34: op1_11_in27 = reg_0957;
    37: op1_11_in27 = reg_0100;
    39: op1_11_in27 = imem04_in[63:60];
    40: op1_11_in27 = reg_0313;
    41: op1_11_in27 = imem05_in[11:8];
    43: op1_11_in27 = reg_0124;
    44: op1_11_in27 = reg_0581;
    45: op1_11_in27 = reg_0721;
    47: op1_11_in27 = reg_0004;
    48: op1_11_in27 = reg_0724;
    50: op1_11_in27 = reg_0144;
    51: op1_11_in27 = reg_0944;
    52: op1_11_in27 = reg_1019;
    53: op1_11_in27 = imem05_in[67:64];
    54: op1_11_in27 = reg_0528;
    55: op1_11_in27 = reg_0250;
    58: op1_11_in27 = reg_0182;
    61: op1_11_in27 = reg_0285;
    62: op1_11_in27 = reg_0509;
    63: op1_11_in27 = reg_0632;
    64: op1_11_in27 = reg_0625;
    65: op1_11_in27 = reg_0717;
    67: op1_11_in27 = reg_0705;
    68: op1_11_in27 = reg_0049;
    69: op1_11_in27 = reg_0407;
    71: op1_11_in27 = reg_0653;
    72: op1_11_in27 = reg_0297;
    75: op1_11_in27 = reg_0501;
    76: op1_11_in27 = reg_0572;
    77: op1_11_in27 = reg_0583;
    78: op1_11_in27 = reg_0438;
    79: op1_11_in27 = reg_0804;
    81: op1_11_in27 = reg_0234;
    83: op1_11_in27 = reg_0647;
    84: op1_11_in27 = reg_0840;
    86: op1_11_in27 = reg_0190;
    87: op1_11_in27 = reg_0489;
    89: op1_11_in27 = reg_0070;
    90: op1_11_in27 = imem07_in[127:124];
    91: op1_11_in27 = reg_0710;
    92: op1_11_in27 = reg_1041;
    93: op1_11_in27 = imem03_in[7:4];
    94: op1_11_in27 = imem03_in[91:88];
    95: op1_11_in27 = reg_0859;
    96: op1_11_in27 = reg_0623;
    default: op1_11_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv27 = 1;
    6: op1_11_inv27 = 1;
    9: op1_11_inv27 = 1;
    10: op1_11_inv27 = 1;
    11: op1_11_inv27 = 1;
    12: op1_11_inv27 = 1;
    13: op1_11_inv27 = 1;
    15: op1_11_inv27 = 1;
    17: op1_11_inv27 = 1;
    18: op1_11_inv27 = 1;
    19: op1_11_inv27 = 1;
    21: op1_11_inv27 = 1;
    24: op1_11_inv27 = 1;
    25: op1_11_inv27 = 1;
    26: op1_11_inv27 = 1;
    27: op1_11_inv27 = 1;
    29: op1_11_inv27 = 1;
    30: op1_11_inv27 = 1;
    31: op1_11_inv27 = 1;
    32: op1_11_inv27 = 1;
    33: op1_11_inv27 = 1;
    40: op1_11_inv27 = 1;
    44: op1_11_inv27 = 1;
    45: op1_11_inv27 = 1;
    47: op1_11_inv27 = 1;
    48: op1_11_inv27 = 1;
    53: op1_11_inv27 = 1;
    55: op1_11_inv27 = 1;
    61: op1_11_inv27 = 1;
    65: op1_11_inv27 = 1;
    67: op1_11_inv27 = 1;
    68: op1_11_inv27 = 1;
    69: op1_11_inv27 = 1;
    71: op1_11_inv27 = 1;
    72: op1_11_inv27 = 1;
    75: op1_11_inv27 = 1;
    76: op1_11_inv27 = 1;
    77: op1_11_inv27 = 1;
    81: op1_11_inv27 = 1;
    83: op1_11_inv27 = 1;
    87: op1_11_inv27 = 1;
    90: op1_11_inv27 = 1;
    93: op1_11_inv27 = 1;
    94: op1_11_inv27 = 1;
    default: op1_11_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in28 = reg_0529;
    6: op1_11_in28 = reg_0823;
    7: op1_11_in28 = imem06_in[75:72];
    9: op1_11_in28 = imem04_in[7:4];
    10: op1_11_in28 = reg_0118;
    11: op1_11_in28 = reg_0265;
    12: op1_11_in28 = reg_0762;
    13: op1_11_in28 = imem06_in[103:100];
    15: op1_11_in28 = imem01_in[91:88];
    16: op1_11_in28 = reg_0283;
    17: op1_11_in28 = reg_0027;
    54: op1_11_in28 = reg_0027;
    18: op1_11_in28 = imem04_in[67:64];
    19: op1_11_in28 = reg_0623;
    20: op1_11_in28 = reg_0755;
    22: op1_11_in28 = reg_0359;
    23: op1_11_in28 = imem04_in[27:24];
    24: op1_11_in28 = reg_0336;
    25: op1_11_in28 = reg_0738;
    26: op1_11_in28 = reg_0500;
    27: op1_11_in28 = reg_0386;
    28: op1_11_in28 = imem06_in[39:36];
    29: op1_11_in28 = reg_0593;
    30: op1_11_in28 = imem04_in[79:76];
    31: op1_11_in28 = reg_0420;
    32: op1_11_in28 = reg_0236;
    33: op1_11_in28 = reg_1034;
    34: op1_11_in28 = reg_0953;
    37: op1_11_in28 = reg_0109;
    39: op1_11_in28 = imem04_in[95:92];
    40: op1_11_in28 = reg_0268;
    41: op1_11_in28 = imem05_in[23:20];
    43: op1_11_in28 = reg_0112;
    44: op1_11_in28 = reg_0923;
    45: op1_11_in28 = reg_0723;
    47: op1_11_in28 = reg_0389;
    48: op1_11_in28 = reg_0718;
    67: op1_11_in28 = reg_0718;
    50: op1_11_in28 = imem06_in[15:12];
    51: op1_11_in28 = reg_0959;
    52: op1_11_in28 = reg_0398;
    53: op1_11_in28 = imem05_in[95:92];
    55: op1_11_in28 = reg_0421;
    58: op1_11_in28 = reg_0183;
    61: op1_11_in28 = reg_0501;
    62: op1_11_in28 = reg_0836;
    63: op1_11_in28 = reg_0348;
    64: op1_11_in28 = reg_0626;
    65: op1_11_in28 = reg_0711;
    68: op1_11_in28 = reg_0840;
    69: op1_11_in28 = reg_0065;
    71: op1_11_in28 = reg_0899;
    72: op1_11_in28 = reg_0895;
    75: op1_11_in28 = reg_0522;
    76: op1_11_in28 = reg_0445;
    77: op1_11_in28 = reg_0935;
    78: op1_11_in28 = reg_0707;
    79: op1_11_in28 = reg_0632;
    81: op1_11_in28 = reg_0496;
    83: op1_11_in28 = reg_0143;
    84: op1_11_in28 = reg_0291;
    86: op1_11_in28 = imem01_in[7:4];
    87: op1_11_in28 = reg_0215;
    89: op1_11_in28 = imem05_in[7:4];
    90: op1_11_in28 = reg_0567;
    91: op1_11_in28 = reg_0361;
    92: op1_11_in28 = reg_0769;
    93: op1_11_in28 = imem03_in[23:20];
    94: op1_11_in28 = imem03_in[123:120];
    95: op1_11_in28 = reg_0620;
    96: op1_11_in28 = reg_0238;
    default: op1_11_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv28 = 1;
    9: op1_11_inv28 = 1;
    11: op1_11_inv28 = 1;
    12: op1_11_inv28 = 1;
    13: op1_11_inv28 = 1;
    15: op1_11_inv28 = 1;
    16: op1_11_inv28 = 1;
    18: op1_11_inv28 = 1;
    25: op1_11_inv28 = 1;
    26: op1_11_inv28 = 1;
    27: op1_11_inv28 = 1;
    28: op1_11_inv28 = 1;
    30: op1_11_inv28 = 1;
    31: op1_11_inv28 = 1;
    33: op1_11_inv28 = 1;
    39: op1_11_inv28 = 1;
    43: op1_11_inv28 = 1;
    45: op1_11_inv28 = 1;
    47: op1_11_inv28 = 1;
    48: op1_11_inv28 = 1;
    50: op1_11_inv28 = 1;
    51: op1_11_inv28 = 1;
    52: op1_11_inv28 = 1;
    54: op1_11_inv28 = 1;
    55: op1_11_inv28 = 1;
    58: op1_11_inv28 = 1;
    61: op1_11_inv28 = 1;
    63: op1_11_inv28 = 1;
    65: op1_11_inv28 = 1;
    68: op1_11_inv28 = 1;
    69: op1_11_inv28 = 1;
    71: op1_11_inv28 = 1;
    72: op1_11_inv28 = 1;
    77: op1_11_inv28 = 1;
    81: op1_11_inv28 = 1;
    83: op1_11_inv28 = 1;
    84: op1_11_inv28 = 1;
    86: op1_11_inv28 = 1;
    87: op1_11_inv28 = 1;
    89: op1_11_inv28 = 1;
    91: op1_11_inv28 = 1;
    95: op1_11_inv28 = 1;
    default: op1_11_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in29 = reg_0539;
    6: op1_11_in29 = reg_0817;
    7: op1_11_in29 = imem06_in[91:88];
    9: op1_11_in29 = imem04_in[47:44];
    10: op1_11_in29 = reg_0120;
    11: op1_11_in29 = reg_0272;
    12: op1_11_in29 = reg_0220;
    13: op1_11_in29 = reg_0629;
    15: op1_11_in29 = imem01_in[99:96];
    16: op1_11_in29 = reg_0289;
    17: op1_11_in29 = reg_0801;
    18: op1_11_in29 = imem04_in[95:92];
    19: op1_11_in29 = reg_0402;
    20: op1_11_in29 = reg_0068;
    22: op1_11_in29 = reg_0329;
    23: op1_11_in29 = imem04_in[59:56];
    24: op1_11_in29 = reg_0007;
    25: op1_11_in29 = reg_0854;
    26: op1_11_in29 = reg_0216;
    27: op1_11_in29 = reg_0399;
    28: op1_11_in29 = imem06_in[55:52];
    29: op1_11_in29 = reg_0597;
    30: op1_11_in29 = imem04_in[87:84];
    31: op1_11_in29 = reg_0175;
    32: op1_11_in29 = reg_0544;
    33: op1_11_in29 = reg_0122;
    34: op1_11_in29 = reg_0960;
    37: op1_11_in29 = imem02_in[11:8];
    39: op1_11_in29 = imem04_in[115:112];
    40: op1_11_in29 = reg_0076;
    41: op1_11_in29 = imem05_in[35:32];
    89: op1_11_in29 = imem05_in[35:32];
    43: op1_11_in29 = reg_0102;
    44: op1_11_in29 = reg_0369;
    45: op1_11_in29 = reg_0714;
    47: op1_11_in29 = reg_0793;
    48: op1_11_in29 = reg_0700;
    50: op1_11_in29 = imem06_in[27:24];
    51: op1_11_in29 = reg_0954;
    52: op1_11_in29 = reg_0396;
    53: op1_11_in29 = imem05_in[115:112];
    54: op1_11_in29 = reg_0529;
    55: op1_11_in29 = reg_0426;
    58: op1_11_in29 = reg_0170;
    61: op1_11_in29 = reg_0829;
    81: op1_11_in29 = reg_0829;
    62: op1_11_in29 = reg_0985;
    63: op1_11_in29 = reg_0241;
    64: op1_11_in29 = reg_0754;
    65: op1_11_in29 = reg_0707;
    77: op1_11_in29 = reg_0707;
    67: op1_11_in29 = reg_0711;
    68: op1_11_in29 = reg_0310;
    69: op1_11_in29 = reg_0027;
    71: op1_11_in29 = reg_0914;
    72: op1_11_in29 = reg_0395;
    75: op1_11_in29 = reg_1043;
    76: op1_11_in29 = reg_0307;
    78: op1_11_in29 = reg_0780;
    79: op1_11_in29 = reg_0222;
    83: op1_11_in29 = reg_0138;
    84: op1_11_in29 = reg_0884;
    86: op1_11_in29 = imem01_in[11:8];
    87: op1_11_in29 = reg_0217;
    90: op1_11_in29 = reg_0165;
    91: op1_11_in29 = reg_0303;
    92: op1_11_in29 = reg_0283;
    93: op1_11_in29 = imem03_in[27:24];
    94: op1_11_in29 = reg_0758;
    95: op1_11_in29 = reg_0301;
    96: op1_11_in29 = reg_0385;
    default: op1_11_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_11_inv29 = 1;
    11: op1_11_inv29 = 1;
    12: op1_11_inv29 = 1;
    16: op1_11_inv29 = 1;
    17: op1_11_inv29 = 1;
    19: op1_11_inv29 = 1;
    22: op1_11_inv29 = 1;
    24: op1_11_inv29 = 1;
    25: op1_11_inv29 = 1;
    32: op1_11_inv29 = 1;
    33: op1_11_inv29 = 1;
    34: op1_11_inv29 = 1;
    37: op1_11_inv29 = 1;
    41: op1_11_inv29 = 1;
    43: op1_11_inv29 = 1;
    44: op1_11_inv29 = 1;
    45: op1_11_inv29 = 1;
    51: op1_11_inv29 = 1;
    52: op1_11_inv29 = 1;
    53: op1_11_inv29 = 1;
    55: op1_11_inv29 = 1;
    58: op1_11_inv29 = 1;
    61: op1_11_inv29 = 1;
    62: op1_11_inv29 = 1;
    64: op1_11_inv29 = 1;
    65: op1_11_inv29 = 1;
    71: op1_11_inv29 = 1;
    75: op1_11_inv29 = 1;
    77: op1_11_inv29 = 1;
    81: op1_11_inv29 = 1;
    83: op1_11_inv29 = 1;
    84: op1_11_inv29 = 1;
    87: op1_11_inv29 = 1;
    91: op1_11_inv29 = 1;
    93: op1_11_inv29 = 1;
    94: op1_11_inv29 = 1;
    95: op1_11_inv29 = 1;
    96: op1_11_inv29 = 1;
    default: op1_11_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_11_in30 = reg_0548;
    6: op1_11_in30 = reg_0820;
    7: op1_11_in30 = imem06_in[99:96];
    9: op1_11_in30 = imem04_in[63:60];
    10: op1_11_in30 = reg_0121;
    11: op1_11_in30 = reg_0261;
    12: op1_11_in30 = reg_0247;
    13: op1_11_in30 = reg_0607;
    15: op1_11_in30 = imem01_in[119:116];
    16: op1_11_in30 = reg_0285;
    17: op1_11_in30 = reg_0754;
    18: op1_11_in30 = imem05_in[11:8];
    19: op1_11_in30 = reg_0381;
    20: op1_11_in30 = reg_0296;
    22: op1_11_in30 = reg_0342;
    23: op1_11_in30 = imem04_in[67:64];
    24: op1_11_in30 = reg_0758;
    25: op1_11_in30 = reg_0774;
    26: op1_11_in30 = reg_1040;
    27: op1_11_in30 = reg_0404;
    28: op1_11_in30 = reg_0628;
    29: op1_11_in30 = reg_0581;
    30: op1_11_in30 = imem04_in[91:88];
    31: op1_11_in30 = reg_0181;
    32: op1_11_in30 = reg_0905;
    33: op1_11_in30 = reg_0118;
    34: op1_11_in30 = reg_1021;
    37: op1_11_in30 = imem02_in[15:12];
    39: op1_11_in30 = imem04_in[119:116];
    40: op1_11_in30 = reg_0014;
    41: op1_11_in30 = imem05_in[43:40];
    43: op1_11_in30 = reg_0114;
    44: op1_11_in30 = reg_0807;
    45: op1_11_in30 = reg_0703;
    47: op1_11_in30 = reg_0795;
    48: op1_11_in30 = reg_0169;
    50: op1_11_in30 = imem06_in[35:32];
    51: op1_11_in30 = reg_0957;
    52: op1_11_in30 = reg_0004;
    53: op1_11_in30 = reg_0966;
    54: op1_11_in30 = reg_0041;
    55: op1_11_in30 = reg_0321;
    58: op1_11_in30 = reg_0158;
    61: op1_11_in30 = reg_0514;
    75: op1_11_in30 = reg_0514;
    81: op1_11_in30 = reg_0514;
    62: op1_11_in30 = reg_0998;
    63: op1_11_in30 = reg_1028;
    64: op1_11_in30 = reg_0692;
    65: op1_11_in30 = reg_0303;
    67: op1_11_in30 = reg_0706;
    68: op1_11_in30 = reg_0884;
    69: op1_11_in30 = reg_0854;
    71: op1_11_in30 = reg_0647;
    72: op1_11_in30 = reg_0617;
    76: op1_11_in30 = reg_0322;
    77: op1_11_in30 = reg_0508;
    78: op1_11_in30 = reg_0806;
    79: op1_11_in30 = reg_0921;
    83: op1_11_in30 = reg_0275;
    84: op1_11_in30 = imem03_in[11:8];
    86: op1_11_in30 = imem01_in[19:16];
    87: op1_11_in30 = reg_0954;
    89: op1_11_in30 = imem05_in[107:104];
    90: op1_11_in30 = reg_0159;
    91: op1_11_in30 = reg_0325;
    92: op1_11_in30 = reg_0860;
    93: op1_11_in30 = imem03_in[31:28];
    94: op1_11_in30 = reg_1050;
    95: op1_11_in30 = reg_0976;
    96: op1_11_in30 = reg_0588;
    default: op1_11_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv30 = 1;
    6: op1_11_inv30 = 1;
    7: op1_11_inv30 = 1;
    10: op1_11_inv30 = 1;
    16: op1_11_inv30 = 1;
    18: op1_11_inv30 = 1;
    20: op1_11_inv30 = 1;
    23: op1_11_inv30 = 1;
    24: op1_11_inv30 = 1;
    28: op1_11_inv30 = 1;
    29: op1_11_inv30 = 1;
    32: op1_11_inv30 = 1;
    37: op1_11_inv30 = 1;
    39: op1_11_inv30 = 1;
    40: op1_11_inv30 = 1;
    44: op1_11_inv30 = 1;
    47: op1_11_inv30 = 1;
    48: op1_11_inv30 = 1;
    50: op1_11_inv30 = 1;
    51: op1_11_inv30 = 1;
    53: op1_11_inv30 = 1;
    54: op1_11_inv30 = 1;
    58: op1_11_inv30 = 1;
    61: op1_11_inv30 = 1;
    62: op1_11_inv30 = 1;
    63: op1_11_inv30 = 1;
    65: op1_11_inv30 = 1;
    67: op1_11_inv30 = 1;
    69: op1_11_inv30 = 1;
    72: op1_11_inv30 = 1;
    75: op1_11_inv30 = 1;
    76: op1_11_inv30 = 1;
    77: op1_11_inv30 = 1;
    78: op1_11_inv30 = 1;
    83: op1_11_inv30 = 1;
    89: op1_11_inv30 = 1;
    96: op1_11_inv30 = 1;
    default: op1_11_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_11_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_11_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in00 = reg_0531;
    6: op1_12_in00 = reg_0833;
    7: op1_12_in00 = imem06_in[111:108];
    8: op1_12_in00 = imem00_in[67:64];
    9: op1_12_in00 = imem04_in[71:68];
    10: op1_12_in00 = reg_0110;
    11: op1_12_in00 = reg_0142;
    12: op1_12_in00 = reg_0248;
    13: op1_12_in00 = reg_0613;
    14: op1_12_in00 = imem00_in[7:4];
    21: op1_12_in00 = imem00_in[7:4];
    35: op1_12_in00 = imem00_in[7:4];
    36: op1_12_in00 = imem00_in[7:4];
    57: op1_12_in00 = imem00_in[7:4];
    66: op1_12_in00 = imem00_in[7:4];
    15: op1_12_in00 = reg_0233;
    16: op1_12_in00 = reg_0307;
    17: op1_12_in00 = reg_0798;
    18: op1_12_in00 = imem05_in[67:64];
    19: op1_12_in00 = reg_0371;
    20: op1_12_in00 = reg_0064;
    22: op1_12_in00 = reg_0355;
    23: op1_12_in00 = imem04_in[75:72];
    24: op1_12_in00 = reg_0016;
    25: op1_12_in00 = reg_0777;
    4: op1_12_in00 = imem07_in[19:16];
    26: op1_12_in00 = reg_0871;
    3: op1_12_in00 = imem07_in[11:8];
    27: op1_12_in00 = reg_0486;
    28: op1_12_in00 = reg_0604;
    29: op1_12_in00 = reg_0543;
    30: op1_12_in00 = imem04_in[119:116];
    31: op1_12_in00 = imem00_in[11:8];
    38: op1_12_in00 = imem00_in[11:8];
    74: op1_12_in00 = imem00_in[11:8];
    2: op1_12_in00 = imem07_in[39:36];
    32: op1_12_in00 = reg_1042;
    33: op1_12_in00 = reg_0120;
    34: op1_12_in00 = reg_0835;
    37: op1_12_in00 = imem02_in[23:20];
    39: op1_12_in00 = reg_0937;
    40: op1_12_in00 = reg_0009;
    41: op1_12_in00 = imem05_in[51:48];
    42: op1_12_in00 = imem00_in[27:24];
    70: op1_12_in00 = imem00_in[27:24];
    43: op1_12_in00 = imem02_in[27:24];
    44: op1_12_in00 = reg_0836;
    45: op1_12_in00 = reg_0729;
    46: op1_12_in00 = imem00_in[31:28];
    47: op1_12_in00 = reg_0509;
    48: op1_12_in00 = reg_0173;
    49: op1_12_in00 = reg_0680;
    50: op1_12_in00 = imem06_in[55:52];
    51: op1_12_in00 = reg_0259;
    52: op1_12_in00 = reg_0824;
    53: op1_12_in00 = reg_0971;
    54: op1_12_in00 = reg_0764;
    55: op1_12_in00 = reg_0868;
    56: op1_12_in00 = imem00_in[59:56];
    58: op1_12_in00 = reg_0184;
    59: op1_12_in00 = imem00_in[23:20];
    60: op1_12_in00 = imem00_in[43:40];
    61: op1_12_in00 = reg_0354;
    81: op1_12_in00 = reg_0354;
    62: op1_12_in00 = reg_0993;
    63: op1_12_in00 = reg_0264;
    64: op1_12_in00 = reg_0614;
    65: op1_12_in00 = reg_0315;
    91: op1_12_in00 = reg_0315;
    67: op1_12_in00 = reg_0422;
    68: op1_12_in00 = imem03_in[11:8];
    69: op1_12_in00 = reg_0070;
    71: op1_12_in00 = reg_0636;
    72: op1_12_in00 = reg_0595;
    73: op1_12_in00 = imem00_in[15:12];
    88: op1_12_in00 = imem00_in[15:12];
    75: op1_12_in00 = reg_0216;
    76: op1_12_in00 = reg_0240;
    77: op1_12_in00 = reg_0706;
    78: op1_12_in00 = reg_0490;
    79: op1_12_in00 = reg_0026;
    80: op1_12_in00 = imem00_in[35:32];
    82: op1_12_in00 = imem00_in[3:0];
    83: op1_12_in00 = reg_0235;
    84: op1_12_in00 = imem03_in[59:56];
    85: op1_12_in00 = imem00_in[19:16];
    86: op1_12_in00 = imem01_in[67:64];
    87: op1_12_in00 = reg_0319;
    89: op1_12_in00 = imem05_in[111:108];
    90: op1_12_in00 = reg_0560;
    92: op1_12_in00 = reg_0821;
    93: op1_12_in00 = imem03_in[43:40];
    94: op1_12_in00 = reg_0761;
    95: op1_12_in00 = reg_0558;
    96: op1_12_in00 = reg_0523;
    default: op1_12_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv00 = 1;
    6: op1_12_inv00 = 1;
    7: op1_12_inv00 = 1;
    8: op1_12_inv00 = 1;
    10: op1_12_inv00 = 1;
    11: op1_12_inv00 = 1;
    15: op1_12_inv00 = 1;
    17: op1_12_inv00 = 1;
    20: op1_12_inv00 = 1;
    21: op1_12_inv00 = 1;
    22: op1_12_inv00 = 1;
    23: op1_12_inv00 = 1;
    25: op1_12_inv00 = 1;
    3: op1_12_inv00 = 1;
    28: op1_12_inv00 = 1;
    30: op1_12_inv00 = 1;
    2: op1_12_inv00 = 1;
    34: op1_12_inv00 = 1;
    36: op1_12_inv00 = 1;
    37: op1_12_inv00 = 1;
    38: op1_12_inv00 = 1;
    41: op1_12_inv00 = 1;
    43: op1_12_inv00 = 1;
    44: op1_12_inv00 = 1;
    45: op1_12_inv00 = 1;
    46: op1_12_inv00 = 1;
    47: op1_12_inv00 = 1;
    48: op1_12_inv00 = 1;
    52: op1_12_inv00 = 1;
    53: op1_12_inv00 = 1;
    56: op1_12_inv00 = 1;
    57: op1_12_inv00 = 1;
    59: op1_12_inv00 = 1;
    64: op1_12_inv00 = 1;
    67: op1_12_inv00 = 1;
    70: op1_12_inv00 = 1;
    72: op1_12_inv00 = 1;
    74: op1_12_inv00 = 1;
    75: op1_12_inv00 = 1;
    78: op1_12_inv00 = 1;
    79: op1_12_inv00 = 1;
    80: op1_12_inv00 = 1;
    81: op1_12_inv00 = 1;
    82: op1_12_inv00 = 1;
    83: op1_12_inv00 = 1;
    85: op1_12_inv00 = 1;
    86: op1_12_inv00 = 1;
    90: op1_12_inv00 = 1;
    94: op1_12_inv00 = 1;
    95: op1_12_inv00 = 1;
    default: op1_12_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in01 = reg_0303;
    6: op1_12_in01 = reg_0825;
    7: op1_12_in01 = reg_0631;
    8: op1_12_in01 = reg_0693;
    9: op1_12_in01 = imem04_in[75:72];
    10: op1_12_in01 = imem02_in[7:4];
    11: op1_12_in01 = reg_0131;
    12: op1_12_in01 = reg_0234;
    13: op1_12_in01 = reg_0620;
    28: op1_12_in01 = reg_0620;
    14: op1_12_in01 = imem00_in[11:8];
    15: op1_12_in01 = reg_1049;
    16: op1_12_in01 = reg_0059;
    40: op1_12_in01 = reg_0059;
    17: op1_12_in01 = imem07_in[7:4];
    18: op1_12_in01 = reg_0963;
    19: op1_12_in01 = reg_0375;
    20: op1_12_in01 = reg_0748;
    21: op1_12_in01 = imem00_in[59:56];
    36: op1_12_in01 = imem00_in[59:56];
    22: op1_12_in01 = reg_0347;
    23: op1_12_in01 = imem04_in[79:76];
    24: op1_12_in01 = imem03_in[3:0];
    25: op1_12_in01 = reg_0285;
    4: op1_12_in01 = imem07_in[47:44];
    26: op1_12_in01 = reg_1017;
    81: op1_12_in01 = reg_1017;
    3: op1_12_in01 = imem07_in[23:20];
    27: op1_12_in01 = reg_0753;
    29: op1_12_in01 = reg_0795;
    30: op1_12_in01 = reg_1004;
    31: op1_12_in01 = imem00_in[23:20];
    73: op1_12_in01 = imem00_in[23:20];
    2: op1_12_in01 = imem07_in[75:72];
    32: op1_12_in01 = reg_0885;
    33: op1_12_in01 = reg_0102;
    34: op1_12_in01 = reg_0256;
    35: op1_12_in01 = imem00_in[27:24];
    38: op1_12_in01 = imem00_in[27:24];
    37: op1_12_in01 = imem02_in[107:104];
    39: op1_12_in01 = reg_0540;
    41: op1_12_in01 = imem05_in[59:56];
    42: op1_12_in01 = imem00_in[39:36];
    66: op1_12_in01 = imem00_in[39:36];
    74: op1_12_in01 = imem00_in[39:36];
    85: op1_12_in01 = imem00_in[39:36];
    88: op1_12_in01 = imem00_in[39:36];
    43: op1_12_in01 = imem02_in[39:36];
    44: op1_12_in01 = reg_0844;
    45: op1_12_in01 = reg_0718;
    46: op1_12_in01 = imem00_in[35:32];
    47: op1_12_in01 = reg_0051;
    49: op1_12_in01 = reg_0688;
    50: op1_12_in01 = imem06_in[67:64];
    51: op1_12_in01 = reg_0032;
    52: op1_12_in01 = reg_0576;
    53: op1_12_in01 = reg_0954;
    54: op1_12_in01 = imem05_in[7:4];
    55: op1_12_in01 = reg_0640;
    56: op1_12_in01 = imem00_in[63:60];
    57: op1_12_in01 = imem00_in[55:52];
    59: op1_12_in01 = imem00_in[87:84];
    60: op1_12_in01 = imem00_in[67:64];
    61: op1_12_in01 = reg_0832;
    62: op1_12_in01 = reg_0981;
    63: op1_12_in01 = imem07_in[27:24];
    64: op1_12_in01 = reg_0395;
    65: op1_12_in01 = reg_0641;
    67: op1_12_in01 = reg_0024;
    68: op1_12_in01 = imem03_in[15:12];
    69: op1_12_in01 = imem05_in[19:16];
    70: op1_12_in01 = imem00_in[51:48];
    71: op1_12_in01 = reg_0394;
    72: op1_12_in01 = reg_0556;
    75: op1_12_in01 = reg_1040;
    76: op1_12_in01 = reg_0662;
    77: op1_12_in01 = reg_0252;
    78: op1_12_in01 = imem06_in[51:48];
    79: op1_12_in01 = reg_0834;
    80: op1_12_in01 = imem00_in[71:68];
    82: op1_12_in01 = imem00_in[7:4];
    83: op1_12_in01 = reg_0448;
    84: op1_12_in01 = reg_0535;
    86: op1_12_in01 = imem01_in[87:84];
    87: op1_12_in01 = reg_0138;
    89: op1_12_in01 = imem05_in[127:124];
    90: op1_12_in01 = reg_0250;
    91: op1_12_in01 = reg_0353;
    92: op1_12_in01 = imem02_in[19:16];
    93: op1_12_in01 = imem03_in[59:56];
    94: op1_12_in01 = reg_0743;
    95: op1_12_in01 = reg_0756;
    96: op1_12_in01 = reg_0975;
    default: op1_12_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv01 = 1;
    6: op1_12_inv01 = 1;
    7: op1_12_inv01 = 1;
    8: op1_12_inv01 = 1;
    11: op1_12_inv01 = 1;
    12: op1_12_inv01 = 1;
    14: op1_12_inv01 = 1;
    15: op1_12_inv01 = 1;
    17: op1_12_inv01 = 1;
    18: op1_12_inv01 = 1;
    19: op1_12_inv01 = 1;
    20: op1_12_inv01 = 1;
    23: op1_12_inv01 = 1;
    25: op1_12_inv01 = 1;
    26: op1_12_inv01 = 1;
    3: op1_12_inv01 = 1;
    27: op1_12_inv01 = 1;
    28: op1_12_inv01 = 1;
    30: op1_12_inv01 = 1;
    31: op1_12_inv01 = 1;
    34: op1_12_inv01 = 1;
    39: op1_12_inv01 = 1;
    41: op1_12_inv01 = 1;
    42: op1_12_inv01 = 1;
    47: op1_12_inv01 = 1;
    51: op1_12_inv01 = 1;
    55: op1_12_inv01 = 1;
    56: op1_12_inv01 = 1;
    57: op1_12_inv01 = 1;
    59: op1_12_inv01 = 1;
    64: op1_12_inv01 = 1;
    68: op1_12_inv01 = 1;
    72: op1_12_inv01 = 1;
    74: op1_12_inv01 = 1;
    76: op1_12_inv01 = 1;
    78: op1_12_inv01 = 1;
    79: op1_12_inv01 = 1;
    81: op1_12_inv01 = 1;
    83: op1_12_inv01 = 1;
    84: op1_12_inv01 = 1;
    85: op1_12_inv01 = 1;
    88: op1_12_inv01 = 1;
    90: op1_12_inv01 = 1;
    91: op1_12_inv01 = 1;
    92: op1_12_inv01 = 1;
    95: op1_12_inv01 = 1;
    96: op1_12_inv01 = 1;
    default: op1_12_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in02 = reg_0304;
    81: op1_12_in02 = reg_0304;
    6: op1_12_in02 = reg_0818;
    7: op1_12_in02 = reg_0577;
    13: op1_12_in02 = reg_0577;
    8: op1_12_in02 = reg_0676;
    9: op1_12_in02 = imem04_in[91:88];
    10: op1_12_in02 = imem02_in[15:12];
    11: op1_12_in02 = imem06_in[19:16];
    12: op1_12_in02 = reg_0238;
    14: op1_12_in02 = imem00_in[35:32];
    15: op1_12_in02 = reg_0234;
    16: op1_12_in02 = reg_0061;
    17: op1_12_in02 = imem07_in[47:44];
    18: op1_12_in02 = reg_0970;
    19: op1_12_in02 = reg_0799;
    20: op1_12_in02 = reg_0736;
    21: op1_12_in02 = imem00_in[63:60];
    22: op1_12_in02 = reg_0007;
    23: op1_12_in02 = imem04_in[95:92];
    24: op1_12_in02 = imem03_in[27:24];
    25: op1_12_in02 = imem05_in[39:36];
    4: op1_12_in02 = imem07_in[103:100];
    26: op1_12_in02 = reg_1034;
    3: op1_12_in02 = reg_0175;
    27: op1_12_in02 = reg_0781;
    28: op1_12_in02 = reg_0608;
    29: op1_12_in02 = reg_0040;
    30: op1_12_in02 = reg_1006;
    31: op1_12_in02 = imem00_in[51:48];
    42: op1_12_in02 = imem00_in[51:48];
    88: op1_12_in02 = imem00_in[51:48];
    2: op1_12_in02 = imem07_in[95:92];
    32: op1_12_in02 = reg_0500;
    33: op1_12_in02 = imem02_in[11:8];
    34: op1_12_in02 = reg_0827;
    35: op1_12_in02 = imem00_in[31:28];
    73: op1_12_in02 = imem00_in[31:28];
    36: op1_12_in02 = imem00_in[107:104];
    37: op1_12_in02 = imem02_in[111:108];
    38: op1_12_in02 = imem00_in[43:40];
    39: op1_12_in02 = reg_0888;
    40: op1_12_in02 = reg_0525;
    41: op1_12_in02 = imem05_in[83:80];
    43: op1_12_in02 = imem02_in[63:60];
    44: op1_12_in02 = reg_0374;
    45: op1_12_in02 = reg_0707;
    46: op1_12_in02 = imem00_in[59:56];
    47: op1_12_in02 = reg_0807;
    49: op1_12_in02 = reg_0687;
    50: op1_12_in02 = reg_0534;
    51: op1_12_in02 = reg_0447;
    52: op1_12_in02 = reg_0373;
    53: op1_12_in02 = reg_0948;
    54: op1_12_in02 = imem05_in[11:8];
    55: op1_12_in02 = reg_0838;
    56: op1_12_in02 = imem00_in[95:92];
    57: op1_12_in02 = imem00_in[83:80];
    59: op1_12_in02 = reg_0671;
    60: op1_12_in02 = imem00_in[75:72];
    80: op1_12_in02 = imem00_in[75:72];
    61: op1_12_in02 = reg_0733;
    62: op1_12_in02 = imem04_in[63:60];
    63: op1_12_in02 = imem07_in[35:32];
    64: op1_12_in02 = reg_0011;
    65: op1_12_in02 = reg_0599;
    66: op1_12_in02 = imem00_in[55:52];
    70: op1_12_in02 = imem00_in[55:52];
    67: op1_12_in02 = reg_0161;
    68: op1_12_in02 = imem03_in[35:32];
    69: op1_12_in02 = imem05_in[27:24];
    71: op1_12_in02 = reg_0368;
    72: op1_12_in02 = reg_0222;
    74: op1_12_in02 = imem00_in[87:84];
    75: op1_12_in02 = reg_0737;
    76: op1_12_in02 = reg_0767;
    77: op1_12_in02 = imem06_in[79:76];
    78: op1_12_in02 = imem06_in[119:116];
    79: op1_12_in02 = reg_0915;
    82: op1_12_in02 = imem00_in[15:12];
    83: op1_12_in02 = reg_0057;
    84: op1_12_in02 = reg_0662;
    85: op1_12_in02 = imem00_in[47:44];
    86: op1_12_in02 = imem01_in[91:88];
    87: op1_12_in02 = reg_0137;
    89: op1_12_in02 = reg_0866;
    90: op1_12_in02 = reg_0047;
    91: op1_12_in02 = reg_0427;
    92: op1_12_in02 = imem02_in[99:96];
    93: op1_12_in02 = imem03_in[79:76];
    94: op1_12_in02 = reg_0578;
    95: op1_12_in02 = reg_0038;
    96: op1_12_in02 = reg_0547;
    default: op1_12_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv02 = 1;
    7: op1_12_inv02 = 1;
    9: op1_12_inv02 = 1;
    10: op1_12_inv02 = 1;
    11: op1_12_inv02 = 1;
    12: op1_12_inv02 = 1;
    14: op1_12_inv02 = 1;
    16: op1_12_inv02 = 1;
    19: op1_12_inv02 = 1;
    20: op1_12_inv02 = 1;
    22: op1_12_inv02 = 1;
    26: op1_12_inv02 = 1;
    3: op1_12_inv02 = 1;
    27: op1_12_inv02 = 1;
    28: op1_12_inv02 = 1;
    30: op1_12_inv02 = 1;
    32: op1_12_inv02 = 1;
    34: op1_12_inv02 = 1;
    39: op1_12_inv02 = 1;
    40: op1_12_inv02 = 1;
    41: op1_12_inv02 = 1;
    42: op1_12_inv02 = 1;
    44: op1_12_inv02 = 1;
    45: op1_12_inv02 = 1;
    47: op1_12_inv02 = 1;
    50: op1_12_inv02 = 1;
    51: op1_12_inv02 = 1;
    52: op1_12_inv02 = 1;
    54: op1_12_inv02 = 1;
    55: op1_12_inv02 = 1;
    56: op1_12_inv02 = 1;
    57: op1_12_inv02 = 1;
    59: op1_12_inv02 = 1;
    60: op1_12_inv02 = 1;
    62: op1_12_inv02 = 1;
    63: op1_12_inv02 = 1;
    65: op1_12_inv02 = 1;
    70: op1_12_inv02 = 1;
    74: op1_12_inv02 = 1;
    75: op1_12_inv02 = 1;
    78: op1_12_inv02 = 1;
    80: op1_12_inv02 = 1;
    85: op1_12_inv02 = 1;
    86: op1_12_inv02 = 1;
    88: op1_12_inv02 = 1;
    90: op1_12_inv02 = 1;
    91: op1_12_inv02 = 1;
    default: op1_12_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in03 = reg_0293;
    6: op1_12_in03 = reg_0582;
    7: op1_12_in03 = reg_0379;
    8: op1_12_in03 = reg_0689;
    9: op1_12_in03 = imem04_in[95:92];
    10: op1_12_in03 = imem02_in[31:28];
    11: op1_12_in03 = imem06_in[75:72];
    12: op1_12_in03 = reg_1050;
    13: op1_12_in03 = reg_0332;
    14: op1_12_in03 = imem00_in[51:48];
    15: op1_12_in03 = reg_0905;
    16: op1_12_in03 = reg_0062;
    17: op1_12_in03 = imem07_in[51:48];
    18: op1_12_in03 = reg_0950;
    19: op1_12_in03 = reg_0027;
    20: op1_12_in03 = reg_0517;
    21: op1_12_in03 = imem00_in[71:68];
    38: op1_12_in03 = imem00_in[71:68];
    73: op1_12_in03 = imem00_in[71:68];
    88: op1_12_in03 = imem00_in[71:68];
    22: op1_12_in03 = reg_0482;
    23: op1_12_in03 = imem04_in[127:124];
    24: op1_12_in03 = imem03_in[107:104];
    25: op1_12_in03 = imem05_in[47:44];
    4: op1_12_in03 = imem07_in[127:124];
    26: op1_12_in03 = reg_0105;
    3: op1_12_in03 = reg_0161;
    27: op1_12_in03 = reg_0798;
    28: op1_12_in03 = reg_0622;
    29: op1_12_in03 = reg_0311;
    30: op1_12_in03 = reg_0536;
    31: op1_12_in03 = imem00_in[67:64];
    2: op1_12_in03 = imem07_in[111:108];
    32: op1_12_in03 = reg_1031;
    33: op1_12_in03 = imem02_in[15:12];
    34: op1_12_in03 = reg_0252;
    35: op1_12_in03 = imem00_in[47:44];
    36: op1_12_in03 = reg_0676;
    37: op1_12_in03 = reg_0653;
    39: op1_12_in03 = reg_0537;
    40: op1_12_in03 = imem05_in[55:52];
    41: op1_12_in03 = reg_0955;
    42: op1_12_in03 = imem00_in[55:52];
    85: op1_12_in03 = imem00_in[55:52];
    43: op1_12_in03 = imem02_in[79:76];
    44: op1_12_in03 = reg_0991;
    45: op1_12_in03 = reg_0805;
    46: op1_12_in03 = imem00_in[75:72];
    70: op1_12_in03 = imem00_in[75:72];
    47: op1_12_in03 = reg_0376;
    49: op1_12_in03 = reg_0453;
    50: op1_12_in03 = reg_0624;
    51: op1_12_in03 = reg_0333;
    52: op1_12_in03 = reg_0051;
    53: op1_12_in03 = reg_0969;
    54: op1_12_in03 = imem05_in[23:20];
    55: op1_12_in03 = reg_0181;
    56: op1_12_in03 = reg_0682;
    57: op1_12_in03 = imem00_in[119:116];
    59: op1_12_in03 = reg_0843;
    60: op1_12_in03 = imem00_in[79:76];
    61: op1_12_in03 = reg_0113;
    62: op1_12_in03 = imem04_in[103:100];
    63: op1_12_in03 = imem07_in[59:56];
    64: op1_12_in03 = reg_0380;
    65: op1_12_in03 = reg_0350;
    66: op1_12_in03 = imem00_in[95:92];
    67: op1_12_in03 = reg_0162;
    68: op1_12_in03 = imem03_in[55:52];
    69: op1_12_in03 = imem05_in[91:88];
    71: op1_12_in03 = reg_0335;
    72: op1_12_in03 = reg_0695;
    74: op1_12_in03 = imem00_in[115:112];
    75: op1_12_in03 = reg_0610;
    76: op1_12_in03 = reg_0581;
    77: op1_12_in03 = reg_0080;
    78: op1_12_in03 = reg_1011;
    79: op1_12_in03 = reg_0755;
    80: op1_12_in03 = reg_0768;
    81: op1_12_in03 = reg_0273;
    82: op1_12_in03 = imem00_in[23:20];
    83: op1_12_in03 = reg_0150;
    84: op1_12_in03 = reg_0281;
    86: op1_12_in03 = imem01_in[119:116];
    87: op1_12_in03 = imem05_in[11:8];
    89: op1_12_in03 = reg_0492;
    90: op1_12_in03 = reg_0419;
    91: op1_12_in03 = reg_0868;
    92: op1_12_in03 = imem02_in[119:116];
    93: op1_12_in03 = reg_0758;
    94: op1_12_in03 = reg_0558;
    95: op1_12_in03 = reg_0239;
    96: op1_12_in03 = imem04_in[11:8];
    default: op1_12_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv03 = 1;
    8: op1_12_inv03 = 1;
    9: op1_12_inv03 = 1;
    12: op1_12_inv03 = 1;
    13: op1_12_inv03 = 1;
    15: op1_12_inv03 = 1;
    16: op1_12_inv03 = 1;
    17: op1_12_inv03 = 1;
    18: op1_12_inv03 = 1;
    20: op1_12_inv03 = 1;
    22: op1_12_inv03 = 1;
    24: op1_12_inv03 = 1;
    4: op1_12_inv03 = 1;
    27: op1_12_inv03 = 1;
    28: op1_12_inv03 = 1;
    2: op1_12_inv03 = 1;
    32: op1_12_inv03 = 1;
    35: op1_12_inv03 = 1;
    36: op1_12_inv03 = 1;
    37: op1_12_inv03 = 1;
    42: op1_12_inv03 = 1;
    43: op1_12_inv03 = 1;
    44: op1_12_inv03 = 1;
    47: op1_12_inv03 = 1;
    49: op1_12_inv03 = 1;
    50: op1_12_inv03 = 1;
    60: op1_12_inv03 = 1;
    61: op1_12_inv03 = 1;
    65: op1_12_inv03 = 1;
    66: op1_12_inv03 = 1;
    69: op1_12_inv03 = 1;
    75: op1_12_inv03 = 1;
    76: op1_12_inv03 = 1;
    78: op1_12_inv03 = 1;
    80: op1_12_inv03 = 1;
    83: op1_12_inv03 = 1;
    84: op1_12_inv03 = 1;
    85: op1_12_inv03 = 1;
    88: op1_12_inv03 = 1;
    90: op1_12_inv03 = 1;
    94: op1_12_inv03 = 1;
    95: op1_12_inv03 = 1;
    96: op1_12_inv03 = 1;
    default: op1_12_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in04 = reg_0290;
    6: op1_12_in04 = reg_0579;
    7: op1_12_in04 = reg_0371;
    8: op1_12_in04 = reg_0684;
    9: op1_12_in04 = reg_0530;
    10: op1_12_in04 = imem02_in[47:44];
    11: op1_12_in04 = reg_0614;
    12: op1_12_in04 = reg_0507;
    13: op1_12_in04 = reg_0375;
    14: op1_12_in04 = imem00_in[111:108];
    73: op1_12_in04 = imem00_in[111:108];
    15: op1_12_in04 = reg_0216;
    16: op1_12_in04 = reg_0065;
    17: op1_12_in04 = imem07_in[95:92];
    18: op1_12_in04 = reg_0945;
    19: op1_12_in04 = reg_1028;
    20: op1_12_in04 = reg_0056;
    21: op1_12_in04 = imem00_in[83:80];
    22: op1_12_in04 = reg_0085;
    23: op1_12_in04 = reg_0303;
    24: op1_12_in04 = imem03_in[119:116];
    25: op1_12_in04 = imem05_in[59:56];
    4: op1_12_in04 = reg_0424;
    26: op1_12_in04 = reg_0116;
    3: op1_12_in04 = reg_0167;
    27: op1_12_in04 = imem07_in[47:44];
    28: op1_12_in04 = reg_0615;
    29: op1_12_in04 = reg_0513;
    30: op1_12_in04 = reg_0301;
    31: op1_12_in04 = imem00_in[75:72];
    88: op1_12_in04 = imem00_in[75:72];
    32: op1_12_in04 = reg_1015;
    33: op1_12_in04 = imem02_in[63:60];
    34: op1_12_in04 = reg_0489;
    35: op1_12_in04 = imem00_in[99:96];
    36: op1_12_in04 = reg_0463;
    37: op1_12_in04 = reg_0639;
    38: op1_12_in04 = imem00_in[79:76];
    39: op1_12_in04 = reg_0764;
    40: op1_12_in04 = imem05_in[123:120];
    41: op1_12_in04 = reg_0956;
    42: op1_12_in04 = imem00_in[107:104];
    43: op1_12_in04 = imem02_in[83:80];
    44: op1_12_in04 = reg_0996;
    45: op1_12_in04 = reg_0361;
    46: op1_12_in04 = imem00_in[91:88];
    47: op1_12_in04 = reg_0518;
    49: op1_12_in04 = reg_0455;
    50: op1_12_in04 = reg_0856;
    51: op1_12_in04 = reg_0149;
    52: op1_12_in04 = reg_0987;
    53: op1_12_in04 = reg_0951;
    54: op1_12_in04 = imem05_in[27:24];
    55: op1_12_in04 = reg_0161;
    56: op1_12_in04 = reg_0685;
    57: op1_12_in04 = imem00_in[123:120];
    59: op1_12_in04 = reg_0680;
    60: op1_12_in04 = imem00_in[87:84];
    61: op1_12_in04 = imem02_in[55:52];
    62: op1_12_in04 = imem04_in[107:104];
    63: op1_12_in04 = imem07_in[107:104];
    64: op1_12_in04 = reg_0293;
    65: op1_12_in04 = reg_0502;
    66: op1_12_in04 = imem00_in[115:112];
    67: op1_12_in04 = reg_0183;
    68: op1_12_in04 = imem03_in[59:56];
    69: op1_12_in04 = imem05_in[107:104];
    70: op1_12_in04 = reg_0001;
    74: op1_12_in04 = reg_0001;
    71: op1_12_in04 = reg_0758;
    72: op1_12_in04 = reg_0857;
    75: op1_12_in04 = reg_0111;
    76: op1_12_in04 = reg_0233;
    77: op1_12_in04 = reg_0696;
    78: op1_12_in04 = reg_0926;
    79: op1_12_in04 = reg_0403;
    80: op1_12_in04 = reg_0523;
    81: op1_12_in04 = reg_0733;
    82: op1_12_in04 = imem00_in[27:24];
    83: op1_12_in04 = reg_0336;
    84: op1_12_in04 = reg_0385;
    85: op1_12_in04 = imem00_in[71:68];
    86: op1_12_in04 = reg_1042;
    87: op1_12_in04 = imem05_in[39:36];
    89: op1_12_in04 = reg_0235;
    90: op1_12_in04 = reg_0589;
    91: op1_12_in04 = reg_0431;
    92: op1_12_in04 = imem02_in[123:120];
    93: op1_12_in04 = reg_0596;
    94: op1_12_in04 = reg_0342;
    95: op1_12_in04 = reg_0230;
    96: op1_12_in04 = imem04_in[39:36];
    default: op1_12_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv04 = 1;
    9: op1_12_inv04 = 1;
    11: op1_12_inv04 = 1;
    13: op1_12_inv04 = 1;
    15: op1_12_inv04 = 1;
    16: op1_12_inv04 = 1;
    18: op1_12_inv04 = 1;
    22: op1_12_inv04 = 1;
    23: op1_12_inv04 = 1;
    24: op1_12_inv04 = 1;
    4: op1_12_inv04 = 1;
    3: op1_12_inv04 = 1;
    27: op1_12_inv04 = 1;
    31: op1_12_inv04 = 1;
    39: op1_12_inv04 = 1;
    40: op1_12_inv04 = 1;
    42: op1_12_inv04 = 1;
    44: op1_12_inv04 = 1;
    47: op1_12_inv04 = 1;
    49: op1_12_inv04 = 1;
    50: op1_12_inv04 = 1;
    51: op1_12_inv04 = 1;
    56: op1_12_inv04 = 1;
    59: op1_12_inv04 = 1;
    60: op1_12_inv04 = 1;
    61: op1_12_inv04 = 1;
    62: op1_12_inv04 = 1;
    63: op1_12_inv04 = 1;
    65: op1_12_inv04 = 1;
    69: op1_12_inv04 = 1;
    71: op1_12_inv04 = 1;
    75: op1_12_inv04 = 1;
    77: op1_12_inv04 = 1;
    79: op1_12_inv04 = 1;
    81: op1_12_inv04 = 1;
    82: op1_12_inv04 = 1;
    83: op1_12_inv04 = 1;
    84: op1_12_inv04 = 1;
    85: op1_12_inv04 = 1;
    86: op1_12_inv04 = 1;
    88: op1_12_inv04 = 1;
    89: op1_12_inv04 = 1;
    90: op1_12_inv04 = 1;
    91: op1_12_inv04 = 1;
    92: op1_12_inv04 = 1;
    94: op1_12_inv04 = 1;
    95: op1_12_inv04 = 1;
    default: op1_12_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in05 = reg_0291;
    6: op1_12_in05 = reg_0569;
    7: op1_12_in05 = reg_0375;
    8: op1_12_in05 = reg_0690;
    9: op1_12_in05 = reg_0539;
    10: op1_12_in05 = imem02_in[75:72];
    11: op1_12_in05 = reg_0610;
    12: op1_12_in05 = reg_0226;
    13: op1_12_in05 = reg_0315;
    14: op1_12_in05 = reg_0670;
    15: op1_12_in05 = reg_0913;
    16: op1_12_in05 = reg_0067;
    17: op1_12_in05 = imem07_in[107:104];
    18: op1_12_in05 = reg_0863;
    19: op1_12_in05 = reg_0018;
    20: op1_12_in05 = reg_0043;
    21: op1_12_in05 = imem00_in[107:104];
    22: op1_12_in05 = reg_0876;
    23: op1_12_in05 = reg_0833;
    24: op1_12_in05 = reg_0582;
    25: op1_12_in05 = imem05_in[119:116];
    4: op1_12_in05 = reg_0430;
    26: op1_12_in05 = reg_0102;
    3: op1_12_in05 = reg_0163;
    27: op1_12_in05 = imem07_in[79:76];
    28: op1_12_in05 = reg_0409;
    29: op1_12_in05 = reg_0246;
    86: op1_12_in05 = reg_0246;
    30: op1_12_in05 = reg_0265;
    31: op1_12_in05 = imem00_in[91:88];
    32: op1_12_in05 = reg_0871;
    33: op1_12_in05 = imem02_in[95:92];
    34: op1_12_in05 = reg_0148;
    35: op1_12_in05 = imem00_in[127:124];
    88: op1_12_in05 = imem00_in[127:124];
    36: op1_12_in05 = reg_0455;
    37: op1_12_in05 = reg_0648;
    38: op1_12_in05 = imem00_in[87:84];
    39: op1_12_in05 = reg_0066;
    40: op1_12_in05 = reg_0973;
    41: op1_12_in05 = reg_0949;
    53: op1_12_in05 = reg_0949;
    42: op1_12_in05 = imem00_in[123:120];
    46: op1_12_in05 = imem00_in[123:120];
    43: op1_12_in05 = imem02_in[87:84];
    44: op1_12_in05 = reg_0989;
    45: op1_12_in05 = reg_0744;
    47: op1_12_in05 = reg_0234;
    49: op1_12_in05 = reg_0476;
    50: op1_12_in05 = reg_0020;
    51: op1_12_in05 = reg_0136;
    52: op1_12_in05 = reg_1002;
    84: op1_12_in05 = reg_1002;
    54: op1_12_in05 = imem05_in[87:84];
    55: op1_12_in05 = reg_0159;
    56: op1_12_in05 = reg_0748;
    57: op1_12_in05 = reg_0685;
    59: op1_12_in05 = reg_0454;
    60: op1_12_in05 = imem00_in[111:108];
    61: op1_12_in05 = imem02_in[71:68];
    62: op1_12_in05 = imem04_in[115:112];
    63: op1_12_in05 = reg_0720;
    64: op1_12_in05 = reg_0946;
    65: op1_12_in05 = reg_0640;
    66: op1_12_in05 = imem00_in[119:116];
    67: op1_12_in05 = reg_0168;
    68: op1_12_in05 = imem03_in[63:60];
    69: op1_12_in05 = imem05_in[115:112];
    70: op1_12_in05 = reg_0519;
    71: op1_12_in05 = reg_0506;
    72: op1_12_in05 = reg_0403;
    73: op1_12_in05 = reg_0682;
    74: op1_12_in05 = reg_0523;
    75: op1_12_in05 = reg_0115;
    76: op1_12_in05 = reg_0266;
    77: op1_12_in05 = reg_1018;
    78: op1_12_in05 = reg_0534;
    79: op1_12_in05 = reg_0369;
    80: op1_12_in05 = reg_0883;
    81: op1_12_in05 = reg_0555;
    82: op1_12_in05 = imem00_in[31:28];
    83: op1_12_in05 = reg_0951;
    85: op1_12_in05 = imem00_in[75:72];
    87: op1_12_in05 = imem05_in[59:56];
    89: op1_12_in05 = reg_0268;
    90: op1_12_in05 = reg_0868;
    91: op1_12_in05 = reg_0175;
    92: op1_12_in05 = reg_0750;
    93: op1_12_in05 = reg_0239;
    94: op1_12_in05 = reg_0397;
    95: op1_12_in05 = reg_0051;
    96: op1_12_in05 = imem04_in[43:40];
    default: op1_12_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv05 = 1;
    6: op1_12_inv05 = 1;
    7: op1_12_inv05 = 1;
    8: op1_12_inv05 = 1;
    9: op1_12_inv05 = 1;
    10: op1_12_inv05 = 1;
    11: op1_12_inv05 = 1;
    12: op1_12_inv05 = 1;
    15: op1_12_inv05 = 1;
    16: op1_12_inv05 = 1;
    17: op1_12_inv05 = 1;
    19: op1_12_inv05 = 1;
    20: op1_12_inv05 = 1;
    23: op1_12_inv05 = 1;
    24: op1_12_inv05 = 1;
    28: op1_12_inv05 = 1;
    29: op1_12_inv05 = 1;
    30: op1_12_inv05 = 1;
    31: op1_12_inv05 = 1;
    32: op1_12_inv05 = 1;
    33: op1_12_inv05 = 1;
    34: op1_12_inv05 = 1;
    35: op1_12_inv05 = 1;
    37: op1_12_inv05 = 1;
    38: op1_12_inv05 = 1;
    40: op1_12_inv05 = 1;
    42: op1_12_inv05 = 1;
    44: op1_12_inv05 = 1;
    47: op1_12_inv05 = 1;
    49: op1_12_inv05 = 1;
    50: op1_12_inv05 = 1;
    52: op1_12_inv05 = 1;
    56: op1_12_inv05 = 1;
    57: op1_12_inv05 = 1;
    64: op1_12_inv05 = 1;
    65: op1_12_inv05 = 1;
    67: op1_12_inv05 = 1;
    70: op1_12_inv05 = 1;
    72: op1_12_inv05 = 1;
    74: op1_12_inv05 = 1;
    75: op1_12_inv05 = 1;
    77: op1_12_inv05 = 1;
    79: op1_12_inv05 = 1;
    81: op1_12_inv05 = 1;
    84: op1_12_inv05 = 1;
    85: op1_12_inv05 = 1;
    88: op1_12_inv05 = 1;
    89: op1_12_inv05 = 1;
    90: op1_12_inv05 = 1;
    96: op1_12_inv05 = 1;
    default: op1_12_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in06 = reg_0062;
    6: op1_12_in06 = reg_0592;
    7: op1_12_in06 = reg_0367;
    13: op1_12_in06 = reg_0367;
    8: op1_12_in06 = reg_0671;
    9: op1_12_in06 = reg_0555;
    10: op1_12_in06 = imem02_in[95:92];
    11: op1_12_in06 = reg_0613;
    12: op1_12_in06 = reg_0216;
    14: op1_12_in06 = reg_0690;
    15: op1_12_in06 = reg_1041;
    16: op1_12_in06 = reg_0057;
    17: op1_12_in06 = reg_0728;
    18: op1_12_in06 = reg_0826;
    19: op1_12_in06 = imem07_in[55:52];
    20: op1_12_in06 = reg_0021;
    21: op1_12_in06 = imem00_in[115:112];
    22: op1_12_in06 = reg_0086;
    23: op1_12_in06 = reg_0046;
    24: op1_12_in06 = reg_0573;
    25: op1_12_in06 = imem05_in[127:124];
    69: op1_12_in06 = imem05_in[127:124];
    4: op1_12_in06 = reg_0447;
    26: op1_12_in06 = reg_0114;
    81: op1_12_in06 = reg_0114;
    3: op1_12_in06 = reg_0164;
    27: op1_12_in06 = imem07_in[87:84];
    28: op1_12_in06 = reg_0401;
    29: op1_12_in06 = reg_0987;
    30: op1_12_in06 = reg_0537;
    31: op1_12_in06 = imem00_in[103:100];
    32: op1_12_in06 = reg_1034;
    33: op1_12_in06 = imem02_in[103:100];
    34: op1_12_in06 = reg_0143;
    35: op1_12_in06 = reg_0682;
    60: op1_12_in06 = reg_0682;
    66: op1_12_in06 = reg_0682;
    36: op1_12_in06 = reg_0464;
    37: op1_12_in06 = reg_0636;
    38: op1_12_in06 = imem00_in[95:92];
    39: op1_12_in06 = reg_0076;
    40: op1_12_in06 = reg_0971;
    41: op1_12_in06 = reg_0806;
    42: op1_12_in06 = reg_0683;
    43: op1_12_in06 = imem02_in[119:116];
    44: op1_12_in06 = reg_0983;
    45: op1_12_in06 = reg_0180;
    91: op1_12_in06 = reg_0180;
    46: op1_12_in06 = reg_0697;
    47: op1_12_in06 = reg_0985;
    49: op1_12_in06 = reg_0467;
    50: op1_12_in06 = reg_0892;
    51: op1_12_in06 = reg_0128;
    52: op1_12_in06 = reg_0991;
    53: op1_12_in06 = reg_0259;
    54: op1_12_in06 = imem05_in[91:88];
    55: op1_12_in06 = reg_0182;
    56: op1_12_in06 = reg_0102;
    57: op1_12_in06 = reg_0686;
    59: op1_12_in06 = reg_0480;
    61: op1_12_in06 = imem02_in[79:76];
    62: op1_12_in06 = reg_1006;
    63: op1_12_in06 = reg_0721;
    64: op1_12_in06 = reg_0264;
    65: op1_12_in06 = reg_0175;
    68: op1_12_in06 = imem03_in[67:64];
    70: op1_12_in06 = reg_0825;
    71: op1_12_in06 = reg_0261;
    72: op1_12_in06 = reg_0022;
    73: op1_12_in06 = reg_0748;
    74: op1_12_in06 = reg_0684;
    75: op1_12_in06 = reg_0110;
    76: op1_12_in06 = reg_0551;
    77: op1_12_in06 = reg_0294;
    78: op1_12_in06 = reg_0297;
    79: op1_12_in06 = reg_0566;
    80: op1_12_in06 = reg_0499;
    82: op1_12_in06 = imem00_in[43:40];
    83: op1_12_in06 = reg_0657;
    84: op1_12_in06 = imem04_in[3:0];
    85: op1_12_in06 = imem00_in[87:84];
    86: op1_12_in06 = reg_0973;
    87: op1_12_in06 = imem05_in[67:64];
    88: op1_12_in06 = reg_0523;
    89: op1_12_in06 = reg_0063;
    90: op1_12_in06 = reg_0024;
    92: op1_12_in06 = reg_0543;
    93: op1_12_in06 = reg_0961;
    94: op1_12_in06 = reg_1049;
    95: op1_12_in06 = reg_0779;
    96: op1_12_in06 = imem04_in[59:56];
    default: op1_12_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_12_inv06 = 1;
    8: op1_12_inv06 = 1;
    9: op1_12_inv06 = 1;
    10: op1_12_inv06 = 1;
    14: op1_12_inv06 = 1;
    15: op1_12_inv06 = 1;
    17: op1_12_inv06 = 1;
    18: op1_12_inv06 = 1;
    19: op1_12_inv06 = 1;
    20: op1_12_inv06 = 1;
    21: op1_12_inv06 = 1;
    22: op1_12_inv06 = 1;
    23: op1_12_inv06 = 1;
    24: op1_12_inv06 = 1;
    4: op1_12_inv06 = 1;
    3: op1_12_inv06 = 1;
    29: op1_12_inv06 = 1;
    35: op1_12_inv06 = 1;
    36: op1_12_inv06 = 1;
    40: op1_12_inv06 = 1;
    42: op1_12_inv06 = 1;
    44: op1_12_inv06 = 1;
    45: op1_12_inv06 = 1;
    46: op1_12_inv06 = 1;
    47: op1_12_inv06 = 1;
    49: op1_12_inv06 = 1;
    57: op1_12_inv06 = 1;
    60: op1_12_inv06 = 1;
    62: op1_12_inv06 = 1;
    63: op1_12_inv06 = 1;
    68: op1_12_inv06 = 1;
    70: op1_12_inv06 = 1;
    71: op1_12_inv06 = 1;
    73: op1_12_inv06 = 1;
    76: op1_12_inv06 = 1;
    78: op1_12_inv06 = 1;
    81: op1_12_inv06 = 1;
    82: op1_12_inv06 = 1;
    83: op1_12_inv06 = 1;
    84: op1_12_inv06 = 1;
    87: op1_12_inv06 = 1;
    89: op1_12_inv06 = 1;
    93: op1_12_inv06 = 1;
    95: op1_12_inv06 = 1;
    default: op1_12_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in07 = reg_0041;
    6: op1_12_in07 = reg_0584;
    7: op1_12_in07 = imem07_in[3:0];
    8: op1_12_in07 = reg_0678;
    9: op1_12_in07 = reg_0549;
    10: op1_12_in07 = reg_0656;
    11: op1_12_in07 = reg_0619;
    12: op1_12_in07 = reg_1035;
    13: op1_12_in07 = reg_0368;
    14: op1_12_in07 = reg_0668;
    15: op1_12_in07 = reg_0871;
    16: op1_12_in07 = imem05_in[23:20];
    17: op1_12_in07 = reg_0730;
    18: op1_12_in07 = reg_0835;
    19: op1_12_in07 = imem07_in[75:72];
    20: op1_12_in07 = reg_0483;
    21: op1_12_in07 = reg_0689;
    22: op1_12_in07 = imem03_in[3:0];
    23: op1_12_in07 = reg_0749;
    24: op1_12_in07 = reg_0587;
    25: op1_12_in07 = reg_0955;
    4: op1_12_in07 = reg_0445;
    93: op1_12_in07 = reg_0445;
    26: op1_12_in07 = reg_0324;
    3: op1_12_in07 = reg_0185;
    27: op1_12_in07 = imem07_in[119:116];
    28: op1_12_in07 = reg_0808;
    29: op1_12_in07 = reg_0995;
    47: op1_12_in07 = reg_0995;
    30: op1_12_in07 = reg_0068;
    31: op1_12_in07 = imem00_in[119:116];
    38: op1_12_in07 = imem00_in[119:116];
    32: op1_12_in07 = reg_0125;
    33: op1_12_in07 = imem02_in[123:120];
    43: op1_12_in07 = imem02_in[123:120];
    34: op1_12_in07 = reg_0140;
    35: op1_12_in07 = reg_0679;
    46: op1_12_in07 = reg_0679;
    36: op1_12_in07 = reg_0476;
    37: op1_12_in07 = reg_0916;
    39: op1_12_in07 = reg_0059;
    40: op1_12_in07 = reg_0948;
    41: op1_12_in07 = reg_0813;
    42: op1_12_in07 = reg_0696;
    44: op1_12_in07 = reg_0994;
    45: op1_12_in07 = reg_0167;
    49: op1_12_in07 = reg_0459;
    50: op1_12_in07 = reg_0781;
    51: op1_12_in07 = reg_0134;
    52: op1_12_in07 = reg_0989;
    53: op1_12_in07 = reg_0446;
    54: op1_12_in07 = imem05_in[111:108];
    55: op1_12_in07 = reg_0160;
    56: op1_12_in07 = reg_0680;
    57: op1_12_in07 = reg_0499;
    59: op1_12_in07 = reg_0210;
    60: op1_12_in07 = reg_0519;
    61: op1_12_in07 = imem02_in[91:88];
    62: op1_12_in07 = reg_0050;
    63: op1_12_in07 = reg_0703;
    64: op1_12_in07 = imem07_in[15:12];
    65: op1_12_in07 = reg_0161;
    66: op1_12_in07 = reg_0683;
    68: op1_12_in07 = imem03_in[71:68];
    69: op1_12_in07 = reg_0365;
    70: op1_12_in07 = reg_0684;
    71: op1_12_in07 = reg_0091;
    72: op1_12_in07 = imem07_in[67:64];
    73: op1_12_in07 = reg_0686;
    74: op1_12_in07 = reg_0753;
    75: op1_12_in07 = imem02_in[95:92];
    76: op1_12_in07 = reg_0998;
    77: op1_12_in07 = reg_0391;
    78: op1_12_in07 = reg_0533;
    79: op1_12_in07 = reg_0704;
    80: op1_12_in07 = reg_0467;
    81: op1_12_in07 = reg_0110;
    82: op1_12_in07 = imem00_in[47:44];
    83: op1_12_in07 = imem06_in[71:68];
    84: op1_12_in07 = imem04_in[115:112];
    85: op1_12_in07 = imem00_in[99:96];
    86: op1_12_in07 = reg_0968;
    87: op1_12_in07 = imem05_in[99:96];
    88: op1_12_in07 = reg_0748;
    89: op1_12_in07 = reg_0646;
    90: op1_12_in07 = reg_0431;
    91: op1_12_in07 = reg_0172;
    92: op1_12_in07 = reg_0277;
    94: op1_12_in07 = reg_0581;
    95: op1_12_in07 = reg_0597;
    96: op1_12_in07 = imem04_in[71:68];
    default: op1_12_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_12_inv07 = 1;
    10: op1_12_inv07 = 1;
    11: op1_12_inv07 = 1;
    13: op1_12_inv07 = 1;
    15: op1_12_inv07 = 1;
    17: op1_12_inv07 = 1;
    19: op1_12_inv07 = 1;
    20: op1_12_inv07 = 1;
    26: op1_12_inv07 = 1;
    3: op1_12_inv07 = 1;
    27: op1_12_inv07 = 1;
    28: op1_12_inv07 = 1;
    29: op1_12_inv07 = 1;
    31: op1_12_inv07 = 1;
    32: op1_12_inv07 = 1;
    33: op1_12_inv07 = 1;
    34: op1_12_inv07 = 1;
    38: op1_12_inv07 = 1;
    41: op1_12_inv07 = 1;
    47: op1_12_inv07 = 1;
    50: op1_12_inv07 = 1;
    52: op1_12_inv07 = 1;
    53: op1_12_inv07 = 1;
    54: op1_12_inv07 = 1;
    55: op1_12_inv07 = 1;
    56: op1_12_inv07 = 1;
    57: op1_12_inv07 = 1;
    65: op1_12_inv07 = 1;
    66: op1_12_inv07 = 1;
    68: op1_12_inv07 = 1;
    69: op1_12_inv07 = 1;
    70: op1_12_inv07 = 1;
    71: op1_12_inv07 = 1;
    73: op1_12_inv07 = 1;
    75: op1_12_inv07 = 1;
    76: op1_12_inv07 = 1;
    78: op1_12_inv07 = 1;
    81: op1_12_inv07 = 1;
    83: op1_12_inv07 = 1;
    84: op1_12_inv07 = 1;
    85: op1_12_inv07 = 1;
    93: op1_12_inv07 = 1;
    94: op1_12_inv07 = 1;
    95: op1_12_inv07 = 1;
    96: op1_12_inv07 = 1;
    default: op1_12_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in08 = imem05_in[3:0];
    6: op1_12_in08 = reg_0593;
    7: op1_12_in08 = imem07_in[27:24];
    8: op1_12_in08 = reg_0476;
    9: op1_12_in08 = reg_0533;
    10: op1_12_in08 = reg_0639;
    11: op1_12_in08 = reg_0608;
    12: op1_12_in08 = reg_0118;
    13: op1_12_in08 = reg_0787;
    14: op1_12_in08 = reg_0675;
    15: op1_12_in08 = reg_1017;
    16: op1_12_in08 = imem05_in[47:44];
    17: op1_12_in08 = reg_0731;
    18: op1_12_in08 = reg_0251;
    19: op1_12_in08 = imem07_in[99:96];
    72: op1_12_in08 = imem07_in[99:96];
    20: op1_12_in08 = reg_0530;
    21: op1_12_in08 = reg_0686;
    22: op1_12_in08 = imem03_in[23:20];
    23: op1_12_in08 = reg_0309;
    24: op1_12_in08 = reg_0360;
    25: op1_12_in08 = reg_0949;
    40: op1_12_in08 = reg_0949;
    4: op1_12_in08 = reg_0443;
    26: op1_12_in08 = reg_0073;
    3: op1_12_in08 = reg_0168;
    27: op1_12_in08 = reg_0710;
    28: op1_12_in08 = reg_0802;
    29: op1_12_in08 = reg_0986;
    30: op1_12_in08 = reg_0074;
    31: op1_12_in08 = reg_0695;
    32: op1_12_in08 = reg_0114;
    33: op1_12_in08 = reg_0645;
    34: op1_12_in08 = imem06_in[15:12];
    35: op1_12_in08 = reg_0674;
    36: op1_12_in08 = reg_0472;
    37: op1_12_in08 = reg_0318;
    38: op1_12_in08 = reg_0685;
    39: op1_12_in08 = reg_0864;
    41: op1_12_in08 = reg_0260;
    42: op1_12_in08 = reg_0698;
    43: op1_12_in08 = reg_0650;
    69: op1_12_in08 = reg_0650;
    44: op1_12_in08 = imem04_in[15:12];
    45: op1_12_in08 = reg_0159;
    46: op1_12_in08 = reg_0669;
    47: op1_12_in08 = reg_1000;
    49: op1_12_in08 = reg_0452;
    50: op1_12_in08 = reg_0556;
    51: op1_12_in08 = reg_0144;
    52: op1_12_in08 = reg_0981;
    53: op1_12_in08 = reg_0493;
    54: op1_12_in08 = reg_0973;
    55: op1_12_in08 = reg_0164;
    56: op1_12_in08 = reg_0828;
    57: op1_12_in08 = reg_0069;
    73: op1_12_in08 = reg_0069;
    59: op1_12_in08 = reg_0193;
    60: op1_12_in08 = reg_0883;
    61: op1_12_in08 = imem02_in[95:92];
    62: op1_12_in08 = reg_0066;
    63: op1_12_in08 = reg_0713;
    64: op1_12_in08 = imem07_in[123:120];
    65: op1_12_in08 = reg_0162;
    66: op1_12_in08 = reg_0825;
    68: op1_12_in08 = imem03_in[111:108];
    70: op1_12_in08 = reg_0842;
    71: op1_12_in08 = imem03_in[31:28];
    74: op1_12_in08 = reg_0450;
    75: op1_12_in08 = imem02_in[115:112];
    76: op1_12_in08 = reg_0996;
    77: op1_12_in08 = reg_0626;
    78: op1_12_in08 = reg_0032;
    79: op1_12_in08 = reg_0719;
    80: op1_12_in08 = reg_0470;
    81: op1_12_in08 = imem02_in[11:8];
    82: op1_12_in08 = imem00_in[51:48];
    83: op1_12_in08 = imem06_in[87:84];
    84: op1_12_in08 = reg_0048;
    85: op1_12_in08 = imem00_in[103:100];
    86: op1_12_in08 = reg_0337;
    87: op1_12_in08 = imem05_in[123:120];
    88: op1_12_in08 = reg_0684;
    89: op1_12_in08 = reg_0935;
    90: op1_12_in08 = reg_0175;
    91: op1_12_in08 = reg_0182;
    92: op1_12_in08 = reg_0090;
    93: op1_12_in08 = reg_0286;
    94: op1_12_in08 = reg_0445;
    95: op1_12_in08 = reg_0266;
    96: op1_12_in08 = imem04_in[79:76];
    default: op1_12_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv08 = 1;
    6: op1_12_inv08 = 1;
    7: op1_12_inv08 = 1;
    8: op1_12_inv08 = 1;
    12: op1_12_inv08 = 1;
    20: op1_12_inv08 = 1;
    22: op1_12_inv08 = 1;
    24: op1_12_inv08 = 1;
    25: op1_12_inv08 = 1;
    26: op1_12_inv08 = 1;
    3: op1_12_inv08 = 1;
    27: op1_12_inv08 = 1;
    32: op1_12_inv08 = 1;
    34: op1_12_inv08 = 1;
    36: op1_12_inv08 = 1;
    37: op1_12_inv08 = 1;
    40: op1_12_inv08 = 1;
    45: op1_12_inv08 = 1;
    46: op1_12_inv08 = 1;
    50: op1_12_inv08 = 1;
    51: op1_12_inv08 = 1;
    52: op1_12_inv08 = 1;
    53: op1_12_inv08 = 1;
    54: op1_12_inv08 = 1;
    55: op1_12_inv08 = 1;
    56: op1_12_inv08 = 1;
    59: op1_12_inv08 = 1;
    60: op1_12_inv08 = 1;
    61: op1_12_inv08 = 1;
    62: op1_12_inv08 = 1;
    63: op1_12_inv08 = 1;
    65: op1_12_inv08 = 1;
    66: op1_12_inv08 = 1;
    69: op1_12_inv08 = 1;
    71: op1_12_inv08 = 1;
    77: op1_12_inv08 = 1;
    79: op1_12_inv08 = 1;
    80: op1_12_inv08 = 1;
    84: op1_12_inv08 = 1;
    87: op1_12_inv08 = 1;
    88: op1_12_inv08 = 1;
    89: op1_12_inv08 = 1;
    90: op1_12_inv08 = 1;
    91: op1_12_inv08 = 1;
    94: op1_12_inv08 = 1;
    95: op1_12_inv08 = 1;
    96: op1_12_inv08 = 1;
    default: op1_12_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in09 = imem05_in[15:12];
    6: op1_12_in09 = reg_0580;
    7: op1_12_in09 = imem07_in[47:44];
    8: op1_12_in09 = reg_0466;
    9: op1_12_in09 = reg_0301;
    10: op1_12_in09 = reg_0651;
    69: op1_12_in09 = reg_0651;
    11: op1_12_in09 = reg_0627;
    12: op1_12_in09 = reg_0119;
    13: op1_12_in09 = reg_0486;
    14: op1_12_in09 = reg_0687;
    15: op1_12_in09 = reg_1038;
    16: op1_12_in09 = imem05_in[51:48];
    17: op1_12_in09 = reg_0714;
    18: op1_12_in09 = reg_0253;
    19: op1_12_in09 = imem07_in[103:100];
    20: op1_12_in09 = reg_0894;
    21: op1_12_in09 = reg_0679;
    22: op1_12_in09 = imem03_in[87:84];
    23: op1_12_in09 = reg_0529;
    24: op1_12_in09 = reg_0343;
    25: op1_12_in09 = reg_0968;
    4: op1_12_in09 = reg_0448;
    26: op1_12_in09 = reg_0793;
    3: op1_12_in09 = reg_0171;
    27: op1_12_in09 = reg_0726;
    28: op1_12_in09 = reg_0753;
    29: op1_12_in09 = reg_0983;
    30: op1_12_in09 = reg_0009;
    31: op1_12_in09 = reg_0697;
    32: op1_12_in09 = reg_0109;
    33: op1_12_in09 = reg_0655;
    34: op1_12_in09 = imem06_in[43:40];
    35: op1_12_in09 = reg_0450;
    36: op1_12_in09 = reg_0456;
    37: op1_12_in09 = reg_0857;
    38: op1_12_in09 = reg_0690;
    39: op1_12_in09 = reg_0963;
    40: op1_12_in09 = reg_0965;
    41: op1_12_in09 = reg_0132;
    42: op1_12_in09 = reg_0684;
    43: op1_12_in09 = reg_0654;
    44: op1_12_in09 = imem04_in[35:32];
    45: op1_12_in09 = reg_0157;
    46: op1_12_in09 = reg_0454;
    47: op1_12_in09 = imem04_in[3:0];
    49: op1_12_in09 = reg_0214;
    50: op1_12_in09 = reg_0889;
    51: op1_12_in09 = imem06_in[15:12];
    52: op1_12_in09 = imem04_in[19:16];
    53: op1_12_in09 = reg_0269;
    54: op1_12_in09 = reg_0957;
    56: op1_12_in09 = reg_0461;
    57: op1_12_in09 = reg_0680;
    60: op1_12_in09 = reg_0680;
    59: op1_12_in09 = reg_0194;
    61: op1_12_in09 = imem02_in[111:108];
    62: op1_12_in09 = reg_0064;
    63: op1_12_in09 = reg_0868;
    64: op1_12_in09 = imem07_in[127:124];
    65: op1_12_in09 = reg_0167;
    66: op1_12_in09 = reg_0670;
    68: op1_12_in09 = imem03_in[127:124];
    70: op1_12_in09 = reg_0356;
    71: op1_12_in09 = imem03_in[79:76];
    72: op1_12_in09 = imem07_in[123:120];
    73: op1_12_in09 = reg_0668;
    74: op1_12_in09 = reg_0469;
    75: op1_12_in09 = reg_0896;
    76: op1_12_in09 = reg_0993;
    77: op1_12_in09 = reg_1011;
    78: op1_12_in09 = reg_0383;
    79: op1_12_in09 = reg_0435;
    80: op1_12_in09 = reg_0478;
    81: op1_12_in09 = imem02_in[43:40];
    82: op1_12_in09 = imem00_in[63:60];
    83: op1_12_in09 = imem06_in[91:88];
    84: op1_12_in09 = reg_0430;
    85: op1_12_in09 = imem00_in[123:120];
    86: op1_12_in09 = reg_1023;
    87: op1_12_in09 = reg_0970;
    88: op1_12_in09 = reg_0686;
    89: op1_12_in09 = reg_0129;
    90: op1_12_in09 = reg_0429;
    91: op1_12_in09 = reg_0539;
    92: op1_12_in09 = reg_0095;
    93: op1_12_in09 = reg_0975;
    94: op1_12_in09 = reg_0988;
    95: op1_12_in09 = reg_0987;
    96: op1_12_in09 = imem04_in[87:84];
    default: op1_12_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv09 = 1;
    12: op1_12_inv09 = 1;
    13: op1_12_inv09 = 1;
    14: op1_12_inv09 = 1;
    15: op1_12_inv09 = 1;
    17: op1_12_inv09 = 1;
    18: op1_12_inv09 = 1;
    19: op1_12_inv09 = 1;
    22: op1_12_inv09 = 1;
    23: op1_12_inv09 = 1;
    24: op1_12_inv09 = 1;
    25: op1_12_inv09 = 1;
    26: op1_12_inv09 = 1;
    3: op1_12_inv09 = 1;
    27: op1_12_inv09 = 1;
    29: op1_12_inv09 = 1;
    30: op1_12_inv09 = 1;
    33: op1_12_inv09 = 1;
    34: op1_12_inv09 = 1;
    37: op1_12_inv09 = 1;
    38: op1_12_inv09 = 1;
    40: op1_12_inv09 = 1;
    44: op1_12_inv09 = 1;
    51: op1_12_inv09 = 1;
    52: op1_12_inv09 = 1;
    54: op1_12_inv09 = 1;
    57: op1_12_inv09 = 1;
    62: op1_12_inv09 = 1;
    63: op1_12_inv09 = 1;
    66: op1_12_inv09 = 1;
    70: op1_12_inv09 = 1;
    71: op1_12_inv09 = 1;
    73: op1_12_inv09 = 1;
    74: op1_12_inv09 = 1;
    75: op1_12_inv09 = 1;
    77: op1_12_inv09 = 1;
    78: op1_12_inv09 = 1;
    79: op1_12_inv09 = 1;
    82: op1_12_inv09 = 1;
    88: op1_12_inv09 = 1;
    89: op1_12_inv09 = 1;
    90: op1_12_inv09 = 1;
    95: op1_12_inv09 = 1;
    default: op1_12_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in10 = imem05_in[55:52];
    6: op1_12_in10 = reg_0578;
    7: op1_12_in10 = imem07_in[63:60];
    8: op1_12_in10 = reg_0471;
    9: op1_12_in10 = reg_0305;
    10: op1_12_in10 = reg_0648;
    11: op1_12_in10 = reg_0601;
    12: op1_12_in10 = reg_0108;
    13: op1_12_in10 = reg_0801;
    14: op1_12_in10 = reg_0460;
    74: op1_12_in10 = reg_0460;
    15: op1_12_in10 = reg_1018;
    16: op1_12_in10 = imem05_in[83:80];
    17: op1_12_in10 = reg_0715;
    18: op1_12_in10 = reg_0132;
    19: op1_12_in10 = imem07_in[111:108];
    20: op1_12_in10 = reg_0955;
    21: op1_12_in10 = reg_0691;
    22: op1_12_in10 = imem03_in[127:124];
    23: op1_12_in10 = reg_0750;
    24: op1_12_in10 = reg_0995;
    25: op1_12_in10 = reg_0953;
    4: op1_12_in10 = reg_0180;
    26: op1_12_in10 = reg_0655;
    27: op1_12_in10 = reg_0714;
    28: op1_12_in10 = reg_0018;
    29: op1_12_in10 = imem04_in[27:24];
    52: op1_12_in10 = imem04_in[27:24];
    30: op1_12_in10 = reg_0015;
    31: op1_12_in10 = reg_0679;
    32: op1_12_in10 = reg_0117;
    33: op1_12_in10 = reg_0637;
    34: op1_12_in10 = imem06_in[79:76];
    35: op1_12_in10 = reg_0451;
    36: op1_12_in10 = reg_0191;
    37: op1_12_in10 = reg_0516;
    38: op1_12_in10 = reg_0699;
    39: op1_12_in10 = reg_0959;
    40: op1_12_in10 = reg_0946;
    41: op1_12_in10 = reg_0140;
    42: op1_12_in10 = reg_0670;
    43: op1_12_in10 = reg_0660;
    44: op1_12_in10 = imem04_in[67:64];
    46: op1_12_in10 = reg_0466;
    47: op1_12_in10 = imem04_in[15:12];
    49: op1_12_in10 = reg_0187;
    50: op1_12_in10 = reg_0495;
    51: op1_12_in10 = imem06_in[27:24];
    53: op1_12_in10 = reg_0145;
    54: op1_12_in10 = reg_0969;
    56: op1_12_in10 = reg_0477;
    57: op1_12_in10 = reg_0476;
    59: op1_12_in10 = reg_0205;
    60: op1_12_in10 = reg_0465;
    61: op1_12_in10 = imem02_in[115:112];
    62: op1_12_in10 = reg_0893;
    63: op1_12_in10 = reg_0165;
    64: op1_12_in10 = reg_0704;
    65: op1_12_in10 = reg_0168;
    66: op1_12_in10 = reg_0883;
    68: op1_12_in10 = reg_0580;
    69: op1_12_in10 = reg_0528;
    70: op1_12_in10 = reg_0749;
    73: op1_12_in10 = reg_0749;
    71: op1_12_in10 = reg_0345;
    72: op1_12_in10 = reg_0721;
    75: op1_12_in10 = reg_0846;
    76: op1_12_in10 = reg_0978;
    77: op1_12_in10 = reg_0735;
    78: op1_12_in10 = reg_0782;
    79: op1_12_in10 = reg_0724;
    80: op1_12_in10 = reg_0214;
    81: op1_12_in10 = imem02_in[55:52];
    82: op1_12_in10 = imem00_in[67:64];
    83: op1_12_in10 = imem06_in[127:124];
    84: op1_12_in10 = reg_0540;
    85: op1_12_in10 = reg_0900;
    86: op1_12_in10 = reg_0592;
    87: op1_12_in10 = reg_0508;
    88: op1_12_in10 = reg_0356;
    89: op1_12_in10 = reg_0023;
    90: op1_12_in10 = reg_0731;
    91: op1_12_in10 = reg_0449;
    92: op1_12_in10 = reg_0425;
    93: op1_12_in10 = reg_0271;
    94: op1_12_in10 = imem04_in[11:8];
    95: op1_12_in10 = reg_0961;
    96: op1_12_in10 = imem04_in[91:88];
    default: op1_12_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv10 = 1;
    6: op1_12_inv10 = 1;
    7: op1_12_inv10 = 1;
    12: op1_12_inv10 = 1;
    13: op1_12_inv10 = 1;
    16: op1_12_inv10 = 1;
    18: op1_12_inv10 = 1;
    19: op1_12_inv10 = 1;
    20: op1_12_inv10 = 1;
    24: op1_12_inv10 = 1;
    25: op1_12_inv10 = 1;
    4: op1_12_inv10 = 1;
    26: op1_12_inv10 = 1;
    27: op1_12_inv10 = 1;
    31: op1_12_inv10 = 1;
    32: op1_12_inv10 = 1;
    33: op1_12_inv10 = 1;
    34: op1_12_inv10 = 1;
    38: op1_12_inv10 = 1;
    41: op1_12_inv10 = 1;
    42: op1_12_inv10 = 1;
    43: op1_12_inv10 = 1;
    46: op1_12_inv10 = 1;
    50: op1_12_inv10 = 1;
    51: op1_12_inv10 = 1;
    52: op1_12_inv10 = 1;
    56: op1_12_inv10 = 1;
    57: op1_12_inv10 = 1;
    62: op1_12_inv10 = 1;
    63: op1_12_inv10 = 1;
    64: op1_12_inv10 = 1;
    66: op1_12_inv10 = 1;
    69: op1_12_inv10 = 1;
    70: op1_12_inv10 = 1;
    73: op1_12_inv10 = 1;
    76: op1_12_inv10 = 1;
    77: op1_12_inv10 = 1;
    78: op1_12_inv10 = 1;
    79: op1_12_inv10 = 1;
    80: op1_12_inv10 = 1;
    83: op1_12_inv10 = 1;
    85: op1_12_inv10 = 1;
    87: op1_12_inv10 = 1;
    88: op1_12_inv10 = 1;
    92: op1_12_inv10 = 1;
    94: op1_12_inv10 = 1;
    95: op1_12_inv10 = 1;
    default: op1_12_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in11 = imem05_in[79:76];
    6: op1_12_in11 = reg_0360;
    7: op1_12_in11 = imem07_in[111:108];
    8: op1_12_in11 = reg_0452;
    9: op1_12_in11 = reg_0282;
    10: op1_12_in11 = reg_0638;
    11: op1_12_in11 = reg_0382;
    12: op1_12_in11 = reg_0102;
    13: op1_12_in11 = reg_0017;
    14: op1_12_in11 = reg_0471;
    15: op1_12_in11 = reg_0103;
    16: op1_12_in11 = imem05_in[95:92];
    17: op1_12_in11 = reg_0442;
    18: op1_12_in11 = reg_0145;
    19: op1_12_in11 = imem07_in[119:116];
    20: op1_12_in11 = reg_0961;
    21: op1_12_in11 = reg_0669;
    85: op1_12_in11 = reg_0669;
    22: op1_12_in11 = reg_0598;
    23: op1_12_in11 = reg_0062;
    24: op1_12_in11 = reg_0994;
    25: op1_12_in11 = reg_0256;
    4: op1_12_in11 = reg_0161;
    63: op1_12_in11 = reg_0161;
    26: op1_12_in11 = reg_0656;
    27: op1_12_in11 = reg_0702;
    28: op1_12_in11 = reg_1010;
    29: op1_12_in11 = imem04_in[31:28];
    30: op1_12_in11 = reg_0278;
    31: op1_12_in11 = reg_0476;
    35: op1_12_in11 = reg_0476;
    32: op1_12_in11 = imem02_in[7:4];
    33: op1_12_in11 = reg_0842;
    34: op1_12_in11 = reg_0631;
    36: op1_12_in11 = reg_0189;
    37: op1_12_in11 = reg_0772;
    38: op1_12_in11 = reg_0455;
    60: op1_12_in11 = reg_0455;
    39: op1_12_in11 = reg_0967;
    40: op1_12_in11 = reg_0947;
    41: op1_12_in11 = reg_0137;
    42: op1_12_in11 = reg_0668;
    43: op1_12_in11 = reg_0657;
    44: op1_12_in11 = imem04_in[75:72];
    46: op1_12_in11 = reg_0470;
    56: op1_12_in11 = reg_0470;
    73: op1_12_in11 = reg_0470;
    47: op1_12_in11 = imem04_in[23:20];
    49: op1_12_in11 = reg_0193;
    50: op1_12_in11 = reg_0356;
    51: op1_12_in11 = imem06_in[31:28];
    52: op1_12_in11 = imem04_in[63:60];
    53: op1_12_in11 = reg_0138;
    54: op1_12_in11 = reg_0950;
    57: op1_12_in11 = reg_0462;
    59: op1_12_in11 = reg_0190;
    61: op1_12_in11 = reg_0651;
    62: op1_12_in11 = reg_0658;
    64: op1_12_in11 = reg_0708;
    66: op1_12_in11 = reg_0828;
    88: op1_12_in11 = reg_0828;
    68: op1_12_in11 = reg_0576;
    69: op1_12_in11 = reg_0030;
    70: op1_12_in11 = reg_0463;
    71: op1_12_in11 = reg_0681;
    72: op1_12_in11 = reg_0714;
    74: op1_12_in11 = reg_0467;
    75: op1_12_in11 = reg_0082;
    76: op1_12_in11 = reg_0974;
    77: op1_12_in11 = reg_0889;
    78: op1_12_in11 = reg_0369;
    79: op1_12_in11 = reg_0729;
    80: op1_12_in11 = reg_0188;
    81: op1_12_in11 = imem02_in[67:64];
    82: op1_12_in11 = imem00_in[71:68];
    83: op1_12_in11 = reg_0625;
    84: op1_12_in11 = reg_0016;
    86: op1_12_in11 = reg_0234;
    87: op1_12_in11 = reg_0490;
    89: op1_12_in11 = reg_0260;
    90: op1_12_in11 = reg_0723;
    91: op1_12_in11 = reg_0529;
    92: op1_12_in11 = reg_0818;
    93: op1_12_in11 = imem04_in[19:16];
    94: op1_12_in11 = imem04_in[43:40];
    95: op1_12_in11 = reg_0523;
    96: op1_12_in11 = imem04_in[107:104];
    default: op1_12_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_12_inv11 = 1;
    8: op1_12_inv11 = 1;
    9: op1_12_inv11 = 1;
    10: op1_12_inv11 = 1;
    13: op1_12_inv11 = 1;
    14: op1_12_inv11 = 1;
    22: op1_12_inv11 = 1;
    23: op1_12_inv11 = 1;
    26: op1_12_inv11 = 1;
    27: op1_12_inv11 = 1;
    29: op1_12_inv11 = 1;
    30: op1_12_inv11 = 1;
    32: op1_12_inv11 = 1;
    34: op1_12_inv11 = 1;
    35: op1_12_inv11 = 1;
    36: op1_12_inv11 = 1;
    37: op1_12_inv11 = 1;
    39: op1_12_inv11 = 1;
    43: op1_12_inv11 = 1;
    47: op1_12_inv11 = 1;
    49: op1_12_inv11 = 1;
    52: op1_12_inv11 = 1;
    53: op1_12_inv11 = 1;
    54: op1_12_inv11 = 1;
    57: op1_12_inv11 = 1;
    61: op1_12_inv11 = 1;
    63: op1_12_inv11 = 1;
    66: op1_12_inv11 = 1;
    68: op1_12_inv11 = 1;
    69: op1_12_inv11 = 1;
    70: op1_12_inv11 = 1;
    72: op1_12_inv11 = 1;
    76: op1_12_inv11 = 1;
    79: op1_12_inv11 = 1;
    80: op1_12_inv11 = 1;
    81: op1_12_inv11 = 1;
    82: op1_12_inv11 = 1;
    85: op1_12_inv11 = 1;
    86: op1_12_inv11 = 1;
    87: op1_12_inv11 = 1;
    88: op1_12_inv11 = 1;
    89: op1_12_inv11 = 1;
    92: op1_12_inv11 = 1;
    95: op1_12_inv11 = 1;
    default: op1_12_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in12 = imem05_in[119:116];
    16: op1_12_in12 = imem05_in[119:116];
    6: op1_12_in12 = reg_0370;
    7: op1_12_in12 = reg_0728;
    8: op1_12_in12 = reg_0187;
    73: op1_12_in12 = reg_0187;
    9: op1_12_in12 = reg_0285;
    10: op1_12_in12 = reg_0667;
    11: op1_12_in12 = reg_0403;
    12: op1_12_in12 = reg_0101;
    13: op1_12_in12 = reg_1010;
    14: op1_12_in12 = reg_0468;
    15: op1_12_in12 = reg_0118;
    17: op1_12_in12 = reg_0443;
    18: op1_12_in12 = reg_0142;
    19: op1_12_in12 = imem07_in[127:124];
    20: op1_12_in12 = imem05_in[63:60];
    21: op1_12_in12 = reg_0454;
    85: op1_12_in12 = reg_0454;
    22: op1_12_in12 = reg_0572;
    23: op1_12_in12 = reg_0071;
    24: op1_12_in12 = reg_0548;
    25: op1_12_in12 = reg_0757;
    4: op1_12_in12 = reg_0169;
    26: op1_12_in12 = reg_0639;
    27: op1_12_in12 = reg_0715;
    28: op1_12_in12 = reg_1011;
    29: op1_12_in12 = imem04_in[43:40];
    30: op1_12_in12 = reg_0059;
    31: op1_12_in12 = reg_0466;
    35: op1_12_in12 = reg_0466;
    32: op1_12_in12 = imem02_in[15:12];
    33: op1_12_in12 = reg_0080;
    34: op1_12_in12 = reg_0622;
    36: op1_12_in12 = reg_0204;
    37: op1_12_in12 = reg_0083;
    38: op1_12_in12 = reg_0462;
    39: op1_12_in12 = reg_0956;
    40: op1_12_in12 = reg_0827;
    41: op1_12_in12 = imem06_in[55:52];
    42: op1_12_in12 = reg_0450;
    43: op1_12_in12 = reg_0334;
    44: op1_12_in12 = imem04_in[83:80];
    46: op1_12_in12 = reg_0456;
    47: op1_12_in12 = imem04_in[67:64];
    49: op1_12_in12 = reg_0207;
    50: op1_12_in12 = reg_0391;
    51: op1_12_in12 = imem06_in[35:32];
    87: op1_12_in12 = imem06_in[35:32];
    52: op1_12_in12 = imem04_in[75:72];
    53: op1_12_in12 = reg_0130;
    54: op1_12_in12 = reg_0951;
    56: op1_12_in12 = reg_0459;
    74: op1_12_in12 = reg_0459;
    57: op1_12_in12 = reg_0480;
    59: op1_12_in12 = imem01_in[55:52];
    60: op1_12_in12 = reg_0464;
    61: op1_12_in12 = reg_0647;
    62: op1_12_in12 = reg_0856;
    63: op1_12_in12 = reg_0162;
    64: op1_12_in12 = reg_0419;
    66: op1_12_in12 = reg_0453;
    68: op1_12_in12 = reg_0038;
    69: op1_12_in12 = reg_0326;
    70: op1_12_in12 = reg_0457;
    71: op1_12_in12 = reg_0046;
    72: op1_12_in12 = reg_0729;
    75: op1_12_in12 = reg_0886;
    76: op1_12_in12 = reg_0988;
    77: op1_12_in12 = reg_0028;
    78: op1_12_in12 = reg_0566;
    79: op1_12_in12 = reg_0789;
    80: op1_12_in12 = reg_0201;
    81: op1_12_in12 = imem02_in[103:100];
    82: op1_12_in12 = imem00_in[103:100];
    83: op1_12_in12 = reg_0393;
    84: op1_12_in12 = reg_0909;
    86: op1_12_in12 = reg_0862;
    88: op1_12_in12 = reg_0753;
    89: op1_12_in12 = reg_0657;
    90: op1_12_in12 = reg_0339;
    92: op1_12_in12 = reg_0087;
    93: op1_12_in12 = imem04_in[55:52];
    94: op1_12_in12 = imem04_in[51:48];
    95: op1_12_in12 = reg_0445;
    96: op1_12_in12 = reg_0405;
    default: op1_12_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_12_inv12 = 1;
    11: op1_12_inv12 = 1;
    12: op1_12_inv12 = 1;
    13: op1_12_inv12 = 1;
    16: op1_12_inv12 = 1;
    18: op1_12_inv12 = 1;
    19: op1_12_inv12 = 1;
    21: op1_12_inv12 = 1;
    22: op1_12_inv12 = 1;
    25: op1_12_inv12 = 1;
    26: op1_12_inv12 = 1;
    29: op1_12_inv12 = 1;
    30: op1_12_inv12 = 1;
    31: op1_12_inv12 = 1;
    32: op1_12_inv12 = 1;
    33: op1_12_inv12 = 1;
    34: op1_12_inv12 = 1;
    38: op1_12_inv12 = 1;
    39: op1_12_inv12 = 1;
    41: op1_12_inv12 = 1;
    46: op1_12_inv12 = 1;
    54: op1_12_inv12 = 1;
    57: op1_12_inv12 = 1;
    63: op1_12_inv12 = 1;
    68: op1_12_inv12 = 1;
    69: op1_12_inv12 = 1;
    70: op1_12_inv12 = 1;
    71: op1_12_inv12 = 1;
    73: op1_12_inv12 = 1;
    75: op1_12_inv12 = 1;
    79: op1_12_inv12 = 1;
    80: op1_12_inv12 = 1;
    81: op1_12_inv12 = 1;
    84: op1_12_inv12 = 1;
    85: op1_12_inv12 = 1;
    89: op1_12_inv12 = 1;
    90: op1_12_inv12 = 1;
    92: op1_12_inv12 = 1;
    93: op1_12_inv12 = 1;
    default: op1_12_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in13 = reg_0490;
    6: op1_12_in13 = reg_0312;
    7: op1_12_in13 = reg_0719;
    19: op1_12_in13 = reg_0719;
    8: op1_12_in13 = reg_0203;
    9: op1_12_in13 = reg_0275;
    10: op1_12_in13 = reg_0352;
    11: op1_12_in13 = reg_0315;
    12: op1_12_in13 = reg_0109;
    13: op1_12_in13 = reg_0805;
    14: op1_12_in13 = reg_0452;
    15: op1_12_in13 = reg_0116;
    16: op1_12_in13 = reg_0944;
    17: op1_12_in13 = reg_0420;
    18: op1_12_in13 = reg_0139;
    20: op1_12_in13 = imem05_in[75:72];
    21: op1_12_in13 = reg_0477;
    42: op1_12_in13 = reg_0477;
    22: op1_12_in13 = reg_0587;
    23: op1_12_in13 = reg_0732;
    24: op1_12_in13 = reg_0546;
    25: op1_12_in13 = reg_0252;
    4: op1_12_in13 = reg_0177;
    26: op1_12_in13 = reg_0644;
    27: op1_12_in13 = reg_0701;
    28: op1_12_in13 = imem07_in[3:0];
    29: op1_12_in13 = imem04_in[59:56];
    93: op1_12_in13 = imem04_in[59:56];
    30: op1_12_in13 = reg_0736;
    31: op1_12_in13 = reg_0462;
    35: op1_12_in13 = reg_0462;
    32: op1_12_in13 = imem02_in[55:52];
    33: op1_12_in13 = reg_0095;
    34: op1_12_in13 = reg_0391;
    36: op1_12_in13 = reg_0188;
    37: op1_12_in13 = reg_0007;
    38: op1_12_in13 = reg_0471;
    39: op1_12_in13 = reg_0950;
    40: op1_12_in13 = reg_0757;
    41: op1_12_in13 = imem06_in[87:84];
    43: op1_12_in13 = reg_0339;
    44: op1_12_in13 = imem04_in[87:84];
    46: op1_12_in13 = reg_0193;
    47: op1_12_in13 = reg_0301;
    49: op1_12_in13 = reg_0186;
    50: op1_12_in13 = reg_0804;
    51: op1_12_in13 = imem06_in[39:36];
    52: op1_12_in13 = imem04_in[111:108];
    53: op1_12_in13 = reg_0131;
    54: op1_12_in13 = reg_0952;
    69: op1_12_in13 = reg_0952;
    56: op1_12_in13 = reg_0208;
    57: op1_12_in13 = reg_0189;
    59: op1_12_in13 = reg_0904;
    86: op1_12_in13 = reg_0904;
    60: op1_12_in13 = reg_0466;
    61: op1_12_in13 = reg_0643;
    62: op1_12_in13 = reg_0044;
    63: op1_12_in13 = reg_0169;
    64: op1_12_in13 = reg_0428;
    66: op1_12_in13 = reg_0455;
    68: op1_12_in13 = reg_0509;
    70: op1_12_in13 = reg_0464;
    71: op1_12_in13 = reg_0396;
    72: op1_12_in13 = reg_0708;
    73: op1_12_in13 = reg_0211;
    74: op1_12_in13 = reg_0200;
    75: op1_12_in13 = reg_0098;
    76: op1_12_in13 = reg_1000;
    77: op1_12_in13 = reg_0534;
    78: op1_12_in13 = imem07_in[23:20];
    79: op1_12_in13 = imem07_in[43:40];
    80: op1_12_in13 = reg_0202;
    81: op1_12_in13 = reg_0666;
    82: op1_12_in13 = imem00_in[107:104];
    83: op1_12_in13 = reg_0338;
    84: op1_12_in13 = reg_0064;
    85: op1_12_in13 = reg_0457;
    87: op1_12_in13 = imem06_in[71:68];
    88: op1_12_in13 = reg_0465;
    89: op1_12_in13 = reg_0046;
    90: op1_12_in13 = reg_0183;
    92: op1_12_in13 = reg_0037;
    94: op1_12_in13 = imem04_in[103:100];
    95: op1_12_in13 = imem04_in[43:40];
    96: op1_12_in13 = reg_0550;
    default: op1_12_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv13 = 1;
    7: op1_12_inv13 = 1;
    9: op1_12_inv13 = 1;
    11: op1_12_inv13 = 1;
    13: op1_12_inv13 = 1;
    15: op1_12_inv13 = 1;
    17: op1_12_inv13 = 1;
    18: op1_12_inv13 = 1;
    19: op1_12_inv13 = 1;
    23: op1_12_inv13 = 1;
    24: op1_12_inv13 = 1;
    25: op1_12_inv13 = 1;
    4: op1_12_inv13 = 1;
    26: op1_12_inv13 = 1;
    27: op1_12_inv13 = 1;
    30: op1_12_inv13 = 1;
    31: op1_12_inv13 = 1;
    34: op1_12_inv13 = 1;
    36: op1_12_inv13 = 1;
    40: op1_12_inv13 = 1;
    42: op1_12_inv13 = 1;
    43: op1_12_inv13 = 1;
    44: op1_12_inv13 = 1;
    47: op1_12_inv13 = 1;
    49: op1_12_inv13 = 1;
    51: op1_12_inv13 = 1;
    52: op1_12_inv13 = 1;
    53: op1_12_inv13 = 1;
    54: op1_12_inv13 = 1;
    57: op1_12_inv13 = 1;
    60: op1_12_inv13 = 1;
    68: op1_12_inv13 = 1;
    69: op1_12_inv13 = 1;
    73: op1_12_inv13 = 1;
    75: op1_12_inv13 = 1;
    79: op1_12_inv13 = 1;
    82: op1_12_inv13 = 1;
    83: op1_12_inv13 = 1;
    84: op1_12_inv13 = 1;
    85: op1_12_inv13 = 1;
    86: op1_12_inv13 = 1;
    89: op1_12_inv13 = 1;
    92: op1_12_inv13 = 1;
    94: op1_12_inv13 = 1;
    96: op1_12_inv13 = 1;
    default: op1_12_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in14 = reg_0491;
    6: op1_12_in14 = reg_0393;
    7: op1_12_in14 = reg_0707;
    72: op1_12_in14 = reg_0707;
    8: op1_12_in14 = reg_0190;
    9: op1_12_in14 = reg_0065;
    10: op1_12_in14 = reg_0364;
    11: op1_12_in14 = reg_0808;
    12: op1_12_in14 = reg_0110;
    13: op1_12_in14 = reg_0783;
    14: op1_12_in14 = reg_0478;
    15: op1_12_in14 = reg_0119;
    16: op1_12_in14 = reg_0955;
    17: op1_12_in14 = reg_0448;
    18: op1_12_in14 = reg_0140;
    19: op1_12_in14 = reg_0717;
    20: op1_12_in14 = imem05_in[87:84];
    21: op1_12_in14 = reg_0469;
    22: op1_12_in14 = reg_0589;
    23: op1_12_in14 = reg_0748;
    24: op1_12_in14 = reg_0297;
    25: op1_12_in14 = reg_0813;
    4: op1_12_in14 = reg_0164;
    26: op1_12_in14 = imem02_in[47:44];
    27: op1_12_in14 = reg_0424;
    28: op1_12_in14 = imem07_in[23:20];
    29: op1_12_in14 = imem04_in[83:80];
    93: op1_12_in14 = imem04_in[83:80];
    30: op1_12_in14 = reg_0738;
    31: op1_12_in14 = reg_0467;
    35: op1_12_in14 = reg_0467;
    32: op1_12_in14 = imem02_in[59:56];
    33: op1_12_in14 = reg_0039;
    75: op1_12_in14 = reg_0039;
    34: op1_12_in14 = reg_0386;
    36: op1_12_in14 = reg_0201;
    37: op1_12_in14 = reg_0088;
    38: op1_12_in14 = reg_0187;
    57: op1_12_in14 = reg_0187;
    39: op1_12_in14 = reg_0947;
    40: op1_12_in14 = reg_0816;
    41: op1_12_in14 = imem06_in[103:100];
    42: op1_12_in14 = reg_0462;
    43: op1_12_in14 = reg_0082;
    44: op1_12_in14 = imem04_in[95:92];
    46: op1_12_in14 = reg_0207;
    47: op1_12_in14 = reg_1003;
    49: op1_12_in14 = reg_0232;
    50: op1_12_in14 = reg_1029;
    51: op1_12_in14 = imem06_in[67:64];
    52: op1_12_in14 = reg_0530;
    53: op1_12_in14 = imem06_in[3:0];
    54: op1_12_in14 = reg_0023;
    56: op1_12_in14 = reg_0191;
    59: op1_12_in14 = reg_0919;
    60: op1_12_in14 = reg_0473;
    61: op1_12_in14 = reg_0645;
    62: op1_12_in14 = imem05_in[47:44];
    63: op1_12_in14 = reg_0168;
    64: op1_12_in14 = reg_0868;
    66: op1_12_in14 = reg_0464;
    68: op1_12_in14 = reg_0377;
    69: op1_12_in14 = reg_0689;
    70: op1_12_in14 = reg_0477;
    85: op1_12_in14 = reg_0477;
    71: op1_12_in14 = reg_0576;
    73: op1_12_in14 = reg_0194;
    74: op1_12_in14 = reg_0208;
    76: op1_12_in14 = imem04_in[35:32];
    77: op1_12_in14 = reg_0439;
    78: op1_12_in14 = imem07_in[27:24];
    79: op1_12_in14 = imem07_in[47:44];
    80: op1_12_in14 = reg_0206;
    81: op1_12_in14 = reg_0803;
    82: op1_12_in14 = imem00_in[111:108];
    83: op1_12_in14 = reg_0817;
    84: op1_12_in14 = reg_0432;
    86: op1_12_in14 = reg_0607;
    87: op1_12_in14 = reg_0080;
    88: op1_12_in14 = reg_0455;
    89: op1_12_in14 = reg_0876;
    90: op1_12_in14 = reg_0184;
    92: op1_12_in14 = reg_0408;
    94: op1_12_in14 = reg_0126;
    95: op1_12_in14 = imem04_in[111:108];
    96: op1_12_in14 = reg_1009;
    default: op1_12_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv14 = 1;
    6: op1_12_inv14 = 1;
    7: op1_12_inv14 = 1;
    9: op1_12_inv14 = 1;
    10: op1_12_inv14 = 1;
    11: op1_12_inv14 = 1;
    12: op1_12_inv14 = 1;
    13: op1_12_inv14 = 1;
    14: op1_12_inv14 = 1;
    16: op1_12_inv14 = 1;
    21: op1_12_inv14 = 1;
    24: op1_12_inv14 = 1;
    28: op1_12_inv14 = 1;
    33: op1_12_inv14 = 1;
    34: op1_12_inv14 = 1;
    35: op1_12_inv14 = 1;
    36: op1_12_inv14 = 1;
    40: op1_12_inv14 = 1;
    41: op1_12_inv14 = 1;
    42: op1_12_inv14 = 1;
    43: op1_12_inv14 = 1;
    44: op1_12_inv14 = 1;
    52: op1_12_inv14 = 1;
    54: op1_12_inv14 = 1;
    57: op1_12_inv14 = 1;
    59: op1_12_inv14 = 1;
    60: op1_12_inv14 = 1;
    61: op1_12_inv14 = 1;
    69: op1_12_inv14 = 1;
    70: op1_12_inv14 = 1;
    72: op1_12_inv14 = 1;
    75: op1_12_inv14 = 1;
    77: op1_12_inv14 = 1;
    78: op1_12_inv14 = 1;
    79: op1_12_inv14 = 1;
    82: op1_12_inv14 = 1;
    83: op1_12_inv14 = 1;
    85: op1_12_inv14 = 1;
    87: op1_12_inv14 = 1;
    93: op1_12_inv14 = 1;
    94: op1_12_inv14 = 1;
    default: op1_12_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in15 = reg_0492;
    6: op1_12_in15 = reg_0331;
    7: op1_12_in15 = reg_0430;
    8: op1_12_in15 = reg_0202;
    38: op1_12_in15 = reg_0202;
    9: op1_12_in15 = reg_0064;
    10: op1_12_in15 = reg_0341;
    11: op1_12_in15 = imem07_in[11:8];
    12: op1_12_in15 = imem02_in[19:16];
    13: op1_12_in15 = imem07_in[3:0];
    14: op1_12_in15 = reg_0193;
    15: op1_12_in15 = imem02_in[11:8];
    16: op1_12_in15 = reg_0969;
    17: op1_12_in15 = reg_0165;
    18: op1_12_in15 = imem06_in[15:12];
    19: op1_12_in15 = reg_0709;
    20: op1_12_in15 = imem05_in[107:104];
    62: op1_12_in15 = imem05_in[107:104];
    21: op1_12_in15 = reg_0460;
    22: op1_12_in15 = reg_0584;
    23: op1_12_in15 = reg_0043;
    24: op1_12_in15 = reg_0559;
    25: op1_12_in15 = reg_0257;
    4: op1_12_in15 = reg_0185;
    26: op1_12_in15 = imem02_in[63:60];
    32: op1_12_in15 = imem02_in[63:60];
    27: op1_12_in15 = reg_0426;
    28: op1_12_in15 = imem07_in[39:36];
    29: op1_12_in15 = reg_0483;
    30: op1_12_in15 = reg_0517;
    31: op1_12_in15 = reg_0191;
    42: op1_12_in15 = reg_0191;
    33: op1_12_in15 = reg_0886;
    34: op1_12_in15 = reg_0741;
    35: op1_12_in15 = reg_0459;
    36: op1_12_in15 = reg_0212;
    37: op1_12_in15 = reg_0867;
    39: op1_12_in15 = reg_0821;
    40: op1_12_in15 = reg_0275;
    41: op1_12_in15 = reg_0624;
    43: op1_12_in15 = reg_0772;
    44: op1_12_in15 = reg_1004;
    46: op1_12_in15 = reg_0199;
    47: op1_12_in15 = reg_1057;
    49: op1_12_in15 = reg_0560;
    50: op1_12_in15 = reg_0629;
    51: op1_12_in15 = imem06_in[107:104];
    52: op1_12_in15 = reg_1003;
    53: op1_12_in15 = imem06_in[43:40];
    54: op1_12_in15 = reg_0436;
    56: op1_12_in15 = reg_0187;
    57: op1_12_in15 = reg_0207;
    59: op1_12_in15 = reg_0798;
    60: op1_12_in15 = reg_0474;
    61: op1_12_in15 = reg_0358;
    63: op1_12_in15 = reg_0171;
    64: op1_12_in15 = reg_0640;
    66: op1_12_in15 = reg_0469;
    85: op1_12_in15 = reg_0469;
    68: op1_12_in15 = reg_0991;
    69: op1_12_in15 = reg_0966;
    70: op1_12_in15 = reg_0473;
    71: op1_12_in15 = reg_0377;
    72: op1_12_in15 = reg_0727;
    73: op1_12_in15 = reg_0205;
    74: op1_12_in15 = imem01_in[35:32];
    75: op1_12_in15 = reg_0389;
    76: op1_12_in15 = imem04_in[87:84];
    77: op1_12_in15 = reg_0591;
    78: op1_12_in15 = imem07_in[31:28];
    79: op1_12_in15 = imem07_in[59:56];
    80: op1_12_in15 = reg_0192;
    81: op1_12_in15 = reg_0096;
    82: op1_12_in15 = reg_0001;
    83: op1_12_in15 = reg_0926;
    84: op1_12_in15 = reg_0407;
    86: op1_12_in15 = reg_0522;
    87: op1_12_in15 = reg_0696;
    88: op1_12_in15 = reg_0477;
    89: op1_12_in15 = reg_0865;
    92: op1_12_in15 = reg_0085;
    93: op1_12_in15 = imem04_in[127:124];
    94: op1_12_in15 = reg_0511;
    95: op1_12_in15 = imem04_in[115:112];
    96: op1_12_in15 = reg_0870;
    default: op1_12_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv15 = 1;
    6: op1_12_inv15 = 1;
    8: op1_12_inv15 = 1;
    10: op1_12_inv15 = 1;
    12: op1_12_inv15 = 1;
    13: op1_12_inv15 = 1;
    15: op1_12_inv15 = 1;
    16: op1_12_inv15 = 1;
    17: op1_12_inv15 = 1;
    19: op1_12_inv15 = 1;
    20: op1_12_inv15 = 1;
    21: op1_12_inv15 = 1;
    22: op1_12_inv15 = 1;
    4: op1_12_inv15 = 1;
    27: op1_12_inv15 = 1;
    35: op1_12_inv15 = 1;
    37: op1_12_inv15 = 1;
    39: op1_12_inv15 = 1;
    42: op1_12_inv15 = 1;
    43: op1_12_inv15 = 1;
    46: op1_12_inv15 = 1;
    50: op1_12_inv15 = 1;
    51: op1_12_inv15 = 1;
    54: op1_12_inv15 = 1;
    56: op1_12_inv15 = 1;
    60: op1_12_inv15 = 1;
    63: op1_12_inv15 = 1;
    64: op1_12_inv15 = 1;
    66: op1_12_inv15 = 1;
    68: op1_12_inv15 = 1;
    70: op1_12_inv15 = 1;
    71: op1_12_inv15 = 1;
    74: op1_12_inv15 = 1;
    75: op1_12_inv15 = 1;
    80: op1_12_inv15 = 1;
    82: op1_12_inv15 = 1;
    84: op1_12_inv15 = 1;
    86: op1_12_inv15 = 1;
    87: op1_12_inv15 = 1;
    88: op1_12_inv15 = 1;
    89: op1_12_inv15 = 1;
    95: op1_12_inv15 = 1;
    default: op1_12_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in16 = reg_0493;
    6: op1_12_in16 = imem03_in[3:0];
    7: op1_12_in16 = reg_0442;
    8: op1_12_in16 = imem01_in[3:0];
    9: op1_12_in16 = reg_0050;
    10: op1_12_in16 = reg_0359;
    11: op1_12_in16 = imem07_in[39:36];
    12: op1_12_in16 = imem02_in[51:48];
    13: op1_12_in16 = imem07_in[23:20];
    14: op1_12_in16 = reg_0211;
    15: op1_12_in16 = imem02_in[39:36];
    16: op1_12_in16 = reg_0951;
    17: op1_12_in16 = reg_0166;
    18: op1_12_in16 = imem06_in[35:32];
    19: op1_12_in16 = reg_0713;
    20: op1_12_in16 = imem05_in[123:120];
    21: op1_12_in16 = reg_0479;
    22: op1_12_in16 = reg_0588;
    23: op1_12_in16 = reg_0854;
    24: op1_12_in16 = reg_0556;
    89: op1_12_in16 = reg_0556;
    25: op1_12_in16 = reg_0260;
    40: op1_12_in16 = reg_0260;
    4: op1_12_in16 = reg_0168;
    26: op1_12_in16 = imem02_in[71:68];
    27: op1_12_in16 = reg_0446;
    28: op1_12_in16 = imem07_in[47:44];
    29: op1_12_in16 = reg_1006;
    30: op1_12_in16 = imem05_in[3:0];
    31: op1_12_in16 = reg_0188;
    32: op1_12_in16 = imem02_in[83:80];
    33: op1_12_in16 = reg_0085;
    34: op1_12_in16 = reg_0382;
    35: op1_12_in16 = reg_0452;
    36: op1_12_in16 = imem01_in[19:16];
    37: op1_12_in16 = reg_0792;
    38: op1_12_in16 = imem01_in[7:4];
    73: op1_12_in16 = imem01_in[7:4];
    80: op1_12_in16 = imem01_in[7:4];
    39: op1_12_in16 = reg_0022;
    41: op1_12_in16 = reg_0533;
    42: op1_12_in16 = reg_0210;
    43: op1_12_in16 = reg_0876;
    44: op1_12_in16 = reg_0536;
    46: op1_12_in16 = imem01_in[63:60];
    47: op1_12_in16 = reg_0932;
    49: op1_12_in16 = reg_0849;
    50: op1_12_in16 = reg_0596;
    51: op1_12_in16 = imem06_in[111:108];
    52: op1_12_in16 = reg_1009;
    53: op1_12_in16 = imem06_in[59:56];
    54: op1_12_in16 = reg_0094;
    56: op1_12_in16 = reg_0209;
    57: op1_12_in16 = reg_0199;
    59: op1_12_in16 = reg_1041;
    60: op1_12_in16 = reg_0458;
    61: op1_12_in16 = reg_0739;
    62: op1_12_in16 = reg_0020;
    64: op1_12_in16 = reg_0175;
    66: op1_12_in16 = reg_0476;
    85: op1_12_in16 = reg_0476;
    68: op1_12_in16 = reg_0992;
    69: op1_12_in16 = reg_0935;
    70: op1_12_in16 = reg_0194;
    71: op1_12_in16 = reg_0820;
    72: op1_12_in16 = reg_0805;
    74: op1_12_in16 = imem01_in[51:48];
    75: op1_12_in16 = reg_0425;
    76: op1_12_in16 = imem04_in[91:88];
    77: op1_12_in16 = reg_0804;
    78: op1_12_in16 = imem07_in[71:68];
    79: op1_12_in16 = imem07_in[67:64];
    81: op1_12_in16 = reg_0886;
    82: op1_12_in16 = reg_0841;
    83: op1_12_in16 = reg_0222;
    84: op1_12_in16 = reg_0041;
    86: op1_12_in16 = reg_0830;
    87: op1_12_in16 = reg_1018;
    88: op1_12_in16 = reg_0473;
    92: op1_12_in16 = reg_0381;
    93: op1_12_in16 = reg_0147;
    94: op1_12_in16 = reg_0802;
    95: op1_12_in16 = imem04_in[119:116];
    96: op1_12_in16 = reg_0048;
    default: op1_12_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv16 = 1;
    7: op1_12_inv16 = 1;
    8: op1_12_inv16 = 1;
    9: op1_12_inv16 = 1;
    11: op1_12_inv16 = 1;
    12: op1_12_inv16 = 1;
    14: op1_12_inv16 = 1;
    16: op1_12_inv16 = 1;
    18: op1_12_inv16 = 1;
    19: op1_12_inv16 = 1;
    22: op1_12_inv16 = 1;
    4: op1_12_inv16 = 1;
    26: op1_12_inv16 = 1;
    29: op1_12_inv16 = 1;
    30: op1_12_inv16 = 1;
    31: op1_12_inv16 = 1;
    33: op1_12_inv16 = 1;
    35: op1_12_inv16 = 1;
    36: op1_12_inv16 = 1;
    38: op1_12_inv16 = 1;
    39: op1_12_inv16 = 1;
    40: op1_12_inv16 = 1;
    41: op1_12_inv16 = 1;
    49: op1_12_inv16 = 1;
    50: op1_12_inv16 = 1;
    51: op1_12_inv16 = 1;
    53: op1_12_inv16 = 1;
    54: op1_12_inv16 = 1;
    57: op1_12_inv16 = 1;
    59: op1_12_inv16 = 1;
    60: op1_12_inv16 = 1;
    62: op1_12_inv16 = 1;
    66: op1_12_inv16 = 1;
    69: op1_12_inv16 = 1;
    71: op1_12_inv16 = 1;
    72: op1_12_inv16 = 1;
    73: op1_12_inv16 = 1;
    74: op1_12_inv16 = 1;
    76: op1_12_inv16 = 1;
    77: op1_12_inv16 = 1;
    79: op1_12_inv16 = 1;
    82: op1_12_inv16 = 1;
    83: op1_12_inv16 = 1;
    84: op1_12_inv16 = 1;
    85: op1_12_inv16 = 1;
    87: op1_12_inv16 = 1;
    92: op1_12_inv16 = 1;
    93: op1_12_inv16 = 1;
    default: op1_12_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in17 = reg_0494;
    6: op1_12_in17 = imem03_in[23:20];
    7: op1_12_in17 = reg_0172;
    64: op1_12_in17 = reg_0172;
    8: op1_12_in17 = imem01_in[27:24];
    38: op1_12_in17 = imem01_in[27:24];
    9: op1_12_in17 = imem05_in[47:44];
    10: op1_12_in17 = reg_0330;
    11: op1_12_in17 = imem07_in[55:52];
    12: op1_12_in17 = imem02_in[59:56];
    13: op1_12_in17 = imem07_in[35:32];
    14: op1_12_in17 = reg_0205;
    15: op1_12_in17 = imem02_in[47:44];
    16: op1_12_in17 = reg_0942;
    17: op1_12_in17 = reg_0164;
    18: op1_12_in17 = imem06_in[39:36];
    19: op1_12_in17 = reg_0429;
    20: op1_12_in17 = reg_0143;
    21: op1_12_in17 = reg_0459;
    22: op1_12_in17 = reg_0576;
    23: op1_12_in17 = reg_0855;
    24: op1_12_in17 = imem04_in[11:8];
    25: op1_12_in17 = reg_1046;
    4: op1_12_in17 = reg_0178;
    26: op1_12_in17 = imem02_in[103:100];
    27: op1_12_in17 = reg_0438;
    28: op1_12_in17 = imem07_in[59:56];
    29: op1_12_in17 = reg_0301;
    30: op1_12_in17 = imem05_in[35:32];
    31: op1_12_in17 = reg_0186;
    32: op1_12_in17 = imem02_in[111:108];
    33: op1_12_in17 = reg_0814;
    37: op1_12_in17 = reg_0814;
    34: op1_12_in17 = reg_0349;
    35: op1_12_in17 = reg_0210;
    36: op1_12_in17 = imem01_in[31:28];
    39: op1_12_in17 = reg_0835;
    40: op1_12_in17 = reg_0831;
    41: op1_12_in17 = reg_0020;
    42: op1_12_in17 = imem01_in[35:32];
    43: op1_12_in17 = reg_0090;
    44: op1_12_in17 = reg_0306;
    52: op1_12_in17 = reg_0306;
    46: op1_12_in17 = reg_0013;
    47: op1_12_in17 = reg_0050;
    49: op1_12_in17 = reg_0272;
    50: op1_12_in17 = reg_0008;
    51: op1_12_in17 = reg_0895;
    53: op1_12_in17 = imem06_in[83:80];
    54: op1_12_in17 = reg_0489;
    56: op1_12_in17 = reg_0188;
    57: op1_12_in17 = imem01_in[15:12];
    59: op1_12_in17 = reg_0116;
    60: op1_12_in17 = reg_0214;
    61: op1_12_in17 = reg_0359;
    62: op1_12_in17 = reg_0237;
    66: op1_12_in17 = reg_0470;
    68: op1_12_in17 = reg_0995;
    69: op1_12_in17 = reg_0675;
    70: op1_12_in17 = reg_0202;
    71: op1_12_in17 = reg_0233;
    72: op1_12_in17 = reg_0361;
    73: op1_12_in17 = imem01_in[23:20];
    74: op1_12_in17 = imem01_in[71:68];
    75: op1_12_in17 = reg_0335;
    76: op1_12_in17 = imem04_in[107:104];
    77: op1_12_in17 = reg_0699;
    78: op1_12_in17 = imem07_in[107:104];
    79: op1_12_in17 = imem07_in[71:68];
    80: op1_12_in17 = imem01_in[11:8];
    81: op1_12_in17 = reg_0323;
    82: op1_12_in17 = reg_0671;
    83: op1_12_in17 = reg_0695;
    84: op1_12_in17 = reg_0065;
    85: op1_12_in17 = reg_0466;
    86: op1_12_in17 = reg_0902;
    87: op1_12_in17 = reg_0384;
    88: op1_12_in17 = reg_0200;
    89: op1_12_in17 = reg_0338;
    92: op1_12_in17 = reg_0778;
    93: op1_12_in17 = reg_0577;
    94: op1_12_in17 = reg_0076;
    95: op1_12_in17 = imem04_in[127:124];
    96: op1_12_in17 = reg_0430;
    default: op1_12_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv17 = 1;
    9: op1_12_inv17 = 1;
    11: op1_12_inv17 = 1;
    15: op1_12_inv17 = 1;
    18: op1_12_inv17 = 1;
    20: op1_12_inv17 = 1;
    25: op1_12_inv17 = 1;
    28: op1_12_inv17 = 1;
    29: op1_12_inv17 = 1;
    32: op1_12_inv17 = 1;
    33: op1_12_inv17 = 1;
    34: op1_12_inv17 = 1;
    36: op1_12_inv17 = 1;
    37: op1_12_inv17 = 1;
    40: op1_12_inv17 = 1;
    42: op1_12_inv17 = 1;
    47: op1_12_inv17 = 1;
    49: op1_12_inv17 = 1;
    50: op1_12_inv17 = 1;
    51: op1_12_inv17 = 1;
    53: op1_12_inv17 = 1;
    54: op1_12_inv17 = 1;
    61: op1_12_inv17 = 1;
    64: op1_12_inv17 = 1;
    68: op1_12_inv17 = 1;
    69: op1_12_inv17 = 1;
    70: op1_12_inv17 = 1;
    71: op1_12_inv17 = 1;
    72: op1_12_inv17 = 1;
    73: op1_12_inv17 = 1;
    74: op1_12_inv17 = 1;
    78: op1_12_inv17 = 1;
    79: op1_12_inv17 = 1;
    80: op1_12_inv17 = 1;
    82: op1_12_inv17 = 1;
    83: op1_12_inv17 = 1;
    85: op1_12_inv17 = 1;
    88: op1_12_inv17 = 1;
    92: op1_12_inv17 = 1;
    94: op1_12_inv17 = 1;
    95: op1_12_inv17 = 1;
    96: op1_12_inv17 = 1;
    default: op1_12_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in18 = reg_0495;
    84: op1_12_in18 = reg_0495;
    6: op1_12_in18 = imem03_in[35:32];
    7: op1_12_in18 = reg_0161;
    8: op1_12_in18 = imem01_in[39:36];
    36: op1_12_in18 = imem01_in[39:36];
    42: op1_12_in18 = imem01_in[39:36];
    9: op1_12_in18 = imem05_in[75:72];
    10: op1_12_in18 = reg_0092;
    11: op1_12_in18 = imem07_in[63:60];
    12: op1_12_in18 = imem02_in[95:92];
    13: op1_12_in18 = imem07_in[39:36];
    14: op1_12_in18 = reg_0199;
    15: op1_12_in18 = imem02_in[51:48];
    16: op1_12_in18 = reg_0945;
    17: op1_12_in18 = reg_0176;
    18: op1_12_in18 = imem06_in[99:96];
    19: op1_12_in18 = reg_0436;
    20: op1_12_in18 = reg_0153;
    21: op1_12_in18 = reg_0214;
    22: op1_12_in18 = reg_0360;
    23: op1_12_in18 = reg_0856;
    24: op1_12_in18 = imem04_in[47:44];
    25: op1_12_in18 = reg_0489;
    26: op1_12_in18 = reg_0088;
    27: op1_12_in18 = reg_0431;
    28: op1_12_in18 = imem07_in[71:68];
    29: op1_12_in18 = reg_0265;
    30: op1_12_in18 = reg_0962;
    31: op1_12_in18 = reg_0196;
    32: op1_12_in18 = reg_0647;
    33: op1_12_in18 = reg_0091;
    34: op1_12_in18 = reg_0599;
    35: op1_12_in18 = reg_0211;
    37: op1_12_in18 = reg_0086;
    38: op1_12_in18 = imem01_in[119:116];
    39: op1_12_in18 = reg_0900;
    40: op1_12_in18 = reg_0135;
    41: op1_12_in18 = reg_0892;
    43: op1_12_in18 = reg_0084;
    44: op1_12_in18 = reg_1057;
    46: op1_12_in18 = reg_0299;
    47: op1_12_in18 = reg_0524;
    49: op1_12_in18 = reg_0224;
    50: op1_12_in18 = imem07_in[87:84];
    51: op1_12_in18 = reg_0220;
    52: op1_12_in18 = reg_0539;
    53: op1_12_in18 = reg_0619;
    54: op1_12_in18 = reg_0152;
    56: op1_12_in18 = reg_0203;
    57: op1_12_in18 = imem01_in[35:32];
    59: op1_12_in18 = reg_0860;
    60: op1_12_in18 = reg_0201;
    61: op1_12_in18 = reg_0394;
    62: op1_12_in18 = reg_0942;
    64: op1_12_in18 = reg_0167;
    66: op1_12_in18 = reg_0458;
    68: op1_12_in18 = reg_0977;
    69: op1_12_in18 = reg_0603;
    70: op1_12_in18 = imem01_in[11:8];
    71: op1_12_in18 = reg_0266;
    72: op1_12_in18 = reg_0419;
    73: op1_12_in18 = imem01_in[51:48];
    74: op1_12_in18 = imem01_in[75:72];
    75: op1_12_in18 = reg_0347;
    76: op1_12_in18 = imem04_in[127:124];
    77: op1_12_in18 = reg_0917;
    78: op1_12_in18 = reg_0529;
    79: op1_12_in18 = imem07_in[83:80];
    80: op1_12_in18 = imem01_in[47:44];
    81: op1_12_in18 = reg_0052;
    82: op1_12_in18 = reg_0685;
    83: op1_12_in18 = reg_0289;
    85: op1_12_in18 = reg_0205;
    86: op1_12_in18 = reg_0111;
    87: op1_12_in18 = reg_0379;
    88: op1_12_in18 = reg_0189;
    89: op1_12_in18 = reg_0926;
    92: op1_12_in18 = reg_0886;
    93: op1_12_in18 = reg_0937;
    94: op1_12_in18 = reg_0056;
    95: op1_12_in18 = reg_0550;
    96: op1_12_in18 = reg_0008;
    default: op1_12_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv18 = 1;
    11: op1_12_inv18 = 1;
    12: op1_12_inv18 = 1;
    13: op1_12_inv18 = 1;
    14: op1_12_inv18 = 1;
    17: op1_12_inv18 = 1;
    18: op1_12_inv18 = 1;
    22: op1_12_inv18 = 1;
    23: op1_12_inv18 = 1;
    24: op1_12_inv18 = 1;
    25: op1_12_inv18 = 1;
    29: op1_12_inv18 = 1;
    33: op1_12_inv18 = 1;
    34: op1_12_inv18 = 1;
    35: op1_12_inv18 = 1;
    36: op1_12_inv18 = 1;
    37: op1_12_inv18 = 1;
    38: op1_12_inv18 = 1;
    39: op1_12_inv18 = 1;
    41: op1_12_inv18 = 1;
    43: op1_12_inv18 = 1;
    47: op1_12_inv18 = 1;
    49: op1_12_inv18 = 1;
    50: op1_12_inv18 = 1;
    51: op1_12_inv18 = 1;
    53: op1_12_inv18 = 1;
    54: op1_12_inv18 = 1;
    60: op1_12_inv18 = 1;
    62: op1_12_inv18 = 1;
    64: op1_12_inv18 = 1;
    68: op1_12_inv18 = 1;
    69: op1_12_inv18 = 1;
    70: op1_12_inv18 = 1;
    72: op1_12_inv18 = 1;
    73: op1_12_inv18 = 1;
    74: op1_12_inv18 = 1;
    75: op1_12_inv18 = 1;
    76: op1_12_inv18 = 1;
    77: op1_12_inv18 = 1;
    78: op1_12_inv18 = 1;
    79: op1_12_inv18 = 1;
    80: op1_12_inv18 = 1;
    81: op1_12_inv18 = 1;
    83: op1_12_inv18 = 1;
    88: op1_12_inv18 = 1;
    93: op1_12_inv18 = 1;
    default: op1_12_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in19 = reg_0262;
    6: op1_12_in19 = imem04_in[7:4];
    7: op1_12_in19 = reg_0163;
    8: op1_12_in19 = imem01_in[83:80];
    9: op1_12_in19 = imem05_in[127:124];
    10: op1_12_in19 = reg_0088;
    11: op1_12_in19 = imem07_in[103:100];
    12: op1_12_in19 = imem02_in[123:120];
    13: op1_12_in19 = imem07_in[75:72];
    14: op1_12_in19 = imem01_in[27:24];
    15: op1_12_in19 = reg_0642;
    16: op1_12_in19 = reg_0952;
    18: op1_12_in19 = reg_0611;
    19: op1_12_in19 = reg_0447;
    20: op1_12_in19 = reg_0155;
    21: op1_12_in19 = reg_0210;
    22: op1_12_in19 = reg_0343;
    23: op1_12_in19 = imem05_in[71:68];
    24: op1_12_in19 = imem04_in[55:52];
    25: op1_12_in19 = reg_0147;
    26: op1_12_in19 = reg_0876;
    27: op1_12_in19 = reg_0179;
    28: op1_12_in19 = imem07_in[83:80];
    29: op1_12_in19 = reg_1009;
    30: op1_12_in19 = reg_0963;
    31: op1_12_in19 = reg_0205;
    32: op1_12_in19 = reg_0640;
    33: op1_12_in19 = reg_0016;
    34: op1_12_in19 = reg_0596;
    35: op1_12_in19 = reg_0201;
    36: op1_12_in19 = imem01_in[71:68];
    37: op1_12_in19 = reg_0090;
    38: op1_12_in19 = reg_0239;
    39: op1_12_in19 = reg_0135;
    40: op1_12_in19 = reg_0133;
    41: op1_12_in19 = reg_0577;
    42: op1_12_in19 = imem01_in[103:100];
    73: op1_12_in19 = imem01_in[103:100];
    43: op1_12_in19 = imem03_in[79:76];
    44: op1_12_in19 = reg_0058;
    46: op1_12_in19 = reg_0544;
    47: op1_12_in19 = reg_0808;
    49: op1_12_in19 = reg_0810;
    50: op1_12_in19 = imem07_in[107:104];
    51: op1_12_in19 = reg_0892;
    52: op1_12_in19 = reg_0540;
    53: op1_12_in19 = reg_0403;
    54: op1_12_in19 = reg_0154;
    56: op1_12_in19 = reg_0196;
    57: op1_12_in19 = imem01_in[55:52];
    59: op1_12_in19 = reg_0117;
    60: op1_12_in19 = reg_0190;
    61: op1_12_in19 = reg_0608;
    62: op1_12_in19 = reg_0333;
    64: op1_12_in19 = reg_0182;
    66: op1_12_in19 = reg_0207;
    68: op1_12_in19 = reg_0990;
    69: op1_12_in19 = reg_0819;
    70: op1_12_in19 = imem01_in[23:20];
    71: op1_12_in19 = reg_0982;
    72: op1_12_in19 = reg_0589;
    74: op1_12_in19 = reg_1042;
    75: op1_12_in19 = reg_0772;
    76: op1_12_in19 = reg_1006;
    77: op1_12_in19 = reg_0619;
    78: op1_12_in19 = reg_0123;
    79: op1_12_in19 = imem07_in[115:112];
    80: op1_12_in19 = reg_0105;
    81: op1_12_in19 = reg_0368;
    82: op1_12_in19 = reg_0825;
    83: op1_12_in19 = reg_0485;
    84: op1_12_in19 = reg_0854;
    85: op1_12_in19 = reg_0195;
    86: op1_12_in19 = reg_0733;
    87: op1_12_in19 = reg_0320;
    88: op1_12_in19 = reg_0187;
    89: op1_12_in19 = reg_0792;
    92: op1_12_in19 = reg_0730;
    93: op1_12_in19 = reg_0306;
    94: op1_12_in19 = reg_0064;
    95: op1_12_in19 = reg_0156;
    96: op1_12_in19 = reg_0586;
    default: op1_12_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_12_inv19 = 1;
    11: op1_12_inv19 = 1;
    12: op1_12_inv19 = 1;
    13: op1_12_inv19 = 1;
    14: op1_12_inv19 = 1;
    18: op1_12_inv19 = 1;
    19: op1_12_inv19 = 1;
    20: op1_12_inv19 = 1;
    21: op1_12_inv19 = 1;
    22: op1_12_inv19 = 1;
    24: op1_12_inv19 = 1;
    25: op1_12_inv19 = 1;
    26: op1_12_inv19 = 1;
    29: op1_12_inv19 = 1;
    31: op1_12_inv19 = 1;
    33: op1_12_inv19 = 1;
    34: op1_12_inv19 = 1;
    37: op1_12_inv19 = 1;
    38: op1_12_inv19 = 1;
    40: op1_12_inv19 = 1;
    42: op1_12_inv19 = 1;
    43: op1_12_inv19 = 1;
    47: op1_12_inv19 = 1;
    54: op1_12_inv19 = 1;
    56: op1_12_inv19 = 1;
    60: op1_12_inv19 = 1;
    61: op1_12_inv19 = 1;
    66: op1_12_inv19 = 1;
    69: op1_12_inv19 = 1;
    72: op1_12_inv19 = 1;
    74: op1_12_inv19 = 1;
    76: op1_12_inv19 = 1;
    77: op1_12_inv19 = 1;
    78: op1_12_inv19 = 1;
    81: op1_12_inv19 = 1;
    82: op1_12_inv19 = 1;
    83: op1_12_inv19 = 1;
    84: op1_12_inv19 = 1;
    85: op1_12_inv19 = 1;
    87: op1_12_inv19 = 1;
    88: op1_12_inv19 = 1;
    89: op1_12_inv19 = 1;
    92: op1_12_inv19 = 1;
    95: op1_12_inv19 = 1;
    default: op1_12_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in20 = reg_0250;
    6: op1_12_in20 = imem04_in[11:8];
    7: op1_12_in20 = reg_0164;
    8: op1_12_in20 = imem01_in[91:88];
    9: op1_12_in20 = reg_0958;
    10: op1_12_in20 = reg_0095;
    11: op1_12_in20 = reg_0712;
    12: op1_12_in20 = reg_0666;
    15: op1_12_in20 = reg_0666;
    13: op1_12_in20 = imem07_in[91:88];
    14: op1_12_in20 = imem01_in[31:28];
    16: op1_12_in20 = reg_0960;
    18: op1_12_in20 = reg_0608;
    19: op1_12_in20 = reg_0444;
    20: op1_12_in20 = reg_0134;
    21: op1_12_in20 = reg_0207;
    22: op1_12_in20 = reg_0369;
    23: op1_12_in20 = imem05_in[107:104];
    24: op1_12_in20 = imem04_in[107:104];
    25: op1_12_in20 = reg_0135;
    26: op1_12_in20 = reg_0506;
    37: op1_12_in20 = reg_0506;
    27: op1_12_in20 = reg_0168;
    28: op1_12_in20 = imem07_in[119:116];
    29: op1_12_in20 = reg_0055;
    30: op1_12_in20 = reg_0973;
    31: op1_12_in20 = reg_0190;
    32: op1_12_in20 = reg_0334;
    33: op1_12_in20 = imem03_in[15:12];
    34: op1_12_in20 = reg_0597;
    35: op1_12_in20 = reg_0213;
    36: op1_12_in20 = imem01_in[83:80];
    38: op1_12_in20 = reg_0224;
    39: op1_12_in20 = reg_0133;
    40: op1_12_in20 = reg_0150;
    41: op1_12_in20 = reg_0495;
    53: op1_12_in20 = reg_0495;
    42: op1_12_in20 = imem01_in[107:104];
    43: op1_12_in20 = reg_0317;
    44: op1_12_in20 = reg_0067;
    46: op1_12_in20 = reg_0221;
    47: op1_12_in20 = reg_0809;
    49: op1_12_in20 = reg_0905;
    50: op1_12_in20 = reg_0720;
    51: op1_12_in20 = reg_0783;
    52: op1_12_in20 = reg_1016;
    54: op1_12_in20 = reg_0143;
    56: op1_12_in20 = reg_0205;
    57: op1_12_in20 = imem01_in[79:76];
    59: op1_12_in20 = imem02_in[119:116];
    60: op1_12_in20 = imem01_in[23:20];
    61: op1_12_in20 = reg_0083;
    62: op1_12_in20 = reg_0145;
    69: op1_12_in20 = reg_0145;
    64: op1_12_in20 = reg_0176;
    66: op1_12_in20 = imem01_in[3:0];
    68: op1_12_in20 = reg_0976;
    70: op1_12_in20 = imem01_in[43:40];
    71: op1_12_in20 = reg_1000;
    72: op1_12_in20 = reg_0180;
    73: op1_12_in20 = imem01_in[111:108];
    74: op1_12_in20 = reg_0120;
    75: op1_12_in20 = reg_0007;
    76: op1_12_in20 = reg_0511;
    77: op1_12_in20 = reg_0270;
    78: op1_12_in20 = reg_0002;
    79: op1_12_in20 = reg_0805;
    80: op1_12_in20 = reg_0225;
    81: op1_12_in20 = reg_0087;
    82: op1_12_in20 = reg_0523;
    83: op1_12_in20 = reg_0022;
    84: op1_12_in20 = reg_0295;
    85: op1_12_in20 = reg_0192;
    86: op1_12_in20 = reg_0827;
    87: op1_12_in20 = reg_0017;
    88: op1_12_in20 = reg_0201;
    89: op1_12_in20 = reg_0011;
    92: op1_12_in20 = imem03_in[7:4];
    93: op1_12_in20 = reg_0048;
    94: op1_12_in20 = reg_0243;
    95: op1_12_in20 = reg_0306;
    96: op1_12_in20 = reg_0537;
    default: op1_12_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv20 = 1;
    6: op1_12_inv20 = 1;
    7: op1_12_inv20 = 1;
    8: op1_12_inv20 = 1;
    11: op1_12_inv20 = 1;
    12: op1_12_inv20 = 1;
    18: op1_12_inv20 = 1;
    19: op1_12_inv20 = 1;
    25: op1_12_inv20 = 1;
    26: op1_12_inv20 = 1;
    31: op1_12_inv20 = 1;
    32: op1_12_inv20 = 1;
    33: op1_12_inv20 = 1;
    34: op1_12_inv20 = 1;
    36: op1_12_inv20 = 1;
    37: op1_12_inv20 = 1;
    38: op1_12_inv20 = 1;
    39: op1_12_inv20 = 1;
    42: op1_12_inv20 = 1;
    47: op1_12_inv20 = 1;
    49: op1_12_inv20 = 1;
    51: op1_12_inv20 = 1;
    52: op1_12_inv20 = 1;
    57: op1_12_inv20 = 1;
    59: op1_12_inv20 = 1;
    68: op1_12_inv20 = 1;
    71: op1_12_inv20 = 1;
    73: op1_12_inv20 = 1;
    76: op1_12_inv20 = 1;
    77: op1_12_inv20 = 1;
    78: op1_12_inv20 = 1;
    79: op1_12_inv20 = 1;
    84: op1_12_inv20 = 1;
    89: op1_12_inv20 = 1;
    94: op1_12_inv20 = 1;
    default: op1_12_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in21 = reg_0251;
    6: op1_12_in21 = imem04_in[15:12];
    8: op1_12_in21 = reg_0500;
    9: op1_12_in21 = reg_0955;
    10: op1_12_in21 = reg_0052;
    11: op1_12_in21 = reg_0701;
    12: op1_12_in21 = reg_0637;
    13: op1_12_in21 = imem07_in[111:108];
    14: op1_12_in21 = imem01_in[43:40];
    15: op1_12_in21 = reg_0654;
    16: op1_12_in21 = reg_0826;
    18: op1_12_in21 = reg_0618;
    19: op1_12_in21 = reg_0435;
    20: op1_12_in21 = imem06_in[87:84];
    21: op1_12_in21 = reg_0211;
    22: op1_12_in21 = reg_0385;
    51: op1_12_in21 = reg_0385;
    23: op1_12_in21 = imem05_in[111:108];
    24: op1_12_in21 = imem04_in[111:108];
    25: op1_12_in21 = reg_0128;
    26: op1_12_in21 = reg_0840;
    27: op1_12_in21 = reg_0157;
    28: op1_12_in21 = imem07_in[123:120];
    29: op1_12_in21 = reg_0537;
    30: op1_12_in21 = reg_0971;
    31: op1_12_in21 = reg_0197;
    32: op1_12_in21 = reg_0318;
    33: op1_12_in21 = imem03_in[87:84];
    34: op1_12_in21 = reg_0595;
    35: op1_12_in21 = reg_0212;
    36: op1_12_in21 = imem01_in[95:92];
    70: op1_12_in21 = imem01_in[95:92];
    37: op1_12_in21 = imem03_in[23:20];
    38: op1_12_in21 = reg_0236;
    39: op1_12_in21 = reg_0151;
    40: op1_12_in21 = reg_0153;
    54: op1_12_in21 = reg_0153;
    41: op1_12_in21 = reg_0914;
    42: op1_12_in21 = reg_0242;
    43: op1_12_in21 = reg_0343;
    44: op1_12_in21 = reg_0064;
    46: op1_12_in21 = reg_0249;
    47: op1_12_in21 = reg_0764;
    49: op1_12_in21 = imem01_in[47:44];
    50: op1_12_in21 = reg_0729;
    52: op1_12_in21 = reg_0524;
    53: op1_12_in21 = reg_0612;
    77: op1_12_in21 = reg_0612;
    56: op1_12_in21 = reg_0202;
    57: op1_12_in21 = imem01_in[119:116];
    59: op1_12_in21 = reg_0363;
    60: op1_12_in21 = imem01_in[35:32];
    61: op1_12_in21 = reg_0089;
    62: op1_12_in21 = reg_0136;
    64: op1_12_in21 = reg_0184;
    66: op1_12_in21 = imem01_in[23:20];
    68: op1_12_in21 = imem04_in[7:4];
    69: op1_12_in21 = reg_0134;
    71: op1_12_in21 = imem04_in[59:56];
    72: op1_12_in21 = reg_0172;
    73: op1_12_in21 = reg_0969;
    74: op1_12_in21 = reg_0487;
    75: op1_12_in21 = reg_0482;
    76: op1_12_in21 = reg_0282;
    78: op1_12_in21 = reg_0428;
    79: op1_12_in21 = reg_0321;
    80: op1_12_in21 = reg_0522;
    81: op1_12_in21 = reg_0037;
    82: op1_12_in21 = reg_0748;
    83: op1_12_in21 = imem07_in[3:0];
    84: op1_12_in21 = reg_0044;
    85: op1_12_in21 = imem01_in[19:16];
    86: op1_12_in21 = reg_0101;
    87: op1_12_in21 = reg_1010;
    88: op1_12_in21 = reg_0213;
    89: op1_12_in21 = imem06_in[35:32];
    92: op1_12_in21 = reg_0033;
    93: op1_12_in21 = reg_0913;
    94: op1_12_in21 = reg_0627;
    95: op1_12_in21 = reg_0390;
    96: op1_12_in21 = reg_0909;
    default: op1_12_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv21 = 1;
    6: op1_12_inv21 = 1;
    8: op1_12_inv21 = 1;
    12: op1_12_inv21 = 1;
    14: op1_12_inv21 = 1;
    15: op1_12_inv21 = 1;
    19: op1_12_inv21 = 1;
    21: op1_12_inv21 = 1;
    22: op1_12_inv21 = 1;
    25: op1_12_inv21 = 1;
    26: op1_12_inv21 = 1;
    27: op1_12_inv21 = 1;
    30: op1_12_inv21 = 1;
    34: op1_12_inv21 = 1;
    35: op1_12_inv21 = 1;
    36: op1_12_inv21 = 1;
    38: op1_12_inv21 = 1;
    39: op1_12_inv21 = 1;
    40: op1_12_inv21 = 1;
    42: op1_12_inv21 = 1;
    43: op1_12_inv21 = 1;
    46: op1_12_inv21 = 1;
    47: op1_12_inv21 = 1;
    49: op1_12_inv21 = 1;
    51: op1_12_inv21 = 1;
    54: op1_12_inv21 = 1;
    61: op1_12_inv21 = 1;
    62: op1_12_inv21 = 1;
    64: op1_12_inv21 = 1;
    66: op1_12_inv21 = 1;
    68: op1_12_inv21 = 1;
    69: op1_12_inv21 = 1;
    70: op1_12_inv21 = 1;
    72: op1_12_inv21 = 1;
    74: op1_12_inv21 = 1;
    75: op1_12_inv21 = 1;
    76: op1_12_inv21 = 1;
    77: op1_12_inv21 = 1;
    78: op1_12_inv21 = 1;
    82: op1_12_inv21 = 1;
    84: op1_12_inv21 = 1;
    86: op1_12_inv21 = 1;
    95: op1_12_inv21 = 1;
    default: op1_12_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in22 = reg_0263;
    6: op1_12_in22 = imem04_in[43:40];
    8: op1_12_in22 = reg_0524;
    9: op1_12_in22 = reg_0967;
    10: op1_12_in22 = reg_0098;
    11: op1_12_in22 = reg_0424;
    12: op1_12_in22 = reg_0646;
    13: op1_12_in22 = reg_0722;
    14: op1_12_in22 = imem01_in[51:48];
    15: op1_12_in22 = reg_0358;
    16: op1_12_in22 = reg_0827;
    18: op1_12_in22 = reg_0623;
    19: op1_12_in22 = reg_0180;
    20: op1_12_in22 = reg_0614;
    21: op1_12_in22 = reg_0198;
    22: op1_12_in22 = reg_0398;
    23: op1_12_in22 = reg_0944;
    24: op1_12_in22 = imem04_in[115:112];
    25: op1_12_in22 = reg_0153;
    26: op1_12_in22 = reg_0310;
    27: op1_12_in22 = reg_0173;
    28: op1_12_in22 = reg_0716;
    29: op1_12_in22 = reg_0062;
    30: op1_12_in22 = reg_0955;
    31: op1_12_in22 = imem01_in[99:96];
    32: op1_12_in22 = reg_0818;
    33: op1_12_in22 = imem03_in[123:120];
    34: op1_12_in22 = imem07_in[3:0];
    35: op1_12_in22 = reg_0199;
    36: op1_12_in22 = imem01_in[123:120];
    37: op1_12_in22 = imem03_in[59:56];
    38: op1_12_in22 = reg_0248;
    39: op1_12_in22 = reg_0152;
    40: op1_12_in22 = reg_0137;
    41: op1_12_in22 = reg_0392;
    42: op1_12_in22 = reg_0240;
    43: op1_12_in22 = reg_0938;
    44: op1_12_in22 = reg_0288;
    46: op1_12_in22 = reg_0769;
    47: op1_12_in22 = reg_0444;
    49: op1_12_in22 = imem01_in[63:60];
    85: op1_12_in22 = imem01_in[63:60];
    50: op1_12_in22 = reg_0718;
    51: op1_12_in22 = reg_0387;
    52: op1_12_in22 = reg_0850;
    53: op1_12_in22 = reg_0294;
    54: op1_12_in22 = reg_0140;
    56: op1_12_in22 = reg_0206;
    57: op1_12_in22 = reg_0786;
    59: op1_12_in22 = reg_0565;
    60: op1_12_in22 = imem01_in[39:36];
    61: op1_12_in22 = reg_0261;
    62: op1_12_in22 = reg_0129;
    66: op1_12_in22 = imem01_in[35:32];
    68: op1_12_in22 = imem04_in[23:20];
    69: op1_12_in22 = imem06_in[15:12];
    70: op1_12_in22 = imem01_in[103:100];
    71: op1_12_in22 = imem04_in[95:92];
    72: op1_12_in22 = reg_0165;
    73: op1_12_in22 = reg_0246;
    74: op1_12_in22 = reg_0962;
    75: op1_12_in22 = reg_0758;
    76: op1_12_in22 = reg_0055;
    77: op1_12_in22 = reg_0018;
    78: op1_12_in22 = reg_0640;
    79: op1_12_in22 = reg_0532;
    80: op1_12_in22 = reg_0829;
    81: op1_12_in22 = reg_0091;
    82: op1_12_in22 = reg_0883;
    83: op1_12_in22 = imem07_in[23:20];
    84: op1_12_in22 = reg_0531;
    86: op1_12_in22 = reg_0115;
    87: op1_12_in22 = reg_0383;
    88: op1_12_in22 = reg_0192;
    89: op1_12_in22 = imem06_in[51:48];
    92: op1_12_in22 = reg_0976;
    93: op1_12_in22 = reg_1005;
    95: op1_12_in22 = reg_1005;
    94: op1_12_in22 = reg_0542;
    96: op1_12_in22 = reg_0848;
    default: op1_12_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv22 = 1;
    11: op1_12_inv22 = 1;
    14: op1_12_inv22 = 1;
    15: op1_12_inv22 = 1;
    16: op1_12_inv22 = 1;
    22: op1_12_inv22 = 1;
    24: op1_12_inv22 = 1;
    25: op1_12_inv22 = 1;
    26: op1_12_inv22 = 1;
    27: op1_12_inv22 = 1;
    29: op1_12_inv22 = 1;
    30: op1_12_inv22 = 1;
    31: op1_12_inv22 = 1;
    32: op1_12_inv22 = 1;
    34: op1_12_inv22 = 1;
    37: op1_12_inv22 = 1;
    40: op1_12_inv22 = 1;
    42: op1_12_inv22 = 1;
    43: op1_12_inv22 = 1;
    47: op1_12_inv22 = 1;
    49: op1_12_inv22 = 1;
    52: op1_12_inv22 = 1;
    53: op1_12_inv22 = 1;
    59: op1_12_inv22 = 1;
    60: op1_12_inv22 = 1;
    66: op1_12_inv22 = 1;
    69: op1_12_inv22 = 1;
    73: op1_12_inv22 = 1;
    74: op1_12_inv22 = 1;
    75: op1_12_inv22 = 1;
    78: op1_12_inv22 = 1;
    79: op1_12_inv22 = 1;
    80: op1_12_inv22 = 1;
    81: op1_12_inv22 = 1;
    82: op1_12_inv22 = 1;
    83: op1_12_inv22 = 1;
    87: op1_12_inv22 = 1;
    88: op1_12_inv22 = 1;
    93: op1_12_inv22 = 1;
    94: op1_12_inv22 = 1;
    96: op1_12_inv22 = 1;
    default: op1_12_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in23 = reg_0145;
    6: op1_12_in23 = imem04_in[55:52];
    8: op1_12_in23 = reg_0517;
    9: op1_12_in23 = reg_0964;
    10: op1_12_in23 = imem03_in[3:0];
    11: op1_12_in23 = reg_0432;
    12: op1_12_in23 = reg_0664;
    13: op1_12_in23 = reg_0728;
    14: op1_12_in23 = imem01_in[63:60];
    15: op1_12_in23 = reg_0359;
    16: op1_12_in23 = reg_0898;
    18: op1_12_in23 = reg_0601;
    19: op1_12_in23 = reg_0172;
    20: op1_12_in23 = reg_0633;
    21: op1_12_in23 = imem01_in[23:20];
    35: op1_12_in23 = imem01_in[23:20];
    22: op1_12_in23 = reg_0396;
    23: op1_12_in23 = reg_0955;
    24: op1_12_in23 = imem04_in[127:124];
    25: op1_12_in23 = reg_0137;
    54: op1_12_in23 = reg_0137;
    26: op1_12_in23 = reg_0484;
    27: op1_12_in23 = reg_0184;
    28: op1_12_in23 = reg_0704;
    29: op1_12_in23 = reg_0067;
    30: op1_12_in23 = reg_0957;
    31: op1_12_in23 = reg_0013;
    32: op1_12_in23 = reg_0037;
    33: op1_12_in23 = imem03_in[127:124];
    34: op1_12_in23 = imem07_in[11:8];
    36: op1_12_in23 = reg_0218;
    37: op1_12_in23 = imem03_in[87:84];
    38: op1_12_in23 = reg_0103;
    39: op1_12_in23 = reg_0134;
    40: op1_12_in23 = imem06_in[11:8];
    41: op1_12_in23 = reg_0264;
    42: op1_12_in23 = reg_0224;
    43: op1_12_in23 = reg_0322;
    44: op1_12_in23 = reg_0059;
    46: op1_12_in23 = reg_1037;
    47: op1_12_in23 = reg_0423;
    49: op1_12_in23 = imem01_in[71:68];
    50: op1_12_in23 = reg_0805;
    51: op1_12_in23 = reg_0356;
    52: op1_12_in23 = reg_0076;
    53: op1_12_in23 = reg_0382;
    56: op1_12_in23 = imem01_in[83:80];
    57: op1_12_in23 = reg_0904;
    59: op1_12_in23 = reg_0279;
    60: op1_12_in23 = imem01_in[51:48];
    61: op1_12_in23 = imem03_in[31:28];
    62: op1_12_in23 = imem06_in[31:28];
    66: op1_12_in23 = imem01_in[47:44];
    68: op1_12_in23 = imem04_in[59:56];
    69: op1_12_in23 = imem06_in[19:16];
    70: op1_12_in23 = imem01_in[107:104];
    71: op1_12_in23 = imem04_in[99:96];
    72: op1_12_in23 = reg_0169;
    73: op1_12_in23 = reg_1014;
    74: op1_12_in23 = reg_1039;
    75: op1_12_in23 = reg_0761;
    76: op1_12_in23 = reg_0931;
    77: op1_12_in23 = reg_0782;
    87: op1_12_in23 = reg_0782;
    78: op1_12_in23 = reg_0175;
    79: op1_12_in23 = reg_0868;
    80: op1_12_in23 = reg_0216;
    81: op1_12_in23 = reg_0049;
    82: op1_12_in23 = reg_0499;
    83: op1_12_in23 = imem07_in[55:52];
    84: op1_12_in23 = imem05_in[31:28];
    85: op1_12_in23 = imem01_in[91:88];
    86: op1_12_in23 = reg_0109;
    88: op1_12_in23 = imem01_in[15:12];
    89: op1_12_in23 = imem06_in[55:52];
    92: op1_12_in23 = reg_0278;
    93: op1_12_in23 = reg_0802;
    94: op1_12_in23 = reg_0070;
    95: op1_12_in23 = reg_0586;
    96: op1_12_in23 = reg_0850;
    default: op1_12_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv23 = 1;
    6: op1_12_inv23 = 1;
    9: op1_12_inv23 = 1;
    12: op1_12_inv23 = 1;
    13: op1_12_inv23 = 1;
    15: op1_12_inv23 = 1;
    16: op1_12_inv23 = 1;
    18: op1_12_inv23 = 1;
    20: op1_12_inv23 = 1;
    24: op1_12_inv23 = 1;
    25: op1_12_inv23 = 1;
    27: op1_12_inv23 = 1;
    31: op1_12_inv23 = 1;
    32: op1_12_inv23 = 1;
    33: op1_12_inv23 = 1;
    35: op1_12_inv23 = 1;
    36: op1_12_inv23 = 1;
    37: op1_12_inv23 = 1;
    38: op1_12_inv23 = 1;
    44: op1_12_inv23 = 1;
    47: op1_12_inv23 = 1;
    50: op1_12_inv23 = 1;
    51: op1_12_inv23 = 1;
    54: op1_12_inv23 = 1;
    56: op1_12_inv23 = 1;
    57: op1_12_inv23 = 1;
    60: op1_12_inv23 = 1;
    62: op1_12_inv23 = 1;
    66: op1_12_inv23 = 1;
    68: op1_12_inv23 = 1;
    69: op1_12_inv23 = 1;
    70: op1_12_inv23 = 1;
    74: op1_12_inv23 = 1;
    76: op1_12_inv23 = 1;
    77: op1_12_inv23 = 1;
    80: op1_12_inv23 = 1;
    86: op1_12_inv23 = 1;
    87: op1_12_inv23 = 1;
    88: op1_12_inv23 = 1;
    93: op1_12_inv23 = 1;
    95: op1_12_inv23 = 1;
    96: op1_12_inv23 = 1;
    default: op1_12_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in24 = reg_0133;
    6: op1_12_in24 = imem04_in[75:72];
    8: op1_12_in24 = reg_0508;
    9: op1_12_in24 = reg_0953;
    10: op1_12_in24 = imem03_in[7:4];
    11: op1_12_in24 = reg_0419;
    12: op1_12_in24 = reg_0656;
    13: op1_12_in24 = reg_0719;
    28: op1_12_in24 = reg_0719;
    14: op1_12_in24 = imem01_in[87:84];
    60: op1_12_in24 = imem01_in[87:84];
    15: op1_12_in24 = reg_0363;
    16: op1_12_in24 = reg_0254;
    18: op1_12_in24 = reg_0381;
    19: op1_12_in24 = reg_0178;
    20: op1_12_in24 = reg_0348;
    21: op1_12_in24 = imem01_in[47:44];
    22: op1_12_in24 = reg_0389;
    23: op1_12_in24 = reg_0942;
    30: op1_12_in24 = reg_0942;
    24: op1_12_in24 = reg_0061;
    25: op1_12_in24 = reg_0144;
    26: op1_12_in24 = reg_0079;
    29: op1_12_in24 = reg_0075;
    31: op1_12_in24 = reg_0218;
    32: op1_12_in24 = reg_0336;
    33: op1_12_in24 = reg_0343;
    34: op1_12_in24 = imem07_in[71:68];
    35: op1_12_in24 = imem01_in[39:36];
    88: op1_12_in24 = imem01_in[39:36];
    36: op1_12_in24 = reg_0239;
    37: op1_12_in24 = imem03_in[119:116];
    38: op1_12_in24 = reg_0102;
    39: op1_12_in24 = reg_0610;
    40: op1_12_in24 = imem06_in[59:56];
    41: op1_12_in24 = reg_0295;
    42: op1_12_in24 = reg_0555;
    43: op1_12_in24 = reg_0833;
    44: op1_12_in24 = reg_0054;
    46: op1_12_in24 = reg_0740;
    47: op1_12_in24 = reg_0445;
    49: op1_12_in24 = imem01_in[79:76];
    66: op1_12_in24 = imem01_in[79:76];
    50: op1_12_in24 = reg_0303;
    51: op1_12_in24 = reg_0344;
    52: op1_12_in24 = reg_0302;
    53: op1_12_in24 = reg_0222;
    54: op1_12_in24 = reg_0134;
    56: op1_12_in24 = imem01_in[107:104];
    57: op1_12_in24 = reg_0242;
    59: op1_12_in24 = reg_0358;
    61: op1_12_in24 = imem03_in[67:64];
    62: op1_12_in24 = imem06_in[63:60];
    68: op1_12_in24 = imem04_in[111:108];
    69: op1_12_in24 = imem06_in[43:40];
    70: op1_12_in24 = imem01_in[127:124];
    71: op1_12_in24 = imem04_in[103:100];
    73: op1_12_in24 = reg_0120;
    74: op1_12_in24 = reg_0501;
    75: op1_12_in24 = reg_0086;
    76: op1_12_in24 = reg_0313;
    77: op1_12_in24 = reg_0566;
    78: op1_12_in24 = reg_0166;
    79: op1_12_in24 = reg_0179;
    80: op1_12_in24 = reg_0737;
    81: op1_12_in24 = reg_0084;
    82: op1_12_in24 = reg_0749;
    83: op1_12_in24 = imem07_in[75:72];
    84: op1_12_in24 = imem05_in[55:52];
    85: op1_12_in24 = imem01_in[111:108];
    86: op1_12_in24 = reg_0110;
    87: op1_12_in24 = reg_0545;
    89: op1_12_in24 = imem06_in[87:84];
    92: op1_12_in24 = reg_0038;
    93: op1_12_in24 = reg_0524;
    94: op1_12_in24 = reg_0332;
    95: op1_12_in24 = reg_0016;
    96: op1_12_in24 = reg_0296;
    default: op1_12_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_12_inv24 = 1;
    11: op1_12_inv24 = 1;
    12: op1_12_inv24 = 1;
    13: op1_12_inv24 = 1;
    15: op1_12_inv24 = 1;
    16: op1_12_inv24 = 1;
    18: op1_12_inv24 = 1;
    24: op1_12_inv24 = 1;
    25: op1_12_inv24 = 1;
    29: op1_12_inv24 = 1;
    32: op1_12_inv24 = 1;
    34: op1_12_inv24 = 1;
    36: op1_12_inv24 = 1;
    41: op1_12_inv24 = 1;
    42: op1_12_inv24 = 1;
    43: op1_12_inv24 = 1;
    44: op1_12_inv24 = 1;
    46: op1_12_inv24 = 1;
    49: op1_12_inv24 = 1;
    52: op1_12_inv24 = 1;
    54: op1_12_inv24 = 1;
    60: op1_12_inv24 = 1;
    61: op1_12_inv24 = 1;
    62: op1_12_inv24 = 1;
    66: op1_12_inv24 = 1;
    69: op1_12_inv24 = 1;
    73: op1_12_inv24 = 1;
    77: op1_12_inv24 = 1;
    78: op1_12_inv24 = 1;
    80: op1_12_inv24 = 1;
    81: op1_12_inv24 = 1;
    85: op1_12_inv24 = 1;
    86: op1_12_inv24 = 1;
    88: op1_12_inv24 = 1;
    92: op1_12_inv24 = 1;
    95: op1_12_inv24 = 1;
    default: op1_12_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in25 = reg_0151;
    6: op1_12_in25 = imem04_in[107:104];
    8: op1_12_in25 = reg_0230;
    9: op1_12_in25 = reg_0256;
    10: op1_12_in25 = imem03_in[15:12];
    11: op1_12_in25 = reg_0434;
    12: op1_12_in25 = reg_0640;
    13: op1_12_in25 = reg_0730;
    14: op1_12_in25 = imem01_in[115:112];
    56: op1_12_in25 = imem01_in[115:112];
    15: op1_12_in25 = reg_0338;
    16: op1_12_in25 = reg_0255;
    18: op1_12_in25 = reg_0349;
    41: op1_12_in25 = reg_0349;
    20: op1_12_in25 = reg_0379;
    21: op1_12_in25 = imem01_in[67:64];
    35: op1_12_in25 = imem01_in[67:64];
    22: op1_12_in25 = reg_0985;
    23: op1_12_in25 = reg_0965;
    24: op1_12_in25 = reg_0763;
    25: op1_12_in25 = reg_0607;
    26: op1_12_in25 = imem03_in[3:0];
    28: op1_12_in25 = reg_0723;
    29: op1_12_in25 = reg_0064;
    30: op1_12_in25 = reg_0949;
    31: op1_12_in25 = reg_0247;
    32: op1_12_in25 = reg_0083;
    33: op1_12_in25 = reg_1019;
    34: op1_12_in25 = imem07_in[83:80];
    36: op1_12_in25 = reg_0860;
    37: op1_12_in25 = reg_1050;
    38: op1_12_in25 = imem02_in[39:36];
    39: op1_12_in25 = reg_0026;
    40: op1_12_in25 = imem06_in[79:76];
    42: op1_12_in25 = reg_0828;
    43: op1_12_in25 = reg_0369;
    44: op1_12_in25 = reg_0283;
    46: op1_12_in25 = reg_0615;
    47: op1_12_in25 = reg_0031;
    49: op1_12_in25 = imem01_in[95:92];
    50: op1_12_in25 = reg_0315;
    51: op1_12_in25 = reg_0295;
    52: op1_12_in25 = reg_0584;
    53: op1_12_in25 = reg_0894;
    54: op1_12_in25 = imem06_in[15:12];
    57: op1_12_in25 = reg_0933;
    59: op1_12_in25 = reg_0424;
    60: op1_12_in25 = imem01_in[99:96];
    61: op1_12_in25 = imem03_in[75:72];
    62: op1_12_in25 = imem06_in[99:96];
    66: op1_12_in25 = imem01_in[83:80];
    68: op1_12_in25 = reg_0282;
    69: op1_12_in25 = imem06_in[59:56];
    70: op1_12_in25 = reg_0969;
    71: op1_12_in25 = imem04_in[111:108];
    73: op1_12_in25 = reg_1024;
    74: op1_12_in25 = reg_0798;
    75: op1_12_in25 = reg_0016;
    76: op1_12_in25 = reg_0909;
    77: op1_12_in25 = imem07_in[11:8];
    79: op1_12_in25 = reg_0168;
    80: op1_12_in25 = reg_0906;
    81: op1_12_in25 = reg_0079;
    82: op1_12_in25 = reg_0663;
    83: op1_12_in25 = imem07_in[95:92];
    84: op1_12_in25 = imem05_in[63:60];
    85: op1_12_in25 = reg_0105;
    86: op1_12_in25 = imem02_in[7:4];
    87: op1_12_in25 = imem07_in[39:36];
    88: op1_12_in25 = imem01_in[43:40];
    89: op1_12_in25 = imem06_in[103:100];
    92: op1_12_in25 = reg_0051;
    93: op1_12_in25 = reg_0067;
    94: op1_12_in25 = imem05_in[3:0];
    95: op1_12_in25 = reg_0848;
    96: op1_12_in25 = reg_0732;
    default: op1_12_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv25 = 1;
    8: op1_12_inv25 = 1;
    9: op1_12_inv25 = 1;
    11: op1_12_inv25 = 1;
    12: op1_12_inv25 = 1;
    13: op1_12_inv25 = 1;
    15: op1_12_inv25 = 1;
    18: op1_12_inv25 = 1;
    25: op1_12_inv25 = 1;
    29: op1_12_inv25 = 1;
    31: op1_12_inv25 = 1;
    32: op1_12_inv25 = 1;
    36: op1_12_inv25 = 1;
    38: op1_12_inv25 = 1;
    40: op1_12_inv25 = 1;
    42: op1_12_inv25 = 1;
    46: op1_12_inv25 = 1;
    47: op1_12_inv25 = 1;
    50: op1_12_inv25 = 1;
    51: op1_12_inv25 = 1;
    52: op1_12_inv25 = 1;
    53: op1_12_inv25 = 1;
    54: op1_12_inv25 = 1;
    56: op1_12_inv25 = 1;
    57: op1_12_inv25 = 1;
    59: op1_12_inv25 = 1;
    60: op1_12_inv25 = 1;
    62: op1_12_inv25 = 1;
    71: op1_12_inv25 = 1;
    74: op1_12_inv25 = 1;
    75: op1_12_inv25 = 1;
    77: op1_12_inv25 = 1;
    85: op1_12_inv25 = 1;
    89: op1_12_inv25 = 1;
    92: op1_12_inv25 = 1;
    default: op1_12_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in26 = reg_0138;
    6: op1_12_in26 = reg_0548;
    8: op1_12_in26 = reg_0247;
    9: op1_12_in26 = reg_0241;
    41: op1_12_in26 = reg_0241;
    10: op1_12_in26 = imem03_in[39:36];
    11: op1_12_in26 = reg_0446;
    12: op1_12_in26 = reg_0665;
    13: op1_12_in26 = reg_0434;
    14: op1_12_in26 = reg_0013;
    15: op1_12_in26 = reg_0049;
    16: op1_12_in26 = reg_0132;
    18: op1_12_in26 = reg_0405;
    20: op1_12_in26 = reg_0351;
    21: op1_12_in26 = imem01_in[91:88];
    35: op1_12_in26 = imem01_in[91:88];
    22: op1_12_in26 = reg_0982;
    23: op1_12_in26 = reg_0251;
    24: op1_12_in26 = reg_0014;
    25: op1_12_in26 = reg_0613;
    26: op1_12_in26 = imem03_in[27:24];
    28: op1_12_in26 = reg_0726;
    29: op1_12_in26 = reg_0072;
    30: op1_12_in26 = reg_0965;
    31: op1_12_in26 = reg_0238;
    57: op1_12_in26 = reg_0238;
    32: op1_12_in26 = reg_0482;
    33: op1_12_in26 = reg_0322;
    34: op1_12_in26 = reg_0728;
    36: op1_12_in26 = reg_0248;
    42: op1_12_in26 = reg_0248;
    37: op1_12_in26 = reg_1008;
    38: op1_12_in26 = imem02_in[51:48];
    39: op1_12_in26 = reg_0621;
    40: op1_12_in26 = imem06_in[83:80];
    43: op1_12_in26 = reg_0509;
    44: op1_12_in26 = imem05_in[3:0];
    47: op1_12_in26 = imem05_in[3:0];
    46: op1_12_in26 = reg_0124;
    49: op1_12_in26 = imem01_in[115:112];
    50: op1_12_in26 = reg_0427;
    51: op1_12_in26 = reg_0384;
    52: op1_12_in26 = reg_0809;
    53: op1_12_in26 = reg_0594;
    54: op1_12_in26 = imem06_in[47:44];
    56: op1_12_in26 = reg_0586;
    59: op1_12_in26 = reg_0335;
    60: op1_12_in26 = reg_0933;
    61: op1_12_in26 = imem03_in[79:76];
    62: op1_12_in26 = imem06_in[119:116];
    66: op1_12_in26 = imem01_in[95:92];
    68: op1_12_in26 = reg_0888;
    69: op1_12_in26 = imem06_in[127:124];
    70: op1_12_in26 = reg_1056;
    71: op1_12_in26 = imem04_in[123:120];
    73: op1_12_in26 = reg_0793;
    74: op1_12_in26 = reg_0604;
    75: op1_12_in26 = reg_0884;
    76: op1_12_in26 = reg_0066;
    77: op1_12_in26 = imem07_in[39:36];
    79: op1_12_in26 = reg_0178;
    80: op1_12_in26 = reg_1051;
    81: op1_12_in26 = imem03_in[7:4];
    82: op1_12_in26 = reg_0453;
    83: op1_12_in26 = reg_0165;
    84: op1_12_in26 = imem05_in[75:72];
    85: op1_12_in26 = reg_0522;
    86: op1_12_in26 = imem02_in[23:20];
    87: op1_12_in26 = imem07_in[51:48];
    88: op1_12_in26 = imem01_in[79:76];
    89: op1_12_in26 = imem06_in[107:104];
    92: op1_12_in26 = reg_0820;
    93: op1_12_in26 = reg_0409;
    94: op1_12_in26 = imem05_in[11:8];
    95: op1_12_in26 = reg_0056;
    96: op1_12_in26 = reg_0061;
    default: op1_12_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_12_inv26 = 1;
    10: op1_12_inv26 = 1;
    11: op1_12_inv26 = 1;
    12: op1_12_inv26 = 1;
    16: op1_12_inv26 = 1;
    20: op1_12_inv26 = 1;
    25: op1_12_inv26 = 1;
    26: op1_12_inv26 = 1;
    34: op1_12_inv26 = 1;
    35: op1_12_inv26 = 1;
    36: op1_12_inv26 = 1;
    37: op1_12_inv26 = 1;
    41: op1_12_inv26 = 1;
    43: op1_12_inv26 = 1;
    46: op1_12_inv26 = 1;
    50: op1_12_inv26 = 1;
    51: op1_12_inv26 = 1;
    52: op1_12_inv26 = 1;
    53: op1_12_inv26 = 1;
    56: op1_12_inv26 = 1;
    57: op1_12_inv26 = 1;
    59: op1_12_inv26 = 1;
    62: op1_12_inv26 = 1;
    68: op1_12_inv26 = 1;
    69: op1_12_inv26 = 1;
    74: op1_12_inv26 = 1;
    76: op1_12_inv26 = 1;
    80: op1_12_inv26 = 1;
    84: op1_12_inv26 = 1;
    85: op1_12_inv26 = 1;
    86: op1_12_inv26 = 1;
    87: op1_12_inv26 = 1;
    88: op1_12_inv26 = 1;
    89: op1_12_inv26 = 1;
    92: op1_12_inv26 = 1;
    95: op1_12_inv26 = 1;
    default: op1_12_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in27 = imem06_in[11:8];
    6: op1_12_in27 = reg_0537;
    68: op1_12_in27 = reg_0537;
    8: op1_12_in27 = reg_0122;
    9: op1_12_in27 = reg_0257;
    10: op1_12_in27 = imem03_in[79:76];
    11: op1_12_in27 = reg_0440;
    12: op1_12_in27 = reg_0667;
    13: op1_12_in27 = reg_0444;
    14: op1_12_in27 = reg_0242;
    15: op1_12_in27 = reg_0087;
    16: op1_12_in27 = reg_0145;
    18: op1_12_in27 = reg_0313;
    20: op1_12_in27 = reg_0313;
    21: op1_12_in27 = imem01_in[107:104];
    22: op1_12_in27 = reg_0979;
    23: op1_12_in27 = reg_0260;
    24: op1_12_in27 = reg_0276;
    25: op1_12_in27 = reg_0631;
    26: op1_12_in27 = imem03_in[43:40];
    28: op1_12_in27 = reg_0717;
    29: op1_12_in27 = reg_0732;
    30: op1_12_in27 = reg_0953;
    31: op1_12_in27 = reg_0219;
    32: op1_12_in27 = reg_0089;
    33: op1_12_in27 = reg_0824;
    34: op1_12_in27 = reg_0710;
    35: op1_12_in27 = reg_0779;
    56: op1_12_in27 = reg_0779;
    36: op1_12_in27 = reg_1039;
    42: op1_12_in27 = reg_1039;
    37: op1_12_in27 = reg_0933;
    38: op1_12_in27 = imem02_in[67:64];
    39: op1_12_in27 = reg_0928;
    40: op1_12_in27 = imem06_in[103:100];
    41: op1_12_in27 = reg_0617;
    43: op1_12_in27 = reg_0807;
    44: op1_12_in27 = imem05_in[35:32];
    46: op1_12_in27 = reg_0109;
    47: op1_12_in27 = imem05_in[71:68];
    49: op1_12_in27 = reg_0522;
    50: op1_12_in27 = reg_0868;
    51: op1_12_in27 = reg_0628;
    52: op1_12_in27 = reg_0554;
    53: op1_12_in27 = reg_0241;
    54: op1_12_in27 = imem06_in[59:56];
    57: op1_12_in27 = reg_0798;
    59: op1_12_in27 = reg_0054;
    60: op1_12_in27 = reg_0919;
    61: op1_12_in27 = imem03_in[127:124];
    62: op1_12_in27 = imem06_in[123:120];
    66: op1_12_in27 = reg_0218;
    69: op1_12_in27 = reg_0344;
    70: op1_12_in27 = reg_0592;
    71: op1_12_in27 = reg_1004;
    73: op1_12_in27 = reg_0520;
    74: op1_12_in27 = reg_0520;
    75: op1_12_in27 = imem03_in[75:72];
    76: op1_12_in27 = reg_0288;
    77: op1_12_in27 = imem07_in[59:56];
    79: op1_12_in27 = reg_0176;
    80: op1_12_in27 = reg_0112;
    81: op1_12_in27 = imem03_in[27:24];
    82: op1_12_in27 = reg_0464;
    83: op1_12_in27 = reg_0721;
    84: op1_12_in27 = imem05_in[91:88];
    85: op1_12_in27 = reg_0496;
    86: op1_12_in27 = imem02_in[27:24];
    87: op1_12_in27 = imem07_in[71:68];
    88: op1_12_in27 = imem01_in[87:84];
    89: op1_12_in27 = imem06_in[111:108];
    92: op1_12_in27 = reg_0613;
    93: op1_12_in27 = reg_0856;
    94: op1_12_in27 = imem05_in[31:28];
    95: op1_12_in27 = reg_0764;
    96: op1_12_in27 = reg_0065;
    default: op1_12_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv27 = 1;
    13: op1_12_inv27 = 1;
    14: op1_12_inv27 = 1;
    15: op1_12_inv27 = 1;
    16: op1_12_inv27 = 1;
    18: op1_12_inv27 = 1;
    21: op1_12_inv27 = 1;
    22: op1_12_inv27 = 1;
    26: op1_12_inv27 = 1;
    31: op1_12_inv27 = 1;
    34: op1_12_inv27 = 1;
    35: op1_12_inv27 = 1;
    38: op1_12_inv27 = 1;
    43: op1_12_inv27 = 1;
    46: op1_12_inv27 = 1;
    47: op1_12_inv27 = 1;
    50: op1_12_inv27 = 1;
    52: op1_12_inv27 = 1;
    53: op1_12_inv27 = 1;
    54: op1_12_inv27 = 1;
    59: op1_12_inv27 = 1;
    60: op1_12_inv27 = 1;
    68: op1_12_inv27 = 1;
    69: op1_12_inv27 = 1;
    70: op1_12_inv27 = 1;
    73: op1_12_inv27 = 1;
    75: op1_12_inv27 = 1;
    76: op1_12_inv27 = 1;
    77: op1_12_inv27 = 1;
    80: op1_12_inv27 = 1;
    85: op1_12_inv27 = 1;
    86: op1_12_inv27 = 1;
    94: op1_12_inv27 = 1;
    default: op1_12_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in28 = imem06_in[19:16];
    6: op1_12_in28 = reg_0549;
    8: op1_12_in28 = reg_0103;
    9: op1_12_in28 = reg_0258;
    10: op1_12_in28 = reg_0582;
    11: op1_12_in28 = reg_0159;
    12: op1_12_in28 = reg_0341;
    13: op1_12_in28 = reg_0437;
    14: op1_12_in28 = reg_0503;
    15: op1_12_in28 = imem03_in[47:44];
    16: op1_12_in28 = reg_0152;
    18: op1_12_in28 = reg_0404;
    20: op1_12_in28 = reg_0404;
    21: op1_12_in28 = reg_0246;
    22: op1_12_in28 = reg_0986;
    23: op1_12_in28 = reg_0497;
    24: op1_12_in28 = reg_0279;
    25: op1_12_in28 = reg_0633;
    26: op1_12_in28 = reg_0602;
    28: op1_12_in28 = reg_0714;
    29: op1_12_in28 = reg_0278;
    30: op1_12_in28 = reg_1021;
    31: op1_12_in28 = reg_1042;
    88: op1_12_in28 = reg_1042;
    32: op1_12_in28 = reg_0291;
    33: op1_12_in28 = reg_0847;
    34: op1_12_in28 = reg_0709;
    35: op1_12_in28 = reg_0224;
    36: op1_12_in28 = reg_0830;
    37: op1_12_in28 = reg_0046;
    38: op1_12_in28 = imem02_in[99:96];
    39: op1_12_in28 = reg_0615;
    40: op1_12_in28 = imem06_in[115:112];
    54: op1_12_in28 = imem06_in[115:112];
    41: op1_12_in28 = reg_0605;
    42: op1_12_in28 = reg_0869;
    57: op1_12_in28 = reg_0869;
    43: op1_12_in28 = reg_1002;
    44: op1_12_in28 = imem05_in[39:36];
    46: op1_12_in28 = imem02_in[63:60];
    47: op1_12_in28 = imem05_in[103:100];
    49: op1_12_in28 = reg_0496;
    50: op1_12_in28 = reg_0174;
    51: op1_12_in28 = reg_0609;
    52: op1_12_in28 = reg_0517;
    53: op1_12_in28 = reg_0545;
    56: op1_12_in28 = reg_0928;
    59: op1_12_in28 = reg_0083;
    60: op1_12_in28 = reg_0274;
    61: op1_12_in28 = reg_0620;
    62: op1_12_in28 = reg_0696;
    66: op1_12_in28 = reg_0592;
    68: op1_12_in28 = reg_0058;
    69: op1_12_in28 = reg_1019;
    70: op1_12_in28 = reg_0793;
    71: op1_12_in28 = reg_1009;
    73: op1_12_in28 = reg_0514;
    74: op1_12_in28 = reg_0610;
    75: op1_12_in28 = imem03_in[91:88];
    76: op1_12_in28 = reg_0732;
    77: op1_12_in28 = imem07_in[67:64];
    80: op1_12_in28 = reg_0117;
    81: op1_12_in28 = imem03_in[75:72];
    82: op1_12_in28 = reg_0469;
    83: op1_12_in28 = reg_0726;
    84: op1_12_in28 = imem05_in[95:92];
    94: op1_12_in28 = imem05_in[95:92];
    85: op1_12_in28 = reg_0604;
    86: op1_12_in28 = imem02_in[55:52];
    87: op1_12_in28 = imem07_in[87:84];
    89: op1_12_in28 = imem07_in[27:24];
    92: op1_12_in28 = reg_0523;
    93: op1_12_in28 = imem05_in[63:60];
    95: op1_12_in28 = reg_0071;
    96: op1_12_in28 = reg_0494;
    default: op1_12_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv28 = 1;
    9: op1_12_inv28 = 1;
    14: op1_12_inv28 = 1;
    15: op1_12_inv28 = 1;
    16: op1_12_inv28 = 1;
    18: op1_12_inv28 = 1;
    20: op1_12_inv28 = 1;
    21: op1_12_inv28 = 1;
    24: op1_12_inv28 = 1;
    25: op1_12_inv28 = 1;
    26: op1_12_inv28 = 1;
    29: op1_12_inv28 = 1;
    32: op1_12_inv28 = 1;
    35: op1_12_inv28 = 1;
    36: op1_12_inv28 = 1;
    39: op1_12_inv28 = 1;
    40: op1_12_inv28 = 1;
    41: op1_12_inv28 = 1;
    42: op1_12_inv28 = 1;
    43: op1_12_inv28 = 1;
    46: op1_12_inv28 = 1;
    47: op1_12_inv28 = 1;
    50: op1_12_inv28 = 1;
    54: op1_12_inv28 = 1;
    56: op1_12_inv28 = 1;
    61: op1_12_inv28 = 1;
    62: op1_12_inv28 = 1;
    66: op1_12_inv28 = 1;
    69: op1_12_inv28 = 1;
    74: op1_12_inv28 = 1;
    75: op1_12_inv28 = 1;
    77: op1_12_inv28 = 1;
    80: op1_12_inv28 = 1;
    84: op1_12_inv28 = 1;
    86: op1_12_inv28 = 1;
    87: op1_12_inv28 = 1;
    88: op1_12_inv28 = 1;
    93: op1_12_inv28 = 1;
    95: op1_12_inv28 = 1;
    default: op1_12_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in29 = imem06_in[27:24];
    6: op1_12_in29 = reg_0554;
    8: op1_12_in29 = reg_0125;
    9: op1_12_in29 = reg_0253;
    10: op1_12_in29 = reg_0571;
    11: op1_12_in29 = reg_0169;
    12: op1_12_in29 = reg_0359;
    13: op1_12_in29 = reg_0420;
    14: op1_12_in29 = reg_0238;
    15: op1_12_in29 = imem03_in[79:76];
    16: op1_12_in29 = imem06_in[39:36];
    18: op1_12_in29 = reg_0406;
    20: op1_12_in29 = reg_0315;
    21: op1_12_in29 = reg_0766;
    22: op1_12_in29 = reg_0974;
    23: op1_12_in29 = reg_0148;
    24: op1_12_in29 = reg_0738;
    25: op1_12_in29 = reg_0632;
    26: op1_12_in29 = reg_0586;
    28: op1_12_in29 = reg_0702;
    29: op1_12_in29 = reg_0774;
    30: op1_12_in29 = reg_0826;
    31: op1_12_in29 = reg_0230;
    32: op1_12_in29 = imem03_in[3:0];
    33: op1_12_in29 = reg_0509;
    34: op1_12_in29 = reg_0711;
    35: op1_12_in29 = reg_0828;
    36: op1_12_in29 = reg_0871;
    60: op1_12_in29 = reg_0871;
    37: op1_12_in29 = reg_0346;
    38: op1_12_in29 = imem02_in[103:100];
    39: op1_12_in29 = imem06_in[31:28];
    40: op1_12_in29 = imem06_in[119:116];
    41: op1_12_in29 = reg_0609;
    42: op1_12_in29 = reg_0829;
    43: op1_12_in29 = reg_0984;
    44: op1_12_in29 = imem05_in[123:120];
    46: op1_12_in29 = imem02_in[87:84];
    47: op1_12_in29 = reg_0962;
    49: op1_12_in29 = reg_0520;
    50: op1_12_in29 = reg_0167;
    51: op1_12_in29 = reg_1010;
    52: op1_12_in29 = reg_0429;
    53: op1_12_in29 = imem07_in[27:24];
    54: op1_12_in29 = reg_0534;
    56: op1_12_in29 = reg_0870;
    57: op1_12_in29 = reg_0514;
    70: op1_12_in29 = reg_0514;
    59: op1_12_in29 = reg_0482;
    61: op1_12_in29 = reg_0572;
    62: op1_12_in29 = reg_0393;
    66: op1_12_in29 = reg_1045;
    68: op1_12_in29 = reg_0517;
    96: op1_12_in29 = reg_0517;
    69: op1_12_in29 = reg_0229;
    71: op1_12_in29 = reg_0888;
    73: op1_12_in29 = reg_0830;
    74: op1_12_in29 = reg_0304;
    75: op1_12_in29 = reg_0099;
    76: op1_12_in29 = reg_0764;
    77: op1_12_in29 = imem07_in[83:80];
    80: op1_12_in29 = imem02_in[47:44];
    81: op1_12_in29 = imem03_in[95:92];
    82: op1_12_in29 = reg_0481;
    83: op1_12_in29 = reg_0717;
    84: op1_12_in29 = reg_0655;
    85: op1_12_in29 = reg_1037;
    86: op1_12_in29 = imem02_in[67:64];
    87: op1_12_in29 = imem07_in[99:96];
    88: op1_12_in29 = reg_0225;
    89: op1_12_in29 = imem07_in[79:76];
    92: op1_12_in29 = reg_0050;
    93: op1_12_in29 = imem05_in[107:104];
    94: op1_12_in29 = imem05_in[119:116];
    95: op1_12_in29 = reg_0777;
    default: op1_12_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv29 = 1;
    6: op1_12_inv29 = 1;
    9: op1_12_inv29 = 1;
    10: op1_12_inv29 = 1;
    11: op1_12_inv29 = 1;
    14: op1_12_inv29 = 1;
    16: op1_12_inv29 = 1;
    18: op1_12_inv29 = 1;
    21: op1_12_inv29 = 1;
    22: op1_12_inv29 = 1;
    24: op1_12_inv29 = 1;
    25: op1_12_inv29 = 1;
    26: op1_12_inv29 = 1;
    31: op1_12_inv29 = 1;
    32: op1_12_inv29 = 1;
    34: op1_12_inv29 = 1;
    36: op1_12_inv29 = 1;
    37: op1_12_inv29 = 1;
    38: op1_12_inv29 = 1;
    39: op1_12_inv29 = 1;
    40: op1_12_inv29 = 1;
    42: op1_12_inv29 = 1;
    44: op1_12_inv29 = 1;
    47: op1_12_inv29 = 1;
    49: op1_12_inv29 = 1;
    50: op1_12_inv29 = 1;
    53: op1_12_inv29 = 1;
    56: op1_12_inv29 = 1;
    57: op1_12_inv29 = 1;
    61: op1_12_inv29 = 1;
    62: op1_12_inv29 = 1;
    66: op1_12_inv29 = 1;
    70: op1_12_inv29 = 1;
    74: op1_12_inv29 = 1;
    76: op1_12_inv29 = 1;
    77: op1_12_inv29 = 1;
    81: op1_12_inv29 = 1;
    82: op1_12_inv29 = 1;
    84: op1_12_inv29 = 1;
    85: op1_12_inv29 = 1;
    86: op1_12_inv29 = 1;
    87: op1_12_inv29 = 1;
    89: op1_12_inv29 = 1;
    93: op1_12_inv29 = 1;
    95: op1_12_inv29 = 1;
    default: op1_12_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_12_in30 = imem06_in[55:52];
    6: op1_12_in30 = reg_0540;
    8: op1_12_in30 = reg_0101;
    9: op1_12_in30 = reg_0136;
    10: op1_12_in30 = reg_0573;
    11: op1_12_in30 = reg_0185;
    12: op1_12_in30 = reg_0328;
    13: op1_12_in30 = imem07_in[23:20];
    14: op1_12_in30 = reg_0507;
    15: op1_12_in30 = imem03_in[127:124];
    16: op1_12_in30 = imem06_in[95:92];
    18: op1_12_in30 = reg_0799;
    20: op1_12_in30 = imem07_in[55:52];
    21: op1_12_in30 = reg_0247;
    22: op1_12_in30 = reg_0977;
    23: op1_12_in30 = reg_0133;
    24: op1_12_in30 = reg_0774;
    25: op1_12_in30 = reg_0622;
    51: op1_12_in30 = reg_0622;
    26: op1_12_in30 = reg_0599;
    28: op1_12_in30 = reg_0729;
    29: op1_12_in30 = reg_0855;
    30: op1_12_in30 = reg_0835;
    31: op1_12_in30 = reg_0500;
    32: op1_12_in30 = imem03_in[23:20];
    33: op1_12_in30 = reg_0836;
    34: op1_12_in30 = reg_0706;
    35: op1_12_in30 = reg_0221;
    36: op1_12_in30 = reg_1017;
    37: op1_12_in30 = reg_0389;
    38: op1_12_in30 = imem02_in[107:104];
    39: op1_12_in30 = imem06_in[47:44];
    40: op1_12_in30 = imem06_in[123:120];
    41: op1_12_in30 = reg_0545;
    42: op1_12_in30 = reg_0216;
    43: op1_12_in30 = reg_0997;
    44: op1_12_in30 = reg_0962;
    46: op1_12_in30 = reg_0642;
    47: op1_12_in30 = reg_0954;
    49: op1_12_in30 = reg_1043;
    88: op1_12_in30 = reg_1043;
    52: op1_12_in30 = reg_0041;
    76: op1_12_in30 = reg_0041;
    53: op1_12_in30 = imem07_in[91:88];
    54: op1_12_in30 = reg_0895;
    56: op1_12_in30 = reg_0592;
    57: op1_12_in30 = reg_0830;
    59: op1_12_in30 = reg_0088;
    60: op1_12_in30 = reg_0253;
    61: op1_12_in30 = reg_0580;
    62: op1_12_in30 = reg_0626;
    66: op1_12_in30 = reg_0238;
    68: op1_12_in30 = reg_0332;
    95: op1_12_in30 = reg_0332;
    69: op1_12_in30 = reg_0395;
    70: op1_12_in30 = reg_0354;
    71: op1_12_in30 = reg_0778;
    73: op1_12_in30 = reg_1055;
    74: op1_12_in30 = reg_0003;
    75: op1_12_in30 = reg_0111;
    77: op1_12_in30 = reg_0710;
    80: op1_12_in30 = imem02_in[111:108];
    81: op1_12_in30 = imem03_in[119:116];
    82: op1_12_in30 = reg_0474;
    83: op1_12_in30 = reg_0715;
    84: op1_12_in30 = reg_0140;
    85: op1_12_in30 = reg_0227;
    86: op1_12_in30 = imem02_in[91:88];
    87: op1_12_in30 = imem07_in[119:116];
    89: op1_12_in30 = imem07_in[107:104];
    92: op1_12_in30 = reg_0986;
    93: op1_12_in30 = reg_0636;
    94: op1_12_in30 = reg_0217;
    96: op1_12_in30 = reg_0777;
    default: op1_12_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    11: op1_12_inv30 = 1;
    14: op1_12_inv30 = 1;
    16: op1_12_inv30 = 1;
    20: op1_12_inv30 = 1;
    21: op1_12_inv30 = 1;
    25: op1_12_inv30 = 1;
    26: op1_12_inv30 = 1;
    28: op1_12_inv30 = 1;
    30: op1_12_inv30 = 1;
    31: op1_12_inv30 = 1;
    32: op1_12_inv30 = 1;
    33: op1_12_inv30 = 1;
    34: op1_12_inv30 = 1;
    36: op1_12_inv30 = 1;
    37: op1_12_inv30 = 1;
    38: op1_12_inv30 = 1;
    41: op1_12_inv30 = 1;
    44: op1_12_inv30 = 1;
    47: op1_12_inv30 = 1;
    52: op1_12_inv30 = 1;
    53: op1_12_inv30 = 1;
    54: op1_12_inv30 = 1;
    56: op1_12_inv30 = 1;
    57: op1_12_inv30 = 1;
    62: op1_12_inv30 = 1;
    66: op1_12_inv30 = 1;
    68: op1_12_inv30 = 1;
    69: op1_12_inv30 = 1;
    70: op1_12_inv30 = 1;
    73: op1_12_inv30 = 1;
    74: op1_12_inv30 = 1;
    75: op1_12_inv30 = 1;
    76: op1_12_inv30 = 1;
    77: op1_12_inv30 = 1;
    80: op1_12_inv30 = 1;
    83: op1_12_inv30 = 1;
    84: op1_12_inv30 = 1;
    85: op1_12_inv30 = 1;
    86: op1_12_inv30 = 1;
    88: op1_12_inv30 = 1;
    92: op1_12_inv30 = 1;
    default: op1_12_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_12_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_12_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in00 = imem06_in[59:56];
    6: op1_13_in00 = reg_0541;
    71: op1_13_in00 = reg_0541;
    7: op1_13_in00 = imem00_in[15:12];
    8: op1_13_in00 = reg_0109;
    9: op1_13_in00 = reg_0146;
    10: op1_13_in00 = reg_0572;
    11: op1_13_in00 = imem00_in[3:0];
    45: op1_13_in00 = imem00_in[3:0];
    12: op1_13_in00 = reg_0045;
    13: op1_13_in00 = imem00_in[47:44];
    28: op1_13_in00 = imem00_in[47:44];
    14: op1_13_in00 = reg_0249;
    66: op1_13_in00 = reg_0249;
    15: op1_13_in00 = reg_0598;
    16: op1_13_in00 = imem06_in[103:100];
    17: op1_13_in00 = imem00_in[55:52];
    18: op1_13_in00 = reg_0800;
    19: op1_13_in00 = imem00_in[75:72];
    20: op1_13_in00 = imem07_in[83:80];
    21: op1_13_in00 = reg_0230;
    22: op1_13_in00 = reg_0282;
    23: op1_13_in00 = reg_0150;
    24: op1_13_in00 = imem05_in[39:36];
    25: op1_13_in00 = reg_0348;
    26: op1_13_in00 = reg_0579;
    4: op1_13_in00 = imem07_in[91:88];
    27: op1_13_in00 = imem00_in[23:20];
    50: op1_13_in00 = imem00_in[23:20];
    65: op1_13_in00 = imem00_in[23:20];
    90: op1_13_in00 = imem00_in[23:20];
    3: op1_13_in00 = imem07_in[19:16];
    29: op1_13_in00 = reg_0773;
    30: op1_13_in00 = reg_0900;
    31: op1_13_in00 = reg_1036;
    32: op1_13_in00 = imem03_in[67:64];
    2: op1_13_in00 = imem07_in[43:40];
    33: op1_13_in00 = reg_0312;
    34: op1_13_in00 = imem00_in[63:60];
    35: op1_13_in00 = reg_0219;
    36: op1_13_in00 = reg_1018;
    37: op1_13_in00 = reg_0923;
    38: op1_13_in00 = reg_0661;
    39: op1_13_in00 = imem06_in[51:48];
    40: op1_13_in00 = reg_0614;
    41: op1_13_in00 = imem07_in[3:0];
    42: op1_13_in00 = reg_0354;
    43: op1_13_in00 = imem04_in[11:8];
    44: op1_13_in00 = reg_0957;
    46: op1_13_in00 = reg_0654;
    47: op1_13_in00 = reg_0965;
    48: op1_13_in00 = imem00_in[59:56];
    49: op1_13_in00 = reg_1031;
    51: op1_13_in00 = imem07_in[7:4];
    52: op1_13_in00 = imem05_in[3:0];
    53: op1_13_in00 = imem07_in[99:96];
    54: op1_13_in00 = reg_0220;
    55: op1_13_in00 = reg_0897;
    56: op1_13_in00 = reg_0503;
    57: op1_13_in00 = reg_1037;
    58: op1_13_in00 = imem00_in[7:4];
    67: op1_13_in00 = imem00_in[7:4];
    79: op1_13_in00 = imem00_in[7:4];
    59: op1_13_in00 = reg_0090;
    60: op1_13_in00 = reg_0522;
    61: op1_13_in00 = reg_0245;
    62: op1_13_in00 = reg_0679;
    63: op1_13_in00 = imem00_in[39:36];
    64: op1_13_in00 = imem00_in[27:24];
    68: op1_13_in00 = reg_0531;
    69: op1_13_in00 = reg_0617;
    70: op1_13_in00 = reg_0610;
    72: op1_13_in00 = imem00_in[19:16];
    73: op1_13_in00 = reg_1033;
    74: op1_13_in00 = reg_0555;
    75: op1_13_in00 = reg_1007;
    76: op1_13_in00 = reg_0065;
    77: op1_13_in00 = reg_0715;
    78: op1_13_in00 = imem00_in[35:32];
    80: op1_13_in00 = imem02_in[123:120];
    81: op1_13_in00 = reg_0434;
    82: op1_13_in00 = reg_0459;
    83: op1_13_in00 = reg_0718;
    84: op1_13_in00 = reg_0958;
    85: op1_13_in00 = reg_0521;
    86: op1_13_in00 = imem02_in[107:104];
    87: op1_13_in00 = reg_0708;
    88: op1_13_in00 = reg_1040;
    89: op1_13_in00 = imem07_in[115:112];
    91: op1_13_in00 = reg_0187;
    92: op1_13_in00 = reg_0988;
    93: op1_13_in00 = reg_0319;
    94: op1_13_in00 = reg_0128;
    95: op1_13_in00 = imem05_in[23:20];
    96: op1_13_in00 = reg_0542;
    default: op1_13_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv00 = 1;
    8: op1_13_inv00 = 1;
    9: op1_13_inv00 = 1;
    13: op1_13_inv00 = 1;
    14: op1_13_inv00 = 1;
    16: op1_13_inv00 = 1;
    17: op1_13_inv00 = 1;
    18: op1_13_inv00 = 1;
    21: op1_13_inv00 = 1;
    22: op1_13_inv00 = 1;
    25: op1_13_inv00 = 1;
    4: op1_13_inv00 = 1;
    29: op1_13_inv00 = 1;
    31: op1_13_inv00 = 1;
    32: op1_13_inv00 = 1;
    2: op1_13_inv00 = 1;
    33: op1_13_inv00 = 1;
    34: op1_13_inv00 = 1;
    35: op1_13_inv00 = 1;
    37: op1_13_inv00 = 1;
    39: op1_13_inv00 = 1;
    41: op1_13_inv00 = 1;
    43: op1_13_inv00 = 1;
    44: op1_13_inv00 = 1;
    45: op1_13_inv00 = 1;
    47: op1_13_inv00 = 1;
    49: op1_13_inv00 = 1;
    50: op1_13_inv00 = 1;
    51: op1_13_inv00 = 1;
    52: op1_13_inv00 = 1;
    53: op1_13_inv00 = 1;
    54: op1_13_inv00 = 1;
    56: op1_13_inv00 = 1;
    57: op1_13_inv00 = 1;
    61: op1_13_inv00 = 1;
    62: op1_13_inv00 = 1;
    63: op1_13_inv00 = 1;
    64: op1_13_inv00 = 1;
    65: op1_13_inv00 = 1;
    66: op1_13_inv00 = 1;
    67: op1_13_inv00 = 1;
    68: op1_13_inv00 = 1;
    72: op1_13_inv00 = 1;
    73: op1_13_inv00 = 1;
    75: op1_13_inv00 = 1;
    77: op1_13_inv00 = 1;
    78: op1_13_inv00 = 1;
    80: op1_13_inv00 = 1;
    81: op1_13_inv00 = 1;
    82: op1_13_inv00 = 1;
    85: op1_13_inv00 = 1;
    87: op1_13_inv00 = 1;
    89: op1_13_inv00 = 1;
    90: op1_13_inv00 = 1;
    91: op1_13_inv00 = 1;
    94: op1_13_inv00 = 1;
    96: op1_13_inv00 = 1;
    default: op1_13_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in01 = imem06_in[83:80];
    6: op1_13_in01 = reg_0281;
    7: op1_13_in01 = imem00_in[55:52];
    8: op1_13_in01 = reg_0107;
    84: op1_13_in01 = reg_0107;
    9: op1_13_in01 = reg_0143;
    10: op1_13_in01 = reg_0395;
    11: op1_13_in01 = imem00_in[23:20];
    12: op1_13_in01 = reg_0089;
    13: op1_13_in01 = imem00_in[79:76];
    14: op1_13_in01 = reg_0230;
    15: op1_13_in01 = reg_0572;
    16: op1_13_in01 = reg_0620;
    17: op1_13_in01 = imem00_in[103:100];
    18: op1_13_in01 = reg_0005;
    19: op1_13_in01 = imem00_in[115:112];
    20: op1_13_in01 = reg_0726;
    21: op1_13_in01 = reg_0885;
    22: op1_13_in01 = reg_0048;
    23: op1_13_in01 = reg_0152;
    24: op1_13_in01 = imem05_in[59:56];
    25: op1_13_in01 = reg_0372;
    26: op1_13_in01 = reg_0568;
    4: op1_13_in01 = imem07_in[111:108];
    27: op1_13_in01 = imem00_in[63:60];
    63: op1_13_in01 = imem00_in[63:60];
    28: op1_13_in01 = imem00_in[95:92];
    3: op1_13_in01 = imem07_in[23:20];
    29: op1_13_in01 = imem05_in[19:16];
    30: op1_13_in01 = reg_0832;
    31: op1_13_in01 = reg_0122;
    32: op1_13_in01 = reg_0573;
    33: op1_13_in01 = reg_0993;
    34: op1_13_in01 = imem00_in[107:104];
    35: op1_13_in01 = reg_0905;
    36: op1_13_in01 = reg_0123;
    37: op1_13_in01 = reg_0373;
    38: op1_13_in01 = reg_0651;
    39: op1_13_in01 = imem06_in[59:56];
    40: op1_13_in01 = reg_0533;
    41: op1_13_in01 = imem07_in[39:36];
    51: op1_13_in01 = imem07_in[39:36];
    42: op1_13_in01 = reg_1017;
    43: op1_13_in01 = imem04_in[39:36];
    92: op1_13_in01 = imem04_in[39:36];
    44: op1_13_in01 = reg_0964;
    45: op1_13_in01 = imem00_in[15:12];
    46: op1_13_in01 = reg_0649;
    47: op1_13_in01 = reg_0943;
    48: op1_13_in01 = reg_0685;
    49: op1_13_in01 = reg_0737;
    88: op1_13_in01 = reg_0737;
    50: op1_13_in01 = imem00_in[47:44];
    65: op1_13_in01 = imem00_in[47:44];
    52: op1_13_in01 = imem05_in[15:12];
    53: op1_13_in01 = imem07_in[127:124];
    89: op1_13_in01 = imem07_in[127:124];
    54: op1_13_in01 = reg_0407;
    55: op1_13_in01 = reg_0375;
    56: op1_13_in01 = reg_0236;
    57: op1_13_in01 = reg_0521;
    58: op1_13_in01 = imem00_in[59:56];
    59: op1_13_in01 = reg_0840;
    60: op1_13_in01 = reg_0829;
    61: op1_13_in01 = reg_0434;
    62: op1_13_in01 = reg_0384;
    64: op1_13_in01 = imem00_in[39:36];
    66: op1_13_in01 = reg_0607;
    67: op1_13_in01 = imem00_in[27:24];
    68: op1_13_in01 = reg_0252;
    69: op1_13_in01 = reg_0619;
    70: op1_13_in01 = reg_1051;
    71: op1_13_in01 = reg_0802;
    72: op1_13_in01 = imem00_in[35:32];
    73: op1_13_in01 = reg_0114;
    74: op1_13_in01 = reg_0114;
    75: op1_13_in01 = reg_0580;
    76: op1_13_in01 = reg_0409;
    77: op1_13_in01 = reg_0563;
    78: op1_13_in01 = imem00_in[75:72];
    79: op1_13_in01 = imem00_in[11:8];
    80: op1_13_in01 = reg_0750;
    81: op1_13_in01 = reg_0298;
    82: op1_13_in01 = reg_0452;
    83: op1_13_in01 = reg_0299;
    85: op1_13_in01 = reg_1041;
    86: op1_13_in01 = reg_0334;
    87: op1_13_in01 = reg_0653;
    90: op1_13_in01 = imem00_in[51:48];
    91: op1_13_in01 = reg_0506;
    93: op1_13_in01 = reg_0057;
    94: op1_13_in01 = reg_0257;
    95: op1_13_in01 = imem05_in[31:28];
    96: op1_13_in01 = imem05_in[3:0];
    default: op1_13_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv01 = 1;
    9: op1_13_inv01 = 1;
    11: op1_13_inv01 = 1;
    12: op1_13_inv01 = 1;
    16: op1_13_inv01 = 1;
    19: op1_13_inv01 = 1;
    21: op1_13_inv01 = 1;
    23: op1_13_inv01 = 1;
    25: op1_13_inv01 = 1;
    27: op1_13_inv01 = 1;
    28: op1_13_inv01 = 1;
    3: op1_13_inv01 = 1;
    29: op1_13_inv01 = 1;
    30: op1_13_inv01 = 1;
    31: op1_13_inv01 = 1;
    33: op1_13_inv01 = 1;
    34: op1_13_inv01 = 1;
    37: op1_13_inv01 = 1;
    39: op1_13_inv01 = 1;
    41: op1_13_inv01 = 1;
    42: op1_13_inv01 = 1;
    43: op1_13_inv01 = 1;
    47: op1_13_inv01 = 1;
    49: op1_13_inv01 = 1;
    50: op1_13_inv01 = 1;
    53: op1_13_inv01 = 1;
    54: op1_13_inv01 = 1;
    55: op1_13_inv01 = 1;
    59: op1_13_inv01 = 1;
    63: op1_13_inv01 = 1;
    67: op1_13_inv01 = 1;
    71: op1_13_inv01 = 1;
    74: op1_13_inv01 = 1;
    82: op1_13_inv01 = 1;
    83: op1_13_inv01 = 1;
    85: op1_13_inv01 = 1;
    86: op1_13_inv01 = 1;
    87: op1_13_inv01 = 1;
    89: op1_13_inv01 = 1;
    90: op1_13_inv01 = 1;
    91: op1_13_inv01 = 1;
    95: op1_13_inv01 = 1;
    96: op1_13_inv01 = 1;
    default: op1_13_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in02 = imem06_in[95:92];
    6: op1_13_in02 = reg_0294;
    7: op1_13_in02 = imem00_in[79:76];
    8: op1_13_in02 = reg_0126;
    9: op1_13_in02 = reg_0153;
    10: op1_13_in02 = reg_0387;
    11: op1_13_in02 = imem00_in[35:32];
    12: op1_13_in02 = reg_0073;
    13: op1_13_in02 = imem00_in[83:80];
    78: op1_13_in02 = imem00_in[83:80];
    14: op1_13_in02 = reg_1044;
    15: op1_13_in02 = reg_0597;
    16: op1_13_in02 = reg_0621;
    17: op1_13_in02 = reg_0695;
    18: op1_13_in02 = reg_0011;
    19: op1_13_in02 = reg_0684;
    48: op1_13_in02 = reg_0684;
    20: op1_13_in02 = reg_0717;
    21: op1_13_in02 = reg_1043;
    22: op1_13_in02 = reg_0292;
    23: op1_13_in02 = reg_0143;
    24: op1_13_in02 = imem05_in[63:60];
    25: op1_13_in02 = reg_0349;
    26: op1_13_in02 = reg_0578;
    4: op1_13_in02 = reg_0425;
    27: op1_13_in02 = imem00_in[71:68];
    50: op1_13_in02 = imem00_in[71:68];
    63: op1_13_in02 = imem00_in[71:68];
    28: op1_13_in02 = imem00_in[127:124];
    3: op1_13_in02 = imem07_in[59:56];
    29: op1_13_in02 = imem05_in[27:24];
    30: op1_13_in02 = reg_0148;
    31: op1_13_in02 = reg_0125;
    32: op1_13_in02 = reg_0492;
    33: op1_13_in02 = reg_0978;
    34: op1_13_in02 = reg_0690;
    35: op1_13_in02 = reg_0869;
    36: op1_13_in02 = reg_0105;
    37: op1_13_in02 = reg_0513;
    38: op1_13_in02 = reg_0638;
    39: op1_13_in02 = imem06_in[91:88];
    40: op1_13_in02 = reg_0856;
    41: op1_13_in02 = imem07_in[87:84];
    42: op1_13_in02 = reg_0099;
    43: op1_13_in02 = imem04_in[55:52];
    44: op1_13_in02 = reg_0943;
    45: op1_13_in02 = reg_0672;
    46: op1_13_in02 = reg_0647;
    47: op1_13_in02 = reg_0900;
    49: op1_13_in02 = reg_0111;
    51: op1_13_in02 = imem07_in[67:64];
    52: op1_13_in02 = imem05_in[43:40];
    53: op1_13_in02 = reg_0727;
    54: op1_13_in02 = reg_0020;
    55: op1_13_in02 = imem00_in[15:12];
    79: op1_13_in02 = imem00_in[15:12];
    56: op1_13_in02 = reg_0274;
    57: op1_13_in02 = reg_0740;
    58: op1_13_in02 = imem00_in[67:64];
    72: op1_13_in02 = imem00_in[67:64];
    59: op1_13_in02 = reg_0484;
    60: op1_13_in02 = reg_0830;
    61: op1_13_in02 = reg_0923;
    62: op1_13_in02 = reg_0439;
    64: op1_13_in02 = imem00_in[43:40];
    65: op1_13_in02 = reg_0825;
    66: op1_13_in02 = reg_0798;
    67: op1_13_in02 = imem00_in[59:56];
    68: op1_13_in02 = reg_0281;
    69: op1_13_in02 = reg_0946;
    70: op1_13_in02 = reg_0769;
    71: op1_13_in02 = reg_0276;
    73: op1_13_in02 = reg_0113;
    74: op1_13_in02 = reg_0113;
    75: op1_13_in02 = reg_0322;
    76: op1_13_in02 = reg_0108;
    77: op1_13_in02 = reg_0123;
    80: op1_13_in02 = reg_0810;
    81: op1_13_in02 = reg_0823;
    82: op1_13_in02 = reg_0208;
    83: op1_13_in02 = reg_0047;
    84: op1_13_in02 = reg_0223;
    85: op1_13_in02 = reg_0283;
    86: op1_13_in02 = reg_0285;
    87: op1_13_in02 = reg_0744;
    88: op1_13_in02 = reg_0354;
    89: op1_13_in02 = reg_0221;
    90: op1_13_in02 = imem00_in[91:88];
    91: op1_13_in02 = reg_0324;
    92: op1_13_in02 = imem04_in[67:64];
    93: op1_13_in02 = reg_0063;
    94: op1_13_in02 = reg_0831;
    95: op1_13_in02 = imem05_in[67:64];
    96: op1_13_in02 = imem05_in[71:68];
    default: op1_13_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv02 = 1;
    9: op1_13_inv02 = 1;
    11: op1_13_inv02 = 1;
    19: op1_13_inv02 = 1;
    20: op1_13_inv02 = 1;
    22: op1_13_inv02 = 1;
    24: op1_13_inv02 = 1;
    27: op1_13_inv02 = 1;
    28: op1_13_inv02 = 1;
    3: op1_13_inv02 = 1;
    29: op1_13_inv02 = 1;
    30: op1_13_inv02 = 1;
    31: op1_13_inv02 = 1;
    35: op1_13_inv02 = 1;
    36: op1_13_inv02 = 1;
    38: op1_13_inv02 = 1;
    40: op1_13_inv02 = 1;
    42: op1_13_inv02 = 1;
    44: op1_13_inv02 = 1;
    45: op1_13_inv02 = 1;
    46: op1_13_inv02 = 1;
    48: op1_13_inv02 = 1;
    49: op1_13_inv02 = 1;
    54: op1_13_inv02 = 1;
    55: op1_13_inv02 = 1;
    56: op1_13_inv02 = 1;
    59: op1_13_inv02 = 1;
    60: op1_13_inv02 = 1;
    61: op1_13_inv02 = 1;
    62: op1_13_inv02 = 1;
    64: op1_13_inv02 = 1;
    66: op1_13_inv02 = 1;
    67: op1_13_inv02 = 1;
    68: op1_13_inv02 = 1;
    69: op1_13_inv02 = 1;
    73: op1_13_inv02 = 1;
    76: op1_13_inv02 = 1;
    80: op1_13_inv02 = 1;
    83: op1_13_inv02 = 1;
    84: op1_13_inv02 = 1;
    87: op1_13_inv02 = 1;
    89: op1_13_inv02 = 1;
    92: op1_13_inv02 = 1;
    93: op1_13_inv02 = 1;
    95: op1_13_inv02 = 1;
    96: op1_13_inv02 = 1;
    default: op1_13_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in03 = imem06_in[111:108];
    6: op1_13_in03 = reg_0277;
    7: op1_13_in03 = reg_0670;
    8: op1_13_in03 = imem02_in[7:4];
    9: op1_13_in03 = reg_0141;
    10: op1_13_in03 = reg_0312;
    11: op1_13_in03 = imem00_in[47:44];
    12: op1_13_in03 = imem03_in[3:0];
    13: op1_13_in03 = imem00_in[95:92];
    14: op1_13_in03 = reg_1040;
    15: op1_13_in03 = reg_0360;
    16: op1_13_in03 = reg_0619;
    17: op1_13_in03 = reg_0696;
    18: op1_13_in03 = imem07_in[3:0];
    19: op1_13_in03 = reg_0679;
    20: op1_13_in03 = reg_0714;
    21: op1_13_in03 = reg_1045;
    22: op1_13_in03 = reg_0537;
    23: op1_13_in03 = imem06_in[7:4];
    24: op1_13_in03 = imem05_in[87:84];
    25: op1_13_in03 = reg_0383;
    26: op1_13_in03 = reg_0590;
    4: op1_13_in03 = reg_0424;
    27: op1_13_in03 = imem00_in[79:76];
    63: op1_13_in03 = imem00_in[79:76];
    67: op1_13_in03 = imem00_in[79:76];
    28: op1_13_in03 = reg_0693;
    3: op1_13_in03 = imem07_in[83:80];
    29: op1_13_in03 = imem05_in[75:72];
    30: op1_13_in03 = reg_0139;
    31: op1_13_in03 = reg_0112;
    32: op1_13_in03 = reg_0343;
    33: op1_13_in03 = reg_0999;
    34: op1_13_in03 = reg_0451;
    35: op1_13_in03 = reg_1033;
    36: op1_13_in03 = reg_0124;
    37: op1_13_in03 = reg_0982;
    38: op1_13_in03 = reg_0662;
    39: op1_13_in03 = imem06_in[99:96];
    40: op1_13_in03 = reg_0577;
    41: op1_13_in03 = imem07_in[95:92];
    42: op1_13_in03 = reg_0115;
    43: op1_13_in03 = imem04_in[123:120];
    44: op1_13_in03 = reg_0972;
    45: op1_13_in03 = reg_0677;
    46: op1_13_in03 = reg_0082;
    47: op1_13_in03 = reg_0229;
    48: op1_13_in03 = reg_0686;
    49: op1_13_in03 = reg_0104;
    91: op1_13_in03 = reg_0104;
    50: op1_13_in03 = reg_0683;
    51: op1_13_in03 = imem07_in[99:96];
    52: op1_13_in03 = imem05_in[47:44];
    53: op1_13_in03 = reg_0361;
    54: op1_13_in03 = reg_0371;
    55: op1_13_in03 = imem00_in[87:84];
    56: op1_13_in03 = reg_0522;
    57: op1_13_in03 = reg_0832;
    88: op1_13_in03 = reg_0832;
    58: op1_13_in03 = imem00_in[71:68];
    72: op1_13_in03 = imem00_in[71:68];
    79: op1_13_in03 = imem00_in[71:68];
    59: op1_13_in03 = reg_0872;
    60: op1_13_in03 = reg_0232;
    61: op1_13_in03 = reg_0038;
    62: op1_13_in03 = reg_0863;
    64: op1_13_in03 = imem00_in[55:52];
    65: op1_13_in03 = reg_0843;
    66: op1_13_in03 = reg_0869;
    68: op1_13_in03 = reg_0435;
    69: op1_13_in03 = reg_0241;
    70: op1_13_in03 = reg_0003;
    71: op1_13_in03 = reg_0584;
    73: op1_13_in03 = reg_0821;
    74: op1_13_in03 = imem02_in[75:72];
    75: op1_13_in03 = reg_0547;
    76: op1_13_in03 = reg_0044;
    77: op1_13_in03 = reg_0805;
    78: op1_13_in03 = imem00_in[115:112];
    80: op1_13_in03 = reg_0637;
    81: op1_13_in03 = reg_0596;
    82: op1_13_in03 = reg_0204;
    83: op1_13_in03 = reg_0744;
    84: op1_13_in03 = reg_0819;
    85: op1_13_in03 = reg_0733;
    86: op1_13_in03 = reg_0075;
    87: op1_13_in03 = reg_0419;
    89: op1_13_in03 = reg_0515;
    90: op1_13_in03 = imem00_in[99:96];
    92: op1_13_in03 = imem04_in[71:68];
    93: op1_13_in03 = reg_0675;
    94: op1_13_in03 = reg_0707;
    95: op1_13_in03 = reg_0866;
    96: op1_13_in03 = imem05_in[91:88];
    default: op1_13_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv03 = 1;
    9: op1_13_inv03 = 1;
    10: op1_13_inv03 = 1;
    14: op1_13_inv03 = 1;
    17: op1_13_inv03 = 1;
    19: op1_13_inv03 = 1;
    20: op1_13_inv03 = 1;
    21: op1_13_inv03 = 1;
    22: op1_13_inv03 = 1;
    24: op1_13_inv03 = 1;
    4: op1_13_inv03 = 1;
    28: op1_13_inv03 = 1;
    3: op1_13_inv03 = 1;
    29: op1_13_inv03 = 1;
    32: op1_13_inv03 = 1;
    33: op1_13_inv03 = 1;
    34: op1_13_inv03 = 1;
    36: op1_13_inv03 = 1;
    39: op1_13_inv03 = 1;
    40: op1_13_inv03 = 1;
    41: op1_13_inv03 = 1;
    42: op1_13_inv03 = 1;
    44: op1_13_inv03 = 1;
    45: op1_13_inv03 = 1;
    46: op1_13_inv03 = 1;
    53: op1_13_inv03 = 1;
    55: op1_13_inv03 = 1;
    56: op1_13_inv03 = 1;
    57: op1_13_inv03 = 1;
    61: op1_13_inv03 = 1;
    62: op1_13_inv03 = 1;
    63: op1_13_inv03 = 1;
    65: op1_13_inv03 = 1;
    66: op1_13_inv03 = 1;
    71: op1_13_inv03 = 1;
    73: op1_13_inv03 = 1;
    75: op1_13_inv03 = 1;
    77: op1_13_inv03 = 1;
    78: op1_13_inv03 = 1;
    79: op1_13_inv03 = 1;
    81: op1_13_inv03 = 1;
    82: op1_13_inv03 = 1;
    84: op1_13_inv03 = 1;
    87: op1_13_inv03 = 1;
    90: op1_13_inv03 = 1;
    92: op1_13_inv03 = 1;
    93: op1_13_inv03 = 1;
    94: op1_13_inv03 = 1;
    95: op1_13_inv03 = 1;
    default: op1_13_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in04 = reg_0610;
    6: op1_13_in04 = reg_0282;
    7: op1_13_in04 = reg_0677;
    8: op1_13_in04 = imem02_in[15:12];
    9: op1_13_in04 = reg_0857;
    10: op1_13_in04 = reg_0331;
    11: op1_13_in04 = imem00_in[75:72];
    72: op1_13_in04 = imem00_in[75:72];
    12: op1_13_in04 = imem03_in[35:32];
    13: op1_13_in04 = imem00_in[107:104];
    14: op1_13_in04 = reg_1038;
    15: op1_13_in04 = reg_0369;
    16: op1_13_in04 = reg_0618;
    17: op1_13_in04 = reg_0676;
    18: op1_13_in04 = imem07_in[43:40];
    19: op1_13_in04 = reg_0671;
    20: op1_13_in04 = reg_0703;
    21: op1_13_in04 = reg_0122;
    22: op1_13_in04 = imem04_in[3:0];
    23: op1_13_in04 = imem06_in[75:72];
    24: op1_13_in04 = reg_0958;
    25: op1_13_in04 = reg_0799;
    26: op1_13_in04 = reg_0576;
    4: op1_13_in04 = reg_0440;
    27: op1_13_in04 = imem00_in[83:80];
    28: op1_13_in04 = reg_0685;
    3: op1_13_in04 = imem07_in[91:88];
    29: op1_13_in04 = imem05_in[79:76];
    30: op1_13_in04 = reg_0153;
    31: op1_13_in04 = reg_0121;
    32: op1_13_in04 = reg_1049;
    33: op1_13_in04 = reg_0977;
    34: op1_13_in04 = reg_0455;
    35: op1_13_in04 = reg_0500;
    36: op1_13_in04 = reg_0118;
    37: op1_13_in04 = reg_0996;
    38: op1_13_in04 = reg_0665;
    39: op1_13_in04 = imem06_in[111:108];
    40: op1_13_in04 = reg_0395;
    41: op1_13_in04 = imem07_in[107:104];
    42: op1_13_in04 = imem02_in[55:52];
    43: op1_13_in04 = imem04_in[127:124];
    44: op1_13_in04 = reg_1021;
    45: op1_13_in04 = reg_0691;
    46: op1_13_in04 = reg_0565;
    47: op1_13_in04 = reg_0251;
    48: op1_13_in04 = reg_0690;
    49: op1_13_in04 = reg_0106;
    50: op1_13_in04 = reg_0681;
    51: op1_13_in04 = imem07_in[127:124];
    52: op1_13_in04 = imem05_in[111:108];
    53: op1_13_in04 = reg_0002;
    54: op1_13_in04 = reg_0556;
    55: op1_13_in04 = imem00_in[95:92];
    56: op1_13_in04 = reg_0798;
    57: op1_13_in04 = reg_0003;
    58: op1_13_in04 = reg_0683;
    59: op1_13_in04 = imem03_in[23:20];
    60: op1_13_in04 = reg_1055;
    61: op1_13_in04 = reg_0807;
    62: op1_13_in04 = reg_0008;
    63: op1_13_in04 = reg_0519;
    90: op1_13_in04 = reg_0519;
    64: op1_13_in04 = imem00_in[103:100];
    65: op1_13_in04 = reg_0069;
    66: op1_13_in04 = reg_0829;
    67: op1_13_in04 = reg_0748;
    68: op1_13_in04 = reg_0390;
    69: op1_13_in04 = reg_0405;
    70: op1_13_in04 = reg_0733;
    71: op1_13_in04 = reg_0815;
    73: op1_13_in04 = reg_0745;
    74: op1_13_in04 = imem02_in[87:84];
    75: op1_13_in04 = reg_0298;
    76: op1_13_in04 = imem05_in[3:0];
    77: op1_13_in04 = reg_0303;
    78: op1_13_in04 = reg_0001;
    79: op1_13_in04 = imem00_in[87:84];
    80: op1_13_in04 = reg_0896;
    81: op1_13_in04 = reg_0239;
    82: op1_13_in04 = reg_0188;
    83: op1_13_in04 = reg_0315;
    84: op1_13_in04 = reg_0019;
    85: op1_13_in04 = reg_0555;
    86: op1_13_in04 = reg_0605;
    87: op1_13_in04 = reg_0599;
    88: op1_13_in04 = reg_1053;
    89: op1_13_in04 = reg_0164;
    91: op1_13_in04 = imem00_in[35:32];
    92: op1_13_in04 = imem04_in[99:96];
    93: op1_13_in04 = reg_0152;
    94: op1_13_in04 = reg_0970;
    95: op1_13_in04 = reg_0492;
    96: op1_13_in04 = imem05_in[127:124];
    default: op1_13_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv04 = 1;
    9: op1_13_inv04 = 1;
    10: op1_13_inv04 = 1;
    12: op1_13_inv04 = 1;
    14: op1_13_inv04 = 1;
    15: op1_13_inv04 = 1;
    19: op1_13_inv04 = 1;
    20: op1_13_inv04 = 1;
    23: op1_13_inv04 = 1;
    26: op1_13_inv04 = 1;
    27: op1_13_inv04 = 1;
    28: op1_13_inv04 = 1;
    3: op1_13_inv04 = 1;
    31: op1_13_inv04 = 1;
    32: op1_13_inv04 = 1;
    33: op1_13_inv04 = 1;
    34: op1_13_inv04 = 1;
    35: op1_13_inv04 = 1;
    36: op1_13_inv04 = 1;
    37: op1_13_inv04 = 1;
    40: op1_13_inv04 = 1;
    42: op1_13_inv04 = 1;
    43: op1_13_inv04 = 1;
    44: op1_13_inv04 = 1;
    45: op1_13_inv04 = 1;
    46: op1_13_inv04 = 1;
    48: op1_13_inv04 = 1;
    49: op1_13_inv04 = 1;
    50: op1_13_inv04 = 1;
    51: op1_13_inv04 = 1;
    53: op1_13_inv04 = 1;
    54: op1_13_inv04 = 1;
    58: op1_13_inv04 = 1;
    61: op1_13_inv04 = 1;
    62: op1_13_inv04 = 1;
    64: op1_13_inv04 = 1;
    65: op1_13_inv04 = 1;
    66: op1_13_inv04 = 1;
    67: op1_13_inv04 = 1;
    68: op1_13_inv04 = 1;
    70: op1_13_inv04 = 1;
    72: op1_13_inv04 = 1;
    73: op1_13_inv04 = 1;
    74: op1_13_inv04 = 1;
    75: op1_13_inv04 = 1;
    80: op1_13_inv04 = 1;
    81: op1_13_inv04 = 1;
    83: op1_13_inv04 = 1;
    84: op1_13_inv04 = 1;
    85: op1_13_inv04 = 1;
    87: op1_13_inv04 = 1;
    88: op1_13_inv04 = 1;
    89: op1_13_inv04 = 1;
    90: op1_13_inv04 = 1;
    91: op1_13_inv04 = 1;
    94: op1_13_inv04 = 1;
    96: op1_13_inv04 = 1;
    default: op1_13_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in05 = reg_0624;
    6: op1_13_in05 = reg_0306;
    7: op1_13_in05 = reg_0678;
    19: op1_13_in05 = reg_0678;
    8: op1_13_in05 = imem02_in[43:40];
    9: op1_13_in05 = reg_0876;
    10: op1_13_in05 = reg_0991;
    11: op1_13_in05 = imem00_in[115:112];
    12: op1_13_in05 = imem03_in[59:56];
    13: op1_13_in05 = reg_0672;
    14: op1_13_in05 = reg_0125;
    15: op1_13_in05 = reg_0385;
    39: op1_13_in05 = reg_0385;
    81: op1_13_in05 = reg_0385;
    16: op1_13_in05 = reg_0601;
    17: op1_13_in05 = reg_0689;
    18: op1_13_in05 = imem07_in[107:104];
    20: op1_13_in05 = reg_0724;
    21: op1_13_in05 = reg_0111;
    22: op1_13_in05 = imem04_in[47:44];
    23: op1_13_in05 = imem06_in[79:76];
    24: op1_13_in05 = reg_0966;
    25: op1_13_in05 = reg_1028;
    26: op1_13_in05 = reg_0395;
    4: op1_13_in05 = reg_0444;
    27: op1_13_in05 = imem00_in[87:84];
    28: op1_13_in05 = reg_0690;
    3: op1_13_in05 = imem07_in[95:92];
    29: op1_13_in05 = imem05_in[87:84];
    30: op1_13_in05 = reg_0140;
    31: op1_13_in05 = imem02_in[7:4];
    32: op1_13_in05 = reg_0046;
    33: op1_13_in05 = imem04_in[23:20];
    34: op1_13_in05 = reg_0469;
    35: op1_13_in05 = reg_1017;
    36: op1_13_in05 = reg_0117;
    37: op1_13_in05 = imem04_in[7:4];
    38: op1_13_in05 = reg_0636;
    40: op1_13_in05 = reg_0391;
    41: op1_13_in05 = imem07_in[111:108];
    42: op1_13_in05 = imem02_in[71:68];
    43: op1_13_in05 = reg_0265;
    44: op1_13_in05 = reg_0215;
    45: op1_13_in05 = reg_0688;
    46: op1_13_in05 = reg_0334;
    47: op1_13_in05 = reg_0816;
    48: op1_13_in05 = reg_0668;
    49: op1_13_in05 = reg_0115;
    50: op1_13_in05 = reg_0694;
    51: op1_13_in05 = reg_0730;
    52: op1_13_in05 = reg_0955;
    53: op1_13_in05 = reg_0250;
    54: op1_13_in05 = reg_0914;
    55: op1_13_in05 = reg_0463;
    56: op1_13_in05 = reg_0514;
    57: op1_13_in05 = reg_1053;
    58: op1_13_in05 = reg_0843;
    59: op1_13_in05 = imem03_in[35:32];
    60: op1_13_in05 = reg_0103;
    61: op1_13_in05 = reg_0836;
    62: op1_13_in05 = reg_0699;
    63: op1_13_in05 = reg_0738;
    64: op1_13_in05 = imem00_in[123:120];
    65: op1_13_in05 = reg_0749;
    66: op1_13_in05 = reg_0830;
    67: op1_13_in05 = reg_0670;
    68: op1_13_in05 = imem05_in[3:0];
    69: op1_13_in05 = reg_0264;
    70: op1_13_in05 = reg_0555;
    88: op1_13_in05 = reg_0555;
    71: op1_13_in05 = reg_0288;
    72: op1_13_in05 = imem00_in[83:80];
    73: op1_13_in05 = imem02_in[3:0];
    74: op1_13_in05 = imem02_in[99:96];
    75: op1_13_in05 = reg_0396;
    76: op1_13_in05 = imem05_in[19:16];
    77: op1_13_in05 = reg_0422;
    78: op1_13_in05 = reg_0682;
    79: op1_13_in05 = imem00_in[95:92];
    80: op1_13_in05 = reg_0096;
    82: op1_13_in05 = reg_0193;
    83: op1_13_in05 = reg_0532;
    84: op1_13_in05 = imem06_in[47:44];
    85: op1_13_in05 = reg_0101;
    86: op1_13_in05 = reg_0639;
    87: op1_13_in05 = reg_0427;
    89: op1_13_in05 = reg_0959;
    90: op1_13_in05 = reg_0685;
    91: op1_13_in05 = imem00_in[51:48];
    92: op1_13_in05 = reg_0577;
    93: op1_13_in05 = reg_0964;
    94: op1_13_in05 = reg_0252;
    95: op1_13_in05 = reg_0954;
    96: op1_13_in05 = reg_1021;
    default: op1_13_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv05 = 1;
    9: op1_13_inv05 = 1;
    10: op1_13_inv05 = 1;
    12: op1_13_inv05 = 1;
    15: op1_13_inv05 = 1;
    16: op1_13_inv05 = 1;
    17: op1_13_inv05 = 1;
    21: op1_13_inv05 = 1;
    22: op1_13_inv05 = 1;
    4: op1_13_inv05 = 1;
    27: op1_13_inv05 = 1;
    28: op1_13_inv05 = 1;
    3: op1_13_inv05 = 1;
    29: op1_13_inv05 = 1;
    30: op1_13_inv05 = 1;
    32: op1_13_inv05 = 1;
    33: op1_13_inv05 = 1;
    34: op1_13_inv05 = 1;
    35: op1_13_inv05 = 1;
    41: op1_13_inv05 = 1;
    43: op1_13_inv05 = 1;
    45: op1_13_inv05 = 1;
    46: op1_13_inv05 = 1;
    47: op1_13_inv05 = 1;
    49: op1_13_inv05 = 1;
    52: op1_13_inv05 = 1;
    54: op1_13_inv05 = 1;
    55: op1_13_inv05 = 1;
    57: op1_13_inv05 = 1;
    59: op1_13_inv05 = 1;
    60: op1_13_inv05 = 1;
    61: op1_13_inv05 = 1;
    62: op1_13_inv05 = 1;
    64: op1_13_inv05 = 1;
    68: op1_13_inv05 = 1;
    69: op1_13_inv05 = 1;
    70: op1_13_inv05 = 1;
    74: op1_13_inv05 = 1;
    75: op1_13_inv05 = 1;
    78: op1_13_inv05 = 1;
    79: op1_13_inv05 = 1;
    80: op1_13_inv05 = 1;
    85: op1_13_inv05 = 1;
    86: op1_13_inv05 = 1;
    88: op1_13_inv05 = 1;
    90: op1_13_inv05 = 1;
    95: op1_13_inv05 = 1;
    default: op1_13_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in06 = reg_0611;
    6: op1_13_in06 = reg_0275;
    7: op1_13_in06 = reg_0450;
    45: op1_13_in06 = reg_0450;
    90: op1_13_in06 = reg_0450;
    8: op1_13_in06 = imem02_in[47:44];
    9: op1_13_in06 = reg_0878;
    10: op1_13_in06 = imem04_in[11:8];
    11: op1_13_in06 = imem00_in[119:116];
    12: op1_13_in06 = imem03_in[103:100];
    13: op1_13_in06 = reg_0698;
    50: op1_13_in06 = reg_0698;
    14: op1_13_in06 = reg_0112;
    21: op1_13_in06 = reg_0112;
    15: op1_13_in06 = reg_0312;
    16: op1_13_in06 = reg_0402;
    17: op1_13_in06 = reg_0677;
    18: op1_13_in06 = reg_0704;
    41: op1_13_in06 = reg_0704;
    19: op1_13_in06 = reg_0476;
    20: op1_13_in06 = reg_0432;
    22: op1_13_in06 = imem04_in[59:56];
    23: op1_13_in06 = imem06_in[95:92];
    24: op1_13_in06 = reg_0957;
    52: op1_13_in06 = reg_0957;
    69: op1_13_in06 = reg_0957;
    25: op1_13_in06 = reg_0025;
    26: op1_13_in06 = reg_0373;
    4: op1_13_in06 = reg_0443;
    27: op1_13_in06 = imem00_in[95:92];
    72: op1_13_in06 = imem00_in[95:92];
    28: op1_13_in06 = reg_0477;
    3: op1_13_in06 = imem07_in[99:96];
    29: op1_13_in06 = reg_0944;
    96: op1_13_in06 = reg_0944;
    30: op1_13_in06 = reg_0155;
    31: op1_13_in06 = imem02_in[39:36];
    73: op1_13_in06 = imem02_in[39:36];
    32: op1_13_in06 = reg_0397;
    33: op1_13_in06 = imem04_in[47:44];
    34: op1_13_in06 = reg_0460;
    35: op1_13_in06 = reg_0105;
    36: op1_13_in06 = imem02_in[7:4];
    70: op1_13_in06 = imem02_in[7:4];
    37: op1_13_in06 = imem04_in[31:28];
    38: op1_13_in06 = reg_0663;
    39: op1_13_in06 = reg_0383;
    40: op1_13_in06 = reg_0386;
    42: op1_13_in06 = imem02_in[91:88];
    43: op1_13_in06 = reg_0540;
    44: op1_13_in06 = reg_0821;
    46: op1_13_in06 = reg_0842;
    47: op1_13_in06 = reg_0896;
    48: op1_13_in06 = reg_0680;
    49: op1_13_in06 = reg_0110;
    88: op1_13_in06 = reg_0110;
    51: op1_13_in06 = reg_0729;
    53: op1_13_in06 = reg_0433;
    54: op1_13_in06 = reg_0295;
    55: op1_13_in06 = reg_0451;
    56: op1_13_in06 = reg_0616;
    57: op1_13_in06 = reg_0114;
    58: op1_13_in06 = reg_0900;
    59: op1_13_in06 = imem03_in[87:84];
    60: op1_13_in06 = reg_0113;
    61: op1_13_in06 = reg_0998;
    62: op1_13_in06 = reg_0011;
    63: op1_13_in06 = reg_0753;
    64: op1_13_in06 = imem00_in[127:124];
    65: op1_13_in06 = reg_0669;
    66: op1_13_in06 = reg_0521;
    67: op1_13_in06 = reg_0883;
    68: op1_13_in06 = imem05_in[7:4];
    71: op1_13_in06 = reg_0444;
    74: op1_13_in06 = imem02_in[111:108];
    75: op1_13_in06 = reg_0596;
    76: op1_13_in06 = imem05_in[27:24];
    77: op1_13_in06 = reg_0421;
    78: op1_13_in06 = reg_0841;
    79: op1_13_in06 = reg_0519;
    80: op1_13_in06 = reg_0783;
    81: op1_13_in06 = reg_0551;
    82: op1_13_in06 = reg_0207;
    83: op1_13_in06 = reg_0350;
    84: op1_13_in06 = imem06_in[59:56];
    85: op1_13_in06 = reg_0115;
    86: op1_13_in06 = reg_0348;
    87: op1_13_in06 = reg_0502;
    89: op1_13_in06 = reg_0442;
    91: op1_13_in06 = imem00_in[63:60];
    92: op1_13_in06 = reg_0405;
    93: op1_13_in06 = reg_0530;
    94: op1_13_in06 = reg_0258;
    95: op1_13_in06 = reg_0139;
    default: op1_13_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv06 = 1;
    6: op1_13_inv06 = 1;
    8: op1_13_inv06 = 1;
    10: op1_13_inv06 = 1;
    12: op1_13_inv06 = 1;
    16: op1_13_inv06 = 1;
    19: op1_13_inv06 = 1;
    21: op1_13_inv06 = 1;
    23: op1_13_inv06 = 1;
    25: op1_13_inv06 = 1;
    26: op1_13_inv06 = 1;
    4: op1_13_inv06 = 1;
    27: op1_13_inv06 = 1;
    28: op1_13_inv06 = 1;
    3: op1_13_inv06 = 1;
    29: op1_13_inv06 = 1;
    35: op1_13_inv06 = 1;
    36: op1_13_inv06 = 1;
    39: op1_13_inv06 = 1;
    40: op1_13_inv06 = 1;
    41: op1_13_inv06 = 1;
    42: op1_13_inv06 = 1;
    44: op1_13_inv06 = 1;
    51: op1_13_inv06 = 1;
    52: op1_13_inv06 = 1;
    54: op1_13_inv06 = 1;
    55: op1_13_inv06 = 1;
    56: op1_13_inv06 = 1;
    59: op1_13_inv06 = 1;
    60: op1_13_inv06 = 1;
    61: op1_13_inv06 = 1;
    62: op1_13_inv06 = 1;
    63: op1_13_inv06 = 1;
    68: op1_13_inv06 = 1;
    69: op1_13_inv06 = 1;
    70: op1_13_inv06 = 1;
    71: op1_13_inv06 = 1;
    74: op1_13_inv06 = 1;
    79: op1_13_inv06 = 1;
    82: op1_13_inv06 = 1;
    86: op1_13_inv06 = 1;
    88: op1_13_inv06 = 1;
    90: op1_13_inv06 = 1;
    95: op1_13_inv06 = 1;
    default: op1_13_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in07 = reg_0623;
    6: op1_13_in07 = reg_0062;
    7: op1_13_in07 = reg_0473;
    8: op1_13_in07 = imem02_in[71:68];
    9: op1_13_in07 = reg_0628;
    10: op1_13_in07 = imem04_in[55:52];
    11: op1_13_in07 = reg_0695;
    62: op1_13_in07 = reg_0695;
    12: op1_13_in07 = reg_0583;
    13: op1_13_in07 = reg_0691;
    14: op1_13_in07 = reg_0106;
    15: op1_13_in07 = reg_0987;
    16: op1_13_in07 = reg_0372;
    17: op1_13_in07 = reg_0671;
    18: op1_13_in07 = reg_0719;
    19: op1_13_in07 = reg_0462;
    20: op1_13_in07 = reg_0183;
    21: op1_13_in07 = reg_0114;
    22: op1_13_in07 = imem04_in[67:64];
    23: op1_13_in07 = reg_0626;
    24: op1_13_in07 = reg_0969;
    25: op1_13_in07 = reg_0805;
    26: op1_13_in07 = reg_0376;
    4: op1_13_in07 = reg_0448;
    27: op1_13_in07 = imem00_in[111:108];
    28: op1_13_in07 = reg_0466;
    3: op1_13_in07 = imem07_in[107:104];
    29: op1_13_in07 = reg_0942;
    30: op1_13_in07 = reg_0137;
    31: op1_13_in07 = imem02_in[43:40];
    32: op1_13_in07 = reg_0004;
    33: op1_13_in07 = imem04_in[51:48];
    34: op1_13_in07 = reg_0458;
    35: op1_13_in07 = reg_0102;
    36: op1_13_in07 = imem02_in[19:16];
    88: op1_13_in07 = imem02_in[19:16];
    37: op1_13_in07 = imem04_in[63:60];
    38: op1_13_in07 = reg_0085;
    39: op1_13_in07 = reg_0399;
    40: op1_13_in07 = reg_0399;
    41: op1_13_in07 = reg_0726;
    42: op1_13_in07 = imem02_in[127:124];
    43: op1_13_in07 = reg_0537;
    44: op1_13_in07 = reg_0806;
    45: op1_13_in07 = reg_0455;
    46: op1_13_in07 = reg_0330;
    47: op1_13_in07 = reg_0831;
    48: op1_13_in07 = reg_0454;
    49: op1_13_in07 = imem02_in[11:8];
    50: op1_13_in07 = reg_0679;
    51: op1_13_in07 = reg_0715;
    52: op1_13_in07 = reg_0950;
    53: op1_13_in07 = reg_0589;
    54: op1_13_in07 = reg_0390;
    55: op1_13_in07 = reg_0464;
    56: op1_13_in07 = reg_0740;
    57: op1_13_in07 = reg_0101;
    58: op1_13_in07 = reg_0670;
    59: op1_13_in07 = imem03_in[119:116];
    60: op1_13_in07 = imem02_in[47:44];
    61: op1_13_in07 = reg_0982;
    81: op1_13_in07 = reg_0982;
    63: op1_13_in07 = reg_0749;
    64: op1_13_in07 = reg_0683;
    79: op1_13_in07 = reg_0683;
    65: op1_13_in07 = reg_0451;
    66: op1_13_in07 = reg_0616;
    67: op1_13_in07 = reg_0481;
    68: op1_13_in07 = imem05_in[35:32];
    69: op1_13_in07 = imem07_in[3:0];
    70: op1_13_in07 = imem02_in[51:48];
    71: op1_13_in07 = reg_0552;
    72: op1_13_in07 = imem00_in[99:96];
    73: op1_13_in07 = imem02_in[55:52];
    74: op1_13_in07 = imem02_in[115:112];
    75: op1_13_in07 = reg_0779;
    76: op1_13_in07 = imem05_in[31:28];
    77: op1_13_in07 = reg_0419;
    78: op1_13_in07 = reg_0900;
    80: op1_13_in07 = reg_0034;
    82: op1_13_in07 = imem01_in[19:16];
    83: op1_13_in07 = reg_0868;
    84: op1_13_in07 = imem06_in[87:84];
    85: op1_13_in07 = reg_0745;
    86: op1_13_in07 = reg_0637;
    87: op1_13_in07 = reg_0174;
    89: op1_13_in07 = reg_0718;
    90: op1_13_in07 = reg_0460;
    91: op1_13_in07 = imem00_in[67:64];
    92: op1_13_in07 = reg_1009;
    93: op1_13_in07 = reg_0960;
    94: op1_13_in07 = reg_0490;
    95: op1_13_in07 = reg_0138;
    96: op1_13_in07 = reg_0652;
    default: op1_13_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv07 = 1;
    6: op1_13_inv07 = 1;
    9: op1_13_inv07 = 1;
    10: op1_13_inv07 = 1;
    11: op1_13_inv07 = 1;
    12: op1_13_inv07 = 1;
    14: op1_13_inv07 = 1;
    15: op1_13_inv07 = 1;
    16: op1_13_inv07 = 1;
    17: op1_13_inv07 = 1;
    20: op1_13_inv07 = 1;
    22: op1_13_inv07 = 1;
    24: op1_13_inv07 = 1;
    26: op1_13_inv07 = 1;
    4: op1_13_inv07 = 1;
    29: op1_13_inv07 = 1;
    35: op1_13_inv07 = 1;
    39: op1_13_inv07 = 1;
    40: op1_13_inv07 = 1;
    41: op1_13_inv07 = 1;
    42: op1_13_inv07 = 1;
    44: op1_13_inv07 = 1;
    45: op1_13_inv07 = 1;
    47: op1_13_inv07 = 1;
    48: op1_13_inv07 = 1;
    49: op1_13_inv07 = 1;
    53: op1_13_inv07 = 1;
    54: op1_13_inv07 = 1;
    55: op1_13_inv07 = 1;
    56: op1_13_inv07 = 1;
    57: op1_13_inv07 = 1;
    58: op1_13_inv07 = 1;
    60: op1_13_inv07 = 1;
    61: op1_13_inv07 = 1;
    62: op1_13_inv07 = 1;
    63: op1_13_inv07 = 1;
    64: op1_13_inv07 = 1;
    66: op1_13_inv07 = 1;
    67: op1_13_inv07 = 1;
    68: op1_13_inv07 = 1;
    71: op1_13_inv07 = 1;
    73: op1_13_inv07 = 1;
    74: op1_13_inv07 = 1;
    76: op1_13_inv07 = 1;
    77: op1_13_inv07 = 1;
    80: op1_13_inv07 = 1;
    83: op1_13_inv07 = 1;
    84: op1_13_inv07 = 1;
    85: op1_13_inv07 = 1;
    90: op1_13_inv07 = 1;
    92: op1_13_inv07 = 1;
    94: op1_13_inv07 = 1;
    95: op1_13_inv07 = 1;
    96: op1_13_inv07 = 1;
    default: op1_13_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in08 = reg_0612;
    6: op1_13_in08 = reg_0067;
    7: op1_13_in08 = reg_0470;
    8: op1_13_in08 = imem02_in[75:72];
    9: op1_13_in08 = reg_0604;
    10: op1_13_in08 = imem04_in[59:56];
    11: op1_13_in08 = reg_0683;
    12: op1_13_in08 = reg_0592;
    13: op1_13_in08 = reg_0678;
    14: op1_13_in08 = reg_0109;
    15: op1_13_in08 = reg_0979;
    16: op1_13_in08 = reg_0368;
    17: op1_13_in08 = reg_0668;
    18: op1_13_in08 = reg_0717;
    19: op1_13_in08 = reg_0481;
    20: op1_13_in08 = reg_0166;
    21: op1_13_in08 = reg_0101;
    22: op1_13_in08 = imem04_in[71:68];
    23: op1_13_in08 = reg_0619;
    24: op1_13_in08 = reg_0942;
    25: op1_13_in08 = reg_0798;
    26: op1_13_in08 = reg_0998;
    4: op1_13_in08 = reg_0182;
    27: op1_13_in08 = imem00_in[119:116];
    28: op1_13_in08 = reg_0462;
    55: op1_13_in08 = reg_0462;
    3: op1_13_in08 = imem07_in[115:112];
    29: op1_13_in08 = reg_0952;
    30: op1_13_in08 = imem06_in[35:32];
    31: op1_13_in08 = imem02_in[59:56];
    32: op1_13_in08 = reg_0824;
    33: op1_13_in08 = imem04_in[87:84];
    34: op1_13_in08 = reg_0191;
    35: op1_13_in08 = reg_0126;
    36: op1_13_in08 = imem02_in[115:112];
    37: op1_13_in08 = imem04_in[111:108];
    38: op1_13_in08 = reg_0090;
    39: op1_13_in08 = reg_0630;
    40: op1_13_in08 = reg_0804;
    41: op1_13_in08 = reg_0729;
    42: op1_13_in08 = reg_0645;
    43: op1_13_in08 = reg_0799;
    44: op1_13_in08 = reg_0816;
    45: op1_13_in08 = reg_0464;
    46: op1_13_in08 = reg_0886;
    47: op1_13_in08 = reg_0147;
    48: op1_13_in08 = reg_0450;
    49: op1_13_in08 = imem02_in[19:16];
    50: op1_13_in08 = reg_0691;
    51: op1_13_in08 = reg_0303;
    52: op1_13_in08 = reg_0964;
    53: op1_13_in08 = reg_0420;
    77: op1_13_in08 = reg_0420;
    54: op1_13_in08 = reg_0222;
    56: op1_13_in08 = reg_0304;
    57: op1_13_in08 = reg_0877;
    58: op1_13_in08 = reg_0356;
    59: op1_13_in08 = reg_0580;
    60: op1_13_in08 = imem02_in[79:76];
    61: op1_13_in08 = reg_0996;
    62: op1_13_in08 = reg_0386;
    63: op1_13_in08 = reg_0463;
    64: op1_13_in08 = reg_0883;
    65: op1_13_in08 = reg_0477;
    66: op1_13_in08 = reg_0610;
    67: op1_13_in08 = reg_0480;
    68: op1_13_in08 = imem05_in[63:60];
    69: op1_13_in08 = imem07_in[19:16];
    70: op1_13_in08 = imem02_in[87:84];
    71: op1_13_in08 = reg_0108;
    72: op1_13_in08 = reg_0519;
    73: op1_13_in08 = imem02_in[111:108];
    74: op1_13_in08 = reg_0750;
    75: op1_13_in08 = reg_0376;
    76: op1_13_in08 = imem05_in[47:44];
    78: op1_13_in08 = reg_0842;
    79: op1_13_in08 = reg_0685;
    80: op1_13_in08 = reg_0763;
    81: op1_13_in08 = reg_0984;
    82: op1_13_in08 = imem01_in[35:32];
    83: op1_13_in08 = reg_0175;
    84: op1_13_in08 = reg_0625;
    85: op1_13_in08 = reg_0810;
    86: op1_13_in08 = reg_0279;
    87: op1_13_in08 = reg_0447;
    88: op1_13_in08 = imem02_in[71:68];
    89: op1_13_in08 = reg_0421;
    90: op1_13_in08 = reg_0214;
    91: op1_13_in08 = imem00_in[71:68];
    92: op1_13_in08 = reg_0390;
    93: op1_13_in08 = reg_0707;
    94: op1_13_in08 = reg_0144;
    95: op1_13_in08 = reg_0448;
    96: op1_13_in08 = reg_0647;
    default: op1_13_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv08 = 1;
    11: op1_13_inv08 = 1;
    12: op1_13_inv08 = 1;
    19: op1_13_inv08 = 1;
    20: op1_13_inv08 = 1;
    22: op1_13_inv08 = 1;
    24: op1_13_inv08 = 1;
    26: op1_13_inv08 = 1;
    4: op1_13_inv08 = 1;
    3: op1_13_inv08 = 1;
    29: op1_13_inv08 = 1;
    30: op1_13_inv08 = 1;
    31: op1_13_inv08 = 1;
    34: op1_13_inv08 = 1;
    35: op1_13_inv08 = 1;
    38: op1_13_inv08 = 1;
    39: op1_13_inv08 = 1;
    40: op1_13_inv08 = 1;
    44: op1_13_inv08 = 1;
    45: op1_13_inv08 = 1;
    46: op1_13_inv08 = 1;
    47: op1_13_inv08 = 1;
    49: op1_13_inv08 = 1;
    53: op1_13_inv08 = 1;
    54: op1_13_inv08 = 1;
    62: op1_13_inv08 = 1;
    64: op1_13_inv08 = 1;
    65: op1_13_inv08 = 1;
    67: op1_13_inv08 = 1;
    68: op1_13_inv08 = 1;
    77: op1_13_inv08 = 1;
    79: op1_13_inv08 = 1;
    80: op1_13_inv08 = 1;
    81: op1_13_inv08 = 1;
    82: op1_13_inv08 = 1;
    83: op1_13_inv08 = 1;
    85: op1_13_inv08 = 1;
    87: op1_13_inv08 = 1;
    89: op1_13_inv08 = 1;
    90: op1_13_inv08 = 1;
    91: op1_13_inv08 = 1;
    default: op1_13_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in09 = reg_0379;
    6: op1_13_in09 = reg_0056;
    7: op1_13_in09 = reg_0479;
    8: op1_13_in09 = imem02_in[119:116];
    9: op1_13_in09 = reg_0607;
    10: op1_13_in09 = imem04_in[115:112];
    11: op1_13_in09 = reg_0690;
    12: op1_13_in09 = reg_0600;
    13: op1_13_in09 = reg_0457;
    14: op1_13_in09 = imem02_in[3:0];
    15: op1_13_in09 = reg_0984;
    16: op1_13_in09 = reg_0808;
    17: op1_13_in09 = reg_0461;
    18: op1_13_in09 = reg_0703;
    19: op1_13_in09 = reg_0472;
    20: op1_13_in09 = reg_0164;
    21: op1_13_in09 = reg_0107;
    22: op1_13_in09 = imem04_in[79:76];
    23: op1_13_in09 = reg_0632;
    24: op1_13_in09 = reg_0949;
    25: op1_13_in09 = imem07_in[3:0];
    26: op1_13_in09 = reg_0991;
    27: op1_13_in09 = reg_0697;
    28: op1_13_in09 = reg_0200;
    3: op1_13_in09 = reg_0159;
    29: op1_13_in09 = reg_0960;
    30: op1_13_in09 = imem06_in[71:68];
    31: op1_13_in09 = imem02_in[87:84];
    60: op1_13_in09 = imem02_in[87:84];
    88: op1_13_in09 = imem02_in[87:84];
    32: op1_13_in09 = reg_0509;
    33: op1_13_in09 = imem04_in[99:96];
    34: op1_13_in09 = imem01_in[3:0];
    35: op1_13_in09 = imem02_in[19:16];
    57: op1_13_in09 = imem02_in[19:16];
    36: op1_13_in09 = imem02_in[127:124];
    37: op1_13_in09 = reg_1003;
    38: op1_13_in09 = reg_0091;
    39: op1_13_in09 = reg_0780;
    40: op1_13_in09 = reg_0332;
    41: op1_13_in09 = reg_0705;
    42: op1_13_in09 = reg_0653;
    70: op1_13_in09 = reg_0653;
    43: op1_13_in09 = reg_0076;
    44: op1_13_in09 = reg_0819;
    45: op1_13_in09 = reg_0460;
    46: op1_13_in09 = reg_0818;
    47: op1_13_in09 = reg_0146;
    48: op1_13_in09 = reg_0474;
    49: op1_13_in09 = imem02_in[43:40];
    50: op1_13_in09 = reg_0671;
    51: op1_13_in09 = reg_0250;
    52: op1_13_in09 = reg_0965;
    53: op1_13_in09 = reg_0024;
    54: op1_13_in09 = reg_0917;
    55: op1_13_in09 = reg_0480;
    56: op1_13_in09 = reg_0860;
    58: op1_13_in09 = reg_0674;
    78: op1_13_in09 = reg_0674;
    59: op1_13_in09 = reg_0874;
    61: op1_13_in09 = reg_0986;
    62: op1_13_in09 = reg_0371;
    63: op1_13_in09 = reg_0450;
    64: op1_13_in09 = reg_0668;
    65: op1_13_in09 = reg_0475;
    66: op1_13_in09 = reg_0304;
    67: op1_13_in09 = reg_0468;
    68: op1_13_in09 = imem05_in[67:64];
    69: op1_13_in09 = imem07_in[23:20];
    71: op1_13_in09 = reg_0542;
    72: op1_13_in09 = reg_0825;
    73: op1_13_in09 = reg_0803;
    74: op1_13_in09 = reg_0643;
    75: op1_13_in09 = reg_0385;
    76: op1_13_in09 = imem05_in[55:52];
    77: op1_13_in09 = reg_0165;
    79: op1_13_in09 = reg_0843;
    80: op1_13_in09 = reg_0341;
    81: op1_13_in09 = reg_0989;
    82: op1_13_in09 = imem01_in[43:40];
    83: op1_13_in09 = reg_0731;
    84: op1_13_in09 = reg_0244;
    85: op1_13_in09 = reg_0914;
    86: op1_13_in09 = reg_0441;
    87: op1_13_in09 = reg_0183;
    89: op1_13_in09 = reg_0406;
    90: op1_13_in09 = reg_0211;
    91: op1_13_in09 = imem00_in[111:108];
    92: op1_13_in09 = reg_0913;
    93: op1_13_in09 = reg_0970;
    94: op1_13_in09 = imem06_in[15:12];
    95: op1_13_in09 = reg_0269;
    96: op1_13_in09 = reg_0139;
    default: op1_13_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv09 = 1;
    6: op1_13_inv09 = 1;
    7: op1_13_inv09 = 1;
    9: op1_13_inv09 = 1;
    10: op1_13_inv09 = 1;
    12: op1_13_inv09 = 1;
    14: op1_13_inv09 = 1;
    18: op1_13_inv09 = 1;
    19: op1_13_inv09 = 1;
    21: op1_13_inv09 = 1;
    23: op1_13_inv09 = 1;
    24: op1_13_inv09 = 1;
    26: op1_13_inv09 = 1;
    28: op1_13_inv09 = 1;
    3: op1_13_inv09 = 1;
    31: op1_13_inv09 = 1;
    32: op1_13_inv09 = 1;
    34: op1_13_inv09 = 1;
    36: op1_13_inv09 = 1;
    38: op1_13_inv09 = 1;
    39: op1_13_inv09 = 1;
    40: op1_13_inv09 = 1;
    42: op1_13_inv09 = 1;
    43: op1_13_inv09 = 1;
    44: op1_13_inv09 = 1;
    48: op1_13_inv09 = 1;
    51: op1_13_inv09 = 1;
    54: op1_13_inv09 = 1;
    55: op1_13_inv09 = 1;
    58: op1_13_inv09 = 1;
    59: op1_13_inv09 = 1;
    60: op1_13_inv09 = 1;
    61: op1_13_inv09 = 1;
    62: op1_13_inv09 = 1;
    64: op1_13_inv09 = 1;
    67: op1_13_inv09 = 1;
    69: op1_13_inv09 = 1;
    71: op1_13_inv09 = 1;
    74: op1_13_inv09 = 1;
    75: op1_13_inv09 = 1;
    76: op1_13_inv09 = 1;
    77: op1_13_inv09 = 1;
    78: op1_13_inv09 = 1;
    79: op1_13_inv09 = 1;
    80: op1_13_inv09 = 1;
    84: op1_13_inv09 = 1;
    85: op1_13_inv09 = 1;
    87: op1_13_inv09 = 1;
    90: op1_13_inv09 = 1;
    92: op1_13_inv09 = 1;
    default: op1_13_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in10 = reg_0381;
    6: op1_13_in10 = reg_0068;
    7: op1_13_in10 = reg_0211;
    8: op1_13_in10 = reg_0658;
    9: op1_13_in10 = reg_0605;
    10: op1_13_in10 = reg_0540;
    11: op1_13_in10 = reg_0678;
    12: op1_13_in10 = reg_0578;
    13: op1_13_in10 = reg_0466;
    14: op1_13_in10 = imem02_in[43:40];
    15: op1_13_in10 = reg_0993;
    16: op1_13_in10 = reg_1028;
    17: op1_13_in10 = reg_0460;
    18: op1_13_in10 = reg_0724;
    19: op1_13_in10 = reg_0204;
    20: op1_13_in10 = reg_0178;
    21: op1_13_in10 = reg_0918;
    22: op1_13_in10 = imem04_in[87:84];
    23: op1_13_in10 = reg_0332;
    24: op1_13_in10 = reg_0965;
    93: op1_13_in10 = reg_0965;
    25: op1_13_in10 = imem07_in[23:20];
    26: op1_13_in10 = reg_0979;
    27: op1_13_in10 = reg_0672;
    28: op1_13_in10 = reg_0188;
    3: op1_13_in10 = reg_0160;
    29: op1_13_in10 = reg_0834;
    30: op1_13_in10 = reg_0610;
    31: op1_13_in10 = imem02_in[91:88];
    32: op1_13_in10 = reg_0820;
    33: op1_13_in10 = imem04_in[111:108];
    34: op1_13_in10 = imem01_in[7:4];
    35: op1_13_in10 = imem02_in[35:32];
    36: op1_13_in10 = reg_0646;
    37: op1_13_in10 = reg_0277;
    38: op1_13_in10 = imem03_in[59:56];
    39: op1_13_in10 = reg_0025;
    40: op1_13_in10 = reg_0241;
    41: op1_13_in10 = reg_0718;
    42: op1_13_in10 = reg_0663;
    43: op1_13_in10 = reg_0276;
    44: op1_13_in10 = reg_0132;
    45: op1_13_in10 = reg_0480;
    46: op1_13_in10 = reg_0762;
    47: op1_13_in10 = reg_0139;
    48: op1_13_in10 = reg_0479;
    49: op1_13_in10 = reg_0657;
    50: op1_13_in10 = reg_0688;
    51: op1_13_in10 = reg_0325;
    52: op1_13_in10 = reg_0961;
    53: op1_13_in10 = reg_0165;
    54: op1_13_in10 = reg_0017;
    55: op1_13_in10 = reg_0473;
    56: op1_13_in10 = reg_0101;
    57: op1_13_in10 = imem02_in[63:60];
    58: op1_13_in10 = reg_0753;
    59: op1_13_in10 = reg_0051;
    60: op1_13_in10 = imem02_in[111:108];
    61: op1_13_in10 = reg_0989;
    62: op1_13_in10 = reg_0916;
    63: op1_13_in10 = reg_0455;
    64: op1_13_in10 = reg_0687;
    65: op1_13_in10 = reg_0472;
    66: op1_13_in10 = reg_0615;
    67: op1_13_in10 = reg_0208;
    68: op1_13_in10 = imem05_in[95:92];
    69: op1_13_in10 = imem07_in[39:36];
    70: op1_13_in10 = reg_0341;
    71: op1_13_in10 = imem05_in[19:16];
    72: op1_13_in10 = reg_0748;
    73: op1_13_in10 = reg_0096;
    74: op1_13_in10 = reg_0908;
    75: op1_13_in10 = reg_1002;
    76: op1_13_in10 = imem05_in[75:72];
    77: op1_13_in10 = reg_0162;
    78: op1_13_in10 = reg_0749;
    79: op1_13_in10 = reg_0523;
    80: op1_13_in10 = reg_0765;
    81: op1_13_in10 = reg_1000;
    82: op1_13_in10 = imem01_in[63:60];
    83: op1_13_in10 = reg_0703;
    84: op1_13_in10 = reg_0614;
    85: op1_13_in10 = reg_0084;
    86: op1_13_in10 = reg_0424;
    87: op1_13_in10 = reg_0690;
    88: op1_13_in10 = imem02_in[115:112];
    89: op1_13_in10 = reg_0641;
    90: op1_13_in10 = reg_0198;
    91: op1_13_in10 = reg_0463;
    92: op1_13_in10 = reg_0430;
    94: op1_13_in10 = imem06_in[35:32];
    95: op1_13_in10 = reg_0063;
    96: op1_13_in10 = reg_0013;
    default: op1_13_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv10 = 1;
    9: op1_13_inv10 = 1;
    13: op1_13_inv10 = 1;
    14: op1_13_inv10 = 1;
    15: op1_13_inv10 = 1;
    16: op1_13_inv10 = 1;
    17: op1_13_inv10 = 1;
    18: op1_13_inv10 = 1;
    20: op1_13_inv10 = 1;
    21: op1_13_inv10 = 1;
    22: op1_13_inv10 = 1;
    23: op1_13_inv10 = 1;
    25: op1_13_inv10 = 1;
    26: op1_13_inv10 = 1;
    27: op1_13_inv10 = 1;
    28: op1_13_inv10 = 1;
    29: op1_13_inv10 = 1;
    30: op1_13_inv10 = 1;
    31: op1_13_inv10 = 1;
    33: op1_13_inv10 = 1;
    36: op1_13_inv10 = 1;
    37: op1_13_inv10 = 1;
    39: op1_13_inv10 = 1;
    41: op1_13_inv10 = 1;
    43: op1_13_inv10 = 1;
    46: op1_13_inv10 = 1;
    47: op1_13_inv10 = 1;
    51: op1_13_inv10 = 1;
    55: op1_13_inv10 = 1;
    56: op1_13_inv10 = 1;
    57: op1_13_inv10 = 1;
    58: op1_13_inv10 = 1;
    59: op1_13_inv10 = 1;
    60: op1_13_inv10 = 1;
    61: op1_13_inv10 = 1;
    67: op1_13_inv10 = 1;
    68: op1_13_inv10 = 1;
    71: op1_13_inv10 = 1;
    76: op1_13_inv10 = 1;
    77: op1_13_inv10 = 1;
    80: op1_13_inv10 = 1;
    83: op1_13_inv10 = 1;
    85: op1_13_inv10 = 1;
    86: op1_13_inv10 = 1;
    89: op1_13_inv10 = 1;
    91: op1_13_inv10 = 1;
    93: op1_13_inv10 = 1;
    94: op1_13_inv10 = 1;
    95: op1_13_inv10 = 1;
    default: op1_13_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in11 = reg_0351;
    6: op1_13_in11 = reg_0071;
    7: op1_13_in11 = reg_0201;
    8: op1_13_in11 = reg_0666;
    9: op1_13_in11 = reg_0408;
    10: op1_13_in11 = reg_0533;
    11: op1_13_in11 = reg_0680;
    12: op1_13_in11 = reg_0581;
    13: op1_13_in11 = reg_0480;
    14: op1_13_in11 = imem02_in[111:108];
    57: op1_13_in11 = imem02_in[111:108];
    15: op1_13_in11 = reg_0980;
    16: op1_13_in11 = reg_0753;
    17: op1_13_in11 = reg_0210;
    18: op1_13_in11 = reg_0708;
    19: op1_13_in11 = reg_0207;
    20: op1_13_in11 = reg_0176;
    21: op1_13_in11 = reg_0052;
    22: op1_13_in11 = imem04_in[119:116];
    23: op1_13_in11 = reg_0344;
    24: op1_13_in11 = reg_0953;
    25: op1_13_in11 = imem07_in[31:28];
    26: op1_13_in11 = reg_0984;
    27: op1_13_in11 = reg_0694;
    28: op1_13_in11 = reg_0203;
    3: op1_13_in11 = reg_0185;
    53: op1_13_in11 = reg_0185;
    29: op1_13_in11 = reg_0022;
    30: op1_13_in11 = reg_0608;
    31: op1_13_in11 = imem02_in[95:92];
    32: op1_13_in11 = reg_0982;
    33: op1_13_in11 = reg_1004;
    34: op1_13_in11 = imem01_in[11:8];
    35: op1_13_in11 = imem02_in[39:36];
    36: op1_13_in11 = reg_0660;
    37: op1_13_in11 = reg_0912;
    38: op1_13_in11 = imem03_in[79:76];
    39: op1_13_in11 = reg_0008;
    40: op1_13_in11 = reg_0017;
    41: op1_13_in11 = reg_0711;
    42: op1_13_in11 = reg_0334;
    43: op1_13_in11 = reg_0808;
    44: op1_13_in11 = reg_0128;
    45: op1_13_in11 = reg_0459;
    46: op1_13_in11 = reg_0083;
    47: op1_13_in11 = reg_0129;
    48: op1_13_in11 = reg_0458;
    49: op1_13_in11 = reg_0655;
    50: op1_13_in11 = reg_0465;
    64: op1_13_in11 = reg_0465;
    78: op1_13_in11 = reg_0465;
    91: op1_13_in11 = reg_0465;
    51: op1_13_in11 = reg_0589;
    52: op1_13_in11 = reg_0233;
    54: op1_13_in11 = reg_0025;
    55: op1_13_in11 = reg_0479;
    56: op1_13_in11 = reg_0109;
    58: op1_13_in11 = reg_0455;
    59: op1_13_in11 = reg_0993;
    60: op1_13_in11 = imem02_in[127:124];
    61: op1_13_in11 = reg_1000;
    62: op1_13_in11 = reg_0633;
    63: op1_13_in11 = reg_0469;
    65: op1_13_in11 = reg_0468;
    66: op1_13_in11 = reg_1051;
    67: op1_13_in11 = reg_0204;
    68: op1_13_in11 = reg_0940;
    69: op1_13_in11 = reg_0719;
    70: op1_13_in11 = reg_0837;
    71: op1_13_in11 = imem05_in[55:52];
    72: op1_13_in11 = reg_0684;
    73: op1_13_in11 = reg_0095;
    74: op1_13_in11 = reg_0323;
    75: op1_13_in11 = reg_0991;
    76: op1_13_in11 = imem05_in[83:80];
    77: op1_13_in11 = reg_0169;
    79: op1_13_in11 = reg_0669;
    80: op1_13_in11 = reg_0279;
    81: op1_13_in11 = reg_0997;
    82: op1_13_in11 = imem01_in[71:68];
    83: op1_13_in11 = reg_0539;
    84: op1_13_in11 = reg_0440;
    85: op1_13_in11 = reg_0308;
    86: op1_13_in11 = reg_0389;
    87: op1_13_in11 = reg_0157;
    88: op1_13_in11 = reg_0750;
    89: op1_13_in11 = reg_0868;
    90: op1_13_in11 = reg_0206;
    92: op1_13_in11 = reg_0864;
    93: op1_13_in11 = reg_0144;
    94: op1_13_in11 = imem06_in[75:72];
    95: op1_13_in11 = reg_0646;
    96: op1_13_in11 = reg_0226;
    default: op1_13_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv11 = 1;
    9: op1_13_inv11 = 1;
    12: op1_13_inv11 = 1;
    13: op1_13_inv11 = 1;
    15: op1_13_inv11 = 1;
    18: op1_13_inv11 = 1;
    19: op1_13_inv11 = 1;
    22: op1_13_inv11 = 1;
    24: op1_13_inv11 = 1;
    26: op1_13_inv11 = 1;
    27: op1_13_inv11 = 1;
    28: op1_13_inv11 = 1;
    3: op1_13_inv11 = 1;
    29: op1_13_inv11 = 1;
    34: op1_13_inv11 = 1;
    35: op1_13_inv11 = 1;
    37: op1_13_inv11 = 1;
    38: op1_13_inv11 = 1;
    39: op1_13_inv11 = 1;
    41: op1_13_inv11 = 1;
    42: op1_13_inv11 = 1;
    44: op1_13_inv11 = 1;
    45: op1_13_inv11 = 1;
    48: op1_13_inv11 = 1;
    50: op1_13_inv11 = 1;
    52: op1_13_inv11 = 1;
    53: op1_13_inv11 = 1;
    56: op1_13_inv11 = 1;
    59: op1_13_inv11 = 1;
    62: op1_13_inv11 = 1;
    63: op1_13_inv11 = 1;
    66: op1_13_inv11 = 1;
    67: op1_13_inv11 = 1;
    68: op1_13_inv11 = 1;
    74: op1_13_inv11 = 1;
    77: op1_13_inv11 = 1;
    78: op1_13_inv11 = 1;
    79: op1_13_inv11 = 1;
    81: op1_13_inv11 = 1;
    83: op1_13_inv11 = 1;
    84: op1_13_inv11 = 1;
    85: op1_13_inv11 = 1;
    86: op1_13_inv11 = 1;
    88: op1_13_inv11 = 1;
    89: op1_13_inv11 = 1;
    91: op1_13_inv11 = 1;
    94: op1_13_inv11 = 1;
    95: op1_13_inv11 = 1;
    default: op1_13_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in12 = reg_0382;
    6: op1_13_in12 = reg_0057;
    7: op1_13_in12 = reg_0205;
    8: op1_13_in12 = reg_0641;
    9: op1_13_in12 = reg_0351;
    10: op1_13_in12 = reg_0294;
    11: op1_13_in12 = reg_0669;
    12: op1_13_in12 = reg_0360;
    85: op1_13_in12 = reg_0360;
    13: op1_13_in12 = reg_0214;
    14: op1_13_in12 = imem02_in[123:120];
    57: op1_13_in12 = imem02_in[123:120];
    15: op1_13_in12 = reg_0977;
    75: op1_13_in12 = reg_0977;
    16: op1_13_in12 = reg_1010;
    17: op1_13_in12 = reg_0204;
    18: op1_13_in12 = reg_0718;
    19: op1_13_in12 = reg_0213;
    21: op1_13_in12 = reg_0881;
    22: op1_13_in12 = reg_0740;
    23: op1_13_in12 = reg_0381;
    24: op1_13_in12 = reg_0835;
    29: op1_13_in12 = reg_0835;
    25: op1_13_in12 = imem07_in[59:56];
    26: op1_13_in12 = reg_0996;
    27: op1_13_in12 = reg_0676;
    28: op1_13_in12 = reg_0186;
    30: op1_13_in12 = reg_0618;
    31: op1_13_in12 = imem02_in[103:100];
    32: op1_13_in12 = reg_0993;
    33: op1_13_in12 = reg_0536;
    34: op1_13_in12 = imem01_in[15:12];
    35: op1_13_in12 = imem02_in[43:40];
    36: op1_13_in12 = reg_0657;
    37: op1_13_in12 = reg_0539;
    38: op1_13_in12 = imem03_in[99:96];
    39: op1_13_in12 = imem07_in[35:32];
    40: op1_13_in12 = reg_0609;
    41: op1_13_in12 = reg_0429;
    42: op1_13_in12 = reg_0045;
    43: op1_13_in12 = reg_0528;
    44: op1_13_in12 = reg_0152;
    45: op1_13_in12 = reg_0203;
    46: op1_13_in12 = reg_0084;
    47: op1_13_in12 = reg_0141;
    48: op1_13_in12 = reg_0189;
    49: op1_13_in12 = reg_0654;
    50: op1_13_in12 = reg_0475;
    58: op1_13_in12 = reg_0475;
    51: op1_13_in12 = reg_0427;
    52: op1_13_in12 = reg_0259;
    53: op1_13_in12 = reg_0168;
    54: op1_13_in12 = reg_0531;
    55: op1_13_in12 = reg_0459;
    56: op1_13_in12 = imem02_in[23:20];
    59: op1_13_in12 = reg_0220;
    60: op1_13_in12 = reg_0363;
    61: op1_13_in12 = reg_0976;
    62: op1_13_in12 = reg_0219;
    63: op1_13_in12 = reg_0474;
    64: op1_13_in12 = reg_0455;
    65: op1_13_in12 = reg_0458;
    66: op1_13_in12 = reg_1055;
    67: op1_13_in12 = reg_0194;
    68: op1_13_in12 = reg_0508;
    69: op1_13_in12 = reg_0725;
    70: op1_13_in12 = reg_0424;
    74: op1_13_in12 = reg_0424;
    71: op1_13_in12 = imem05_in[59:56];
    72: op1_13_in12 = reg_0842;
    73: op1_13_in12 = reg_0081;
    76: op1_13_in12 = imem05_in[123:120];
    77: op1_13_in12 = reg_0182;
    78: op1_13_in12 = reg_0454;
    91: op1_13_in12 = reg_0454;
    79: op1_13_in12 = reg_0453;
    80: op1_13_in12 = reg_0052;
    81: op1_13_in12 = imem04_in[11:8];
    82: op1_13_in12 = imem01_in[99:96];
    83: op1_13_in12 = reg_0449;
    84: op1_13_in12 = reg_0297;
    86: op1_13_in12 = reg_0087;
    88: op1_13_in12 = reg_0334;
    89: op1_13_in12 = reg_0172;
    90: op1_13_in12 = reg_0199;
    92: op1_13_in12 = reg_0008;
    93: op1_13_in12 = imem06_in[3:0];
    94: op1_13_in12 = imem06_in[83:80];
    95: op1_13_in12 = reg_0695;
    96: op1_13_in12 = reg_0648;
    default: op1_13_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_13_inv12 = 1;
    10: op1_13_inv12 = 1;
    11: op1_13_inv12 = 1;
    12: op1_13_inv12 = 1;
    13: op1_13_inv12 = 1;
    15: op1_13_inv12 = 1;
    16: op1_13_inv12 = 1;
    21: op1_13_inv12 = 1;
    22: op1_13_inv12 = 1;
    25: op1_13_inv12 = 1;
    26: op1_13_inv12 = 1;
    28: op1_13_inv12 = 1;
    29: op1_13_inv12 = 1;
    31: op1_13_inv12 = 1;
    35: op1_13_inv12 = 1;
    36: op1_13_inv12 = 1;
    37: op1_13_inv12 = 1;
    38: op1_13_inv12 = 1;
    40: op1_13_inv12 = 1;
    41: op1_13_inv12 = 1;
    48: op1_13_inv12 = 1;
    49: op1_13_inv12 = 1;
    50: op1_13_inv12 = 1;
    51: op1_13_inv12 = 1;
    53: op1_13_inv12 = 1;
    56: op1_13_inv12 = 1;
    58: op1_13_inv12 = 1;
    61: op1_13_inv12 = 1;
    62: op1_13_inv12 = 1;
    63: op1_13_inv12 = 1;
    65: op1_13_inv12 = 1;
    67: op1_13_inv12 = 1;
    68: op1_13_inv12 = 1;
    70: op1_13_inv12 = 1;
    72: op1_13_inv12 = 1;
    73: op1_13_inv12 = 1;
    74: op1_13_inv12 = 1;
    75: op1_13_inv12 = 1;
    82: op1_13_inv12 = 1;
    83: op1_13_inv12 = 1;
    85: op1_13_inv12 = 1;
    86: op1_13_inv12 = 1;
    88: op1_13_inv12 = 1;
    89: op1_13_inv12 = 1;
    90: op1_13_inv12 = 1;
    93: op1_13_inv12 = 1;
    95: op1_13_inv12 = 1;
    default: op1_13_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in13 = reg_0383;
    6: op1_13_in13 = reg_0072;
    7: op1_13_in13 = imem01_in[99:96];
    8: op1_13_in13 = reg_0665;
    9: op1_13_in13 = reg_0409;
    10: op1_13_in13 = reg_0297;
    11: op1_13_in13 = reg_0457;
    12: op1_13_in13 = reg_0317;
    13: op1_13_in13 = reg_0194;
    48: op1_13_in13 = reg_0194;
    14: op1_13_in13 = imem02_in[127:124];
    15: op1_13_in13 = reg_1000;
    16: op1_13_in13 = imem07_in[19:16];
    17: op1_13_in13 = reg_0198;
    18: op1_13_in13 = reg_0727;
    19: op1_13_in13 = reg_0196;
    21: op1_13_in13 = reg_0655;
    22: op1_13_in13 = reg_0078;
    23: op1_13_in13 = reg_0408;
    24: op1_13_in13 = reg_0900;
    29: op1_13_in13 = reg_0900;
    25: op1_13_in13 = imem07_in[71:68];
    26: op1_13_in13 = reg_1001;
    27: op1_13_in13 = reg_0686;
    28: op1_13_in13 = reg_0195;
    30: op1_13_in13 = reg_0622;
    31: op1_13_in13 = reg_0666;
    32: op1_13_in13 = reg_0981;
    33: op1_13_in13 = reg_0540;
    34: op1_13_in13 = imem01_in[31:28];
    35: op1_13_in13 = imem02_in[123:120];
    36: op1_13_in13 = reg_0661;
    37: op1_13_in13 = reg_1057;
    38: op1_13_in13 = imem03_in[119:116];
    39: op1_13_in13 = imem07_in[103:100];
    40: op1_13_in13 = reg_0633;
    41: op1_13_in13 = reg_0448;
    42: op1_13_in13 = reg_0080;
    43: op1_13_in13 = reg_0053;
    44: op1_13_in13 = reg_0142;
    45: op1_13_in13 = reg_0211;
    46: op1_13_in13 = imem03_in[87:84];
    47: op1_13_in13 = imem06_in[3:0];
    49: op1_13_in13 = reg_0359;
    73: op1_13_in13 = reg_0359;
    50: op1_13_in13 = reg_0480;
    51: op1_13_in13 = reg_0868;
    52: op1_13_in13 = reg_0252;
    54: op1_13_in13 = imem07_in[23:20];
    55: op1_13_in13 = reg_0193;
    56: op1_13_in13 = imem02_in[43:40];
    57: op1_13_in13 = reg_0650;
    58: op1_13_in13 = reg_0468;
    59: op1_13_in13 = reg_0123;
    60: op1_13_in13 = reg_0646;
    61: op1_13_in13 = imem04_in[19:16];
    62: op1_13_in13 = imem07_in[39:36];
    63: op1_13_in13 = reg_0214;
    64: op1_13_in13 = reg_0477;
    91: op1_13_in13 = reg_0477;
    65: op1_13_in13 = reg_0204;
    66: op1_13_in13 = reg_0112;
    67: op1_13_in13 = reg_0206;
    68: op1_13_in13 = reg_0956;
    69: op1_13_in13 = reg_0718;
    70: op1_13_in13 = reg_0052;
    71: op1_13_in13 = reg_0217;
    72: op1_13_in13 = reg_0669;
    74: op1_13_in13 = reg_0423;
    75: op1_13_in13 = reg_0975;
    76: op1_13_in13 = reg_0215;
    77: op1_13_in13 = reg_0164;
    78: op1_13_in13 = reg_0451;
    79: op1_13_in13 = reg_0455;
    80: op1_13_in13 = reg_0329;
    81: op1_13_in13 = imem04_in[51:48];
    82: op1_13_in13 = imem01_in[107:104];
    83: op1_13_in13 = reg_0157;
    84: op1_13_in13 = reg_0698;
    85: op1_13_in13 = reg_0639;
    86: op1_13_in13 = reg_0608;
    88: op1_13_in13 = reg_0090;
    89: op1_13_in13 = reg_0179;
    90: op1_13_in13 = imem01_in[19:16];
    92: op1_13_in13 = reg_0752;
    93: op1_13_in13 = reg_1019;
    94: op1_13_in13 = imem06_in[103:100];
    95: op1_13_in13 = reg_0813;
    96: op1_13_in13 = reg_0259;
    default: op1_13_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv13 = 1;
    7: op1_13_inv13 = 1;
    8: op1_13_inv13 = 1;
    12: op1_13_inv13 = 1;
    13: op1_13_inv13 = 1;
    15: op1_13_inv13 = 1;
    16: op1_13_inv13 = 1;
    17: op1_13_inv13 = 1;
    19: op1_13_inv13 = 1;
    21: op1_13_inv13 = 1;
    23: op1_13_inv13 = 1;
    24: op1_13_inv13 = 1;
    26: op1_13_inv13 = 1;
    27: op1_13_inv13 = 1;
    28: op1_13_inv13 = 1;
    31: op1_13_inv13 = 1;
    32: op1_13_inv13 = 1;
    36: op1_13_inv13 = 1;
    38: op1_13_inv13 = 1;
    42: op1_13_inv13 = 1;
    46: op1_13_inv13 = 1;
    48: op1_13_inv13 = 1;
    50: op1_13_inv13 = 1;
    51: op1_13_inv13 = 1;
    54: op1_13_inv13 = 1;
    56: op1_13_inv13 = 1;
    59: op1_13_inv13 = 1;
    60: op1_13_inv13 = 1;
    61: op1_13_inv13 = 1;
    62: op1_13_inv13 = 1;
    65: op1_13_inv13 = 1;
    70: op1_13_inv13 = 1;
    71: op1_13_inv13 = 1;
    73: op1_13_inv13 = 1;
    78: op1_13_inv13 = 1;
    79: op1_13_inv13 = 1;
    84: op1_13_inv13 = 1;
    88: op1_13_inv13 = 1;
    90: op1_13_inv13 = 1;
    92: op1_13_inv13 = 1;
    94: op1_13_inv13 = 1;
    96: op1_13_inv13 = 1;
    default: op1_13_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in14 = reg_0315;
    6: op1_13_in14 = reg_0834;
    7: op1_13_in14 = reg_0523;
    8: op1_13_in14 = reg_0652;
    9: op1_13_in14 = reg_0401;
    10: op1_13_in14 = reg_0047;
    11: op1_13_in14 = reg_0459;
    12: op1_13_in14 = reg_0327;
    13: op1_13_in14 = imem01_in[55:52];
    14: op1_13_in14 = reg_0654;
    15: op1_13_in14 = reg_0997;
    16: op1_13_in14 = imem07_in[43:40];
    17: op1_13_in14 = reg_0212;
    18: op1_13_in14 = reg_0425;
    19: op1_13_in14 = reg_0195;
    21: op1_13_in14 = reg_0651;
    22: op1_13_in14 = reg_0259;
    23: op1_13_in14 = reg_0406;
    24: op1_13_in14 = reg_0757;
    29: op1_13_in14 = reg_0757;
    25: op1_13_in14 = imem07_in[79:76];
    26: op1_13_in14 = reg_0986;
    27: op1_13_in14 = reg_0670;
    28: op1_13_in14 = imem01_in[11:8];
    30: op1_13_in14 = reg_0623;
    31: op1_13_in14 = reg_0660;
    32: op1_13_in14 = reg_0977;
    33: op1_13_in14 = reg_0932;
    34: op1_13_in14 = imem01_in[35:32];
    35: op1_13_in14 = reg_0657;
    36: op1_13_in14 = reg_0662;
    37: op1_13_in14 = reg_0540;
    38: op1_13_in14 = reg_1007;
    39: op1_13_in14 = imem07_in[119:116];
    40: op1_13_in14 = reg_0029;
    41: op1_13_in14 = reg_0169;
    42: op1_13_in14 = reg_0817;
    43: op1_13_in14 = reg_0854;
    44: op1_13_in14 = reg_0134;
    45: op1_13_in14 = reg_0186;
    46: op1_13_in14 = reg_0580;
    47: op1_13_in14 = imem06_in[27:24];
    48: op1_13_in14 = reg_0192;
    67: op1_13_in14 = reg_0192;
    49: op1_13_in14 = reg_0082;
    50: op1_13_in14 = reg_0473;
    51: op1_13_in14 = reg_0164;
    52: op1_13_in14 = reg_0446;
    54: op1_13_in14 = imem07_in[39:36];
    55: op1_13_in14 = reg_0201;
    56: op1_13_in14 = imem02_in[91:88];
    57: op1_13_in14 = reg_0363;
    58: op1_13_in14 = reg_0452;
    59: op1_13_in14 = reg_0483;
    60: op1_13_in14 = reg_0639;
    61: op1_13_in14 = imem04_in[23:20];
    62: op1_13_in14 = imem07_in[67:64];
    63: op1_13_in14 = reg_0200;
    64: op1_13_in14 = reg_0472;
    65: op1_13_in14 = reg_0188;
    66: op1_13_in14 = reg_0109;
    68: op1_13_in14 = reg_0436;
    69: op1_13_in14 = reg_0433;
    70: op1_13_in14 = reg_0423;
    73: op1_13_in14 = reg_0423;
    80: op1_13_in14 = reg_0423;
    71: op1_13_in14 = reg_0951;
    72: op1_13_in14 = reg_0451;
    74: op1_13_in14 = reg_0331;
    75: op1_13_in14 = imem04_in[15:12];
    76: op1_13_in14 = reg_0136;
    77: op1_13_in14 = reg_0170;
    78: op1_13_in14 = reg_0461;
    79: op1_13_in14 = reg_0477;
    81: op1_13_in14 = imem04_in[71:68];
    82: op1_13_in14 = reg_0122;
    83: op1_13_in14 = reg_0697;
    84: op1_13_in14 = reg_0556;
    85: op1_13_in14 = reg_0077;
    86: op1_13_in14 = reg_0775;
    88: op1_13_in14 = reg_0887;
    89: op1_13_in14 = reg_0161;
    90: op1_13_in14 = imem01_in[75:72];
    91: op1_13_in14 = reg_0476;
    92: op1_13_in14 = reg_0584;
    93: op1_13_in14 = reg_0338;
    94: op1_13_in14 = imem06_in[111:108];
    95: op1_13_in14 = reg_0892;
    96: op1_13_in14 = reg_0152;
    default: op1_13_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv14 = 1;
    10: op1_13_inv14 = 1;
    12: op1_13_inv14 = 1;
    13: op1_13_inv14 = 1;
    16: op1_13_inv14 = 1;
    17: op1_13_inv14 = 1;
    18: op1_13_inv14 = 1;
    19: op1_13_inv14 = 1;
    24: op1_13_inv14 = 1;
    25: op1_13_inv14 = 1;
    27: op1_13_inv14 = 1;
    28: op1_13_inv14 = 1;
    37: op1_13_inv14 = 1;
    39: op1_13_inv14 = 1;
    42: op1_13_inv14 = 1;
    43: op1_13_inv14 = 1;
    46: op1_13_inv14 = 1;
    47: op1_13_inv14 = 1;
    48: op1_13_inv14 = 1;
    50: op1_13_inv14 = 1;
    54: op1_13_inv14 = 1;
    57: op1_13_inv14 = 1;
    62: op1_13_inv14 = 1;
    64: op1_13_inv14 = 1;
    67: op1_13_inv14 = 1;
    73: op1_13_inv14 = 1;
    75: op1_13_inv14 = 1;
    80: op1_13_inv14 = 1;
    82: op1_13_inv14 = 1;
    83: op1_13_inv14 = 1;
    86: op1_13_inv14 = 1;
    90: op1_13_inv14 = 1;
    91: op1_13_inv14 = 1;
    92: op1_13_inv14 = 1;
    94: op1_13_inv14 = 1;
    default: op1_13_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in15 = reg_0367;
    6: op1_13_in15 = reg_0821;
    7: op1_13_in15 = reg_0501;
    8: op1_13_in15 = reg_0320;
    9: op1_13_in15 = imem06_in[7:4];
    10: op1_13_in15 = reg_0066;
    11: op1_13_in15 = reg_0186;
    12: op1_13_in15 = reg_0312;
    13: op1_13_in15 = imem01_in[63:60];
    14: op1_13_in15 = reg_0661;
    15: op1_13_in15 = imem04_in[43:40];
    75: op1_13_in15 = imem04_in[43:40];
    16: op1_13_in15 = imem07_in[47:44];
    17: op1_13_in15 = reg_0190;
    18: op1_13_in15 = reg_0441;
    19: op1_13_in15 = reg_0197;
    21: op1_13_in15 = reg_0640;
    22: op1_13_in15 = reg_0755;
    23: op1_13_in15 = reg_0799;
    24: op1_13_in15 = reg_1046;
    25: op1_13_in15 = imem07_in[107:104];
    26: op1_13_in15 = reg_0990;
    27: op1_13_in15 = reg_0679;
    28: op1_13_in15 = imem01_in[27:24];
    29: op1_13_in15 = reg_0252;
    30: op1_13_in15 = reg_0615;
    31: op1_13_in15 = reg_0656;
    71: op1_13_in15 = reg_0656;
    32: op1_13_in15 = reg_0988;
    33: op1_13_in15 = reg_0537;
    34: op1_13_in15 = imem01_in[71:68];
    35: op1_13_in15 = reg_0662;
    36: op1_13_in15 = reg_0667;
    37: op1_13_in15 = reg_1016;
    38: op1_13_in15 = reg_1008;
    39: op1_13_in15 = imem07_in[123:120];
    40: op1_13_in15 = reg_0622;
    41: op1_13_in15 = reg_0183;
    42: op1_13_in15 = reg_0093;
    43: op1_13_in15 = reg_0773;
    44: op1_13_in15 = reg_0144;
    45: op1_13_in15 = reg_0198;
    46: op1_13_in15 = reg_0397;
    47: op1_13_in15 = imem06_in[39:36];
    48: op1_13_in15 = reg_1051;
    49: op1_13_in15 = reg_0637;
    50: op1_13_in15 = reg_0470;
    64: op1_13_in15 = reg_0470;
    51: op1_13_in15 = reg_0168;
    52: op1_13_in15 = reg_0438;
    54: op1_13_in15 = imem07_in[51:48];
    55: op1_13_in15 = reg_0205;
    56: op1_13_in15 = imem02_in[119:116];
    57: op1_13_in15 = reg_0657;
    58: op1_13_in15 = reg_0458;
    59: op1_13_in15 = reg_0530;
    60: op1_13_in15 = reg_0652;
    61: op1_13_in15 = imem04_in[55:52];
    62: op1_13_in15 = imem07_in[83:80];
    63: op1_13_in15 = reg_0210;
    65: op1_13_in15 = reg_0207;
    66: op1_13_in15 = reg_0103;
    67: op1_13_in15 = imem01_in[15:12];
    68: op1_13_in15 = reg_0447;
    69: op1_13_in15 = reg_0321;
    70: op1_13_in15 = reg_0087;
    72: op1_13_in15 = reg_0455;
    73: op1_13_in15 = reg_0368;
    74: op1_13_in15 = reg_0818;
    76: op1_13_in15 = reg_0944;
    78: op1_13_in15 = reg_0466;
    91: op1_13_in15 = reg_0466;
    79: op1_13_in15 = reg_0469;
    80: op1_13_in15 = reg_0389;
    81: op1_13_in15 = imem04_in[75:72];
    82: op1_13_in15 = reg_1042;
    84: op1_13_in15 = reg_0591;
    85: op1_13_in15 = reg_0095;
    86: op1_13_in15 = reg_0155;
    88: op1_13_in15 = reg_0323;
    89: op1_13_in15 = reg_0731;
    90: op1_13_in15 = imem01_in[83:80];
    92: op1_13_in15 = reg_0494;
    93: op1_13_in15 = reg_0754;
    94: op1_13_in15 = reg_0010;
    95: op1_13_in15 = reg_0964;
    96: op1_13_in15 = reg_0260;
    default: op1_13_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv15 = 1;
    7: op1_13_inv15 = 1;
    11: op1_13_inv15 = 1;
    12: op1_13_inv15 = 1;
    13: op1_13_inv15 = 1;
    15: op1_13_inv15 = 1;
    16: op1_13_inv15 = 1;
    18: op1_13_inv15 = 1;
    19: op1_13_inv15 = 1;
    24: op1_13_inv15 = 1;
    26: op1_13_inv15 = 1;
    27: op1_13_inv15 = 1;
    28: op1_13_inv15 = 1;
    29: op1_13_inv15 = 1;
    30: op1_13_inv15 = 1;
    31: op1_13_inv15 = 1;
    35: op1_13_inv15 = 1;
    36: op1_13_inv15 = 1;
    37: op1_13_inv15 = 1;
    38: op1_13_inv15 = 1;
    41: op1_13_inv15 = 1;
    44: op1_13_inv15 = 1;
    45: op1_13_inv15 = 1;
    46: op1_13_inv15 = 1;
    47: op1_13_inv15 = 1;
    49: op1_13_inv15 = 1;
    50: op1_13_inv15 = 1;
    51: op1_13_inv15 = 1;
    54: op1_13_inv15 = 1;
    55: op1_13_inv15 = 1;
    59: op1_13_inv15 = 1;
    61: op1_13_inv15 = 1;
    63: op1_13_inv15 = 1;
    65: op1_13_inv15 = 1;
    66: op1_13_inv15 = 1;
    67: op1_13_inv15 = 1;
    68: op1_13_inv15 = 1;
    71: op1_13_inv15 = 1;
    73: op1_13_inv15 = 1;
    74: op1_13_inv15 = 1;
    75: op1_13_inv15 = 1;
    76: op1_13_inv15 = 1;
    82: op1_13_inv15 = 1;
    85: op1_13_inv15 = 1;
    86: op1_13_inv15 = 1;
    94: op1_13_inv15 = 1;
    default: op1_13_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in16 = reg_0368;
    6: op1_13_in16 = reg_0835;
    7: op1_13_in16 = reg_0502;
    8: op1_13_in16 = reg_0330;
    9: op1_13_in16 = imem06_in[19:16];
    10: op1_13_in16 = reg_0076;
    11: op1_13_in16 = reg_0196;
    12: op1_13_in16 = reg_0397;
    13: op1_13_in16 = imem01_in[119:116];
    14: op1_13_in16 = reg_0665;
    15: op1_13_in16 = imem04_in[47:44];
    16: op1_13_in16 = imem07_in[75:72];
    17: op1_13_in16 = reg_0199;
    18: op1_13_in16 = reg_0428;
    19: op1_13_in16 = imem01_in[3:0];
    21: op1_13_in16 = reg_0334;
    22: op1_13_in16 = reg_0070;
    23: op1_13_in16 = reg_0752;
    24: op1_13_in16 = reg_0819;
    25: op1_13_in16 = imem07_in[119:116];
    26: op1_13_in16 = reg_1000;
    27: op1_13_in16 = reg_0678;
    28: op1_13_in16 = imem01_in[63:60];
    29: op1_13_in16 = reg_0260;
    95: op1_13_in16 = reg_0260;
    30: op1_13_in16 = reg_0914;
    31: op1_13_in16 = reg_0638;
    32: op1_13_in16 = reg_0990;
    33: op1_13_in16 = reg_0764;
    34: op1_13_in16 = reg_0235;
    35: op1_13_in16 = reg_0643;
    36: op1_13_in16 = reg_0045;
    37: op1_13_in16 = reg_0061;
    38: op1_13_in16 = reg_1019;
    39: op1_13_in16 = reg_0714;
    40: op1_13_in16 = imem07_in[3:0];
    41: op1_13_in16 = reg_0177;
    42: op1_13_in16 = reg_0083;
    43: op1_13_in16 = imem05_in[3:0];
    44: op1_13_in16 = imem06_in[3:0];
    45: op1_13_in16 = reg_0190;
    46: op1_13_in16 = reg_0389;
    47: op1_13_in16 = imem06_in[43:40];
    48: op1_13_in16 = reg_0623;
    49: op1_13_in16 = reg_0558;
    50: op1_13_in16 = reg_0471;
    51: op1_13_in16 = reg_0178;
    52: op1_13_in16 = reg_0148;
    54: op1_13_in16 = imem07_in[79:76];
    55: op1_13_in16 = imem01_in[35:32];
    56: op1_13_in16 = reg_0326;
    57: op1_13_in16 = reg_0326;
    58: op1_13_in16 = reg_0187;
    63: op1_13_in16 = reg_0187;
    59: op1_13_in16 = reg_0937;
    60: op1_13_in16 = reg_0837;
    61: op1_13_in16 = imem04_in[59:56];
    62: op1_13_in16 = imem07_in[103:100];
    64: op1_13_in16 = reg_0459;
    65: op1_13_in16 = reg_0186;
    66: op1_13_in16 = imem02_in[15:12];
    67: op1_13_in16 = imem01_in[79:76];
    68: op1_13_in16 = reg_0960;
    69: op1_13_in16 = reg_0315;
    70: op1_13_in16 = reg_0644;
    71: op1_13_in16 = reg_0486;
    72: op1_13_in16 = reg_0191;
    73: op1_13_in16 = reg_0248;
    74: op1_13_in16 = reg_0088;
    75: op1_13_in16 = imem04_in[91:88];
    76: op1_13_in16 = reg_0647;
    78: op1_13_in16 = reg_0452;
    79: op1_13_in16 = reg_0480;
    91: op1_13_in16 = reg_0480;
    80: op1_13_in16 = reg_0087;
    81: op1_13_in16 = imem04_in[79:76];
    82: op1_13_in16 = reg_0973;
    84: op1_13_in16 = reg_0380;
    85: op1_13_in16 = reg_0423;
    86: op1_13_in16 = reg_0086;
    88: op1_13_in16 = reg_0052;
    89: op1_13_in16 = reg_0182;
    90: op1_13_in16 = imem01_in[87:84];
    92: op1_13_in16 = reg_0071;
    93: op1_13_in16 = reg_0889;
    94: op1_13_in16 = reg_0895;
    96: op1_13_in16 = reg_0272;
    default: op1_13_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv16 = 1;
    6: op1_13_inv16 = 1;
    10: op1_13_inv16 = 1;
    14: op1_13_inv16 = 1;
    16: op1_13_inv16 = 1;
    17: op1_13_inv16 = 1;
    18: op1_13_inv16 = 1;
    19: op1_13_inv16 = 1;
    21: op1_13_inv16 = 1;
    24: op1_13_inv16 = 1;
    25: op1_13_inv16 = 1;
    26: op1_13_inv16 = 1;
    27: op1_13_inv16 = 1;
    30: op1_13_inv16 = 1;
    31: op1_13_inv16 = 1;
    33: op1_13_inv16 = 1;
    34: op1_13_inv16 = 1;
    37: op1_13_inv16 = 1;
    41: op1_13_inv16 = 1;
    42: op1_13_inv16 = 1;
    43: op1_13_inv16 = 1;
    44: op1_13_inv16 = 1;
    45: op1_13_inv16 = 1;
    48: op1_13_inv16 = 1;
    52: op1_13_inv16 = 1;
    56: op1_13_inv16 = 1;
    57: op1_13_inv16 = 1;
    59: op1_13_inv16 = 1;
    61: op1_13_inv16 = 1;
    64: op1_13_inv16 = 1;
    67: op1_13_inv16 = 1;
    68: op1_13_inv16 = 1;
    69: op1_13_inv16 = 1;
    71: op1_13_inv16 = 1;
    72: op1_13_inv16 = 1;
    80: op1_13_inv16 = 1;
    85: op1_13_inv16 = 1;
    86: op1_13_inv16 = 1;
    88: op1_13_inv16 = 1;
    93: op1_13_inv16 = 1;
    95: op1_13_inv16 = 1;
    default: op1_13_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in17 = reg_0031;
    6: op1_13_in17 = reg_0836;
    7: op1_13_in17 = reg_0515;
    8: op1_13_in17 = reg_0353;
    9: op1_13_in17 = imem06_in[23:20];
    10: op1_13_in17 = reg_0067;
    11: op1_13_in17 = reg_0197;
    12: op1_13_in17 = reg_0361;
    13: op1_13_in17 = imem01_in[123:120];
    14: op1_13_in17 = reg_0333;
    15: op1_13_in17 = imem04_in[59:56];
    16: op1_13_in17 = imem07_in[107:104];
    17: op1_13_in17 = imem01_in[71:68];
    18: op1_13_in17 = reg_0175;
    19: op1_13_in17 = imem01_in[11:8];
    65: op1_13_in17 = imem01_in[11:8];
    21: op1_13_in17 = reg_0341;
    22: op1_13_in17 = reg_0525;
    23: op1_13_in17 = reg_0801;
    24: op1_13_in17 = reg_0831;
    25: op1_13_in17 = imem07_in[123:120];
    26: op1_13_in17 = reg_0997;
    27: op1_13_in17 = reg_0687;
    28: op1_13_in17 = imem01_in[83:80];
    29: op1_13_in17 = reg_1046;
    30: op1_13_in17 = reg_0392;
    31: op1_13_in17 = reg_0663;
    32: op1_13_in17 = reg_0994;
    33: op1_13_in17 = reg_0061;
    34: op1_13_in17 = reg_0786;
    35: op1_13_in17 = reg_0886;
    36: op1_13_in17 = reg_0516;
    37: op1_13_in17 = reg_0268;
    38: op1_13_in17 = reg_1049;
    39: op1_13_in17 = reg_0715;
    40: op1_13_in17 = imem07_in[87:84];
    54: op1_13_in17 = imem07_in[87:84];
    41: op1_13_in17 = reg_0185;
    42: op1_13_in17 = reg_0007;
    80: op1_13_in17 = reg_0007;
    43: op1_13_in17 = imem05_in[51:48];
    44: op1_13_in17 = imem06_in[123:120];
    45: op1_13_in17 = reg_0195;
    46: op1_13_in17 = reg_0576;
    47: op1_13_in17 = imem06_in[55:52];
    48: op1_13_in17 = reg_0645;
    60: op1_13_in17 = reg_0645;
    49: op1_13_in17 = reg_0418;
    50: op1_13_in17 = reg_0200;
    64: op1_13_in17 = reg_0200;
    51: op1_13_in17 = reg_0173;
    52: op1_13_in17 = reg_0151;
    55: op1_13_in17 = imem01_in[59:56];
    56: op1_13_in17 = reg_0082;
    57: op1_13_in17 = reg_0646;
    58: op1_13_in17 = reg_0193;
    59: op1_13_in17 = reg_0912;
    61: op1_13_in17 = imem04_in[63:60];
    62: op1_13_in17 = imem07_in[115:112];
    63: op1_13_in17 = reg_0204;
    72: op1_13_in17 = reg_0204;
    66: op1_13_in17 = imem02_in[91:88];
    67: op1_13_in17 = imem01_in[91:88];
    68: op1_13_in17 = reg_0145;
    69: op1_13_in17 = reg_0589;
    70: op1_13_in17 = reg_0772;
    71: op1_13_in17 = reg_0941;
    73: op1_13_in17 = reg_0087;
    74: op1_13_in17 = reg_0761;
    75: op1_13_in17 = imem04_in[111:108];
    76: op1_13_in17 = reg_0137;
    78: op1_13_in17 = reg_0458;
    79: op1_13_in17 = reg_0468;
    81: op1_13_in17 = reg_0306;
    82: op1_13_in17 = reg_1014;
    84: op1_13_in17 = reg_0807;
    85: op1_13_in17 = reg_0818;
    86: op1_13_in17 = reg_0624;
    88: op1_13_in17 = reg_0423;
    89: op1_13_in17 = reg_0565;
    90: op1_13_in17 = reg_0105;
    91: op1_13_in17 = reg_0473;
    92: op1_13_in17 = imem05_in[23:20];
    93: op1_13_in17 = reg_0814;
    94: op1_13_in17 = reg_0792;
    95: op1_13_in17 = reg_0272;
    96: op1_13_in17 = reg_0530;
    default: op1_13_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv17 = 1;
    6: op1_13_inv17 = 1;
    7: op1_13_inv17 = 1;
    10: op1_13_inv17 = 1;
    12: op1_13_inv17 = 1;
    13: op1_13_inv17 = 1;
    14: op1_13_inv17 = 1;
    16: op1_13_inv17 = 1;
    18: op1_13_inv17 = 1;
    19: op1_13_inv17 = 1;
    21: op1_13_inv17 = 1;
    22: op1_13_inv17 = 1;
    24: op1_13_inv17 = 1;
    25: op1_13_inv17 = 1;
    26: op1_13_inv17 = 1;
    27: op1_13_inv17 = 1;
    28: op1_13_inv17 = 1;
    30: op1_13_inv17 = 1;
    32: op1_13_inv17 = 1;
    33: op1_13_inv17 = 1;
    34: op1_13_inv17 = 1;
    35: op1_13_inv17 = 1;
    36: op1_13_inv17 = 1;
    38: op1_13_inv17 = 1;
    39: op1_13_inv17 = 1;
    40: op1_13_inv17 = 1;
    41: op1_13_inv17 = 1;
    44: op1_13_inv17 = 1;
    45: op1_13_inv17 = 1;
    46: op1_13_inv17 = 1;
    48: op1_13_inv17 = 1;
    55: op1_13_inv17 = 1;
    56: op1_13_inv17 = 1;
    57: op1_13_inv17 = 1;
    62: op1_13_inv17 = 1;
    63: op1_13_inv17 = 1;
    64: op1_13_inv17 = 1;
    69: op1_13_inv17 = 1;
    71: op1_13_inv17 = 1;
    72: op1_13_inv17 = 1;
    75: op1_13_inv17 = 1;
    79: op1_13_inv17 = 1;
    80: op1_13_inv17 = 1;
    88: op1_13_inv17 = 1;
    91: op1_13_inv17 = 1;
    94: op1_13_inv17 = 1;
    95: op1_13_inv17 = 1;
    default: op1_13_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in18 = reg_0032;
    6: op1_13_in18 = reg_0837;
    49: op1_13_in18 = reg_0837;
    7: op1_13_in18 = reg_0505;
    8: op1_13_in18 = reg_0310;
    9: op1_13_in18 = imem06_in[71:68];
    10: op1_13_in18 = imem05_in[51:48];
    11: op1_13_in18 = reg_0790;
    12: op1_13_in18 = reg_0309;
    13: op1_13_in18 = reg_1051;
    14: op1_13_in18 = reg_0364;
    15: op1_13_in18 = imem04_in[71:68];
    16: op1_13_in18 = reg_0731;
    17: op1_13_in18 = imem01_in[75:72];
    18: op1_13_in18 = reg_0161;
    69: op1_13_in18 = reg_0161;
    19: op1_13_in18 = imem01_in[31:28];
    21: op1_13_in18 = reg_0359;
    22: op1_13_in18 = reg_0738;
    23: op1_13_in18 = reg_0025;
    24: op1_13_in18 = reg_0132;
    25: op1_13_in18 = reg_0719;
    26: op1_13_in18 = imem04_in[7:4];
    27: op1_13_in18 = reg_0669;
    28: op1_13_in18 = imem01_in[115:112];
    29: op1_13_in18 = reg_0832;
    30: op1_13_in18 = reg_0243;
    31: op1_13_in18 = reg_0842;
    32: op1_13_in18 = imem04_in[11:8];
    33: op1_13_in18 = reg_0063;
    34: op1_13_in18 = reg_0487;
    35: op1_13_in18 = reg_0339;
    36: op1_13_in18 = reg_0007;
    37: op1_13_in18 = reg_0071;
    38: op1_13_in18 = reg_0046;
    39: op1_13_in18 = reg_0436;
    40: op1_13_in18 = imem07_in[111:108];
    54: op1_13_in18 = imem07_in[111:108];
    41: op1_13_in18 = reg_0157;
    42: op1_13_in18 = reg_0814;
    43: op1_13_in18 = imem05_in[63:60];
    44: op1_13_in18 = reg_0407;
    45: op1_13_in18 = reg_0197;
    46: op1_13_in18 = reg_0823;
    47: op1_13_in18 = imem06_in[75:72];
    48: op1_13_in18 = imem01_in[3:0];
    50: op1_13_in18 = reg_0193;
    52: op1_13_in18 = reg_0138;
    55: op1_13_in18 = imem01_in[71:68];
    56: op1_13_in18 = reg_0300;
    57: op1_13_in18 = reg_0515;
    58: op1_13_in18 = reg_0205;
    59: op1_13_in18 = reg_0055;
    60: op1_13_in18 = reg_0441;
    61: op1_13_in18 = imem04_in[67:64];
    62: op1_13_in18 = imem07_in[127:124];
    63: op1_13_in18 = reg_0186;
    72: op1_13_in18 = reg_0186;
    64: op1_13_in18 = reg_0208;
    78: op1_13_in18 = reg_0208;
    65: op1_13_in18 = imem01_in[63:60];
    66: op1_13_in18 = imem02_in[127:124];
    67: op1_13_in18 = imem01_in[111:108];
    68: op1_13_in18 = reg_0130;
    70: op1_13_in18 = reg_0088;
    71: op1_13_in18 = reg_0948;
    73: op1_13_in18 = reg_0644;
    74: op1_13_in18 = reg_0484;
    75: op1_13_in18 = reg_1004;
    76: op1_13_in18 = reg_0648;
    79: op1_13_in18 = reg_0191;
    80: op1_13_in18 = reg_0482;
    81: op1_13_in18 = reg_1020;
    82: op1_13_in18 = reg_0337;
    84: op1_13_in18 = reg_0017;
    85: op1_13_in18 = reg_0087;
    86: op1_13_in18 = reg_0341;
    88: op1_13_in18 = reg_0516;
    89: op1_13_in18 = reg_0690;
    90: op1_13_in18 = reg_0968;
    91: op1_13_in18 = reg_0467;
    92: op1_13_in18 = imem05_in[35:32];
    93: op1_13_in18 = reg_0895;
    94: op1_13_in18 = reg_0698;
    95: op1_13_in18 = reg_0617;
    96: op1_13_in18 = reg_0972;
    default: op1_13_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv18 = 1;
    7: op1_13_inv18 = 1;
    8: op1_13_inv18 = 1;
    9: op1_13_inv18 = 1;
    15: op1_13_inv18 = 1;
    17: op1_13_inv18 = 1;
    21: op1_13_inv18 = 1;
    22: op1_13_inv18 = 1;
    24: op1_13_inv18 = 1;
    26: op1_13_inv18 = 1;
    27: op1_13_inv18 = 1;
    28: op1_13_inv18 = 1;
    31: op1_13_inv18 = 1;
    35: op1_13_inv18 = 1;
    37: op1_13_inv18 = 1;
    38: op1_13_inv18 = 1;
    40: op1_13_inv18 = 1;
    41: op1_13_inv18 = 1;
    42: op1_13_inv18 = 1;
    43: op1_13_inv18 = 1;
    46: op1_13_inv18 = 1;
    49: op1_13_inv18 = 1;
    50: op1_13_inv18 = 1;
    52: op1_13_inv18 = 1;
    55: op1_13_inv18 = 1;
    57: op1_13_inv18 = 1;
    58: op1_13_inv18 = 1;
    59: op1_13_inv18 = 1;
    60: op1_13_inv18 = 1;
    67: op1_13_inv18 = 1;
    70: op1_13_inv18 = 1;
    73: op1_13_inv18 = 1;
    75: op1_13_inv18 = 1;
    78: op1_13_inv18 = 1;
    79: op1_13_inv18 = 1;
    80: op1_13_inv18 = 1;
    84: op1_13_inv18 = 1;
    90: op1_13_inv18 = 1;
    91: op1_13_inv18 = 1;
    default: op1_13_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in19 = reg_0017;
    6: op1_13_in19 = imem05_in[3:0];
    7: op1_13_in19 = reg_0232;
    8: op1_13_in19 = reg_0355;
    9: op1_13_in19 = imem07_in[23:20];
    10: op1_13_in19 = imem05_in[75:72];
    11: op1_13_in19 = reg_0792;
    12: op1_13_in19 = reg_0374;
    13: op1_13_in19 = reg_0247;
    14: op1_13_in19 = reg_0320;
    15: op1_13_in19 = imem04_in[91:88];
    61: op1_13_in19 = imem04_in[91:88];
    16: op1_13_in19 = reg_0714;
    17: op1_13_in19 = imem01_in[95:92];
    18: op1_13_in19 = reg_0169;
    19: op1_13_in19 = imem01_in[47:44];
    21: op1_13_in19 = reg_0329;
    22: op1_13_in19 = reg_0751;
    23: op1_13_in19 = reg_0018;
    24: op1_13_in19 = reg_0136;
    25: op1_13_in19 = reg_0730;
    26: op1_13_in19 = imem04_in[15:12];
    32: op1_13_in19 = imem04_in[15:12];
    27: op1_13_in19 = reg_0453;
    28: op1_13_in19 = reg_0013;
    29: op1_13_in19 = reg_0819;
    30: op1_13_in19 = reg_0222;
    31: op1_13_in19 = reg_0080;
    33: op1_13_in19 = reg_0296;
    34: op1_13_in19 = reg_1039;
    35: op1_13_in19 = reg_0817;
    36: op1_13_in19 = reg_0761;
    80: op1_13_in19 = reg_0761;
    37: op1_13_in19 = reg_0882;
    38: op1_13_in19 = reg_0793;
    39: op1_13_in19 = reg_0422;
    40: op1_13_in19 = imem07_in[119:116];
    54: op1_13_in19 = imem07_in[119:116];
    41: op1_13_in19 = reg_0158;
    42: op1_13_in19 = reg_0084;
    43: op1_13_in19 = imem05_in[115:112];
    44: op1_13_in19 = reg_0556;
    45: op1_13_in19 = imem01_in[7:4];
    46: op1_13_in19 = reg_0038;
    47: op1_13_in19 = imem06_in[107:104];
    48: op1_13_in19 = imem01_in[79:76];
    49: op1_13_in19 = reg_0096;
    50: op1_13_in19 = reg_0202;
    52: op1_13_in19 = reg_0141;
    55: op1_13_in19 = reg_0586;
    56: op1_13_in19 = reg_0652;
    57: op1_13_in19 = reg_0637;
    58: op1_13_in19 = imem01_in[11:8];
    59: op1_13_in19 = reg_0048;
    60: op1_13_in19 = reg_0039;
    62: op1_13_in19 = reg_0719;
    63: op1_13_in19 = reg_0194;
    64: op1_13_in19 = reg_0203;
    65: op1_13_in19 = imem01_in[91:88];
    66: op1_13_in19 = reg_0290;
    67: op1_13_in19 = imem01_in[115:112];
    68: op1_13_in19 = reg_0140;
    69: op1_13_in19 = reg_0162;
    70: op1_13_in19 = reg_0089;
    71: op1_13_in19 = reg_0436;
    72: op1_13_in19 = reg_0196;
    73: op1_13_in19 = reg_0335;
    74: op1_13_in19 = imem03_in[15:12];
    75: op1_13_in19 = reg_0483;
    76: op1_13_in19 = reg_0966;
    78: op1_13_in19 = reg_0210;
    79: op1_13_in19 = reg_0210;
    81: op1_13_in19 = reg_0540;
    82: op1_13_in19 = reg_0971;
    84: op1_13_in19 = reg_0835;
    85: op1_13_in19 = reg_0644;
    86: op1_13_in19 = reg_0367;
    88: op1_13_in19 = reg_0347;
    90: op1_13_in19 = reg_0337;
    91: op1_13_in19 = reg_0471;
    92: op1_13_in19 = imem05_in[39:36];
    93: op1_13_in19 = reg_0698;
    94: op1_13_in19 = reg_0918;
    95: op1_13_in19 = reg_0530;
    96: op1_13_in19 = reg_0806;
    default: op1_13_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_13_inv19 = 1;
    12: op1_13_inv19 = 1;
    13: op1_13_inv19 = 1;
    14: op1_13_inv19 = 1;
    16: op1_13_inv19 = 1;
    17: op1_13_inv19 = 1;
    18: op1_13_inv19 = 1;
    19: op1_13_inv19 = 1;
    22: op1_13_inv19 = 1;
    23: op1_13_inv19 = 1;
    31: op1_13_inv19 = 1;
    32: op1_13_inv19 = 1;
    35: op1_13_inv19 = 1;
    37: op1_13_inv19 = 1;
    43: op1_13_inv19 = 1;
    44: op1_13_inv19 = 1;
    45: op1_13_inv19 = 1;
    46: op1_13_inv19 = 1;
    49: op1_13_inv19 = 1;
    54: op1_13_inv19 = 1;
    55: op1_13_inv19 = 1;
    56: op1_13_inv19 = 1;
    57: op1_13_inv19 = 1;
    59: op1_13_inv19 = 1;
    60: op1_13_inv19 = 1;
    61: op1_13_inv19 = 1;
    62: op1_13_inv19 = 1;
    64: op1_13_inv19 = 1;
    65: op1_13_inv19 = 1;
    67: op1_13_inv19 = 1;
    68: op1_13_inv19 = 1;
    70: op1_13_inv19 = 1;
    71: op1_13_inv19 = 1;
    73: op1_13_inv19 = 1;
    76: op1_13_inv19 = 1;
    79: op1_13_inv19 = 1;
    81: op1_13_inv19 = 1;
    84: op1_13_inv19 = 1;
    86: op1_13_inv19 = 1;
    91: op1_13_inv19 = 1;
    93: op1_13_inv19 = 1;
    95: op1_13_inv19 = 1;
    default: op1_13_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in20 = reg_0020;
    6: op1_13_in20 = imem05_in[7:4];
    7: op1_13_in20 = reg_0222;
    8: op1_13_in20 = reg_0095;
    9: op1_13_in20 = imem07_in[71:68];
    10: op1_13_in20 = imem05_in[103:100];
    11: op1_13_in20 = imem01_in[7:4];
    12: op1_13_in20 = reg_0389;
    13: op1_13_in20 = reg_0503;
    14: op1_13_in20 = reg_0346;
    15: op1_13_in20 = reg_0545;
    16: op1_13_in20 = reg_0724;
    17: op1_13_in20 = imem01_in[103:100];
    48: op1_13_in20 = imem01_in[103:100];
    18: op1_13_in20 = reg_0182;
    19: op1_13_in20 = imem01_in[67:64];
    21: op1_13_in20 = reg_0318;
    22: op1_13_in20 = reg_0773;
    23: op1_13_in20 = imem07_in[11:8];
    24: op1_13_in20 = reg_0129;
    25: op1_13_in20 = reg_0710;
    26: op1_13_in20 = imem04_in[19:16];
    32: op1_13_in20 = imem04_in[19:16];
    27: op1_13_in20 = reg_0469;
    28: op1_13_in20 = reg_0560;
    29: op1_13_in20 = reg_0497;
    30: op1_13_in20 = reg_0787;
    31: op1_13_in20 = reg_0290;
    33: op1_13_in20 = reg_0009;
    34: op1_13_in20 = reg_0230;
    35: op1_13_in20 = reg_0261;
    36: op1_13_in20 = reg_0261;
    37: op1_13_in20 = reg_0528;
    38: op1_13_in20 = reg_0765;
    39: op1_13_in20 = reg_0447;
    40: op1_13_in20 = imem07_in[127:124];
    42: op1_13_in20 = reg_0291;
    43: op1_13_in20 = reg_0962;
    44: op1_13_in20 = reg_0403;
    45: op1_13_in20 = imem01_in[11:8];
    46: op1_13_in20 = reg_0311;
    47: op1_13_in20 = reg_0883;
    49: op1_13_in20 = reg_0097;
    50: op1_13_in20 = imem01_in[3:0];
    52: op1_13_in20 = reg_0137;
    54: op1_13_in20 = reg_0716;
    55: op1_13_in20 = reg_0904;
    56: op1_13_in20 = reg_0837;
    57: op1_13_in20 = reg_0279;
    58: op1_13_in20 = reg_0933;
    59: op1_13_in20 = reg_1057;
    60: op1_13_in20 = reg_0372;
    61: op1_13_in20 = imem04_in[99:96];
    62: op1_13_in20 = reg_0730;
    63: op1_13_in20 = reg_0213;
    64: op1_13_in20 = reg_0194;
    65: op1_13_in20 = imem01_in[95:92];
    66: op1_13_in20 = reg_0914;
    67: op1_13_in20 = reg_0586;
    68: op1_13_in20 = imem06_in[11:8];
    69: op1_13_in20 = reg_0167;
    70: op1_13_in20 = reg_0876;
    71: op1_13_in20 = reg_0150;
    72: op1_13_in20 = reg_0192;
    73: op1_13_in20 = reg_0083;
    74: op1_13_in20 = imem03_in[83:80];
    75: op1_13_in20 = reg_1006;
    76: op1_13_in20 = reg_0786;
    78: op1_13_in20 = reg_0189;
    79: op1_13_in20 = reg_0207;
    80: op1_13_in20 = reg_0049;
    81: op1_13_in20 = reg_1016;
    82: op1_13_in20 = reg_1023;
    84: op1_13_in20 = reg_0369;
    85: op1_13_in20 = reg_0037;
    86: op1_13_in20 = imem03_in[3:0];
    88: op1_13_in20 = reg_0045;
    90: op1_13_in20 = reg_0592;
    91: op1_13_in20 = reg_0456;
    92: op1_13_in20 = imem05_in[43:40];
    93: op1_13_in20 = reg_0611;
    94: op1_13_in20 = reg_0133;
    95: op1_13_in20 = reg_0972;
    96: op1_13_in20 = reg_0252;
    default: op1_13_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv20 = 1;
    13: op1_13_inv20 = 1;
    15: op1_13_inv20 = 1;
    18: op1_13_inv20 = 1;
    19: op1_13_inv20 = 1;
    25: op1_13_inv20 = 1;
    26: op1_13_inv20 = 1;
    28: op1_13_inv20 = 1;
    36: op1_13_inv20 = 1;
    37: op1_13_inv20 = 1;
    38: op1_13_inv20 = 1;
    39: op1_13_inv20 = 1;
    42: op1_13_inv20 = 1;
    45: op1_13_inv20 = 1;
    47: op1_13_inv20 = 1;
    49: op1_13_inv20 = 1;
    54: op1_13_inv20 = 1;
    55: op1_13_inv20 = 1;
    56: op1_13_inv20 = 1;
    58: op1_13_inv20 = 1;
    61: op1_13_inv20 = 1;
    63: op1_13_inv20 = 1;
    64: op1_13_inv20 = 1;
    66: op1_13_inv20 = 1;
    67: op1_13_inv20 = 1;
    69: op1_13_inv20 = 1;
    70: op1_13_inv20 = 1;
    71: op1_13_inv20 = 1;
    72: op1_13_inv20 = 1;
    74: op1_13_inv20 = 1;
    75: op1_13_inv20 = 1;
    76: op1_13_inv20 = 1;
    79: op1_13_inv20 = 1;
    84: op1_13_inv20 = 1;
    85: op1_13_inv20 = 1;
    88: op1_13_inv20 = 1;
    93: op1_13_inv20 = 1;
    94: op1_13_inv20 = 1;
    95: op1_13_inv20 = 1;
    default: op1_13_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in21 = reg_0018;
    6: op1_13_in21 = imem05_in[71:68];
    7: op1_13_in21 = reg_0246;
    8: op1_13_in21 = reg_0082;
    9: op1_13_in21 = imem07_in[75:72];
    10: op1_13_in21 = imem05_in[111:108];
    11: op1_13_in21 = imem01_in[11:8];
    12: op1_13_in21 = reg_0985;
    13: op1_13_in21 = reg_0236;
    14: op1_13_in21 = reg_0092;
    15: op1_13_in21 = reg_0536;
    16: op1_13_in21 = reg_0708;
    17: op1_13_in21 = imem01_in[127:124];
    18: op1_13_in21 = reg_0160;
    19: op1_13_in21 = imem01_in[91:88];
    21: op1_13_in21 = reg_0342;
    22: op1_13_in21 = reg_0044;
    23: op1_13_in21 = imem07_in[23:20];
    24: op1_13_in21 = imem06_in[19:16];
    25: op1_13_in21 = reg_0731;
    54: op1_13_in21 = reg_0731;
    26: op1_13_in21 = imem04_in[43:40];
    27: op1_13_in21 = reg_0472;
    28: op1_13_in21 = reg_0239;
    29: op1_13_in21 = reg_0132;
    30: op1_13_in21 = reg_0027;
    31: op1_13_in21 = reg_0086;
    32: op1_13_in21 = imem04_in[39:36];
    33: op1_13_in21 = reg_0278;
    34: op1_13_in21 = reg_1036;
    35: op1_13_in21 = reg_0077;
    36: op1_13_in21 = reg_0049;
    37: op1_13_in21 = reg_0517;
    38: op1_13_in21 = reg_0820;
    39: op1_13_in21 = reg_0428;
    40: op1_13_in21 = reg_0728;
    42: op1_13_in21 = imem03_in[11:8];
    80: op1_13_in21 = imem03_in[11:8];
    86: op1_13_in21 = imem03_in[11:8];
    43: op1_13_in21 = reg_0970;
    44: op1_13_in21 = reg_0783;
    45: op1_13_in21 = imem01_in[35:32];
    50: op1_13_in21 = imem01_in[35:32];
    46: op1_13_in21 = reg_0767;
    47: op1_13_in21 = reg_0915;
    48: op1_13_in21 = reg_0520;
    49: op1_13_in21 = reg_0083;
    52: op1_13_in21 = imem06_in[7:4];
    55: op1_13_in21 = reg_0933;
    56: op1_13_in21 = reg_0359;
    57: op1_13_in21 = reg_0358;
    58: op1_13_in21 = reg_0870;
    59: op1_13_in21 = reg_0932;
    60: op1_13_in21 = reg_0818;
    61: op1_13_in21 = imem04_in[111:108];
    62: op1_13_in21 = reg_0717;
    63: op1_13_in21 = imem01_in[31:28];
    64: op1_13_in21 = reg_0202;
    65: op1_13_in21 = imem01_in[115:112];
    66: op1_13_in21 = reg_0036;
    67: op1_13_in21 = reg_0285;
    68: op1_13_in21 = imem06_in[67:64];
    69: op1_13_in21 = reg_0170;
    70: op1_13_in21 = reg_0261;
    71: op1_13_in21 = reg_0151;
    72: op1_13_in21 = imem01_in[3:0];
    73: op1_13_in21 = reg_0007;
    74: op1_13_in21 = imem03_in[107:104];
    75: op1_13_in21 = reg_0301;
    76: op1_13_in21 = reg_0438;
    78: op1_13_in21 = reg_0193;
    79: op1_13_in21 = reg_0186;
    81: op1_13_in21 = reg_0752;
    82: op1_13_in21 = reg_1056;
    84: op1_13_in21 = imem07_in[79:76];
    85: op1_13_in21 = imem02_in[7:4];
    88: op1_13_in21 = reg_0355;
    90: op1_13_in21 = reg_1035;
    91: op1_13_in21 = reg_0458;
    92: op1_13_in21 = imem05_in[99:96];
    93: op1_13_in21 = reg_0403;
    94: op1_13_in21 = reg_0124;
    95: op1_13_in21 = reg_0707;
    96: op1_13_in21 = reg_0816;
    default: op1_13_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv21 = 1;
    13: op1_13_inv21 = 1;
    14: op1_13_inv21 = 1;
    17: op1_13_inv21 = 1;
    18: op1_13_inv21 = 1;
    19: op1_13_inv21 = 1;
    21: op1_13_inv21 = 1;
    23: op1_13_inv21 = 1;
    24: op1_13_inv21 = 1;
    25: op1_13_inv21 = 1;
    30: op1_13_inv21 = 1;
    31: op1_13_inv21 = 1;
    33: op1_13_inv21 = 1;
    35: op1_13_inv21 = 1;
    36: op1_13_inv21 = 1;
    37: op1_13_inv21 = 1;
    39: op1_13_inv21 = 1;
    42: op1_13_inv21 = 1;
    45: op1_13_inv21 = 1;
    46: op1_13_inv21 = 1;
    48: op1_13_inv21 = 1;
    49: op1_13_inv21 = 1;
    55: op1_13_inv21 = 1;
    58: op1_13_inv21 = 1;
    59: op1_13_inv21 = 1;
    60: op1_13_inv21 = 1;
    64: op1_13_inv21 = 1;
    66: op1_13_inv21 = 1;
    74: op1_13_inv21 = 1;
    79: op1_13_inv21 = 1;
    80: op1_13_inv21 = 1;
    88: op1_13_inv21 = 1;
    91: op1_13_inv21 = 1;
    92: op1_13_inv21 = 1;
    93: op1_13_inv21 = 1;
    94: op1_13_inv21 = 1;
    95: op1_13_inv21 = 1;
    default: op1_13_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in22 = imem07_in[3:0];
    94: op1_13_in22 = imem07_in[3:0];
    6: op1_13_in22 = imem05_in[95:92];
    7: op1_13_in22 = reg_0224;
    8: op1_13_in22 = reg_0055;
    9: op1_13_in22 = imem07_in[79:76];
    10: op1_13_in22 = imem05_in[123:120];
    11: op1_13_in22 = imem01_in[27:24];
    12: op1_13_in22 = reg_1002;
    13: op1_13_in22 = reg_0234;
    90: op1_13_in22 = reg_0234;
    14: op1_13_in22 = reg_0084;
    15: op1_13_in22 = reg_0550;
    16: op1_13_in22 = reg_0707;
    17: op1_13_in22 = reg_0235;
    18: op1_13_in22 = reg_0183;
    19: op1_13_in22 = reg_0508;
    21: op1_13_in22 = reg_0336;
    22: op1_13_in22 = imem05_in[35:32];
    23: op1_13_in22 = imem07_in[123:120];
    24: op1_13_in22 = imem06_in[87:84];
    25: op1_13_in22 = reg_0703;
    26: op1_13_in22 = imem04_in[59:56];
    27: op1_13_in22 = reg_0200;
    28: op1_13_in22 = reg_0555;
    29: op1_13_in22 = reg_0145;
    95: op1_13_in22 = reg_0145;
    30: op1_13_in22 = reg_0808;
    31: op1_13_in22 = reg_0090;
    32: op1_13_in22 = imem04_in[63:60];
    33: op1_13_in22 = reg_0059;
    34: op1_13_in22 = reg_0111;
    35: op1_13_in22 = reg_0872;
    36: op1_13_in22 = reg_0840;
    37: op1_13_in22 = reg_0856;
    38: op1_13_in22 = reg_0844;
    39: op1_13_in22 = reg_0443;
    40: op1_13_in22 = reg_0719;
    42: op1_13_in22 = imem03_in[71:68];
    43: op1_13_in22 = reg_0955;
    44: op1_13_in22 = reg_0042;
    45: op1_13_in22 = imem01_in[39:36];
    46: op1_13_in22 = reg_0374;
    47: op1_13_in22 = reg_0892;
    48: op1_13_in22 = reg_1043;
    49: op1_13_in22 = reg_0007;
    50: op1_13_in22 = imem01_in[47:44];
    52: op1_13_in22 = imem06_in[47:44];
    54: op1_13_in22 = reg_0713;
    55: op1_13_in22 = reg_1056;
    56: op1_13_in22 = reg_0248;
    57: op1_13_in22 = reg_0039;
    58: op1_13_in22 = reg_0919;
    59: op1_13_in22 = reg_0541;
    60: op1_13_in22 = reg_0037;
    61: op1_13_in22 = reg_0483;
    62: op1_13_in22 = reg_0575;
    63: op1_13_in22 = imem01_in[35:32];
    64: op1_13_in22 = imem01_in[19:16];
    65: op1_13_in22 = reg_0242;
    66: op1_13_in22 = reg_0087;
    67: op1_13_in22 = reg_0520;
    68: op1_13_in22 = imem06_in[75:72];
    70: op1_13_in22 = reg_0091;
    71: op1_13_in22 = reg_0142;
    72: op1_13_in22 = imem01_in[63:60];
    73: op1_13_in22 = reg_0758;
    74: op1_13_in22 = imem03_in[123:120];
    75: op1_13_in22 = reg_0530;
    76: op1_13_in22 = reg_0651;
    78: op1_13_in22 = reg_0194;
    79: op1_13_in22 = reg_0192;
    80: op1_13_in22 = imem03_in[35:32];
    81: op1_13_in22 = reg_0568;
    82: op1_13_in22 = reg_1024;
    84: op1_13_in22 = reg_0515;
    85: op1_13_in22 = imem02_in[91:88];
    86: op1_13_in22 = imem03_in[15:12];
    88: op1_13_in22 = reg_0778;
    91: op1_13_in22 = reg_0198;
    92: op1_13_in22 = imem05_in[115:112];
    93: op1_13_in22 = reg_0222;
    96: op1_13_in22 = reg_0949;
    default: op1_13_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv22 = 1;
    6: op1_13_inv22 = 1;
    7: op1_13_inv22 = 1;
    9: op1_13_inv22 = 1;
    10: op1_13_inv22 = 1;
    11: op1_13_inv22 = 1;
    14: op1_13_inv22 = 1;
    15: op1_13_inv22 = 1;
    16: op1_13_inv22 = 1;
    17: op1_13_inv22 = 1;
    21: op1_13_inv22 = 1;
    24: op1_13_inv22 = 1;
    25: op1_13_inv22 = 1;
    26: op1_13_inv22 = 1;
    27: op1_13_inv22 = 1;
    32: op1_13_inv22 = 1;
    34: op1_13_inv22 = 1;
    36: op1_13_inv22 = 1;
    37: op1_13_inv22 = 1;
    38: op1_13_inv22 = 1;
    43: op1_13_inv22 = 1;
    45: op1_13_inv22 = 1;
    46: op1_13_inv22 = 1;
    47: op1_13_inv22 = 1;
    54: op1_13_inv22 = 1;
    55: op1_13_inv22 = 1;
    58: op1_13_inv22 = 1;
    59: op1_13_inv22 = 1;
    62: op1_13_inv22 = 1;
    65: op1_13_inv22 = 1;
    66: op1_13_inv22 = 1;
    67: op1_13_inv22 = 1;
    70: op1_13_inv22 = 1;
    71: op1_13_inv22 = 1;
    72: op1_13_inv22 = 1;
    86: op1_13_inv22 = 1;
    88: op1_13_inv22 = 1;
    93: op1_13_inv22 = 1;
    94: op1_13_inv22 = 1;
    95: op1_13_inv22 = 1;
    default: op1_13_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in23 = imem07_in[27:24];
    6: op1_13_in23 = imem05_in[107:104];
    7: op1_13_in23 = reg_0220;
    8: op1_13_in23 = reg_0077;
    9: op1_13_in23 = reg_0719;
    10: op1_13_in23 = imem05_in[127:124];
    92: op1_13_in23 = imem05_in[127:124];
    11: op1_13_in23 = imem01_in[115:112];
    12: op1_13_in23 = reg_0994;
    13: op1_13_in23 = reg_1052;
    14: op1_13_in23 = reg_0098;
    15: op1_13_in23 = reg_0548;
    16: op1_13_in23 = reg_0700;
    17: op1_13_in23 = reg_0508;
    18: op1_13_in23 = reg_0170;
    19: op1_13_in23 = reg_0226;
    21: op1_13_in23 = imem02_in[27:24];
    22: op1_13_in23 = imem05_in[39:36];
    23: op1_13_in23 = reg_0723;
    24: op1_13_in23 = reg_0625;
    25: op1_13_in23 = reg_0712;
    26: op1_13_in23 = imem04_in[71:68];
    27: op1_13_in23 = reg_0197;
    28: op1_13_in23 = reg_0828;
    29: op1_13_in23 = reg_0135;
    30: op1_13_in23 = reg_1028;
    31: op1_13_in23 = reg_0049;
    32: op1_13_in23 = imem04_in[75:72];
    33: op1_13_in23 = reg_0054;
    34: op1_13_in23 = reg_0118;
    35: op1_13_in23 = imem03_in[3:0];
    36: op1_13_in23 = reg_0484;
    37: op1_13_in23 = imem05_in[7:4];
    38: op1_13_in23 = reg_0979;
    39: op1_13_in23 = reg_0448;
    40: op1_13_in23 = reg_0725;
    42: op1_13_in23 = imem03_in[115:112];
    43: op1_13_in23 = reg_0956;
    44: op1_13_in23 = reg_0393;
    45: op1_13_in23 = imem01_in[47:44];
    46: op1_13_in23 = reg_0987;
    47: op1_13_in23 = reg_0403;
    48: op1_13_in23 = reg_0829;
    49: op1_13_in23 = reg_0776;
    50: op1_13_in23 = reg_0586;
    52: op1_13_in23 = imem06_in[51:48];
    54: op1_13_in23 = reg_0744;
    55: op1_13_in23 = reg_0487;
    56: op1_13_in23 = reg_0644;
    57: op1_13_in23 = reg_0347;
    58: op1_13_in23 = reg_0238;
    59: op1_13_in23 = reg_0313;
    60: op1_13_in23 = reg_0335;
    61: op1_13_in23 = reg_1003;
    62: op1_13_in23 = reg_0002;
    63: op1_13_in23 = imem01_in[39:36];
    64: op1_13_in23 = imem01_in[35:32];
    65: op1_13_in23 = reg_1056;
    66: op1_13_in23 = reg_0007;
    67: op1_13_in23 = reg_0521;
    68: op1_13_in23 = imem06_in[95:92];
    70: op1_13_in23 = reg_0840;
    71: op1_13_in23 = reg_0156;
    72: op1_13_in23 = reg_1042;
    73: op1_13_in23 = imem03_in[11:8];
    74: op1_13_in23 = reg_0572;
    75: op1_13_in23 = reg_0937;
    76: op1_13_in23 = reg_0741;
    96: op1_13_in23 = reg_0741;
    78: op1_13_in23 = imem01_in[19:16];
    79: op1_13_in23 = imem01_in[3:0];
    80: op1_13_in23 = imem03_in[39:36];
    81: op1_13_in23 = reg_0067;
    82: op1_13_in23 = reg_0862;
    84: op1_13_in23 = reg_0299;
    85: op1_13_in23 = imem02_in[95:92];
    86: op1_13_in23 = imem03_in[35:32];
    88: op1_13_in23 = reg_0656;
    90: op1_13_in23 = reg_0607;
    91: op1_13_in23 = reg_0190;
    93: op1_13_in23 = reg_0566;
    94: op1_13_in23 = imem07_in[11:8];
    95: op1_13_in23 = reg_0709;
    default: op1_13_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv23 = 1;
    11: op1_13_inv23 = 1;
    13: op1_13_inv23 = 1;
    14: op1_13_inv23 = 1;
    17: op1_13_inv23 = 1;
    21: op1_13_inv23 = 1;
    23: op1_13_inv23 = 1;
    25: op1_13_inv23 = 1;
    28: op1_13_inv23 = 1;
    30: op1_13_inv23 = 1;
    31: op1_13_inv23 = 1;
    32: op1_13_inv23 = 1;
    34: op1_13_inv23 = 1;
    35: op1_13_inv23 = 1;
    36: op1_13_inv23 = 1;
    37: op1_13_inv23 = 1;
    39: op1_13_inv23 = 1;
    40: op1_13_inv23 = 1;
    42: op1_13_inv23 = 1;
    45: op1_13_inv23 = 1;
    46: op1_13_inv23 = 1;
    47: op1_13_inv23 = 1;
    49: op1_13_inv23 = 1;
    59: op1_13_inv23 = 1;
    62: op1_13_inv23 = 1;
    64: op1_13_inv23 = 1;
    66: op1_13_inv23 = 1;
    68: op1_13_inv23 = 1;
    70: op1_13_inv23 = 1;
    71: op1_13_inv23 = 1;
    72: op1_13_inv23 = 1;
    75: op1_13_inv23 = 1;
    78: op1_13_inv23 = 1;
    79: op1_13_inv23 = 1;
    80: op1_13_inv23 = 1;
    81: op1_13_inv23 = 1;
    88: op1_13_inv23 = 1;
    90: op1_13_inv23 = 1;
    91: op1_13_inv23 = 1;
    92: op1_13_inv23 = 1;
    96: op1_13_inv23 = 1;
    default: op1_13_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in24 = reg_0722;
    6: op1_13_in24 = imem05_in[119:116];
    7: op1_13_in24 = reg_0247;
    8: op1_13_in24 = reg_0093;
    9: op1_13_in24 = reg_0726;
    10: op1_13_in24 = reg_0954;
    11: op1_13_in24 = imem01_in[119:116];
    12: op1_13_in24 = imem04_in[55:52];
    13: op1_13_in24 = reg_1042;
    19: op1_13_in24 = reg_1042;
    14: op1_13_in24 = reg_0055;
    15: op1_13_in24 = reg_0558;
    16: op1_13_in24 = reg_0423;
    17: op1_13_in24 = reg_1032;
    18: op1_13_in24 = reg_0176;
    21: op1_13_in24 = imem02_in[47:44];
    22: op1_13_in24 = imem05_in[55:52];
    23: op1_13_in24 = reg_0711;
    24: op1_13_in24 = reg_0604;
    90: op1_13_in24 = reg_0604;
    25: op1_13_in24 = reg_0707;
    26: op1_13_in24 = imem04_in[87:84];
    27: op1_13_in24 = imem01_in[7:4];
    28: op1_13_in24 = reg_0248;
    29: op1_13_in24 = reg_0151;
    30: op1_13_in24 = reg_0025;
    31: op1_13_in24 = reg_0531;
    32: op1_13_in24 = imem04_in[115:112];
    33: op1_13_in24 = reg_0058;
    34: op1_13_in24 = imem02_in[35:32];
    35: op1_13_in24 = imem03_in[15:12];
    36: op1_13_in24 = imem03_in[7:4];
    37: op1_13_in24 = imem05_in[31:28];
    38: op1_13_in24 = reg_0993;
    39: op1_13_in24 = reg_0431;
    40: op1_13_in24 = reg_0706;
    42: op1_13_in24 = imem03_in[127:124];
    43: op1_13_in24 = reg_0948;
    44: op1_13_in24 = reg_0295;
    45: op1_13_in24 = imem01_in[55:52];
    46: op1_13_in24 = reg_0983;
    47: op1_13_in24 = reg_0632;
    48: op1_13_in24 = reg_1037;
    49: op1_13_in24 = reg_0086;
    50: op1_13_in24 = reg_0779;
    52: op1_13_in24 = imem06_in[87:84];
    54: op1_13_in24 = reg_0428;
    55: op1_13_in24 = reg_0514;
    56: op1_13_in24 = reg_0608;
    57: op1_13_in24 = reg_0085;
    58: op1_13_in24 = reg_0520;
    59: op1_13_in24 = reg_0799;
    60: op1_13_in24 = reg_0482;
    61: op1_13_in24 = reg_0937;
    62: op1_13_in24 = reg_0406;
    63: op1_13_in24 = imem01_in[107:104];
    64: op1_13_in24 = imem01_in[59:56];
    65: op1_13_in24 = reg_0285;
    66: op1_13_in24 = reg_0867;
    67: op1_13_in24 = reg_0740;
    68: op1_13_in24 = imem06_in[119:116];
    70: op1_13_in24 = reg_0291;
    71: op1_13_in24 = reg_0154;
    72: op1_13_in24 = reg_0971;
    73: op1_13_in24 = imem03_in[47:44];
    74: op1_13_in24 = reg_1007;
    75: op1_13_in24 = reg_0912;
    76: op1_13_in24 = imem06_in[3:0];
    78: op1_13_in24 = imem01_in[27:24];
    79: op1_13_in24 = imem01_in[23:20];
    80: op1_13_in24 = imem03_in[59:56];
    81: op1_13_in24 = reg_0276;
    82: op1_13_in24 = reg_0607;
    84: op1_13_in24 = reg_0805;
    85: op1_13_in24 = imem02_in[115:112];
    86: op1_13_in24 = imem03_in[39:36];
    88: op1_13_in24 = reg_0365;
    91: op1_13_in24 = imem01_in[35:32];
    92: op1_13_in24 = reg_0215;
    93: op1_13_in24 = imem07_in[31:28];
    94: op1_13_in24 = imem07_in[71:68];
    95: op1_13_in24 = reg_0651;
    96: op1_13_in24 = reg_0657;
    default: op1_13_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv24 = 1;
    10: op1_13_inv24 = 1;
    15: op1_13_inv24 = 1;
    16: op1_13_inv24 = 1;
    17: op1_13_inv24 = 1;
    23: op1_13_inv24 = 1;
    24: op1_13_inv24 = 1;
    25: op1_13_inv24 = 1;
    26: op1_13_inv24 = 1;
    27: op1_13_inv24 = 1;
    28: op1_13_inv24 = 1;
    29: op1_13_inv24 = 1;
    32: op1_13_inv24 = 1;
    33: op1_13_inv24 = 1;
    34: op1_13_inv24 = 1;
    36: op1_13_inv24 = 1;
    37: op1_13_inv24 = 1;
    38: op1_13_inv24 = 1;
    39: op1_13_inv24 = 1;
    42: op1_13_inv24 = 1;
    46: op1_13_inv24 = 1;
    52: op1_13_inv24 = 1;
    55: op1_13_inv24 = 1;
    57: op1_13_inv24 = 1;
    60: op1_13_inv24 = 1;
    63: op1_13_inv24 = 1;
    65: op1_13_inv24 = 1;
    72: op1_13_inv24 = 1;
    74: op1_13_inv24 = 1;
    78: op1_13_inv24 = 1;
    79: op1_13_inv24 = 1;
    81: op1_13_inv24 = 1;
    86: op1_13_inv24 = 1;
    88: op1_13_inv24 = 1;
    92: op1_13_inv24 = 1;
    93: op1_13_inv24 = 1;
    94: op1_13_inv24 = 1;
    95: op1_13_inv24 = 1;
    default: op1_13_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in25 = reg_0710;
    6: op1_13_in25 = reg_0215;
    7: op1_13_in25 = reg_0236;
    8: op1_13_in25 = imem03_in[15:12];
    9: op1_13_in25 = reg_0725;
    10: op1_13_in25 = reg_0946;
    11: op1_13_in25 = reg_0905;
    12: op1_13_in25 = imem04_in[59:56];
    13: op1_13_in25 = reg_0496;
    65: op1_13_in25 = reg_0496;
    14: op1_13_in25 = imem03_in[19:16];
    85: op1_13_in25 = imem03_in[19:16];
    15: op1_13_in25 = reg_0531;
    44: op1_13_in25 = reg_0531;
    16: op1_13_in25 = reg_0439;
    17: op1_13_in25 = reg_0869;
    19: op1_13_in25 = reg_0230;
    21: op1_13_in25 = imem02_in[55:52];
    22: op1_13_in25 = imem05_in[79:76];
    23: op1_13_in25 = reg_0425;
    24: op1_13_in25 = reg_0607;
    25: op1_13_in25 = reg_0701;
    26: op1_13_in25 = imem04_in[95:92];
    27: op1_13_in25 = imem01_in[39:36];
    28: op1_13_in25 = reg_0811;
    29: op1_13_in25 = reg_0146;
    30: op1_13_in25 = reg_0781;
    31: op1_13_in25 = reg_0360;
    32: op1_13_in25 = imem04_in[119:116];
    33: op1_13_in25 = reg_0875;
    34: op1_13_in25 = imem02_in[51:48];
    35: op1_13_in25 = imem03_in[35:32];
    36: op1_13_in25 = imem03_in[11:8];
    60: op1_13_in25 = imem03_in[11:8];
    37: op1_13_in25 = imem05_in[67:64];
    38: op1_13_in25 = reg_0997;
    39: op1_13_in25 = reg_0180;
    40: op1_13_in25 = reg_0436;
    42: op1_13_in25 = reg_0847;
    43: op1_13_in25 = reg_0942;
    45: op1_13_in25 = imem01_in[115:112];
    63: op1_13_in25 = imem01_in[115:112];
    46: op1_13_in25 = reg_0877;
    47: op1_13_in25 = reg_0612;
    48: op1_13_in25 = reg_0227;
    49: op1_13_in25 = reg_0261;
    66: op1_13_in25 = reg_0261;
    50: op1_13_in25 = reg_0904;
    52: op1_13_in25 = imem06_in[103:100];
    54: op1_13_in25 = reg_0167;
    55: op1_13_in25 = reg_0740;
    56: op1_13_in25 = reg_0516;
    57: op1_13_in25 = reg_0310;
    58: op1_13_in25 = reg_1043;
    90: op1_13_in25 = reg_1043;
    59: op1_13_in25 = reg_0067;
    61: op1_13_in25 = reg_0541;
    62: op1_13_in25 = reg_0589;
    64: op1_13_in25 = imem01_in[67:64];
    67: op1_13_in25 = reg_1017;
    68: op1_13_in25 = imem06_in[123:120];
    70: op1_13_in25 = reg_0743;
    71: op1_13_in25 = reg_0144;
    72: op1_13_in25 = reg_1024;
    73: op1_13_in25 = imem03_in[79:76];
    74: op1_13_in25 = reg_0240;
    75: op1_13_in25 = reg_0050;
    76: op1_13_in25 = imem06_in[23:20];
    78: op1_13_in25 = imem01_in[35:32];
    79: op1_13_in25 = imem01_in[27:24];
    80: op1_13_in25 = imem03_in[123:120];
    81: op1_13_in25 = reg_0584;
    82: op1_13_in25 = reg_0500;
    84: op1_13_in25 = reg_0421;
    86: op1_13_in25 = imem03_in[67:64];
    88: op1_13_in25 = reg_0894;
    91: op1_13_in25 = imem01_in[103:100];
    92: op1_13_in25 = reg_0655;
    93: op1_13_in25 = imem07_in[87:84];
    94: op1_13_in25 = imem07_in[99:96];
    95: op1_13_in25 = reg_0951;
    96: op1_13_in25 = imem06_in[3:0];
    default: op1_13_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv25 = 1;
    6: op1_13_inv25 = 1;
    8: op1_13_inv25 = 1;
    11: op1_13_inv25 = 1;
    12: op1_13_inv25 = 1;
    14: op1_13_inv25 = 1;
    19: op1_13_inv25 = 1;
    24: op1_13_inv25 = 1;
    25: op1_13_inv25 = 1;
    26: op1_13_inv25 = 1;
    27: op1_13_inv25 = 1;
    28: op1_13_inv25 = 1;
    34: op1_13_inv25 = 1;
    35: op1_13_inv25 = 1;
    36: op1_13_inv25 = 1;
    37: op1_13_inv25 = 1;
    38: op1_13_inv25 = 1;
    40: op1_13_inv25 = 1;
    42: op1_13_inv25 = 1;
    45: op1_13_inv25 = 1;
    47: op1_13_inv25 = 1;
    49: op1_13_inv25 = 1;
    50: op1_13_inv25 = 1;
    52: op1_13_inv25 = 1;
    54: op1_13_inv25 = 1;
    60: op1_13_inv25 = 1;
    61: op1_13_inv25 = 1;
    64: op1_13_inv25 = 1;
    65: op1_13_inv25 = 1;
    66: op1_13_inv25 = 1;
    72: op1_13_inv25 = 1;
    82: op1_13_inv25 = 1;
    85: op1_13_inv25 = 1;
    86: op1_13_inv25 = 1;
    90: op1_13_inv25 = 1;
    92: op1_13_inv25 = 1;
    default: op1_13_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in26 = reg_0723;
    6: op1_13_in26 = reg_0259;
    7: op1_13_in26 = reg_0248;
    8: op1_13_in26 = imem03_in[23:20];
    14: op1_13_in26 = imem03_in[23:20];
    9: op1_13_in26 = reg_0714;
    10: op1_13_in26 = reg_0268;
    11: op1_13_in26 = reg_1033;
    12: op1_13_in26 = imem04_in[63:60];
    13: op1_13_in26 = reg_0869;
    65: op1_13_in26 = reg_0869;
    15: op1_13_in26 = reg_0547;
    16: op1_13_in26 = reg_0427;
    17: op1_13_in26 = reg_1043;
    19: op1_13_in26 = reg_0885;
    21: op1_13_in26 = imem02_in[59:56];
    22: op1_13_in26 = imem05_in[83:80];
    37: op1_13_in26 = imem05_in[83:80];
    23: op1_13_in26 = reg_0424;
    24: op1_13_in26 = reg_0631;
    25: op1_13_in26 = reg_0706;
    26: op1_13_in26 = imem04_in[119:116];
    27: op1_13_in26 = imem01_in[67:64];
    28: op1_13_in26 = reg_0221;
    29: op1_13_in26 = reg_0154;
    30: op1_13_in26 = reg_1011;
    31: op1_13_in26 = reg_0568;
    32: op1_13_in26 = reg_0301;
    33: op1_13_in26 = reg_0285;
    34: op1_13_in26 = imem02_in[67:64];
    35: op1_13_in26 = imem03_in[39:36];
    36: op1_13_in26 = imem03_in[39:36];
    38: op1_13_in26 = imem04_in[83:80];
    39: op1_13_in26 = reg_0165;
    40: op1_13_in26 = reg_0434;
    42: op1_13_in26 = reg_0923;
    43: op1_13_in26 = reg_0946;
    44: op1_13_in26 = reg_0008;
    45: op1_13_in26 = reg_0779;
    46: op1_13_in26 = reg_0546;
    47: op1_13_in26 = reg_0264;
    48: op1_13_in26 = reg_0610;
    49: op1_13_in26 = reg_0016;
    50: op1_13_in26 = reg_0933;
    52: op1_13_in26 = imem06_in[119:116];
    54: op1_13_in26 = reg_0160;
    55: op1_13_in26 = reg_1017;
    56: op1_13_in26 = reg_0083;
    57: op1_13_in26 = imem03_in[11:8];
    58: op1_13_in26 = reg_0521;
    59: op1_13_in26 = reg_0074;
    60: op1_13_in26 = imem03_in[31:28];
    61: op1_13_in26 = reg_0848;
    62: op1_13_in26 = reg_0868;
    63: op1_13_in26 = imem01_in[119:116];
    64: op1_13_in26 = imem01_in[91:88];
    66: op1_13_in26 = reg_0840;
    67: op1_13_in26 = reg_0832;
    68: op1_13_in26 = reg_0696;
    70: op1_13_in26 = reg_0676;
    71: op1_13_in26 = reg_0629;
    72: op1_13_in26 = reg_0904;
    73: op1_13_in26 = reg_0006;
    74: op1_13_in26 = reg_0661;
    75: op1_13_in26 = reg_0850;
    76: op1_13_in26 = imem06_in[27:24];
    78: op1_13_in26 = imem01_in[75:72];
    79: op1_13_in26 = imem01_in[39:36];
    80: op1_13_in26 = reg_0620;
    81: op1_13_in26 = reg_0809;
    82: op1_13_in26 = reg_0902;
    84: op1_13_in26 = reg_0744;
    85: op1_13_in26 = imem03_in[99:96];
    86: op1_13_in26 = imem03_in[87:84];
    88: op1_13_in26 = reg_0874;
    90: op1_13_in26 = reg_0830;
    91: op1_13_in26 = imem01_in[111:108];
    92: op1_13_in26 = reg_0275;
    93: op1_13_in26 = imem07_in[99:96];
    94: op1_13_in26 = reg_0726;
    95: op1_13_in26 = reg_0741;
    96: op1_13_in26 = imem06_in[47:44];
    default: op1_13_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv26 = 1;
    13: op1_13_inv26 = 1;
    16: op1_13_inv26 = 1;
    17: op1_13_inv26 = 1;
    19: op1_13_inv26 = 1;
    27: op1_13_inv26 = 1;
    29: op1_13_inv26 = 1;
    30: op1_13_inv26 = 1;
    31: op1_13_inv26 = 1;
    32: op1_13_inv26 = 1;
    33: op1_13_inv26 = 1;
    34: op1_13_inv26 = 1;
    38: op1_13_inv26 = 1;
    43: op1_13_inv26 = 1;
    44: op1_13_inv26 = 1;
    45: op1_13_inv26 = 1;
    48: op1_13_inv26 = 1;
    49: op1_13_inv26 = 1;
    54: op1_13_inv26 = 1;
    55: op1_13_inv26 = 1;
    58: op1_13_inv26 = 1;
    59: op1_13_inv26 = 1;
    61: op1_13_inv26 = 1;
    62: op1_13_inv26 = 1;
    64: op1_13_inv26 = 1;
    65: op1_13_inv26 = 1;
    68: op1_13_inv26 = 1;
    70: op1_13_inv26 = 1;
    73: op1_13_inv26 = 1;
    75: op1_13_inv26 = 1;
    76: op1_13_inv26 = 1;
    78: op1_13_inv26 = 1;
    80: op1_13_inv26 = 1;
    81: op1_13_inv26 = 1;
    84: op1_13_inv26 = 1;
    90: op1_13_inv26 = 1;
    91: op1_13_inv26 = 1;
    92: op1_13_inv26 = 1;
    93: op1_13_inv26 = 1;
    default: op1_13_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in27 = reg_0724;
    6: op1_13_in27 = reg_0270;
    7: op1_13_in27 = reg_0245;
    8: op1_13_in27 = imem03_in[27:24];
    9: op1_13_in27 = reg_0701;
    10: op1_13_in27 = reg_0250;
    11: op1_13_in27 = reg_1041;
    12: op1_13_in27 = imem04_in[83:80];
    13: op1_13_in27 = reg_0885;
    14: op1_13_in27 = imem03_in[111:108];
    15: op1_13_in27 = reg_0281;
    16: op1_13_in27 = reg_0420;
    17: op1_13_in27 = reg_0830;
    19: op1_13_in27 = reg_1043;
    21: op1_13_in27 = imem02_in[67:64];
    22: op1_13_in27 = imem05_in[103:100];
    37: op1_13_in27 = imem05_in[103:100];
    23: op1_13_in27 = reg_0429;
    24: op1_13_in27 = reg_0626;
    68: op1_13_in27 = reg_0626;
    25: op1_13_in27 = reg_0424;
    26: op1_13_in27 = imem04_in[127:124];
    27: op1_13_in27 = imem01_in[71:68];
    28: op1_13_in27 = reg_0500;
    72: op1_13_in27 = reg_0500;
    29: op1_13_in27 = reg_0139;
    30: op1_13_in27 = reg_0011;
    31: op1_13_in27 = reg_0569;
    32: op1_13_in27 = reg_0530;
    33: op1_13_in27 = reg_0044;
    34: op1_13_in27 = imem02_in[83:80];
    35: op1_13_in27 = imem03_in[43:40];
    36: op1_13_in27 = imem03_in[67:64];
    38: op1_13_in27 = imem04_in[123:120];
    39: op1_13_in27 = reg_0179;
    40: op1_13_in27 = reg_0438;
    42: op1_13_in27 = reg_0040;
    43: op1_13_in27 = reg_0835;
    44: op1_13_in27 = reg_0622;
    45: op1_13_in27 = reg_0560;
    46: op1_13_in27 = reg_0579;
    47: op1_13_in27 = reg_0399;
    48: op1_13_in27 = reg_0925;
    49: op1_13_in27 = imem03_in[3:0];
    50: op1_13_in27 = reg_0592;
    52: op1_13_in27 = reg_0624;
    54: op1_13_in27 = reg_0163;
    55: op1_13_in27 = reg_0232;
    82: op1_13_in27 = reg_0232;
    56: op1_13_in27 = reg_0007;
    57: op1_13_in27 = imem03_in[15:12];
    58: op1_13_in27 = reg_0906;
    59: op1_13_in27 = imem04_in[11:8];
    60: op1_13_in27 = imem03_in[39:36];
    61: op1_13_in27 = reg_0067;
    62: op1_13_in27 = reg_0161;
    63: op1_13_in27 = reg_0933;
    64: op1_13_in27 = imem01_in[107:104];
    65: op1_13_in27 = reg_1040;
    66: op1_13_in27 = reg_0310;
    67: op1_13_in27 = reg_0860;
    70: op1_13_in27 = reg_0099;
    71: op1_13_in27 = reg_0128;
    73: op1_13_in27 = reg_0620;
    74: op1_13_in27 = reg_0038;
    75: op1_13_in27 = reg_0056;
    76: op1_13_in27 = imem06_in[63:60];
    78: op1_13_in27 = imem01_in[95:92];
    79: op1_13_in27 = reg_0122;
    80: op1_13_in27 = reg_0012;
    81: op1_13_in27 = reg_0288;
    84: op1_13_in27 = reg_0406;
    85: op1_13_in27 = reg_0535;
    86: op1_13_in27 = imem03_in[103:100];
    88: op1_13_in27 = reg_0050;
    90: op1_13_in27 = reg_1037;
    91: op1_13_in27 = imem01_in[115:112];
    92: op1_13_in27 = reg_0141;
    93: op1_13_in27 = reg_0726;
    94: op1_13_in27 = reg_0164;
    95: op1_13_in27 = imem06_in[75:72];
    96: op1_13_in27 = imem06_in[75:72];
    default: op1_13_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv27 = 1;
    8: op1_13_inv27 = 1;
    9: op1_13_inv27 = 1;
    11: op1_13_inv27 = 1;
    14: op1_13_inv27 = 1;
    15: op1_13_inv27 = 1;
    17: op1_13_inv27 = 1;
    19: op1_13_inv27 = 1;
    21: op1_13_inv27 = 1;
    22: op1_13_inv27 = 1;
    24: op1_13_inv27 = 1;
    25: op1_13_inv27 = 1;
    30: op1_13_inv27 = 1;
    31: op1_13_inv27 = 1;
    33: op1_13_inv27 = 1;
    34: op1_13_inv27 = 1;
    36: op1_13_inv27 = 1;
    37: op1_13_inv27 = 1;
    38: op1_13_inv27 = 1;
    42: op1_13_inv27 = 1;
    43: op1_13_inv27 = 1;
    44: op1_13_inv27 = 1;
    45: op1_13_inv27 = 1;
    47: op1_13_inv27 = 1;
    48: op1_13_inv27 = 1;
    49: op1_13_inv27 = 1;
    54: op1_13_inv27 = 1;
    56: op1_13_inv27 = 1;
    57: op1_13_inv27 = 1;
    59: op1_13_inv27 = 1;
    60: op1_13_inv27 = 1;
    63: op1_13_inv27 = 1;
    65: op1_13_inv27 = 1;
    66: op1_13_inv27 = 1;
    68: op1_13_inv27 = 1;
    72: op1_13_inv27 = 1;
    73: op1_13_inv27 = 1;
    78: op1_13_inv27 = 1;
    82: op1_13_inv27 = 1;
    84: op1_13_inv27 = 1;
    85: op1_13_inv27 = 1;
    86: op1_13_inv27 = 1;
    88: op1_13_inv27 = 1;
    90: op1_13_inv27 = 1;
    93: op1_13_inv27 = 1;
    94: op1_13_inv27 = 1;
    95: op1_13_inv27 = 1;
    96: op1_13_inv27 = 1;
    default: op1_13_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in28 = reg_0707;
    6: op1_13_in28 = reg_0253;
    10: op1_13_in28 = reg_0253;
    7: op1_13_in28 = reg_0238;
    8: op1_13_in28 = imem03_in[51:48];
    9: op1_13_in28 = reg_0422;
    11: op1_13_in28 = reg_1038;
    12: op1_13_in28 = imem04_in[87:84];
    13: op1_13_in28 = reg_0830;
    14: op1_13_in28 = imem03_in[123:120];
    15: op1_13_in28 = reg_0295;
    16: op1_13_in28 = reg_0169;
    62: op1_13_in28 = reg_0169;
    17: op1_13_in28 = reg_1037;
    19: op1_13_in28 = reg_1044;
    21: op1_13_in28 = imem02_in[83:80];
    22: op1_13_in28 = imem05_in[111:108];
    23: op1_13_in28 = reg_0434;
    24: op1_13_in28 = reg_0615;
    25: op1_13_in28 = reg_0436;
    26: op1_13_in28 = reg_1006;
    46: op1_13_in28 = reg_1006;
    27: op1_13_in28 = imem01_in[111:108];
    28: op1_13_in28 = reg_0118;
    29: op1_13_in28 = reg_0153;
    30: op1_13_in28 = imem07_in[23:20];
    31: op1_13_in28 = reg_0532;
    32: op1_13_in28 = reg_0292;
    33: op1_13_in28 = imem05_in[31:28];
    34: op1_13_in28 = imem02_in[107:104];
    35: op1_13_in28 = imem03_in[47:44];
    60: op1_13_in28 = imem03_in[47:44];
    36: op1_13_in28 = imem03_in[79:76];
    37: op1_13_in28 = reg_0962;
    38: op1_13_in28 = imem04_in[127:124];
    39: op1_13_in28 = reg_0166;
    40: op1_13_in28 = reg_0448;
    42: op1_13_in28 = reg_0373;
    43: op1_13_in28 = reg_0816;
    44: op1_13_in28 = imem07_in[35:32];
    45: op1_13_in28 = reg_0218;
    47: op1_13_in28 = reg_0390;
    48: op1_13_in28 = reg_0906;
    49: op1_13_in28 = imem03_in[39:36];
    50: op1_13_in28 = reg_0216;
    72: op1_13_in28 = reg_0216;
    52: op1_13_in28 = reg_0220;
    54: op1_13_in28 = reg_0178;
    55: op1_13_in28 = reg_0003;
    56: op1_13_in28 = reg_0761;
    57: op1_13_in28 = imem03_in[31:28];
    58: op1_13_in28 = reg_1055;
    59: op1_13_in28 = imem04_in[67:64];
    61: op1_13_in28 = reg_0072;
    63: op1_13_in28 = reg_0503;
    64: op1_13_in28 = imem01_in[127:124];
    65: op1_13_in28 = reg_1041;
    66: op1_13_in28 = reg_0884;
    67: op1_13_in28 = reg_0821;
    68: op1_13_in28 = reg_0384;
    70: op1_13_in28 = reg_0245;
    71: op1_13_in28 = reg_0510;
    73: op1_13_in28 = reg_0345;
    74: op1_13_in28 = reg_0376;
    75: op1_13_in28 = reg_0809;
    76: op1_13_in28 = imem06_in[95:92];
    78: op1_13_in28 = imem01_in[107:104];
    79: op1_13_in28 = reg_1042;
    80: op1_13_in28 = reg_0445;
    81: op1_13_in28 = reg_0893;
    82: op1_13_in28 = reg_0769;
    84: op1_13_in28 = reg_0350;
    85: op1_13_in28 = reg_0585;
    86: op1_13_in28 = imem03_in[107:104];
    88: op1_13_in28 = reg_0574;
    90: op1_13_in28 = reg_0832;
    91: op1_13_in28 = reg_0488;
    92: op1_13_in28 = reg_0947;
    93: op1_13_in28 = reg_0374;
    94: op1_13_in28 = reg_0442;
    95: op1_13_in28 = imem06_in[123:120];
    96: op1_13_in28 = imem06_in[127:124];
    default: op1_13_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv28 = 1;
    8: op1_13_inv28 = 1;
    9: op1_13_inv28 = 1;
    10: op1_13_inv28 = 1;
    12: op1_13_inv28 = 1;
    13: op1_13_inv28 = 1;
    14: op1_13_inv28 = 1;
    17: op1_13_inv28 = 1;
    22: op1_13_inv28 = 1;
    25: op1_13_inv28 = 1;
    28: op1_13_inv28 = 1;
    31: op1_13_inv28 = 1;
    32: op1_13_inv28 = 1;
    33: op1_13_inv28 = 1;
    35: op1_13_inv28 = 1;
    40: op1_13_inv28 = 1;
    42: op1_13_inv28 = 1;
    47: op1_13_inv28 = 1;
    50: op1_13_inv28 = 1;
    52: op1_13_inv28 = 1;
    54: op1_13_inv28 = 1;
    60: op1_13_inv28 = 1;
    66: op1_13_inv28 = 1;
    67: op1_13_inv28 = 1;
    70: op1_13_inv28 = 1;
    71: op1_13_inv28 = 1;
    73: op1_13_inv28 = 1;
    74: op1_13_inv28 = 1;
    75: op1_13_inv28 = 1;
    76: op1_13_inv28 = 1;
    79: op1_13_inv28 = 1;
    80: op1_13_inv28 = 1;
    81: op1_13_inv28 = 1;
    82: op1_13_inv28 = 1;
    84: op1_13_inv28 = 1;
    86: op1_13_inv28 = 1;
    88: op1_13_inv28 = 1;
    90: op1_13_inv28 = 1;
    91: op1_13_inv28 = 1;
    92: op1_13_inv28 = 1;
    93: op1_13_inv28 = 1;
    94: op1_13_inv28 = 1;
    default: op1_13_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in29 = reg_0700;
    6: op1_13_in29 = reg_0263;
    7: op1_13_in29 = reg_0219;
    8: op1_13_in29 = imem03_in[75:72];
    9: op1_13_in29 = reg_0447;
    10: op1_13_in29 = reg_0147;
    11: op1_13_in29 = reg_0112;
    12: op1_13_in29 = imem04_in[99:96];
    13: op1_13_in29 = reg_1037;
    14: op1_13_in29 = reg_0586;
    15: op1_13_in29 = reg_0286;
    16: op1_13_in29 = reg_0163;
    17: op1_13_in29 = reg_1035;
    19: op1_13_in29 = reg_1033;
    21: op1_13_in29 = imem02_in[95:92];
    22: op1_13_in29 = imem05_in[115:112];
    23: op1_13_in29 = reg_0449;
    24: op1_13_in29 = reg_0406;
    25: op1_13_in29 = reg_0421;
    26: op1_13_in29 = reg_1009;
    27: op1_13_in29 = imem01_in[123:120];
    28: op1_13_in29 = reg_0119;
    29: op1_13_in29 = reg_0130;
    30: op1_13_in29 = imem07_in[47:44];
    44: op1_13_in29 = imem07_in[47:44];
    31: op1_13_in29 = imem03_in[19:16];
    32: op1_13_in29 = reg_0541;
    33: op1_13_in29 = imem05_in[75:72];
    34: op1_13_in29 = reg_0650;
    35: op1_13_in29 = imem03_in[67:64];
    36: op1_13_in29 = imem03_in[95:92];
    37: op1_13_in29 = reg_0973;
    38: op1_13_in29 = reg_0277;
    39: op1_13_in29 = reg_0164;
    40: op1_13_in29 = reg_0431;
    42: op1_13_in29 = reg_0509;
    43: op1_13_in29 = reg_0149;
    45: op1_13_in29 = reg_0299;
    46: op1_13_in29 = reg_0055;
    47: op1_13_in29 = reg_0594;
    48: op1_13_in29 = reg_0105;
    49: op1_13_in29 = imem03_in[43:40];
    50: op1_13_in29 = reg_0737;
    52: op1_13_in29 = reg_0611;
    54: op1_13_in29 = reg_0158;
    55: op1_13_in29 = reg_1053;
    56: op1_13_in29 = reg_0084;
    57: op1_13_in29 = imem03_in[39:36];
    58: op1_13_in29 = reg_0003;
    82: op1_13_in29 = reg_0003;
    59: op1_13_in29 = imem04_in[95:92];
    60: op1_13_in29 = imem03_in[51:48];
    61: op1_13_in29 = reg_0284;
    62: op1_13_in29 = reg_0166;
    63: op1_13_in29 = reg_0249;
    64: op1_13_in29 = reg_0762;
    65: op1_13_in29 = reg_1017;
    66: op1_13_in29 = imem03_in[27:24];
    67: op1_13_in29 = imem02_in[7:4];
    68: op1_13_in29 = reg_0692;
    70: op1_13_in29 = reg_0327;
    71: op1_13_in29 = reg_1021;
    72: op1_13_in29 = reg_0232;
    73: op1_13_in29 = reg_0681;
    74: op1_13_in29 = reg_1002;
    75: op1_13_in29 = reg_0061;
    76: op1_13_in29 = reg_0010;
    78: op1_13_in29 = imem01_in[111:108];
    79: op1_13_in29 = reg_0106;
    80: op1_13_in29 = reg_0298;
    81: op1_13_in29 = reg_0041;
    84: op1_13_in29 = reg_0172;
    85: op1_13_in29 = reg_0046;
    86: op1_13_in29 = reg_0060;
    88: op1_13_in29 = reg_0576;
    90: op1_13_in29 = reg_0283;
    91: op1_13_in29 = reg_1039;
    92: op1_13_in29 = reg_0964;
    93: op1_13_in29 = reg_0805;
    94: op1_13_in29 = reg_0563;
    95: op1_13_in29 = reg_1018;
    96: op1_13_in29 = reg_0660;
    default: op1_13_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv29 = 1;
    8: op1_13_inv29 = 1;
    9: op1_13_inv29 = 1;
    10: op1_13_inv29 = 1;
    11: op1_13_inv29 = 1;
    12: op1_13_inv29 = 1;
    13: op1_13_inv29 = 1;
    19: op1_13_inv29 = 1;
    21: op1_13_inv29 = 1;
    24: op1_13_inv29 = 1;
    25: op1_13_inv29 = 1;
    28: op1_13_inv29 = 1;
    30: op1_13_inv29 = 1;
    31: op1_13_inv29 = 1;
    32: op1_13_inv29 = 1;
    33: op1_13_inv29 = 1;
    34: op1_13_inv29 = 1;
    37: op1_13_inv29 = 1;
    38: op1_13_inv29 = 1;
    39: op1_13_inv29 = 1;
    46: op1_13_inv29 = 1;
    47: op1_13_inv29 = 1;
    48: op1_13_inv29 = 1;
    50: op1_13_inv29 = 1;
    55: op1_13_inv29 = 1;
    56: op1_13_inv29 = 1;
    58: op1_13_inv29 = 1;
    62: op1_13_inv29 = 1;
    64: op1_13_inv29 = 1;
    67: op1_13_inv29 = 1;
    68: op1_13_inv29 = 1;
    70: op1_13_inv29 = 1;
    71: op1_13_inv29 = 1;
    72: op1_13_inv29 = 1;
    73: op1_13_inv29 = 1;
    74: op1_13_inv29 = 1;
    78: op1_13_inv29 = 1;
    79: op1_13_inv29 = 1;
    80: op1_13_inv29 = 1;
    84: op1_13_inv29 = 1;
    86: op1_13_inv29 = 1;
    88: op1_13_inv29 = 1;
    90: op1_13_inv29 = 1;
    91: op1_13_inv29 = 1;
    94: op1_13_inv29 = 1;
    96: op1_13_inv29 = 1;
    default: op1_13_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_13_in30 = reg_0434;
    6: op1_13_in30 = reg_0151;
    7: op1_13_in30 = reg_0225;
    8: op1_13_in30 = imem03_in[87:84];
    9: op1_13_in30 = reg_0419;
    10: op1_13_in30 = reg_0143;
    11: op1_13_in30 = reg_0115;
    12: op1_13_in30 = imem04_in[111:108];
    13: op1_13_in30 = reg_0216;
    14: op1_13_in30 = reg_0587;
    15: op1_13_in30 = reg_0298;
    16: op1_13_in30 = reg_0183;
    17: op1_13_in30 = reg_1015;
    19: op1_13_in30 = reg_1036;
    21: op1_13_in30 = imem03_in[63:60];
    49: op1_13_in30 = imem03_in[63:60];
    22: op1_13_in30 = imem05_in[119:116];
    23: op1_13_in30 = reg_0448;
    24: op1_13_in30 = reg_0367;
    25: op1_13_in30 = reg_0418;
    26: op1_13_in30 = reg_0539;
    27: op1_13_in30 = reg_0786;
    28: op1_13_in30 = reg_0108;
    29: op1_13_in30 = reg_0140;
    30: op1_13_in30 = imem07_in[55:52];
    31: op1_13_in30 = imem03_in[23:20];
    32: op1_13_in30 = reg_0067;
    33: op1_13_in30 = imem05_in[83:80];
    34: op1_13_in30 = reg_0645;
    35: op1_13_in30 = imem03_in[75:72];
    36: op1_13_in30 = imem03_in[127:124];
    37: op1_13_in30 = reg_0960;
    38: op1_13_in30 = reg_0306;
    39: op1_13_in30 = reg_0185;
    40: op1_13_in30 = reg_0174;
    42: op1_13_in30 = reg_0820;
    43: op1_13_in30 = reg_0145;
    44: op1_13_in30 = imem07_in[71:68];
    45: op1_13_in30 = reg_0810;
    46: op1_13_in30 = reg_0537;
    47: op1_13_in30 = reg_0309;
    48: op1_13_in30 = reg_0122;
    50: op1_13_in30 = reg_0616;
    52: op1_13_in30 = reg_0612;
    55: op1_13_in30 = reg_0101;
    56: op1_13_in30 = reg_0310;
    57: op1_13_in30 = imem03_in[47:44];
    58: op1_13_in30 = reg_0283;
    59: op1_13_in30 = imem04_in[103:100];
    60: op1_13_in30 = imem03_in[67:64];
    61: op1_13_in30 = reg_0444;
    62: op1_13_in30 = reg_0173;
    63: op1_13_in30 = reg_0829;
    64: op1_13_in30 = reg_0936;
    65: op1_13_in30 = reg_0304;
    66: op1_13_in30 = imem03_in[51:48];
    67: op1_13_in30 = imem02_in[11:8];
    68: op1_13_in30 = reg_0297;
    70: op1_13_in30 = reg_0590;
    71: op1_13_in30 = reg_0787;
    72: op1_13_in30 = reg_0512;
    73: op1_13_in30 = reg_0228;
    74: op1_13_in30 = reg_0995;
    75: op1_13_in30 = reg_0658;
    76: op1_13_in30 = reg_0625;
    78: op1_13_in30 = reg_0487;
    79: op1_13_in30 = reg_1044;
    80: op1_13_in30 = reg_0396;
    85: op1_13_in30 = reg_0396;
    81: op1_13_in30 = reg_0065;
    82: op1_13_in30 = reg_0273;
    84: op1_13_in30 = reg_0429;
    86: op1_13_in30 = reg_0535;
    88: op1_13_in30 = imem03_in[31:28];
    90: op1_13_in30 = reg_0821;
    91: op1_13_in30 = reg_0610;
    92: op1_13_in30 = reg_0436;
    93: op1_13_in30 = reg_0303;
    94: op1_13_in30 = reg_0759;
    95: op1_13_in30 = reg_0393;
    96: op1_13_in30 = reg_0080;
    default: op1_13_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv30 = 1;
    8: op1_13_inv30 = 1;
    9: op1_13_inv30 = 1;
    10: op1_13_inv30 = 1;
    12: op1_13_inv30 = 1;
    13: op1_13_inv30 = 1;
    14: op1_13_inv30 = 1;
    17: op1_13_inv30 = 1;
    19: op1_13_inv30 = 1;
    21: op1_13_inv30 = 1;
    22: op1_13_inv30 = 1;
    24: op1_13_inv30 = 1;
    25: op1_13_inv30 = 1;
    26: op1_13_inv30 = 1;
    27: op1_13_inv30 = 1;
    29: op1_13_inv30 = 1;
    30: op1_13_inv30 = 1;
    32: op1_13_inv30 = 1;
    34: op1_13_inv30 = 1;
    35: op1_13_inv30 = 1;
    38: op1_13_inv30 = 1;
    39: op1_13_inv30 = 1;
    40: op1_13_inv30 = 1;
    43: op1_13_inv30 = 1;
    44: op1_13_inv30 = 1;
    45: op1_13_inv30 = 1;
    47: op1_13_inv30 = 1;
    48: op1_13_inv30 = 1;
    59: op1_13_inv30 = 1;
    60: op1_13_inv30 = 1;
    63: op1_13_inv30 = 1;
    65: op1_13_inv30 = 1;
    66: op1_13_inv30 = 1;
    68: op1_13_inv30 = 1;
    73: op1_13_inv30 = 1;
    75: op1_13_inv30 = 1;
    76: op1_13_inv30 = 1;
    78: op1_13_inv30 = 1;
    80: op1_13_inv30 = 1;
    81: op1_13_inv30 = 1;
    82: op1_13_inv30 = 1;
    84: op1_13_inv30 = 1;
    85: op1_13_inv30 = 1;
    86: op1_13_inv30 = 1;
    88: op1_13_inv30 = 1;
    90: op1_13_inv30 = 1;
    92: op1_13_inv30 = 1;
    93: op1_13_inv30 = 1;
    default: op1_13_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_13_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_13_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in00 = imem00_in[3:0];
    20: op1_14_in00 = imem00_in[3:0];
    23: op1_14_in00 = imem00_in[3:0];
    77: op1_14_in00 = imem00_in[3:0];
    6: op1_14_in00 = reg_0142;
    7: op1_14_in00 = reg_0112;
    58: op1_14_in00 = reg_0112;
    82: op1_14_in00 = reg_0112;
    8: op1_14_in00 = imem03_in[103:100];
    9: op1_14_in00 = imem00_in[7:4];
    83: op1_14_in00 = imem00_in[7:4];
    10: op1_14_in00 = reg_0130;
    11: op1_14_in00 = reg_0117;
    12: op1_14_in00 = imem04_in[119:116];
    13: op1_14_in00 = reg_1038;
    14: op1_14_in00 = reg_0591;
    15: op1_14_in00 = reg_0061;
    16: op1_14_in00 = imem00_in[27:24];
    17: op1_14_in00 = reg_1041;
    18: op1_14_in00 = imem00_in[23:20];
    19: op1_14_in00 = reg_1015;
    21: op1_14_in00 = imem03_in[99:96];
    22: op1_14_in00 = reg_0955;
    24: op1_14_in00 = reg_1029;
    25: op1_14_in00 = imem00_in[39:36];
    87: op1_14_in00 = imem00_in[39:36];
    26: op1_14_in00 = reg_1057;
    27: op1_14_in00 = reg_0224;
    4: op1_14_in00 = imem07_in[95:92];
    2: op1_14_in00 = imem07_in[95:92];
    28: op1_14_in00 = reg_0114;
    29: op1_14_in00 = reg_0131;
    30: op1_14_in00 = imem00_in[79:76];
    31: op1_14_in00 = imem03_in[67:64];
    66: op1_14_in00 = imem03_in[67:64];
    32: op1_14_in00 = reg_0068;
    33: op1_14_in00 = imem05_in[119:116];
    3: op1_14_in00 = imem07_in[15:12];
    34: op1_14_in00 = reg_0662;
    80: op1_14_in00 = reg_0662;
    35: op1_14_in00 = imem03_in[111:108];
    36: op1_14_in00 = reg_1019;
    37: op1_14_in00 = reg_0821;
    38: op1_14_in00 = reg_0733;
    39: op1_14_in00 = reg_0157;
    40: op1_14_in00 = reg_0175;
    41: op1_14_in00 = imem00_in[11:8];
    53: op1_14_in00 = imem00_in[11:8];
    54: op1_14_in00 = imem00_in[11:8];
    42: op1_14_in00 = reg_0985;
    43: op1_14_in00 = reg_0139;
    44: op1_14_in00 = imem07_in[79:76];
    45: op1_14_in00 = reg_0247;
    46: op1_14_in00 = reg_0067;
    47: op1_14_in00 = reg_0017;
    48: op1_14_in00 = reg_0111;
    49: op1_14_in00 = imem03_in[95:92];
    50: op1_14_in00 = reg_0610;
    51: op1_14_in00 = imem00_in[35:32];
    52: op1_14_in00 = reg_0381;
    55: op1_14_in00 = reg_0109;
    56: op1_14_in00 = imem03_in[11:8];
    57: op1_14_in00 = imem03_in[59:56];
    59: op1_14_in00 = imem05_in[11:8];
    60: op1_14_in00 = imem03_in[83:80];
    61: op1_14_in00 = reg_0552;
    62: op1_14_in00 = reg_0171;
    63: op1_14_in00 = reg_0830;
    64: op1_14_in00 = reg_0218;
    65: op1_14_in00 = reg_0832;
    67: op1_14_in00 = imem02_in[15:12];
    68: op1_14_in00 = reg_0395;
    69: op1_14_in00 = imem00_in[19:16];
    70: op1_14_in00 = imem03_in[3:0];
    71: op1_14_in00 = reg_0215;
    72: op1_14_in00 = reg_0116;
    73: op1_14_in00 = reg_0307;
    74: op1_14_in00 = reg_0989;
    75: op1_14_in00 = reg_0517;
    76: op1_14_in00 = reg_0344;
    78: op1_14_in00 = reg_0904;
    79: op1_14_in00 = reg_1031;
    81: op1_14_in00 = reg_0027;
    84: op1_14_in00 = reg_0701;
    85: op1_14_in00 = reg_0590;
    86: op1_14_in00 = reg_0012;
    88: op1_14_in00 = imem03_in[39:36];
    89: op1_14_in00 = imem00_in[55:52];
    90: op1_14_in00 = imem02_in[35:32];
    91: op1_14_in00 = reg_1033;
    92: op1_14_in00 = reg_0330;
    93: op1_14_in00 = reg_0421;
    94: op1_14_in00 = reg_0433;
    95: op1_14_in00 = reg_0021;
    96: op1_14_in00 = reg_0625;
    default: op1_14_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv00 = 1;
    10: op1_14_inv00 = 1;
    11: op1_14_inv00 = 1;
    13: op1_14_inv00 = 1;
    16: op1_14_inv00 = 1;
    17: op1_14_inv00 = 1;
    19: op1_14_inv00 = 1;
    21: op1_14_inv00 = 1;
    23: op1_14_inv00 = 1;
    24: op1_14_inv00 = 1;
    4: op1_14_inv00 = 1;
    28: op1_14_inv00 = 1;
    29: op1_14_inv00 = 1;
    32: op1_14_inv00 = 1;
    33: op1_14_inv00 = 1;
    34: op1_14_inv00 = 1;
    37: op1_14_inv00 = 1;
    38: op1_14_inv00 = 1;
    40: op1_14_inv00 = 1;
    44: op1_14_inv00 = 1;
    46: op1_14_inv00 = 1;
    48: op1_14_inv00 = 1;
    50: op1_14_inv00 = 1;
    53: op1_14_inv00 = 1;
    55: op1_14_inv00 = 1;
    58: op1_14_inv00 = 1;
    63: op1_14_inv00 = 1;
    65: op1_14_inv00 = 1;
    68: op1_14_inv00 = 1;
    70: op1_14_inv00 = 1;
    71: op1_14_inv00 = 1;
    74: op1_14_inv00 = 1;
    75: op1_14_inv00 = 1;
    76: op1_14_inv00 = 1;
    78: op1_14_inv00 = 1;
    83: op1_14_inv00 = 1;
    84: op1_14_inv00 = 1;
    85: op1_14_inv00 = 1;
    88: op1_14_inv00 = 1;
    89: op1_14_inv00 = 1;
    90: op1_14_inv00 = 1;
    92: op1_14_inv00 = 1;
    93: op1_14_inv00 = 1;
    94: op1_14_inv00 = 1;
    95: op1_14_inv00 = 1;
    96: op1_14_inv00 = 1;
    default: op1_14_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in01 = imem00_in[55:52];
    6: op1_14_in01 = reg_0141;
    7: op1_14_in01 = reg_0109;
    8: op1_14_in01 = imem03_in[119:116];
    9: op1_14_in01 = imem00_in[47:44];
    23: op1_14_in01 = imem00_in[47:44];
    10: op1_14_in01 = imem06_in[3:0];
    43: op1_14_in01 = imem06_in[3:0];
    11: op1_14_in01 = reg_0113;
    12: op1_14_in01 = reg_0545;
    13: op1_14_in01 = reg_0105;
    14: op1_14_in01 = reg_0563;
    15: op1_14_in01 = reg_0075;
    16: op1_14_in01 = imem00_in[31:28];
    17: op1_14_in01 = reg_1018;
    18: op1_14_in01 = imem00_in[51:48];
    51: op1_14_in01 = imem00_in[51:48];
    19: op1_14_in01 = reg_0871;
    20: op1_14_in01 = imem00_in[99:96];
    21: op1_14_in01 = reg_0573;
    22: op1_14_in01 = reg_0956;
    24: op1_14_in01 = reg_0027;
    25: op1_14_in01 = imem00_in[59:56];
    26: op1_14_in01 = reg_0292;
    27: op1_14_in01 = reg_0769;
    4: op1_14_in01 = reg_0441;
    28: op1_14_in01 = imem02_in[35:32];
    29: op1_14_in01 = reg_0144;
    30: op1_14_in01 = reg_0698;
    31: op1_14_in01 = imem03_in[87:84];
    57: op1_14_in01 = imem03_in[87:84];
    32: op1_14_in01 = reg_0071;
    33: op1_14_in01 = reg_0971;
    3: op1_14_in01 = imem07_in[71:68];
    34: op1_14_in01 = reg_0837;
    35: op1_14_in01 = imem03_in[123:120];
    49: op1_14_in01 = imem03_in[123:120];
    36: op1_14_in01 = reg_0245;
    73: op1_14_in01 = reg_0245;
    37: op1_14_in01 = reg_0806;
    38: op1_14_in01 = reg_0062;
    40: op1_14_in01 = reg_0179;
    41: op1_14_in01 = imem00_in[19:16];
    42: op1_14_in01 = reg_0982;
    44: op1_14_in01 = imem07_in[95:92];
    45: op1_14_in01 = reg_0487;
    46: op1_14_in01 = reg_0015;
    47: op1_14_in01 = imem07_in[63:60];
    48: op1_14_in01 = reg_0100;
    50: op1_14_in01 = reg_1017;
    52: op1_14_in01 = reg_0391;
    53: op1_14_in01 = imem00_in[23:20];
    83: op1_14_in01 = imem00_in[23:20];
    54: op1_14_in01 = imem00_in[27:24];
    55: op1_14_in01 = reg_0117;
    91: op1_14_in01 = reg_0117;
    56: op1_14_in01 = imem03_in[27:24];
    58: op1_14_in01 = reg_0860;
    59: op1_14_in01 = imem05_in[31:28];
    60: op1_14_in01 = imem03_in[91:88];
    61: op1_14_in01 = reg_0542;
    63: op1_14_in01 = reg_0737;
    64: op1_14_in01 = reg_0242;
    65: op1_14_in01 = reg_0283;
    66: op1_14_in01 = reg_0060;
    67: op1_14_in01 = imem02_in[63:60];
    68: op1_14_in01 = reg_0613;
    69: op1_14_in01 = imem00_in[39:36];
    70: op1_14_in01 = imem03_in[15:12];
    71: op1_14_in01 = reg_0351;
    72: op1_14_in01 = reg_0733;
    74: op1_14_in01 = reg_0981;
    75: op1_14_in01 = reg_0777;
    76: op1_14_in01 = reg_0691;
    77: op1_14_in01 = imem00_in[7:4];
    78: op1_14_in01 = reg_0111;
    79: op1_14_in01 = reg_0610;
    80: op1_14_in01 = reg_0576;
    81: op1_14_in01 = reg_0517;
    82: op1_14_in01 = reg_0877;
    84: op1_14_in01 = reg_0185;
    85: op1_14_in01 = reg_0397;
    86: op1_14_in01 = reg_0760;
    87: op1_14_in01 = imem00_in[87:84];
    88: op1_14_in01 = imem03_in[43:40];
    89: op1_14_in01 = imem00_in[83:80];
    90: op1_14_in01 = reg_0844;
    92: op1_14_in01 = reg_0587;
    93: op1_14_in01 = reg_0641;
    94: op1_14_in01 = reg_0315;
    95: op1_14_in01 = reg_0817;
    96: op1_14_in01 = reg_1019;
    default: op1_14_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv01 = 1;
    7: op1_14_inv01 = 1;
    8: op1_14_inv01 = 1;
    10: op1_14_inv01 = 1;
    13: op1_14_inv01 = 1;
    14: op1_14_inv01 = 1;
    16: op1_14_inv01 = 1;
    17: op1_14_inv01 = 1;
    19: op1_14_inv01 = 1;
    26: op1_14_inv01 = 1;
    27: op1_14_inv01 = 1;
    28: op1_14_inv01 = 1;
    29: op1_14_inv01 = 1;
    32: op1_14_inv01 = 1;
    34: op1_14_inv01 = 1;
    35: op1_14_inv01 = 1;
    36: op1_14_inv01 = 1;
    37: op1_14_inv01 = 1;
    38: op1_14_inv01 = 1;
    40: op1_14_inv01 = 1;
    44: op1_14_inv01 = 1;
    45: op1_14_inv01 = 1;
    47: op1_14_inv01 = 1;
    48: op1_14_inv01 = 1;
    51: op1_14_inv01 = 1;
    52: op1_14_inv01 = 1;
    53: op1_14_inv01 = 1;
    54: op1_14_inv01 = 1;
    56: op1_14_inv01 = 1;
    57: op1_14_inv01 = 1;
    59: op1_14_inv01 = 1;
    60: op1_14_inv01 = 1;
    61: op1_14_inv01 = 1;
    66: op1_14_inv01 = 1;
    67: op1_14_inv01 = 1;
    70: op1_14_inv01 = 1;
    71: op1_14_inv01 = 1;
    72: op1_14_inv01 = 1;
    73: op1_14_inv01 = 1;
    74: op1_14_inv01 = 1;
    78: op1_14_inv01 = 1;
    81: op1_14_inv01 = 1;
    83: op1_14_inv01 = 1;
    86: op1_14_inv01 = 1;
    90: op1_14_inv01 = 1;
    94: op1_14_inv01 = 1;
    95: op1_14_inv01 = 1;
    default: op1_14_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in02 = imem00_in[91:88];
    51: op1_14_in02 = imem00_in[91:88];
    87: op1_14_in02 = imem00_in[91:88];
    89: op1_14_in02 = imem00_in[91:88];
    6: op1_14_in02 = reg_0137;
    7: op1_14_in02 = imem02_in[7:4];
    8: op1_14_in02 = reg_0586;
    9: op1_14_in02 = imem00_in[51:48];
    10: op1_14_in02 = imem06_in[7:4];
    11: op1_14_in02 = imem02_in[19:16];
    55: op1_14_in02 = imem02_in[19:16];
    12: op1_14_in02 = reg_0557;
    13: op1_14_in02 = reg_0124;
    14: op1_14_in02 = reg_0373;
    15: op1_14_in02 = imem05_in[43:40];
    16: op1_14_in02 = imem00_in[43:40];
    17: op1_14_in02 = reg_0102;
    18: op1_14_in02 = imem00_in[95:92];
    19: op1_14_in02 = reg_0105;
    20: op1_14_in02 = imem00_in[103:100];
    21: op1_14_in02 = reg_0583;
    22: op1_14_in02 = reg_0957;
    23: op1_14_in02 = imem00_in[87:84];
    24: op1_14_in02 = reg_0801;
    25: op1_14_in02 = imem00_in[83:80];
    26: op1_14_in02 = reg_0540;
    27: op1_14_in02 = reg_0496;
    4: op1_14_in02 = reg_0419;
    28: op1_14_in02 = imem02_in[47:44];
    29: op1_14_in02 = reg_0800;
    30: op1_14_in02 = reg_0690;
    31: op1_14_in02 = imem03_in[103:100];
    32: op1_14_in02 = reg_0063;
    33: op1_14_in02 = reg_0972;
    92: op1_14_in02 = reg_0972;
    3: op1_14_in02 = imem07_in[87:84];
    34: op1_14_in02 = reg_0334;
    35: op1_14_in02 = reg_0317;
    36: op1_14_in02 = reg_0327;
    73: op1_14_in02 = reg_0327;
    37: op1_14_in02 = reg_0244;
    96: op1_14_in02 = reg_0244;
    38: op1_14_in02 = reg_0066;
    40: op1_14_in02 = reg_0162;
    41: op1_14_in02 = imem00_in[67:64];
    42: op1_14_in02 = reg_0990;
    43: op1_14_in02 = imem06_in[59:56];
    44: op1_14_in02 = imem07_in[107:104];
    47: op1_14_in02 = imem07_in[107:104];
    45: op1_14_in02 = reg_0798;
    46: op1_14_in02 = reg_0288;
    48: op1_14_in02 = reg_0115;
    49: op1_14_in02 = imem03_in[127:124];
    50: op1_14_in02 = reg_0925;
    63: op1_14_in02 = reg_0925;
    52: op1_14_in02 = reg_0264;
    53: op1_14_in02 = imem00_in[35:32];
    54: op1_14_in02 = imem00_in[39:36];
    56: op1_14_in02 = imem03_in[55:52];
    57: op1_14_in02 = imem03_in[91:88];
    58: op1_14_in02 = imem02_in[15:12];
    59: op1_14_in02 = imem05_in[55:52];
    60: op1_14_in02 = imem03_in[107:104];
    61: op1_14_in02 = reg_0531;
    64: op1_14_in02 = reg_0919;
    65: op1_14_in02 = reg_0555;
    66: op1_14_in02 = reg_0760;
    67: op1_14_in02 = imem02_in[103:100];
    68: op1_14_in02 = reg_0698;
    69: op1_14_in02 = imem00_in[55:52];
    70: op1_14_in02 = imem03_in[39:36];
    71: op1_14_in02 = reg_0393;
    72: op1_14_in02 = reg_0109;
    74: op1_14_in02 = reg_0988;
    75: op1_14_in02 = reg_0044;
    76: op1_14_in02 = reg_0391;
    77: op1_14_in02 = imem00_in[27:24];
    78: op1_14_in02 = reg_0827;
    79: op1_14_in02 = reg_0111;
    80: op1_14_in02 = reg_0238;
    81: op1_14_in02 = reg_0108;
    82: op1_14_in02 = reg_0110;
    83: op1_14_in02 = imem00_in[31:28];
    85: op1_14_in02 = reg_0281;
    86: op1_14_in02 = reg_0228;
    88: op1_14_in02 = imem03_in[79:76];
    90: op1_14_in02 = reg_0605;
    91: op1_14_in02 = imem02_in[23:20];
    93: op1_14_in02 = reg_0868;
    94: op1_14_in02 = reg_0429;
    95: op1_14_in02 = reg_0926;
    default: op1_14_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_14_inv02 = 1;
    9: op1_14_inv02 = 1;
    11: op1_14_inv02 = 1;
    12: op1_14_inv02 = 1;
    13: op1_14_inv02 = 1;
    14: op1_14_inv02 = 1;
    16: op1_14_inv02 = 1;
    17: op1_14_inv02 = 1;
    18: op1_14_inv02 = 1;
    19: op1_14_inv02 = 1;
    20: op1_14_inv02 = 1;
    22: op1_14_inv02 = 1;
    23: op1_14_inv02 = 1;
    26: op1_14_inv02 = 1;
    27: op1_14_inv02 = 1;
    4: op1_14_inv02 = 1;
    28: op1_14_inv02 = 1;
    30: op1_14_inv02 = 1;
    31: op1_14_inv02 = 1;
    32: op1_14_inv02 = 1;
    3: op1_14_inv02 = 1;
    36: op1_14_inv02 = 1;
    38: op1_14_inv02 = 1;
    41: op1_14_inv02 = 1;
    42: op1_14_inv02 = 1;
    43: op1_14_inv02 = 1;
    45: op1_14_inv02 = 1;
    46: op1_14_inv02 = 1;
    47: op1_14_inv02 = 1;
    50: op1_14_inv02 = 1;
    52: op1_14_inv02 = 1;
    54: op1_14_inv02 = 1;
    55: op1_14_inv02 = 1;
    57: op1_14_inv02 = 1;
    59: op1_14_inv02 = 1;
    60: op1_14_inv02 = 1;
    61: op1_14_inv02 = 1;
    63: op1_14_inv02 = 1;
    65: op1_14_inv02 = 1;
    66: op1_14_inv02 = 1;
    67: op1_14_inv02 = 1;
    68: op1_14_inv02 = 1;
    72: op1_14_inv02 = 1;
    73: op1_14_inv02 = 1;
    74: op1_14_inv02 = 1;
    77: op1_14_inv02 = 1;
    78: op1_14_inv02 = 1;
    80: op1_14_inv02 = 1;
    82: op1_14_inv02 = 1;
    83: op1_14_inv02 = 1;
    85: op1_14_inv02 = 1;
    86: op1_14_inv02 = 1;
    90: op1_14_inv02 = 1;
    91: op1_14_inv02 = 1;
    92: op1_14_inv02 = 1;
    94: op1_14_inv02 = 1;
    default: op1_14_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in03 = reg_0670;
    6: op1_14_in03 = imem06_in[35:32];
    7: op1_14_in03 = imem02_in[11:8];
    8: op1_14_in03 = reg_0573;
    49: op1_14_in03 = reg_0573;
    9: op1_14_in03 = imem00_in[55:52];
    16: op1_14_in03 = imem00_in[55:52];
    10: op1_14_in03 = imem06_in[11:8];
    11: op1_14_in03 = reg_0655;
    12: op1_14_in03 = reg_0552;
    13: op1_14_in03 = reg_0111;
    14: op1_14_in03 = reg_0322;
    15: op1_14_in03 = imem05_in[51:48];
    17: op1_14_in03 = imem02_in[39:36];
    58: op1_14_in03 = imem02_in[39:36];
    18: op1_14_in03 = reg_0684;
    19: op1_14_in03 = reg_0107;
    20: op1_14_in03 = imem00_in[127:124];
    21: op1_14_in03 = reg_0568;
    22: op1_14_in03 = reg_0969;
    23: op1_14_in03 = reg_0695;
    24: op1_14_in03 = reg_1010;
    25: op1_14_in03 = imem00_in[99:96];
    51: op1_14_in03 = imem00_in[99:96];
    26: op1_14_in03 = reg_0541;
    27: op1_14_in03 = reg_0230;
    4: op1_14_in03 = reg_0434;
    28: op1_14_in03 = imem02_in[99:96];
    29: op1_14_in03 = reg_0371;
    30: op1_14_in03 = reg_0668;
    31: op1_14_in03 = imem03_in[127:124];
    88: op1_14_in03 = imem03_in[127:124];
    32: op1_14_in03 = reg_0070;
    33: op1_14_in03 = reg_0826;
    3: op1_14_in03 = imem07_in[107:104];
    34: op1_14_in03 = reg_0097;
    35: op1_14_in03 = reg_0938;
    36: op1_14_in03 = reg_0933;
    37: op1_14_in03 = reg_0489;
    38: op1_14_in03 = reg_0075;
    40: op1_14_in03 = reg_0183;
    41: op1_14_in03 = imem00_in[75:72];
    42: op1_14_in03 = reg_1000;
    43: op1_14_in03 = imem06_in[83:80];
    44: op1_14_in03 = imem07_in[111:108];
    45: op1_14_in03 = reg_0869;
    46: op1_14_in03 = imem04_in[3:0];
    47: op1_14_in03 = imem07_in[123:120];
    48: op1_14_in03 = reg_0109;
    50: op1_14_in03 = reg_0123;
    52: op1_14_in03 = reg_0383;
    53: op1_14_in03 = imem00_in[47:44];
    54: op1_14_in03 = imem00_in[47:44];
    55: op1_14_in03 = imem02_in[27:24];
    56: op1_14_in03 = imem03_in[99:96];
    57: op1_14_in03 = reg_0012;
    59: op1_14_in03 = reg_0957;
    60: op1_14_in03 = reg_0345;
    61: op1_14_in03 = reg_0270;
    63: op1_14_in03 = reg_0906;
    64: op1_14_in03 = reg_0592;
    65: op1_14_in03 = reg_0827;
    66: op1_14_in03 = reg_1007;
    67: op1_14_in03 = imem02_in[111:108];
    68: op1_14_in03 = reg_0804;
    69: op1_14_in03 = imem00_in[71:68];
    70: op1_14_in03 = imem03_in[47:44];
    71: op1_14_in03 = reg_0895;
    72: op1_14_in03 = reg_0103;
    73: op1_14_in03 = reg_0238;
    74: op1_14_in03 = imem04_in[15:12];
    75: op1_14_in03 = imem05_in[35:32];
    76: op1_14_in03 = reg_0926;
    77: op1_14_in03 = imem00_in[35:32];
    78: op1_14_in03 = reg_0115;
    79: op1_14_in03 = reg_0745;
    80: op1_14_in03 = reg_0278;
    81: op1_14_in03 = reg_0332;
    82: op1_14_in03 = imem02_in[7:4];
    83: op1_14_in03 = imem00_in[43:40];
    85: op1_14_in03 = reg_0239;
    86: op1_14_in03 = reg_0307;
    87: op1_14_in03 = reg_0001;
    89: op1_14_in03 = imem00_in[115:112];
    90: op1_14_in03 = reg_0090;
    91: op1_14_in03 = imem02_in[35:32];
    92: op1_14_in03 = reg_0970;
    93: op1_14_in03 = reg_0339;
    94: op1_14_in03 = reg_0179;
    95: op1_14_in03 = reg_0735;
    96: op1_14_in03 = reg_0267;
    default: op1_14_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv03 = 1;
    8: op1_14_inv03 = 1;
    10: op1_14_inv03 = 1;
    13: op1_14_inv03 = 1;
    14: op1_14_inv03 = 1;
    15: op1_14_inv03 = 1;
    21: op1_14_inv03 = 1;
    22: op1_14_inv03 = 1;
    25: op1_14_inv03 = 1;
    26: op1_14_inv03 = 1;
    4: op1_14_inv03 = 1;
    28: op1_14_inv03 = 1;
    29: op1_14_inv03 = 1;
    30: op1_14_inv03 = 1;
    3: op1_14_inv03 = 1;
    34: op1_14_inv03 = 1;
    36: op1_14_inv03 = 1;
    37: op1_14_inv03 = 1;
    43: op1_14_inv03 = 1;
    44: op1_14_inv03 = 1;
    46: op1_14_inv03 = 1;
    51: op1_14_inv03 = 1;
    53: op1_14_inv03 = 1;
    56: op1_14_inv03 = 1;
    57: op1_14_inv03 = 1;
    61: op1_14_inv03 = 1;
    67: op1_14_inv03 = 1;
    68: op1_14_inv03 = 1;
    72: op1_14_inv03 = 1;
    74: op1_14_inv03 = 1;
    75: op1_14_inv03 = 1;
    76: op1_14_inv03 = 1;
    77: op1_14_inv03 = 1;
    78: op1_14_inv03 = 1;
    79: op1_14_inv03 = 1;
    86: op1_14_inv03 = 1;
    88: op1_14_inv03 = 1;
    89: op1_14_inv03 = 1;
    91: op1_14_inv03 = 1;
    92: op1_14_inv03 = 1;
    94: op1_14_inv03 = 1;
    default: op1_14_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in04 = reg_0679;
    6: op1_14_in04 = imem06_in[63:60];
    10: op1_14_in04 = imem06_in[63:60];
    7: op1_14_in04 = imem02_in[51:48];
    8: op1_14_in04 = reg_0569;
    9: op1_14_in04 = imem00_in[59:56];
    16: op1_14_in04 = imem00_in[59:56];
    11: op1_14_in04 = reg_0653;
    12: op1_14_in04 = reg_0542;
    13: op1_14_in04 = reg_0125;
    14: op1_14_in04 = reg_0376;
    15: op1_14_in04 = imem05_in[75:72];
    17: op1_14_in04 = imem02_in[43:40];
    18: op1_14_in04 = reg_0691;
    19: op1_14_in04 = imem02_in[23:20];
    20: op1_14_in04 = reg_0683;
    21: op1_14_in04 = reg_0370;
    22: op1_14_in04 = reg_0942;
    23: op1_14_in04 = reg_0690;
    24: op1_14_in04 = reg_0805;
    25: op1_14_in04 = imem00_in[123:120];
    26: op1_14_in04 = reg_0062;
    27: op1_14_in04 = reg_0830;
    4: op1_14_in04 = reg_0444;
    28: op1_14_in04 = imem02_in[103:100];
    29: op1_14_in04 = reg_0754;
    30: op1_14_in04 = reg_0675;
    31: op1_14_in04 = reg_0767;
    32: op1_14_in04 = reg_0882;
    33: op1_14_in04 = reg_0813;
    3: op1_14_in04 = imem07_in[115:112];
    34: op1_14_in04 = reg_0817;
    35: op1_14_in04 = reg_1049;
    36: op1_14_in04 = reg_0398;
    37: op1_14_in04 = reg_0156;
    38: op1_14_in04 = reg_0072;
    40: op1_14_in04 = reg_0166;
    41: op1_14_in04 = imem00_in[87:84];
    54: op1_14_in04 = imem00_in[87:84];
    42: op1_14_in04 = reg_0593;
    43: op1_14_in04 = imem06_in[95:92];
    44: op1_14_in04 = reg_0720;
    45: op1_14_in04 = reg_0514;
    46: op1_14_in04 = imem04_in[43:40];
    47: op1_14_in04 = reg_0704;
    48: op1_14_in04 = imem02_in[7:4];
    49: op1_14_in04 = reg_0317;
    50: op1_14_in04 = reg_0111;
    51: op1_14_in04 = reg_0693;
    52: op1_14_in04 = reg_0390;
    53: op1_14_in04 = imem00_in[99:96];
    55: op1_14_in04 = imem02_in[47:44];
    56: op1_14_in04 = imem03_in[111:108];
    57: op1_14_in04 = reg_0099;
    58: op1_14_in04 = imem02_in[63:60];
    59: op1_14_in04 = reg_0035;
    60: op1_14_in04 = reg_0228;
    61: op1_14_in04 = reg_0490;
    63: op1_14_in04 = reg_0232;
    64: op1_14_in04 = reg_1036;
    65: op1_14_in04 = reg_0877;
    66: op1_14_in04 = reg_0245;
    67: op1_14_in04 = reg_0810;
    68: op1_14_in04 = reg_0222;
    69: op1_14_in04 = imem00_in[119:116];
    89: op1_14_in04 = imem00_in[119:116];
    70: op1_14_in04 = imem03_in[51:48];
    71: op1_14_in04 = reg_0624;
    72: op1_14_in04 = reg_0113;
    73: op1_14_in04 = reg_0579;
    80: op1_14_in04 = reg_0579;
    74: op1_14_in04 = imem04_in[19:16];
    75: op1_14_in04 = imem05_in[55:52];
    76: op1_14_in04 = reg_0028;
    77: op1_14_in04 = imem00_in[47:44];
    78: op1_14_in04 = imem02_in[31:28];
    79: op1_14_in04 = imem02_in[27:24];
    81: op1_14_in04 = reg_0856;
    82: op1_14_in04 = imem02_in[39:36];
    83: op1_14_in04 = imem00_in[63:60];
    85: op1_14_in04 = reg_1008;
    86: op1_14_in04 = reg_0434;
    87: op1_14_in04 = reg_0682;
    88: op1_14_in04 = reg_0756;
    90: op1_14_in04 = reg_0639;
    91: op1_14_in04 = imem02_in[99:96];
    92: op1_14_in04 = reg_0326;
    93: op1_14_in04 = reg_0539;
    94: op1_14_in04 = reg_0723;
    95: op1_14_in04 = reg_0384;
    96: op1_14_in04 = reg_0926;
    default: op1_14_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv04 = 1;
    6: op1_14_inv04 = 1;
    7: op1_14_inv04 = 1;
    10: op1_14_inv04 = 1;
    12: op1_14_inv04 = 1;
    13: op1_14_inv04 = 1;
    15: op1_14_inv04 = 1;
    17: op1_14_inv04 = 1;
    18: op1_14_inv04 = 1;
    19: op1_14_inv04 = 1;
    20: op1_14_inv04 = 1;
    21: op1_14_inv04 = 1;
    22: op1_14_inv04 = 1;
    25: op1_14_inv04 = 1;
    30: op1_14_inv04 = 1;
    37: op1_14_inv04 = 1;
    38: op1_14_inv04 = 1;
    40: op1_14_inv04 = 1;
    41: op1_14_inv04 = 1;
    42: op1_14_inv04 = 1;
    44: op1_14_inv04 = 1;
    46: op1_14_inv04 = 1;
    48: op1_14_inv04 = 1;
    50: op1_14_inv04 = 1;
    52: op1_14_inv04 = 1;
    55: op1_14_inv04 = 1;
    59: op1_14_inv04 = 1;
    60: op1_14_inv04 = 1;
    61: op1_14_inv04 = 1;
    63: op1_14_inv04 = 1;
    64: op1_14_inv04 = 1;
    65: op1_14_inv04 = 1;
    66: op1_14_inv04 = 1;
    69: op1_14_inv04 = 1;
    71: op1_14_inv04 = 1;
    72: op1_14_inv04 = 1;
    76: op1_14_inv04 = 1;
    77: op1_14_inv04 = 1;
    78: op1_14_inv04 = 1;
    79: op1_14_inv04 = 1;
    80: op1_14_inv04 = 1;
    82: op1_14_inv04 = 1;
    85: op1_14_inv04 = 1;
    86: op1_14_inv04 = 1;
    87: op1_14_inv04 = 1;
    88: op1_14_inv04 = 1;
    91: op1_14_inv04 = 1;
    93: op1_14_inv04 = 1;
    94: op1_14_inv04 = 1;
    95: op1_14_inv04 = 1;
    96: op1_14_inv04 = 1;
    default: op1_14_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in05 = reg_0465;
    6: op1_14_in05 = imem06_in[67:64];
    7: op1_14_in05 = imem02_in[79:76];
    8: op1_14_in05 = reg_0591;
    71: op1_14_in05 = reg_0591;
    9: op1_14_in05 = imem00_in[115:112];
    41: op1_14_in05 = imem00_in[115:112];
    10: op1_14_in05 = imem06_in[87:84];
    11: op1_14_in05 = reg_0661;
    12: op1_14_in05 = reg_0548;
    13: op1_14_in05 = reg_0116;
    50: op1_14_in05 = reg_0116;
    14: op1_14_in05 = reg_0374;
    15: op1_14_in05 = imem05_in[103:100];
    16: op1_14_in05 = imem00_in[91:88];
    17: op1_14_in05 = imem02_in[75:72];
    18: op1_14_in05 = reg_0674;
    19: op1_14_in05 = imem02_in[47:44];
    78: op1_14_in05 = imem02_in[47:44];
    20: op1_14_in05 = reg_0694;
    21: op1_14_in05 = reg_0362;
    22: op1_14_in05 = reg_0943;
    23: op1_14_in05 = reg_0481;
    24: op1_14_in05 = reg_1011;
    25: op1_14_in05 = reg_0693;
    26: op1_14_in05 = reg_0268;
    27: op1_14_in05 = reg_0871;
    4: op1_14_in05 = reg_0181;
    3: op1_14_in05 = reg_0181;
    28: op1_14_in05 = reg_0647;
    29: op1_14_in05 = reg_0545;
    30: op1_14_in05 = reg_0450;
    31: op1_14_in05 = reg_0513;
    32: op1_14_in05 = reg_0773;
    33: op1_14_in05 = reg_0816;
    34: op1_14_in05 = reg_0338;
    35: op1_14_in05 = reg_0322;
    36: op1_14_in05 = reg_0580;
    37: op1_14_in05 = reg_0130;
    38: op1_14_in05 = reg_0058;
    40: op1_14_in05 = reg_0185;
    42: op1_14_in05 = reg_0511;
    43: op1_14_in05 = reg_0220;
    44: op1_14_in05 = reg_0725;
    45: op1_14_in05 = reg_1040;
    46: op1_14_in05 = imem04_in[59:56];
    47: op1_14_in05 = reg_0730;
    48: op1_14_in05 = imem02_in[19:16];
    49: op1_14_in05 = reg_0343;
    51: op1_14_in05 = reg_0684;
    52: op1_14_in05 = reg_0380;
    53: op1_14_in05 = imem00_in[111:108];
    54: op1_14_in05 = imem00_in[107:104];
    55: op1_14_in05 = imem02_in[55:52];
    56: op1_14_in05 = reg_0572;
    57: op1_14_in05 = reg_0228;
    58: op1_14_in05 = imem02_in[115:112];
    59: op1_14_in05 = reg_0785;
    60: op1_14_in05 = reg_0445;
    61: op1_14_in05 = reg_0260;
    63: op1_14_in05 = reg_0555;
    64: op1_14_in05 = reg_0238;
    65: op1_14_in05 = imem02_in[23:20];
    66: op1_14_in05 = reg_0585;
    67: op1_14_in05 = reg_0741;
    92: op1_14_in05 = reg_0741;
    68: op1_14_in05 = reg_0605;
    69: op1_14_in05 = imem00_in[123:120];
    70: op1_14_in05 = imem03_in[99:96];
    72: op1_14_in05 = reg_0364;
    73: op1_14_in05 = reg_0040;
    74: op1_14_in05 = imem04_in[31:28];
    75: op1_14_in05 = imem05_in[59:56];
    76: op1_14_in05 = reg_0534;
    77: op1_14_in05 = imem00_in[75:72];
    79: op1_14_in05 = imem02_in[35:32];
    80: op1_14_in05 = reg_0609;
    81: op1_14_in05 = imem05_in[19:16];
    82: op1_14_in05 = imem02_in[51:48];
    83: op1_14_in05 = imem00_in[71:68];
    85: op1_14_in05 = reg_0377;
    86: op1_14_in05 = reg_0298;
    87: op1_14_in05 = reg_0685;
    88: op1_14_in05 = reg_0281;
    89: op1_14_in05 = reg_0669;
    90: op1_14_in05 = reg_0621;
    91: op1_14_in05 = reg_0536;
    93: op1_14_in05 = reg_0565;
    94: op1_14_in05 = reg_0714;
    95: op1_14_in05 = reg_0533;
    96: op1_14_in05 = reg_0328;
    default: op1_14_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv05 = 1;
    6: op1_14_inv05 = 1;
    7: op1_14_inv05 = 1;
    11: op1_14_inv05 = 1;
    12: op1_14_inv05 = 1;
    13: op1_14_inv05 = 1;
    17: op1_14_inv05 = 1;
    19: op1_14_inv05 = 1;
    21: op1_14_inv05 = 1;
    22: op1_14_inv05 = 1;
    30: op1_14_inv05 = 1;
    31: op1_14_inv05 = 1;
    32: op1_14_inv05 = 1;
    35: op1_14_inv05 = 1;
    36: op1_14_inv05 = 1;
    38: op1_14_inv05 = 1;
    40: op1_14_inv05 = 1;
    42: op1_14_inv05 = 1;
    46: op1_14_inv05 = 1;
    48: op1_14_inv05 = 1;
    49: op1_14_inv05 = 1;
    50: op1_14_inv05 = 1;
    51: op1_14_inv05 = 1;
    53: op1_14_inv05 = 1;
    54: op1_14_inv05 = 1;
    55: op1_14_inv05 = 1;
    56: op1_14_inv05 = 1;
    58: op1_14_inv05 = 1;
    59: op1_14_inv05 = 1;
    61: op1_14_inv05 = 1;
    65: op1_14_inv05 = 1;
    67: op1_14_inv05 = 1;
    70: op1_14_inv05 = 1;
    71: op1_14_inv05 = 1;
    72: op1_14_inv05 = 1;
    75: op1_14_inv05 = 1;
    79: op1_14_inv05 = 1;
    81: op1_14_inv05 = 1;
    85: op1_14_inv05 = 1;
    89: op1_14_inv05 = 1;
    91: op1_14_inv05 = 1;
    default: op1_14_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in06 = reg_0455;
    6: op1_14_in06 = imem06_in[83:80];
    7: op1_14_in06 = imem02_in[99:96];
    19: op1_14_in06 = imem02_in[99:96];
    8: op1_14_in06 = reg_0593;
    9: op1_14_in06 = imem00_in[119:116];
    10: op1_14_in06 = reg_0625;
    11: op1_14_in06 = reg_0640;
    28: op1_14_in06 = reg_0640;
    12: op1_14_in06 = reg_0549;
    13: op1_14_in06 = reg_0119;
    14: op1_14_in06 = reg_0389;
    15: op1_14_in06 = reg_0944;
    16: op1_14_in06 = imem00_in[103:100];
    17: op1_14_in06 = imem02_in[87:84];
    48: op1_14_in06 = imem02_in[87:84];
    18: op1_14_in06 = reg_0699;
    20: op1_14_in06 = reg_0676;
    21: op1_14_in06 = reg_0398;
    22: op1_14_in06 = reg_0953;
    23: op1_14_in06 = reg_0471;
    24: op1_14_in06 = reg_0798;
    25: op1_14_in06 = reg_0690;
    26: op1_14_in06 = reg_0066;
    27: op1_14_in06 = reg_1017;
    4: op1_14_in06 = reg_0182;
    29: op1_14_in06 = reg_0607;
    30: op1_14_in06 = reg_0464;
    31: op1_14_in06 = reg_0234;
    32: op1_14_in06 = reg_0286;
    33: op1_14_in06 = reg_0275;
    3: op1_14_in06 = reg_0162;
    34: op1_14_in06 = reg_0083;
    35: op1_14_in06 = reg_0046;
    36: op1_14_in06 = reg_0576;
    37: op1_14_in06 = reg_0759;
    38: op1_14_in06 = reg_0285;
    41: op1_14_in06 = imem00_in[123:120];
    42: op1_14_in06 = reg_0912;
    43: op1_14_in06 = reg_0782;
    44: op1_14_in06 = reg_0703;
    45: op1_14_in06 = reg_0906;
    46: op1_14_in06 = imem04_in[87:84];
    47: op1_14_in06 = reg_0731;
    49: op1_14_in06 = reg_1007;
    50: op1_14_in06 = reg_0104;
    51: op1_14_in06 = reg_0679;
    52: op1_14_in06 = reg_0917;
    53: op1_14_in06 = reg_0693;
    54: op1_14_in06 = reg_0695;
    55: op1_14_in06 = imem02_in[63:60];
    56: op1_14_in06 = reg_0245;
    57: op1_14_in06 = reg_0396;
    58: op1_14_in06 = reg_0363;
    59: op1_14_in06 = reg_0057;
    60: op1_14_in06 = reg_0327;
    61: op1_14_in06 = imem05_in[3:0];
    63: op1_14_in06 = reg_0120;
    64: op1_14_in06 = reg_0500;
    65: op1_14_in06 = imem02_in[35:32];
    66: op1_14_in06 = reg_0434;
    67: op1_14_in06 = reg_0336;
    68: op1_14_in06 = imem07_in[11:8];
    69: op1_14_in06 = reg_0682;
    70: op1_14_in06 = imem03_in[107:104];
    71: op1_14_in06 = reg_0863;
    72: op1_14_in06 = reg_0873;
    73: op1_14_in06 = reg_0773;
    88: op1_14_in06 = reg_0773;
    74: op1_14_in06 = imem04_in[39:36];
    75: op1_14_in06 = imem05_in[71:68];
    76: op1_14_in06 = reg_1030;
    77: op1_14_in06 = imem00_in[79:76];
    78: op1_14_in06 = imem02_in[119:116];
    79: op1_14_in06 = imem02_in[43:40];
    80: op1_14_in06 = reg_0779;
    81: op1_14_in06 = imem05_in[27:24];
    82: op1_14_in06 = imem02_in[67:64];
    83: op1_14_in06 = imem00_in[127:124];
    85: op1_14_in06 = reg_0993;
    86: op1_14_in06 = reg_0662;
    87: op1_14_in06 = reg_0684;
    89: op1_14_in06 = reg_0469;
    90: op1_14_in06 = reg_0418;
    91: op1_14_in06 = reg_0605;
    92: op1_14_in06 = imem06_in[3:0];
    93: op1_14_in06 = reg_0185;
    94: op1_14_in06 = reg_0701;
    95: op1_14_in06 = reg_0928;
    96: op1_14_in06 = reg_0754;
    default: op1_14_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv06 = 1;
    6: op1_14_inv06 = 1;
    7: op1_14_inv06 = 1;
    8: op1_14_inv06 = 1;
    15: op1_14_inv06 = 1;
    17: op1_14_inv06 = 1;
    18: op1_14_inv06 = 1;
    19: op1_14_inv06 = 1;
    20: op1_14_inv06 = 1;
    21: op1_14_inv06 = 1;
    22: op1_14_inv06 = 1;
    23: op1_14_inv06 = 1;
    26: op1_14_inv06 = 1;
    27: op1_14_inv06 = 1;
    28: op1_14_inv06 = 1;
    30: op1_14_inv06 = 1;
    31: op1_14_inv06 = 1;
    33: op1_14_inv06 = 1;
    34: op1_14_inv06 = 1;
    37: op1_14_inv06 = 1;
    38: op1_14_inv06 = 1;
    42: op1_14_inv06 = 1;
    43: op1_14_inv06 = 1;
    45: op1_14_inv06 = 1;
    46: op1_14_inv06 = 1;
    48: op1_14_inv06 = 1;
    49: op1_14_inv06 = 1;
    50: op1_14_inv06 = 1;
    52: op1_14_inv06 = 1;
    54: op1_14_inv06 = 1;
    56: op1_14_inv06 = 1;
    57: op1_14_inv06 = 1;
    61: op1_14_inv06 = 1;
    64: op1_14_inv06 = 1;
    65: op1_14_inv06 = 1;
    66: op1_14_inv06 = 1;
    67: op1_14_inv06 = 1;
    68: op1_14_inv06 = 1;
    69: op1_14_inv06 = 1;
    72: op1_14_inv06 = 1;
    74: op1_14_inv06 = 1;
    75: op1_14_inv06 = 1;
    77: op1_14_inv06 = 1;
    78: op1_14_inv06 = 1;
    79: op1_14_inv06 = 1;
    82: op1_14_inv06 = 1;
    86: op1_14_inv06 = 1;
    87: op1_14_inv06 = 1;
    89: op1_14_inv06 = 1;
    90: op1_14_inv06 = 1;
    93: op1_14_inv06 = 1;
    94: op1_14_inv06 = 1;
    default: op1_14_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in07 = reg_0475;
    6: op1_14_in07 = imem06_in[119:116];
    7: op1_14_in07 = imem02_in[115:112];
    19: op1_14_in07 = imem02_in[115:112];
    8: op1_14_in07 = reg_0384;
    9: op1_14_in07 = reg_0683;
    10: op1_14_in07 = reg_0604;
    11: op1_14_in07 = reg_0352;
    12: op1_14_in07 = reg_0546;
    13: op1_14_in07 = reg_0102;
    14: op1_14_in07 = reg_0987;
    15: op1_14_in07 = reg_0967;
    16: op1_14_in07 = imem00_in[115:112];
    17: op1_14_in07 = reg_0650;
    18: op1_14_in07 = reg_0454;
    20: op1_14_in07 = reg_0689;
    41: op1_14_in07 = reg_0689;
    53: op1_14_in07 = reg_0689;
    21: op1_14_in07 = reg_0397;
    22: op1_14_in07 = reg_0960;
    23: op1_14_in07 = reg_0479;
    24: op1_14_in07 = imem07_in[39:36];
    25: op1_14_in07 = reg_0674;
    26: op1_14_in07 = reg_0259;
    27: op1_14_in07 = reg_1018;
    4: op1_14_in07 = reg_0160;
    28: op1_14_in07 = reg_0644;
    29: op1_14_in07 = reg_0608;
    30: op1_14_in07 = reg_0477;
    31: op1_14_in07 = reg_0984;
    32: op1_14_in07 = imem05_in[3:0];
    33: op1_14_in07 = reg_0831;
    3: op1_14_in07 = reg_0159;
    34: op1_14_in07 = reg_0085;
    35: op1_14_in07 = reg_0824;
    36: op1_14_in07 = reg_0543;
    37: op1_14_in07 = reg_0486;
    38: op1_14_in07 = imem05_in[7:4];
    42: op1_14_in07 = reg_1016;
    43: op1_14_in07 = reg_0632;
    44: op1_14_in07 = reg_0705;
    45: op1_14_in07 = reg_0105;
    46: op1_14_in07 = imem05_in[47:44];
    81: op1_14_in07 = imem05_in[47:44];
    47: op1_14_in07 = reg_0725;
    48: op1_14_in07 = imem02_in[95:92];
    82: op1_14_in07 = imem02_in[95:92];
    49: op1_14_in07 = reg_0327;
    56: op1_14_in07 = reg_0327;
    50: op1_14_in07 = reg_0119;
    51: op1_14_in07 = reg_0690;
    52: op1_14_in07 = reg_0000;
    54: op1_14_in07 = reg_0697;
    94: op1_14_in07 = reg_0697;
    55: op1_14_in07 = imem02_in[79:76];
    57: op1_14_in07 = reg_0661;
    58: op1_14_in07 = reg_0657;
    59: op1_14_in07 = reg_0215;
    60: op1_14_in07 = reg_0577;
    61: op1_14_in07 = imem05_in[75:72];
    63: op1_14_in07 = reg_0364;
    64: op1_14_in07 = reg_1041;
    65: op1_14_in07 = imem02_in[43:40];
    66: op1_14_in07 = reg_0547;
    67: op1_14_in07 = reg_0279;
    68: op1_14_in07 = imem07_in[15:12];
    69: op1_14_in07 = reg_0825;
    70: op1_14_in07 = imem03_in[127:124];
    71: op1_14_in07 = reg_0222;
    72: op1_14_in07 = reg_0330;
    73: op1_14_in07 = reg_0609;
    74: op1_14_in07 = imem04_in[67:64];
    75: op1_14_in07 = imem05_in[79:76];
    76: op1_14_in07 = reg_0895;
    77: op1_14_in07 = imem00_in[91:88];
    78: op1_14_in07 = imem02_in[127:124];
    79: op1_14_in07 = imem02_in[67:64];
    80: op1_14_in07 = reg_0312;
    83: op1_14_in07 = reg_0768;
    85: op1_14_in07 = imem04_in[51:48];
    86: op1_14_in07 = reg_0823;
    87: op1_14_in07 = reg_0749;
    88: op1_14_in07 = reg_0672;
    89: op1_14_in07 = reg_0462;
    90: op1_14_in07 = reg_0837;
    91: op1_14_in07 = reg_0090;
    92: op1_14_in07 = imem06_in[59:56];
    93: op1_14_in07 = reg_0371;
    95: op1_14_in07 = reg_0783;
    96: op1_14_in07 = reg_0889;
    default: op1_14_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv07 = 1;
    6: op1_14_inv07 = 1;
    9: op1_14_inv07 = 1;
    10: op1_14_inv07 = 1;
    12: op1_14_inv07 = 1;
    15: op1_14_inv07 = 1;
    25: op1_14_inv07 = 1;
    27: op1_14_inv07 = 1;
    4: op1_14_inv07 = 1;
    30: op1_14_inv07 = 1;
    31: op1_14_inv07 = 1;
    32: op1_14_inv07 = 1;
    33: op1_14_inv07 = 1;
    3: op1_14_inv07 = 1;
    35: op1_14_inv07 = 1;
    37: op1_14_inv07 = 1;
    44: op1_14_inv07 = 1;
    46: op1_14_inv07 = 1;
    47: op1_14_inv07 = 1;
    49: op1_14_inv07 = 1;
    51: op1_14_inv07 = 1;
    55: op1_14_inv07 = 1;
    56: op1_14_inv07 = 1;
    57: op1_14_inv07 = 1;
    60: op1_14_inv07 = 1;
    72: op1_14_inv07 = 1;
    73: op1_14_inv07 = 1;
    74: op1_14_inv07 = 1;
    75: op1_14_inv07 = 1;
    77: op1_14_inv07 = 1;
    82: op1_14_inv07 = 1;
    83: op1_14_inv07 = 1;
    86: op1_14_inv07 = 1;
    87: op1_14_inv07 = 1;
    90: op1_14_inv07 = 1;
    91: op1_14_inv07 = 1;
    93: op1_14_inv07 = 1;
    94: op1_14_inv07 = 1;
    95: op1_14_inv07 = 1;
    96: op1_14_inv07 = 1;
    default: op1_14_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in08 = reg_0460;
    6: op1_14_in08 = imem06_in[123:120];
    7: op1_14_in08 = imem02_in[127:124];
    8: op1_14_in08 = reg_0362;
    9: op1_14_in08 = reg_0696;
    10: op1_14_in08 = reg_0616;
    11: op1_14_in08 = reg_0357;
    12: op1_14_in08 = reg_0540;
    13: op1_14_in08 = imem02_in[7:4];
    14: op1_14_in08 = reg_0984;
    15: op1_14_in08 = reg_0950;
    16: op1_14_in08 = reg_0682;
    17: op1_14_in08 = reg_0645;
    18: op1_14_in08 = reg_0455;
    19: op1_14_in08 = reg_0642;
    20: op1_14_in08 = reg_0686;
    21: op1_14_in08 = reg_0393;
    22: op1_14_in08 = reg_0757;
    23: op1_14_in08 = reg_0210;
    24: op1_14_in08 = imem07_in[87:84];
    25: op1_14_in08 = reg_0678;
    26: op1_14_in08 = reg_0068;
    27: op1_14_in08 = reg_0111;
    4: op1_14_in08 = reg_0163;
    3: op1_14_in08 = reg_0163;
    28: op1_14_in08 = reg_0659;
    29: op1_14_in08 = reg_0615;
    30: op1_14_in08 = reg_0480;
    31: op1_14_in08 = reg_0986;
    32: op1_14_in08 = imem05_in[19:16];
    33: op1_14_in08 = reg_0489;
    34: op1_14_in08 = reg_0884;
    35: op1_14_in08 = reg_0874;
    36: op1_14_in08 = reg_0311;
    37: op1_14_in08 = reg_0787;
    96: op1_14_in08 = reg_0787;
    38: op1_14_in08 = imem05_in[87:84];
    41: op1_14_in08 = reg_0668;
    42: op1_14_in08 = reg_0932;
    43: op1_14_in08 = reg_0754;
    44: op1_14_in08 = reg_0421;
    45: op1_14_in08 = reg_0116;
    46: op1_14_in08 = imem05_in[63:60];
    47: op1_14_in08 = reg_0705;
    48: op1_14_in08 = reg_0647;
    49: op1_14_in08 = reg_0397;
    50: op1_14_in08 = reg_0117;
    51: op1_14_in08 = reg_0677;
    52: op1_14_in08 = reg_1029;
    95: op1_14_in08 = reg_1029;
    53: op1_14_in08 = reg_0463;
    54: op1_14_in08 = reg_0694;
    55: op1_14_in08 = imem02_in[107:104];
    56: op1_14_in08 = reg_0434;
    57: op1_14_in08 = reg_0662;
    58: op1_14_in08 = reg_0651;
    59: op1_14_in08 = reg_0023;
    60: op1_14_in08 = reg_0240;
    61: op1_14_in08 = imem05_in[99:96];
    63: op1_14_in08 = reg_0314;
    64: op1_14_in08 = reg_0610;
    65: op1_14_in08 = reg_0759;
    66: op1_14_in08 = reg_0298;
    67: op1_14_in08 = reg_0424;
    68: op1_14_in08 = imem07_in[47:44];
    69: op1_14_in08 = reg_0900;
    70: op1_14_in08 = reg_0998;
    71: op1_14_in08 = imem06_in[43:40];
    72: op1_14_in08 = reg_0365;
    73: op1_14_in08 = reg_0672;
    74: op1_14_in08 = imem04_in[103:100];
    75: op1_14_in08 = imem05_in[95:92];
    76: op1_14_in08 = reg_0439;
    77: op1_14_in08 = imem00_in[99:96];
    78: op1_14_in08 = reg_0650;
    79: op1_14_in08 = imem02_in[103:100];
    80: op1_14_in08 = reg_0581;
    81: op1_14_in08 = imem05_in[55:52];
    82: op1_14_in08 = imem02_in[115:112];
    83: op1_14_in08 = reg_0883;
    85: op1_14_in08 = imem04_in[79:76];
    86: op1_14_in08 = reg_0278;
    87: op1_14_in08 = reg_0451;
    88: op1_14_in08 = reg_0376;
    89: op1_14_in08 = reg_0481;
    90: op1_14_in08 = reg_0358;
    91: op1_14_in08 = reg_0554;
    92: op1_14_in08 = imem06_in[83:80];
    94: op1_14_in08 = reg_0184;
    default: op1_14_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv08 = 1;
    6: op1_14_inv08 = 1;
    10: op1_14_inv08 = 1;
    12: op1_14_inv08 = 1;
    13: op1_14_inv08 = 1;
    14: op1_14_inv08 = 1;
    17: op1_14_inv08 = 1;
    19: op1_14_inv08 = 1;
    20: op1_14_inv08 = 1;
    22: op1_14_inv08 = 1;
    23: op1_14_inv08 = 1;
    24: op1_14_inv08 = 1;
    26: op1_14_inv08 = 1;
    28: op1_14_inv08 = 1;
    32: op1_14_inv08 = 1;
    33: op1_14_inv08 = 1;
    34: op1_14_inv08 = 1;
    36: op1_14_inv08 = 1;
    37: op1_14_inv08 = 1;
    41: op1_14_inv08 = 1;
    44: op1_14_inv08 = 1;
    46: op1_14_inv08 = 1;
    49: op1_14_inv08 = 1;
    50: op1_14_inv08 = 1;
    52: op1_14_inv08 = 1;
    54: op1_14_inv08 = 1;
    56: op1_14_inv08 = 1;
    61: op1_14_inv08 = 1;
    63: op1_14_inv08 = 1;
    65: op1_14_inv08 = 1;
    67: op1_14_inv08 = 1;
    72: op1_14_inv08 = 1;
    74: op1_14_inv08 = 1;
    76: op1_14_inv08 = 1;
    77: op1_14_inv08 = 1;
    80: op1_14_inv08 = 1;
    81: op1_14_inv08 = 1;
    82: op1_14_inv08 = 1;
    85: op1_14_inv08 = 1;
    89: op1_14_inv08 = 1;
    94: op1_14_inv08 = 1;
    95: op1_14_inv08 = 1;
    default: op1_14_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in09 = reg_0468;
    53: op1_14_in09 = reg_0468;
    6: op1_14_in09 = reg_0614;
    7: op1_14_in09 = reg_0658;
    8: op1_14_in09 = reg_0373;
    9: op1_14_in09 = reg_0685;
    10: op1_14_in09 = reg_0609;
    11: op1_14_in09 = reg_0338;
    12: op1_14_in09 = reg_0532;
    13: op1_14_in09 = imem02_in[31:28];
    14: op1_14_in09 = reg_1001;
    70: op1_14_in09 = reg_1001;
    15: op1_14_in09 = reg_0964;
    16: op1_14_in09 = reg_0690;
    17: op1_14_in09 = reg_0655;
    18: op1_14_in09 = reg_0469;
    19: op1_14_in09 = reg_0661;
    56: op1_14_in09 = reg_0661;
    60: op1_14_in09 = reg_0661;
    20: op1_14_in09 = reg_0677;
    21: op1_14_in09 = reg_0998;
    22: op1_14_in09 = reg_0260;
    23: op1_14_in09 = reg_0202;
    24: op1_14_in09 = imem07_in[119:116];
    25: op1_14_in09 = reg_0692;
    26: op1_14_in09 = reg_0071;
    27: op1_14_in09 = reg_0119;
    45: op1_14_in09 = reg_0119;
    4: op1_14_in09 = reg_0183;
    28: op1_14_in09 = reg_0339;
    29: op1_14_in09 = imem06_in[7:4];
    30: op1_14_in09 = reg_0471;
    31: op1_14_in09 = reg_0994;
    32: op1_14_in09 = imem05_in[39:36];
    33: op1_14_in09 = reg_0145;
    34: op1_14_in09 = imem03_in[7:4];
    35: op1_14_in09 = reg_0793;
    66: op1_14_in09 = reg_0793;
    36: op1_14_in09 = reg_0374;
    37: op1_14_in09 = reg_0073;
    38: op1_14_in09 = imem05_in[115:112];
    41: op1_14_in09 = reg_0680;
    42: op1_14_in09 = imem04_in[19:16];
    43: op1_14_in09 = reg_0293;
    44: op1_14_in09 = reg_0321;
    46: op1_14_in09 = imem05_in[71:68];
    47: op1_14_in09 = reg_0706;
    48: op1_14_in09 = reg_0082;
    49: op1_14_in09 = reg_0581;
    73: op1_14_in09 = reg_0581;
    50: op1_14_in09 = reg_0126;
    51: op1_14_in09 = reg_0673;
    52: op1_14_in09 = reg_0594;
    54: op1_14_in09 = reg_0698;
    76: op1_14_in09 = reg_0698;
    55: op1_14_in09 = reg_0642;
    57: op1_14_in09 = reg_0795;
    58: op1_14_in09 = reg_0647;
    59: op1_14_in09 = reg_0435;
    61: op1_14_in09 = reg_0233;
    63: op1_14_in09 = reg_0026;
    64: op1_14_in09 = reg_1053;
    65: op1_14_in09 = reg_0899;
    67: op1_14_in09 = reg_0329;
    68: op1_14_in09 = imem07_in[67:64];
    69: op1_14_in09 = reg_0670;
    71: op1_14_in09 = imem06_in[87:84];
    72: op1_14_in09 = reg_0094;
    74: op1_14_in09 = reg_0530;
    75: op1_14_in09 = imem05_in[103:100];
    77: op1_14_in09 = imem00_in[119:116];
    78: op1_14_in09 = reg_0810;
    79: op1_14_in09 = reg_0885;
    80: op1_14_in09 = reg_0985;
    81: op1_14_in09 = imem05_in[59:56];
    82: op1_14_in09 = imem02_in[127:124];
    83: op1_14_in09 = reg_0674;
    85: op1_14_in09 = imem04_in[91:88];
    86: op1_14_in09 = reg_0596;
    87: op1_14_in09 = reg_0477;
    88: op1_14_in09 = reg_0385;
    89: op1_14_in09 = reg_0472;
    90: op1_14_in09 = reg_0368;
    91: op1_14_in09 = reg_0372;
    92: op1_14_in09 = reg_0691;
    95: op1_14_in09 = reg_0169;
    96: op1_14_in09 = reg_0630;
    default: op1_14_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv09 = 1;
    6: op1_14_inv09 = 1;
    7: op1_14_inv09 = 1;
    8: op1_14_inv09 = 1;
    10: op1_14_inv09 = 1;
    11: op1_14_inv09 = 1;
    17: op1_14_inv09 = 1;
    19: op1_14_inv09 = 1;
    20: op1_14_inv09 = 1;
    22: op1_14_inv09 = 1;
    23: op1_14_inv09 = 1;
    24: op1_14_inv09 = 1;
    25: op1_14_inv09 = 1;
    27: op1_14_inv09 = 1;
    28: op1_14_inv09 = 1;
    30: op1_14_inv09 = 1;
    31: op1_14_inv09 = 1;
    33: op1_14_inv09 = 1;
    35: op1_14_inv09 = 1;
    37: op1_14_inv09 = 1;
    41: op1_14_inv09 = 1;
    42: op1_14_inv09 = 1;
    43: op1_14_inv09 = 1;
    45: op1_14_inv09 = 1;
    48: op1_14_inv09 = 1;
    51: op1_14_inv09 = 1;
    53: op1_14_inv09 = 1;
    64: op1_14_inv09 = 1;
    65: op1_14_inv09 = 1;
    66: op1_14_inv09 = 1;
    67: op1_14_inv09 = 1;
    68: op1_14_inv09 = 1;
    69: op1_14_inv09 = 1;
    71: op1_14_inv09 = 1;
    76: op1_14_inv09 = 1;
    77: op1_14_inv09 = 1;
    79: op1_14_inv09 = 1;
    80: op1_14_inv09 = 1;
    83: op1_14_inv09 = 1;
    85: op1_14_inv09 = 1;
    86: op1_14_inv09 = 1;
    90: op1_14_inv09 = 1;
    91: op1_14_inv09 = 1;
    92: op1_14_inv09 = 1;
    95: op1_14_inv09 = 1;
    default: op1_14_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in10 = reg_0192;
    6: op1_14_in10 = reg_0625;
    7: op1_14_in10 = reg_0664;
    8: op1_14_in10 = reg_0322;
    9: op1_14_in10 = reg_0672;
    10: op1_14_in10 = reg_0611;
    11: op1_14_in10 = reg_0350;
    12: op1_14_in10 = reg_0558;
    13: op1_14_in10 = imem02_in[51:48];
    14: op1_14_in10 = reg_0978;
    15: op1_14_in10 = reg_0946;
    16: op1_14_in10 = reg_0671;
    17: op1_14_in10 = reg_0661;
    18: op1_14_in10 = reg_0472;
    19: op1_14_in10 = reg_0647;
    20: op1_14_in10 = reg_0678;
    21: op1_14_in10 = reg_0982;
    22: op1_14_in10 = reg_0825;
    23: op1_14_in10 = reg_0197;
    24: op1_14_in10 = imem07_in[127:124];
    25: op1_14_in10 = reg_0465;
    26: op1_14_in10 = reg_0296;
    27: op1_14_in10 = reg_0115;
    4: op1_14_in10 = reg_0185;
    28: op1_14_in10 = reg_0776;
    29: op1_14_in10 = imem06_in[19:16];
    30: op1_14_in10 = reg_0479;
    31: op1_14_in10 = imem04_in[11:8];
    32: op1_14_in10 = imem05_in[63:60];
    33: op1_14_in10 = imem06_in[11:8];
    34: op1_14_in10 = imem03_in[59:56];
    35: op1_14_in10 = reg_0543;
    36: op1_14_in10 = reg_0234;
    37: op1_14_in10 = reg_0533;
    38: op1_14_in10 = reg_0959;
    41: op1_14_in10 = reg_0455;
    42: op1_14_in10 = imem04_in[43:40];
    43: op1_14_in10 = reg_0387;
    44: op1_14_in10 = reg_0744;
    45: op1_14_in10 = reg_0100;
    46: op1_14_in10 = imem05_in[79:76];
    81: op1_14_in10 = imem05_in[79:76];
    47: op1_14_in10 = reg_0250;
    48: op1_14_in10 = reg_0637;
    49: op1_14_in10 = reg_0396;
    50: op1_14_in10 = reg_0110;
    51: op1_14_in10 = reg_0699;
    54: op1_14_in10 = reg_0699;
    52: op1_14_in10 = reg_0630;
    53: op1_14_in10 = reg_0209;
    55: op1_14_in10 = reg_0515;
    56: op1_14_in10 = reg_0847;
    57: op1_14_in10 = reg_0246;
    58: op1_14_in10 = reg_0026;
    59: op1_14_in10 = reg_0336;
    60: op1_14_in10 = reg_0590;
    61: op1_14_in10 = reg_0757;
    63: op1_14_in10 = reg_0857;
    64: op1_14_in10 = reg_0114;
    65: op1_14_in10 = reg_0873;
    66: op1_14_in10 = reg_0513;
    67: op1_14_in10 = reg_0644;
    68: op1_14_in10 = imem07_in[71:68];
    69: op1_14_in10 = reg_0470;
    70: op1_14_in10 = reg_0975;
    71: op1_14_in10 = imem06_in[111:108];
    72: op1_14_in10 = reg_0360;
    73: op1_14_in10 = reg_0588;
    74: op1_14_in10 = reg_1020;
    75: op1_14_in10 = imem05_in[107:104];
    76: op1_14_in10 = reg_0915;
    77: op1_14_in10 = imem00_in[127:124];
    78: op1_14_in10 = reg_0700;
    79: op1_14_in10 = reg_0082;
    80: op1_14_in10 = reg_0992;
    82: op1_14_in10 = reg_0916;
    83: op1_14_in10 = reg_0463;
    85: op1_14_in10 = imem04_in[103:100];
    86: op1_14_in10 = reg_0239;
    87: op1_14_in10 = reg_0469;
    88: op1_14_in10 = reg_0551;
    89: op1_14_in10 = reg_0474;
    90: op1_14_in10 = reg_0155;
    91: op1_14_in10 = reg_0037;
    92: op1_14_in10 = reg_0439;
    95: op1_14_in10 = reg_0392;
    96: op1_14_in10 = reg_0510;
    default: op1_14_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv10 = 1;
    6: op1_14_inv10 = 1;
    7: op1_14_inv10 = 1;
    9: op1_14_inv10 = 1;
    12: op1_14_inv10 = 1;
    14: op1_14_inv10 = 1;
    15: op1_14_inv10 = 1;
    19: op1_14_inv10 = 1;
    20: op1_14_inv10 = 1;
    21: op1_14_inv10 = 1;
    24: op1_14_inv10 = 1;
    25: op1_14_inv10 = 1;
    26: op1_14_inv10 = 1;
    4: op1_14_inv10 = 1;
    28: op1_14_inv10 = 1;
    31: op1_14_inv10 = 1;
    33: op1_14_inv10 = 1;
    34: op1_14_inv10 = 1;
    35: op1_14_inv10 = 1;
    41: op1_14_inv10 = 1;
    42: op1_14_inv10 = 1;
    43: op1_14_inv10 = 1;
    44: op1_14_inv10 = 1;
    45: op1_14_inv10 = 1;
    47: op1_14_inv10 = 1;
    48: op1_14_inv10 = 1;
    49: op1_14_inv10 = 1;
    51: op1_14_inv10 = 1;
    53: op1_14_inv10 = 1;
    55: op1_14_inv10 = 1;
    57: op1_14_inv10 = 1;
    59: op1_14_inv10 = 1;
    60: op1_14_inv10 = 1;
    61: op1_14_inv10 = 1;
    63: op1_14_inv10 = 1;
    66: op1_14_inv10 = 1;
    69: op1_14_inv10 = 1;
    72: op1_14_inv10 = 1;
    73: op1_14_inv10 = 1;
    76: op1_14_inv10 = 1;
    77: op1_14_inv10 = 1;
    78: op1_14_inv10 = 1;
    79: op1_14_inv10 = 1;
    80: op1_14_inv10 = 1;
    82: op1_14_inv10 = 1;
    86: op1_14_inv10 = 1;
    87: op1_14_inv10 = 1;
    88: op1_14_inv10 = 1;
    91: op1_14_inv10 = 1;
    default: op1_14_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in11 = imem01_in[43:40];
    6: op1_14_in11 = reg_0605;
    7: op1_14_in11 = reg_0661;
    8: op1_14_in11 = reg_0361;
    9: op1_14_in11 = reg_0676;
    10: op1_14_in11 = reg_0618;
    11: op1_14_in11 = reg_0042;
    12: op1_14_in11 = reg_0533;
    96: op1_14_in11 = reg_0533;
    13: op1_14_in11 = imem02_in[79:76];
    14: op1_14_in11 = reg_0989;
    15: op1_14_in11 = reg_0952;
    16: op1_14_in11 = reg_0680;
    17: op1_14_in11 = reg_0639;
    18: op1_14_in11 = reg_0471;
    19: op1_14_in11 = reg_0649;
    20: op1_14_in11 = reg_0688;
    21: op1_14_in11 = reg_0984;
    22: op1_14_in11 = reg_0896;
    23: op1_14_in11 = imem01_in[63:60];
    24: op1_14_in11 = reg_0716;
    25: op1_14_in11 = reg_0454;
    26: op1_14_in11 = reg_0070;
    27: op1_14_in11 = reg_0121;
    4: op1_14_in11 = reg_0157;
    28: op1_14_in11 = reg_0761;
    29: op1_14_in11 = imem06_in[43:40];
    30: op1_14_in11 = reg_0459;
    31: op1_14_in11 = imem04_in[19:16];
    32: op1_14_in11 = imem05_in[75:72];
    33: op1_14_in11 = imem06_in[47:44];
    34: op1_14_in11 = imem03_in[83:80];
    35: op1_14_in11 = reg_0370;
    36: op1_14_in11 = reg_0991;
    88: op1_14_in11 = reg_0991;
    37: op1_14_in11 = reg_0403;
    38: op1_14_in11 = reg_0968;
    41: op1_14_in11 = reg_0461;
    42: op1_14_in11 = imem04_in[55:52];
    43: op1_14_in11 = reg_0294;
    44: op1_14_in11 = reg_0599;
    45: op1_14_in11 = reg_0101;
    64: op1_14_in11 = reg_0101;
    46: op1_14_in11 = imem05_in[95:92];
    47: op1_14_in11 = reg_0422;
    48: op1_14_in11 = reg_0621;
    49: op1_14_in11 = reg_0824;
    50: op1_14_in11 = imem02_in[7:4];
    51: op1_14_in11 = reg_0464;
    52: op1_14_in11 = reg_0596;
    53: op1_14_in11 = reg_0204;
    54: op1_14_in11 = reg_0451;
    55: op1_14_in11 = reg_0647;
    56: op1_14_in11 = reg_0038;
    57: op1_14_in11 = reg_0822;
    58: op1_14_in11 = reg_0279;
    59: op1_14_in11 = reg_0404;
    60: op1_14_in11 = reg_0784;
    61: op1_14_in11 = reg_0252;
    63: op1_14_in11 = reg_0673;
    65: op1_14_in11 = reg_0565;
    66: op1_14_in11 = reg_0987;
    67: op1_14_in11 = reg_0037;
    68: op1_14_in11 = imem07_in[87:84];
    69: op1_14_in11 = reg_0474;
    70: op1_14_in11 = reg_0994;
    71: op1_14_in11 = imem07_in[39:36];
    72: op1_14_in11 = imem02_in[27:24];
    73: op1_14_in11 = reg_0266;
    74: op1_14_in11 = reg_0778;
    75: op1_14_in11 = imem05_in[115:112];
    76: op1_14_in11 = reg_0782;
    77: op1_14_in11 = reg_0670;
    78: op1_14_in11 = reg_0885;
    79: op1_14_in11 = reg_0887;
    80: op1_14_in11 = reg_0981;
    81: op1_14_in11 = imem05_in[91:88];
    82: op1_14_in11 = reg_0637;
    83: op1_14_in11 = reg_0450;
    85: op1_14_in11 = imem04_in[107:104];
    86: op1_14_in11 = reg_0767;
    87: op1_14_in11 = reg_0473;
    89: op1_14_in11 = reg_0479;
    90: op1_14_in11 = reg_0082;
    91: op1_14_in11 = reg_0335;
    92: op1_14_in11 = reg_0606;
    95: op1_14_in11 = reg_0040;
    default: op1_14_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_14_inv11 = 1;
    8: op1_14_inv11 = 1;
    11: op1_14_inv11 = 1;
    12: op1_14_inv11 = 1;
    13: op1_14_inv11 = 1;
    14: op1_14_inv11 = 1;
    17: op1_14_inv11 = 1;
    18: op1_14_inv11 = 1;
    19: op1_14_inv11 = 1;
    25: op1_14_inv11 = 1;
    26: op1_14_inv11 = 1;
    27: op1_14_inv11 = 1;
    30: op1_14_inv11 = 1;
    31: op1_14_inv11 = 1;
    32: op1_14_inv11 = 1;
    35: op1_14_inv11 = 1;
    37: op1_14_inv11 = 1;
    41: op1_14_inv11 = 1;
    42: op1_14_inv11 = 1;
    43: op1_14_inv11 = 1;
    44: op1_14_inv11 = 1;
    45: op1_14_inv11 = 1;
    46: op1_14_inv11 = 1;
    48: op1_14_inv11 = 1;
    50: op1_14_inv11 = 1;
    51: op1_14_inv11 = 1;
    52: op1_14_inv11 = 1;
    55: op1_14_inv11 = 1;
    57: op1_14_inv11 = 1;
    60: op1_14_inv11 = 1;
    61: op1_14_inv11 = 1;
    64: op1_14_inv11 = 1;
    66: op1_14_inv11 = 1;
    67: op1_14_inv11 = 1;
    71: op1_14_inv11 = 1;
    72: op1_14_inv11 = 1;
    73: op1_14_inv11 = 1;
    77: op1_14_inv11 = 1;
    79: op1_14_inv11 = 1;
    80: op1_14_inv11 = 1;
    81: op1_14_inv11 = 1;
    82: op1_14_inv11 = 1;
    85: op1_14_inv11 = 1;
    86: op1_14_inv11 = 1;
    87: op1_14_inv11 = 1;
    88: op1_14_inv11 = 1;
    90: op1_14_inv11 = 1;
    91: op1_14_inv11 = 1;
    default: op1_14_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in12 = imem01_in[59:56];
    6: op1_14_in12 = reg_0626;
    52: op1_14_in12 = reg_0626;
    7: op1_14_in12 = reg_0656;
    8: op1_14_in12 = reg_0992;
    9: op1_14_in12 = reg_0698;
    10: op1_14_in12 = reg_0356;
    11: op1_14_in12 = reg_0055;
    12: op1_14_in12 = reg_0556;
    13: op1_14_in12 = reg_0646;
    14: op1_14_in12 = reg_0981;
    15: op1_14_in12 = reg_0972;
    16: op1_14_in12 = reg_0699;
    17: op1_14_in12 = reg_0651;
    18: op1_14_in12 = reg_0452;
    19: op1_14_in12 = reg_0352;
    20: op1_14_in12 = reg_0669;
    21: op1_14_in12 = reg_0999;
    22: op1_14_in12 = reg_0489;
    23: op1_14_in12 = imem01_in[71:68];
    24: op1_14_in12 = reg_0719;
    92: op1_14_in12 = reg_0719;
    25: op1_14_in12 = reg_0451;
    26: op1_14_in12 = reg_0059;
    27: op1_14_in12 = reg_0126;
    4: op1_14_in12 = reg_0173;
    28: op1_14_in12 = reg_0085;
    29: op1_14_in12 = imem06_in[47:44];
    30: op1_14_in12 = reg_0191;
    31: op1_14_in12 = imem04_in[23:20];
    32: op1_14_in12 = imem05_in[103:100];
    33: op1_14_in12 = imem06_in[55:52];
    34: op1_14_in12 = imem03_in[87:84];
    35: op1_14_in12 = reg_0836;
    36: op1_14_in12 = reg_0980;
    37: op1_14_in12 = reg_0566;
    38: op1_14_in12 = reg_1021;
    41: op1_14_in12 = reg_0476;
    54: op1_14_in12 = reg_0476;
    42: op1_14_in12 = imem04_in[59:56];
    80: op1_14_in12 = imem04_in[59:56];
    43: op1_14_in12 = reg_0264;
    44: op1_14_in12 = reg_0589;
    45: op1_14_in12 = reg_0109;
    46: op1_14_in12 = imem05_in[127:124];
    47: op1_14_in12 = reg_0047;
    48: op1_14_in12 = reg_0643;
    49: op1_14_in12 = reg_0389;
    50: op1_14_in12 = imem02_in[27:24];
    51: op1_14_in12 = reg_0466;
    53: op1_14_in12 = reg_0188;
    55: op1_14_in12 = reg_0652;
    56: op1_14_in12 = reg_0377;
    57: op1_14_in12 = reg_0987;
    73: op1_14_in12 = reg_0987;
    58: op1_14_in12 = reg_0323;
    59: op1_14_in12 = reg_0135;
    60: op1_14_in12 = reg_0518;
    61: op1_14_in12 = reg_0023;
    63: op1_14_in12 = reg_0281;
    64: op1_14_in12 = imem02_in[23:20];
    65: op1_14_in12 = reg_0645;
    66: op1_14_in12 = reg_1001;
    67: op1_14_in12 = reg_0054;
    68: op1_14_in12 = imem07_in[107:104];
    69: op1_14_in12 = reg_0456;
    70: op1_14_in12 = imem04_in[7:4];
    71: op1_14_in12 = imem07_in[55:52];
    72: op1_14_in12 = imem02_in[47:44];
    74: op1_14_in12 = reg_0909;
    75: op1_14_in12 = reg_0136;
    76: op1_14_in12 = reg_0022;
    77: op1_14_in12 = reg_0687;
    78: op1_14_in12 = reg_0034;
    79: op1_14_in12 = reg_0762;
    81: op1_14_in12 = imem05_in[99:96];
    82: op1_14_in12 = reg_0833;
    83: op1_14_in12 = reg_0481;
    85: op1_14_in12 = imem04_in[115:112];
    86: op1_14_in12 = reg_0597;
    87: op1_14_in12 = reg_0459;
    89: op1_14_in12 = reg_0459;
    88: op1_14_in12 = reg_0995;
    90: op1_14_in12 = reg_0713;
    91: op1_14_in12 = reg_0045;
    95: op1_14_in12 = reg_0628;
    96: op1_14_in12 = reg_0289;
    default: op1_14_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv12 = 1;
    7: op1_14_inv12 = 1;
    9: op1_14_inv12 = 1;
    10: op1_14_inv12 = 1;
    11: op1_14_inv12 = 1;
    12: op1_14_inv12 = 1;
    13: op1_14_inv12 = 1;
    16: op1_14_inv12 = 1;
    17: op1_14_inv12 = 1;
    18: op1_14_inv12 = 1;
    20: op1_14_inv12 = 1;
    22: op1_14_inv12 = 1;
    27: op1_14_inv12 = 1;
    4: op1_14_inv12 = 1;
    28: op1_14_inv12 = 1;
    29: op1_14_inv12 = 1;
    33: op1_14_inv12 = 1;
    34: op1_14_inv12 = 1;
    36: op1_14_inv12 = 1;
    38: op1_14_inv12 = 1;
    41: op1_14_inv12 = 1;
    44: op1_14_inv12 = 1;
    45: op1_14_inv12 = 1;
    47: op1_14_inv12 = 1;
    48: op1_14_inv12 = 1;
    52: op1_14_inv12 = 1;
    55: op1_14_inv12 = 1;
    56: op1_14_inv12 = 1;
    58: op1_14_inv12 = 1;
    59: op1_14_inv12 = 1;
    65: op1_14_inv12 = 1;
    66: op1_14_inv12 = 1;
    67: op1_14_inv12 = 1;
    68: op1_14_inv12 = 1;
    70: op1_14_inv12 = 1;
    79: op1_14_inv12 = 1;
    86: op1_14_inv12 = 1;
    88: op1_14_inv12 = 1;
    91: op1_14_inv12 = 1;
    95: op1_14_inv12 = 1;
    default: op1_14_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in13 = imem01_in[67:64];
    6: op1_14_in13 = reg_0618;
    7: op1_14_in13 = reg_0651;
    8: op1_14_in13 = reg_0995;
    9: op1_14_in13 = reg_0679;
    10: op1_14_in13 = reg_0381;
    11: op1_14_in13 = imem03_in[23:20];
    12: op1_14_in13 = reg_0299;
    13: op1_14_in13 = reg_0363;
    14: op1_14_in13 = reg_0975;
    15: op1_14_in13 = reg_0900;
    16: op1_14_in13 = reg_0451;
    17: op1_14_in13 = reg_0640;
    18: op1_14_in13 = reg_0196;
    19: op1_14_in13 = reg_0357;
    20: op1_14_in13 = reg_0464;
    21: op1_14_in13 = reg_0988;
    22: op1_14_in13 = reg_0132;
    23: op1_14_in13 = reg_1053;
    24: op1_14_in13 = reg_0721;
    25: op1_14_in13 = reg_0475;
    26: op1_14_in13 = reg_0738;
    27: op1_14_in13 = reg_0110;
    28: op1_14_in13 = reg_0484;
    29: op1_14_in13 = imem06_in[55:52];
    30: op1_14_in13 = reg_0211;
    31: op1_14_in13 = imem04_in[103:100];
    32: op1_14_in13 = imem05_in[119:116];
    33: op1_14_in13 = imem06_in[95:92];
    34: op1_14_in13 = imem03_in[91:88];
    35: op1_14_in13 = reg_0513;
    60: op1_14_in13 = reg_0513;
    36: op1_14_in13 = imem04_in[3:0];
    37: op1_14_in13 = reg_0588;
    38: op1_14_in13 = reg_0491;
    41: op1_14_in13 = reg_0479;
    42: op1_14_in13 = imem04_in[63:60];
    43: op1_14_in13 = reg_0594;
    44: op1_14_in13 = reg_0868;
    45: op1_14_in13 = reg_0035;
    46: op1_14_in13 = reg_0970;
    47: op1_14_in13 = reg_0321;
    48: op1_14_in13 = reg_0648;
    49: op1_14_in13 = reg_0874;
    50: op1_14_in13 = imem02_in[51:48];
    51: op1_14_in13 = reg_0470;
    52: op1_14_in13 = imem07_in[55:52];
    53: op1_14_in13 = reg_0307;
    54: op1_14_in13 = reg_0466;
    55: op1_14_in13 = reg_0359;
    56: op1_14_in13 = reg_0376;
    57: op1_14_in13 = reg_0996;
    58: op1_14_in13 = reg_0358;
    59: op1_14_in13 = reg_0154;
    61: op1_14_in13 = reg_0436;
    63: op1_14_in13 = reg_0667;
    64: op1_14_in13 = imem02_in[111:108];
    65: op1_14_in13 = reg_0516;
    66: op1_14_in13 = reg_0986;
    67: op1_14_in13 = reg_0776;
    68: op1_14_in13 = reg_0719;
    69: op1_14_in13 = reg_0189;
    70: op1_14_in13 = imem04_in[11:8];
    71: op1_14_in13 = imem07_in[79:76];
    72: op1_14_in13 = imem02_in[63:60];
    73: op1_14_in13 = reg_0992;
    74: op1_14_in13 = reg_0524;
    75: op1_14_in13 = reg_0142;
    76: op1_14_in13 = imem07_in[3:0];
    77: op1_14_in13 = reg_0465;
    78: op1_14_in13 = reg_0643;
    79: op1_14_in13 = reg_0389;
    80: op1_14_in13 = reg_1004;
    81: op1_14_in13 = imem05_in[127:124];
    82: op1_14_in13 = reg_0846;
    83: op1_14_in13 = reg_0456;
    85: op1_14_in13 = imem04_in[119:116];
    86: op1_14_in13 = reg_0998;
    87: op1_14_in13 = reg_0204;
    88: op1_14_in13 = reg_0993;
    89: op1_14_in13 = reg_0188;
    90: op1_14_in13 = reg_0573;
    91: op1_14_in13 = reg_0355;
    92: op1_14_in13 = reg_1020;
    95: op1_14_in13 = reg_0403;
    96: op1_14_in13 = reg_0040;
    default: op1_14_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv13 = 1;
    6: op1_14_inv13 = 1;
    7: op1_14_inv13 = 1;
    8: op1_14_inv13 = 1;
    9: op1_14_inv13 = 1;
    11: op1_14_inv13 = 1;
    14: op1_14_inv13 = 1;
    17: op1_14_inv13 = 1;
    26: op1_14_inv13 = 1;
    27: op1_14_inv13 = 1;
    29: op1_14_inv13 = 1;
    30: op1_14_inv13 = 1;
    31: op1_14_inv13 = 1;
    33: op1_14_inv13 = 1;
    34: op1_14_inv13 = 1;
    37: op1_14_inv13 = 1;
    42: op1_14_inv13 = 1;
    43: op1_14_inv13 = 1;
    44: op1_14_inv13 = 1;
    45: op1_14_inv13 = 1;
    48: op1_14_inv13 = 1;
    49: op1_14_inv13 = 1;
    51: op1_14_inv13 = 1;
    59: op1_14_inv13 = 1;
    60: op1_14_inv13 = 1;
    63: op1_14_inv13 = 1;
    64: op1_14_inv13 = 1;
    67: op1_14_inv13 = 1;
    69: op1_14_inv13 = 1;
    72: op1_14_inv13 = 1;
    73: op1_14_inv13 = 1;
    79: op1_14_inv13 = 1;
    80: op1_14_inv13 = 1;
    82: op1_14_inv13 = 1;
    89: op1_14_inv13 = 1;
    96: op1_14_inv13 = 1;
    default: op1_14_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in14 = imem01_in[75:72];
    6: op1_14_in14 = reg_0356;
    7: op1_14_in14 = reg_0636;
    8: op1_14_in14 = reg_0986;
    9: op1_14_in14 = reg_0677;
    10: op1_14_in14 = reg_0408;
    11: op1_14_in14 = imem03_in[59:56];
    12: op1_14_in14 = reg_0282;
    13: op1_14_in14 = reg_0328;
    14: op1_14_in14 = reg_1000;
    21: op1_14_in14 = reg_1000;
    15: op1_14_in14 = reg_0229;
    16: op1_14_in14 = reg_0464;
    77: op1_14_in14 = reg_0464;
    17: op1_14_in14 = reg_0663;
    18: op1_14_in14 = reg_0202;
    19: op1_14_in14 = reg_0320;
    20: op1_14_in14 = reg_0461;
    22: op1_14_in14 = reg_0148;
    23: op1_14_in14 = reg_0236;
    24: op1_14_in14 = reg_0717;
    25: op1_14_in14 = reg_0472;
    26: op1_14_in14 = reg_0773;
    27: op1_14_in14 = imem02_in[27:24];
    28: op1_14_in14 = reg_0077;
    29: op1_14_in14 = imem06_in[75:72];
    30: op1_14_in14 = reg_0201;
    31: op1_14_in14 = reg_0483;
    32: op1_14_in14 = reg_0963;
    33: op1_14_in14 = imem06_in[123:120];
    34: op1_14_in14 = imem03_in[95:92];
    35: op1_14_in14 = reg_0374;
    36: op1_14_in14 = imem04_in[95:92];
    37: op1_14_in14 = reg_0385;
    38: op1_14_in14 = reg_0275;
    41: op1_14_in14 = reg_0452;
    51: op1_14_in14 = reg_0452;
    42: op1_14_in14 = imem04_in[71:68];
    43: op1_14_in14 = reg_0309;
    44: op1_14_in14 = reg_0159;
    45: op1_14_in14 = reg_0517;
    46: op1_14_in14 = reg_0957;
    47: op1_14_in14 = reg_0599;
    48: op1_14_in14 = reg_0652;
    49: op1_14_in14 = reg_0376;
    50: op1_14_in14 = imem02_in[63:60];
    52: op1_14_in14 = imem07_in[67:64];
    53: op1_14_in14 = reg_0106;
    54: op1_14_in14 = reg_0481;
    55: op1_14_in14 = reg_0329;
    56: op1_14_in14 = reg_0312;
    57: op1_14_in14 = reg_0990;
    58: op1_14_in14 = reg_0039;
    59: op1_14_in14 = reg_0141;
    60: op1_14_in14 = reg_0996;
    61: op1_14_in14 = reg_0404;
    63: op1_14_in14 = imem02_in[3:0];
    64: op1_14_in14 = reg_0355;
    65: op1_14_in14 = reg_0772;
    79: op1_14_in14 = reg_0772;
    66: op1_14_in14 = reg_0976;
    67: op1_14_in14 = reg_0761;
    68: op1_14_in14 = reg_0710;
    69: op1_14_in14 = reg_0207;
    70: op1_14_in14 = imem04_in[35:32];
    71: op1_14_in14 = imem07_in[103:100];
    72: op1_14_in14 = imem02_in[75:72];
    73: op1_14_in14 = reg_0984;
    74: op1_14_in14 = reg_0284;
    75: op1_14_in14 = reg_0013;
    76: op1_14_in14 = imem07_in[11:8];
    78: op1_14_in14 = reg_0341;
    80: op1_14_in14 = reg_1003;
    81: op1_14_in14 = reg_0215;
    82: op1_14_in14 = reg_0885;
    83: op1_14_in14 = reg_0200;
    85: op1_14_in14 = reg_0577;
    86: op1_14_in14 = reg_0991;
    87: op1_14_in14 = reg_0194;
    88: op1_14_in14 = reg_0989;
    89: op1_14_in14 = reg_0211;
    90: op1_14_in14 = reg_0311;
    91: op1_14_in14 = reg_0155;
    92: op1_14_in14 = reg_0036;
    95: op1_14_in14 = reg_0782;
    96: op1_14_in14 = reg_0020;
    default: op1_14_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv14 = 1;
    6: op1_14_inv14 = 1;
    7: op1_14_inv14 = 1;
    9: op1_14_inv14 = 1;
    11: op1_14_inv14 = 1;
    13: op1_14_inv14 = 1;
    14: op1_14_inv14 = 1;
    15: op1_14_inv14 = 1;
    16: op1_14_inv14 = 1;
    17: op1_14_inv14 = 1;
    18: op1_14_inv14 = 1;
    23: op1_14_inv14 = 1;
    25: op1_14_inv14 = 1;
    26: op1_14_inv14 = 1;
    27: op1_14_inv14 = 1;
    31: op1_14_inv14 = 1;
    32: op1_14_inv14 = 1;
    33: op1_14_inv14 = 1;
    34: op1_14_inv14 = 1;
    36: op1_14_inv14 = 1;
    38: op1_14_inv14 = 1;
    41: op1_14_inv14 = 1;
    43: op1_14_inv14 = 1;
    45: op1_14_inv14 = 1;
    46: op1_14_inv14 = 1;
    49: op1_14_inv14 = 1;
    53: op1_14_inv14 = 1;
    54: op1_14_inv14 = 1;
    55: op1_14_inv14 = 1;
    56: op1_14_inv14 = 1;
    58: op1_14_inv14 = 1;
    64: op1_14_inv14 = 1;
    65: op1_14_inv14 = 1;
    66: op1_14_inv14 = 1;
    69: op1_14_inv14 = 1;
    70: op1_14_inv14 = 1;
    71: op1_14_inv14 = 1;
    74: op1_14_inv14 = 1;
    75: op1_14_inv14 = 1;
    78: op1_14_inv14 = 1;
    80: op1_14_inv14 = 1;
    81: op1_14_inv14 = 1;
    82: op1_14_inv14 = 1;
    86: op1_14_inv14 = 1;
    88: op1_14_inv14 = 1;
    90: op1_14_inv14 = 1;
    92: op1_14_inv14 = 1;
    95: op1_14_inv14 = 1;
    96: op1_14_inv14 = 1;
    default: op1_14_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in15 = imem01_in[83:80];
    6: op1_14_in15 = reg_0372;
    7: op1_14_in15 = reg_0333;
    8: op1_14_in15 = reg_0978;
    9: op1_14_in15 = reg_0691;
    10: op1_14_in15 = reg_0392;
    11: op1_14_in15 = imem03_in[87:84];
    12: op1_14_in15 = reg_0296;
    13: op1_14_in15 = reg_0086;
    67: op1_14_in15 = reg_0086;
    14: op1_14_in15 = imem04_in[47:44];
    15: op1_14_in15 = reg_0253;
    16: op1_14_in15 = reg_0474;
    17: op1_14_in15 = reg_0334;
    18: op1_14_in15 = reg_0197;
    19: op1_14_in15 = reg_0318;
    20: op1_14_in15 = reg_0472;
    21: op1_14_in15 = imem04_in[27:24];
    57: op1_14_in15 = imem04_in[27:24];
    22: op1_14_in15 = reg_0142;
    23: op1_14_in15 = reg_0238;
    24: op1_14_in15 = reg_0715;
    25: op1_14_in15 = reg_0471;
    26: op1_14_in15 = reg_0021;
    27: op1_14_in15 = imem02_in[47:44];
    28: op1_14_in15 = reg_0321;
    29: op1_14_in15 = imem06_in[79:76];
    30: op1_14_in15 = reg_0196;
    31: op1_14_in15 = reg_0265;
    32: op1_14_in15 = reg_0973;
    33: op1_14_in15 = reg_0610;
    34: op1_14_in15 = imem03_in[103:100];
    35: op1_14_in15 = reg_0234;
    36: op1_14_in15 = imem04_in[111:108];
    37: op1_14_in15 = reg_0293;
    38: op1_14_in15 = reg_0130;
    41: op1_14_in15 = reg_0458;
    42: op1_14_in15 = imem04_in[99:96];
    43: op1_14_in15 = reg_0633;
    44: op1_14_in15 = reg_0160;
    45: op1_14_in15 = reg_0036;
    96: op1_14_in15 = reg_0036;
    46: op1_14_in15 = reg_0022;
    47: op1_14_in15 = reg_0502;
    48: op1_14_in15 = reg_0916;
    49: op1_14_in15 = reg_0985;
    50: op1_14_in15 = imem02_in[67:64];
    51: op1_14_in15 = reg_0214;
    52: op1_14_in15 = imem07_in[87:84];
    53: op1_14_in15 = reg_0018;
    54: op1_14_in15 = reg_0459;
    55: op1_14_in15 = reg_0423;
    56: op1_14_in15 = reg_0822;
    58: op1_14_in15 = reg_0368;
    59: op1_14_in15 = reg_0140;
    60: op1_14_in15 = reg_1001;
    61: op1_14_in15 = reg_0447;
    63: op1_14_in15 = imem02_in[19:16];
    64: op1_14_in15 = reg_0666;
    65: op1_14_in15 = reg_0776;
    66: op1_14_in15 = imem04_in[3:0];
    68: op1_14_in15 = reg_0731;
    69: op1_14_in15 = reg_0124;
    70: op1_14_in15 = imem04_in[115:112];
    71: op1_14_in15 = imem07_in[127:124];
    72: op1_14_in15 = reg_0279;
    73: op1_14_in15 = reg_0989;
    74: op1_14_in15 = reg_0432;
    75: op1_14_in15 = reg_0259;
    76: op1_14_in15 = imem07_in[51:48];
    77: op1_14_in15 = reg_0481;
    78: op1_14_in15 = reg_0425;
    79: op1_14_in15 = reg_0761;
    80: op1_14_in15 = reg_0061;
    81: op1_14_in15 = reg_0319;
    82: op1_14_in15 = reg_0082;
    83: op1_14_in15 = reg_0208;
    85: op1_14_in15 = reg_0942;
    86: op1_14_in15 = reg_0979;
    87: op1_14_in15 = reg_0195;
    88: op1_14_in15 = reg_0988;
    89: op1_14_in15 = reg_0199;
    90: op1_14_in15 = reg_0984;
    91: op1_14_in15 = reg_0085;
    92: op1_14_in15 = imem07_in[7:4];
    95: op1_14_in15 = reg_0084;
    default: op1_14_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_14_inv15 = 1;
    8: op1_14_inv15 = 1;
    9: op1_14_inv15 = 1;
    10: op1_14_inv15 = 1;
    12: op1_14_inv15 = 1;
    14: op1_14_inv15 = 1;
    16: op1_14_inv15 = 1;
    18: op1_14_inv15 = 1;
    19: op1_14_inv15 = 1;
    20: op1_14_inv15 = 1;
    21: op1_14_inv15 = 1;
    22: op1_14_inv15 = 1;
    23: op1_14_inv15 = 1;
    24: op1_14_inv15 = 1;
    30: op1_14_inv15 = 1;
    32: op1_14_inv15 = 1;
    34: op1_14_inv15 = 1;
    35: op1_14_inv15 = 1;
    42: op1_14_inv15 = 1;
    44: op1_14_inv15 = 1;
    45: op1_14_inv15 = 1;
    48: op1_14_inv15 = 1;
    49: op1_14_inv15 = 1;
    53: op1_14_inv15 = 1;
    54: op1_14_inv15 = 1;
    61: op1_14_inv15 = 1;
    66: op1_14_inv15 = 1;
    67: op1_14_inv15 = 1;
    68: op1_14_inv15 = 1;
    69: op1_14_inv15 = 1;
    72: op1_14_inv15 = 1;
    73: op1_14_inv15 = 1;
    75: op1_14_inv15 = 1;
    78: op1_14_inv15 = 1;
    79: op1_14_inv15 = 1;
    82: op1_14_inv15 = 1;
    86: op1_14_inv15 = 1;
    87: op1_14_inv15 = 1;
    88: op1_14_inv15 = 1;
    89: op1_14_inv15 = 1;
    92: op1_14_inv15 = 1;
    95: op1_14_inv15 = 1;
    default: op1_14_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in16 = imem01_in[95:92];
    6: op1_14_in16 = reg_0313;
    7: op1_14_in16 = reg_0326;
    8: op1_14_in16 = reg_0997;
    9: op1_14_in16 = reg_0673;
    10: op1_14_in16 = reg_0409;
    11: op1_14_in16 = imem03_in[99:96];
    12: op1_14_in16 = reg_0286;
    13: op1_14_in16 = reg_0090;
    14: op1_14_in16 = imem04_in[63:60];
    15: op1_14_in16 = reg_0148;
    61: op1_14_in16 = reg_0148;
    16: op1_14_in16 = reg_0189;
    17: op1_14_in16 = reg_0320;
    18: op1_14_in16 = imem01_in[27:24];
    19: op1_14_in16 = reg_0310;
    20: op1_14_in16 = reg_0467;
    77: op1_14_in16 = reg_0467;
    21: op1_14_in16 = imem04_in[35:32];
    22: op1_14_in16 = reg_0139;
    23: op1_14_in16 = reg_1050;
    24: op1_14_in16 = reg_0701;
    25: op1_14_in16 = reg_0468;
    26: op1_14_in16 = imem05_in[83:80];
    27: op1_14_in16 = imem02_in[51:48];
    28: op1_14_in16 = reg_0323;
    29: op1_14_in16 = imem06_in[87:84];
    30: op1_14_in16 = reg_0212;
    31: op1_14_in16 = reg_0539;
    32: op1_14_in16 = reg_0944;
    33: op1_14_in16 = reg_0613;
    34: op1_14_in16 = imem03_in[115:112];
    35: op1_14_in16 = reg_0982;
    36: op1_14_in16 = reg_0483;
    37: op1_14_in16 = reg_0356;
    38: op1_14_in16 = imem06_in[3:0];
    41: op1_14_in16 = reg_0200;
    42: op1_14_in16 = imem04_in[103:100];
    43: op1_14_in16 = reg_0008;
    44: op1_14_in16 = reg_0183;
    45: op1_14_in16 = reg_0449;
    46: op1_14_in16 = reg_0252;
    47: op1_14_in16 = reg_0640;
    48: op1_14_in16 = reg_0081;
    49: op1_14_in16 = reg_1002;
    50: op1_14_in16 = imem02_in[99:96];
    51: op1_14_in16 = reg_0191;
    52: op1_14_in16 = reg_0720;
    53: op1_14_in16 = reg_0240;
    54: op1_14_in16 = reg_0478;
    55: op1_14_in16 = reg_0772;
    56: op1_14_in16 = reg_0991;
    57: op1_14_in16 = imem04_in[39:36];
    58: op1_14_in16 = reg_0335;
    59: op1_14_in16 = reg_0131;
    60: op1_14_in16 = imem04_in[7:4];
    63: op1_14_in16 = imem02_in[31:28];
    64: op1_14_in16 = reg_0224;
    65: op1_14_in16 = reg_0761;
    66: op1_14_in16 = imem04_in[11:8];
    67: op1_14_in16 = reg_0091;
    68: op1_14_in16 = reg_0708;
    71: op1_14_in16 = reg_0708;
    69: op1_14_in16 = reg_0247;
    70: op1_14_in16 = imem04_in[119:116];
    72: op1_14_in16 = reg_0441;
    73: op1_14_in16 = reg_0974;
    74: op1_14_in16 = reg_0552;
    75: op1_14_in16 = reg_0935;
    76: op1_14_in16 = imem07_in[59:56];
    78: op1_14_in16 = reg_0331;
    79: op1_14_in16 = reg_0085;
    80: op1_14_in16 = reg_0777;
    81: op1_14_in16 = reg_0143;
    82: op1_14_in16 = reg_0098;
    83: op1_14_in16 = reg_0186;
    85: op1_14_in16 = reg_0292;
    86: op1_14_in16 = reg_0984;
    87: op1_14_in16 = imem01_in[19:16];
    88: op1_14_in16 = imem04_in[23:20];
    89: op1_14_in16 = imem01_in[7:4];
    90: op1_14_in16 = reg_0228;
    91: op1_14_in16 = reg_0656;
    92: op1_14_in16 = imem07_in[19:16];
    95: op1_14_in16 = reg_0566;
    96: op1_14_in16 = reg_0403;
    default: op1_14_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv16 = 1;
    8: op1_14_inv16 = 1;
    9: op1_14_inv16 = 1;
    13: op1_14_inv16 = 1;
    14: op1_14_inv16 = 1;
    15: op1_14_inv16 = 1;
    16: op1_14_inv16 = 1;
    18: op1_14_inv16 = 1;
    22: op1_14_inv16 = 1;
    24: op1_14_inv16 = 1;
    27: op1_14_inv16 = 1;
    28: op1_14_inv16 = 1;
    29: op1_14_inv16 = 1;
    30: op1_14_inv16 = 1;
    32: op1_14_inv16 = 1;
    33: op1_14_inv16 = 1;
    35: op1_14_inv16 = 1;
    36: op1_14_inv16 = 1;
    37: op1_14_inv16 = 1;
    41: op1_14_inv16 = 1;
    43: op1_14_inv16 = 1;
    46: op1_14_inv16 = 1;
    47: op1_14_inv16 = 1;
    48: op1_14_inv16 = 1;
    51: op1_14_inv16 = 1;
    53: op1_14_inv16 = 1;
    56: op1_14_inv16 = 1;
    60: op1_14_inv16 = 1;
    61: op1_14_inv16 = 1;
    68: op1_14_inv16 = 1;
    69: op1_14_inv16 = 1;
    70: op1_14_inv16 = 1;
    72: op1_14_inv16 = 1;
    74: op1_14_inv16 = 1;
    77: op1_14_inv16 = 1;
    78: op1_14_inv16 = 1;
    79: op1_14_inv16 = 1;
    80: op1_14_inv16 = 1;
    81: op1_14_inv16 = 1;
    85: op1_14_inv16 = 1;
    86: op1_14_inv16 = 1;
    88: op1_14_inv16 = 1;
    89: op1_14_inv16 = 1;
    91: op1_14_inv16 = 1;
    92: op1_14_inv16 = 1;
    95: op1_14_inv16 = 1;
    96: op1_14_inv16 = 1;
    default: op1_14_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in17 = imem01_in[123:120];
    6: op1_14_in17 = reg_0404;
    7: op1_14_in17 = reg_0354;
    8: op1_14_in17 = imem04_in[119:116];
    9: op1_14_in17 = reg_0463;
    10: op1_14_in17 = reg_0315;
    11: op1_14_in17 = reg_0573;
    12: op1_14_in17 = reg_0019;
    13: op1_14_in17 = reg_0087;
    14: op1_14_in17 = imem04_in[111:108];
    42: op1_14_in17 = imem04_in[111:108];
    15: op1_14_in17 = reg_0149;
    16: op1_14_in17 = reg_0204;
    17: op1_14_in17 = reg_0330;
    18: op1_14_in17 = imem01_in[43:40];
    19: op1_14_in17 = reg_0328;
    20: op1_14_in17 = reg_0471;
    77: op1_14_in17 = reg_0471;
    21: op1_14_in17 = imem04_in[43:40];
    22: op1_14_in17 = reg_0129;
    23: op1_14_in17 = reg_0249;
    24: op1_14_in17 = reg_0700;
    25: op1_14_in17 = reg_0208;
    26: op1_14_in17 = imem05_in[91:88];
    27: op1_14_in17 = imem02_in[55:52];
    28: op1_14_in17 = reg_0744;
    29: op1_14_in17 = imem06_in[99:96];
    30: op1_14_in17 = imem01_in[3:0];
    31: op1_14_in17 = reg_0888;
    32: op1_14_in17 = reg_0956;
    33: op1_14_in17 = reg_0620;
    34: op1_14_in17 = imem03_in[127:124];
    35: op1_14_in17 = reg_0986;
    86: op1_14_in17 = reg_0986;
    36: op1_14_in17 = reg_0265;
    37: op1_14_in17 = reg_0386;
    38: op1_14_in17 = imem06_in[11:8];
    41: op1_14_in17 = reg_0188;
    43: op1_14_in17 = reg_0263;
    44: op1_14_in17 = reg_0166;
    45: op1_14_in17 = reg_0644;
    46: op1_14_in17 = reg_0491;
    47: op1_14_in17 = reg_0175;
    48: op1_14_in17 = reg_0080;
    49: op1_14_in17 = reg_0991;
    50: op1_14_in17 = reg_0653;
    51: op1_14_in17 = reg_0189;
    52: op1_14_in17 = reg_0710;
    53: op1_14_in17 = reg_0928;
    54: op1_14_in17 = reg_0458;
    55: op1_14_in17 = reg_0792;
    56: op1_14_in17 = imem04_in[51:48];
    57: op1_14_in17 = imem04_in[79:76];
    58: op1_14_in17 = reg_0772;
    59: op1_14_in17 = reg_0134;
    60: op1_14_in17 = imem04_in[19:16];
    66: op1_14_in17 = imem04_in[19:16];
    61: op1_14_in17 = reg_0135;
    63: op1_14_in17 = reg_0279;
    64: op1_14_in17 = reg_0648;
    65: op1_14_in17 = reg_0086;
    79: op1_14_in17 = reg_0086;
    67: op1_14_in17 = reg_0291;
    68: op1_14_in17 = reg_0715;
    69: op1_14_in17 = imem01_in[15:12];
    70: op1_14_in17 = reg_0530;
    71: op1_14_in17 = reg_0711;
    72: op1_14_in17 = reg_0052;
    82: op1_14_in17 = reg_0052;
    73: op1_14_in17 = reg_0977;
    74: op1_14_in17 = reg_0027;
    75: op1_14_in17 = reg_0447;
    76: op1_14_in17 = imem07_in[67:64];
    78: op1_14_in17 = reg_0089;
    80: op1_14_in17 = reg_0295;
    81: op1_14_in17 = reg_0139;
    83: op1_14_in17 = reg_0198;
    85: op1_14_in17 = reg_0031;
    87: op1_14_in17 = imem01_in[27:24];
    88: op1_14_in17 = imem04_in[59:56];
    89: op1_14_in17 = imem01_in[35:32];
    90: op1_14_in17 = reg_0585;
    91: op1_14_in17 = reg_0082;
    92: op1_14_in17 = imem07_in[35:32];
    95: op1_14_in17 = imem07_in[31:28];
    96: op1_14_in17 = reg_0804;
    default: op1_14_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_14_inv17 = 1;
    10: op1_14_inv17 = 1;
    12: op1_14_inv17 = 1;
    13: op1_14_inv17 = 1;
    15: op1_14_inv17 = 1;
    16: op1_14_inv17 = 1;
    17: op1_14_inv17 = 1;
    19: op1_14_inv17 = 1;
    21: op1_14_inv17 = 1;
    23: op1_14_inv17 = 1;
    24: op1_14_inv17 = 1;
    25: op1_14_inv17 = 1;
    26: op1_14_inv17 = 1;
    28: op1_14_inv17 = 1;
    30: op1_14_inv17 = 1;
    32: op1_14_inv17 = 1;
    33: op1_14_inv17 = 1;
    36: op1_14_inv17 = 1;
    37: op1_14_inv17 = 1;
    38: op1_14_inv17 = 1;
    41: op1_14_inv17 = 1;
    42: op1_14_inv17 = 1;
    44: op1_14_inv17 = 1;
    46: op1_14_inv17 = 1;
    48: op1_14_inv17 = 1;
    50: op1_14_inv17 = 1;
    53: op1_14_inv17 = 1;
    56: op1_14_inv17 = 1;
    58: op1_14_inv17 = 1;
    59: op1_14_inv17 = 1;
    60: op1_14_inv17 = 1;
    61: op1_14_inv17 = 1;
    63: op1_14_inv17 = 1;
    66: op1_14_inv17 = 1;
    68: op1_14_inv17 = 1;
    69: op1_14_inv17 = 1;
    70: op1_14_inv17 = 1;
    71: op1_14_inv17 = 1;
    74: op1_14_inv17 = 1;
    78: op1_14_inv17 = 1;
    79: op1_14_inv17 = 1;
    81: op1_14_inv17 = 1;
    82: op1_14_inv17 = 1;
    87: op1_14_inv17 = 1;
    88: op1_14_inv17 = 1;
    90: op1_14_inv17 = 1;
    91: op1_14_inv17 = 1;
    92: op1_14_inv17 = 1;
    95: op1_14_inv17 = 1;
    96: op1_14_inv17 = 1;
    default: op1_14_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in18 = reg_0517;
    6: op1_14_in18 = reg_0315;
    7: op1_14_in18 = reg_0359;
    8: op1_14_in18 = reg_0530;
    9: op1_14_in18 = reg_0465;
    10: op1_14_in18 = reg_0780;
    11: op1_14_in18 = reg_0395;
    12: op1_14_in18 = reg_0488;
    13: op1_14_in18 = reg_0073;
    14: op1_14_in18 = reg_0528;
    42: op1_14_in18 = reg_0528;
    15: op1_14_in18 = reg_0145;
    16: op1_14_in18 = reg_0205;
    17: op1_14_in18 = reg_0089;
    18: op1_14_in18 = reg_0239;
    19: op1_14_in18 = reg_0083;
    58: op1_14_in18 = reg_0083;
    72: op1_14_in18 = reg_0083;
    20: op1_14_in18 = reg_0478;
    21: op1_14_in18 = imem04_in[47:44];
    22: op1_14_in18 = reg_0134;
    23: op1_14_in18 = reg_0230;
    24: op1_14_in18 = reg_0441;
    25: op1_14_in18 = reg_0191;
    26: op1_14_in18 = reg_0944;
    27: op1_14_in18 = imem02_in[91:88];
    28: op1_14_in18 = reg_0266;
    29: op1_14_in18 = imem06_in[103:100];
    30: op1_14_in18 = imem01_in[63:60];
    31: op1_14_in18 = reg_1016;
    32: op1_14_in18 = reg_0951;
    33: op1_14_in18 = reg_0616;
    34: op1_14_in18 = reg_0394;
    35: op1_14_in18 = reg_1000;
    36: op1_14_in18 = reg_0277;
    37: op1_14_in18 = reg_0388;
    38: op1_14_in18 = imem06_in[31:28];
    41: op1_14_in18 = reg_0196;
    77: op1_14_in18 = reg_0196;
    83: op1_14_in18 = reg_0196;
    43: op1_14_in18 = reg_0270;
    44: op1_14_in18 = reg_0185;
    45: op1_14_in18 = imem02_in[59:56];
    46: op1_14_in18 = reg_0257;
    47: op1_14_in18 = reg_0180;
    48: op1_14_in18 = reg_0516;
    49: op1_14_in18 = reg_0980;
    50: op1_14_in18 = reg_0654;
    51: op1_14_in18 = reg_0211;
    52: op1_14_in18 = reg_0717;
    53: op1_14_in18 = reg_0919;
    54: op1_14_in18 = reg_0210;
    55: op1_14_in18 = reg_0940;
    56: op1_14_in18 = imem04_in[71:68];
    57: op1_14_in18 = reg_0306;
    59: op1_14_in18 = imem06_in[7:4];
    60: op1_14_in18 = imem04_in[31:28];
    61: op1_14_in18 = reg_0146;
    63: op1_14_in18 = reg_0358;
    64: op1_14_in18 = reg_0837;
    65: op1_14_in18 = reg_0840;
    66: op1_14_in18 = imem04_in[39:36];
    67: op1_14_in18 = imem03_in[123:120];
    68: op1_14_in18 = reg_0711;
    69: op1_14_in18 = imem01_in[43:40];
    70: op1_14_in18 = reg_1003;
    71: op1_14_in18 = reg_0433;
    73: op1_14_in18 = reg_0983;
    74: op1_14_in18 = reg_0777;
    75: op1_14_in18 = reg_0819;
    76: op1_14_in18 = imem07_in[87:84];
    78: op1_14_in18 = reg_0776;
    79: op1_14_in18 = reg_0506;
    80: op1_14_in18 = imem05_in[3:0];
    81: op1_14_in18 = reg_0448;
    82: op1_14_in18 = reg_0608;
    85: op1_14_in18 = reg_0507;
    86: op1_14_in18 = reg_0978;
    87: op1_14_in18 = imem01_in[95:92];
    88: op1_14_in18 = imem04_in[67:64];
    89: op1_14_in18 = imem01_in[103:100];
    90: op1_14_in18 = reg_0092;
    91: op1_14_in18 = reg_0713;
    92: op1_14_in18 = reg_0720;
    95: op1_14_in18 = imem07_in[95:92];
    96: op1_14_in18 = imem07_in[23:20];
    default: op1_14_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_14_inv18 = 1;
    9: op1_14_inv18 = 1;
    15: op1_14_inv18 = 1;
    16: op1_14_inv18 = 1;
    17: op1_14_inv18 = 1;
    21: op1_14_inv18 = 1;
    22: op1_14_inv18 = 1;
    26: op1_14_inv18 = 1;
    28: op1_14_inv18 = 1;
    29: op1_14_inv18 = 1;
    31: op1_14_inv18 = 1;
    32: op1_14_inv18 = 1;
    34: op1_14_inv18 = 1;
    38: op1_14_inv18 = 1;
    42: op1_14_inv18 = 1;
    45: op1_14_inv18 = 1;
    47: op1_14_inv18 = 1;
    49: op1_14_inv18 = 1;
    50: op1_14_inv18 = 1;
    51: op1_14_inv18 = 1;
    52: op1_14_inv18 = 1;
    53: op1_14_inv18 = 1;
    56: op1_14_inv18 = 1;
    58: op1_14_inv18 = 1;
    59: op1_14_inv18 = 1;
    63: op1_14_inv18 = 1;
    66: op1_14_inv18 = 1;
    72: op1_14_inv18 = 1;
    73: op1_14_inv18 = 1;
    78: op1_14_inv18 = 1;
    79: op1_14_inv18 = 1;
    80: op1_14_inv18 = 1;
    83: op1_14_inv18 = 1;
    86: op1_14_inv18 = 1;
    87: op1_14_inv18 = 1;
    88: op1_14_inv18 = 1;
    90: op1_14_inv18 = 1;
    default: op1_14_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in19 = reg_0518;
    6: op1_14_in19 = reg_0337;
    7: op1_14_in19 = reg_0318;
    8: op1_14_in19 = reg_0528;
    9: op1_14_in19 = reg_0464;
    10: op1_14_in19 = reg_0783;
    11: op1_14_in19 = reg_0360;
    12: op1_14_in19 = reg_0785;
    13: op1_14_in19 = reg_0079;
    14: op1_14_in19 = reg_0555;
    15: op1_14_in19 = reg_0140;
    16: op1_14_in19 = reg_0202;
    17: op1_14_in19 = reg_0085;
    18: op1_14_in19 = reg_0766;
    19: op1_14_in19 = reg_0088;
    20: op1_14_in19 = reg_0214;
    21: op1_14_in19 = imem04_in[55:52];
    22: op1_14_in19 = imem06_in[39:36];
    23: op1_14_in19 = reg_1015;
    24: op1_14_in19 = reg_0430;
    25: op1_14_in19 = reg_0209;
    26: op1_14_in19 = reg_0900;
    27: op1_14_in19 = imem02_in[107:104];
    28: op1_14_in19 = reg_0586;
    29: op1_14_in19 = imem06_in[127:124];
    30: op1_14_in19 = imem01_in[67:64];
    31: op1_14_in19 = reg_0537;
    32: op1_14_in19 = reg_0942;
    33: op1_14_in19 = reg_0611;
    34: op1_14_in19 = reg_0576;
    35: op1_14_in19 = reg_0994;
    36: op1_14_in19 = reg_0055;
    37: op1_14_in19 = reg_0000;
    38: op1_14_in19 = imem06_in[47:44];
    41: op1_14_in19 = reg_0195;
    83: op1_14_in19 = reg_0195;
    42: op1_14_in19 = reg_0517;
    43: op1_14_in19 = reg_0637;
    45: op1_14_in19 = reg_0863;
    46: op1_14_in19 = reg_0489;
    47: op1_14_in19 = reg_0177;
    48: op1_14_in19 = reg_0772;
    49: op1_14_in19 = reg_0974;
    50: op1_14_in19 = reg_0359;
    63: op1_14_in19 = reg_0359;
    51: op1_14_in19 = reg_0201;
    52: op1_14_in19 = reg_0718;
    53: op1_14_in19 = reg_1056;
    54: op1_14_in19 = reg_0204;
    55: op1_14_in19 = reg_0678;
    56: op1_14_in19 = imem04_in[83:80];
    57: op1_14_in19 = reg_0539;
    58: op1_14_in19 = reg_0482;
    59: op1_14_in19 = imem06_in[55:52];
    60: op1_14_in19 = imem04_in[39:36];
    61: op1_14_in19 = reg_0154;
    64: op1_14_in19 = reg_0052;
    65: op1_14_in19 = reg_0872;
    66: op1_14_in19 = imem04_in[47:44];
    67: op1_14_in19 = imem03_in[127:124];
    68: op1_14_in19 = reg_0701;
    69: op1_14_in19 = imem01_in[71:68];
    70: op1_14_in19 = reg_0048;
    71: op1_14_in19 = reg_0315;
    72: op1_14_in19 = reg_0261;
    73: op1_14_in19 = reg_0997;
    74: op1_14_in19 = reg_0251;
    75: op1_14_in19 = reg_0972;
    76: op1_14_in19 = imem07_in[91:88];
    77: op1_14_in19 = imem01_in[19:16];
    78: op1_14_in19 = reg_0506;
    79: op1_14_in19 = imem03_in[19:16];
    80: op1_14_in19 = imem05_in[23:20];
    81: op1_14_in19 = reg_0963;
    82: op1_14_in19 = reg_0776;
    85: op1_14_in19 = reg_0909;
    86: op1_14_in19 = reg_1000;
    87: op1_14_in19 = reg_1014;
    88: op1_14_in19 = imem04_in[91:88];
    89: op1_14_in19 = imem01_in[127:124];
    90: op1_14_in19 = reg_0761;
    91: op1_14_in19 = reg_0367;
    92: op1_14_in19 = reg_0726;
    95: op1_14_in19 = imem07_in[119:116];
    96: op1_14_in19 = imem07_in[79:76];
    default: op1_14_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv19 = 1;
    7: op1_14_inv19 = 1;
    8: op1_14_inv19 = 1;
    10: op1_14_inv19 = 1;
    11: op1_14_inv19 = 1;
    12: op1_14_inv19 = 1;
    15: op1_14_inv19 = 1;
    16: op1_14_inv19 = 1;
    17: op1_14_inv19 = 1;
    21: op1_14_inv19 = 1;
    22: op1_14_inv19 = 1;
    23: op1_14_inv19 = 1;
    25: op1_14_inv19 = 1;
    26: op1_14_inv19 = 1;
    29: op1_14_inv19 = 1;
    30: op1_14_inv19 = 1;
    31: op1_14_inv19 = 1;
    34: op1_14_inv19 = 1;
    37: op1_14_inv19 = 1;
    38: op1_14_inv19 = 1;
    41: op1_14_inv19 = 1;
    42: op1_14_inv19 = 1;
    45: op1_14_inv19 = 1;
    47: op1_14_inv19 = 1;
    48: op1_14_inv19 = 1;
    49: op1_14_inv19 = 1;
    50: op1_14_inv19 = 1;
    51: op1_14_inv19 = 1;
    53: op1_14_inv19 = 1;
    54: op1_14_inv19 = 1;
    57: op1_14_inv19 = 1;
    58: op1_14_inv19 = 1;
    65: op1_14_inv19 = 1;
    66: op1_14_inv19 = 1;
    70: op1_14_inv19 = 1;
    71: op1_14_inv19 = 1;
    72: op1_14_inv19 = 1;
    79: op1_14_inv19 = 1;
    80: op1_14_inv19 = 1;
    83: op1_14_inv19 = 1;
    88: op1_14_inv19 = 1;
    89: op1_14_inv19 = 1;
    90: op1_14_inv19 = 1;
    91: op1_14_inv19 = 1;
    92: op1_14_inv19 = 1;
    default: op1_14_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in20 = reg_0498;
    6: op1_14_in20 = reg_0027;
    29: op1_14_in20 = reg_0027;
    7: op1_14_in20 = reg_0330;
    8: op1_14_in20 = reg_0546;
    9: op1_14_in20 = reg_0469;
    10: op1_14_in20 = reg_0754;
    11: op1_14_in20 = reg_0319;
    12: op1_14_in20 = reg_0973;
    13: op1_14_in20 = imem03_in[19:16];
    14: op1_14_in20 = reg_0304;
    15: op1_14_in20 = reg_0134;
    16: op1_14_in20 = reg_0199;
    17: op1_14_in20 = reg_0077;
    18: op1_14_in20 = reg_1052;
    19: op1_14_in20 = reg_0089;
    48: op1_14_in20 = reg_0089;
    20: op1_14_in20 = reg_0191;
    21: op1_14_in20 = imem04_in[59:56];
    22: op1_14_in20 = imem06_in[59:56];
    23: op1_14_in20 = reg_0228;
    24: op1_14_in20 = reg_0436;
    25: op1_14_in20 = reg_0207;
    26: op1_14_in20 = reg_0256;
    27: op1_14_in20 = reg_0642;
    28: op1_14_in20 = reg_0592;
    30: op1_14_in20 = imem01_in[87:84];
    31: op1_14_in20 = reg_0061;
    32: op1_14_in20 = reg_0952;
    33: op1_14_in20 = reg_0627;
    34: op1_14_in20 = reg_0051;
    35: op1_14_in20 = imem04_in[11:8];
    36: op1_14_in20 = reg_1057;
    56: op1_14_in20 = reg_1057;
    57: op1_14_in20 = reg_1057;
    37: op1_14_in20 = imem06_in[3:0];
    38: op1_14_in20 = imem06_in[115:112];
    41: op1_14_in20 = reg_1034;
    42: op1_14_in20 = reg_0773;
    43: op1_14_in20 = reg_0704;
    45: op1_14_in20 = reg_0095;
    46: op1_14_in20 = reg_0132;
    47: op1_14_in20 = reg_0185;
    49: op1_14_in20 = reg_0663;
    50: op1_14_in20 = reg_0656;
    51: op1_14_in20 = reg_0213;
    54: op1_14_in20 = reg_0213;
    52: op1_14_in20 = reg_0701;
    53: op1_14_in20 = reg_1036;
    55: op1_14_in20 = reg_0734;
    58: op1_14_in20 = reg_0876;
    82: op1_14_in20 = reg_0876;
    59: op1_14_in20 = imem06_in[79:76];
    60: op1_14_in20 = imem04_in[43:40];
    61: op1_14_in20 = reg_0387;
    63: op1_14_in20 = reg_0087;
    64: op1_14_in20 = reg_0329;
    65: op1_14_in20 = imem03_in[35:32];
    66: op1_14_in20 = imem04_in[79:76];
    67: op1_14_in20 = reg_0099;
    68: op1_14_in20 = reg_0575;
    69: op1_14_in20 = imem01_in[79:76];
    70: op1_14_in20 = reg_0888;
    71: op1_14_in20 = reg_0838;
    72: op1_14_in20 = reg_0872;
    73: op1_14_in20 = imem04_in[15:12];
    74: op1_14_in20 = reg_0542;
    75: op1_14_in20 = reg_0780;
    76: op1_14_in20 = imem07_in[103:100];
    77: op1_14_in20 = imem01_in[39:36];
    78: op1_14_in20 = reg_0484;
    79: op1_14_in20 = imem03_in[43:40];
    80: op1_14_in20 = imem05_in[35:32];
    81: op1_14_in20 = reg_0525;
    83: op1_14_in20 = imem01_in[7:4];
    85: op1_14_in20 = reg_0524;
    86: op1_14_in20 = imem04_in[27:24];
    87: op1_14_in20 = reg_1022;
    88: op1_14_in20 = imem04_in[127:124];
    89: op1_14_in20 = reg_0610;
    90: op1_14_in20 = reg_0007;
    91: op1_14_in20 = imem03_in[15:12];
    92: op1_14_in20 = reg_0560;
    95: op1_14_in20 = reg_0721;
    96: op1_14_in20 = imem07_in[111:108];
    default: op1_14_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv20 = 1;
    8: op1_14_inv20 = 1;
    11: op1_14_inv20 = 1;
    12: op1_14_inv20 = 1;
    18: op1_14_inv20 = 1;
    19: op1_14_inv20 = 1;
    20: op1_14_inv20 = 1;
    22: op1_14_inv20 = 1;
    26: op1_14_inv20 = 1;
    27: op1_14_inv20 = 1;
    29: op1_14_inv20 = 1;
    31: op1_14_inv20 = 1;
    34: op1_14_inv20 = 1;
    35: op1_14_inv20 = 1;
    36: op1_14_inv20 = 1;
    38: op1_14_inv20 = 1;
    41: op1_14_inv20 = 1;
    42: op1_14_inv20 = 1;
    45: op1_14_inv20 = 1;
    47: op1_14_inv20 = 1;
    51: op1_14_inv20 = 1;
    53: op1_14_inv20 = 1;
    54: op1_14_inv20 = 1;
    58: op1_14_inv20 = 1;
    59: op1_14_inv20 = 1;
    60: op1_14_inv20 = 1;
    61: op1_14_inv20 = 1;
    63: op1_14_inv20 = 1;
    66: op1_14_inv20 = 1;
    67: op1_14_inv20 = 1;
    68: op1_14_inv20 = 1;
    69: op1_14_inv20 = 1;
    70: op1_14_inv20 = 1;
    71: op1_14_inv20 = 1;
    74: op1_14_inv20 = 1;
    75: op1_14_inv20 = 1;
    79: op1_14_inv20 = 1;
    80: op1_14_inv20 = 1;
    81: op1_14_inv20 = 1;
    82: op1_14_inv20 = 1;
    85: op1_14_inv20 = 1;
    86: op1_14_inv20 = 1;
    87: op1_14_inv20 = 1;
    89: op1_14_inv20 = 1;
    90: op1_14_inv20 = 1;
    91: op1_14_inv20 = 1;
    92: op1_14_inv20 = 1;
    95: op1_14_inv20 = 1;
    default: op1_14_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in21 = reg_0233;
    6: op1_14_in21 = reg_0020;
    7: op1_14_in21 = reg_0363;
    8: op1_14_in21 = reg_0559;
    9: op1_14_in21 = reg_0476;
    10: op1_14_in21 = imem07_in[11:8];
    11: op1_14_in21 = reg_0312;
    12: op1_14_in21 = reg_0955;
    13: op1_14_in21 = imem03_in[31:28];
    17: op1_14_in21 = imem03_in[31:28];
    14: op1_14_in21 = reg_0061;
    36: op1_14_in21 = reg_0061;
    15: op1_14_in21 = imem06_in[39:36];
    16: op1_14_in21 = imem01_in[15:12];
    18: op1_14_in21 = reg_1039;
    19: op1_14_in21 = reg_0090;
    20: op1_14_in21 = reg_0189;
    21: op1_14_in21 = imem04_in[87:84];
    66: op1_14_in21 = imem04_in[87:84];
    22: op1_14_in21 = imem06_in[103:100];
    23: op1_14_in21 = reg_1038;
    24: op1_14_in21 = reg_0423;
    25: op1_14_in21 = reg_0197;
    26: op1_14_in21 = reg_0251;
    27: op1_14_in21 = reg_0654;
    28: op1_14_in21 = reg_0591;
    29: op1_14_in21 = reg_0801;
    30: op1_14_in21 = reg_0786;
    31: op1_14_in21 = reg_0733;
    32: op1_14_in21 = reg_0215;
    33: op1_14_in21 = reg_0615;
    34: op1_14_in21 = reg_0376;
    35: op1_14_in21 = imem04_in[19:16];
    37: op1_14_in21 = imem06_in[51:48];
    38: op1_14_in21 = reg_0027;
    41: op1_14_in21 = reg_0235;
    42: op1_14_in21 = reg_0286;
    43: op1_14_in21 = reg_0726;
    45: op1_14_in21 = reg_0096;
    46: op1_14_in21 = reg_0147;
    47: op1_14_in21 = reg_0176;
    48: op1_14_in21 = reg_0867;
    49: op1_14_in21 = reg_0012;
    50: op1_14_in21 = reg_0082;
    51: op1_14_in21 = reg_0196;
    52: op1_14_in21 = reg_0805;
    53: op1_14_in21 = reg_0285;
    54: op1_14_in21 = reg_0205;
    55: op1_14_in21 = imem03_in[3:0];
    72: op1_14_in21 = imem03_in[3:0];
    56: op1_14_in21 = reg_0541;
    57: op1_14_in21 = reg_0888;
    58: op1_14_in21 = reg_0084;
    59: op1_14_in21 = imem06_in[111:108];
    60: op1_14_in21 = imem04_in[67:64];
    61: op1_14_in21 = reg_0787;
    63: op1_14_in21 = reg_0516;
    64: op1_14_in21 = reg_0347;
    65: op1_14_in21 = imem03_in[39:36];
    67: op1_14_in21 = reg_0228;
    68: op1_14_in21 = reg_0250;
    69: op1_14_in21 = imem01_in[95:92];
    70: op1_14_in21 = reg_0931;
    71: op1_14_in21 = reg_0185;
    73: op1_14_in21 = imem04_in[27:24];
    74: op1_14_in21 = reg_0042;
    75: op1_14_in21 = reg_0135;
    76: op1_14_in21 = imem07_in[107:104];
    77: op1_14_in21 = imem01_in[83:80];
    78: op1_14_in21 = reg_0291;
    79: op1_14_in21 = imem03_in[71:68];
    80: op1_14_in21 = imem05_in[115:112];
    81: op1_14_in21 = reg_0314;
    82: op1_14_in21 = reg_0086;
    83: op1_14_in21 = imem01_in[19:16];
    85: op1_14_in21 = reg_0401;
    86: op1_14_in21 = imem04_in[35:32];
    87: op1_14_in21 = reg_0234;
    88: op1_14_in21 = reg_0430;
    89: op1_14_in21 = reg_1017;
    90: op1_14_in21 = reg_0301;
    91: op1_14_in21 = imem03_in[27:24];
    92: op1_14_in21 = reg_0164;
    95: op1_14_in21 = reg_0374;
    96: op1_14_in21 = imem07_in[115:112];
    default: op1_14_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv21 = 1;
    7: op1_14_inv21 = 1;
    9: op1_14_inv21 = 1;
    11: op1_14_inv21 = 1;
    13: op1_14_inv21 = 1;
    15: op1_14_inv21 = 1;
    16: op1_14_inv21 = 1;
    18: op1_14_inv21 = 1;
    19: op1_14_inv21 = 1;
    20: op1_14_inv21 = 1;
    21: op1_14_inv21 = 1;
    23: op1_14_inv21 = 1;
    24: op1_14_inv21 = 1;
    25: op1_14_inv21 = 1;
    29: op1_14_inv21 = 1;
    30: op1_14_inv21 = 1;
    32: op1_14_inv21 = 1;
    34: op1_14_inv21 = 1;
    35: op1_14_inv21 = 1;
    37: op1_14_inv21 = 1;
    43: op1_14_inv21 = 1;
    48: op1_14_inv21 = 1;
    54: op1_14_inv21 = 1;
    55: op1_14_inv21 = 1;
    56: op1_14_inv21 = 1;
    57: op1_14_inv21 = 1;
    60: op1_14_inv21 = 1;
    61: op1_14_inv21 = 1;
    63: op1_14_inv21 = 1;
    64: op1_14_inv21 = 1;
    65: op1_14_inv21 = 1;
    66: op1_14_inv21 = 1;
    68: op1_14_inv21 = 1;
    69: op1_14_inv21 = 1;
    74: op1_14_inv21 = 1;
    75: op1_14_inv21 = 1;
    76: op1_14_inv21 = 1;
    77: op1_14_inv21 = 1;
    78: op1_14_inv21 = 1;
    79: op1_14_inv21 = 1;
    81: op1_14_inv21 = 1;
    82: op1_14_inv21 = 1;
    83: op1_14_inv21 = 1;
    86: op1_14_inv21 = 1;
    89: op1_14_inv21 = 1;
    91: op1_14_inv21 = 1;
    default: op1_14_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in22 = reg_0228;
    6: op1_14_in22 = reg_0024;
    7: op1_14_in22 = reg_0086;
    8: op1_14_in22 = reg_0531;
    9: op1_14_in22 = reg_0466;
    10: op1_14_in22 = imem07_in[43:40];
    11: op1_14_in22 = reg_0985;
    12: op1_14_in22 = reg_0957;
    13: op1_14_in22 = imem03_in[35:32];
    14: op1_14_in22 = reg_0047;
    15: op1_14_in22 = imem06_in[87:84];
    16: op1_14_in22 = imem01_in[59:56];
    17: op1_14_in22 = imem03_in[87:84];
    18: op1_14_in22 = reg_1042;
    19: op1_14_in22 = reg_0091;
    20: op1_14_in22 = reg_0211;
    21: op1_14_in22 = imem04_in[91:88];
    22: op1_14_in22 = imem06_in[123:120];
    23: op1_14_in22 = reg_0122;
    24: op1_14_in22 = reg_0440;
    25: op1_14_in22 = reg_0307;
    26: op1_14_in22 = reg_0257;
    27: op1_14_in22 = reg_0656;
    28: op1_14_in22 = reg_0585;
    29: op1_14_in22 = reg_0781;
    30: op1_14_in22 = reg_0563;
    31: op1_14_in22 = reg_0078;
    32: op1_14_in22 = reg_0900;
    33: op1_14_in22 = reg_0612;
    34: op1_14_in22 = reg_0312;
    35: op1_14_in22 = imem04_in[99:96];
    36: op1_14_in22 = reg_0760;
    37: op1_14_in22 = imem07_in[31:28];
    38: op1_14_in22 = reg_0408;
    41: op1_14_in22 = reg_0544;
    42: op1_14_in22 = imem05_in[15:12];
    43: op1_14_in22 = reg_0714;
    45: op1_14_in22 = reg_0097;
    46: op1_14_in22 = reg_0150;
    47: op1_14_in22 = reg_0184;
    48: op1_14_in22 = reg_0814;
    49: op1_14_in22 = reg_0855;
    50: op1_14_in22 = reg_0045;
    51: op1_14_in22 = imem01_in[39:36];
    52: op1_14_in22 = reg_0361;
    53: op1_14_in22 = reg_0253;
    54: op1_14_in22 = reg_0192;
    55: op1_14_in22 = imem03_in[7:4];
    56: op1_14_in22 = reg_0507;
    57: op1_14_in22 = reg_0799;
    58: op1_14_in22 = imem03_in[11:8];
    59: op1_14_in22 = reg_0660;
    60: op1_14_in22 = imem04_in[95:92];
    61: op1_14_in22 = reg_0783;
    63: op1_14_in22 = reg_0007;
    64: op1_14_in22 = reg_0758;
    65: op1_14_in22 = imem03_in[43:40];
    66: op1_14_in22 = imem04_in[107:104];
    67: op1_14_in22 = reg_1007;
    68: op1_14_in22 = reg_0353;
    69: op1_14_in22 = reg_0798;
    70: op1_14_in22 = reg_0541;
    71: op1_14_in22 = reg_0171;
    72: op1_14_in22 = imem03_in[83:80];
    79: op1_14_in22 = imem03_in[83:80];
    73: op1_14_in22 = imem04_in[59:56];
    74: op1_14_in22 = reg_0958;
    75: op1_14_in22 = reg_0965;
    76: op1_14_in22 = imem07_in[119:116];
    96: op1_14_in22 = imem07_in[119:116];
    77: op1_14_in22 = imem01_in[115:112];
    78: op1_14_in22 = imem03_in[3:0];
    80: op1_14_in22 = reg_0217;
    81: op1_14_in22 = reg_0892;
    82: op1_14_in22 = reg_0090;
    83: op1_14_in22 = imem01_in[23:20];
    85: op1_14_in22 = reg_0015;
    86: op1_14_in22 = imem04_in[43:40];
    87: op1_14_in22 = reg_0225;
    88: op1_14_in22 = reg_0848;
    89: op1_14_in22 = reg_0304;
    90: op1_14_in22 = reg_0331;
    91: op1_14_in22 = imem03_in[47:44];
    92: op1_14_in22 = reg_0653;
    95: op1_14_in22 = reg_0708;
    default: op1_14_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv22 = 1;
    6: op1_14_inv22 = 1;
    7: op1_14_inv22 = 1;
    10: op1_14_inv22 = 1;
    13: op1_14_inv22 = 1;
    15: op1_14_inv22 = 1;
    17: op1_14_inv22 = 1;
    25: op1_14_inv22 = 1;
    27: op1_14_inv22 = 1;
    30: op1_14_inv22 = 1;
    31: op1_14_inv22 = 1;
    32: op1_14_inv22 = 1;
    35: op1_14_inv22 = 1;
    36: op1_14_inv22 = 1;
    37: op1_14_inv22 = 1;
    46: op1_14_inv22 = 1;
    47: op1_14_inv22 = 1;
    52: op1_14_inv22 = 1;
    53: op1_14_inv22 = 1;
    55: op1_14_inv22 = 1;
    58: op1_14_inv22 = 1;
    61: op1_14_inv22 = 1;
    63: op1_14_inv22 = 1;
    64: op1_14_inv22 = 1;
    65: op1_14_inv22 = 1;
    66: op1_14_inv22 = 1;
    68: op1_14_inv22 = 1;
    70: op1_14_inv22 = 1;
    75: op1_14_inv22 = 1;
    82: op1_14_inv22 = 1;
    88: op1_14_inv22 = 1;
    89: op1_14_inv22 = 1;
    90: op1_14_inv22 = 1;
    91: op1_14_inv22 = 1;
    95: op1_14_inv22 = 1;
    96: op1_14_inv22 = 1;
    default: op1_14_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in23 = reg_0221;
    6: op1_14_in23 = reg_0023;
    7: op1_14_in23 = reg_0090;
    8: op1_14_in23 = reg_0556;
    9: op1_14_in23 = reg_0472;
    10: op1_14_in23 = imem07_in[55:52];
    11: op1_14_in23 = reg_0978;
    12: op1_14_in23 = reg_0964;
    13: op1_14_in23 = imem03_in[83:80];
    14: op1_14_in23 = reg_0078;
    15: op1_14_in23 = imem06_in[123:120];
    16: op1_14_in23 = imem01_in[63:60];
    17: op1_14_in23 = imem03_in[99:96];
    18: op1_14_in23 = reg_1045;
    19: op1_14_in23 = reg_0084;
    20: op1_14_in23 = reg_0196;
    21: op1_14_in23 = reg_0543;
    67: op1_14_in23 = reg_0543;
    22: op1_14_in23 = reg_0614;
    23: op1_14_in23 = reg_0125;
    24: op1_14_in23 = reg_0444;
    25: op1_14_in23 = reg_0926;
    26: op1_14_in23 = reg_1046;
    27: op1_14_in23 = reg_0640;
    28: op1_14_in23 = reg_0576;
    29: op1_14_in23 = reg_1010;
    30: op1_14_in23 = reg_0811;
    31: op1_14_in23 = reg_0760;
    32: op1_14_in23 = reg_0229;
    33: op1_14_in23 = reg_0914;
    34: op1_14_in23 = reg_0246;
    35: op1_14_in23 = reg_0536;
    36: op1_14_in23 = reg_0755;
    37: op1_14_in23 = imem07_in[51:48];
    38: op1_14_in23 = reg_0558;
    41: op1_14_in23 = imem01_in[95:92];
    42: op1_14_in23 = imem05_in[35:32];
    43: op1_14_in23 = reg_0707;
    45: op1_14_in23 = reg_0335;
    46: op1_14_in23 = reg_0128;
    47: op1_14_in23 = reg_0502;
    48: op1_14_in23 = reg_0506;
    49: op1_14_in23 = reg_0512;
    50: op1_14_in23 = reg_0842;
    51: op1_14_in23 = imem01_in[43:40];
    52: op1_14_in23 = reg_0420;
    53: op1_14_in23 = reg_0607;
    54: op1_14_in23 = imem01_in[3:0];
    55: op1_14_in23 = imem03_in[15:12];
    56: op1_14_in23 = reg_0524;
    57: op1_14_in23 = reg_0802;
    58: op1_14_in23 = imem03_in[23:20];
    59: op1_14_in23 = reg_0384;
    60: op1_14_in23 = imem04_in[119:116];
    61: op1_14_in23 = reg_0320;
    63: op1_14_in23 = reg_0758;
    64: op1_14_in23 = reg_0876;
    65: op1_14_in23 = imem03_in[51:48];
    66: op1_14_in23 = imem04_in[127:124];
    68: op1_14_in23 = reg_0350;
    69: op1_14_in23 = reg_0604;
    70: op1_14_in23 = reg_0537;
    72: op1_14_in23 = imem03_in[87:84];
    73: op1_14_in23 = imem04_in[67:64];
    74: op1_14_in23 = reg_0131;
    75: op1_14_in23 = imem06_in[63:60];
    76: op1_14_in23 = imem07_in[123:120];
    96: op1_14_in23 = imem07_in[123:120];
    77: op1_14_in23 = reg_0969;
    78: op1_14_in23 = imem03_in[63:60];
    79: op1_14_in23 = reg_0535;
    80: op1_14_in23 = reg_0655;
    81: op1_14_in23 = reg_0153;
    82: op1_14_in23 = reg_0091;
    83: op1_14_in23 = imem01_in[27:24];
    85: op1_14_in23 = reg_0064;
    86: op1_14_in23 = imem04_in[63:60];
    87: op1_14_in23 = reg_0869;
    88: op1_14_in23 = reg_0808;
    89: op1_14_in23 = reg_0615;
    90: op1_14_in23 = reg_0397;
    91: op1_14_in23 = reg_0859;
    92: op1_14_in23 = reg_0744;
    95: op1_14_in23 = reg_0718;
    default: op1_14_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_14_inv23 = 1;
    8: op1_14_inv23 = 1;
    9: op1_14_inv23 = 1;
    11: op1_14_inv23 = 1;
    12: op1_14_inv23 = 1;
    13: op1_14_inv23 = 1;
    14: op1_14_inv23 = 1;
    15: op1_14_inv23 = 1;
    16: op1_14_inv23 = 1;
    17: op1_14_inv23 = 1;
    19: op1_14_inv23 = 1;
    21: op1_14_inv23 = 1;
    27: op1_14_inv23 = 1;
    29: op1_14_inv23 = 1;
    30: op1_14_inv23 = 1;
    33: op1_14_inv23 = 1;
    36: op1_14_inv23 = 1;
    37: op1_14_inv23 = 1;
    41: op1_14_inv23 = 1;
    42: op1_14_inv23 = 1;
    45: op1_14_inv23 = 1;
    51: op1_14_inv23 = 1;
    52: op1_14_inv23 = 1;
    53: op1_14_inv23 = 1;
    55: op1_14_inv23 = 1;
    56: op1_14_inv23 = 1;
    57: op1_14_inv23 = 1;
    58: op1_14_inv23 = 1;
    60: op1_14_inv23 = 1;
    63: op1_14_inv23 = 1;
    64: op1_14_inv23 = 1;
    65: op1_14_inv23 = 1;
    69: op1_14_inv23 = 1;
    70: op1_14_inv23 = 1;
    72: op1_14_inv23 = 1;
    77: op1_14_inv23 = 1;
    79: op1_14_inv23 = 1;
    80: op1_14_inv23 = 1;
    81: op1_14_inv23 = 1;
    83: op1_14_inv23 = 1;
    85: op1_14_inv23 = 1;
    86: op1_14_inv23 = 1;
    88: op1_14_inv23 = 1;
    89: op1_14_inv23 = 1;
    90: op1_14_inv23 = 1;
    91: op1_14_inv23 = 1;
    default: op1_14_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in24 = reg_0219;
    30: op1_14_in24 = reg_0219;
    6: op1_14_in24 = imem07_in[3:0];
    7: op1_14_in24 = reg_0051;
    8: op1_14_in24 = reg_0282;
    9: op1_14_in24 = reg_0467;
    10: op1_14_in24 = imem07_in[71:68];
    37: op1_14_in24 = imem07_in[71:68];
    11: op1_14_in24 = reg_0983;
    12: op1_14_in24 = reg_0953;
    13: op1_14_in24 = imem03_in[115:112];
    14: op1_14_in24 = reg_0058;
    15: op1_14_in24 = reg_0617;
    16: op1_14_in24 = imem01_in[91:88];
    17: op1_14_in24 = reg_0579;
    90: op1_14_in24 = reg_0579;
    18: op1_14_in24 = reg_0102;
    19: op1_14_in24 = reg_0087;
    20: op1_14_in24 = reg_0199;
    21: op1_14_in24 = reg_0557;
    22: op1_14_in24 = reg_0604;
    23: op1_14_in24 = reg_0120;
    24: op1_14_in24 = reg_0443;
    25: op1_14_in24 = reg_0928;
    26: op1_14_in24 = reg_0896;
    27: op1_14_in24 = reg_0636;
    28: op1_14_in24 = imem03_in[75:72];
    29: op1_14_in24 = reg_0783;
    31: op1_14_in24 = reg_0276;
    32: op1_14_in24 = reg_0251;
    33: op1_14_in24 = reg_0391;
    34: op1_14_in24 = reg_0374;
    35: op1_14_in24 = reg_0277;
    36: op1_14_in24 = reg_0069;
    38: op1_14_in24 = reg_0593;
    41: op1_14_in24 = imem01_in[115:112];
    42: op1_14_in24 = imem05_in[47:44];
    43: op1_14_in24 = reg_0701;
    45: op1_14_in24 = reg_0091;
    46: op1_14_in24 = reg_0138;
    48: op1_14_in24 = reg_0049;
    82: op1_14_in24 = reg_0049;
    49: op1_14_in24 = reg_0547;
    50: op1_14_in24 = reg_0039;
    51: op1_14_in24 = imem01_in[95:92];
    52: op1_14_in24 = reg_0640;
    53: op1_14_in24 = reg_0522;
    54: op1_14_in24 = imem01_in[19:16];
    55: op1_14_in24 = imem03_in[35:32];
    56: op1_14_in24 = reg_0850;
    57: op1_14_in24 = reg_0056;
    58: op1_14_in24 = imem03_in[31:28];
    59: op1_14_in24 = reg_0613;
    60: op1_14_in24 = reg_1003;
    61: op1_14_in24 = reg_0660;
    63: op1_14_in24 = reg_0089;
    64: op1_14_in24 = reg_0090;
    65: op1_14_in24 = imem03_in[67:64];
    78: op1_14_in24 = imem03_in[67:64];
    66: op1_14_in24 = reg_0530;
    67: op1_14_in24 = reg_0833;
    68: op1_14_in24 = reg_0172;
    69: op1_14_in24 = reg_0520;
    87: op1_14_in24 = reg_0520;
    70: op1_14_in24 = reg_0507;
    72: op1_14_in24 = reg_0006;
    73: op1_14_in24 = imem04_in[83:80];
    74: op1_14_in24 = reg_0944;
    75: op1_14_in24 = imem06_in[83:80];
    76: op1_14_in24 = reg_0667;
    77: op1_14_in24 = reg_1032;
    79: op1_14_in24 = reg_0681;
    80: op1_14_in24 = reg_0139;
    81: op1_14_in24 = reg_0952;
    83: op1_14_in24 = imem01_in[51:48];
    85: op1_14_in24 = reg_0027;
    86: op1_14_in24 = imem04_in[75:72];
    88: op1_14_in24 = reg_0041;
    89: op1_14_in24 = reg_0555;
    91: op1_14_in24 = reg_0317;
    92: op1_14_in24 = reg_0502;
    95: op1_14_in24 = reg_0759;
    96: op1_14_in24 = reg_0165;
    default: op1_14_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv24 = 1;
    7: op1_14_inv24 = 1;
    10: op1_14_inv24 = 1;
    12: op1_14_inv24 = 1;
    13: op1_14_inv24 = 1;
    16: op1_14_inv24 = 1;
    18: op1_14_inv24 = 1;
    19: op1_14_inv24 = 1;
    22: op1_14_inv24 = 1;
    24: op1_14_inv24 = 1;
    25: op1_14_inv24 = 1;
    29: op1_14_inv24 = 1;
    30: op1_14_inv24 = 1;
    31: op1_14_inv24 = 1;
    33: op1_14_inv24 = 1;
    34: op1_14_inv24 = 1;
    35: op1_14_inv24 = 1;
    36: op1_14_inv24 = 1;
    38: op1_14_inv24 = 1;
    41: op1_14_inv24 = 1;
    43: op1_14_inv24 = 1;
    46: op1_14_inv24 = 1;
    49: op1_14_inv24 = 1;
    50: op1_14_inv24 = 1;
    51: op1_14_inv24 = 1;
    58: op1_14_inv24 = 1;
    59: op1_14_inv24 = 1;
    60: op1_14_inv24 = 1;
    64: op1_14_inv24 = 1;
    66: op1_14_inv24 = 1;
    73: op1_14_inv24 = 1;
    74: op1_14_inv24 = 1;
    75: op1_14_inv24 = 1;
    76: op1_14_inv24 = 1;
    78: op1_14_inv24 = 1;
    79: op1_14_inv24 = 1;
    81: op1_14_inv24 = 1;
    83: op1_14_inv24 = 1;
    86: op1_14_inv24 = 1;
    87: op1_14_inv24 = 1;
    89: op1_14_inv24 = 1;
    91: op1_14_inv24 = 1;
    92: op1_14_inv24 = 1;
    95: op1_14_inv24 = 1;
    96: op1_14_inv24 = 1;
    default: op1_14_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in25 = reg_0122;
    6: op1_14_in25 = imem07_in[23:20];
    7: op1_14_in25 = reg_0060;
    8: op1_14_in25 = reg_0306;
    9: op1_14_in25 = reg_0471;
    10: op1_14_in25 = imem07_in[95:92];
    11: op1_14_in25 = reg_0976;
    12: op1_14_in25 = imem05_in[15:12];
    13: op1_14_in25 = reg_0583;
    17: op1_14_in25 = reg_0583;
    14: op1_14_in25 = reg_0057;
    15: op1_14_in25 = reg_0612;
    16: op1_14_in25 = imem01_in[103:100];
    18: op1_14_in25 = reg_0101;
    89: op1_14_in25 = reg_0101;
    19: op1_14_in25 = reg_0093;
    20: op1_14_in25 = imem01_in[3:0];
    21: op1_14_in25 = reg_0553;
    22: op1_14_in25 = reg_0630;
    23: op1_14_in25 = reg_0113;
    24: op1_14_in25 = reg_0448;
    25: op1_14_in25 = reg_0521;
    26: op1_14_in25 = reg_0143;
    27: op1_14_in25 = reg_0663;
    28: op1_14_in25 = imem03_in[79:76];
    55: op1_14_in25 = imem03_in[79:76];
    29: op1_14_in25 = imem07_in[7:4];
    30: op1_14_in25 = reg_0249;
    31: op1_14_in25 = reg_0278;
    32: op1_14_in25 = reg_0489;
    33: op1_14_in25 = reg_0741;
    34: op1_14_in25 = reg_0996;
    35: op1_14_in25 = reg_0055;
    36: op1_14_in25 = reg_0009;
    37: op1_14_in25 = imem07_in[79:76];
    38: op1_14_in25 = reg_0925;
    41: op1_14_in25 = reg_0112;
    42: op1_14_in25 = imem05_in[67:64];
    43: op1_14_in25 = reg_0727;
    45: op1_14_in25 = reg_0016;
    46: op1_14_in25 = imem06_in[7:4];
    48: op1_14_in25 = imem03_in[35:32];
    49: op1_14_in25 = reg_1006;
    50: op1_14_in25 = reg_0096;
    51: op1_14_in25 = imem01_in[127:124];
    52: op1_14_in25 = reg_0838;
    53: op1_14_in25 = reg_0604;
    54: op1_14_in25 = imem01_in[55:52];
    56: op1_14_in25 = reg_0302;
    57: op1_14_in25 = reg_0815;
    58: op1_14_in25 = imem03_in[43:40];
    59: op1_14_in25 = reg_0533;
    60: op1_14_in25 = reg_1009;
    61: op1_14_in25 = reg_0692;
    63: op1_14_in25 = reg_0086;
    64: op1_14_in25 = imem03_in[3:0];
    65: op1_14_in25 = imem03_in[75:72];
    66: op1_14_in25 = reg_0511;
    67: op1_14_in25 = reg_0795;
    68: op1_14_in25 = reg_0179;
    69: op1_14_in25 = reg_0514;
    70: op1_14_in25 = reg_0752;
    72: op1_14_in25 = reg_0681;
    73: op1_14_in25 = imem04_in[91:88];
    74: op1_14_in25 = reg_0655;
    75: op1_14_in25 = imem06_in[99:96];
    76: op1_14_in25 = reg_0339;
    77: op1_14_in25 = reg_1014;
    78: op1_14_in25 = reg_0357;
    79: op1_14_in25 = reg_0445;
    80: op1_14_in25 = reg_0892;
    81: op1_14_in25 = reg_0819;
    82: op1_14_in25 = imem03_in[7:4];
    83: op1_14_in25 = imem01_in[87:84];
    85: op1_14_in25 = reg_0044;
    86: op1_14_in25 = reg_0147;
    87: op1_14_in25 = reg_0227;
    88: op1_14_in25 = reg_0108;
    90: op1_14_in25 = reg_0597;
    91: op1_14_in25 = reg_0307;
    92: op1_14_in25 = reg_0429;
    95: op1_14_in25 = reg_0805;
    96: op1_14_in25 = reg_0715;
    default: op1_14_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_14_inv25 = 1;
    9: op1_14_inv25 = 1;
    11: op1_14_inv25 = 1;
    12: op1_14_inv25 = 1;
    19: op1_14_inv25 = 1;
    22: op1_14_inv25 = 1;
    23: op1_14_inv25 = 1;
    24: op1_14_inv25 = 1;
    25: op1_14_inv25 = 1;
    26: op1_14_inv25 = 1;
    27: op1_14_inv25 = 1;
    28: op1_14_inv25 = 1;
    30: op1_14_inv25 = 1;
    36: op1_14_inv25 = 1;
    37: op1_14_inv25 = 1;
    41: op1_14_inv25 = 1;
    42: op1_14_inv25 = 1;
    46: op1_14_inv25 = 1;
    48: op1_14_inv25 = 1;
    49: op1_14_inv25 = 1;
    50: op1_14_inv25 = 1;
    51: op1_14_inv25 = 1;
    53: op1_14_inv25 = 1;
    61: op1_14_inv25 = 1;
    65: op1_14_inv25 = 1;
    66: op1_14_inv25 = 1;
    67: op1_14_inv25 = 1;
    69: op1_14_inv25 = 1;
    74: op1_14_inv25 = 1;
    79: op1_14_inv25 = 1;
    80: op1_14_inv25 = 1;
    81: op1_14_inv25 = 1;
    85: op1_14_inv25 = 1;
    90: op1_14_inv25 = 1;
    91: op1_14_inv25 = 1;
    95: op1_14_inv25 = 1;
    default: op1_14_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in26 = reg_0111;
    6: op1_14_in26 = imem07_in[39:36];
    7: op1_14_in26 = reg_0087;
    8: op1_14_in26 = reg_0293;
    9: op1_14_in26 = reg_0478;
    10: op1_14_in26 = reg_0721;
    11: op1_14_in26 = imem04_in[7:4];
    12: op1_14_in26 = imem05_in[31:28];
    85: op1_14_in26 = imem05_in[31:28];
    13: op1_14_in26 = reg_0587;
    14: op1_14_in26 = imem05_in[3:0];
    15: op1_14_in26 = reg_0348;
    16: op1_14_in26 = imem01_in[111:108];
    17: op1_14_in26 = reg_0563;
    18: op1_14_in26 = imem02_in[23:20];
    19: op1_14_in26 = imem03_in[11:8];
    20: op1_14_in26 = imem01_in[19:16];
    21: op1_14_in26 = reg_0550;
    86: op1_14_in26 = reg_0550;
    22: op1_14_in26 = reg_0611;
    23: op1_14_in26 = imem02_in[11:8];
    24: op1_14_in26 = reg_0175;
    25: op1_14_in26 = reg_0245;
    78: op1_14_in26 = reg_0245;
    26: op1_14_in26 = reg_0138;
    27: op1_14_in26 = reg_0045;
    28: op1_14_in26 = imem03_in[119:116];
    29: op1_14_in26 = imem07_in[11:8];
    30: op1_14_in26 = reg_0905;
    31: op1_14_in26 = reg_0054;
    32: op1_14_in26 = reg_0148;
    33: op1_14_in26 = reg_0388;
    34: op1_14_in26 = reg_0981;
    35: op1_14_in26 = reg_1057;
    36: op1_14_in26 = reg_0015;
    37: op1_14_in26 = imem07_in[83:80];
    38: op1_14_in26 = reg_0585;
    41: op1_14_in26 = reg_0115;
    42: op1_14_in26 = reg_0948;
    43: op1_14_in26 = imem07_in[15:12];
    45: op1_14_in26 = imem03_in[67:64];
    46: op1_14_in26 = imem06_in[19:16];
    48: op1_14_in26 = imem03_in[71:68];
    49: op1_14_in26 = reg_0265;
    66: op1_14_in26 = reg_0265;
    50: op1_14_in26 = reg_0330;
    51: op1_14_in26 = reg_0586;
    53: op1_14_in26 = reg_1043;
    54: op1_14_in26 = imem01_in[67:64];
    55: op1_14_in26 = imem03_in[103:100];
    56: op1_14_in26 = reg_0584;
    57: op1_14_in26 = reg_0064;
    58: op1_14_in26 = imem03_in[59:56];
    59: op1_14_in26 = reg_0382;
    60: op1_14_in26 = reg_0048;
    61: op1_14_in26 = reg_0534;
    63: op1_14_in26 = reg_0084;
    64: op1_14_in26 = imem03_in[99:96];
    65: op1_14_in26 = imem03_in[115:112];
    67: op1_14_in26 = reg_0807;
    68: op1_14_in26 = reg_0183;
    69: op1_14_in26 = reg_1017;
    70: op1_14_in26 = reg_0076;
    72: op1_14_in26 = reg_0760;
    73: op1_14_in26 = imem04_in[95:92];
    74: op1_14_in26 = reg_0143;
    75: op1_14_in26 = imem06_in[103:100];
    76: op1_14_in26 = reg_0677;
    77: op1_14_in26 = reg_0968;
    79: op1_14_in26 = reg_0307;
    80: op1_14_in26 = reg_0486;
    81: op1_14_in26 = reg_0972;
    82: op1_14_in26 = imem03_in[51:48];
    83: op1_14_in26 = imem01_in[91:88];
    87: op1_14_in26 = reg_1040;
    88: op1_14_in26 = reg_0542;
    89: op1_14_in26 = reg_0113;
    90: op1_14_in26 = reg_0588;
    91: op1_14_in26 = reg_0007;
    92: op1_14_in26 = reg_0181;
    95: op1_14_in26 = reg_0641;
    96: op1_14_in26 = reg_0361;
    default: op1_14_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv26 = 1;
    6: op1_14_inv26 = 1;
    8: op1_14_inv26 = 1;
    10: op1_14_inv26 = 1;
    11: op1_14_inv26 = 1;
    12: op1_14_inv26 = 1;
    13: op1_14_inv26 = 1;
    17: op1_14_inv26 = 1;
    18: op1_14_inv26 = 1;
    19: op1_14_inv26 = 1;
    20: op1_14_inv26 = 1;
    21: op1_14_inv26 = 1;
    23: op1_14_inv26 = 1;
    24: op1_14_inv26 = 1;
    25: op1_14_inv26 = 1;
    26: op1_14_inv26 = 1;
    27: op1_14_inv26 = 1;
    29: op1_14_inv26 = 1;
    30: op1_14_inv26 = 1;
    31: op1_14_inv26 = 1;
    32: op1_14_inv26 = 1;
    33: op1_14_inv26 = 1;
    37: op1_14_inv26 = 1;
    41: op1_14_inv26 = 1;
    46: op1_14_inv26 = 1;
    49: op1_14_inv26 = 1;
    50: op1_14_inv26 = 1;
    54: op1_14_inv26 = 1;
    56: op1_14_inv26 = 1;
    58: op1_14_inv26 = 1;
    60: op1_14_inv26 = 1;
    65: op1_14_inv26 = 1;
    68: op1_14_inv26 = 1;
    69: op1_14_inv26 = 1;
    70: op1_14_inv26 = 1;
    73: op1_14_inv26 = 1;
    74: op1_14_inv26 = 1;
    75: op1_14_inv26 = 1;
    77: op1_14_inv26 = 1;
    78: op1_14_inv26 = 1;
    81: op1_14_inv26 = 1;
    82: op1_14_inv26 = 1;
    85: op1_14_inv26 = 1;
    88: op1_14_inv26 = 1;
    89: op1_14_inv26 = 1;
    90: op1_14_inv26 = 1;
    92: op1_14_inv26 = 1;
    96: op1_14_inv26 = 1;
    default: op1_14_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in27 = reg_0112;
    6: op1_14_in27 = imem07_in[63:60];
    7: op1_14_in27 = imem03_in[23:20];
    8: op1_14_in27 = reg_0296;
    70: op1_14_in27 = reg_0296;
    9: op1_14_in27 = reg_0200;
    10: op1_14_in27 = reg_0715;
    11: op1_14_in27 = imem04_in[99:96];
    73: op1_14_in27 = imem04_in[99:96];
    12: op1_14_in27 = imem05_in[47:44];
    13: op1_14_in27 = reg_0360;
    14: op1_14_in27 = imem05_in[43:40];
    85: op1_14_in27 = imem05_in[43:40];
    15: op1_14_in27 = reg_0332;
    88: op1_14_in27 = reg_0332;
    16: op1_14_in27 = imem01_in[119:116];
    17: op1_14_in27 = reg_0585;
    18: op1_14_in27 = imem02_in[67:64];
    19: op1_14_in27 = imem03_in[27:24];
    20: op1_14_in27 = imem01_in[27:24];
    21: op1_14_in27 = reg_0549;
    22: op1_14_in27 = reg_0622;
    23: op1_14_in27 = imem02_in[19:16];
    89: op1_14_in27 = imem02_in[19:16];
    24: op1_14_in27 = reg_0180;
    25: op1_14_in27 = reg_0304;
    69: op1_14_in27 = reg_0304;
    26: op1_14_in27 = reg_0129;
    27: op1_14_in27 = reg_0916;
    28: op1_14_in27 = imem03_in[123:120];
    48: op1_14_in27 = imem03_in[123:120];
    29: op1_14_in27 = imem07_in[19:16];
    43: op1_14_in27 = imem07_in[19:16];
    30: op1_14_in27 = reg_0230;
    31: op1_14_in27 = reg_0751;
    32: op1_14_in27 = reg_0145;
    33: op1_14_in27 = reg_0222;
    34: op1_14_in27 = reg_0988;
    35: op1_14_in27 = reg_1020;
    36: op1_14_in27 = reg_0054;
    37: op1_14_in27 = imem07_in[103:100];
    38: op1_14_in27 = reg_0293;
    41: op1_14_in27 = imem02_in[71:68];
    42: op1_14_in27 = reg_0950;
    45: op1_14_in27 = imem03_in[103:100];
    46: op1_14_in27 = imem06_in[47:44];
    49: op1_14_in27 = reg_1009;
    50: op1_14_in27 = reg_0083;
    51: op1_14_in27 = reg_0762;
    53: op1_14_in27 = reg_1031;
    54: op1_14_in27 = imem01_in[127:124];
    55: op1_14_in27 = imem03_in[115:112];
    56: op1_14_in27 = reg_0015;
    57: op1_14_in27 = reg_0578;
    58: op1_14_in27 = imem03_in[71:68];
    59: op1_14_in27 = reg_0591;
    60: op1_14_in27 = reg_0537;
    61: op1_14_in27 = reg_1030;
    63: op1_14_in27 = reg_0840;
    64: op1_14_in27 = imem03_in[127:124];
    65: op1_14_in27 = reg_0006;
    66: op1_14_in27 = reg_0277;
    67: op1_14_in27 = reg_0844;
    68: op1_14_in27 = reg_0176;
    72: op1_14_in27 = reg_0580;
    74: op1_14_in27 = reg_0275;
    75: op1_14_in27 = imem06_in[115:112];
    76: op1_14_in27 = reg_0250;
    77: op1_14_in27 = reg_1044;
    78: op1_14_in27 = reg_0327;
    79: op1_14_in27 = reg_0327;
    80: op1_14_in27 = reg_0651;
    81: op1_14_in27 = reg_0780;
    82: op1_14_in27 = imem03_in[55:52];
    83: op1_14_in27 = imem01_in[95:92];
    86: op1_14_in27 = reg_0390;
    87: op1_14_in27 = reg_0737;
    90: op1_14_in27 = reg_0266;
    91: op1_14_in27 = reg_0331;
    92: op1_14_in27 = reg_0179;
    95: op1_14_in27 = reg_0431;
    96: op1_14_in27 = reg_0303;
    default: op1_14_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv27 = 1;
    6: op1_14_inv27 = 1;
    7: op1_14_inv27 = 1;
    9: op1_14_inv27 = 1;
    11: op1_14_inv27 = 1;
    12: op1_14_inv27 = 1;
    14: op1_14_inv27 = 1;
    16: op1_14_inv27 = 1;
    17: op1_14_inv27 = 1;
    19: op1_14_inv27 = 1;
    21: op1_14_inv27 = 1;
    22: op1_14_inv27 = 1;
    23: op1_14_inv27 = 1;
    24: op1_14_inv27 = 1;
    28: op1_14_inv27 = 1;
    29: op1_14_inv27 = 1;
    31: op1_14_inv27 = 1;
    32: op1_14_inv27 = 1;
    33: op1_14_inv27 = 1;
    34: op1_14_inv27 = 1;
    37: op1_14_inv27 = 1;
    43: op1_14_inv27 = 1;
    45: op1_14_inv27 = 1;
    50: op1_14_inv27 = 1;
    53: op1_14_inv27 = 1;
    55: op1_14_inv27 = 1;
    57: op1_14_inv27 = 1;
    59: op1_14_inv27 = 1;
    60: op1_14_inv27 = 1;
    61: op1_14_inv27 = 1;
    64: op1_14_inv27 = 1;
    65: op1_14_inv27 = 1;
    67: op1_14_inv27 = 1;
    68: op1_14_inv27 = 1;
    69: op1_14_inv27 = 1;
    70: op1_14_inv27 = 1;
    72: op1_14_inv27 = 1;
    73: op1_14_inv27 = 1;
    77: op1_14_inv27 = 1;
    78: op1_14_inv27 = 1;
    82: op1_14_inv27 = 1;
    83: op1_14_inv27 = 1;
    85: op1_14_inv27 = 1;
    86: op1_14_inv27 = 1;
    90: op1_14_inv27 = 1;
    91: op1_14_inv27 = 1;
    92: op1_14_inv27 = 1;
    96: op1_14_inv27 = 1;
    default: op1_14_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in28 = reg_0113;
    6: op1_14_in28 = imem07_in[79:76];
    7: op1_14_in28 = imem03_in[35:32];
    8: op1_14_in28 = reg_0297;
    9: op1_14_in28 = reg_0208;
    10: op1_14_in28 = reg_0701;
    11: op1_14_in28 = reg_0543;
    12: op1_14_in28 = imem05_in[59:56];
    13: op1_14_in28 = reg_0319;
    14: op1_14_in28 = imem05_in[119:116];
    15: op1_14_in28 = reg_0344;
    16: op1_14_in28 = reg_0249;
    17: op1_14_in28 = reg_0578;
    18: op1_14_in28 = imem02_in[91:88];
    19: op1_14_in28 = imem03_in[63:60];
    20: op1_14_in28 = imem01_in[55:52];
    21: op1_14_in28 = reg_0554;
    22: op1_14_in28 = reg_0407;
    23: op1_14_in28 = imem02_in[23:20];
    24: op1_14_in28 = reg_0165;
    25: op1_14_in28 = reg_0906;
    69: op1_14_in28 = reg_0906;
    26: op1_14_in28 = imem06_in[15:12];
    27: op1_14_in28 = reg_0096;
    28: op1_14_in28 = reg_0987;
    29: op1_14_in28 = imem07_in[27:24];
    30: op1_14_in28 = reg_1043;
    31: op1_14_in28 = reg_0043;
    32: op1_14_in28 = reg_0135;
    33: op1_14_in28 = reg_0380;
    34: op1_14_in28 = reg_0983;
    35: op1_14_in28 = reg_1016;
    36: op1_14_in28 = reg_0738;
    37: op1_14_in28 = imem07_in[107:104];
    38: op1_14_in28 = reg_0356;
    41: op1_14_in28 = imem02_in[95:92];
    42: op1_14_in28 = reg_0972;
    43: op1_14_in28 = imem07_in[35:32];
    45: op1_14_in28 = reg_0535;
    46: op1_14_in28 = imem06_in[79:76];
    48: op1_14_in28 = reg_0492;
    49: op1_14_in28 = reg_0277;
    50: op1_14_in28 = reg_0007;
    51: op1_14_in28 = reg_0870;
    53: op1_14_in28 = reg_0521;
    54: op1_14_in28 = reg_0918;
    55: op1_14_in28 = reg_0765;
    56: op1_14_in28 = reg_0064;
    57: op1_14_in28 = reg_0075;
    58: op1_14_in28 = reg_0006;
    59: op1_14_in28 = reg_0894;
    60: op1_14_in28 = reg_0752;
    61: op1_14_in28 = reg_0804;
    63: op1_14_in28 = reg_0016;
    64: op1_14_in28 = reg_0620;
    65: op1_14_in28 = reg_0620;
    66: op1_14_in28 = reg_0282;
    67: op1_14_in28 = reg_0374;
    70: op1_14_in28 = reg_0808;
    72: op1_14_in28 = reg_0322;
    73: op1_14_in28 = imem04_in[119:116];
    74: op1_14_in28 = reg_0235;
    75: op1_14_in28 = reg_0338;
    76: op1_14_in28 = reg_0325;
    77: op1_14_in28 = reg_0971;
    78: op1_14_in28 = reg_0585;
    79: op1_14_in28 = reg_0046;
    80: op1_14_in28 = reg_0508;
    81: op1_14_in28 = reg_0970;
    82: op1_14_in28 = imem03_in[59:56];
    83: op1_14_in28 = imem01_in[99:96];
    85: op1_14_in28 = imem05_in[67:64];
    86: op1_14_in28 = reg_0586;
    87: op1_14_in28 = reg_0354;
    88: op1_14_in28 = imem05_in[7:4];
    89: op1_14_in28 = imem02_in[31:28];
    90: op1_14_in28 = imem03_in[23:20];
    91: op1_14_in28 = reg_0820;
    92: op1_14_in28 = reg_0184;
    95: op1_14_in28 = reg_0182;
    96: op1_14_in28 = reg_0315;
    default: op1_14_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv28 = 1;
    7: op1_14_inv28 = 1;
    8: op1_14_inv28 = 1;
    13: op1_14_inv28 = 1;
    14: op1_14_inv28 = 1;
    17: op1_14_inv28 = 1;
    20: op1_14_inv28 = 1;
    21: op1_14_inv28 = 1;
    22: op1_14_inv28 = 1;
    23: op1_14_inv28 = 1;
    24: op1_14_inv28 = 1;
    26: op1_14_inv28 = 1;
    29: op1_14_inv28 = 1;
    30: op1_14_inv28 = 1;
    33: op1_14_inv28 = 1;
    35: op1_14_inv28 = 1;
    41: op1_14_inv28 = 1;
    45: op1_14_inv28 = 1;
    51: op1_14_inv28 = 1;
    53: op1_14_inv28 = 1;
    54: op1_14_inv28 = 1;
    55: op1_14_inv28 = 1;
    56: op1_14_inv28 = 1;
    59: op1_14_inv28 = 1;
    60: op1_14_inv28 = 1;
    61: op1_14_inv28 = 1;
    64: op1_14_inv28 = 1;
    65: op1_14_inv28 = 1;
    66: op1_14_inv28 = 1;
    67: op1_14_inv28 = 1;
    70: op1_14_inv28 = 1;
    72: op1_14_inv28 = 1;
    74: op1_14_inv28 = 1;
    75: op1_14_inv28 = 1;
    76: op1_14_inv28 = 1;
    78: op1_14_inv28 = 1;
    81: op1_14_inv28 = 1;
    82: op1_14_inv28 = 1;
    86: op1_14_inv28 = 1;
    87: op1_14_inv28 = 1;
    88: op1_14_inv28 = 1;
    89: op1_14_inv28 = 1;
    92: op1_14_inv28 = 1;
    95: op1_14_inv28 = 1;
    default: op1_14_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in29 = reg_0121;
    6: op1_14_in29 = imem07_in[91:88];
    7: op1_14_in29 = imem03_in[47:44];
    8: op1_14_in29 = reg_0275;
    9: op1_14_in29 = reg_0191;
    10: op1_14_in29 = reg_0430;
    11: op1_14_in29 = reg_0552;
    12: op1_14_in29 = imem05_in[107:104];
    13: op1_14_in29 = reg_0385;
    14: op1_14_in29 = reg_0959;
    15: op1_14_in29 = reg_0372;
    16: op1_14_in29 = reg_0216;
    30: op1_14_in29 = reg_0216;
    17: op1_14_in29 = reg_0576;
    18: op1_14_in29 = imem02_in[99:96];
    19: op1_14_in29 = imem03_in[79:76];
    20: op1_14_in29 = imem01_in[59:56];
    21: op1_14_in29 = reg_0556;
    22: op1_14_in29 = reg_0409;
    23: op1_14_in29 = reg_0653;
    24: op1_14_in29 = reg_0162;
    25: op1_14_in29 = imem01_in[15:12];
    26: op1_14_in29 = imem06_in[83:80];
    27: op1_14_in29 = reg_0865;
    28: op1_14_in29 = reg_1002;
    29: op1_14_in29 = imem07_in[31:28];
    31: op1_14_in29 = reg_0854;
    32: op1_14_in29 = reg_0143;
    33: op1_14_in29 = reg_0402;
    34: op1_14_in29 = imem04_in[15:12];
    35: op1_14_in29 = reg_0313;
    36: op1_14_in29 = reg_0021;
    37: op1_14_in29 = imem07_in[115:112];
    38: op1_14_in29 = reg_0332;
    41: op1_14_in29 = reg_0640;
    42: op1_14_in29 = reg_0229;
    43: op1_14_in29 = imem07_in[47:44];
    45: op1_14_in29 = reg_1049;
    46: op1_14_in29 = imem06_in[115:112];
    48: op1_14_in29 = reg_1050;
    49: op1_14_in29 = reg_0055;
    50: op1_14_in29 = reg_0761;
    51: op1_14_in29 = reg_0919;
    53: op1_14_in29 = reg_0304;
    54: op1_14_in29 = reg_0762;
    55: op1_14_in29 = reg_0370;
    56: op1_14_in29 = reg_0809;
    57: op1_14_in29 = imem05_in[35:32];
    58: op1_14_in29 = reg_0620;
    59: op1_14_in29 = reg_0241;
    60: op1_14_in29 = reg_0015;
    61: op1_14_in29 = reg_0632;
    63: op1_14_in29 = reg_0077;
    64: op1_14_in29 = reg_0535;
    65: op1_14_in29 = reg_0760;
    66: op1_14_in29 = reg_0912;
    67: op1_14_in29 = reg_0822;
    69: op1_14_in29 = reg_0114;
    70: op1_14_in29 = reg_0815;
    72: op1_14_in29 = reg_0238;
    73: op1_14_in29 = reg_1004;
    74: op1_14_in29 = reg_0057;
    75: op1_14_in29 = reg_0624;
    76: op1_14_in29 = reg_0321;
    77: op1_14_in29 = reg_1022;
    78: op1_14_in29 = reg_0298;
    79: op1_14_in29 = reg_0547;
    80: op1_14_in29 = reg_0949;
    81: op1_14_in29 = reg_0508;
    82: op1_14_in29 = imem03_in[75:72];
    83: op1_14_in29 = reg_1042;
    85: op1_14_in29 = imem05_in[79:76];
    86: op1_14_in29 = reg_0123;
    87: op1_14_in29 = reg_0610;
    88: op1_14_in29 = imem05_in[55:52];
    89: op1_14_in29 = imem02_in[43:40];
    90: op1_14_in29 = imem03_in[31:28];
    91: op1_14_in29 = reg_0233;
    95: op1_14_in29 = reg_0449;
    96: op1_14_in29 = reg_0428;
    default: op1_14_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_14_inv29 = 1;
    8: op1_14_inv29 = 1;
    9: op1_14_inv29 = 1;
    14: op1_14_inv29 = 1;
    17: op1_14_inv29 = 1;
    18: op1_14_inv29 = 1;
    19: op1_14_inv29 = 1;
    23: op1_14_inv29 = 1;
    27: op1_14_inv29 = 1;
    29: op1_14_inv29 = 1;
    31: op1_14_inv29 = 1;
    33: op1_14_inv29 = 1;
    42: op1_14_inv29 = 1;
    46: op1_14_inv29 = 1;
    50: op1_14_inv29 = 1;
    51: op1_14_inv29 = 1;
    53: op1_14_inv29 = 1;
    54: op1_14_inv29 = 1;
    56: op1_14_inv29 = 1;
    58: op1_14_inv29 = 1;
    60: op1_14_inv29 = 1;
    61: op1_14_inv29 = 1;
    66: op1_14_inv29 = 1;
    69: op1_14_inv29 = 1;
    72: op1_14_inv29 = 1;
    73: op1_14_inv29 = 1;
    74: op1_14_inv29 = 1;
    75: op1_14_inv29 = 1;
    76: op1_14_inv29 = 1;
    77: op1_14_inv29 = 1;
    78: op1_14_inv29 = 1;
    79: op1_14_inv29 = 1;
    80: op1_14_inv29 = 1;
    81: op1_14_inv29 = 1;
    85: op1_14_inv29 = 1;
    86: op1_14_inv29 = 1;
    87: op1_14_inv29 = 1;
    89: op1_14_inv29 = 1;
    90: op1_14_inv29 = 1;
    default: op1_14_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_14_in30 = imem02_in[23:20];
    6: op1_14_in30 = imem07_in[107:104];
    7: op1_14_in30 = imem03_in[51:48];
    8: op1_14_in30 = reg_0278;
    9: op1_14_in30 = reg_0187;
    10: op1_14_in30 = reg_0432;
    60: op1_14_in30 = reg_0432;
    11: op1_14_in30 = reg_0548;
    12: op1_14_in30 = reg_0132;
    13: op1_14_in30 = reg_0398;
    45: op1_14_in30 = reg_0398;
    14: op1_14_in30 = reg_0955;
    15: op1_14_in30 = reg_0408;
    16: op1_14_in30 = reg_1040;
    17: op1_14_in30 = reg_0319;
    18: op1_14_in30 = imem02_in[127:124];
    19: op1_14_in30 = imem03_in[99:96];
    20: op1_14_in30 = imem01_in[83:80];
    21: op1_14_in30 = reg_0547;
    22: op1_14_in30 = reg_0399;
    23: op1_14_in30 = reg_0661;
    24: op1_14_in30 = reg_0159;
    25: op1_14_in30 = imem01_in[19:16];
    26: op1_14_in30 = imem06_in[115:112];
    27: op1_14_in30 = reg_0338;
    28: op1_14_in30 = reg_0995;
    29: op1_14_in30 = imem07_in[47:44];
    30: op1_14_in30 = reg_0871;
    31: op1_14_in30 = imem05_in[11:8];
    36: op1_14_in30 = imem05_in[11:8];
    32: op1_14_in30 = reg_0153;
    33: op1_14_in30 = reg_0599;
    34: op1_14_in30 = imem04_in[27:24];
    35: op1_14_in30 = reg_0760;
    37: op1_14_in30 = reg_0722;
    38: op1_14_in30 = reg_0626;
    41: op1_14_in30 = reg_0641;
    42: op1_14_in30 = reg_0275;
    43: op1_14_in30 = reg_0162;
    46: op1_14_in30 = reg_0073;
    48: op1_14_in30 = reg_0317;
    49: op1_14_in30 = reg_1057;
    50: op1_14_in30 = reg_0792;
    51: op1_14_in30 = reg_0592;
    53: op1_14_in30 = imem01_in[15:12];
    54: op1_14_in30 = reg_0933;
    55: op1_14_in30 = reg_1002;
    56: op1_14_in30 = reg_0284;
    57: op1_14_in30 = imem05_in[39:36];
    58: op1_14_in30 = reg_0345;
    59: op1_14_in30 = reg_0605;
    61: op1_14_in30 = reg_0917;
    63: op1_14_in30 = reg_0079;
    64: op1_14_in30 = reg_1007;
    65: op1_14_in30 = reg_1007;
    66: op1_14_in30 = reg_1020;
    67: op1_14_in30 = reg_0985;
    69: op1_14_in30 = reg_0113;
    70: op1_14_in30 = reg_0288;
    72: op1_14_in30 = reg_0376;
    73: op1_14_in30 = reg_0282;
    74: op1_14_in30 = reg_0941;
    75: op1_14_in30 = reg_0533;
    76: op1_14_in30 = reg_0428;
    77: op1_14_in30 = reg_0862;
    78: op1_14_in30 = reg_0240;
    79: op1_14_in30 = reg_0823;
    80: op1_14_in30 = reg_0490;
    81: op1_14_in30 = imem06_in[27:24];
    82: op1_14_in30 = imem03_in[79:76];
    83: op1_14_in30 = reg_1014;
    85: op1_14_in30 = imem05_in[83:80];
    86: op1_14_in30 = reg_0524;
    87: op1_14_in30 = reg_0740;
    88: op1_14_in30 = imem05_in[99:96];
    89: op1_14_in30 = imem02_in[47:44];
    90: op1_14_in30 = imem03_in[87:84];
    91: op1_14_in30 = reg_0978;
    95: op1_14_in30 = reg_0697;
    96: op1_14_in30 = reg_0350;
    default: op1_14_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv30 = 1;
    7: op1_14_inv30 = 1;
    8: op1_14_inv30 = 1;
    9: op1_14_inv30 = 1;
    10: op1_14_inv30 = 1;
    11: op1_14_inv30 = 1;
    12: op1_14_inv30 = 1;
    16: op1_14_inv30 = 1;
    19: op1_14_inv30 = 1;
    20: op1_14_inv30 = 1;
    22: op1_14_inv30 = 1;
    24: op1_14_inv30 = 1;
    28: op1_14_inv30 = 1;
    29: op1_14_inv30 = 1;
    37: op1_14_inv30 = 1;
    38: op1_14_inv30 = 1;
    42: op1_14_inv30 = 1;
    45: op1_14_inv30 = 1;
    49: op1_14_inv30 = 1;
    53: op1_14_inv30 = 1;
    55: op1_14_inv30 = 1;
    57: op1_14_inv30 = 1;
    59: op1_14_inv30 = 1;
    63: op1_14_inv30 = 1;
    65: op1_14_inv30 = 1;
    67: op1_14_inv30 = 1;
    70: op1_14_inv30 = 1;
    72: op1_14_inv30 = 1;
    75: op1_14_inv30 = 1;
    77: op1_14_inv30 = 1;
    78: op1_14_inv30 = 1;
    79: op1_14_inv30 = 1;
    82: op1_14_inv30 = 1;
    83: op1_14_inv30 = 1;
    85: op1_14_inv30 = 1;
    86: op1_14_inv30 = 1;
    89: op1_14_inv30 = 1;
    90: op1_14_inv30 = 1;
    91: op1_14_inv30 = 1;
    95: op1_14_inv30 = 1;
    96: op1_14_inv30 = 1;
    default: op1_14_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_14_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_14_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in00 = imem02_in[31:28];
    6: op1_15_in00 = imem07_in[123:120];
    7: op1_15_in00 = imem03_in[75:72];
    8: op1_15_in00 = reg_0046;
    9: op1_15_in00 = reg_0188;
    10: op1_15_in00 = imem00_in[35:32];
    52: op1_15_in00 = imem00_in[35:32];
    11: op1_15_in00 = reg_0541;
    12: op1_15_in00 = reg_0148;
    13: op1_15_in00 = reg_0389;
    14: op1_15_in00 = reg_0217;
    15: op1_15_in00 = reg_0403;
    16: op1_15_in00 = reg_1031;
    17: op1_15_in00 = reg_0327;
    18: op1_15_in00 = reg_0666;
    89: op1_15_in00 = reg_0666;
    19: op1_15_in00 = reg_0578;
    20: op1_15_in00 = imem01_in[99:96];
    21: op1_15_in00 = reg_0065;
    22: op1_15_in00 = reg_0367;
    23: op1_15_in00 = reg_0640;
    24: op1_15_in00 = imem00_in[51:48];
    25: op1_15_in00 = imem01_in[39:36];
    26: op1_15_in00 = reg_0610;
    27: op1_15_in00 = reg_0762;
    28: op1_15_in00 = reg_0993;
    29: op1_15_in00 = imem07_in[119:116];
    4: op1_15_in00 = imem07_in[47:44];
    30: op1_15_in00 = reg_0123;
    31: op1_15_in00 = imem05_in[27:24];
    32: op1_15_in00 = reg_0130;
    33: op1_15_in00 = reg_0026;
    2: op1_15_in00 = imem07_in[99:96];
    34: op1_15_in00 = imem04_in[35:32];
    3: op1_15_in00 = reg_0170;
    35: op1_15_in00 = reg_0268;
    36: op1_15_in00 = imem05_in[23:20];
    37: op1_15_in00 = reg_0723;
    38: op1_15_in00 = reg_1010;
    39: op1_15_in00 = imem00_in[67:64];
    40: op1_15_in00 = imem00_in[23:20];
    92: op1_15_in00 = imem00_in[23:20];
    41: op1_15_in00 = reg_0665;
    42: op1_15_in00 = reg_0155;
    43: op1_15_in00 = reg_0169;
    44: op1_15_in00 = imem00_in[3:0];
    68: op1_15_in00 = imem00_in[3:0];
    93: op1_15_in00 = imem00_in[3:0];
    45: op1_15_in00 = reg_0346;
    46: op1_15_in00 = reg_0759;
    47: op1_15_in00 = imem00_in[7:4];
    62: op1_15_in00 = imem00_in[7:4];
    48: op1_15_in00 = reg_0343;
    49: op1_15_in00 = reg_1020;
    50: op1_15_in00 = reg_0086;
    51: op1_15_in00 = reg_1035;
    53: op1_15_in00 = imem01_in[55:52];
    54: op1_15_in00 = reg_0503;
    55: op1_15_in00 = reg_0979;
    56: op1_15_in00 = reg_0756;
    57: op1_15_in00 = imem05_in[71:68];
    58: op1_15_in00 = reg_0099;
    59: op1_15_in00 = reg_0017;
    60: op1_15_in00 = imem05_in[11:8];
    61: op1_15_in00 = imem06_in[27:24];
    63: op1_15_in00 = imem03_in[3:0];
    64: op1_15_in00 = reg_0245;
    65: op1_15_in00 = reg_0240;
    66: op1_15_in00 = reg_0050;
    67: op1_15_in00 = reg_0996;
    69: op1_15_in00 = reg_0821;
    70: op1_15_in00 = reg_0732;
    71: op1_15_in00 = imem00_in[43:40];
    72: op1_15_in00 = reg_0385;
    73: op1_15_in00 = reg_0888;
    74: op1_15_in00 = reg_0675;
    75: op1_15_in00 = reg_0439;
    76: op1_15_in00 = reg_0353;
    77: op1_15_in00 = reg_0607;
    78: op1_15_in00 = reg_0661;
    79: op1_15_in00 = reg_0278;
    80: op1_15_in00 = imem06_in[11:8];
    81: op1_15_in00 = imem06_in[47:44];
    82: op1_15_in00 = imem03_in[83:80];
    83: op1_15_in00 = reg_0546;
    84: op1_15_in00 = imem00_in[31:28];
    85: op1_15_in00 = imem05_in[127:124];
    86: op1_15_in00 = reg_0067;
    87: op1_15_in00 = reg_0615;
    88: op1_15_in00 = reg_0866;
    90: op1_15_in00 = imem03_in[111:108];
    91: op1_15_in00 = reg_0509;
    94: op1_15_in00 = imem00_in[15:12];
    95: op1_15_in00 = reg_0171;
    96: op1_15_in00 = reg_0868;
    default: op1_15_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv00 = 1;
    8: op1_15_inv00 = 1;
    11: op1_15_inv00 = 1;
    17: op1_15_inv00 = 1;
    19: op1_15_inv00 = 1;
    21: op1_15_inv00 = 1;
    22: op1_15_inv00 = 1;
    24: op1_15_inv00 = 1;
    25: op1_15_inv00 = 1;
    26: op1_15_inv00 = 1;
    29: op1_15_inv00 = 1;
    4: op1_15_inv00 = 1;
    32: op1_15_inv00 = 1;
    2: op1_15_inv00 = 1;
    34: op1_15_inv00 = 1;
    36: op1_15_inv00 = 1;
    39: op1_15_inv00 = 1;
    41: op1_15_inv00 = 1;
    44: op1_15_inv00 = 1;
    45: op1_15_inv00 = 1;
    46: op1_15_inv00 = 1;
    47: op1_15_inv00 = 1;
    48: op1_15_inv00 = 1;
    49: op1_15_inv00 = 1;
    51: op1_15_inv00 = 1;
    53: op1_15_inv00 = 1;
    54: op1_15_inv00 = 1;
    55: op1_15_inv00 = 1;
    57: op1_15_inv00 = 1;
    58: op1_15_inv00 = 1;
    59: op1_15_inv00 = 1;
    61: op1_15_inv00 = 1;
    63: op1_15_inv00 = 1;
    66: op1_15_inv00 = 1;
    68: op1_15_inv00 = 1;
    70: op1_15_inv00 = 1;
    71: op1_15_inv00 = 1;
    73: op1_15_inv00 = 1;
    75: op1_15_inv00 = 1;
    78: op1_15_inv00 = 1;
    79: op1_15_inv00 = 1;
    80: op1_15_inv00 = 1;
    81: op1_15_inv00 = 1;
    83: op1_15_inv00 = 1;
    84: op1_15_inv00 = 1;
    85: op1_15_inv00 = 1;
    86: op1_15_inv00 = 1;
    87: op1_15_inv00 = 1;
    88: op1_15_inv00 = 1;
    91: op1_15_inv00 = 1;
    92: op1_15_inv00 = 1;
    94: op1_15_inv00 = 1;
    95: op1_15_inv00 = 1;
    default: op1_15_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in01 = imem02_in[43:40];
    6: op1_15_in01 = reg_0704;
    7: op1_15_in01 = imem03_in[87:84];
    8: op1_15_in01 = imem05_in[3:0];
    9: op1_15_in01 = reg_0203;
    10: op1_15_in01 = imem00_in[47:44];
    52: op1_15_in01 = imem00_in[47:44];
    11: op1_15_in01 = reg_0547;
    12: op1_15_in01 = reg_0136;
    13: op1_15_in01 = reg_0998;
    14: op1_15_in01 = reg_0250;
    15: op1_15_in01 = reg_0390;
    16: op1_15_in01 = reg_1038;
    17: op1_15_in01 = reg_0377;
    18: op1_15_in01 = reg_0664;
    19: op1_15_in01 = reg_0581;
    20: op1_15_in01 = imem01_in[127:124];
    21: op1_15_in01 = reg_0067;
    22: op1_15_in01 = reg_0401;
    23: op1_15_in01 = reg_0667;
    24: op1_15_in01 = imem00_in[83:80];
    25: op1_15_in01 = imem01_in[59:56];
    26: op1_15_in01 = reg_0625;
    27: op1_15_in01 = reg_0336;
    28: op1_15_in01 = imem04_in[31:28];
    29: op1_15_in01 = reg_0720;
    4: op1_15_in01 = imem07_in[51:48];
    30: op1_15_in01 = reg_0105;
    31: op1_15_in01 = imem05_in[67:64];
    32: op1_15_in01 = reg_0131;
    33: op1_15_in01 = reg_0753;
    34: op1_15_in01 = imem04_in[39:36];
    35: op1_15_in01 = reg_0069;
    36: op1_15_in01 = imem05_in[43:40];
    37: op1_15_in01 = reg_0703;
    38: op1_15_in01 = reg_0008;
    39: op1_15_in01 = imem00_in[71:68];
    40: op1_15_in01 = imem00_in[67:64];
    41: op1_15_in01 = reg_0837;
    42: op1_15_in01 = imem06_in[15:12];
    43: op1_15_in01 = reg_0163;
    44: op1_15_in01 = imem00_in[15:12];
    45: op1_15_in01 = reg_0874;
    46: op1_15_in01 = reg_0624;
    47: op1_15_in01 = imem00_in[23:20];
    48: op1_15_in01 = reg_0938;
    49: op1_15_in01 = reg_0050;
    50: op1_15_in01 = reg_0090;
    51: op1_15_in01 = reg_0503;
    53: op1_15_in01 = imem01_in[75:72];
    54: op1_15_in01 = reg_0607;
    55: op1_15_in01 = reg_0993;
    56: op1_15_in01 = reg_0864;
    57: op1_15_in01 = imem05_in[127:124];
    58: op1_15_in01 = reg_0445;
    59: op1_15_in01 = reg_0633;
    60: op1_15_in01 = imem05_in[31:28];
    61: op1_15_in01 = imem06_in[115:112];
    62: op1_15_in01 = imem00_in[51:48];
    71: op1_15_in01 = imem00_in[51:48];
    84: op1_15_in01 = imem00_in[51:48];
    92: op1_15_in01 = imem00_in[51:48];
    63: op1_15_in01 = imem03_in[11:8];
    64: op1_15_in01 = reg_0434;
    65: op1_15_in01 = reg_0576;
    66: op1_15_in01 = reg_0537;
    67: op1_15_in01 = reg_1001;
    68: op1_15_in01 = imem00_in[7:4];
    69: op1_15_in01 = imem02_in[35:32];
    70: op1_15_in01 = reg_0284;
    72: op1_15_in01 = reg_1002;
    73: op1_15_in01 = reg_1016;
    74: op1_15_in01 = reg_0125;
    75: op1_15_in01 = reg_0804;
    76: op1_15_in01 = reg_0589;
    77: op1_15_in01 = reg_0604;
    78: op1_15_in01 = reg_0662;
    79: op1_15_in01 = reg_0281;
    80: op1_15_in01 = imem06_in[35:32];
    81: op1_15_in01 = imem06_in[103:100];
    82: op1_15_in01 = imem03_in[107:104];
    83: op1_15_in01 = reg_0234;
    85: op1_15_in01 = reg_1021;
    86: op1_15_in01 = reg_0074;
    87: op1_15_in01 = reg_1055;
    88: op1_15_in01 = reg_0217;
    89: op1_15_in01 = reg_0605;
    90: op1_15_in01 = imem03_in[115:112];
    91: op1_15_in01 = imem04_in[47:44];
    93: op1_15_in01 = imem00_in[11:8];
    94: op1_15_in01 = imem00_in[63:60];
    96: op1_15_in01 = reg_0024;
    default: op1_15_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv01 = 1;
    9: op1_15_inv01 = 1;
    10: op1_15_inv01 = 1;
    11: op1_15_inv01 = 1;
    12: op1_15_inv01 = 1;
    13: op1_15_inv01 = 1;
    19: op1_15_inv01 = 1;
    20: op1_15_inv01 = 1;
    22: op1_15_inv01 = 1;
    23: op1_15_inv01 = 1;
    25: op1_15_inv01 = 1;
    28: op1_15_inv01 = 1;
    29: op1_15_inv01 = 1;
    4: op1_15_inv01 = 1;
    32: op1_15_inv01 = 1;
    33: op1_15_inv01 = 1;
    34: op1_15_inv01 = 1;
    35: op1_15_inv01 = 1;
    38: op1_15_inv01 = 1;
    40: op1_15_inv01 = 1;
    42: op1_15_inv01 = 1;
    43: op1_15_inv01 = 1;
    47: op1_15_inv01 = 1;
    48: op1_15_inv01 = 1;
    51: op1_15_inv01 = 1;
    53: op1_15_inv01 = 1;
    56: op1_15_inv01 = 1;
    58: op1_15_inv01 = 1;
    59: op1_15_inv01 = 1;
    61: op1_15_inv01 = 1;
    62: op1_15_inv01 = 1;
    63: op1_15_inv01 = 1;
    64: op1_15_inv01 = 1;
    65: op1_15_inv01 = 1;
    66: op1_15_inv01 = 1;
    68: op1_15_inv01 = 1;
    69: op1_15_inv01 = 1;
    73: op1_15_inv01 = 1;
    77: op1_15_inv01 = 1;
    78: op1_15_inv01 = 1;
    80: op1_15_inv01 = 1;
    81: op1_15_inv01 = 1;
    82: op1_15_inv01 = 1;
    85: op1_15_inv01 = 1;
    86: op1_15_inv01 = 1;
    87: op1_15_inv01 = 1;
    89: op1_15_inv01 = 1;
    92: op1_15_inv01 = 1;
    93: op1_15_inv01 = 1;
    94: op1_15_inv01 = 1;
    96: op1_15_inv01 = 1;
    default: op1_15_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in02 = imem02_in[51:48];
    6: op1_15_in02 = reg_0721;
    7: op1_15_in02 = imem03_in[95:92];
    8: op1_15_in02 = imem05_in[47:44];
    9: op1_15_in02 = reg_0196;
    10: op1_15_in02 = imem00_in[51:48];
    11: op1_15_in02 = reg_0282;
    12: op1_15_in02 = reg_0151;
    13: op1_15_in02 = reg_1002;
    14: op1_15_in02 = reg_0258;
    15: op1_15_in02 = reg_0367;
    16: op1_15_in02 = reg_1034;
    51: op1_15_in02 = reg_1034;
    17: op1_15_in02 = reg_0393;
    18: op1_15_in02 = reg_0656;
    19: op1_15_in02 = reg_0588;
    20: op1_15_in02 = reg_1055;
    21: op1_15_in02 = reg_0072;
    22: op1_15_in02 = reg_0027;
    23: op1_15_in02 = reg_0663;
    24: op1_15_in02 = imem00_in[99:96];
    25: op1_15_in02 = imem01_in[87:84];
    26: op1_15_in02 = reg_0604;
    27: op1_15_in02 = reg_0083;
    28: op1_15_in02 = imem04_in[35:32];
    29: op1_15_in02 = reg_0730;
    4: op1_15_in02 = imem07_in[91:88];
    30: op1_15_in02 = reg_0124;
    31: op1_15_in02 = imem05_in[87:84];
    32: op1_15_in02 = reg_0144;
    33: op1_15_in02 = reg_0030;
    34: op1_15_in02 = imem04_in[127:124];
    35: op1_15_in02 = reg_0058;
    36: op1_15_in02 = imem05_in[71:68];
    37: op1_15_in02 = reg_0440;
    38: op1_15_in02 = imem07_in[27:24];
    39: op1_15_in02 = imem00_in[107:104];
    52: op1_15_in02 = imem00_in[107:104];
    40: op1_15_in02 = imem00_in[71:68];
    41: op1_15_in02 = reg_0818;
    42: op1_15_in02 = imem06_in[23:20];
    43: op1_15_in02 = reg_0183;
    44: op1_15_in02 = imem00_in[91:88];
    45: op1_15_in02 = reg_0543;
    46: op1_15_in02 = reg_0577;
    47: op1_15_in02 = imem00_in[75:72];
    48: op1_15_in02 = reg_1049;
    49: op1_15_in02 = reg_0802;
    50: op1_15_in02 = reg_0506;
    53: op1_15_in02 = imem01_in[83:80];
    54: op1_15_in02 = reg_0869;
    55: op1_15_in02 = reg_1000;
    56: op1_15_in02 = imem05_in[3:0];
    57: op1_15_in02 = reg_0569;
    58: op1_15_in02 = reg_0547;
    59: op1_15_in02 = reg_0029;
    60: op1_15_in02 = imem05_in[55:52];
    61: op1_15_in02 = imem07_in[79:76];
    62: op1_15_in02 = imem00_in[67:64];
    63: op1_15_in02 = imem03_in[15:12];
    64: op1_15_in02 = reg_0346;
    65: op1_15_in02 = reg_0509;
    66: op1_15_in02 = reg_0507;
    67: op1_15_in02 = reg_0983;
    68: op1_15_in02 = imem00_in[35:32];
    69: op1_15_in02 = imem02_in[59:56];
    70: op1_15_in02 = reg_0777;
    71: op1_15_in02 = imem00_in[103:100];
    72: op1_15_in02 = reg_0992;
    73: op1_15_in02 = reg_0541;
    74: op1_15_in02 = reg_0004;
    75: op1_15_in02 = reg_0695;
    76: op1_15_in02 = reg_0640;
    77: op1_15_in02 = reg_1043;
    78: op1_15_in02 = reg_0238;
    79: op1_15_in02 = reg_0239;
    80: op1_15_in02 = imem06_in[43:40];
    81: op1_15_in02 = reg_0626;
    82: op1_15_in02 = reg_0345;
    83: op1_15_in02 = reg_0225;
    84: op1_15_in02 = reg_0684;
    85: op1_15_in02 = reg_0215;
    86: op1_15_in02 = reg_0288;
    87: op1_15_in02 = reg_0273;
    88: op1_15_in02 = reg_0652;
    89: op1_15_in02 = reg_0069;
    90: op1_15_in02 = imem04_in[3:0];
    91: op1_15_in02 = imem04_in[55:52];
    92: op1_15_in02 = imem00_in[115:112];
    93: op1_15_in02 = imem00_in[27:24];
    94: op1_15_in02 = reg_0682;
    96: op1_15_in02 = reg_0431;
    default: op1_15_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv02 = 1;
    6: op1_15_inv02 = 1;
    8: op1_15_inv02 = 1;
    10: op1_15_inv02 = 1;
    11: op1_15_inv02 = 1;
    14: op1_15_inv02 = 1;
    19: op1_15_inv02 = 1;
    20: op1_15_inv02 = 1;
    21: op1_15_inv02 = 1;
    23: op1_15_inv02 = 1;
    24: op1_15_inv02 = 1;
    26: op1_15_inv02 = 1;
    28: op1_15_inv02 = 1;
    4: op1_15_inv02 = 1;
    30: op1_15_inv02 = 1;
    36: op1_15_inv02 = 1;
    38: op1_15_inv02 = 1;
    39: op1_15_inv02 = 1;
    40: op1_15_inv02 = 1;
    43: op1_15_inv02 = 1;
    45: op1_15_inv02 = 1;
    46: op1_15_inv02 = 1;
    48: op1_15_inv02 = 1;
    49: op1_15_inv02 = 1;
    51: op1_15_inv02 = 1;
    53: op1_15_inv02 = 1;
    54: op1_15_inv02 = 1;
    56: op1_15_inv02 = 1;
    57: op1_15_inv02 = 1;
    61: op1_15_inv02 = 1;
    64: op1_15_inv02 = 1;
    65: op1_15_inv02 = 1;
    67: op1_15_inv02 = 1;
    69: op1_15_inv02 = 1;
    72: op1_15_inv02 = 1;
    73: op1_15_inv02 = 1;
    74: op1_15_inv02 = 1;
    75: op1_15_inv02 = 1;
    76: op1_15_inv02 = 1;
    79: op1_15_inv02 = 1;
    80: op1_15_inv02 = 1;
    84: op1_15_inv02 = 1;
    87: op1_15_inv02 = 1;
    90: op1_15_inv02 = 1;
    94: op1_15_inv02 = 1;
    96: op1_15_inv02 = 1;
    default: op1_15_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in03 = imem02_in[71:68];
    6: op1_15_in03 = reg_0724;
    7: op1_15_in03 = imem03_in[107:104];
    8: op1_15_in03 = imem05_in[51:48];
    9: op1_15_in03 = reg_0205;
    10: op1_15_in03 = imem00_in[83:80];
    40: op1_15_in03 = imem00_in[83:80];
    11: op1_15_in03 = reg_0306;
    12: op1_15_in03 = reg_0152;
    13: op1_15_in03 = reg_0991;
    14: op1_15_in03 = reg_0865;
    15: op1_15_in03 = reg_0787;
    16: op1_15_in03 = reg_0105;
    17: op1_15_in03 = reg_0361;
    18: op1_15_in03 = reg_0652;
    19: op1_15_in03 = reg_0387;
    20: op1_15_in03 = reg_0239;
    21: op1_15_in03 = reg_0009;
    22: op1_15_in03 = reg_0026;
    23: op1_15_in03 = reg_0320;
    24: op1_15_in03 = reg_0695;
    25: op1_15_in03 = imem01_in[103:100];
    26: op1_15_in03 = reg_0629;
    27: op1_15_in03 = reg_0792;
    28: op1_15_in03 = imem04_in[99:96];
    91: op1_15_in03 = imem04_in[99:96];
    29: op1_15_in03 = reg_0721;
    4: op1_15_in03 = imem07_in[99:96];
    30: op1_15_in03 = reg_0100;
    31: op1_15_in03 = imem05_in[99:96];
    32: op1_15_in03 = reg_0919;
    33: op1_15_in03 = imem07_in[43:40];
    34: op1_15_in03 = reg_1009;
    35: op1_15_in03 = reg_0528;
    36: op1_15_in03 = reg_0973;
    37: op1_15_in03 = reg_0442;
    38: op1_15_in03 = imem07_in[35:32];
    39: op1_15_in03 = reg_0696;
    41: op1_15_in03 = reg_0817;
    42: op1_15_in03 = imem06_in[31:28];
    43: op1_15_in03 = reg_0166;
    44: op1_15_in03 = reg_0686;
    45: op1_15_in03 = reg_0038;
    46: op1_15_in03 = reg_0889;
    47: op1_15_in03 = imem00_in[79:76];
    62: op1_15_in03 = imem00_in[79:76];
    48: op1_15_in03 = reg_0245;
    49: op1_15_in03 = reg_0568;
    50: op1_15_in03 = reg_0884;
    51: op1_15_in03 = reg_0522;
    83: op1_15_in03 = reg_0522;
    52: op1_15_in03 = reg_0694;
    53: op1_15_in03 = imem02_in[11:8];
    54: op1_15_in03 = reg_0830;
    55: op1_15_in03 = imem04_in[63:60];
    56: op1_15_in03 = imem05_in[87:84];
    57: op1_15_in03 = reg_0944;
    58: op1_15_in03 = reg_0346;
    59: op1_15_in03 = imem07_in[7:4];
    60: op1_15_in03 = imem05_in[103:100];
    61: op1_15_in03 = imem07_in[87:84];
    63: op1_15_in03 = imem03_in[27:24];
    64: op1_15_in03 = reg_0240;
    65: op1_15_in03 = reg_0513;
    66: op1_15_in03 = reg_0524;
    67: op1_15_in03 = imem04_in[11:8];
    68: op1_15_in03 = imem00_in[43:40];
    69: op1_15_in03 = imem02_in[63:60];
    70: op1_15_in03 = reg_0044;
    71: op1_15_in03 = reg_0842;
    72: op1_15_in03 = reg_0979;
    73: op1_15_in03 = reg_0909;
    74: op1_15_in03 = reg_0786;
    75: op1_15_in03 = reg_0289;
    76: op1_15_in03 = reg_0167;
    77: op1_15_in03 = reg_0829;
    78: op1_15_in03 = reg_0377;
    79: op1_15_in03 = reg_0040;
    80: op1_15_in03 = imem06_in[63:60];
    81: op1_15_in03 = reg_0338;
    82: op1_15_in03 = reg_0099;
    84: op1_15_in03 = reg_0738;
    85: op1_15_in03 = reg_0866;
    86: op1_15_in03 = reg_0284;
    87: op1_15_in03 = reg_0877;
    88: op1_15_in03 = reg_0128;
    89: op1_15_in03 = reg_0554;
    90: op1_15_in03 = imem04_in[51:48];
    92: op1_15_in03 = reg_0310;
    93: op1_15_in03 = imem00_in[47:44];
    94: op1_15_in03 = reg_0572;
    96: op1_15_in03 = reg_0174;
    default: op1_15_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv03 = 1;
    8: op1_15_inv03 = 1;
    9: op1_15_inv03 = 1;
    11: op1_15_inv03 = 1;
    17: op1_15_inv03 = 1;
    19: op1_15_inv03 = 1;
    20: op1_15_inv03 = 1;
    21: op1_15_inv03 = 1;
    25: op1_15_inv03 = 1;
    27: op1_15_inv03 = 1;
    31: op1_15_inv03 = 1;
    33: op1_15_inv03 = 1;
    34: op1_15_inv03 = 1;
    35: op1_15_inv03 = 1;
    36: op1_15_inv03 = 1;
    38: op1_15_inv03 = 1;
    39: op1_15_inv03 = 1;
    40: op1_15_inv03 = 1;
    44: op1_15_inv03 = 1;
    45: op1_15_inv03 = 1;
    46: op1_15_inv03 = 1;
    49: op1_15_inv03 = 1;
    52: op1_15_inv03 = 1;
    53: op1_15_inv03 = 1;
    57: op1_15_inv03 = 1;
    62: op1_15_inv03 = 1;
    64: op1_15_inv03 = 1;
    65: op1_15_inv03 = 1;
    66: op1_15_inv03 = 1;
    73: op1_15_inv03 = 1;
    74: op1_15_inv03 = 1;
    77: op1_15_inv03 = 1;
    78: op1_15_inv03 = 1;
    81: op1_15_inv03 = 1;
    82: op1_15_inv03 = 1;
    83: op1_15_inv03 = 1;
    84: op1_15_inv03 = 1;
    86: op1_15_inv03 = 1;
    88: op1_15_inv03 = 1;
    89: op1_15_inv03 = 1;
    90: op1_15_inv03 = 1;
    92: op1_15_inv03 = 1;
    93: op1_15_inv03 = 1;
    96: op1_15_inv03 = 1;
    default: op1_15_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in04 = imem02_in[87:84];
    6: op1_15_in04 = reg_0706;
    7: op1_15_in04 = reg_0582;
    8: op1_15_in04 = imem05_in[67:64];
    9: op1_15_in04 = imem01_in[11:8];
    10: op1_15_in04 = imem00_in[107:104];
    62: op1_15_in04 = imem00_in[107:104];
    11: op1_15_in04 = reg_0276;
    12: op1_15_in04 = reg_0144;
    13: op1_15_in04 = reg_0996;
    14: op1_15_in04 = reg_0254;
    15: op1_15_in04 = reg_0027;
    16: op1_15_in04 = reg_0107;
    17: op1_15_in04 = reg_0396;
    18: op1_15_in04 = reg_0325;
    19: op1_15_in04 = reg_0362;
    20: op1_15_in04 = reg_0735;
    21: op1_15_in04 = reg_0738;
    22: op1_15_in04 = reg_0781;
    23: op1_15_in04 = reg_0354;
    24: op1_15_in04 = reg_0682;
    25: op1_15_in04 = imem01_in[123:120];
    26: op1_15_in04 = reg_0607;
    27: op1_15_in04 = reg_0086;
    28: op1_15_in04 = reg_0063;
    29: op1_15_in04 = reg_0714;
    4: op1_15_in04 = imem07_in[107:104];
    30: op1_15_in04 = reg_0101;
    31: op1_15_in04 = reg_0944;
    32: op1_15_in04 = reg_0928;
    33: op1_15_in04 = imem07_in[51:48];
    34: op1_15_in04 = reg_0888;
    35: op1_15_in04 = reg_0056;
    36: op1_15_in04 = reg_0970;
    37: op1_15_in04 = reg_0438;
    38: op1_15_in04 = imem07_in[39:36];
    39: op1_15_in04 = reg_0694;
    40: op1_15_in04 = imem00_in[119:116];
    41: op1_15_in04 = reg_0338;
    42: op1_15_in04 = imem06_in[71:68];
    43: op1_15_in04 = reg_0170;
    44: op1_15_in04 = reg_0691;
    45: op1_15_in04 = reg_0795;
    46: op1_15_in04 = reg_0293;
    47: op1_15_in04 = imem00_in[83:80];
    48: op1_15_in04 = reg_0576;
    64: op1_15_in04 = reg_0576;
    49: op1_15_in04 = reg_0401;
    50: op1_15_in04 = reg_0872;
    51: op1_15_in04 = reg_0520;
    52: op1_15_in04 = reg_0689;
    53: op1_15_in04 = imem02_in[31:28];
    54: op1_15_in04 = reg_0232;
    55: op1_15_in04 = imem04_in[75:72];
    56: op1_15_in04 = imem05_in[119:116];
    57: op1_15_in04 = reg_0225;
    58: op1_15_in04 = reg_0661;
    59: op1_15_in04 = imem07_in[15:12];
    60: op1_15_in04 = reg_0951;
    61: op1_15_in04 = imem07_in[127:124];
    63: op1_15_in04 = imem03_in[47:44];
    65: op1_15_in04 = reg_0822;
    66: op1_15_in04 = reg_0584;
    67: op1_15_in04 = imem04_in[19:16];
    68: op1_15_in04 = imem00_in[75:72];
    69: op1_15_in04 = imem02_in[71:68];
    70: op1_15_in04 = imem05_in[59:56];
    71: op1_15_in04 = reg_0749;
    72: op1_15_in04 = reg_1001;
    73: op1_15_in04 = reg_0524;
    74: op1_15_in04 = imem05_in[55:52];
    75: op1_15_in04 = reg_0807;
    76: op1_15_in04 = reg_0176;
    77: op1_15_in04 = reg_0514;
    78: op1_15_in04 = reg_0820;
    79: op1_15_in04 = reg_0377;
    80: op1_15_in04 = imem06_in[87:84];
    81: op1_15_in04 = reg_0614;
    82: op1_15_in04 = reg_0760;
    83: op1_15_in04 = reg_0869;
    84: op1_15_in04 = reg_0674;
    85: op1_15_in04 = reg_0954;
    86: op1_15_in04 = reg_0764;
    87: op1_15_in04 = reg_0117;
    88: op1_15_in04 = reg_0142;
    89: op1_15_in04 = reg_0483;
    90: op1_15_in04 = imem04_in[59:56];
    91: op1_15_in04 = imem04_in[115:112];
    92: op1_15_in04 = reg_0453;
    93: op1_15_in04 = imem00_in[51:48];
    94: op1_15_in04 = reg_0867;
    96: op1_15_in04 = reg_0175;
    default: op1_15_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv04 = 1;
    7: op1_15_inv04 = 1;
    8: op1_15_inv04 = 1;
    12: op1_15_inv04 = 1;
    14: op1_15_inv04 = 1;
    15: op1_15_inv04 = 1;
    16: op1_15_inv04 = 1;
    20: op1_15_inv04 = 1;
    22: op1_15_inv04 = 1;
    26: op1_15_inv04 = 1;
    27: op1_15_inv04 = 1;
    31: op1_15_inv04 = 1;
    32: op1_15_inv04 = 1;
    34: op1_15_inv04 = 1;
    35: op1_15_inv04 = 1;
    36: op1_15_inv04 = 1;
    38: op1_15_inv04 = 1;
    42: op1_15_inv04 = 1;
    43: op1_15_inv04 = 1;
    45: op1_15_inv04 = 1;
    46: op1_15_inv04 = 1;
    49: op1_15_inv04 = 1;
    52: op1_15_inv04 = 1;
    54: op1_15_inv04 = 1;
    56: op1_15_inv04 = 1;
    57: op1_15_inv04 = 1;
    59: op1_15_inv04 = 1;
    60: op1_15_inv04 = 1;
    62: op1_15_inv04 = 1;
    65: op1_15_inv04 = 1;
    67: op1_15_inv04 = 1;
    71: op1_15_inv04 = 1;
    72: op1_15_inv04 = 1;
    74: op1_15_inv04 = 1;
    75: op1_15_inv04 = 1;
    76: op1_15_inv04 = 1;
    80: op1_15_inv04 = 1;
    81: op1_15_inv04 = 1;
    82: op1_15_inv04 = 1;
    83: op1_15_inv04 = 1;
    85: op1_15_inv04 = 1;
    88: op1_15_inv04 = 1;
    94: op1_15_inv04 = 1;
    default: op1_15_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の5番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in05 = reg_0651;
    6: op1_15_in05 = reg_0436;
    7: op1_15_in05 = reg_0596;
    8: op1_15_in05 = imem05_in[75:72];
    9: op1_15_in05 = imem01_in[23:20];
    10: op1_15_in05 = reg_0672;
    11: op1_15_in05 = reg_0295;
    12: op1_15_in05 = imem06_in[7:4];
    13: op1_15_in05 = reg_0980;
    79: op1_15_in05 = reg_0980;
    14: op1_15_in05 = reg_0132;
    15: op1_15_in05 = reg_0486;
    16: op1_15_in05 = reg_0126;
    90: op1_15_in05 = reg_0126;
    17: op1_15_in05 = reg_0331;
    18: op1_15_in05 = reg_0347;
    19: op1_15_in05 = reg_0369;
    45: op1_15_in05 = reg_0369;
    75: op1_15_in05 = reg_0369;
    20: op1_15_in05 = reg_0240;
    21: op1_15_in05 = reg_0751;
    22: op1_15_in05 = imem07_in[15:12];
    23: op1_15_in05 = reg_0324;
    24: op1_15_in05 = reg_0693;
    25: op1_15_in05 = reg_1039;
    26: op1_15_in05 = reg_0620;
    27: op1_15_in05 = reg_0090;
    28: op1_15_in05 = reg_0070;
    29: op1_15_in05 = reg_0703;
    4: op1_15_in05 = reg_0441;
    30: op1_15_in05 = reg_0109;
    31: op1_15_in05 = reg_0959;
    32: op1_15_in05 = reg_0754;
    33: op1_15_in05 = imem07_in[95:92];
    34: op1_15_in05 = reg_0541;
    35: op1_15_in05 = reg_0053;
    36: op1_15_in05 = reg_0969;
    37: op1_15_in05 = reg_0179;
    38: op1_15_in05 = imem07_in[47:44];
    39: op1_15_in05 = reg_0679;
    52: op1_15_in05 = reg_0679;
    40: op1_15_in05 = imem00_in[127:124];
    41: op1_15_in05 = reg_0037;
    42: op1_15_in05 = imem06_in[87:84];
    44: op1_15_in05 = reg_0668;
    46: op1_15_in05 = reg_0395;
    47: op1_15_in05 = imem00_in[107:104];
    48: op1_15_in05 = reg_0874;
    64: op1_15_in05 = reg_0874;
    49: op1_15_in05 = reg_0015;
    50: op1_15_in05 = imem03_in[39:36];
    51: op1_15_in05 = reg_0829;
    53: op1_15_in05 = imem02_in[67:64];
    54: op1_15_in05 = reg_1053;
    55: op1_15_in05 = reg_1006;
    56: op1_15_in05 = reg_0215;
    57: op1_15_in05 = reg_0492;
    58: op1_15_in05 = reg_0662;
    59: op1_15_in05 = imem07_in[31:28];
    60: op1_15_in05 = reg_0689;
    61: op1_15_in05 = reg_0718;
    62: op1_15_in05 = reg_0883;
    63: op1_15_in05 = imem03_in[51:48];
    65: op1_15_in05 = reg_0996;
    66: op1_15_in05 = reg_0296;
    67: op1_15_in05 = imem04_in[47:44];
    68: op1_15_in05 = imem00_in[79:76];
    69: op1_15_in05 = imem02_in[91:88];
    70: op1_15_in05 = imem05_in[79:76];
    71: op1_15_in05 = reg_0463;
    72: op1_15_in05 = reg_0986;
    73: op1_15_in05 = reg_0850;
    74: op1_15_in05 = imem05_in[83:80];
    77: op1_15_in05 = reg_0500;
    78: op1_15_in05 = reg_0385;
    80: op1_15_in05 = imem06_in[99:96];
    81: op1_15_in05 = reg_0440;
    82: op1_15_in05 = reg_1007;
    83: op1_15_in05 = reg_0604;
    84: op1_15_in05 = reg_0457;
    85: op1_15_in05 = reg_0143;
    86: op1_15_in05 = reg_0407;
    87: op1_15_in05 = imem02_in[15:12];
    88: op1_15_in05 = reg_0137;
    89: op1_15_in05 = reg_0642;
    91: op1_15_in05 = reg_0147;
    92: op1_15_in05 = reg_0451;
    93: op1_15_in05 = imem00_in[75:72];
    94: op1_15_in05 = reg_0684;
    96: op1_15_in05 = reg_0172;
    default: op1_15_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv05 = 1;
    7: op1_15_inv05 = 1;
    9: op1_15_inv05 = 1;
    11: op1_15_inv05 = 1;
    12: op1_15_inv05 = 1;
    13: op1_15_inv05 = 1;
    15: op1_15_inv05 = 1;
    16: op1_15_inv05 = 1;
    18: op1_15_inv05 = 1;
    20: op1_15_inv05 = 1;
    21: op1_15_inv05 = 1;
    22: op1_15_inv05 = 1;
    23: op1_15_inv05 = 1;
    25: op1_15_inv05 = 1;
    26: op1_15_inv05 = 1;
    27: op1_15_inv05 = 1;
    4: op1_15_inv05 = 1;
    30: op1_15_inv05 = 1;
    31: op1_15_inv05 = 1;
    33: op1_15_inv05 = 1;
    35: op1_15_inv05 = 1;
    38: op1_15_inv05 = 1;
    41: op1_15_inv05 = 1;
    42: op1_15_inv05 = 1;
    44: op1_15_inv05 = 1;
    46: op1_15_inv05 = 1;
    48: op1_15_inv05 = 1;
    50: op1_15_inv05 = 1;
    51: op1_15_inv05 = 1;
    52: op1_15_inv05 = 1;
    54: op1_15_inv05 = 1;
    60: op1_15_inv05 = 1;
    62: op1_15_inv05 = 1;
    63: op1_15_inv05 = 1;
    66: op1_15_inv05 = 1;
    67: op1_15_inv05 = 1;
    69: op1_15_inv05 = 1;
    70: op1_15_inv05 = 1;
    74: op1_15_inv05 = 1;
    75: op1_15_inv05 = 1;
    78: op1_15_inv05 = 1;
    80: op1_15_inv05 = 1;
    81: op1_15_inv05 = 1;
    83: op1_15_inv05 = 1;
    84: op1_15_inv05 = 1;
    86: op1_15_inv05 = 1;
    87: op1_15_inv05 = 1;
    88: op1_15_inv05 = 1;
    96: op1_15_inv05 = 1;
    default: op1_15_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の6番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in06 = reg_0636;
    6: op1_15_in06 = reg_0422;
    4: op1_15_in06 = reg_0422;
    7: op1_15_in06 = reg_0583;
    8: op1_15_in06 = imem05_in[99:96];
    9: op1_15_in06 = imem01_in[35:32];
    10: op1_15_in06 = reg_0686;
    11: op1_15_in06 = reg_0298;
    12: op1_15_in06 = imem06_in[43:40];
    13: op1_15_in06 = reg_0988;
    14: op1_15_in06 = reg_0147;
    15: op1_15_in06 = reg_0753;
    16: op1_15_in06 = imem02_in[11:8];
    17: op1_15_in06 = reg_0984;
    18: op1_15_in06 = reg_0336;
    19: op1_15_in06 = reg_0322;
    20: op1_15_in06 = reg_0502;
    21: op1_15_in06 = reg_0043;
    22: op1_15_in06 = imem07_in[39:36];
    23: op1_15_in06 = reg_0342;
    24: op1_15_in06 = reg_0672;
    25: op1_15_in06 = reg_0216;
    26: op1_15_in06 = reg_0615;
    27: op1_15_in06 = reg_0840;
    28: op1_15_in06 = imem05_in[19:16];
    29: op1_15_in06 = reg_0705;
    30: op1_15_in06 = reg_0127;
    31: op1_15_in06 = reg_0955;
    32: op1_15_in06 = reg_0621;
    33: op1_15_in06 = reg_0702;
    34: op1_15_in06 = reg_0074;
    35: op1_15_in06 = imem05_in[3:0];
    36: op1_15_in06 = reg_0896;
    37: op1_15_in06 = reg_0169;
    38: op1_15_in06 = imem07_in[51:48];
    39: op1_15_in06 = reg_0675;
    40: op1_15_in06 = reg_0695;
    41: op1_15_in06 = imem03_in[35:32];
    42: op1_15_in06 = imem06_in[119:116];
    44: op1_15_in06 = reg_0669;
    45: op1_15_in06 = reg_0509;
    46: op1_15_in06 = reg_0042;
    47: op1_15_in06 = imem00_in[115:112];
    48: op1_15_in06 = reg_0923;
    49: op1_15_in06 = imem04_in[35:32];
    50: op1_15_in06 = imem03_in[63:60];
    51: op1_15_in06 = reg_0514;
    83: op1_15_in06 = reg_0514;
    52: op1_15_in06 = reg_0477;
    53: op1_15_in06 = imem02_in[71:68];
    54: op1_15_in06 = reg_0555;
    55: op1_15_in06 = reg_0306;
    56: op1_15_in06 = reg_0032;
    57: op1_15_in06 = reg_0689;
    58: op1_15_in06 = reg_0576;
    59: op1_15_in06 = imem07_in[67:64];
    60: op1_15_in06 = reg_0943;
    61: op1_15_in06 = reg_0002;
    62: op1_15_in06 = reg_0828;
    63: op1_15_in06 = imem03_in[83:80];
    64: op1_15_in06 = reg_0311;
    65: op1_15_in06 = reg_0986;
    66: op1_15_in06 = reg_0808;
    73: op1_15_in06 = reg_0808;
    67: op1_15_in06 = imem04_in[63:60];
    68: op1_15_in06 = imem00_in[95:92];
    69: op1_15_in06 = imem02_in[107:104];
    70: op1_15_in06 = reg_0970;
    71: op1_15_in06 = reg_0457;
    72: op1_15_in06 = reg_0981;
    74: op1_15_in06 = imem05_in[87:84];
    75: op1_15_in06 = reg_0573;
    77: op1_15_in06 = reg_1037;
    78: op1_15_in06 = reg_0987;
    79: op1_15_in06 = imem04_in[3:0];
    80: op1_15_in06 = imem06_in[111:108];
    81: op1_15_in06 = reg_0395;
    82: op1_15_in06 = reg_0445;
    84: op1_15_in06 = reg_0475;
    85: op1_15_in06 = reg_0057;
    86: op1_15_in06 = reg_0444;
    87: op1_15_in06 = imem02_in[27:24];
    88: op1_15_in06 = reg_0646;
    89: op1_15_in06 = reg_0052;
    90: op1_15_in06 = reg_0405;
    91: op1_15_in06 = reg_0577;
    92: op1_15_in06 = reg_0461;
    93: op1_15_in06 = imem00_in[83:80];
    94: op1_15_in06 = reg_0186;
    96: op1_15_in06 = reg_0731;
    default: op1_15_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv06 = 1;
    9: op1_15_inv06 = 1;
    11: op1_15_inv06 = 1;
    12: op1_15_inv06 = 1;
    20: op1_15_inv06 = 1;
    21: op1_15_inv06 = 1;
    23: op1_15_inv06 = 1;
    24: op1_15_inv06 = 1;
    25: op1_15_inv06 = 1;
    27: op1_15_inv06 = 1;
    28: op1_15_inv06 = 1;
    32: op1_15_inv06 = 1;
    33: op1_15_inv06 = 1;
    34: op1_15_inv06 = 1;
    35: op1_15_inv06 = 1;
    36: op1_15_inv06 = 1;
    37: op1_15_inv06 = 1;
    39: op1_15_inv06 = 1;
    40: op1_15_inv06 = 1;
    44: op1_15_inv06 = 1;
    45: op1_15_inv06 = 1;
    46: op1_15_inv06 = 1;
    50: op1_15_inv06 = 1;
    51: op1_15_inv06 = 1;
    52: op1_15_inv06 = 1;
    53: op1_15_inv06 = 1;
    57: op1_15_inv06 = 1;
    59: op1_15_inv06 = 1;
    60: op1_15_inv06 = 1;
    62: op1_15_inv06 = 1;
    63: op1_15_inv06 = 1;
    64: op1_15_inv06 = 1;
    65: op1_15_inv06 = 1;
    67: op1_15_inv06 = 1;
    68: op1_15_inv06 = 1;
    69: op1_15_inv06 = 1;
    71: op1_15_inv06 = 1;
    72: op1_15_inv06 = 1;
    75: op1_15_inv06 = 1;
    77: op1_15_inv06 = 1;
    79: op1_15_inv06 = 1;
    80: op1_15_inv06 = 1;
    81: op1_15_inv06 = 1;
    82: op1_15_inv06 = 1;
    89: op1_15_inv06 = 1;
    96: op1_15_inv06 = 1;
    default: op1_15_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の7番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in07 = reg_0652;
    6: op1_15_in07 = reg_0440;
    7: op1_15_in07 = reg_0568;
    8: op1_15_in07 = reg_0962;
    9: op1_15_in07 = imem01_in[43:40];
    10: op1_15_in07 = reg_0691;
    11: op1_15_in07 = reg_0061;
    12: op1_15_in07 = imem06_in[67:64];
    13: op1_15_in07 = reg_0997;
    14: op1_15_in07 = reg_0149;
    15: op1_15_in07 = reg_0025;
    16: op1_15_in07 = imem02_in[31:28];
    17: op1_15_in07 = reg_0993;
    78: op1_15_in07 = reg_0993;
    18: op1_15_in07 = reg_0097;
    19: op1_15_in07 = reg_0312;
    20: op1_15_in07 = reg_0248;
    21: op1_15_in07 = imem05_in[75:72];
    22: op1_15_in07 = imem07_in[111:108];
    23: op1_15_in07 = reg_0328;
    24: op1_15_in07 = reg_0676;
    25: op1_15_in07 = reg_1035;
    26: op1_15_in07 = reg_0379;
    27: op1_15_in07 = reg_0484;
    28: op1_15_in07 = imem05_in[95:92];
    29: op1_15_in07 = reg_0424;
    4: op1_15_in07 = reg_0433;
    30: op1_15_in07 = imem02_in[35:32];
    87: op1_15_in07 = imem02_in[35:32];
    31: op1_15_in07 = reg_0954;
    32: op1_15_in07 = reg_0616;
    33: op1_15_in07 = reg_0703;
    96: op1_15_in07 = reg_0703;
    34: op1_15_in07 = reg_0009;
    35: op1_15_in07 = imem05_in[15:12];
    36: op1_15_in07 = reg_0132;
    38: op1_15_in07 = imem07_in[79:76];
    39: op1_15_in07 = reg_0688;
    40: op1_15_in07 = reg_0697;
    41: op1_15_in07 = imem03_in[71:68];
    42: op1_15_in07 = reg_0613;
    44: op1_15_in07 = reg_0478;
    45: op1_15_in07 = reg_0376;
    46: op1_15_in07 = reg_0388;
    47: op1_15_in07 = reg_0693;
    48: op1_15_in07 = reg_0844;
    49: op1_15_in07 = imem04_in[43:40];
    50: op1_15_in07 = imem03_in[67:64];
    51: op1_15_in07 = reg_0830;
    83: op1_15_in07 = reg_0830;
    52: op1_15_in07 = reg_0479;
    53: op1_15_in07 = imem02_in[91:88];
    54: op1_15_in07 = reg_0101;
    55: op1_15_in07 = reg_0539;
    56: op1_15_in07 = reg_0023;
    57: op1_15_in07 = reg_0435;
    58: op1_15_in07 = reg_0370;
    59: op1_15_in07 = imem07_in[123:120];
    60: op1_15_in07 = reg_0022;
    61: op1_15_in07 = reg_0303;
    62: op1_15_in07 = reg_0465;
    63: op1_15_in07 = reg_0012;
    64: op1_15_in07 = reg_0767;
    65: op1_15_in07 = reg_0980;
    66: op1_15_in07 = reg_0074;
    67: op1_15_in07 = imem04_in[79:76];
    68: op1_15_in07 = imem00_in[119:116];
    69: op1_15_in07 = imem02_in[119:116];
    70: op1_15_in07 = reg_0945;
    71: op1_15_in07 = reg_0466;
    72: op1_15_in07 = reg_0988;
    73: op1_15_in07 = reg_0288;
    74: op1_15_in07 = imem05_in[103:100];
    75: op1_15_in07 = reg_0678;
    77: op1_15_in07 = reg_0521;
    79: op1_15_in07 = imem04_in[11:8];
    80: op1_15_in07 = reg_0889;
    81: op1_15_in07 = reg_0008;
    82: op1_15_in07 = reg_0307;
    84: op1_15_in07 = reg_0458;
    85: op1_15_in07 = reg_0667;
    86: op1_15_in07 = reg_0041;
    88: op1_15_in07 = reg_0675;
    89: op1_15_in07 = reg_0423;
    90: op1_15_in07 = reg_0937;
    91: op1_15_in07 = reg_0306;
    92: op1_15_in07 = reg_0477;
    93: op1_15_in07 = imem00_in[107:104];
    94: op1_15_in07 = reg_0310;
    default: op1_15_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv07 = 1;
    8: op1_15_inv07 = 1;
    11: op1_15_inv07 = 1;
    18: op1_15_inv07 = 1;
    20: op1_15_inv07 = 1;
    21: op1_15_inv07 = 1;
    22: op1_15_inv07 = 1;
    24: op1_15_inv07 = 1;
    25: op1_15_inv07 = 1;
    28: op1_15_inv07 = 1;
    29: op1_15_inv07 = 1;
    4: op1_15_inv07 = 1;
    31: op1_15_inv07 = 1;
    39: op1_15_inv07 = 1;
    42: op1_15_inv07 = 1;
    44: op1_15_inv07 = 1;
    45: op1_15_inv07 = 1;
    46: op1_15_inv07 = 1;
    48: op1_15_inv07 = 1;
    49: op1_15_inv07 = 1;
    50: op1_15_inv07 = 1;
    51: op1_15_inv07 = 1;
    53: op1_15_inv07 = 1;
    54: op1_15_inv07 = 1;
    56: op1_15_inv07 = 1;
    58: op1_15_inv07 = 1;
    59: op1_15_inv07 = 1;
    60: op1_15_inv07 = 1;
    66: op1_15_inv07 = 1;
    67: op1_15_inv07 = 1;
    69: op1_15_inv07 = 1;
    71: op1_15_inv07 = 1;
    73: op1_15_inv07 = 1;
    79: op1_15_inv07 = 1;
    80: op1_15_inv07 = 1;
    81: op1_15_inv07 = 1;
    83: op1_15_inv07 = 1;
    84: op1_15_inv07 = 1;
    85: op1_15_inv07 = 1;
    87: op1_15_inv07 = 1;
    88: op1_15_inv07 = 1;
    90: op1_15_inv07 = 1;
    94: op1_15_inv07 = 1;
    default: op1_15_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の8番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in08 = reg_0352;
    6: op1_15_in08 = reg_0444;
    7: op1_15_in08 = reg_0587;
    8: op1_15_in08 = reg_0958;
    9: op1_15_in08 = imem01_in[47:44];
    10: op1_15_in08 = reg_0688;
    11: op1_15_in08 = reg_0046;
    12: op1_15_in08 = imem06_in[111:108];
    13: op1_15_in08 = imem04_in[3:0];
    14: op1_15_in08 = reg_0145;
    15: op1_15_in08 = reg_0805;
    16: op1_15_in08 = imem02_in[39:36];
    17: op1_15_in08 = reg_0975;
    18: op1_15_in08 = reg_0087;
    19: op1_15_in08 = reg_0998;
    20: op1_15_in08 = reg_0507;
    21: op1_15_in08 = imem05_in[91:88];
    22: op1_15_in08 = reg_0716;
    23: op1_15_in08 = reg_0336;
    56: op1_15_in08 = reg_0336;
    24: op1_15_in08 = reg_0670;
    25: op1_15_in08 = reg_1017;
    77: op1_15_in08 = reg_1017;
    26: op1_15_in08 = reg_0405;
    27: op1_15_in08 = reg_0077;
    28: op1_15_in08 = reg_0964;
    29: op1_15_in08 = reg_0432;
    4: op1_15_in08 = reg_0448;
    30: op1_15_in08 = imem02_in[59:56];
    31: op1_15_in08 = reg_0949;
    32: op1_15_in08 = reg_0633;
    33: op1_15_in08 = reg_0709;
    34: op1_15_in08 = reg_0278;
    35: op1_15_in08 = imem05_in[67:64];
    36: op1_15_in08 = reg_0133;
    38: op1_15_in08 = imem07_in[107:104];
    39: op1_15_in08 = reg_0673;
    40: op1_15_in08 = reg_0681;
    47: op1_15_in08 = reg_0681;
    41: op1_15_in08 = imem03_in[95:92];
    42: op1_15_in08 = reg_0220;
    44: op1_15_in08 = reg_0196;
    45: op1_15_in08 = reg_0820;
    46: op1_15_in08 = reg_0894;
    48: op1_15_in08 = reg_0822;
    49: op1_15_in08 = imem04_in[47:44];
    50: op1_15_in08 = imem03_in[83:80];
    51: op1_15_in08 = reg_0227;
    52: op1_15_in08 = reg_0459;
    53: op1_15_in08 = imem02_in[95:92];
    54: op1_15_in08 = reg_0117;
    55: op1_15_in08 = reg_1057;
    57: op1_15_in08 = reg_0094;
    58: op1_15_in08 = reg_0051;
    59: op1_15_in08 = reg_0720;
    60: op1_15_in08 = reg_0757;
    61: op1_15_in08 = reg_0325;
    62: op1_15_in08 = reg_0451;
    63: op1_15_in08 = reg_0099;
    64: op1_15_in08 = reg_0518;
    65: op1_15_in08 = reg_0994;
    78: op1_15_in08 = reg_0994;
    66: op1_15_in08 = reg_0288;
    67: op1_15_in08 = imem04_in[115:112];
    68: op1_15_in08 = reg_0519;
    69: op1_15_in08 = reg_0759;
    70: op1_15_in08 = reg_0343;
    71: op1_15_in08 = reg_0473;
    72: op1_15_in08 = reg_0976;
    73: op1_15_in08 = reg_0027;
    74: op1_15_in08 = imem06_in[87:84];
    75: op1_15_in08 = reg_0569;
    79: op1_15_in08 = imem04_in[79:76];
    80: op1_15_in08 = reg_0392;
    81: op1_15_in08 = reg_0804;
    82: op1_15_in08 = reg_0322;
    83: op1_15_in08 = reg_1037;
    84: op1_15_in08 = reg_0187;
    85: op1_15_in08 = reg_0953;
    86: op1_15_in08 = reg_0065;
    87: op1_15_in08 = imem02_in[43:40];
    88: op1_15_in08 = reg_0152;
    89: op1_15_in08 = reg_0394;
    90: op1_15_in08 = reg_0870;
    91: op1_15_in08 = reg_0864;
    92: op1_15_in08 = reg_0469;
    93: op1_15_in08 = imem00_in[115:112];
    94: op1_15_in08 = reg_0344;
    96: op1_15_in08 = reg_0447;
    default: op1_15_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv08 = 1;
    8: op1_15_inv08 = 1;
    13: op1_15_inv08 = 1;
    15: op1_15_inv08 = 1;
    16: op1_15_inv08 = 1;
    17: op1_15_inv08 = 1;
    20: op1_15_inv08 = 1;
    28: op1_15_inv08 = 1;
    31: op1_15_inv08 = 1;
    32: op1_15_inv08 = 1;
    34: op1_15_inv08 = 1;
    35: op1_15_inv08 = 1;
    44: op1_15_inv08 = 1;
    47: op1_15_inv08 = 1;
    48: op1_15_inv08 = 1;
    50: op1_15_inv08 = 1;
    51: op1_15_inv08 = 1;
    52: op1_15_inv08 = 1;
    53: op1_15_inv08 = 1;
    54: op1_15_inv08 = 1;
    56: op1_15_inv08 = 1;
    59: op1_15_inv08 = 1;
    65: op1_15_inv08 = 1;
    68: op1_15_inv08 = 1;
    69: op1_15_inv08 = 1;
    70: op1_15_inv08 = 1;
    71: op1_15_inv08 = 1;
    74: op1_15_inv08 = 1;
    77: op1_15_inv08 = 1;
    80: op1_15_inv08 = 1;
    81: op1_15_inv08 = 1;
    82: op1_15_inv08 = 1;
    83: op1_15_inv08 = 1;
    85: op1_15_inv08 = 1;
    86: op1_15_inv08 = 1;
    87: op1_15_inv08 = 1;
    89: op1_15_inv08 = 1;
    91: op1_15_inv08 = 1;
    92: op1_15_inv08 = 1;
    93: op1_15_inv08 = 1;
    default: op1_15_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の9番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in09 = reg_0324;
    6: op1_15_in09 = reg_0427;
    7: op1_15_in09 = reg_0592;
    8: op1_15_in09 = reg_0971;
    9: op1_15_in09 = imem01_in[87:84];
    10: op1_15_in09 = reg_0453;
    11: op1_15_in09 = reg_0065;
    12: op1_15_in09 = reg_0630;
    13: op1_15_in09 = imem04_in[7:4];
    14: op1_15_in09 = reg_0136;
    15: op1_15_in09 = imem07_in[23:20];
    16: op1_15_in09 = imem02_in[59:56];
    17: op1_15_in09 = reg_0976;
    18: op1_15_in09 = imem03_in[11:8];
    19: op1_15_in09 = reg_0991;
    20: op1_15_in09 = reg_1032;
    21: op1_15_in09 = reg_0973;
    22: op1_15_in09 = reg_0719;
    23: op1_15_in09 = reg_0776;
    24: op1_15_in09 = reg_0691;
    25: op1_15_in09 = reg_1018;
    26: op1_15_in09 = reg_0375;
    27: op1_15_in09 = reg_0079;
    28: op1_15_in09 = reg_0945;
    29: op1_15_in09 = reg_0426;
    4: op1_15_in09 = reg_0167;
    30: op1_15_in09 = imem02_in[83:80];
    31: op1_15_in09 = reg_0821;
    54: op1_15_in09 = reg_0821;
    32: op1_15_in09 = reg_0632;
    33: op1_15_in09 = reg_0711;
    34: op1_15_in09 = reg_0047;
    35: op1_15_in09 = reg_0966;
    36: op1_15_in09 = reg_0139;
    38: op1_15_in09 = imem07_in[123:120];
    39: op1_15_in09 = reg_0450;
    40: op1_15_in09 = reg_0679;
    41: op1_15_in09 = reg_0938;
    42: op1_15_in09 = reg_0782;
    44: op1_15_in09 = reg_0212;
    45: op1_15_in09 = reg_0246;
    46: op1_15_in09 = reg_0017;
    47: op1_15_in09 = reg_0672;
    48: op1_15_in09 = reg_0988;
    49: op1_15_in09 = imem04_in[55:52];
    50: op1_15_in09 = imem03_in[95:92];
    51: op1_15_in09 = reg_0521;
    52: op1_15_in09 = reg_0200;
    53: op1_15_in09 = imem02_in[99:96];
    55: op1_15_in09 = reg_1005;
    56: op1_15_in09 = reg_0436;
    57: op1_15_in09 = reg_0489;
    58: op1_15_in09 = reg_0376;
    59: op1_15_in09 = reg_0731;
    60: op1_15_in09 = reg_0435;
    61: op1_15_in09 = reg_0350;
    62: op1_15_in09 = reg_0455;
    63: op1_15_in09 = reg_0445;
    64: op1_15_in09 = reg_0822;
    65: op1_15_in09 = imem04_in[11:8];
    66: op1_15_in09 = reg_0764;
    67: op1_15_in09 = imem04_in[123:120];
    68: op1_15_in09 = reg_0686;
    69: op1_15_in09 = reg_0036;
    70: op1_15_in09 = reg_0259;
    71: op1_15_in09 = reg_0474;
    72: op1_15_in09 = imem04_in[35:32];
    73: op1_15_in09 = reg_0251;
    74: op1_15_in09 = imem06_in[115:112];
    75: op1_15_in09 = imem07_in[31:28];
    77: op1_15_in09 = reg_0304;
    78: op1_15_in09 = imem04_in[3:0];
    79: op1_15_in09 = imem04_in[91:88];
    80: op1_15_in09 = reg_0556;
    81: op1_15_in09 = reg_0857;
    93: op1_15_in09 = reg_0857;
    82: op1_15_in09 = reg_0585;
    83: op1_15_in09 = reg_0216;
    84: op1_15_in09 = imem01_in[43:40];
    85: op1_15_in09 = reg_0314;
    86: op1_15_in09 = reg_0027;
    87: op1_15_in09 = imem02_in[91:88];
    88: op1_15_in09 = reg_0023;
    89: op1_15_in09 = reg_0425;
    90: op1_15_in09 = reg_0888;
    91: op1_15_in09 = reg_0799;
    92: op1_15_in09 = reg_0466;
    94: op1_15_in09 = reg_0760;
    96: op1_15_in09 = reg_0182;
    default: op1_15_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv09 = 1;
    6: op1_15_inv09 = 1;
    7: op1_15_inv09 = 1;
    8: op1_15_inv09 = 1;
    10: op1_15_inv09 = 1;
    12: op1_15_inv09 = 1;
    14: op1_15_inv09 = 1;
    16: op1_15_inv09 = 1;
    17: op1_15_inv09 = 1;
    20: op1_15_inv09 = 1;
    23: op1_15_inv09 = 1;
    26: op1_15_inv09 = 1;
    28: op1_15_inv09 = 1;
    29: op1_15_inv09 = 1;
    30: op1_15_inv09 = 1;
    32: op1_15_inv09 = 1;
    38: op1_15_inv09 = 1;
    41: op1_15_inv09 = 1;
    44: op1_15_inv09 = 1;
    46: op1_15_inv09 = 1;
    47: op1_15_inv09 = 1;
    51: op1_15_inv09 = 1;
    55: op1_15_inv09 = 1;
    57: op1_15_inv09 = 1;
    58: op1_15_inv09 = 1;
    59: op1_15_inv09 = 1;
    61: op1_15_inv09 = 1;
    65: op1_15_inv09 = 1;
    68: op1_15_inv09 = 1;
    73: op1_15_inv09 = 1;
    78: op1_15_inv09 = 1;
    83: op1_15_inv09 = 1;
    84: op1_15_inv09 = 1;
    85: op1_15_inv09 = 1;
    88: op1_15_inv09 = 1;
    89: op1_15_inv09 = 1;
    90: op1_15_inv09 = 1;
    92: op1_15_inv09 = 1;
    default: op1_15_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の10番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in10 = reg_0353;
    6: op1_15_in10 = reg_0420;
    7: op1_15_in10 = reg_0591;
    8: op1_15_in10 = reg_0956;
    35: op1_15_in10 = reg_0956;
    9: op1_15_in10 = imem01_in[95:92];
    10: op1_15_in10 = reg_0466;
    11: op1_15_in10 = reg_0058;
    12: op1_15_in10 = reg_0624;
    13: op1_15_in10 = imem04_in[55:52];
    72: op1_15_in10 = imem04_in[55:52];
    14: op1_15_in10 = reg_0150;
    15: op1_15_in10 = imem07_in[95:92];
    16: op1_15_in10 = imem02_in[91:88];
    17: op1_15_in10 = reg_0994;
    18: op1_15_in10 = imem03_in[35:32];
    19: op1_15_in10 = reg_0979;
    20: op1_15_in10 = reg_1040;
    83: op1_15_in10 = reg_1040;
    21: op1_15_in10 = reg_0958;
    22: op1_15_in10 = reg_0731;
    23: op1_15_in10 = reg_0079;
    24: op1_15_in10 = reg_0465;
    25: op1_15_in10 = reg_0123;
    26: op1_15_in10 = reg_0399;
    27: op1_15_in10 = imem03_in[3:0];
    28: op1_15_in10 = reg_0946;
    29: op1_15_in10 = reg_0418;
    4: op1_15_in10 = reg_0183;
    30: op1_15_in10 = imem02_in[87:84];
    31: op1_15_in10 = reg_0831;
    32: op1_15_in10 = reg_0627;
    33: op1_15_in10 = reg_0432;
    34: op1_15_in10 = reg_0875;
    36: op1_15_in10 = reg_0140;
    38: op1_15_in10 = reg_0730;
    39: op1_15_in10 = reg_0471;
    40: op1_15_in10 = reg_0677;
    41: op1_15_in10 = reg_0833;
    42: op1_15_in10 = reg_0385;
    44: op1_15_in10 = imem01_in[59:56];
    45: op1_15_in10 = reg_0234;
    46: op1_15_in10 = reg_1010;
    47: op1_15_in10 = reg_0680;
    48: op1_15_in10 = reg_0976;
    49: op1_15_in10 = imem04_in[95:92];
    50: op1_15_in10 = imem03_in[99:96];
    51: op1_15_in10 = reg_0354;
    52: op1_15_in10 = reg_0203;
    53: op1_15_in10 = imem02_in[107:104];
    54: op1_15_in10 = imem02_in[47:44];
    55: op1_15_in10 = reg_0292;
    56: op1_15_in10 = reg_1046;
    57: op1_15_in10 = reg_0151;
    58: op1_15_in10 = reg_0984;
    59: op1_15_in10 = reg_0721;
    60: op1_15_in10 = reg_0497;
    61: op1_15_in10 = reg_0868;
    62: op1_15_in10 = reg_0200;
    63: op1_15_in10 = reg_0434;
    64: op1_15_in10 = reg_0980;
    65: op1_15_in10 = imem04_in[79:76];
    66: op1_15_in10 = reg_0243;
    67: op1_15_in10 = reg_0265;
    68: op1_15_in10 = reg_0753;
    69: op1_15_in10 = reg_0837;
    70: op1_15_in10 = reg_0125;
    71: op1_15_in10 = reg_0478;
    73: op1_15_in10 = reg_0542;
    74: op1_15_in10 = imem06_in[123:120];
    75: op1_15_in10 = imem07_in[83:80];
    77: op1_15_in10 = reg_1051;
    78: op1_15_in10 = imem04_in[7:4];
    79: op1_15_in10 = imem04_in[103:100];
    80: op1_15_in10 = reg_0863;
    81: op1_15_in10 = reg_0293;
    82: op1_15_in10 = reg_0298;
    84: op1_15_in10 = imem01_in[63:60];
    85: op1_15_in10 = reg_0892;
    86: op1_15_in10 = reg_0777;
    87: op1_15_in10 = imem02_in[95:92];
    88: op1_15_in10 = reg_0272;
    89: op1_15_in10 = reg_0045;
    90: op1_15_in10 = reg_0008;
    91: op1_15_in10 = reg_0802;
    92: op1_15_in10 = reg_0475;
    93: op1_15_in10 = reg_0166;
    94: op1_15_in10 = reg_0132;
    96: op1_15_in10 = reg_0339;
    default: op1_15_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv10 = 1;
    8: op1_15_inv10 = 1;
    11: op1_15_inv10 = 1;
    12: op1_15_inv10 = 1;
    13: op1_15_inv10 = 1;
    14: op1_15_inv10 = 1;
    15: op1_15_inv10 = 1;
    16: op1_15_inv10 = 1;
    17: op1_15_inv10 = 1;
    18: op1_15_inv10 = 1;
    20: op1_15_inv10 = 1;
    21: op1_15_inv10 = 1;
    22: op1_15_inv10 = 1;
    26: op1_15_inv10 = 1;
    4: op1_15_inv10 = 1;
    33: op1_15_inv10 = 1;
    34: op1_15_inv10 = 1;
    36: op1_15_inv10 = 1;
    38: op1_15_inv10 = 1;
    39: op1_15_inv10 = 1;
    42: op1_15_inv10 = 1;
    45: op1_15_inv10 = 1;
    46: op1_15_inv10 = 1;
    47: op1_15_inv10 = 1;
    49: op1_15_inv10 = 1;
    50: op1_15_inv10 = 1;
    55: op1_15_inv10 = 1;
    56: op1_15_inv10 = 1;
    57: op1_15_inv10 = 1;
    60: op1_15_inv10 = 1;
    63: op1_15_inv10 = 1;
    65: op1_15_inv10 = 1;
    70: op1_15_inv10 = 1;
    77: op1_15_inv10 = 1;
    79: op1_15_inv10 = 1;
    80: op1_15_inv10 = 1;
    83: op1_15_inv10 = 1;
    84: op1_15_inv10 = 1;
    88: op1_15_inv10 = 1;
    89: op1_15_inv10 = 1;
    90: op1_15_inv10 = 1;
    94: op1_15_inv10 = 1;
    default: op1_15_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in11 = reg_0342;
    6: op1_15_in11 = reg_0174;
    7: op1_15_in11 = reg_0597;
    8: op1_15_in11 = reg_0948;
    9: op1_15_in11 = imem01_in[111:108];
    10: op1_15_in11 = reg_0480;
    11: op1_15_in11 = reg_0076;
    12: op1_15_in11 = reg_0621;
    13: op1_15_in11 = imem04_in[59:56];
    72: op1_15_in11 = imem04_in[59:56];
    14: op1_15_in11 = reg_0143;
    15: op1_15_in11 = imem07_in[127:124];
    16: op1_15_in11 = imem02_in[111:108];
    17: op1_15_in11 = imem04_in[39:36];
    18: op1_15_in11 = imem03_in[43:40];
    19: op1_15_in11 = reg_0980;
    58: op1_15_in11 = reg_0980;
    20: op1_15_in11 = reg_0913;
    21: op1_15_in11 = reg_0969;
    22: op1_15_in11 = reg_0721;
    23: op1_15_in11 = imem03_in[67:64];
    24: op1_15_in11 = reg_0453;
    25: op1_15_in11 = reg_0105;
    26: op1_15_in11 = reg_0406;
    27: op1_15_in11 = imem03_in[11:8];
    28: op1_15_in11 = reg_0961;
    29: op1_15_in11 = reg_0437;
    4: op1_15_in11 = reg_0166;
    30: op1_15_in11 = imem02_in[95:92];
    31: op1_15_in11 = reg_0136;
    32: op1_15_in11 = reg_0385;
    33: op1_15_in11 = reg_0427;
    34: op1_15_in11 = reg_0021;
    35: op1_15_in11 = reg_0946;
    36: op1_15_in11 = reg_0155;
    38: op1_15_in11 = reg_0710;
    39: op1_15_in11 = reg_0200;
    40: op1_15_in11 = reg_0678;
    41: op1_15_in11 = reg_0373;
    42: op1_15_in11 = reg_0351;
    44: op1_15_in11 = imem01_in[103:100];
    45: op1_15_in11 = reg_0977;
    46: op1_15_in11 = reg_0633;
    47: op1_15_in11 = reg_0673;
    48: op1_15_in11 = imem04_in[7:4];
    49: op1_15_in11 = imem05_in[27:24];
    50: op1_15_in11 = imem03_in[103:100];
    51: op1_15_in11 = reg_0610;
    52: op1_15_in11 = reg_0201;
    53: op1_15_in11 = imem02_in[119:116];
    54: op1_15_in11 = imem02_in[87:84];
    55: op1_15_in11 = reg_0888;
    56: op1_15_in11 = reg_0148;
    57: op1_15_in11 = reg_0156;
    59: op1_15_in11 = reg_0705;
    60: op1_15_in11 = reg_0133;
    61: op1_15_in11 = reg_0172;
    62: op1_15_in11 = reg_0187;
    63: op1_15_in11 = reg_0346;
    64: op1_15_in11 = reg_1000;
    65: op1_15_in11 = imem04_in[91:88];
    66: op1_15_in11 = reg_0041;
    67: op1_15_in11 = reg_0277;
    68: op1_15_in11 = reg_0687;
    69: op1_15_in11 = reg_0052;
    70: op1_15_in11 = reg_0865;
    71: op1_15_in11 = reg_0211;
    73: op1_15_in11 = reg_0531;
    74: op1_15_in11 = reg_0694;
    75: op1_15_in11 = reg_0361;
    77: op1_15_in11 = reg_0769;
    78: op1_15_in11 = imem04_in[11:8];
    79: op1_15_in11 = imem04_in[107:104];
    80: op1_15_in11 = reg_0222;
    81: op1_15_in11 = reg_0485;
    82: op1_15_in11 = reg_0396;
    83: op1_15_in11 = reg_1041;
    84: op1_15_in11 = imem01_in[119:116];
    85: op1_15_in11 = reg_0486;
    86: op1_15_in11 = reg_0251;
    87: op1_15_in11 = imem02_in[103:100];
    88: op1_15_in11 = reg_0736;
    89: op1_15_in11 = reg_0776;
    90: op1_15_in11 = reg_0882;
    91: op1_15_in11 = reg_0848;
    92: op1_15_in11 = reg_0203;
    93: op1_15_in11 = reg_0899;
    94: op1_15_in11 = reg_0810;
    96: op1_15_in11 = reg_0183;
    default: op1_15_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv11 = 1;
    6: op1_15_inv11 = 1;
    7: op1_15_inv11 = 1;
    8: op1_15_inv11 = 1;
    9: op1_15_inv11 = 1;
    10: op1_15_inv11 = 1;
    11: op1_15_inv11 = 1;
    12: op1_15_inv11 = 1;
    14: op1_15_inv11 = 1;
    16: op1_15_inv11 = 1;
    18: op1_15_inv11 = 1;
    22: op1_15_inv11 = 1;
    23: op1_15_inv11 = 1;
    24: op1_15_inv11 = 1;
    26: op1_15_inv11 = 1;
    30: op1_15_inv11 = 1;
    32: op1_15_inv11 = 1;
    33: op1_15_inv11 = 1;
    34: op1_15_inv11 = 1;
    35: op1_15_inv11 = 1;
    38: op1_15_inv11 = 1;
    40: op1_15_inv11 = 1;
    49: op1_15_inv11 = 1;
    51: op1_15_inv11 = 1;
    53: op1_15_inv11 = 1;
    54: op1_15_inv11 = 1;
    55: op1_15_inv11 = 1;
    57: op1_15_inv11 = 1;
    58: op1_15_inv11 = 1;
    61: op1_15_inv11 = 1;
    64: op1_15_inv11 = 1;
    66: op1_15_inv11 = 1;
    67: op1_15_inv11 = 1;
    68: op1_15_inv11 = 1;
    71: op1_15_inv11 = 1;
    74: op1_15_inv11 = 1;
    75: op1_15_inv11 = 1;
    78: op1_15_inv11 = 1;
    79: op1_15_inv11 = 1;
    80: op1_15_inv11 = 1;
    81: op1_15_inv11 = 1;
    82: op1_15_inv11 = 1;
    84: op1_15_inv11 = 1;
    85: op1_15_inv11 = 1;
    86: op1_15_inv11 = 1;
    88: op1_15_inv11 = 1;
    89: op1_15_inv11 = 1;
    91: op1_15_inv11 = 1;
    92: op1_15_inv11 = 1;
    96: op1_15_inv11 = 1;
    default: op1_15_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in12 = reg_0083;
    6: op1_15_in12 = reg_0181;
    7: op1_15_in12 = reg_0588;
    8: op1_15_in12 = reg_0267;
    9: op1_15_in12 = imem01_in[127:124];
    10: op1_15_in12 = reg_0473;
    11: op1_15_in12 = reg_0043;
    12: op1_15_in12 = reg_0619;
    13: op1_15_in12 = imem04_in[67:64];
    14: op1_15_in12 = reg_0155;
    15: op1_15_in12 = reg_0719;
    16: op1_15_in12 = reg_0642;
    17: op1_15_in12 = imem04_in[99:96];
    18: op1_15_in12 = imem03_in[91:88];
    19: op1_15_in12 = reg_0899;
    20: op1_15_in12 = reg_1038;
    21: op1_15_in12 = reg_0968;
    22: op1_15_in12 = reg_0729;
    23: op1_15_in12 = imem03_in[119:116];
    24: op1_15_in12 = reg_0469;
    25: op1_15_in12 = reg_0108;
    26: op1_15_in12 = reg_0380;
    27: op1_15_in12 = imem03_in[15:12];
    28: op1_15_in12 = reg_0960;
    29: op1_15_in12 = reg_0420;
    4: op1_15_in12 = reg_0178;
    30: op1_15_in12 = reg_0653;
    31: op1_15_in12 = reg_0133;
    32: op1_15_in12 = reg_0387;
    33: op1_15_in12 = reg_0431;
    34: op1_15_in12 = imem05_in[7:4];
    35: op1_15_in12 = reg_0952;
    36: op1_15_in12 = reg_0137;
    57: op1_15_in12 = reg_0137;
    38: op1_15_in12 = reg_0724;
    39: op1_15_in12 = reg_0210;
    40: op1_15_in12 = reg_0468;
    41: op1_15_in12 = reg_0807;
    42: op1_15_in12 = reg_0388;
    44: op1_15_in12 = imem01_in[111:108];
    45: op1_15_in12 = reg_0975;
    46: op1_15_in12 = reg_0005;
    47: op1_15_in12 = reg_0669;
    48: op1_15_in12 = imem04_in[15:12];
    49: op1_15_in12 = imem05_in[39:36];
    50: op1_15_in12 = reg_0940;
    51: op1_15_in12 = reg_1017;
    83: op1_15_in12 = reg_1017;
    52: op1_15_in12 = reg_0192;
    53: op1_15_in12 = reg_0355;
    54: op1_15_in12 = imem02_in[91:88];
    55: op1_15_in12 = reg_0931;
    56: op1_15_in12 = reg_0135;
    58: op1_15_in12 = reg_0974;
    59: op1_15_in12 = reg_0325;
    60: op1_15_in12 = reg_0139;
    61: op1_15_in12 = reg_0170;
    62: op1_15_in12 = reg_0194;
    92: op1_15_in12 = reg_0194;
    63: op1_15_in12 = reg_0847;
    64: op1_15_in12 = reg_0983;
    65: op1_15_in12 = imem04_in[111:108];
    66: op1_15_in12 = reg_0065;
    67: op1_15_in12 = reg_0306;
    68: op1_15_in12 = reg_0749;
    69: op1_15_in12 = reg_0329;
    70: op1_15_in12 = reg_0004;
    71: op1_15_in12 = reg_0206;
    72: op1_15_in12 = imem04_in[87:84];
    73: op1_15_in12 = reg_0042;
    74: op1_15_in12 = reg_0696;
    75: op1_15_in12 = reg_0575;
    77: op1_15_in12 = reg_0111;
    78: op1_15_in12 = imem04_in[27:24];
    79: op1_15_in12 = reg_1005;
    80: op1_15_in12 = reg_0857;
    81: op1_15_in12 = reg_0403;
    82: op1_15_in12 = reg_0823;
    84: op1_15_in12 = reg_1023;
    85: op1_15_in12 = reg_0146;
    86: op1_15_in12 = imem05_in[11:8];
    87: op1_15_in12 = imem02_in[119:116];
    88: op1_15_in12 = reg_0831;
    89: op1_15_in12 = reg_0656;
    90: op1_15_in12 = reg_0586;
    91: op1_15_in12 = reg_0568;
    93: op1_15_in12 = reg_0344;
    94: op1_15_in12 = reg_0455;
    96: op1_15_in12 = reg_0701;
    default: op1_15_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv12 = 1;
    7: op1_15_inv12 = 1;
    10: op1_15_inv12 = 1;
    13: op1_15_inv12 = 1;
    14: op1_15_inv12 = 1;
    15: op1_15_inv12 = 1;
    17: op1_15_inv12 = 1;
    19: op1_15_inv12 = 1;
    20: op1_15_inv12 = 1;
    22: op1_15_inv12 = 1;
    23: op1_15_inv12 = 1;
    24: op1_15_inv12 = 1;
    26: op1_15_inv12 = 1;
    27: op1_15_inv12 = 1;
    4: op1_15_inv12 = 1;
    34: op1_15_inv12 = 1;
    35: op1_15_inv12 = 1;
    36: op1_15_inv12 = 1;
    38: op1_15_inv12 = 1;
    41: op1_15_inv12 = 1;
    48: op1_15_inv12 = 1;
    49: op1_15_inv12 = 1;
    50: op1_15_inv12 = 1;
    54: op1_15_inv12 = 1;
    55: op1_15_inv12 = 1;
    60: op1_15_inv12 = 1;
    62: op1_15_inv12 = 1;
    63: op1_15_inv12 = 1;
    66: op1_15_inv12 = 1;
    68: op1_15_inv12 = 1;
    70: op1_15_inv12 = 1;
    72: op1_15_inv12 = 1;
    73: op1_15_inv12 = 1;
    74: op1_15_inv12 = 1;
    75: op1_15_inv12 = 1;
    77: op1_15_inv12 = 1;
    82: op1_15_inv12 = 1;
    84: op1_15_inv12 = 1;
    85: op1_15_inv12 = 1;
    86: op1_15_inv12 = 1;
    87: op1_15_inv12 = 1;
    88: op1_15_inv12 = 1;
    default: op1_15_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in13 = reg_0081;
    6: op1_15_in13 = reg_0160;
    7: op1_15_in13 = reg_0384;
    42: op1_15_in13 = reg_0384;
    8: op1_15_in13 = reg_0241;
    9: op1_15_in13 = reg_0504;
    10: op1_15_in13 = reg_0470;
    11: op1_15_in13 = reg_0072;
    12: op1_15_in13 = reg_0612;
    13: op1_15_in13 = imem04_in[71:68];
    14: op1_15_in13 = imem06_in[31:28];
    15: op1_15_in13 = reg_0705;
    38: op1_15_in13 = reg_0705;
    16: op1_15_in13 = reg_0658;
    17: op1_15_in13 = imem04_in[119:116];
    78: op1_15_in13 = imem04_in[119:116];
    18: op1_15_in13 = imem03_in[115:112];
    19: op1_15_in13 = reg_0282;
    65: op1_15_in13 = reg_0282;
    20: op1_15_in13 = reg_0123;
    21: op1_15_in13 = reg_0953;
    22: op1_15_in13 = reg_0713;
    23: op1_15_in13 = reg_0571;
    24: op1_15_in13 = reg_0473;
    25: op1_15_in13 = reg_0100;
    26: op1_15_in13 = reg_1030;
    27: op1_15_in13 = imem03_in[31:28];
    28: op1_15_in13 = reg_0827;
    29: op1_15_in13 = reg_0172;
    30: op1_15_in13 = reg_0637;
    31: op1_15_in13 = reg_0150;
    32: op1_15_in13 = reg_0042;
    33: op1_15_in13 = reg_0179;
    34: op1_15_in13 = imem05_in[15:12];
    35: op1_15_in13 = reg_0972;
    36: op1_15_in13 = reg_0613;
    39: op1_15_in13 = reg_0187;
    40: op1_15_in13 = reg_0452;
    41: op1_15_in13 = reg_0234;
    44: op1_15_in13 = reg_0786;
    45: op1_15_in13 = reg_0988;
    46: op1_15_in13 = imem07_in[11:8];
    47: op1_15_in13 = reg_0465;
    48: op1_15_in13 = imem04_in[19:16];
    49: op1_15_in13 = imem05_in[47:44];
    50: op1_15_in13 = reg_1050;
    51: op1_15_in13 = reg_0304;
    52: op1_15_in13 = imem01_in[3:0];
    53: op1_15_in13 = reg_0646;
    54: op1_15_in13 = imem02_in[127:124];
    55: op1_15_in13 = reg_0799;
    56: op1_15_in13 = reg_0128;
    57: op1_15_in13 = reg_0071;
    58: op1_15_in13 = reg_0977;
    59: op1_15_in13 = reg_0426;
    60: op1_15_in13 = reg_0129;
    62: op1_15_in13 = reg_0201;
    63: op1_15_in13 = reg_0543;
    64: op1_15_in13 = reg_0976;
    66: op1_15_in13 = reg_0517;
    67: op1_15_in13 = reg_1005;
    68: op1_15_in13 = reg_0463;
    69: op1_15_in13 = reg_0394;
    70: op1_15_in13 = reg_0947;
    71: op1_15_in13 = imem01_in[59:56];
    72: op1_15_in13 = imem04_in[111:108];
    73: op1_15_in13 = reg_0509;
    74: op1_15_in13 = reg_0391;
    75: op1_15_in13 = reg_0315;
    77: op1_15_in13 = reg_0860;
    79: op1_15_in13 = reg_0292;
    80: op1_15_in13 = reg_0289;
    81: op1_15_in13 = reg_0369;
    82: op1_15_in13 = reg_0756;
    83: op1_15_in13 = reg_0906;
    84: op1_15_in13 = reg_0503;
    85: op1_15_in13 = reg_0528;
    86: op1_15_in13 = imem05_in[27:24];
    87: op1_15_in13 = reg_0090;
    88: op1_15_in13 = reg_0486;
    89: op1_15_in13 = reg_0365;
    90: op1_15_in13 = reg_0752;
    91: op1_15_in13 = reg_0524;
    92: op1_15_in13 = reg_0213;
    93: op1_15_in13 = reg_0680;
    94: op1_15_in13 = reg_0474;
    96: op1_15_in13 = reg_0529;
    default: op1_15_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv13 = 1;
    10: op1_15_inv13 = 1;
    11: op1_15_inv13 = 1;
    12: op1_15_inv13 = 1;
    13: op1_15_inv13 = 1;
    14: op1_15_inv13 = 1;
    15: op1_15_inv13 = 1;
    16: op1_15_inv13 = 1;
    18: op1_15_inv13 = 1;
    20: op1_15_inv13 = 1;
    21: op1_15_inv13 = 1;
    24: op1_15_inv13 = 1;
    30: op1_15_inv13 = 1;
    32: op1_15_inv13 = 1;
    33: op1_15_inv13 = 1;
    36: op1_15_inv13 = 1;
    38: op1_15_inv13 = 1;
    39: op1_15_inv13 = 1;
    40: op1_15_inv13 = 1;
    44: op1_15_inv13 = 1;
    45: op1_15_inv13 = 1;
    46: op1_15_inv13 = 1;
    47: op1_15_inv13 = 1;
    52: op1_15_inv13 = 1;
    53: op1_15_inv13 = 1;
    55: op1_15_inv13 = 1;
    56: op1_15_inv13 = 1;
    57: op1_15_inv13 = 1;
    58: op1_15_inv13 = 1;
    59: op1_15_inv13 = 1;
    60: op1_15_inv13 = 1;
    62: op1_15_inv13 = 1;
    63: op1_15_inv13 = 1;
    64: op1_15_inv13 = 1;
    65: op1_15_inv13 = 1;
    66: op1_15_inv13 = 1;
    67: op1_15_inv13 = 1;
    68: op1_15_inv13 = 1;
    70: op1_15_inv13 = 1;
    71: op1_15_inv13 = 1;
    72: op1_15_inv13 = 1;
    73: op1_15_inv13 = 1;
    74: op1_15_inv13 = 1;
    77: op1_15_inv13 = 1;
    84: op1_15_inv13 = 1;
    91: op1_15_inv13 = 1;
    92: op1_15_inv13 = 1;
    94: op1_15_inv13 = 1;
    default: op1_15_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in14 = reg_0086;
    6: op1_15_in14 = reg_0183;
    7: op1_15_in14 = reg_0362;
    8: op1_15_in14 = reg_0148;
    9: op1_15_in14 = reg_0512;
    10: op1_15_in14 = reg_0452;
    11: op1_15_in14 = imem05_in[43:40];
    12: op1_15_in14 = reg_0408;
    13: op1_15_in14 = imem04_in[75:72];
    14: op1_15_in14 = imem06_in[51:48];
    15: op1_15_in14 = reg_0713;
    38: op1_15_in14 = reg_0713;
    16: op1_15_in14 = reg_0653;
    17: op1_15_in14 = reg_0552;
    18: op1_15_in14 = reg_0586;
    19: op1_15_in14 = reg_0041;
    20: op1_15_in14 = reg_0127;
    21: op1_15_in14 = reg_0821;
    22: op1_15_in14 = reg_0430;
    23: op1_15_in14 = reg_0580;
    24: op1_15_in14 = reg_0456;
    25: op1_15_in14 = reg_0101;
    26: op1_15_in14 = reg_0800;
    27: op1_15_in14 = imem03_in[51:48];
    28: op1_15_in14 = reg_0254;
    29: op1_15_in14 = reg_0160;
    30: op1_15_in14 = reg_0649;
    31: op1_15_in14 = reg_0151;
    32: op1_15_in14 = reg_0392;
    33: op1_15_in14 = reg_0167;
    34: op1_15_in14 = imem05_in[39:36];
    35: op1_15_in14 = reg_0960;
    36: op1_15_in14 = reg_1030;
    39: op1_15_in14 = reg_0193;
    40: op1_15_in14 = reg_0200;
    41: op1_15_in14 = reg_1001;
    42: op1_15_in14 = reg_0625;
    44: op1_15_in14 = reg_0487;
    45: op1_15_in14 = reg_1000;
    46: op1_15_in14 = imem07_in[23:20];
    47: op1_15_in14 = reg_0461;
    48: op1_15_in14 = imem04_in[23:20];
    49: op1_15_in14 = imem05_in[67:64];
    50: op1_15_in14 = reg_0317;
    51: op1_15_in14 = reg_0111;
    52: op1_15_in14 = imem01_in[55:52];
    53: op1_15_in14 = reg_0082;
    54: op1_15_in14 = reg_0642;
    55: op1_15_in14 = reg_0076;
    56: op1_15_in14 = reg_0140;
    57: op1_15_in14 = reg_0915;
    58: op1_15_in14 = reg_0988;
    59: op1_15_in14 = reg_0599;
    60: op1_15_in14 = reg_0144;
    62: op1_15_in14 = reg_0213;
    63: op1_15_in14 = reg_0795;
    64: op1_15_in14 = imem04_in[7:4];
    65: op1_15_in14 = reg_0306;
    66: op1_15_in14 = reg_0973;
    67: op1_15_in14 = reg_1016;
    68: op1_15_in14 = reg_0465;
    69: op1_15_in14 = reg_0368;
    70: op1_15_in14 = reg_0438;
    71: op1_15_in14 = imem01_in[63:60];
    72: op1_15_in14 = reg_0931;
    73: op1_15_in14 = reg_0892;
    74: op1_15_in14 = reg_0262;
    75: op1_15_in14 = reg_0868;
    77: op1_15_in14 = reg_0109;
    78: op1_15_in14 = reg_1009;
    79: op1_15_in14 = reg_0050;
    80: op1_15_in14 = reg_0026;
    81: op1_15_in14 = reg_0095;
    82: op1_15_in14 = reg_0596;
    83: op1_15_in14 = reg_1055;
    84: op1_15_in14 = reg_1024;
    85: op1_15_in14 = reg_0950;
    86: op1_15_in14 = imem05_in[79:76];
    87: op1_15_in14 = reg_0348;
    88: op1_15_in14 = reg_0651;
    89: op1_15_in14 = reg_0367;
    90: op1_15_in14 = reg_0014;
    91: op1_15_in14 = reg_0850;
    92: op1_15_in14 = reg_0190;
    93: op1_15_in14 = reg_0453;
    94: op1_15_in14 = reg_0468;
    96: op1_15_in14 = reg_0171;
    default: op1_15_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv14 = 1;
    14: op1_15_inv14 = 1;
    15: op1_15_inv14 = 1;
    17: op1_15_inv14 = 1;
    22: op1_15_inv14 = 1;
    23: op1_15_inv14 = 1;
    27: op1_15_inv14 = 1;
    28: op1_15_inv14 = 1;
    30: op1_15_inv14 = 1;
    31: op1_15_inv14 = 1;
    32: op1_15_inv14 = 1;
    33: op1_15_inv14 = 1;
    34: op1_15_inv14 = 1;
    38: op1_15_inv14 = 1;
    39: op1_15_inv14 = 1;
    40: op1_15_inv14 = 1;
    41: op1_15_inv14 = 1;
    42: op1_15_inv14 = 1;
    45: op1_15_inv14 = 1;
    50: op1_15_inv14 = 1;
    51: op1_15_inv14 = 1;
    55: op1_15_inv14 = 1;
    57: op1_15_inv14 = 1;
    62: op1_15_inv14 = 1;
    63: op1_15_inv14 = 1;
    64: op1_15_inv14 = 1;
    66: op1_15_inv14 = 1;
    67: op1_15_inv14 = 1;
    68: op1_15_inv14 = 1;
    72: op1_15_inv14 = 1;
    73: op1_15_inv14 = 1;
    78: op1_15_inv14 = 1;
    79: op1_15_inv14 = 1;
    80: op1_15_inv14 = 1;
    82: op1_15_inv14 = 1;
    83: op1_15_inv14 = 1;
    85: op1_15_inv14 = 1;
    87: op1_15_inv14 = 1;
    88: op1_15_inv14 = 1;
    89: op1_15_inv14 = 1;
    91: op1_15_inv14 = 1;
    92: op1_15_inv14 = 1;
    93: op1_15_inv14 = 1;
    96: op1_15_inv14 = 1;
    default: op1_15_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in15 = reg_0087;
    44: op1_15_in15 = reg_0087;
    7: op1_15_in15 = reg_0322;
    8: op1_15_in15 = reg_0154;
    9: op1_15_in15 = reg_0511;
    10: op1_15_in15 = reg_0200;
    11: op1_15_in15 = imem05_in[59:56];
    12: op1_15_in15 = reg_0386;
    13: op1_15_in15 = imem04_in[127:124];
    14: op1_15_in15 = reg_0613;
    15: op1_15_in15 = reg_0707;
    16: op1_15_in15 = reg_0664;
    17: op1_15_in15 = reg_0529;
    18: op1_15_in15 = reg_0585;
    19: op1_15_in15 = reg_0559;
    20: op1_15_in15 = reg_0126;
    21: op1_15_in15 = reg_0835;
    22: op1_15_in15 = reg_0419;
    23: op1_15_in15 = reg_0387;
    24: op1_15_in15 = reg_0214;
    25: op1_15_in15 = reg_0115;
    26: op1_15_in15 = reg_0753;
    27: op1_15_in15 = imem03_in[67:64];
    28: op1_15_in15 = reg_0132;
    29: op1_15_in15 = reg_0163;
    30: op1_15_in15 = reg_0652;
    31: op1_15_in15 = reg_0144;
    32: op1_15_in15 = reg_0351;
    33: op1_15_in15 = reg_0177;
    34: op1_15_in15 = imem05_in[43:40];
    35: op1_15_in15 = reg_0826;
    36: op1_15_in15 = reg_0026;
    38: op1_15_in15 = reg_0718;
    39: op1_15_in15 = reg_0207;
    40: op1_15_in15 = reg_0210;
    41: op1_15_in15 = reg_0976;
    42: op1_15_in15 = reg_0017;
    45: op1_15_in15 = imem04_in[35:32];
    46: op1_15_in15 = imem07_in[39:36];
    47: op1_15_in15 = reg_0481;
    48: op1_15_in15 = imem04_in[39:36];
    49: op1_15_in15 = imem05_in[95:92];
    50: op1_15_in15 = reg_1019;
    51: op1_15_in15 = reg_0116;
    52: op1_15_in15 = imem01_in[67:64];
    53: op1_15_in15 = reg_0637;
    54: op1_15_in15 = reg_0657;
    55: op1_15_in15 = reg_0014;
    56: op1_15_in15 = reg_0155;
    57: op1_15_in15 = reg_0612;
    58: op1_15_in15 = reg_0994;
    59: op1_15_in15 = reg_0838;
    75: op1_15_in15 = reg_0838;
    60: op1_15_in15 = imem06_in[63:60];
    62: op1_15_in15 = imem01_in[43:40];
    63: op1_15_in15 = reg_0311;
    64: op1_15_in15 = imem04_in[11:8];
    65: op1_15_in15 = reg_0048;
    66: op1_15_in15 = reg_0806;
    67: op1_15_in15 = reg_0050;
    68: op1_15_in15 = reg_0475;
    69: op1_15_in15 = reg_0867;
    70: op1_15_in15 = reg_0151;
    71: op1_15_in15 = imem01_in[111:108];
    72: op1_15_in15 = reg_0537;
    73: op1_15_in15 = reg_0946;
    74: op1_15_in15 = reg_0384;
    77: op1_15_in15 = imem02_in[123:120];
    78: op1_15_in15 = reg_1005;
    79: op1_15_in15 = reg_0313;
    80: op1_15_in15 = reg_0834;
    81: op1_15_in15 = reg_0716;
    82: op1_15_in15 = reg_0281;
    83: op1_15_in15 = reg_1053;
    84: op1_15_in15 = reg_0604;
    85: op1_15_in15 = reg_0945;
    86: op1_15_in15 = imem05_in[99:96];
    87: op1_15_in15 = reg_0483;
    88: op1_15_in15 = reg_0706;
    89: op1_15_in15 = imem03_in[43:40];
    90: op1_15_in15 = reg_0015;
    91: op1_15_in15 = reg_0076;
    92: op1_15_in15 = imem01_in[15:12];
    93: op1_15_in15 = reg_0451;
    94: op1_15_in15 = reg_0456;
    default: op1_15_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_15_inv15 = 1;
    12: op1_15_inv15 = 1;
    13: op1_15_inv15 = 1;
    15: op1_15_inv15 = 1;
    16: op1_15_inv15 = 1;
    18: op1_15_inv15 = 1;
    19: op1_15_inv15 = 1;
    21: op1_15_inv15 = 1;
    23: op1_15_inv15 = 1;
    25: op1_15_inv15 = 1;
    26: op1_15_inv15 = 1;
    29: op1_15_inv15 = 1;
    31: op1_15_inv15 = 1;
    33: op1_15_inv15 = 1;
    34: op1_15_inv15 = 1;
    36: op1_15_inv15 = 1;
    38: op1_15_inv15 = 1;
    40: op1_15_inv15 = 1;
    45: op1_15_inv15 = 1;
    51: op1_15_inv15 = 1;
    52: op1_15_inv15 = 1;
    53: op1_15_inv15 = 1;
    54: op1_15_inv15 = 1;
    55: op1_15_inv15 = 1;
    56: op1_15_inv15 = 1;
    57: op1_15_inv15 = 1;
    58: op1_15_inv15 = 1;
    59: op1_15_inv15 = 1;
    63: op1_15_inv15 = 1;
    64: op1_15_inv15 = 1;
    67: op1_15_inv15 = 1;
    68: op1_15_inv15 = 1;
    70: op1_15_inv15 = 1;
    71: op1_15_inv15 = 1;
    73: op1_15_inv15 = 1;
    74: op1_15_inv15 = 1;
    77: op1_15_inv15 = 1;
    78: op1_15_inv15 = 1;
    79: op1_15_inv15 = 1;
    81: op1_15_inv15 = 1;
    83: op1_15_inv15 = 1;
    88: op1_15_inv15 = 1;
    91: op1_15_inv15 = 1;
    default: op1_15_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in16 = imem03_in[3:0];
    7: op1_15_in16 = reg_0396;
    8: op1_15_in16 = reg_0138;
    9: op1_15_in16 = reg_0520;
    10: op1_15_in16 = reg_0208;
    11: op1_15_in16 = imem05_in[63:60];
    12: op1_15_in16 = reg_0406;
    13: op1_15_in16 = reg_0534;
    14: op1_15_in16 = reg_0609;
    15: op1_15_in16 = reg_0706;
    16: op1_15_in16 = reg_0652;
    17: op1_15_in16 = reg_0535;
    18: op1_15_in16 = reg_0595;
    19: op1_15_in16 = imem04_in[7:4];
    20: op1_15_in16 = imem02_in[55:52];
    21: op1_15_in16 = reg_0827;
    22: op1_15_in16 = reg_0446;
    23: op1_15_in16 = reg_0327;
    24: op1_15_in16 = reg_0191;
    25: op1_15_in16 = reg_0117;
    26: op1_15_in16 = reg_0781;
    27: op1_15_in16 = imem03_in[95:92];
    28: op1_15_in16 = reg_0145;
    29: op1_15_in16 = reg_0166;
    30: op1_15_in16 = reg_0916;
    31: op1_15_in16 = imem06_in[15:12];
    32: op1_15_in16 = imem06_in[35:32];
    34: op1_15_in16 = imem05_in[87:84];
    35: op1_15_in16 = reg_0252;
    36: op1_15_in16 = reg_0805;
    38: op1_15_in16 = reg_0711;
    39: op1_15_in16 = reg_0201;
    40: op1_15_in16 = reg_0187;
    41: op1_15_in16 = reg_0997;
    42: op1_15_in16 = imem07_in[27:24];
    44: op1_15_in16 = reg_1039;
    45: op1_15_in16 = imem04_in[51:48];
    46: op1_15_in16 = imem07_in[115:112];
    47: op1_15_in16 = reg_0456;
    48: op1_15_in16 = imem04_in[71:68];
    49: op1_15_in16 = imem05_in[115:112];
    50: op1_15_in16 = reg_0576;
    51: op1_15_in16 = reg_0119;
    52: op1_15_in16 = imem01_in[71:68];
    53: op1_15_in16 = reg_0565;
    54: op1_15_in16 = reg_0326;
    55: op1_15_in16 = reg_0302;
    56: op1_15_in16 = imem06_in[51:48];
    57: op1_15_in16 = reg_0093;
    58: op1_15_in16 = imem04_in[31:28];
    59: op1_15_in16 = reg_0164;
    60: op1_15_in16 = imem06_in[79:76];
    62: op1_15_in16 = imem01_in[47:44];
    63: op1_15_in16 = reg_0369;
    64: op1_15_in16 = imem04_in[35:32];
    65: op1_15_in16 = reg_0568;
    66: op1_15_in16 = reg_0655;
    67: op1_15_in16 = reg_0541;
    68: op1_15_in16 = reg_0462;
    69: op1_15_in16 = reg_0506;
    70: op1_15_in16 = reg_0139;
    71: op1_15_in16 = imem01_in[115:112];
    72: op1_15_in16 = reg_0909;
    73: op1_15_in16 = reg_0952;
    74: op1_15_in16 = reg_0297;
    75: op1_15_in16 = reg_0175;
    77: op1_15_in16 = reg_0844;
    78: op1_15_in16 = reg_0276;
    79: op1_15_in16 = reg_0507;
    80: op1_15_in16 = reg_0022;
    81: op1_15_in16 = reg_0677;
    82: op1_15_in16 = reg_0040;
    83: op1_15_in16 = reg_0555;
    84: op1_15_in16 = reg_1040;
    85: op1_15_in16 = reg_0490;
    86: op1_15_in16 = imem05_in[111:108];
    87: op1_15_in16 = reg_0621;
    88: op1_15_in16 = reg_0951;
    89: op1_15_in16 = imem03_in[115:112];
    90: op1_15_in16 = reg_0064;
    91: op1_15_in16 = reg_0401;
    92: op1_15_in16 = imem01_in[51:48];
    93: op1_15_in16 = reg_0476;
    94: op1_15_in16 = reg_0200;
    default: op1_15_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_15_inv16 = 1;
    12: op1_15_inv16 = 1;
    15: op1_15_inv16 = 1;
    16: op1_15_inv16 = 1;
    21: op1_15_inv16 = 1;
    22: op1_15_inv16 = 1;
    23: op1_15_inv16 = 1;
    24: op1_15_inv16 = 1;
    25: op1_15_inv16 = 1;
    26: op1_15_inv16 = 1;
    27: op1_15_inv16 = 1;
    29: op1_15_inv16 = 1;
    31: op1_15_inv16 = 1;
    34: op1_15_inv16 = 1;
    38: op1_15_inv16 = 1;
    40: op1_15_inv16 = 1;
    45: op1_15_inv16 = 1;
    46: op1_15_inv16 = 1;
    48: op1_15_inv16 = 1;
    49: op1_15_inv16 = 1;
    56: op1_15_inv16 = 1;
    57: op1_15_inv16 = 1;
    60: op1_15_inv16 = 1;
    64: op1_15_inv16 = 1;
    65: op1_15_inv16 = 1;
    67: op1_15_inv16 = 1;
    71: op1_15_inv16 = 1;
    72: op1_15_inv16 = 1;
    78: op1_15_inv16 = 1;
    82: op1_15_inv16 = 1;
    85: op1_15_inv16 = 1;
    86: op1_15_inv16 = 1;
    88: op1_15_inv16 = 1;
    91: op1_15_inv16 = 1;
    default: op1_15_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in17 = imem03_in[87:84];
    7: op1_15_in17 = reg_0374;
    8: op1_15_in17 = reg_0130;
    9: op1_15_in17 = reg_0509;
    10: op1_15_in17 = reg_0204;
    11: op1_15_in17 = imem05_in[75:72];
    12: op1_15_in17 = reg_0799;
    13: op1_15_in17 = reg_0535;
    14: op1_15_in17 = reg_0619;
    15: op1_15_in17 = reg_0423;
    16: op1_15_in17 = reg_0333;
    17: op1_15_in17 = reg_0532;
    18: op1_15_in17 = reg_0394;
    19: op1_15_in17 = imem04_in[15:12];
    20: op1_15_in17 = imem02_in[75:72];
    21: op1_15_in17 = reg_0757;
    22: op1_15_in17 = reg_0443;
    23: op1_15_in17 = reg_0322;
    24: op1_15_in17 = reg_0210;
    25: op1_15_in17 = reg_0121;
    26: op1_15_in17 = reg_1010;
    27: op1_15_in17 = imem03_in[111:108];
    28: op1_15_in17 = reg_0135;
    29: op1_15_in17 = reg_0164;
    30: op1_15_in17 = reg_0081;
    31: op1_15_in17 = imem06_in[23:20];
    32: op1_15_in17 = imem07_in[27:24];
    34: op1_15_in17 = imem05_in[103:100];
    35: op1_15_in17 = reg_0813;
    36: op1_15_in17 = reg_0735;
    38: op1_15_in17 = reg_0422;
    39: op1_15_in17 = reg_0212;
    40: op1_15_in17 = reg_0198;
    41: op1_15_in17 = imem04_in[47:44];
    42: op1_15_in17 = imem07_in[35:32];
    44: op1_15_in17 = reg_0496;
    45: op1_15_in17 = imem04_in[59:56];
    46: op1_15_in17 = reg_0728;
    47: op1_15_in17 = reg_0458;
    48: op1_15_in17 = imem04_in[83:80];
    49: op1_15_in17 = imem05_in[123:120];
    50: op1_15_in17 = reg_0874;
    51: op1_15_in17 = reg_0112;
    52: op1_15_in17 = imem01_in[111:108];
    53: op1_15_in17 = reg_0365;
    54: op1_15_in17 = reg_0656;
    55: op1_15_in17 = reg_0808;
    91: op1_15_in17 = reg_0808;
    56: op1_15_in17 = imem06_in[83:80];
    57: op1_15_in17 = reg_0673;
    58: op1_15_in17 = imem04_in[39:36];
    59: op1_15_in17 = reg_0173;
    60: op1_15_in17 = imem06_in[87:84];
    62: op1_15_in17 = reg_0786;
    63: op1_15_in17 = reg_0807;
    64: op1_15_in17 = imem04_in[43:40];
    65: op1_15_in17 = reg_0076;
    66: op1_15_in17 = reg_0689;
    67: op1_15_in17 = reg_0064;
    68: op1_15_in17 = reg_0472;
    69: op1_15_in17 = reg_0884;
    70: op1_15_in17 = reg_0138;
    71: op1_15_in17 = reg_0488;
    72: op1_15_in17 = reg_0524;
    73: op1_15_in17 = reg_0943;
    74: op1_15_in17 = reg_0895;
    75: op1_15_in17 = reg_0167;
    77: op1_15_in17 = reg_0916;
    78: op1_15_in17 = reg_0288;
    90: op1_15_in17 = reg_0288;
    79: op1_15_in17 = reg_0909;
    80: op1_15_in17 = imem07_in[3:0];
    81: op1_15_in17 = reg_0678;
    82: op1_15_in17 = reg_0609;
    83: op1_15_in17 = reg_0860;
    84: op1_15_in17 = reg_0116;
    85: op1_15_in17 = reg_0144;
    86: op1_15_in17 = reg_0866;
    87: op1_15_in17 = reg_0073;
    88: op1_15_in17 = imem06_in[7:4];
    89: op1_15_in17 = imem03_in[123:120];
    92: op1_15_in17 = imem01_in[55:52];
    93: op1_15_in17 = reg_0460;
    94: op1_15_in17 = reg_0205;
    default: op1_15_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv17 = 1;
    8: op1_15_inv17 = 1;
    9: op1_15_inv17 = 1;
    10: op1_15_inv17 = 1;
    11: op1_15_inv17 = 1;
    16: op1_15_inv17 = 1;
    17: op1_15_inv17 = 1;
    19: op1_15_inv17 = 1;
    22: op1_15_inv17 = 1;
    23: op1_15_inv17 = 1;
    25: op1_15_inv17 = 1;
    27: op1_15_inv17 = 1;
    31: op1_15_inv17 = 1;
    34: op1_15_inv17 = 1;
    39: op1_15_inv17 = 1;
    40: op1_15_inv17 = 1;
    42: op1_15_inv17 = 1;
    45: op1_15_inv17 = 1;
    48: op1_15_inv17 = 1;
    51: op1_15_inv17 = 1;
    52: op1_15_inv17 = 1;
    54: op1_15_inv17 = 1;
    55: op1_15_inv17 = 1;
    56: op1_15_inv17 = 1;
    59: op1_15_inv17 = 1;
    60: op1_15_inv17 = 1;
    63: op1_15_inv17 = 1;
    66: op1_15_inv17 = 1;
    67: op1_15_inv17 = 1;
    70: op1_15_inv17 = 1;
    73: op1_15_inv17 = 1;
    77: op1_15_inv17 = 1;
    78: op1_15_inv17 = 1;
    79: op1_15_inv17 = 1;
    80: op1_15_inv17 = 1;
    81: op1_15_inv17 = 1;
    82: op1_15_inv17 = 1;
    84: op1_15_inv17 = 1;
    85: op1_15_inv17 = 1;
    87: op1_15_inv17 = 1;
    88: op1_15_inv17 = 1;
    89: op1_15_inv17 = 1;
    90: op1_15_inv17 = 1;
    91: op1_15_inv17 = 1;
    92: op1_15_inv17 = 1;
    94: op1_15_inv17 = 1;
    default: op1_15_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in18 = imem03_in[119:116];
    7: op1_15_in18 = reg_0987;
    8: op1_15_in18 = reg_0155;
    9: op1_15_in18 = reg_0502;
    10: op1_15_in18 = reg_0193;
    11: op1_15_in18 = imem05_in[111:108];
    12: op1_15_in18 = reg_0800;
    13: op1_15_in18 = reg_0549;
    14: op1_15_in18 = reg_0633;
    15: op1_15_in18 = reg_0162;
    16: op1_15_in18 = reg_0088;
    17: op1_15_in18 = reg_0551;
    18: op1_15_in18 = reg_0395;
    19: op1_15_in18 = imem04_in[31:28];
    20: op1_15_in18 = imem02_in[115:112];
    21: op1_15_in18 = reg_0252;
    22: op1_15_in18 = reg_0420;
    23: op1_15_in18 = reg_0389;
    24: op1_15_in18 = reg_0187;
    25: op1_15_in18 = imem02_in[15:12];
    26: op1_15_in18 = reg_1011;
    27: op1_15_in18 = reg_0599;
    28: op1_15_in18 = reg_0136;
    30: op1_15_in18 = reg_0225;
    31: op1_15_in18 = imem06_in[63:60];
    32: op1_15_in18 = imem07_in[95:92];
    34: op1_15_in18 = imem05_in[123:120];
    35: op1_15_in18 = reg_0275;
    36: op1_15_in18 = reg_0615;
    38: op1_15_in18 = reg_0447;
    39: op1_15_in18 = reg_0205;
    40: op1_15_in18 = reg_0190;
    41: op1_15_in18 = imem04_in[79:76];
    42: op1_15_in18 = imem07_in[43:40];
    44: op1_15_in18 = reg_1043;
    45: op1_15_in18 = imem04_in[63:60];
    46: op1_15_in18 = reg_0321;
    47: op1_15_in18 = reg_0188;
    48: op1_15_in18 = imem04_in[91:88];
    49: op1_15_in18 = reg_0955;
    50: op1_15_in18 = reg_0051;
    82: op1_15_in18 = reg_0051;
    51: op1_15_in18 = reg_0114;
    52: op1_15_in18 = imem01_in[123:120];
    53: op1_15_in18 = reg_0739;
    54: op1_15_in18 = reg_0621;
    55: op1_15_in18 = reg_0074;
    56: op1_15_in18 = imem06_in[111:108];
    57: op1_15_in18 = reg_0597;
    58: op1_15_in18 = imem04_in[59:56];
    59: op1_15_in18 = reg_0184;
    60: op1_15_in18 = imem06_in[115:112];
    62: op1_15_in18 = reg_0223;
    63: op1_15_in18 = reg_0820;
    64: op1_15_in18 = imem04_in[55:52];
    65: op1_15_in18 = reg_0014;
    66: op1_15_in18 = reg_0266;
    67: op1_15_in18 = reg_0809;
    68: op1_15_in18 = reg_0474;
    69: op1_15_in18 = imem03_in[7:4];
    70: op1_15_in18 = imem06_in[39:36];
    88: op1_15_in18 = imem06_in[39:36];
    71: op1_15_in18 = reg_0234;
    72: op1_15_in18 = reg_0066;
    73: op1_15_in18 = reg_0953;
    74: op1_15_in18 = reg_0556;
    75: op1_15_in18 = reg_0183;
    77: op1_15_in18 = reg_0803;
    78: op1_15_in18 = reg_0658;
    79: op1_15_in18 = reg_0068;
    80: op1_15_in18 = imem07_in[19:16];
    81: op1_15_in18 = reg_0167;
    83: op1_15_in18 = reg_0827;
    84: op1_15_in18 = reg_0761;
    85: op1_15_in18 = imem06_in[23:20];
    86: op1_15_in18 = reg_0142;
    87: op1_15_in18 = reg_0358;
    89: op1_15_in18 = imem03_in[127:124];
    90: op1_15_in18 = reg_0284;
    91: op1_15_in18 = reg_0432;
    92: op1_15_in18 = imem01_in[71:68];
    93: op1_15_in18 = reg_0481;
    94: op1_15_in18 = reg_0607;
    default: op1_15_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_15_inv18 = 1;
    10: op1_15_inv18 = 1;
    12: op1_15_inv18 = 1;
    13: op1_15_inv18 = 1;
    15: op1_15_inv18 = 1;
    16: op1_15_inv18 = 1;
    20: op1_15_inv18 = 1;
    22: op1_15_inv18 = 1;
    23: op1_15_inv18 = 1;
    27: op1_15_inv18 = 1;
    28: op1_15_inv18 = 1;
    30: op1_15_inv18 = 1;
    34: op1_15_inv18 = 1;
    38: op1_15_inv18 = 1;
    41: op1_15_inv18 = 1;
    42: op1_15_inv18 = 1;
    44: op1_15_inv18 = 1;
    45: op1_15_inv18 = 1;
    46: op1_15_inv18 = 1;
    47: op1_15_inv18 = 1;
    49: op1_15_inv18 = 1;
    51: op1_15_inv18 = 1;
    52: op1_15_inv18 = 1;
    53: op1_15_inv18 = 1;
    55: op1_15_inv18 = 1;
    62: op1_15_inv18 = 1;
    63: op1_15_inv18 = 1;
    65: op1_15_inv18 = 1;
    66: op1_15_inv18 = 1;
    67: op1_15_inv18 = 1;
    69: op1_15_inv18 = 1;
    71: op1_15_inv18 = 1;
    72: op1_15_inv18 = 1;
    73: op1_15_inv18 = 1;
    75: op1_15_inv18 = 1;
    80: op1_15_inv18 = 1;
    83: op1_15_inv18 = 1;
    84: op1_15_inv18 = 1;
    91: op1_15_inv18 = 1;
    92: op1_15_inv18 = 1;
    94: op1_15_inv18 = 1;
    default: op1_15_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in19 = reg_0579;
    7: op1_15_in19 = reg_0982;
    8: op1_15_in19 = imem06_in[23:20];
    9: op1_15_in19 = reg_0524;
    10: op1_15_in19 = reg_0213;
    11: op1_15_in19 = imem05_in[115:112];
    12: op1_15_in19 = reg_0808;
    65: op1_15_in19 = reg_0808;
    13: op1_15_in19 = reg_0532;
    14: op1_15_in19 = reg_0349;
    16: op1_15_in19 = reg_0089;
    17: op1_15_in19 = reg_0531;
    18: op1_15_in19 = reg_0387;
    19: op1_15_in19 = imem04_in[59:56];
    20: op1_15_in19 = reg_0645;
    21: op1_15_in19 = reg_0813;
    22: op1_15_in19 = reg_0175;
    23: op1_15_in19 = reg_0998;
    50: op1_15_in19 = reg_0998;
    24: op1_15_in19 = reg_0193;
    25: op1_15_in19 = imem02_in[31:28];
    26: op1_15_in19 = reg_0754;
    27: op1_15_in19 = reg_0583;
    28: op1_15_in19 = reg_0138;
    30: op1_15_in19 = reg_0082;
    31: op1_15_in19 = reg_0610;
    32: op1_15_in19 = reg_0720;
    34: op1_15_in19 = reg_0944;
    35: op1_15_in19 = reg_0825;
    36: op1_15_in19 = imem06_in[7:4];
    38: op1_15_in19 = reg_0439;
    39: op1_15_in19 = reg_0190;
    40: op1_15_in19 = reg_0905;
    41: op1_15_in19 = imem04_in[87:84];
    42: op1_15_in19 = imem07_in[47:44];
    44: op1_15_in19 = reg_0829;
    45: op1_15_in19 = imem04_in[107:104];
    46: op1_15_in19 = reg_0744;
    47: op1_15_in19 = reg_0207;
    48: op1_15_in19 = reg_0530;
    58: op1_15_in19 = reg_0530;
    49: op1_15_in19 = reg_0954;
    51: op1_15_in19 = reg_0109;
    52: op1_15_in19 = reg_1044;
    53: op1_15_in19 = reg_0424;
    54: op1_15_in19 = reg_0652;
    55: op1_15_in19 = reg_0893;
    56: op1_15_in19 = reg_0759;
    57: op1_15_in19 = reg_0566;
    60: op1_15_in19 = reg_0010;
    62: op1_15_in19 = reg_1036;
    63: op1_15_in19 = reg_0518;
    64: op1_15_in19 = imem04_in[83:80];
    66: op1_15_in19 = reg_0022;
    67: op1_15_in19 = reg_0243;
    68: op1_15_in19 = reg_0479;
    69: op1_15_in19 = imem03_in[19:16];
    70: op1_15_in19 = imem06_in[115:112];
    71: op1_15_in19 = reg_1024;
    72: op1_15_in19 = reg_0302;
    73: op1_15_in19 = reg_0734;
    74: op1_15_in19 = reg_0382;
    77: op1_15_in19 = reg_0846;
    78: op1_15_in19 = reg_0065;
    79: op1_15_in19 = reg_0401;
    80: op1_15_in19 = imem07_in[91:88];
    81: op1_15_in19 = reg_0757;
    82: op1_15_in19 = reg_0385;
    83: op1_15_in19 = reg_0101;
    84: op1_15_in19 = reg_0290;
    85: op1_15_in19 = imem06_in[39:36];
    86: op1_15_in19 = reg_0647;
    87: op1_15_in19 = reg_0052;
    88: op1_15_in19 = imem06_in[71:68];
    89: op1_15_in19 = reg_0307;
    90: op1_15_in19 = reg_0764;
    91: op1_15_in19 = reg_0444;
    92: op1_15_in19 = imem01_in[103:100];
    93: op1_15_in19 = reg_0467;
    94: op1_15_in19 = reg_0369;
    default: op1_15_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv19 = 1;
    8: op1_15_inv19 = 1;
    10: op1_15_inv19 = 1;
    11: op1_15_inv19 = 1;
    12: op1_15_inv19 = 1;
    13: op1_15_inv19 = 1;
    16: op1_15_inv19 = 1;
    18: op1_15_inv19 = 1;
    21: op1_15_inv19 = 1;
    22: op1_15_inv19 = 1;
    24: op1_15_inv19 = 1;
    27: op1_15_inv19 = 1;
    28: op1_15_inv19 = 1;
    30: op1_15_inv19 = 1;
    34: op1_15_inv19 = 1;
    35: op1_15_inv19 = 1;
    36: op1_15_inv19 = 1;
    38: op1_15_inv19 = 1;
    39: op1_15_inv19 = 1;
    40: op1_15_inv19 = 1;
    42: op1_15_inv19 = 1;
    45: op1_15_inv19 = 1;
    46: op1_15_inv19 = 1;
    50: op1_15_inv19 = 1;
    53: op1_15_inv19 = 1;
    54: op1_15_inv19 = 1;
    56: op1_15_inv19 = 1;
    57: op1_15_inv19 = 1;
    58: op1_15_inv19 = 1;
    60: op1_15_inv19 = 1;
    62: op1_15_inv19 = 1;
    63: op1_15_inv19 = 1;
    64: op1_15_inv19 = 1;
    65: op1_15_inv19 = 1;
    67: op1_15_inv19 = 1;
    70: op1_15_inv19 = 1;
    72: op1_15_inv19 = 1;
    74: op1_15_inv19 = 1;
    77: op1_15_inv19 = 1;
    80: op1_15_inv19 = 1;
    81: op1_15_inv19 = 1;
    86: op1_15_inv19 = 1;
    87: op1_15_inv19 = 1;
    91: op1_15_inv19 = 1;
    92: op1_15_inv19 = 1;
    93: op1_15_inv19 = 1;
    default: op1_15_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in20 = reg_0589;
    7: op1_15_in20 = reg_0996;
    8: op1_15_in20 = imem06_in[43:40];
    85: op1_15_in20 = imem06_in[43:40];
    9: op1_15_in20 = reg_0503;
    10: op1_15_in20 = reg_0190;
    11: op1_15_in20 = reg_0970;
    12: op1_15_in20 = reg_0486;
    13: op1_15_in20 = reg_0531;
    14: op1_15_in20 = reg_1029;
    16: op1_15_in20 = reg_0095;
    17: op1_15_in20 = reg_0541;
    18: op1_15_in20 = reg_0385;
    19: op1_15_in20 = imem04_in[67:64];
    20: op1_15_in20 = reg_0658;
    21: op1_15_in20 = reg_0257;
    22: op1_15_in20 = reg_0162;
    23: op1_15_in20 = reg_1001;
    24: op1_15_in20 = reg_0198;
    47: op1_15_in20 = reg_0198;
    25: op1_15_in20 = imem02_in[83:80];
    26: op1_15_in20 = imem07_in[3:0];
    27: op1_15_in20 = reg_0572;
    28: op1_15_in20 = reg_0141;
    30: op1_15_in20 = reg_0817;
    31: op1_15_in20 = reg_0620;
    32: op1_15_in20 = reg_0721;
    34: op1_15_in20 = reg_0959;
    35: op1_15_in20 = reg_0244;
    36: op1_15_in20 = imem06_in[35:32];
    38: op1_15_in20 = reg_0179;
    39: op1_15_in20 = imem01_in[51:48];
    40: op1_15_in20 = reg_1051;
    41: op1_15_in20 = reg_0511;
    42: op1_15_in20 = imem07_in[71:68];
    44: op1_15_in20 = reg_0521;
    45: op1_15_in20 = imem04_in[123:120];
    46: op1_15_in20 = reg_0428;
    48: op1_15_in20 = reg_0282;
    49: op1_15_in20 = reg_0969;
    50: op1_15_in20 = reg_1002;
    51: op1_15_in20 = reg_0117;
    52: op1_15_in20 = reg_0242;
    53: op1_15_in20 = reg_0394;
    54: op1_15_in20 = reg_0739;
    55: op1_15_in20 = reg_0899;
    56: op1_15_in20 = reg_0624;
    57: op1_15_in20 = imem06_in[31:28];
    58: op1_15_in20 = reg_1009;
    60: op1_15_in20 = reg_0025;
    62: op1_15_in20 = reg_0522;
    63: op1_15_in20 = reg_0987;
    64: op1_15_in20 = imem04_in[115:112];
    65: op1_15_in20 = reg_0815;
    66: op1_15_in20 = reg_0968;
    67: op1_15_in20 = reg_0444;
    68: op1_15_in20 = reg_0214;
    69: op1_15_in20 = imem03_in[23:20];
    70: op1_15_in20 = reg_0391;
    71: op1_15_in20 = reg_0225;
    72: op1_15_in20 = reg_0015;
    73: op1_15_in20 = imem05_in[39:36];
    74: op1_15_in20 = reg_0008;
    77: op1_15_in20 = reg_0082;
    78: op1_15_in20 = imem05_in[23:20];
    79: op1_15_in20 = reg_0288;
    80: op1_15_in20 = imem07_in[107:104];
    81: op1_15_in20 = reg_0127;
    82: op1_15_in20 = reg_0588;
    83: op1_15_in20 = reg_0115;
    84: op1_15_in20 = reg_0261;
    86: op1_15_in20 = reg_0143;
    87: op1_15_in20 = reg_0087;
    88: op1_15_in20 = imem06_in[103:100];
    89: op1_15_in20 = reg_0149;
    90: op1_15_in20 = reg_0432;
    91: op1_15_in20 = imem05_in[47:44];
    92: op1_15_in20 = imem01_in[119:116];
    93: op1_15_in20 = reg_0470;
    94: op1_15_in20 = reg_0849;
    default: op1_15_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv20 = 1;
    11: op1_15_inv20 = 1;
    17: op1_15_inv20 = 1;
    18: op1_15_inv20 = 1;
    20: op1_15_inv20 = 1;
    21: op1_15_inv20 = 1;
    25: op1_15_inv20 = 1;
    26: op1_15_inv20 = 1;
    27: op1_15_inv20 = 1;
    28: op1_15_inv20 = 1;
    31: op1_15_inv20 = 1;
    32: op1_15_inv20 = 1;
    34: op1_15_inv20 = 1;
    35: op1_15_inv20 = 1;
    38: op1_15_inv20 = 1;
    40: op1_15_inv20 = 1;
    41: op1_15_inv20 = 1;
    42: op1_15_inv20 = 1;
    44: op1_15_inv20 = 1;
    46: op1_15_inv20 = 1;
    48: op1_15_inv20 = 1;
    50: op1_15_inv20 = 1;
    51: op1_15_inv20 = 1;
    53: op1_15_inv20 = 1;
    55: op1_15_inv20 = 1;
    56: op1_15_inv20 = 1;
    57: op1_15_inv20 = 1;
    58: op1_15_inv20 = 1;
    62: op1_15_inv20 = 1;
    63: op1_15_inv20 = 1;
    64: op1_15_inv20 = 1;
    65: op1_15_inv20 = 1;
    67: op1_15_inv20 = 1;
    68: op1_15_inv20 = 1;
    69: op1_15_inv20 = 1;
    72: op1_15_inv20 = 1;
    74: op1_15_inv20 = 1;
    78: op1_15_inv20 = 1;
    80: op1_15_inv20 = 1;
    81: op1_15_inv20 = 1;
    83: op1_15_inv20 = 1;
    84: op1_15_inv20 = 1;
    86: op1_15_inv20 = 1;
    89: op1_15_inv20 = 1;
    90: op1_15_inv20 = 1;
    93: op1_15_inv20 = 1;
    default: op1_15_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in21 = reg_0576;
    7: op1_15_in21 = reg_0980;
    8: op1_15_in21 = imem06_in[91:88];
    9: op1_15_in21 = reg_0515;
    10: op1_15_in21 = reg_0195;
    11: op1_15_in21 = reg_0971;
    12: op1_15_in21 = reg_1010;
    13: op1_15_in21 = reg_0547;
    14: op1_15_in21 = reg_0808;
    16: op1_15_in21 = reg_0085;
    17: op1_15_in21 = reg_0305;
    18: op1_15_in21 = reg_0396;
    19: op1_15_in21 = reg_0854;
    20: op1_15_in21 = reg_0637;
    21: op1_15_in21 = reg_0896;
    22: op1_15_in21 = reg_0170;
    23: op1_15_in21 = reg_0994;
    24: op1_15_in21 = reg_0190;
    25: op1_15_in21 = imem02_in[87:84];
    26: op1_15_in21 = imem07_in[39:36];
    27: op1_15_in21 = reg_0592;
    28: op1_15_in21 = reg_0155;
    30: op1_15_in21 = reg_0037;
    31: op1_15_in21 = reg_0626;
    32: op1_15_in21 = reg_0726;
    34: op1_15_in21 = reg_0949;
    35: op1_15_in21 = reg_1046;
    36: op1_15_in21 = imem06_in[47:44];
    85: op1_15_in21 = imem06_in[47:44];
    38: op1_15_in21 = reg_0161;
    39: op1_15_in21 = imem01_in[115:112];
    40: op1_15_in21 = reg_0276;
    41: op1_15_in21 = reg_0282;
    42: op1_15_in21 = imem07_in[119:116];
    44: op1_15_in21 = reg_0122;
    45: op1_15_in21 = reg_0265;
    46: op1_15_in21 = reg_0350;
    47: op1_15_in21 = reg_0205;
    48: op1_15_in21 = reg_0539;
    49: op1_15_in21 = reg_0964;
    50: op1_15_in21 = reg_0992;
    51: op1_15_in21 = reg_0110;
    83: op1_15_in21 = reg_0110;
    52: op1_15_in21 = reg_1035;
    53: op1_15_in21 = reg_0368;
    54: op1_15_in21 = reg_0329;
    55: op1_15_in21 = reg_0529;
    56: op1_15_in21 = reg_0556;
    57: op1_15_in21 = imem06_in[39:36];
    58: op1_15_in21 = reg_0912;
    60: op1_15_in21 = reg_0028;
    62: op1_15_in21 = reg_1043;
    63: op1_15_in21 = reg_0996;
    64: op1_15_in21 = reg_0536;
    65: op1_15_in21 = reg_0809;
    66: op1_15_in21 = imem05_in[11:8];
    67: op1_15_in21 = reg_0065;
    68: op1_15_in21 = reg_0200;
    69: op1_15_in21 = imem03_in[35:32];
    70: op1_15_in21 = reg_0025;
    71: op1_15_in21 = reg_0607;
    72: op1_15_in21 = reg_0296;
    73: op1_15_in21 = imem05_in[51:48];
    74: op1_15_in21 = reg_0026;
    77: op1_15_in21 = reg_0887;
    78: op1_15_in21 = imem05_in[99:96];
    79: op1_15_in21 = reg_0284;
    80: op1_15_in21 = imem07_in[111:108];
    81: op1_15_in21 = reg_0436;
    82: op1_15_in21 = reg_0991;
    84: op1_15_in21 = imem02_in[7:4];
    86: op1_15_in21 = reg_0138;
    87: op1_15_in21 = reg_0608;
    88: op1_15_in21 = imem06_in[123:120];
    89: op1_15_in21 = reg_0346;
    90: op1_15_in21 = reg_0027;
    91: op1_15_in21 = imem05_in[111:108];
    92: op1_15_in21 = reg_1042;
    93: op1_15_in21 = reg_0479;
    94: op1_15_in21 = reg_0968;
    default: op1_15_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_15_inv21 = 1;
    10: op1_15_inv21 = 1;
    14: op1_15_inv21 = 1;
    18: op1_15_inv21 = 1;
    19: op1_15_inv21 = 1;
    21: op1_15_inv21 = 1;
    23: op1_15_inv21 = 1;
    24: op1_15_inv21 = 1;
    25: op1_15_inv21 = 1;
    27: op1_15_inv21 = 1;
    28: op1_15_inv21 = 1;
    30: op1_15_inv21 = 1;
    32: op1_15_inv21 = 1;
    36: op1_15_inv21 = 1;
    39: op1_15_inv21 = 1;
    41: op1_15_inv21 = 1;
    42: op1_15_inv21 = 1;
    44: op1_15_inv21 = 1;
    46: op1_15_inv21 = 1;
    47: op1_15_inv21 = 1;
    48: op1_15_inv21 = 1;
    50: op1_15_inv21 = 1;
    55: op1_15_inv21 = 1;
    56: op1_15_inv21 = 1;
    58: op1_15_inv21 = 1;
    60: op1_15_inv21 = 1;
    66: op1_15_inv21 = 1;
    67: op1_15_inv21 = 1;
    68: op1_15_inv21 = 1;
    73: op1_15_inv21 = 1;
    77: op1_15_inv21 = 1;
    79: op1_15_inv21 = 1;
    82: op1_15_inv21 = 1;
    84: op1_15_inv21 = 1;
    87: op1_15_inv21 = 1;
    90: op1_15_inv21 = 1;
    92: op1_15_inv21 = 1;
    default: op1_15_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in22 = reg_0384;
    7: op1_15_in22 = reg_0988;
    8: op1_15_in22 = imem06_in[95:92];
    9: op1_15_in22 = reg_0232;
    10: op1_15_in22 = reg_0772;
    11: op1_15_in22 = reg_0957;
    12: op1_15_in22 = reg_1011;
    13: op1_15_in22 = reg_0292;
    14: op1_15_in22 = reg_0780;
    16: op1_15_in22 = reg_0052;
    17: op1_15_in22 = reg_0300;
    18: op1_15_in22 = reg_0309;
    19: op1_15_in22 = reg_0875;
    20: op1_15_in22 = reg_0646;
    21: op1_15_in22 = reg_0145;
    23: op1_15_in22 = imem04_in[59:56];
    24: op1_15_in22 = reg_0206;
    25: op1_15_in22 = imem02_in[115:112];
    26: op1_15_in22 = reg_0730;
    27: op1_15_in22 = reg_0591;
    28: op1_15_in22 = imem06_in[27:24];
    30: op1_15_in22 = reg_0093;
    31: op1_15_in22 = reg_0633;
    32: op1_15_in22 = reg_0715;
    34: op1_15_in22 = reg_0821;
    35: op1_15_in22 = reg_0831;
    36: op1_15_in22 = imem06_in[111:108];
    38: op1_15_in22 = reg_0168;
    39: op1_15_in22 = reg_0013;
    40: op1_15_in22 = reg_1034;
    52: op1_15_in22 = reg_1034;
    41: op1_15_in22 = reg_0055;
    58: op1_15_in22 = reg_0055;
    42: op1_15_in22 = imem07_in[127:124];
    80: op1_15_in22 = imem07_in[127:124];
    44: op1_15_in22 = reg_0099;
    45: op1_15_in22 = reg_0277;
    46: op1_15_in22 = reg_0431;
    47: op1_15_in22 = reg_0192;
    48: op1_15_in22 = reg_0931;
    49: op1_15_in22 = reg_0945;
    50: op1_15_in22 = reg_0995;
    51: op1_15_in22 = imem02_in[51:48];
    53: op1_15_in22 = reg_0876;
    54: op1_15_in22 = reg_0389;
    55: op1_15_in22 = reg_0053;
    56: op1_15_in22 = reg_0619;
    57: op1_15_in22 = imem06_in[47:44];
    60: op1_15_in22 = reg_0297;
    62: op1_15_in22 = reg_0500;
    63: op1_15_in22 = reg_0993;
    64: op1_15_in22 = reg_0511;
    65: op1_15_in22 = reg_0444;
    66: op1_15_in22 = imem05_in[55:52];
    67: op1_15_in22 = reg_0494;
    68: op1_15_in22 = reg_0193;
    69: op1_15_in22 = imem03_in[47:44];
    70: op1_15_in22 = reg_0679;
    71: op1_15_in22 = reg_0829;
    72: op1_15_in22 = reg_0072;
    73: op1_15_in22 = imem05_in[67:64];
    74: op1_15_in22 = reg_0370;
    77: op1_15_in22 = reg_0645;
    78: op1_15_in22 = imem05_in[115:112];
    79: op1_15_in22 = reg_0065;
    81: op1_15_in22 = reg_0000;
    82: op1_15_in22 = reg_0984;
    83: op1_15_in22 = imem02_in[43:40];
    84: op1_15_in22 = imem02_in[59:56];
    85: op1_15_in22 = imem06_in[115:112];
    86: op1_15_in22 = reg_0140;
    87: op1_15_in22 = reg_0347;
    88: op1_15_in22 = reg_0010;
    89: op1_15_in22 = reg_0342;
    90: op1_15_in22 = reg_0495;
    91: op1_15_in22 = reg_0268;
    92: op1_15_in22 = reg_0246;
    93: op1_15_in22 = reg_0459;
    94: op1_15_in22 = reg_0240;
    default: op1_15_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv22 = 1;
    10: op1_15_inv22 = 1;
    11: op1_15_inv22 = 1;
    14: op1_15_inv22 = 1;
    16: op1_15_inv22 = 1;
    19: op1_15_inv22 = 1;
    20: op1_15_inv22 = 1;
    23: op1_15_inv22 = 1;
    24: op1_15_inv22 = 1;
    25: op1_15_inv22 = 1;
    30: op1_15_inv22 = 1;
    34: op1_15_inv22 = 1;
    42: op1_15_inv22 = 1;
    45: op1_15_inv22 = 1;
    46: op1_15_inv22 = 1;
    48: op1_15_inv22 = 1;
    50: op1_15_inv22 = 1;
    55: op1_15_inv22 = 1;
    56: op1_15_inv22 = 1;
    58: op1_15_inv22 = 1;
    62: op1_15_inv22 = 1;
    63: op1_15_inv22 = 1;
    64: op1_15_inv22 = 1;
    65: op1_15_inv22 = 1;
    68: op1_15_inv22 = 1;
    69: op1_15_inv22 = 1;
    70: op1_15_inv22 = 1;
    73: op1_15_inv22 = 1;
    77: op1_15_inv22 = 1;
    78: op1_15_inv22 = 1;
    79: op1_15_inv22 = 1;
    82: op1_15_inv22 = 1;
    85: op1_15_inv22 = 1;
    87: op1_15_inv22 = 1;
    88: op1_15_inv22 = 1;
    89: op1_15_inv22 = 1;
    94: op1_15_inv22 = 1;
    default: op1_15_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in23 = reg_0343;
    7: op1_15_in23 = reg_0976;
    8: op1_15_in23 = reg_0628;
    9: op1_15_in23 = reg_0235;
    10: op1_15_in23 = reg_0778;
    11: op1_15_in23 = reg_0965;
    12: op1_15_in23 = reg_0783;
    13: op1_15_in23 = reg_0047;
    14: op1_15_in23 = reg_0805;
    16: op1_15_in23 = reg_0086;
    30: op1_15_in23 = reg_0086;
    17: op1_15_in23 = reg_0289;
    18: op1_15_in23 = reg_0389;
    19: op1_15_in23 = imem05_in[79:76];
    20: op1_15_in23 = reg_0657;
    21: op1_15_in23 = reg_0152;
    23: op1_15_in23 = imem04_in[63:60];
    24: op1_15_in23 = reg_0199;
    25: op1_15_in23 = reg_0650;
    87: op1_15_in23 = reg_0650;
    26: op1_15_in23 = reg_0721;
    27: op1_15_in23 = reg_0581;
    28: op1_15_in23 = imem06_in[103:100];
    31: op1_15_in23 = reg_0618;
    32: op1_15_in23 = reg_0707;
    34: op1_15_in23 = reg_0256;
    35: op1_15_in23 = reg_0129;
    36: op1_15_in23 = imem06_in[123:120];
    38: op1_15_in23 = reg_0184;
    39: op1_15_in23 = reg_0239;
    40: op1_15_in23 = reg_0013;
    41: op1_15_in23 = reg_1057;
    58: op1_15_in23 = reg_1057;
    42: op1_15_in23 = reg_0702;
    44: op1_15_in23 = reg_0106;
    45: op1_15_in23 = reg_0282;
    46: op1_15_in23 = reg_0167;
    47: op1_15_in23 = imem01_in[19:16];
    48: op1_15_in23 = reg_0524;
    49: op1_15_in23 = reg_0952;
    50: op1_15_in23 = reg_0979;
    51: op1_15_in23 = imem02_in[75:72];
    52: op1_15_in23 = reg_0501;
    53: op1_15_in23 = reg_0291;
    54: op1_15_in23 = reg_0248;
    55: op1_15_in23 = reg_0041;
    56: op1_15_in23 = reg_0914;
    57: op1_15_in23 = imem06_in[59:56];
    60: op1_15_in23 = reg_0392;
    62: op1_15_in23 = reg_0740;
    63: op1_15_in23 = reg_0994;
    64: op1_15_in23 = reg_0584;
    65: op1_15_in23 = reg_0251;
    67: op1_15_in23 = reg_0251;
    66: op1_15_in23 = imem05_in[59:56];
    68: op1_15_in23 = reg_0190;
    69: op1_15_in23 = imem03_in[111:108];
    70: op1_15_in23 = reg_0021;
    71: op1_15_in23 = reg_0514;
    72: op1_15_in23 = reg_0893;
    73: op1_15_in23 = reg_0221;
    74: op1_15_in23 = reg_0018;
    77: op1_15_in23 = reg_0358;
    78: op1_15_in23 = reg_0866;
    79: op1_15_in23 = reg_0409;
    80: op1_15_in23 = reg_0722;
    81: op1_15_in23 = reg_0438;
    82: op1_15_in23 = reg_0986;
    83: op1_15_in23 = imem02_in[67:64];
    84: op1_15_in23 = imem02_in[95:92];
    85: op1_15_in23 = reg_0694;
    86: op1_15_in23 = reg_0269;
    88: op1_15_in23 = reg_0391;
    89: op1_15_in23 = reg_0571;
    90: op1_15_in23 = reg_0824;
    91: op1_15_in23 = reg_0695;
    92: op1_15_in23 = reg_0337;
    93: op1_15_in23 = reg_0207;
    94: op1_15_in23 = reg_0519;
    default: op1_15_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv23 = 1;
    7: op1_15_inv23 = 1;
    11: op1_15_inv23 = 1;
    13: op1_15_inv23 = 1;
    14: op1_15_inv23 = 1;
    16: op1_15_inv23 = 1;
    21: op1_15_inv23 = 1;
    23: op1_15_inv23 = 1;
    24: op1_15_inv23 = 1;
    26: op1_15_inv23 = 1;
    30: op1_15_inv23 = 1;
    31: op1_15_inv23 = 1;
    32: op1_15_inv23 = 1;
    34: op1_15_inv23 = 1;
    36: op1_15_inv23 = 1;
    40: op1_15_inv23 = 1;
    41: op1_15_inv23 = 1;
    44: op1_15_inv23 = 1;
    45: op1_15_inv23 = 1;
    52: op1_15_inv23 = 1;
    54: op1_15_inv23 = 1;
    55: op1_15_inv23 = 1;
    56: op1_15_inv23 = 1;
    58: op1_15_inv23 = 1;
    60: op1_15_inv23 = 1;
    62: op1_15_inv23 = 1;
    63: op1_15_inv23 = 1;
    64: op1_15_inv23 = 1;
    67: op1_15_inv23 = 1;
    68: op1_15_inv23 = 1;
    70: op1_15_inv23 = 1;
    72: op1_15_inv23 = 1;
    73: op1_15_inv23 = 1;
    74: op1_15_inv23 = 1;
    77: op1_15_inv23 = 1;
    78: op1_15_inv23 = 1;
    83: op1_15_inv23 = 1;
    84: op1_15_inv23 = 1;
    87: op1_15_inv23 = 1;
    92: op1_15_inv23 = 1;
    default: op1_15_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in24 = reg_0369;
    7: op1_15_in24 = imem04_in[35:32];
    8: op1_15_in24 = reg_0577;
    9: op1_15_in24 = reg_0246;
    10: op1_15_in24 = reg_0777;
    11: op1_15_in24 = reg_0961;
    12: op1_15_in24 = imem07_in[23:20];
    13: op1_15_in24 = reg_0058;
    14: op1_15_in24 = imem07_in[31:28];
    16: op1_15_in24 = reg_0051;
    17: op1_15_in24 = reg_0297;
    18: op1_15_in24 = reg_0985;
    19: op1_15_in24 = imem05_in[83:80];
    20: op1_15_in24 = reg_0661;
    21: op1_15_in24 = reg_0142;
    23: op1_15_in24 = imem04_in[71:68];
    24: op1_15_in24 = reg_0197;
    25: op1_15_in24 = reg_0666;
    26: op1_15_in24 = reg_0717;
    27: op1_15_in24 = reg_0595;
    60: op1_15_in24 = reg_0595;
    28: op1_15_in24 = imem06_in[107:104];
    30: op1_15_in24 = reg_0291;
    31: op1_15_in24 = reg_0042;
    32: op1_15_in24 = reg_0706;
    34: op1_15_in24 = reg_0497;
    35: op1_15_in24 = reg_0141;
    36: op1_15_in24 = reg_0914;
    39: op1_15_in24 = reg_0810;
    40: op1_15_in24 = reg_0779;
    41: op1_15_in24 = reg_1020;
    58: op1_15_in24 = reg_1020;
    42: op1_15_in24 = reg_0729;
    44: op1_15_in24 = reg_0127;
    45: op1_15_in24 = reg_0539;
    46: op1_15_in24 = reg_0182;
    47: op1_15_in24 = imem01_in[31:28];
    48: op1_15_in24 = reg_0808;
    49: op1_15_in24 = reg_0947;
    50: op1_15_in24 = reg_1001;
    51: op1_15_in24 = imem02_in[83:80];
    52: op1_15_in24 = reg_0520;
    53: op1_15_in24 = imem03_in[3:0];
    54: op1_15_in24 = reg_0088;
    55: op1_15_in24 = reg_0882;
    56: op1_15_in24 = reg_0386;
    57: op1_15_in24 = imem06_in[71:68];
    62: op1_15_in24 = reg_1053;
    63: op1_15_in24 = imem04_in[3:0];
    64: op1_15_in24 = reg_0815;
    65: op1_15_in24 = reg_0319;
    66: op1_15_in24 = imem05_in[79:76];
    67: op1_15_in24 = reg_0295;
    68: op1_15_in24 = reg_0195;
    69: op1_15_in24 = reg_0760;
    70: op1_15_in24 = reg_0338;
    71: op1_15_in24 = reg_0832;
    72: op1_15_in24 = reg_0407;
    73: op1_15_in24 = reg_0784;
    74: op1_15_in24 = imem07_in[11:8];
    77: op1_15_in24 = reg_0248;
    78: op1_15_in24 = reg_0217;
    79: op1_15_in24 = reg_0108;
    80: op1_15_in24 = reg_0726;
    81: op1_15_in24 = reg_0688;
    82: op1_15_in24 = reg_0997;
    83: op1_15_in24 = imem02_in[71:68];
    84: op1_15_in24 = reg_0394;
    85: op1_15_in24 = reg_1018;
    86: op1_15_in24 = reg_0057;
    87: op1_15_in24 = reg_0734;
    88: op1_15_in24 = reg_0267;
    89: op1_15_in24 = reg_0038;
    90: op1_15_in24 = reg_0332;
    91: op1_15_in24 = reg_0152;
    92: op1_15_in24 = reg_1023;
    93: op1_15_in24 = reg_0194;
    94: op1_15_in24 = reg_0544;
    default: op1_15_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv24 = 1;
    7: op1_15_inv24 = 1;
    8: op1_15_inv24 = 1;
    9: op1_15_inv24 = 1;
    10: op1_15_inv24 = 1;
    12: op1_15_inv24 = 1;
    13: op1_15_inv24 = 1;
    14: op1_15_inv24 = 1;
    18: op1_15_inv24 = 1;
    20: op1_15_inv24 = 1;
    24: op1_15_inv24 = 1;
    27: op1_15_inv24 = 1;
    28: op1_15_inv24 = 1;
    30: op1_15_inv24 = 1;
    31: op1_15_inv24 = 1;
    39: op1_15_inv24 = 1;
    41: op1_15_inv24 = 1;
    45: op1_15_inv24 = 1;
    49: op1_15_inv24 = 1;
    52: op1_15_inv24 = 1;
    53: op1_15_inv24 = 1;
    54: op1_15_inv24 = 1;
    60: op1_15_inv24 = 1;
    63: op1_15_inv24 = 1;
    66: op1_15_inv24 = 1;
    67: op1_15_inv24 = 1;
    68: op1_15_inv24 = 1;
    69: op1_15_inv24 = 1;
    71: op1_15_inv24 = 1;
    77: op1_15_inv24 = 1;
    80: op1_15_inv24 = 1;
    82: op1_15_inv24 = 1;
    83: op1_15_inv24 = 1;
    84: op1_15_inv24 = 1;
    85: op1_15_inv24 = 1;
    88: op1_15_inv24 = 1;
    89: op1_15_inv24 = 1;
    90: op1_15_inv24 = 1;
    91: op1_15_inv24 = 1;
    93: op1_15_inv24 = 1;
    94: op1_15_inv24 = 1;
    default: op1_15_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in25 = reg_0385;
    7: op1_15_in25 = imem04_in[43:40];
    8: op1_15_in25 = reg_0622;
    9: op1_15_in25 = reg_0239;
    10: op1_15_in25 = reg_0812;
    11: op1_15_in25 = reg_0267;
    12: op1_15_in25 = imem07_in[55:52];
    13: op1_15_in25 = reg_0066;
    14: op1_15_in25 = imem07_in[71:68];
    16: op1_15_in25 = reg_0084;
    17: op1_15_in25 = reg_0076;
    18: op1_15_in25 = reg_0046;
    19: op1_15_in25 = imem05_in[123:120];
    20: op1_15_in25 = reg_0649;
    21: op1_15_in25 = reg_0138;
    23: op1_15_in25 = imem04_in[115:112];
    24: op1_15_in25 = imem01_in[15:12];
    25: op1_15_in25 = reg_0654;
    26: op1_15_in25 = reg_0703;
    27: op1_15_in25 = reg_0590;
    28: op1_15_in25 = imem06_in[111:108];
    30: op1_15_in25 = imem03_in[31:28];
    31: op1_15_in25 = reg_0294;
    32: op1_15_in25 = reg_0433;
    34: op1_15_in25 = reg_0128;
    35: op1_15_in25 = reg_0140;
    36: op1_15_in25 = reg_0042;
    39: op1_15_in25 = reg_0248;
    40: op1_15_in25 = reg_0247;
    41: op1_15_in25 = reg_0778;
    42: op1_15_in25 = reg_0708;
    44: op1_15_in25 = reg_0117;
    45: op1_15_in25 = reg_0055;
    46: op1_15_in25 = reg_0166;
    47: op1_15_in25 = imem01_in[67:64];
    48: op1_15_in25 = reg_0732;
    49: op1_15_in25 = reg_0953;
    50: op1_15_in25 = reg_0980;
    51: op1_15_in25 = reg_0363;
    52: op1_15_in25 = reg_1043;
    53: op1_15_in25 = imem03_in[51:48];
    54: op1_15_in25 = reg_0776;
    55: op1_15_in25 = imem05_in[7:4];
    56: op1_15_in25 = reg_0633;
    57: op1_15_in25 = imem06_in[87:84];
    58: op1_15_in25 = reg_1005;
    60: op1_15_in25 = reg_0781;
    62: op1_15_in25 = imem02_in[39:36];
    63: op1_15_in25 = imem04_in[11:8];
    64: op1_15_in25 = reg_0432;
    65: op1_15_in25 = reg_0581;
    66: op1_15_in25 = imem05_in[107:104];
    67: op1_15_in25 = imem05_in[83:80];
    68: op1_15_in25 = imem01_in[7:4];
    69: op1_15_in25 = reg_0445;
    70: op1_15_in25 = reg_1011;
    71: op1_15_in25 = reg_0283;
    72: op1_15_in25 = reg_0517;
    73: op1_15_in25 = reg_0819;
    74: op1_15_in25 = imem07_in[31:28];
    77: op1_15_in25 = reg_0335;
    78: op1_15_in25 = reg_0652;
    79: op1_15_in25 = reg_0586;
    80: op1_15_in25 = reg_0718;
    81: op1_15_in25 = reg_0165;
    82: op1_15_in25 = imem04_in[3:0];
    83: op1_15_in25 = imem02_in[103:100];
    84: op1_15_in25 = reg_0368;
    85: op1_15_in25 = reg_0391;
    86: op1_15_in25 = reg_0525;
    87: op1_15_in25 = reg_0624;
    88: op1_15_in25 = reg_0926;
    89: op1_15_in25 = reg_1008;
    90: op1_15_in25 = reg_0044;
    91: op1_15_in25 = reg_0970;
    92: op1_15_in25 = reg_0234;
    93: op1_15_in25 = reg_0201;
    94: op1_15_in25 = imem01_in[11:8];
    default: op1_15_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv25 = 1;
    9: op1_15_inv25 = 1;
    11: op1_15_inv25 = 1;
    13: op1_15_inv25 = 1;
    19: op1_15_inv25 = 1;
    21: op1_15_inv25 = 1;
    25: op1_15_inv25 = 1;
    26: op1_15_inv25 = 1;
    27: op1_15_inv25 = 1;
    32: op1_15_inv25 = 1;
    34: op1_15_inv25 = 1;
    36: op1_15_inv25 = 1;
    39: op1_15_inv25 = 1;
    42: op1_15_inv25 = 1;
    44: op1_15_inv25 = 1;
    45: op1_15_inv25 = 1;
    46: op1_15_inv25 = 1;
    48: op1_15_inv25 = 1;
    50: op1_15_inv25 = 1;
    51: op1_15_inv25 = 1;
    52: op1_15_inv25 = 1;
    55: op1_15_inv25 = 1;
    56: op1_15_inv25 = 1;
    58: op1_15_inv25 = 1;
    60: op1_15_inv25 = 1;
    63: op1_15_inv25 = 1;
    70: op1_15_inv25 = 1;
    71: op1_15_inv25 = 1;
    73: op1_15_inv25 = 1;
    78: op1_15_inv25 = 1;
    82: op1_15_inv25 = 1;
    83: op1_15_inv25 = 1;
    84: op1_15_inv25 = 1;
    85: op1_15_inv25 = 1;
    86: op1_15_inv25 = 1;
    87: op1_15_inv25 = 1;
    89: op1_15_inv25 = 1;
    92: op1_15_inv25 = 1;
    93: op1_15_inv25 = 1;
    default: op1_15_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in26 = reg_0006;
    7: op1_15_in26 = imem04_in[51:48];
    8: op1_15_in26 = reg_0372;
    9: op1_15_in26 = reg_0242;
    10: op1_15_in26 = reg_0523;
    11: op1_15_in26 = reg_0262;
    12: op1_15_in26 = imem07_in[59:56];
    13: op1_15_in26 = imem05_in[7:4];
    90: op1_15_in26 = imem05_in[7:4];
    14: op1_15_in26 = imem07_in[111:108];
    16: op1_15_in26 = reg_0094;
    17: op1_15_in26 = reg_0068;
    18: op1_15_in26 = reg_0742;
    19: op1_15_in26 = reg_0955;
    20: op1_15_in26 = reg_0663;
    21: op1_15_in26 = reg_0153;
    23: op1_15_in26 = reg_0281;
    24: op1_15_in26 = reg_0762;
    25: op1_15_in26 = reg_0639;
    51: op1_15_in26 = reg_0639;
    26: op1_15_in26 = reg_0712;
    27: op1_15_in26 = reg_0387;
    28: op1_15_in26 = imem06_in[127:124];
    30: op1_15_in26 = imem03_in[55:52];
    31: op1_15_in26 = reg_0391;
    32: op1_15_in26 = reg_0420;
    34: op1_15_in26 = reg_0139;
    35: op1_15_in26 = imem06_in[15:12];
    36: op1_15_in26 = reg_0264;
    39: op1_15_in26 = reg_0487;
    40: op1_15_in26 = reg_0828;
    41: op1_15_in26 = reg_0931;
    42: op1_15_in26 = reg_0709;
    44: op1_15_in26 = imem02_in[7:4];
    45: op1_15_in26 = reg_0537;
    46: op1_15_in26 = reg_0157;
    47: op1_15_in26 = imem01_in[75:72];
    48: op1_15_in26 = reg_0308;
    49: op1_15_in26 = reg_0835;
    50: op1_15_in26 = imem04_in[19:16];
    63: op1_15_in26 = imem04_in[19:16];
    52: op1_15_in26 = reg_0829;
    53: op1_15_in26 = imem03_in[83:80];
    54: op1_15_in26 = reg_0484;
    55: op1_15_in26 = imem05_in[11:8];
    56: op1_15_in26 = reg_0008;
    57: op1_15_in26 = imem06_in[107:104];
    58: op1_15_in26 = reg_0752;
    60: op1_15_in26 = reg_0863;
    62: op1_15_in26 = imem02_in[43:40];
    64: op1_15_in26 = reg_0407;
    65: op1_15_in26 = reg_0235;
    66: op1_15_in26 = reg_0132;
    67: op1_15_in26 = imem05_in[95:92];
    68: op1_15_in26 = imem01_in[39:36];
    69: op1_15_in26 = reg_0434;
    70: op1_15_in26 = reg_1030;
    71: op1_15_in26 = imem02_in[19:16];
    72: op1_15_in26 = reg_0251;
    73: op1_15_in26 = reg_0148;
    74: op1_15_in26 = imem07_in[55:52];
    77: op1_15_in26 = reg_0761;
    78: op1_15_in26 = reg_0128;
    79: op1_15_in26 = reg_0676;
    80: op1_15_in26 = reg_0563;
    81: op1_15_in26 = reg_0162;
    82: op1_15_in26 = imem04_in[7:4];
    83: op1_15_in26 = imem02_in[119:116];
    84: op1_15_in26 = reg_0425;
    85: op1_15_in26 = reg_0021;
    86: op1_15_in26 = reg_0948;
    87: op1_15_in26 = imem03_in[23:20];
    88: op1_15_in26 = reg_0379;
    89: op1_15_in26 = reg_0773;
    91: op1_15_in26 = reg_0145;
    92: op1_15_in26 = reg_1039;
    93: op1_15_in26 = reg_0369;
    94: op1_15_in26 = imem01_in[71:68];
    default: op1_15_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv26 = 1;
    8: op1_15_inv26 = 1;
    10: op1_15_inv26 = 1;
    12: op1_15_inv26 = 1;
    14: op1_15_inv26 = 1;
    16: op1_15_inv26 = 1;
    17: op1_15_inv26 = 1;
    18: op1_15_inv26 = 1;
    20: op1_15_inv26 = 1;
    23: op1_15_inv26 = 1;
    27: op1_15_inv26 = 1;
    28: op1_15_inv26 = 1;
    30: op1_15_inv26 = 1;
    31: op1_15_inv26 = 1;
    32: op1_15_inv26 = 1;
    34: op1_15_inv26 = 1;
    35: op1_15_inv26 = 1;
    40: op1_15_inv26 = 1;
    41: op1_15_inv26 = 1;
    45: op1_15_inv26 = 1;
    49: op1_15_inv26 = 1;
    52: op1_15_inv26 = 1;
    53: op1_15_inv26 = 1;
    54: op1_15_inv26 = 1;
    57: op1_15_inv26 = 1;
    58: op1_15_inv26 = 1;
    64: op1_15_inv26 = 1;
    66: op1_15_inv26 = 1;
    67: op1_15_inv26 = 1;
    68: op1_15_inv26 = 1;
    70: op1_15_inv26 = 1;
    71: op1_15_inv26 = 1;
    77: op1_15_inv26 = 1;
    78: op1_15_inv26 = 1;
    80: op1_15_inv26 = 1;
    81: op1_15_inv26 = 1;
    82: op1_15_inv26 = 1;
    83: op1_15_inv26 = 1;
    85: op1_15_inv26 = 1;
    91: op1_15_inv26 = 1;
    93: op1_15_inv26 = 1;
    default: op1_15_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in27 = reg_0019;
    7: op1_15_in27 = imem04_in[55:52];
    8: op1_15_in27 = reg_0407;
    9: op1_15_in27 = reg_0240;
    10: op1_15_in27 = reg_0522;
    92: op1_15_in27 = reg_0522;
    11: op1_15_in27 = reg_0270;
    12: op1_15_in27 = imem07_in[91:88];
    13: op1_15_in27 = imem05_in[43:40];
    14: op1_15_in27 = imem07_in[115:112];
    16: op1_15_in27 = imem03_in[7:4];
    17: op1_15_in27 = reg_0063;
    18: op1_15_in27 = reg_0819;
    19: op1_15_in27 = reg_0956;
    20: op1_15_in27 = reg_0364;
    21: op1_15_in27 = reg_0131;
    23: op1_15_in27 = reg_0749;
    24: op1_15_in27 = reg_0246;
    25: op1_15_in27 = reg_0641;
    26: op1_15_in27 = reg_0708;
    27: op1_15_in27 = reg_0385;
    28: op1_15_in27 = reg_0628;
    30: op1_15_in27 = imem03_in[99:96];
    31: op1_15_in27 = reg_0393;
    32: op1_15_in27 = reg_0172;
    34: op1_15_in27 = reg_0140;
    35: op1_15_in27 = imem06_in[47:44];
    36: op1_15_in27 = reg_0399;
    39: op1_15_in27 = reg_1043;
    40: op1_15_in27 = reg_0544;
    41: op1_15_in27 = reg_0763;
    48: op1_15_in27 = reg_0763;
    42: op1_15_in27 = reg_0718;
    44: op1_15_in27 = imem02_in[27:24];
    45: op1_15_in27 = reg_0584;
    46: op1_15_in27 = reg_0158;
    47: op1_15_in27 = imem01_in[87:84];
    49: op1_15_in27 = reg_0900;
    50: op1_15_in27 = imem04_in[27:24];
    63: op1_15_in27 = imem04_in[27:24];
    51: op1_15_in27 = reg_0651;
    52: op1_15_in27 = reg_0740;
    53: op1_15_in27 = imem03_in[91:88];
    54: op1_15_in27 = reg_0675;
    55: op1_15_in27 = imem05_in[67:64];
    56: op1_15_in27 = reg_0263;
    57: op1_15_in27 = imem06_in[119:116];
    58: op1_15_in27 = reg_0850;
    60: op1_15_in27 = reg_0380;
    62: op1_15_in27 = imem02_in[51:48];
    64: op1_15_in27 = reg_0517;
    65: op1_15_in27 = reg_0689;
    66: op1_15_in27 = reg_0143;
    67: op1_15_in27 = imem05_in[127:124];
    68: op1_15_in27 = imem01_in[51:48];
    69: op1_15_in27 = reg_0847;
    70: op1_15_in27 = reg_0624;
    71: op1_15_in27 = imem02_in[23:20];
    72: op1_15_in27 = imem05_in[19:16];
    73: op1_15_in27 = reg_0151;
    74: op1_15_in27 = reg_0722;
    77: op1_15_in27 = reg_0085;
    78: op1_15_in27 = reg_0319;
    79: op1_15_in27 = reg_0955;
    80: op1_15_in27 = reg_0047;
    81: op1_15_in27 = reg_0726;
    82: op1_15_in27 = imem04_in[43:40];
    83: op1_15_in27 = imem02_in[127:124];
    84: op1_15_in27 = reg_0516;
    85: op1_15_in27 = reg_0338;
    86: op1_15_in27 = reg_0336;
    87: op1_15_in27 = imem03_in[55:52];
    88: op1_15_in27 = reg_0729;
    89: op1_15_in27 = reg_1049;
    90: op1_15_in27 = imem05_in[95:92];
    91: op1_15_in27 = reg_0486;
    93: op1_15_in27 = reg_0789;
    94: op1_15_in27 = imem01_in[95:92];
    default: op1_15_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv27 = 1;
    8: op1_15_inv27 = 1;
    9: op1_15_inv27 = 1;
    11: op1_15_inv27 = 1;
    12: op1_15_inv27 = 1;
    14: op1_15_inv27 = 1;
    18: op1_15_inv27 = 1;
    19: op1_15_inv27 = 1;
    20: op1_15_inv27 = 1;
    21: op1_15_inv27 = 1;
    24: op1_15_inv27 = 1;
    25: op1_15_inv27 = 1;
    27: op1_15_inv27 = 1;
    28: op1_15_inv27 = 1;
    30: op1_15_inv27 = 1;
    32: op1_15_inv27 = 1;
    35: op1_15_inv27 = 1;
    39: op1_15_inv27 = 1;
    40: op1_15_inv27 = 1;
    41: op1_15_inv27 = 1;
    42: op1_15_inv27 = 1;
    44: op1_15_inv27 = 1;
    46: op1_15_inv27 = 1;
    47: op1_15_inv27 = 1;
    48: op1_15_inv27 = 1;
    50: op1_15_inv27 = 1;
    51: op1_15_inv27 = 1;
    55: op1_15_inv27 = 1;
    57: op1_15_inv27 = 1;
    58: op1_15_inv27 = 1;
    62: op1_15_inv27 = 1;
    63: op1_15_inv27 = 1;
    64: op1_15_inv27 = 1;
    65: op1_15_inv27 = 1;
    68: op1_15_inv27 = 1;
    69: op1_15_inv27 = 1;
    70: op1_15_inv27 = 1;
    71: op1_15_inv27 = 1;
    72: op1_15_inv27 = 1;
    73: op1_15_inv27 = 1;
    83: op1_15_inv27 = 1;
    84: op1_15_inv27 = 1;
    85: op1_15_inv27 = 1;
    87: op1_15_inv27 = 1;
    89: op1_15_inv27 = 1;
    90: op1_15_inv27 = 1;
    91: op1_15_inv27 = 1;
    default: op1_15_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in28 = reg_0014;
    7: op1_15_in28 = imem04_in[59:56];
    8: op1_15_in28 = reg_0404;
    9: op1_15_in28 = reg_0237;
    10: op1_15_in28 = reg_0513;
    11: op1_15_in28 = reg_0274;
    12: op1_15_in28 = imem07_in[107:104];
    13: op1_15_in28 = imem05_in[47:44];
    14: op1_15_in28 = reg_0723;
    16: op1_15_in28 = imem03_in[23:20];
    17: op1_15_in28 = reg_0075;
    18: op1_15_in28 = reg_0843;
    19: op1_15_in28 = reg_0948;
    20: op1_15_in28 = reg_0320;
    21: op1_15_in28 = imem06_in[3:0];
    23: op1_15_in28 = reg_0829;
    24: op1_15_in28 = reg_0502;
    25: op1_15_in28 = reg_0662;
    26: op1_15_in28 = reg_0709;
    27: op1_15_in28 = reg_0398;
    28: op1_15_in28 = reg_0626;
    30: op1_15_in28 = reg_0583;
    31: op1_15_in28 = reg_0399;
    32: op1_15_in28 = reg_0181;
    34: op1_15_in28 = reg_0134;
    35: op1_15_in28 = imem06_in[79:76];
    36: op1_15_in28 = reg_0804;
    39: op1_15_in28 = reg_1044;
    40: op1_15_in28 = imem01_in[11:8];
    41: op1_15_in28 = reg_0062;
    42: op1_15_in28 = reg_0706;
    44: op1_15_in28 = imem02_in[51:48];
    45: op1_15_in28 = reg_0815;
    58: op1_15_in28 = reg_0815;
    47: op1_15_in28 = imem01_in[123:120];
    48: op1_15_in28 = reg_0446;
    49: op1_15_in28 = reg_0229;
    50: op1_15_in28 = imem04_in[67:64];
    51: op1_15_in28 = reg_0648;
    52: op1_15_in28 = reg_0304;
    53: op1_15_in28 = imem03_in[103:100];
    54: op1_15_in28 = reg_0673;
    55: op1_15_in28 = imem05_in[107:104];
    56: op1_15_in28 = imem07_in[3:0];
    57: op1_15_in28 = reg_0293;
    60: op1_15_in28 = reg_0695;
    62: op1_15_in28 = imem02_in[59:56];
    63: op1_15_in28 = imem04_in[39:36];
    64: op1_15_in28 = reg_0495;
    65: op1_15_in28 = imem05_in[51:48];
    66: op1_15_in28 = reg_0141;
    67: op1_15_in28 = reg_0962;
    68: op1_15_in28 = imem01_in[55:52];
    69: op1_15_in28 = reg_0543;
    70: op1_15_in28 = reg_0382;
    71: op1_15_in28 = imem02_in[31:28];
    72: op1_15_in28 = imem05_in[119:116];
    73: op1_15_in28 = reg_0152;
    74: op1_15_in28 = reg_0720;
    77: op1_15_in28 = reg_0049;
    78: op1_15_in28 = reg_0655;
    79: op1_15_in28 = reg_0129;
    80: op1_15_in28 = reg_0406;
    81: op1_15_in28 = reg_0717;
    82: op1_15_in28 = imem04_in[55:52];
    83: op1_15_in28 = reg_0650;
    84: op1_15_in28 = reg_0867;
    85: op1_15_in28 = reg_0817;
    86: op1_15_in28 = reg_0153;
    87: op1_15_in28 = imem03_in[59:56];
    88: op1_15_in28 = reg_0698;
    89: op1_15_in28 = reg_0820;
    90: op1_15_in28 = imem05_in[103:100];
    91: op1_15_in28 = reg_0806;
    92: op1_15_in28 = reg_1043;
    93: op1_15_in28 = reg_0968;
    94: op1_15_in28 = imem01_in[111:108];
    default: op1_15_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv28 = 1;
    8: op1_15_inv28 = 1;
    16: op1_15_inv28 = 1;
    17: op1_15_inv28 = 1;
    20: op1_15_inv28 = 1;
    23: op1_15_inv28 = 1;
    24: op1_15_inv28 = 1;
    25: op1_15_inv28 = 1;
    27: op1_15_inv28 = 1;
    28: op1_15_inv28 = 1;
    30: op1_15_inv28 = 1;
    41: op1_15_inv28 = 1;
    42: op1_15_inv28 = 1;
    44: op1_15_inv28 = 1;
    45: op1_15_inv28 = 1;
    47: op1_15_inv28 = 1;
    48: op1_15_inv28 = 1;
    50: op1_15_inv28 = 1;
    54: op1_15_inv28 = 1;
    55: op1_15_inv28 = 1;
    58: op1_15_inv28 = 1;
    62: op1_15_inv28 = 1;
    63: op1_15_inv28 = 1;
    65: op1_15_inv28 = 1;
    69: op1_15_inv28 = 1;
    71: op1_15_inv28 = 1;
    77: op1_15_inv28 = 1;
    80: op1_15_inv28 = 1;
    84: op1_15_inv28 = 1;
    85: op1_15_inv28 = 1;
    86: op1_15_inv28 = 1;
    90: op1_15_inv28 = 1;
    91: op1_15_inv28 = 1;
    94: op1_15_inv28 = 1;
    default: op1_15_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in29 = reg_0008;
    7: op1_15_in29 = imem04_in[71:68];
    8: op1_15_in29 = reg_0039;
    9: op1_15_in29 = reg_0234;
    10: op1_15_in29 = reg_0514;
    11: op1_15_in29 = reg_0264;
    12: op1_15_in29 = reg_0719;
    13: op1_15_in29 = imem05_in[71:68];
    14: op1_15_in29 = reg_0703;
    16: op1_15_in29 = imem03_in[27:24];
    17: op1_15_in29 = reg_0064;
    58: op1_15_in29 = reg_0064;
    18: op1_15_in29 = reg_0535;
    19: op1_15_in29 = reg_0942;
    20: op1_15_in29 = reg_0341;
    21: op1_15_in29 = imem06_in[39:36];
    23: op1_15_in29 = reg_0892;
    24: op1_15_in29 = reg_1056;
    25: op1_15_in29 = reg_0665;
    26: op1_15_in29 = reg_0718;
    27: op1_15_in29 = reg_0396;
    28: op1_15_in29 = reg_0622;
    30: op1_15_in29 = reg_0584;
    31: op1_15_in29 = reg_0390;
    32: op1_15_in29 = reg_0162;
    34: op1_15_in29 = imem06_in[7:4];
    35: op1_15_in29 = imem06_in[95:92];
    36: op1_15_in29 = reg_0599;
    39: op1_15_in29 = reg_0500;
    40: op1_15_in29 = imem01_in[43:40];
    41: op1_15_in29 = reg_0760;
    42: op1_15_in29 = reg_0434;
    44: op1_15_in29 = reg_0658;
    45: op1_15_in29 = reg_0809;
    47: op1_15_in29 = reg_0003;
    48: op1_15_in29 = reg_0279;
    49: op1_15_in29 = reg_0251;
    50: op1_15_in29 = imem04_in[87:84];
    63: op1_15_in29 = imem04_in[87:84];
    51: op1_15_in29 = reg_0558;
    52: op1_15_in29 = reg_0123;
    53: op1_15_in29 = reg_0006;
    54: op1_15_in29 = reg_0342;
    55: op1_15_in29 = imem05_in[111:108];
    56: op1_15_in29 = imem07_in[15:12];
    57: op1_15_in29 = reg_0741;
    60: op1_15_in29 = reg_0629;
    62: op1_15_in29 = imem02_in[75:72];
    64: op1_15_in29 = imem05_in[11:8];
    65: op1_15_in29 = imem05_in[99:96];
    66: op1_15_in29 = reg_0130;
    79: op1_15_in29 = reg_0130;
    67: op1_15_in29 = reg_0488;
    68: op1_15_in29 = imem01_in[87:84];
    69: op1_15_in29 = reg_0373;
    70: op1_15_in29 = reg_0695;
    71: op1_15_in29 = reg_0759;
    72: op1_15_in29 = reg_0690;
    73: op1_15_in29 = reg_0154;
    74: op1_15_in29 = reg_0731;
    77: op1_15_in29 = reg_0077;
    78: op1_15_in29 = reg_0226;
    80: op1_15_in29 = reg_0350;
    81: op1_15_in29 = reg_0247;
    82: op1_15_in29 = imem04_in[107:104];
    83: op1_15_in29 = reg_0896;
    84: op1_15_in29 = reg_0876;
    85: op1_15_in29 = reg_1011;
    86: op1_15_in29 = reg_0148;
    87: op1_15_in29 = reg_0681;
    88: op1_15_in29 = reg_0121;
    89: op1_15_in29 = reg_0385;
    90: op1_15_in29 = imem05_in[115:112];
    91: op1_15_in29 = reg_0706;
    92: op1_15_in29 = reg_0829;
    93: op1_15_in29 = reg_0120;
    94: op1_15_in29 = reg_0520;
    default: op1_15_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_15_inv29 = 1;
    13: op1_15_inv29 = 1;
    14: op1_15_inv29 = 1;
    17: op1_15_inv29 = 1;
    18: op1_15_inv29 = 1;
    19: op1_15_inv29 = 1;
    21: op1_15_inv29 = 1;
    23: op1_15_inv29 = 1;
    24: op1_15_inv29 = 1;
    30: op1_15_inv29 = 1;
    31: op1_15_inv29 = 1;
    35: op1_15_inv29 = 1;
    36: op1_15_inv29 = 1;
    39: op1_15_inv29 = 1;
    41: op1_15_inv29 = 1;
    47: op1_15_inv29 = 1;
    49: op1_15_inv29 = 1;
    51: op1_15_inv29 = 1;
    54: op1_15_inv29 = 1;
    55: op1_15_inv29 = 1;
    56: op1_15_inv29 = 1;
    62: op1_15_inv29 = 1;
    64: op1_15_inv29 = 1;
    67: op1_15_inv29 = 1;
    72: op1_15_inv29 = 1;
    78: op1_15_inv29 = 1;
    79: op1_15_inv29 = 1;
    81: op1_15_inv29 = 1;
    82: op1_15_inv29 = 1;
    83: op1_15_inv29 = 1;
    85: op1_15_inv29 = 1;
    87: op1_15_inv29 = 1;
    88: op1_15_inv29 = 1;
    89: op1_15_inv29 = 1;
    90: op1_15_inv29 = 1;
    92: op1_15_inv29 = 1;
    93: op1_15_inv29 = 1;
    default: op1_15_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_15_in30 = reg_0015;
    7: op1_15_in30 = imem04_in[83:80];
    8: op1_15_in30 = reg_0036;
    9: op1_15_in30 = reg_0245;
    10: op1_15_in30 = reg_0524;
    11: op1_15_in30 = reg_0269;
    12: op1_15_in30 = reg_0710;
    13: op1_15_in30 = imem05_in[87:84];
    14: op1_15_in30 = reg_0708;
    16: op1_15_in30 = imem03_in[39:36];
    17: op1_15_in30 = reg_0072;
    18: op1_15_in30 = reg_0541;
    19: op1_15_in30 = reg_0947;
    20: op1_15_in30 = reg_0329;
    21: op1_15_in30 = imem06_in[71:68];
    23: op1_15_in30 = reg_0533;
    24: op1_15_in30 = reg_0503;
    25: op1_15_in30 = reg_0341;
    26: op1_15_in30 = reg_0711;
    27: op1_15_in30 = reg_0389;
    28: op1_15_in30 = reg_0601;
    30: op1_15_in30 = reg_0585;
    31: op1_15_in30 = reg_0000;
    32: op1_15_in30 = reg_0167;
    34: op1_15_in30 = imem06_in[15:12];
    35: op1_15_in30 = imem06_in[103:100];
    36: op1_15_in30 = reg_1028;
    39: op1_15_in30 = reg_1038;
    40: op1_15_in30 = imem01_in[67:64];
    41: op1_15_in30 = reg_0259;
    42: op1_15_in30 = reg_0440;
    44: op1_15_in30 = reg_0666;
    45: op1_15_in30 = reg_0059;
    47: op1_15_in30 = reg_0510;
    48: op1_15_in30 = reg_0873;
    49: op1_15_in30 = reg_0785;
    50: op1_15_in30 = imem04_in[91:88];
    51: op1_15_in30 = reg_0080;
    52: op1_15_in30 = reg_0118;
    53: op1_15_in30 = reg_0535;
    54: op1_15_in30 = imem03_in[23:20];
    55: op1_15_in30 = reg_0970;
    56: op1_15_in30 = imem07_in[83:80];
    57: op1_15_in30 = reg_0264;
    58: op1_15_in30 = reg_0528;
    60: op1_15_in30 = reg_0594;
    62: op1_15_in30 = imem02_in[91:88];
    63: op1_15_in30 = imem04_in[95:92];
    64: op1_15_in30 = imem05_in[23:20];
    65: op1_15_in30 = reg_0215;
    66: op1_15_in30 = reg_0131;
    67: op1_15_in30 = reg_0800;
    68: op1_15_in30 = imem01_in[91:88];
    69: op1_15_in30 = reg_0836;
    70: op1_15_in30 = reg_0386;
    71: op1_15_in30 = reg_0741;
    72: op1_15_in30 = reg_0967;
    73: op1_15_in30 = reg_0153;
    74: op1_15_in30 = reg_0721;
    77: op1_15_in30 = reg_0884;
    78: op1_15_in30 = reg_0956;
    79: op1_15_in30 = reg_0447;
    80: op1_15_in30 = reg_0180;
    81: op1_15_in30 = reg_0641;
    82: op1_15_in30 = imem04_in[127:124];
    83: op1_15_in30 = reg_0885;
    84: op1_15_in30 = reg_0792;
    85: op1_15_in30 = reg_0692;
    86: op1_15_in30 = reg_1046;
    87: op1_15_in30 = reg_0228;
    88: op1_15_in30 = reg_0918;
    89: op1_15_in30 = reg_0233;
    90: op1_15_in30 = imem05_in[119:116];
    91: op1_15_in30 = reg_0951;
    92: op1_15_in30 = reg_0830;
    93: op1_15_in30 = reg_0106;
    94: op1_15_in30 = reg_0134;
    default: op1_15_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_15_inv30 = 1;
    11: op1_15_inv30 = 1;
    12: op1_15_inv30 = 1;
    13: op1_15_inv30 = 1;
    14: op1_15_inv30 = 1;
    16: op1_15_inv30 = 1;
    18: op1_15_inv30 = 1;
    19: op1_15_inv30 = 1;
    21: op1_15_inv30 = 1;
    24: op1_15_inv30 = 1;
    25: op1_15_inv30 = 1;
    27: op1_15_inv30 = 1;
    30: op1_15_inv30 = 1;
    31: op1_15_inv30 = 1;
    32: op1_15_inv30 = 1;
    35: op1_15_inv30 = 1;
    36: op1_15_inv30 = 1;
    42: op1_15_inv30 = 1;
    44: op1_15_inv30 = 1;
    47: op1_15_inv30 = 1;
    48: op1_15_inv30 = 1;
    49: op1_15_inv30 = 1;
    51: op1_15_inv30 = 1;
    52: op1_15_inv30 = 1;
    54: op1_15_inv30 = 1;
    55: op1_15_inv30 = 1;
    56: op1_15_inv30 = 1;
    62: op1_15_inv30 = 1;
    63: op1_15_inv30 = 1;
    71: op1_15_inv30 = 1;
    73: op1_15_inv30 = 1;
    74: op1_15_inv30 = 1;
    77: op1_15_inv30 = 1;
    78: op1_15_inv30 = 1;
    79: op1_15_inv30 = 1;
    85: op1_15_inv30 = 1;
    86: op1_15_inv30 = 1;
    87: op1_15_inv30 = 1;
    91: op1_15_inv30 = 1;
    94: op1_15_inv30 = 1;
    default: op1_15_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_15_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_15_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の0番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_00_in00 = reg_0926;
    7: op2_00_in00 = reg_0940;
    22: op2_00_in00 = reg_0940;
    25: op2_00_in00 = reg_0940;
    8: op2_00_in00 = reg_0497;
    9: op2_00_in00 = reg_0939;
    19: op2_00_in00 = reg_0939;
    10: op2_00_in00 = reg_1008;
    59: op2_00_in00 = reg_1008;
    11: op2_00_in00 = reg_0909;
    18: op2_00_in00 = reg_0909;
    12: op2_00_in00 = reg_1023;
    13: op2_00_in00 = reg_1009;
    14: op2_00_in00 = reg_0231;
    16: op2_00_in00 = reg_0231;
    24: op2_00_in00 = reg_0231;
    28: op2_00_in00 = reg_0231;
    34: op2_00_in00 = reg_0231;
    40: op2_00_in00 = reg_0231;
    48: op2_00_in00 = reg_0231;
    78: op2_00_in00 = reg_0231;
    98: op2_00_in00 = reg_0231;
    15: op2_00_in00 = reg_0889;
    30: op2_00_in00 = reg_0889;
    17: op2_00_in00 = reg_0838;
    31: op2_00_in00 = reg_0838;
    20: op2_00_in00 = reg_1022;
    27: op2_00_in00 = reg_1022;
    21: op2_00_in00 = reg_0907;
    29: op2_00_in00 = reg_0907;
    52: op2_00_in00 = reg_0907;
    67: op2_00_in00 = reg_0907;
    92: op2_00_in00 = reg_0907;
    23: op2_00_in00 = reg_0938;
    62: op2_00_in00 = reg_0938;
    68: op2_00_in00 = reg_0938;
    72: op2_00_in00 = reg_0938;
    84: op2_00_in00 = reg_0938;
    26: op2_00_in00 = reg_0795;
    32: op2_00_in00 = reg_0852;
    89: op2_00_in00 = reg_0852;
    33: op2_00_in00 = reg_0850;
    37: op2_00_in00 = reg_0850;
    35: op2_00_in00 = reg_0803;
    39: op2_00_in00 = reg_0803;
    45: op2_00_in00 = reg_0803;
    61: op2_00_in00 = reg_0803;
    63: op2_00_in00 = reg_0803;
    97: op2_00_in00 = reg_0803;
    36: op2_00_in00 = reg_0415;
    47: op2_00_in00 = reg_0415;
    50: op2_00_in00 = reg_0415;
    57: op2_00_in00 = reg_0415;
    60: op2_00_in00 = reg_0415;
    65: op2_00_in00 = reg_0415;
    80: op2_00_in00 = reg_0415;
    93: op2_00_in00 = reg_0415;
    38: op2_00_in00 = reg_0414;
    51: op2_00_in00 = reg_0414;
    58: op2_00_in00 = reg_0414;
    75: op2_00_in00 = reg_0414;
    82: op2_00_in00 = reg_0414;
    87: op2_00_in00 = reg_0414;
    90: op2_00_in00 = reg_0414;
    41: op2_00_in00 = reg_0417;
    94: op2_00_in00 = reg_0417;
    42: op2_00_in00 = reg_0635;
    96: op2_00_in00 = reg_0635;
    43: op2_00_in00 = reg_0634;
    55: op2_00_in00 = reg_0634;
    44: op2_00_in00 = reg_0873;
    46: op2_00_in00 = reg_0853;
    49: op2_00_in00 = reg_0853;
    54: op2_00_in00 = reg_0853;
    64: op2_00_in00 = reg_0853;
    70: op2_00_in00 = reg_0853;
    73: op2_00_in00 = reg_0853;
    86: op2_00_in00 = reg_0853;
    95: op2_00_in00 = reg_0853;
    53: op2_00_in00 = reg_0416;
    56: op2_00_in00 = reg_0416;
    71: op2_00_in00 = reg_0416;
    79: op2_00_in00 = reg_0416;
    85: op2_00_in00 = reg_0416;
    91: op2_00_in00 = reg_0416;
    66: op2_00_in00 = reg_0851;
    69: op2_00_in00 = reg_0851;
    74: op2_00_in00 = reg_0594;
    76: op2_00_in00 = reg_0593;
    77: op2_00_in00 = reg_0493;
    81: op2_00_in00 = reg_0603;
    83: op2_00_in00 = reg_0574;
    88: op2_00_in00 = reg_0413;
    default: op2_00_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の1番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_00_in01 = reg_0927;
    8: op2_00_in01 = reg_0927;
    31: op2_00_in01 = reg_0927;
    35: op2_00_in01 = reg_0927;
    39: op2_00_in01 = reg_0927;
    45: op2_00_in01 = reg_0927;
    61: op2_00_in01 = reg_0927;
    77: op2_00_in01 = reg_0927;
    7: op2_00_in01 = reg_0941;
    22: op2_00_in01 = reg_0941;
    25: op2_00_in01 = reg_0941;
    55: op2_00_in01 = reg_0941;
    9: op2_00_in01 = reg_1022;
    15: op2_00_in01 = reg_1022;
    10: op2_00_in01 = reg_1009;
    11: op2_00_in01 = reg_0917;
    18: op2_00_in01 = reg_0917;
    27: op2_00_in01 = reg_0917;
    12: op2_00_in01 = reg_0231;
    26: op2_00_in01 = reg_0231;
    42: op2_00_in01 = reg_0231;
    46: op2_00_in01 = reg_0231;
    54: op2_00_in01 = reg_0231;
    64: op2_00_in01 = reg_0231;
    70: op2_00_in01 = reg_0231;
    86: op2_00_in01 = reg_0231;
    94: op2_00_in01 = reg_0231;
    96: op2_00_in01 = reg_0231;
    13: op2_00_in01 = reg_0940;
    19: op2_00_in01 = reg_0940;
    29: op2_00_in01 = reg_0940;
    81: op2_00_in01 = reg_0940;
    14: op2_00_in01 = reg_0525;
    63: op2_00_in01 = reg_0525;
    97: op2_00_in01 = reg_0525;
    16: op2_00_in01 = reg_0280;
    24: op2_00_in01 = reg_0280;
    28: op2_00_in01 = reg_0280;
    34: op2_00_in01 = reg_0280;
    40: op2_00_in01 = reg_0280;
    48: op2_00_in01 = reg_0280;
    78: op2_00_in01 = reg_0280;
    98: op2_00_in01 = reg_0280;
    17: op2_00_in01 = reg_0839;
    20: op2_00_in01 = reg_1023;
    32: op2_00_in01 = reg_1023;
    21: op2_00_in01 = reg_0909;
    30: op2_00_in01 = reg_0909;
    36: op2_00_in01 = reg_0909;
    23: op2_00_in01 = reg_0939;
    33: op2_00_in01 = reg_0603;
    38: op2_00_in01 = reg_0603;
    44: op2_00_in01 = reg_0603;
    58: op2_00_in01 = reg_0603;
    37: op2_00_in01 = reg_0851;
    51: op2_00_in01 = reg_0851;
    59: op2_00_in01 = reg_0851;
    62: op2_00_in01 = reg_0851;
    72: op2_00_in01 = reg_0851;
    41: op2_00_in01 = reg_0803;
    49: op2_00_in01 = reg_0803;
    95: op2_00_in01 = reg_0803;
    43: op2_00_in01 = reg_0853;
    89: op2_00_in01 = reg_0853;
    47: op2_00_in01 = reg_0416;
    50: op2_00_in01 = reg_0416;
    65: op2_00_in01 = reg_0416;
    74: op2_00_in01 = reg_0416;
    52: op2_00_in01 = reg_0634;
    66: op2_00_in01 = reg_0634;
    69: op2_00_in01 = reg_0634;
    92: op2_00_in01 = reg_0634;
    53: op2_00_in01 = reg_0417;
    56: op2_00_in01 = reg_0417;
    71: op2_00_in01 = reg_0417;
    79: op2_00_in01 = reg_0417;
    85: op2_00_in01 = reg_0417;
    91: op2_00_in01 = reg_0417;
    57: op2_00_in01 = reg_0852;
    60: op2_00_in01 = reg_0852;
    67: op2_00_in01 = reg_0852;
    80: op2_00_in01 = reg_0852;
    93: op2_00_in01 = reg_0852;
    68: op2_00_in01 = reg_0415;
    75: op2_00_in01 = reg_0415;
    73: op2_00_in01 = reg_0493;
    76: op2_00_in01 = reg_0711;
    82: op2_00_in01 = reg_0170;
    83: op2_00_in01 = reg_0593;
    88: op2_00_in01 = reg_0593;
    84: op2_00_in01 = reg_0907;
    87: op2_00_in01 = reg_0594;
    90: op2_00_in01 = reg_0594;
    default: op2_00_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の2番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_00_in02 = reg_0928;
    8: op2_00_in02 = reg_0928;
    7: op2_00_in02 = reg_0803;
    43: op2_00_in02 = reg_0803;
    53: op2_00_in02 = reg_0803;
    55: op2_00_in02 = reg_0803;
    85: op2_00_in02 = reg_0803;
    89: op2_00_in02 = reg_0803;
    91: op2_00_in02 = reg_0803;
    9: op2_00_in02 = reg_1023;
    15: op2_00_in02 = reg_1023;
    29: op2_00_in02 = reg_1023;
    66: op2_00_in02 = reg_1023;
    10: op2_00_in02 = reg_0940;
    84: op2_00_in02 = reg_0940;
    11: op2_00_in02 = reg_0838;
    25: op2_00_in02 = reg_0838;
    27: op2_00_in02 = reg_0838;
    12: op2_00_in02 = reg_0525;
    73: op2_00_in02 = reg_0525;
    13: op2_00_in02 = reg_0941;
    19: op2_00_in02 = reg_0941;
    30: op2_00_in02 = reg_0941;
    81: op2_00_in02 = reg_0941;
    14: op2_00_in02 = reg_0840;
    16: op2_00_in02 = reg_0807;
    17: op2_00_in02 = reg_0526;
    31: op2_00_in02 = reg_0526;
    35: op2_00_in02 = reg_0526;
    39: op2_00_in02 = reg_0526;
    45: op2_00_in02 = reg_0526;
    61: op2_00_in02 = reg_0526;
    63: op2_00_in02 = reg_0526;
    77: op2_00_in02 = reg_0526;
    97: op2_00_in02 = reg_0526;
    18: op2_00_in02 = reg_0231;
    20: op2_00_in02 = reg_0231;
    22: op2_00_in02 = reg_0231;
    32: op2_00_in02 = reg_0231;
    56: op2_00_in02 = reg_0231;
    21: op2_00_in02 = reg_0795;
    23: op2_00_in02 = reg_1022;
    24: op2_00_in02 = reg_0287;
    28: op2_00_in02 = reg_0287;
    34: op2_00_in02 = reg_0287;
    40: op2_00_in02 = reg_0287;
    48: op2_00_in02 = reg_0287;
    78: op2_00_in02 = reg_0287;
    98: op2_00_in02 = reg_0287;
    26: op2_00_in02 = reg_0280;
    42: op2_00_in02 = reg_0280;
    46: op2_00_in02 = reg_0280;
    54: op2_00_in02 = reg_0280;
    64: op2_00_in02 = reg_0280;
    70: op2_00_in02 = reg_0280;
    86: op2_00_in02 = reg_0280;
    94: op2_00_in02 = reg_0280;
    96: op2_00_in02 = reg_0280;
    33: op2_00_in02 = reg_0909;
    36: op2_00_in02 = reg_0853;
    67: op2_00_in02 = reg_0853;
    80: op2_00_in02 = reg_0853;
    92: op2_00_in02 = reg_0853;
    37: op2_00_in02 = reg_0416;
    44: op2_00_in02 = reg_0416;
    59: op2_00_in02 = reg_0416;
    62: op2_00_in02 = reg_0416;
    68: op2_00_in02 = reg_0416;
    82: op2_00_in02 = reg_0416;
    38: op2_00_in02 = reg_0634;
    58: op2_00_in02 = reg_0634;
    72: op2_00_in02 = reg_0634;
    75: op2_00_in02 = reg_0634;
    87: op2_00_in02 = reg_0634;
    41: op2_00_in02 = reg_0927;
    49: op2_00_in02 = reg_0927;
    95: op2_00_in02 = reg_0927;
    47: op2_00_in02 = reg_0417;
    50: op2_00_in02 = reg_0417;
    65: op2_00_in02 = reg_0417;
    74: op2_00_in02 = reg_0417;
    51: op2_00_in02 = reg_0852;
    76: op2_00_in02 = reg_0852;
    52: op2_00_in02 = reg_0635;
    57: op2_00_in02 = reg_0635;
    60: op2_00_in02 = reg_0635;
    69: op2_00_in02 = reg_0635;
    93: op2_00_in02 = reg_0635;
    71: op2_00_in02 = reg_0497;
    79: op2_00_in02 = reg_0493;
    83: op2_00_in02 = reg_0415;
    88: op2_00_in02 = reg_0415;
    90: op2_00_in02 = reg_1010;
    default: op2_00_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の3番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_00_in03 = reg_0929;
    8: op2_00_in03 = reg_0929;
    7: op2_00_in03 = reg_0804;
    11: op2_00_in03 = reg_0804;
    25: op2_00_in03 = reg_0804;
    9: op2_00_in03 = reg_0838;
    13: op2_00_in03 = reg_0838;
    15: op2_00_in03 = reg_0838;
    19: op2_00_in03 = reg_0838;
    21: op2_00_in03 = reg_0838;
    29: op2_00_in03 = reg_0838;
    10: op2_00_in03 = reg_0941;
    33: op2_00_in03 = reg_0941;
    37: op2_00_in03 = reg_0941;
    51: op2_00_in03 = reg_0941;
    84: op2_00_in03 = reg_0941;
    12: op2_00_in03 = reg_0840;
    14: op2_00_in03 = reg_0841;
    16: op2_00_in03 = reg_0809;
    24: op2_00_in03 = reg_0809;
    28: op2_00_in03 = reg_0809;
    34: op2_00_in03 = reg_0809;
    17: op2_00_in03 = reg_0527;
    18: op2_00_in03 = reg_0280;
    20: op2_00_in03 = reg_0280;
    22: op2_00_in03 = reg_0280;
    32: op2_00_in03 = reg_0280;
    56: op2_00_in03 = reg_0280;
    23: op2_00_in03 = reg_1023;
    26: op2_00_in03 = reg_0287;
    42: op2_00_in03 = reg_0287;
    46: op2_00_in03 = reg_0287;
    54: op2_00_in03 = reg_0287;
    64: op2_00_in03 = reg_0287;
    70: op2_00_in03 = reg_0287;
    94: op2_00_in03 = reg_0287;
    96: op2_00_in03 = reg_0287;
    27: op2_00_in03 = reg_0927;
    43: op2_00_in03 = reg_0927;
    53: op2_00_in03 = reg_0927;
    55: op2_00_in03 = reg_0927;
    79: op2_00_in03 = reg_0927;
    85: op2_00_in03 = reg_0927;
    89: op2_00_in03 = reg_0927;
    91: op2_00_in03 = reg_0927;
    30: op2_00_in03 = reg_0231;
    36: op2_00_in03 = reg_0231;
    50: op2_00_in03 = reg_0231;
    52: op2_00_in03 = reg_0231;
    60: op2_00_in03 = reg_0231;
    66: op2_00_in03 = reg_0231;
    74: op2_00_in03 = reg_0231;
    80: op2_00_in03 = reg_0231;
    92: op2_00_in03 = reg_0231;
    31: op2_00_in03 = reg_0316;
    35: op2_00_in03 = reg_0316;
    39: op2_00_in03 = reg_0316;
    45: op2_00_in03 = reg_0316;
    61: op2_00_in03 = reg_0316;
    63: op2_00_in03 = reg_0316;
    77: op2_00_in03 = reg_0316;
    97: op2_00_in03 = reg_0316;
    38: op2_00_in03 = reg_0417;
    44: op2_00_in03 = reg_0417;
    59: op2_00_in03 = reg_0417;
    62: op2_00_in03 = reg_0417;
    68: op2_00_in03 = reg_0417;
    82: op2_00_in03 = reg_0417;
    40: op2_00_in03 = reg_0590;
    41: op2_00_in03 = reg_0526;
    49: op2_00_in03 = reg_0526;
    73: op2_00_in03 = reg_0526;
    95: op2_00_in03 = reg_0526;
    47: op2_00_in03 = reg_0803;
    57: op2_00_in03 = reg_0803;
    65: op2_00_in03 = reg_0803;
    67: op2_00_in03 = reg_0803;
    93: op2_00_in03 = reg_0803;
    48: op2_00_in03 = reg_0443;
    98: op2_00_in03 = reg_0443;
    58: op2_00_in03 = reg_0853;
    76: op2_00_in03 = reg_0853;
    69: op2_00_in03 = reg_0497;
    71: op2_00_in03 = reg_0525;
    72: op2_00_in03 = reg_0635;
    75: op2_00_in03 = reg_0635;
    87: op2_00_in03 = reg_0635;
    78: op2_00_in03 = reg_0725;
    81: op2_00_in03 = reg_0493;
    83: op2_00_in03 = reg_0852;
    88: op2_00_in03 = reg_0416;
    90: op2_00_in03 = reg_0917;
    default: op2_00_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の4番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_00_in04 = reg_0930;
    8: op2_00_in04 = reg_0231;
    10: op2_00_in04 = reg_0231;
    38: op2_00_in04 = reg_0231;
    44: op2_00_in04 = reg_0231;
    58: op2_00_in04 = reg_0231;
    62: op2_00_in04 = reg_0231;
    68: op2_00_in04 = reg_0231;
    72: op2_00_in04 = reg_0231;
    76: op2_00_in04 = reg_0231;
    82: op2_00_in04 = reg_0231;
    84: op2_00_in04 = reg_0231;
    90: op2_00_in04 = reg_0231;
    9: op2_00_in04 = reg_0804;
    11: op2_00_in04 = reg_0914;
    12: op2_00_in04 = reg_0929;
    14: op2_00_in04 = reg_0844;
    15: op2_00_in04 = reg_0839;
    16: op2_00_in04 = reg_0842;
    24: op2_00_in04 = reg_0842;
    17: op2_00_in04 = reg_0846;
    18: op2_00_in04 = reg_0287;
    22: op2_00_in04 = reg_0287;
    32: op2_00_in04 = reg_0287;
    56: op2_00_in04 = reg_0287;
    19: op2_00_in04 = reg_0538;
    31: op2_00_in04 = reg_0538;
    39: op2_00_in04 = reg_0538;
    45: op2_00_in04 = reg_0538;
    61: op2_00_in04 = reg_0538;
    63: op2_00_in04 = reg_0538;
    77: op2_00_in04 = reg_0538;
    97: op2_00_in04 = reg_0538;
    21: op2_00_in04 = reg_0561;
    23: op2_00_in04 = reg_0838;
    26: op2_00_in04 = reg_0809;
    27: op2_00_in04 = reg_0526;
    53: op2_00_in04 = reg_0526;
    55: op2_00_in04 = reg_0526;
    71: op2_00_in04 = reg_0526;
    79: op2_00_in04 = reg_0526;
    85: op2_00_in04 = reg_0526;
    89: op2_00_in04 = reg_0526;
    28: op2_00_in04 = reg_0851;
    29: op2_00_in04 = reg_0927;
    47: op2_00_in04 = reg_0927;
    57: op2_00_in04 = reg_0927;
    65: op2_00_in04 = reg_0927;
    67: op2_00_in04 = reg_0927;
    69: op2_00_in04 = reg_0927;
    81: op2_00_in04 = reg_0927;
    33: op2_00_in04 = reg_0803;
    37: op2_00_in04 = reg_0803;
    51: op2_00_in04 = reg_0803;
    59: op2_00_in04 = reg_0803;
    87: op2_00_in04 = reg_0803;
    34: op2_00_in04 = reg_0340;
    40: op2_00_in04 = reg_0340;
    48: op2_00_in04 = reg_0340;
    78: op2_00_in04 = reg_0340;
    98: op2_00_in04 = reg_0340;
    35: op2_00_in04 = reg_0417;
    88: op2_00_in04 = reg_0417;
    36: op2_00_in04 = reg_0635;
    41: op2_00_in04 = reg_0316;
    49: op2_00_in04 = reg_0316;
    95: op2_00_in04 = reg_0316;
    42: op2_00_in04 = reg_0590;
    94: op2_00_in04 = reg_0590;
    96: op2_00_in04 = reg_0590;
    50: op2_00_in04 = reg_0280;
    52: op2_00_in04 = reg_0280;
    60: op2_00_in04 = reg_0280;
    66: op2_00_in04 = reg_0280;
    74: op2_00_in04 = reg_0280;
    80: op2_00_in04 = reg_0280;
    92: op2_00_in04 = reg_0280;
    54: op2_00_in04 = reg_0443;
    70: op2_00_in04 = reg_0443;
    75: op2_00_in04 = reg_0493;
    83: op2_00_in04 = reg_0853;
    93: op2_00_in04 = reg_0525;
    default: op2_00_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の5番目の入力
  always @ ( * ) begin
    case ( state )
    9: op2_00_in05 = reg_0839;
    11: op2_00_in05 = reg_0809;
    12: op2_00_in05 = reg_0930;
    16: op2_00_in05 = reg_0931;
    22: op2_00_in05 = reg_0849;
    23: op2_00_in05 = reg_0564;
    26: op2_00_in05 = reg_0566;
    27: op2_00_in05 = reg_0400;
    29: op2_00_in05 = reg_0526;
    65: op2_00_in05 = reg_0526;
    34: op2_00_in05 = reg_0416;
    37: op2_00_in05 = reg_0927;
    51: op2_00_in05 = reg_0927;
    39: op2_00_in05 = reg_0366;
    42: op2_00_in05 = reg_0340;
    94: op2_00_in05 = reg_0340;
    96: op2_00_in05 = reg_0340;
    52: op2_00_in05 = reg_0287;
    53: op2_00_in05 = reg_0316;
    79: op2_00_in05 = reg_0316;
    85: op2_00_in05 = reg_0316;
    68: op2_00_in05 = reg_0280;
    84: op2_00_in05 = reg_0280;
    75: op2_00_in05 = reg_0525;
    83: op2_00_in05 = reg_0803;
    88: op2_00_in05 = reg_0231;
    95: op2_00_in05 = reg_0538;
    98: op2_00_in05 = reg_0702;
    default: op2_00_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の6番目の入力
  always @ ( * ) begin
    case ( state )
    11: op2_00_in06 = reg_0810;
    53: op2_00_in06 = reg_0538;
    85: op2_00_in06 = reg_0538;
    84: op2_00_in06 = reg_0287;
    88: op2_00_in06 = reg_0280;
    default: op2_00_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の7番目の入力
  always @ ( * ) begin
    case ( state )
    11: op2_00_in07 = reg_0811;
    84: op2_00_in07 = reg_0725;
    88: op2_00_in07 = reg_0287;
    default: op2_00_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の8番目の入力
  always @ ( * ) begin
    case ( state )
    11: op2_00_in08 = reg_0841;
    default: op2_00_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#0のバイアス入力
  always @ ( * ) begin
    case ( state )
    6: op2_00_bias = 80;
    7: op2_00_bias = 57;
    8: op2_00_bias = 62;
    9: op2_00_bias = 81;
    10: op2_00_bias = 72;
    11: op2_00_bias = 131;
    12: op2_00_bias = 87;
    13: op2_00_bias = 59;
    14: op2_00_bias = 70;
    15: op2_00_bias = 70;
    16: op2_00_bias = 93;
    17: op2_00_bias = 62;
    18: op2_00_bias = 75;
    19: op2_00_bias = 77;
    20: op2_00_bias = 51;
    21: op2_00_bias = 75;
    22: op2_00_bias = 82;
    23: op2_00_bias = 78;
    24: op2_00_bias = 77;
    25: op2_00_bias = 68;
    26: op2_00_bias = 79;
    27: op2_00_bias = 72;
    28: op2_00_bias = 65;
    29: op2_00_bias = 101;
    30: op2_00_bias = 67;
    31: op2_00_bias = 65;
    32: op2_00_bias = 71;
    33: op2_00_bias = 76;
    34: op2_00_bias = 72;
    35: op2_00_bias = 61;
    36: op2_00_bias = 68;
    37: op2_00_bias = 73;
    38: op2_00_bias = 75;
    39: op2_00_bias = 85;
    40: op2_00_bias = 68;
    41: op2_00_bias = 69;
    42: op2_00_bias = 92;
    43: op2_00_bias = 53;
    44: op2_00_bias = 75;
    45: op2_00_bias = 66;
    46: op2_00_bias = 60;
    47: op2_00_bias = 84;
    48: op2_00_bias = 69;
    49: op2_00_bias = 64;
    50: op2_00_bias = 75;
    51: op2_00_bias = 83;
    52: op2_00_bias = 78;
    53: op2_00_bias = 83;
    54: op2_00_bias = 65;
    55: op2_00_bias = 78;
    56: op2_00_bias = 79;
    57: op2_00_bias = 81;
    58: op2_00_bias = 72;
    59: op2_00_bias = 75;
    60: op2_00_bias = 68;
    61: op2_00_bias = 84;
    62: op2_00_bias = 72;
    63: op2_00_bias = 64;
    64: op2_00_bias = 55;
    65: op2_00_bias = 74;
    66: op2_00_bias = 74;
    67: op2_00_bias = 71;
    68: op2_00_bias = 98;
    69: op2_00_bias = 79;
    70: op2_00_bias = 78;
    71: op2_00_bias = 66;
    72: op2_00_bias = 70;
    73: op2_00_bias = 63;
    74: op2_00_bias = 63;
    75: op2_00_bias = 84;
    76: op2_00_bias = 71;
    77: op2_00_bias = 69;
    78: op2_00_bias = 63;
    79: op2_00_bias = 73;
    80: op2_00_bias = 71;
    81: op2_00_bias = 75;
    82: op2_00_bias = 69;
    83: op2_00_bias = 73;
    84: op2_00_bias = 107;
    85: op2_00_bias = 102;
    86: op2_00_bias = 57;
    87: op2_00_bias = 84;
    88: op2_00_bias = 119;
    89: op2_00_bias = 74;
    90: op2_00_bias = 78;
    91: op2_00_bias = 72;
    92: op2_00_bias = 78;
    93: op2_00_bias = 65;
    94: op2_00_bias = 88;
    95: op2_00_bias = 72;
    96: op2_00_bias = 78;
    97: op2_00_bias = 67;
    98: op2_00_bias = 89;
    default: op2_00_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#1の0番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_01_in00 = reg_0931;
    12: op2_01_in00 = reg_0931;
    7: op2_01_in00 = reg_0807;
    9: op2_01_in00 = reg_0807;
    8: op2_01_in00 = reg_0930;
    17: op2_01_in00 = reg_0930;
    10: op2_01_in00 = reg_0927;
    23: op2_01_in00 = reg_0927;
    33: op2_01_in00 = reg_0927;
    59: op2_01_in00 = reg_0927;
    83: op2_01_in00 = reg_0927;
    87: op2_01_in00 = reg_0927;
    11: op2_01_in00 = reg_0815;
    13: op2_01_in00 = reg_0839;
    14: op2_01_in00 = reg_0842;
    15: op2_01_in00 = reg_0526;
    25: op2_01_in00 = reg_0526;
    37: op2_01_in00 = reg_0526;
    43: op2_01_in00 = reg_0526;
    47: op2_01_in00 = reg_0526;
    51: op2_01_in00 = reg_0526;
    57: op2_01_in00 = reg_0526;
    67: op2_01_in00 = reg_0526;
    69: op2_01_in00 = reg_0526;
    75: op2_01_in00 = reg_0526;
    81: op2_01_in00 = reg_0526;
    91: op2_01_in00 = reg_0526;
    93: op2_01_in00 = reg_0526;
    16: op2_01_in00 = reg_0844;
    18: op2_01_in00 = reg_0841;
    19: op2_01_in00 = reg_0804;
    21: op2_01_in00 = reg_0804;
    20: op2_01_in00 = reg_0287;
    50: op2_01_in00 = reg_0287;
    60: op2_01_in00 = reg_0287;
    66: op2_01_in00 = reg_0287;
    68: op2_01_in00 = reg_0287;
    74: op2_01_in00 = reg_0287;
    80: op2_01_in00 = reg_0287;
    86: op2_01_in00 = reg_0287;
    92: op2_01_in00 = reg_0287;
    22: op2_01_in00 = reg_0809;
    24: op2_01_in00 = reg_0843;
    34: op2_01_in00 = reg_0843;
    40: op2_01_in00 = reg_0843;
    42: op2_01_in00 = reg_0843;
    48: op2_01_in00 = reg_0843;
    26: op2_01_in00 = reg_0340;
    28: op2_01_in00 = reg_0340;
    54: op2_01_in00 = reg_0340;
    70: op2_01_in00 = reg_0340;
    84: op2_01_in00 = reg_0340;
    27: op2_01_in00 = reg_0316;
    29: op2_01_in00 = reg_0316;
    55: op2_01_in00 = reg_0316;
    65: op2_01_in00 = reg_0316;
    71: op2_01_in00 = reg_0316;
    73: op2_01_in00 = reg_0316;
    89: op2_01_in00 = reg_0316;
    30: op2_01_in00 = reg_0280;
    36: op2_01_in00 = reg_0280;
    38: op2_01_in00 = reg_0280;
    44: op2_01_in00 = reg_0280;
    58: op2_01_in00 = reg_0280;
    62: op2_01_in00 = reg_0280;
    72: op2_01_in00 = reg_0280;
    76: op2_01_in00 = reg_0280;
    82: op2_01_in00 = reg_0280;
    90: op2_01_in00 = reg_0280;
    31: op2_01_in00 = reg_0366;
    45: op2_01_in00 = reg_0366;
    53: op2_01_in00 = reg_0366;
    61: op2_01_in00 = reg_0366;
    63: op2_01_in00 = reg_0366;
    77: op2_01_in00 = reg_0366;
    85: op2_01_in00 = reg_0366;
    95: op2_01_in00 = reg_0366;
    97: op2_01_in00 = reg_0366;
    32: op2_01_in00 = reg_0590;
    46: op2_01_in00 = reg_0590;
    52: op2_01_in00 = reg_0590;
    35: op2_01_in00 = reg_0538;
    41: op2_01_in00 = reg_0538;
    49: op2_01_in00 = reg_0538;
    79: op2_01_in00 = reg_0538;
    39: op2_01_in00 = reg_0562;
    56: op2_01_in00 = reg_0443;
    64: op2_01_in00 = reg_0443;
    88: op2_01_in00 = reg_0443;
    78: op2_01_in00 = reg_0702;
    94: op2_01_in00 = reg_0702;
    96: op2_01_in00 = reg_0702;
    98: op2_01_in00 = reg_0378;
    default: op2_01_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の1番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_01_in01 = reg_0932;
    12: op2_01_in01 = reg_0932;
    7: op2_01_in01 = reg_0809;
    9: op2_01_in01 = reg_0809;
    20: op2_01_in01 = reg_0809;
    8: op2_01_in01 = reg_0931;
    14: op2_01_in01 = reg_0931;
    10: op2_01_in01 = reg_0928;
    11: op2_01_in01 = reg_1003;
    13: op2_01_in01 = reg_0526;
    19: op2_01_in01 = reg_0526;
    21: op2_01_in01 = reg_0526;
    23: op2_01_in01 = reg_0526;
    33: op2_01_in01 = reg_0526;
    59: op2_01_in01 = reg_0526;
    83: op2_01_in01 = reg_0526;
    87: op2_01_in01 = reg_0526;
    15: op2_01_in01 = reg_0527;
    16: op2_01_in01 = reg_0933;
    17: op2_01_in01 = reg_0811;
    54: op2_01_in01 = reg_0811;
    70: op2_01_in01 = reg_0811;
    18: op2_01_in01 = reg_0842;
    22: op2_01_in01 = reg_0842;
    24: op2_01_in01 = reg_0844;
    25: op2_01_in01 = reg_0316;
    37: op2_01_in01 = reg_0316;
    43: op2_01_in01 = reg_0316;
    47: op2_01_in01 = reg_0316;
    51: op2_01_in01 = reg_0316;
    57: op2_01_in01 = reg_0316;
    67: op2_01_in01 = reg_0316;
    69: op2_01_in01 = reg_0316;
    75: op2_01_in01 = reg_0316;
    81: op2_01_in01 = reg_0316;
    91: op2_01_in01 = reg_0316;
    93: op2_01_in01 = reg_0316;
    26: op2_01_in01 = reg_0843;
    28: op2_01_in01 = reg_0843;
    27: op2_01_in01 = reg_0538;
    29: op2_01_in01 = reg_0538;
    55: op2_01_in01 = reg_0538;
    65: op2_01_in01 = reg_0538;
    71: op2_01_in01 = reg_0538;
    73: op2_01_in01 = reg_0538;
    89: op2_01_in01 = reg_0538;
    30: op2_01_in01 = reg_0287;
    36: op2_01_in01 = reg_0287;
    38: op2_01_in01 = reg_0287;
    44: op2_01_in01 = reg_0287;
    58: op2_01_in01 = reg_0287;
    62: op2_01_in01 = reg_0287;
    72: op2_01_in01 = reg_0287;
    76: op2_01_in01 = reg_0287;
    82: op2_01_in01 = reg_0287;
    90: op2_01_in01 = reg_0287;
    31: op2_01_in01 = reg_0562;
    45: op2_01_in01 = reg_0562;
    53: op2_01_in01 = reg_0562;
    61: op2_01_in01 = reg_0562;
    63: op2_01_in01 = reg_0562;
    77: op2_01_in01 = reg_0562;
    85: op2_01_in01 = reg_0562;
    95: op2_01_in01 = reg_0562;
    97: op2_01_in01 = reg_0562;
    32: op2_01_in01 = reg_0340;
    46: op2_01_in01 = reg_0340;
    52: op2_01_in01 = reg_0340;
    56: op2_01_in01 = reg_0340;
    64: op2_01_in01 = reg_0340;
    88: op2_01_in01 = reg_0340;
    34: op2_01_in01 = reg_0378;
    40: op2_01_in01 = reg_0378;
    42: op2_01_in01 = reg_0378;
    48: op2_01_in01 = reg_0378;
    78: op2_01_in01 = reg_0378;
    94: op2_01_in01 = reg_0378;
    96: op2_01_in01 = reg_0378;
    35: op2_01_in01 = reg_0366;
    41: op2_01_in01 = reg_0366;
    49: op2_01_in01 = reg_0366;
    79: op2_01_in01 = reg_0366;
    39: op2_01_in01 = reg_0400;
    50: op2_01_in01 = reg_0443;
    60: op2_01_in01 = reg_0443;
    68: op2_01_in01 = reg_0443;
    74: op2_01_in01 = reg_0443;
    80: op2_01_in01 = reg_0443;
    86: op2_01_in01 = reg_0443;
    92: op2_01_in01 = reg_0443;
    66: op2_01_in01 = reg_0929;
    84: op2_01_in01 = reg_0702;
    98: op2_01_in01 = reg_0564;
    default: op2_01_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の2番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_01_in02 = reg_0933;
    12: op2_01_in02 = reg_0933;
    24: op2_01_in02 = reg_0933;
    7: op2_01_in02 = reg_0810;
    9: op2_01_in02 = reg_0810;
    15: op2_01_in02 = reg_0810;
    8: op2_01_in02 = reg_0932;
    14: op2_01_in02 = reg_0932;
    17: op2_01_in02 = reg_0932;
    10: op2_01_in02 = reg_0929;
    11: op2_01_in02 = reg_1004;
    13: op2_01_in02 = reg_0527;
    19: op2_01_in02 = reg_0527;
    21: op2_01_in02 = reg_0527;
    16: op2_01_in02 = reg_0934;
    18: op2_01_in02 = reg_0931;
    20: op2_01_in02 = reg_0842;
    22: op2_01_in02 = reg_0843;
    32: op2_01_in02 = reg_0843;
    46: op2_01_in02 = reg_0843;
    23: op2_01_in02 = reg_0316;
    33: op2_01_in02 = reg_0316;
    59: op2_01_in02 = reg_0316;
    83: op2_01_in02 = reg_0316;
    87: op2_01_in02 = reg_0316;
    25: op2_01_in02 = reg_0538;
    37: op2_01_in02 = reg_0538;
    43: op2_01_in02 = reg_0538;
    47: op2_01_in02 = reg_0538;
    51: op2_01_in02 = reg_0538;
    57: op2_01_in02 = reg_0538;
    67: op2_01_in02 = reg_0538;
    69: op2_01_in02 = reg_0538;
    75: op2_01_in02 = reg_0538;
    81: op2_01_in02 = reg_0538;
    91: op2_01_in02 = reg_0538;
    93: op2_01_in02 = reg_0538;
    26: op2_01_in02 = reg_0844;
    27: op2_01_in02 = reg_0366;
    29: op2_01_in02 = reg_0366;
    55: op2_01_in02 = reg_0366;
    65: op2_01_in02 = reg_0366;
    71: op2_01_in02 = reg_0366;
    73: op2_01_in02 = reg_0366;
    89: op2_01_in02 = reg_0366;
    28: op2_01_in02 = reg_0378;
    54: op2_01_in02 = reg_0378;
    70: op2_01_in02 = reg_0378;
    84: op2_01_in02 = reg_0378;
    30: op2_01_in02 = reg_0809;
    31: op2_01_in02 = reg_0400;
    45: op2_01_in02 = reg_0400;
    53: op2_01_in02 = reg_0400;
    61: op2_01_in02 = reg_0400;
    63: op2_01_in02 = reg_0400;
    77: op2_01_in02 = reg_0400;
    85: op2_01_in02 = reg_0400;
    95: op2_01_in02 = reg_0400;
    97: op2_01_in02 = reg_0400;
    34: op2_01_in02 = reg_0564;
    40: op2_01_in02 = reg_0564;
    42: op2_01_in02 = reg_0564;
    48: op2_01_in02 = reg_0564;
    78: op2_01_in02 = reg_0564;
    94: op2_01_in02 = reg_0564;
    96: op2_01_in02 = reg_0564;
    35: op2_01_in02 = reg_0562;
    41: op2_01_in02 = reg_0562;
    49: op2_01_in02 = reg_0562;
    79: op2_01_in02 = reg_0562;
    36: op2_01_in02 = reg_0590;
    38: op2_01_in02 = reg_0590;
    44: op2_01_in02 = reg_0590;
    39: op2_01_in02 = reg_0410;
    50: op2_01_in02 = reg_0340;
    60: op2_01_in02 = reg_0340;
    66: op2_01_in02 = reg_0340;
    68: op2_01_in02 = reg_0340;
    74: op2_01_in02 = reg_0340;
    80: op2_01_in02 = reg_0340;
    86: op2_01_in02 = reg_0340;
    92: op2_01_in02 = reg_0340;
    52: op2_01_in02 = reg_0811;
    56: op2_01_in02 = reg_0811;
    64: op2_01_in02 = reg_0811;
    58: op2_01_in02 = reg_0443;
    62: op2_01_in02 = reg_0443;
    72: op2_01_in02 = reg_0443;
    82: op2_01_in02 = reg_0443;
    90: op2_01_in02 = reg_0443;
    76: op2_01_in02 = reg_0725;
    88: op2_01_in02 = reg_0702;
    98: op2_01_in02 = reg_0846;
    default: op2_01_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の3番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_01_in03 = reg_0934;
    12: op2_01_in03 = reg_0934;
    24: op2_01_in03 = reg_0934;
    7: op2_01_in03 = reg_0811;
    9: op2_01_in03 = reg_0811;
    60: op2_01_in03 = reg_0811;
    66: op2_01_in03 = reg_0811;
    68: op2_01_in03 = reg_0811;
    8: op2_01_in03 = reg_0933;
    14: op2_01_in03 = reg_0933;
    10: op2_01_in03 = reg_0930;
    19: op2_01_in03 = reg_0930;
    11: op2_01_in03 = reg_1005;
    13: op2_01_in03 = reg_0810;
    15: op2_01_in03 = reg_0843;
    50: op2_01_in03 = reg_0843;
    16: op2_01_in03 = reg_0935;
    39: op2_01_in03 = reg_0935;
    17: op2_01_in03 = reg_0845;
    26: op2_01_in03 = reg_0845;
    28: op2_01_in03 = reg_0845;
    18: op2_01_in03 = reg_0844;
    22: op2_01_in03 = reg_0844;
    20: op2_01_in03 = reg_0931;
    21: op2_01_in03 = reg_0538;
    23: op2_01_in03 = reg_0538;
    33: op2_01_in03 = reg_0538;
    59: op2_01_in03 = reg_0538;
    83: op2_01_in03 = reg_0538;
    87: op2_01_in03 = reg_0538;
    25: op2_01_in03 = reg_0561;
    27: op2_01_in03 = reg_0562;
    29: op2_01_in03 = reg_0562;
    55: op2_01_in03 = reg_0562;
    65: op2_01_in03 = reg_0562;
    71: op2_01_in03 = reg_0562;
    73: op2_01_in03 = reg_0562;
    89: op2_01_in03 = reg_0562;
    30: op2_01_in03 = reg_0340;
    36: op2_01_in03 = reg_0340;
    38: op2_01_in03 = reg_0340;
    44: op2_01_in03 = reg_0340;
    58: op2_01_in03 = reg_0340;
    62: op2_01_in03 = reg_0340;
    72: op2_01_in03 = reg_0340;
    76: op2_01_in03 = reg_0340;
    82: op2_01_in03 = reg_0340;
    90: op2_01_in03 = reg_0340;
    31: op2_01_in03 = reg_0410;
    45: op2_01_in03 = reg_0410;
    53: op2_01_in03 = reg_0410;
    61: op2_01_in03 = reg_0410;
    63: op2_01_in03 = reg_0410;
    77: op2_01_in03 = reg_0410;
    85: op2_01_in03 = reg_0410;
    95: op2_01_in03 = reg_0410;
    97: op2_01_in03 = reg_0410;
    32: op2_01_in03 = reg_0378;
    46: op2_01_in03 = reg_0378;
    52: op2_01_in03 = reg_0378;
    56: op2_01_in03 = reg_0378;
    64: op2_01_in03 = reg_0378;
    88: op2_01_in03 = reg_0378;
    34: op2_01_in03 = reg_0846;
    40: op2_01_in03 = reg_0846;
    42: op2_01_in03 = reg_0846;
    48: op2_01_in03 = reg_0846;
    94: op2_01_in03 = reg_0846;
    96: op2_01_in03 = reg_0846;
    35: op2_01_in03 = reg_0400;
    41: op2_01_in03 = reg_0400;
    49: op2_01_in03 = reg_0400;
    79: op2_01_in03 = reg_0400;
    37: op2_01_in03 = reg_0366;
    43: op2_01_in03 = reg_0366;
    47: op2_01_in03 = reg_0366;
    51: op2_01_in03 = reg_0366;
    57: op2_01_in03 = reg_0366;
    67: op2_01_in03 = reg_0366;
    69: op2_01_in03 = reg_0366;
    75: op2_01_in03 = reg_0366;
    81: op2_01_in03 = reg_0366;
    91: op2_01_in03 = reg_0366;
    93: op2_01_in03 = reg_0366;
    54: op2_01_in03 = reg_0564;
    70: op2_01_in03 = reg_0564;
    84: op2_01_in03 = reg_0564;
    74: op2_01_in03 = reg_0702;
    80: op2_01_in03 = reg_0702;
    86: op2_01_in03 = reg_0702;
    92: op2_01_in03 = reg_0702;
    78: op2_01_in03 = reg_0565;
    98: op2_01_in03 = reg_0411;
    default: op2_01_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の4番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_01_in04 = reg_0935;
    45: op2_01_in04 = reg_0935;
    53: op2_01_in04 = reg_0935;
    8: op2_01_in04 = reg_0934;
    9: op2_01_in04 = reg_0815;
    15: op2_01_in04 = reg_0815;
    10: op2_01_in04 = reg_0840;
    11: op2_01_in04 = reg_1006;
    12: op2_01_in04 = reg_0842;
    13: op2_01_in04 = reg_0811;
    58: op2_01_in04 = reg_0811;
    62: op2_01_in04 = reg_0811;
    72: op2_01_in04 = reg_0811;
    16: op2_01_in04 = reg_0936;
    17: op2_01_in04 = reg_1004;
    18: op2_01_in04 = reg_0933;
    22: op2_01_in04 = reg_0933;
    20: op2_01_in04 = reg_0844;
    21: op2_01_in04 = reg_0562;
    37: op2_01_in04 = reg_0562;
    43: op2_01_in04 = reg_0562;
    47: op2_01_in04 = reg_0562;
    51: op2_01_in04 = reg_0562;
    57: op2_01_in04 = reg_0562;
    67: op2_01_in04 = reg_0562;
    75: op2_01_in04 = reg_0562;
    81: op2_01_in04 = reg_0562;
    91: op2_01_in04 = reg_0562;
    93: op2_01_in04 = reg_0562;
    23: op2_01_in04 = reg_0565;
    24: op2_01_in04 = reg_0847;
    26: op2_01_in04 = reg_0846;
    28: op2_01_in04 = reg_0846;
    54: op2_01_in04 = reg_0846;
    70: op2_01_in04 = reg_0846;
    27: op2_01_in04 = reg_0850;
    29: op2_01_in04 = reg_0400;
    55: op2_01_in04 = reg_0400;
    65: op2_01_in04 = reg_0400;
    73: op2_01_in04 = reg_0400;
    89: op2_01_in04 = reg_0400;
    30: op2_01_in04 = reg_0411;
    34: op2_01_in04 = reg_0411;
    40: op2_01_in04 = reg_0411;
    48: op2_01_in04 = reg_0411;
    94: op2_01_in04 = reg_0411;
    96: op2_01_in04 = reg_0411;
    32: op2_01_in04 = reg_0564;
    46: op2_01_in04 = reg_0564;
    52: op2_01_in04 = reg_0564;
    56: op2_01_in04 = reg_0564;
    64: op2_01_in04 = reg_0564;
    88: op2_01_in04 = reg_0564;
    33: op2_01_in04 = reg_0366;
    59: op2_01_in04 = reg_0366;
    83: op2_01_in04 = reg_0366;
    87: op2_01_in04 = reg_0366;
    35: op2_01_in04 = reg_0410;
    41: op2_01_in04 = reg_0410;
    79: op2_01_in04 = reg_0410;
    36: op2_01_in04 = reg_0843;
    38: op2_01_in04 = reg_0843;
    44: op2_01_in04 = reg_0843;
    39: op2_01_in04 = reg_0848;
    50: op2_01_in04 = reg_0378;
    60: op2_01_in04 = reg_0378;
    66: op2_01_in04 = reg_0378;
    68: op2_01_in04 = reg_0378;
    74: op2_01_in04 = reg_0378;
    80: op2_01_in04 = reg_0378;
    86: op2_01_in04 = reg_0378;
    92: op2_01_in04 = reg_0378;
    61: op2_01_in04 = reg_0566;
    63: op2_01_in04 = reg_0566;
    85: op2_01_in04 = reg_0566;
    76: op2_01_in04 = reg_0702;
    82: op2_01_in04 = reg_0702;
    77: op2_01_in04 = reg_0958;
    95: op2_01_in04 = reg_0612;
    98: op2_01_in04 = reg_0412;
    default: op2_01_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の5番目の入力
  always @ ( * ) begin
    case ( state )
    11: op2_01_in05 = reg_0526;
    16: op2_01_in05 = reg_0287;
    18: op2_01_in05 = reg_0847;
    20: op2_01_in05 = reg_0933;
    26: op2_01_in05 = reg_0378;
    58: op2_01_in05 = reg_0378;
    29: op2_01_in05 = reg_0410;
    55: op2_01_in05 = reg_0410;
    33: op2_01_in05 = reg_0413;
    39: op2_01_in05 = reg_0413;
    34: op2_01_in05 = reg_0412;
    51: op2_01_in05 = reg_0400;
    57: op2_01_in05 = reg_0400;
    52: op2_01_in05 = reg_0846;
    88: op2_01_in05 = reg_0846;
    61: op2_01_in05 = reg_0550;
    80: op2_01_in05 = reg_0564;
    83: op2_01_in05 = reg_0562;
    default: op2_01_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の6番目の入力
  always @ ( * ) begin
    case ( state )
    61: op2_01_in06 = reg_0413;
    default: op2_01_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#1のバイアス入力
  always @ ( * ) begin
    case ( state )
    6: op2_01_bias = 67;
    7: op2_01_bias = 55;
    8: op2_01_bias = 63;
    9: op2_01_bias = 83;
    10: op2_01_bias = 62;
    11: op2_01_bias = 67;
    12: op2_01_bias = 74;
    13: op2_01_bias = 64;
    14: op2_01_bias = 60;
    15: op2_01_bias = 74;
    16: op2_01_bias = 89;
    17: op2_01_bias = 71;
    18: op2_01_bias = 79;
    19: op2_01_bias = 58;
    20: op2_01_bias = 86;
    21: op2_01_bias = 53;
    22: op2_01_bias = 79;
    23: op2_01_bias = 65;
    24: op2_01_bias = 70;
    25: op2_01_bias = 63;
    26: op2_01_bias = 90;
    27: op2_01_bias = 72;
    28: op2_01_bias = 74;
    29: op2_01_bias = 70;
    30: op2_01_bias = 62;
    31: op2_01_bias = 55;
    32: op2_01_bias = 82;
    33: op2_01_bias = 70;
    34: op2_01_bias = 82;
    35: op2_01_bias = 67;
    36: op2_01_bias = 69;
    37: op2_01_bias = 62;
    38: op2_01_bias = 71;
    39: op2_01_bias = 84;
    40: op2_01_bias = 71;
    41: op2_01_bias = 69;
    42: op2_01_bias = 64;
    43: op2_01_bias = 73;
    44: op2_01_bias = 66;
    45: op2_01_bias = 65;
    46: op2_01_bias = 56;
    47: op2_01_bias = 64;
    48: op2_01_bias = 76;
    49: op2_01_bias = 65;
    50: op2_01_bias = 58;
    51: op2_01_bias = 80;
    52: op2_01_bias = 90;
    53: op2_01_bias = 72;
    54: op2_01_bias = 77;
    55: op2_01_bias = 86;
    56: op2_01_bias = 64;
    57: op2_01_bias = 81;
    58: op2_01_bias = 79;
    59: op2_01_bias = 77;
    60: op2_01_bias = 84;
    61: op2_01_bias = 118;
    62: op2_01_bias = 69;
    63: op2_01_bias = 68;
    64: op2_01_bias = 73;
    65: op2_01_bias = 69;
    66: op2_01_bias = 71;
    67: op2_01_bias = 64;
    68: op2_01_bias = 64;
    69: op2_01_bias = 64;
    70: op2_01_bias = 72;
    71: op2_01_bias = 51;
    72: op2_01_bias = 78;
    73: op2_01_bias = 68;
    74: op2_01_bias = 74;
    75: op2_01_bias = 61;
    76: op2_01_bias = 82;
    77: op2_01_bias = 57;
    78: op2_01_bias = 61;
    79: op2_01_bias = 58;
    80: op2_01_bias = 81;
    81: op2_01_bias = 56;
    82: op2_01_bias = 72;
    83: op2_01_bias = 84;
    84: op2_01_bias = 57;
    85: op2_01_bias = 61;
    86: op2_01_bias = 74;
    87: op2_01_bias = 71;
    88: op2_01_bias = 86;
    89: op2_01_bias = 61;
    90: op2_01_bias = 64;
    91: op2_01_bias = 87;
    92: op2_01_bias = 63;
    93: op2_01_bias = 72;
    94: op2_01_bias = 72;
    95: op2_01_bias = 84;
    96: op2_01_bias = 83;
    97: op2_01_bias = 50;
    98: op2_01_bias = 64;
    default: op2_01_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#2の0番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_02_in00 = reg_0936;
    24: op2_02_in00 = reg_0936;
    7: op2_02_in00 = reg_0815;
    13: op2_02_in00 = reg_0815;
    8: op2_02_in00 = reg_0935;
    12: op2_02_in00 = reg_0935;
    31: op2_02_in00 = reg_0935;
    35: op2_02_in00 = reg_0935;
    41: op2_02_in00 = reg_0935;
    55: op2_02_in00 = reg_0935;
    9: op2_02_in00 = reg_1003;
    15: op2_02_in00 = reg_1003;
    10: op2_02_in00 = reg_0931;
    11: op2_02_in00 = reg_1007;
    14: op2_02_in00 = reg_0934;
    18: op2_02_in00 = reg_0934;
    20: op2_02_in00 = reg_0934;
    22: op2_02_in00 = reg_0934;
    16: op2_02_in00 = reg_0937;
    17: op2_02_in00 = reg_1005;
    19: op2_02_in00 = reg_0811;
    21: op2_02_in00 = reg_0811;
    23: op2_02_in00 = reg_0561;
    25: op2_02_in00 = reg_0562;
    33: op2_02_in00 = reg_0562;
    59: op2_02_in00 = reg_0562;
    69: op2_02_in00 = reg_0562;
    87: op2_02_in00 = reg_0562;
    26: op2_02_in00 = reg_0847;
    79: op2_02_in00 = reg_0847;
    27: op2_02_in00 = reg_0564;
    50: op2_02_in00 = reg_0564;
    58: op2_02_in00 = reg_0564;
    60: op2_02_in00 = reg_0564;
    66: op2_02_in00 = reg_0564;
    68: op2_02_in00 = reg_0564;
    74: op2_02_in00 = reg_0564;
    86: op2_02_in00 = reg_0564;
    92: op2_02_in00 = reg_0564;
    28: op2_02_in00 = reg_0566;
    97: op2_02_in00 = reg_0566;
    29: op2_02_in00 = reg_0565;
    80: op2_02_in00 = reg_0565;
    30: op2_02_in00 = reg_0843;
    32: op2_02_in00 = reg_0846;
    46: op2_02_in00 = reg_0846;
    56: op2_02_in00 = reg_0846;
    64: op2_02_in00 = reg_0846;
    84: op2_02_in00 = reg_0846;
    34: op2_02_in00 = reg_0849;
    36: op2_02_in00 = reg_0378;
    38: op2_02_in00 = reg_0378;
    44: op2_02_in00 = reg_0378;
    62: op2_02_in00 = reg_0378;
    72: op2_02_in00 = reg_0378;
    76: op2_02_in00 = reg_0378;
    82: op2_02_in00 = reg_0378;
    37: op2_02_in00 = reg_0400;
    43: op2_02_in00 = reg_0400;
    47: op2_02_in00 = reg_0400;
    67: op2_02_in00 = reg_0400;
    71: op2_02_in00 = reg_0400;
    75: op2_02_in00 = reg_0400;
    81: op2_02_in00 = reg_0400;
    83: op2_02_in00 = reg_0400;
    91: op2_02_in00 = reg_0400;
    93: op2_02_in00 = reg_0400;
    39: op2_02_in00 = reg_0850;
    40: op2_02_in00 = reg_0412;
    48: op2_02_in00 = reg_0412;
    94: op2_02_in00 = reg_0412;
    96: op2_02_in00 = reg_0412;
    42: op2_02_in00 = reg_0411;
    52: op2_02_in00 = reg_0411;
    54: op2_02_in00 = reg_0411;
    70: op2_02_in00 = reg_0411;
    78: op2_02_in00 = reg_0411;
    88: op2_02_in00 = reg_0411;
    45: op2_02_in00 = reg_0550;
    53: op2_02_in00 = reg_0550;
    77: op2_02_in00 = reg_0550;
    49: op2_02_in00 = reg_0410;
    51: op2_02_in00 = reg_0410;
    57: op2_02_in00 = reg_0410;
    65: op2_02_in00 = reg_0410;
    73: op2_02_in00 = reg_0410;
    89: op2_02_in00 = reg_0410;
    63: op2_02_in00 = reg_0567;
    85: op2_02_in00 = reg_1006;
    95: op2_02_in00 = reg_1006;
    90: op2_02_in00 = reg_0702;
    default: op2_02_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の1番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_02_in01 = reg_0937;
    7: op2_02_in01 = reg_1003;
    13: op2_02_in01 = reg_1003;
    8: op2_02_in01 = reg_0936;
    12: op2_02_in01 = reg_0936;
    26: op2_02_in01 = reg_0936;
    9: op2_02_in01 = reg_1004;
    15: op2_02_in01 = reg_1004;
    10: op2_02_in01 = reg_0932;
    11: op2_02_in01 = reg_1019;
    14: op2_02_in01 = reg_0935;
    18: op2_02_in01 = reg_0935;
    29: op2_02_in01 = reg_0935;
    49: op2_02_in01 = reg_0935;
    51: op2_02_in01 = reg_0935;
    57: op2_02_in01 = reg_0935;
    16: op2_02_in01 = reg_0938;
    17: op2_02_in01 = reg_1006;
    19: op2_02_in01 = reg_0815;
    21: op2_02_in01 = reg_0815;
    20: op2_02_in01 = reg_0847;
    22: op2_02_in01 = reg_0847;
    73: op2_02_in01 = reg_0847;
    89: op2_02_in01 = reg_0847;
    23: op2_02_in01 = reg_0562;
    24: op2_02_in01 = reg_0849;
    25: op2_02_in01 = reg_0564;
    36: op2_02_in01 = reg_0564;
    38: op2_02_in01 = reg_0564;
    44: op2_02_in01 = reg_0564;
    62: op2_02_in01 = reg_0564;
    72: op2_02_in01 = reg_0564;
    76: op2_02_in01 = reg_0564;
    82: op2_02_in01 = reg_0564;
    27: op2_02_in01 = reg_0565;
    74: op2_02_in01 = reg_0565;
    28: op2_02_in01 = reg_0567;
    41: op2_02_in01 = reg_0567;
    97: op2_02_in01 = reg_0567;
    30: op2_02_in01 = reg_0378;
    90: op2_02_in01 = reg_0378;
    31: op2_02_in01 = reg_0848;
    35: op2_02_in01 = reg_0848;
    32: op2_02_in01 = reg_0411;
    46: op2_02_in01 = reg_0411;
    56: op2_02_in01 = reg_0411;
    64: op2_02_in01 = reg_0411;
    80: op2_02_in01 = reg_0411;
    84: op2_02_in01 = reg_0411;
    33: op2_02_in01 = reg_0400;
    59: op2_02_in01 = reg_0400;
    69: op2_02_in01 = reg_0400;
    87: op2_02_in01 = reg_0400;
    34: op2_02_in01 = reg_0873;
    37: op2_02_in01 = reg_0410;
    43: op2_02_in01 = reg_0410;
    47: op2_02_in01 = reg_0410;
    67: op2_02_in01 = reg_0410;
    71: op2_02_in01 = reg_0410;
    75: op2_02_in01 = reg_0410;
    81: op2_02_in01 = reg_0410;
    83: op2_02_in01 = reg_0410;
    91: op2_02_in01 = reg_0410;
    93: op2_02_in01 = reg_0410;
    39: op2_02_in01 = reg_0851;
    40: op2_02_in01 = reg_0574;
    48: op2_02_in01 = reg_0574;
    42: op2_02_in01 = reg_0412;
    52: op2_02_in01 = reg_0412;
    54: op2_02_in01 = reg_0412;
    70: op2_02_in01 = reg_0412;
    78: op2_02_in01 = reg_0412;
    88: op2_02_in01 = reg_0412;
    45: op2_02_in01 = reg_0413;
    53: op2_02_in01 = reg_0413;
    63: op2_02_in01 = reg_0413;
    77: op2_02_in01 = reg_0413;
    85: op2_02_in01 = reg_0413;
    94: op2_02_in01 = reg_0413;
    96: op2_02_in01 = reg_0413;
    50: op2_02_in01 = reg_0846;
    58: op2_02_in01 = reg_0846;
    60: op2_02_in01 = reg_0846;
    66: op2_02_in01 = reg_0846;
    68: op2_02_in01 = reg_0846;
    86: op2_02_in01 = reg_0846;
    92: op2_02_in01 = reg_0846;
    55: op2_02_in01 = reg_0550;
    79: op2_02_in01 = reg_0550;
    65: op2_02_in01 = reg_0566;
    95: op2_02_in01 = reg_0687;
    default: op2_02_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の2番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_02_in02 = reg_0938;
    7: op2_02_in02 = reg_1004;
    13: op2_02_in02 = reg_1004;
    82: op2_02_in02 = reg_1004;
    8: op2_02_in02 = reg_0937;
    12: op2_02_in02 = reg_0937;
    9: op2_02_in02 = reg_1005;
    15: op2_02_in02 = reg_1005;
    10: op2_02_in02 = reg_0933;
    11: op2_02_in02 = reg_0939;
    14: op2_02_in02 = reg_0936;
    18: op2_02_in02 = reg_0936;
    20: op2_02_in02 = reg_0936;
    22: op2_02_in02 = reg_0936;
    16: op2_02_in02 = reg_0907;
    17: op2_02_in02 = reg_1007;
    19: op2_02_in02 = reg_0845;
    21: op2_02_in02 = reg_0845;
    23: op2_02_in02 = reg_0845;
    24: op2_02_in02 = reg_1019;
    25: op2_02_in02 = reg_0565;
    72: op2_02_in02 = reg_0565;
    76: op2_02_in02 = reg_0565;
    26: op2_02_in02 = reg_0849;
    28: op2_02_in02 = reg_0849;
    52: op2_02_in02 = reg_0849;
    54: op2_02_in02 = reg_0849;
    27: op2_02_in02 = reg_0935;
    37: op2_02_in02 = reg_0935;
    43: op2_02_in02 = reg_0935;
    29: op2_02_in02 = reg_0848;
    30: op2_02_in02 = reg_0564;
    90: op2_02_in02 = reg_0564;
    31: op2_02_in02 = reg_0574;
    42: op2_02_in02 = reg_0574;
    70: op2_02_in02 = reg_0574;
    78: op2_02_in02 = reg_0574;
    97: op2_02_in02 = reg_0574;
    32: op2_02_in02 = reg_0567;
    65: op2_02_in02 = reg_0567;
    33: op2_02_in02 = reg_0410;
    59: op2_02_in02 = reg_0410;
    69: op2_02_in02 = reg_0410;
    87: op2_02_in02 = reg_0410;
    34: op2_02_in02 = reg_0889;
    35: op2_02_in02 = reg_0413;
    41: op2_02_in02 = reg_0413;
    55: op2_02_in02 = reg_0413;
    79: op2_02_in02 = reg_0413;
    36: op2_02_in02 = reg_0846;
    38: op2_02_in02 = reg_0846;
    44: op2_02_in02 = reg_0846;
    62: op2_02_in02 = reg_0846;
    39: op2_02_in02 = reg_0416;
    40: op2_02_in02 = reg_0414;
    48: op2_02_in02 = reg_0414;
    53: op2_02_in02 = reg_0414;
    77: op2_02_in02 = reg_0414;
    94: op2_02_in02 = reg_0414;
    96: op2_02_in02 = reg_0414;
    45: op2_02_in02 = reg_0572;
    46: op2_02_in02 = reg_0412;
    56: op2_02_in02 = reg_0412;
    64: op2_02_in02 = reg_0412;
    80: op2_02_in02 = reg_0412;
    84: op2_02_in02 = reg_0412;
    47: op2_02_in02 = reg_0566;
    67: op2_02_in02 = reg_0566;
    83: op2_02_in02 = reg_0566;
    49: op2_02_in02 = reg_0550;
    51: op2_02_in02 = reg_0550;
    57: op2_02_in02 = reg_0550;
    73: op2_02_in02 = reg_0550;
    50: op2_02_in02 = reg_0411;
    58: op2_02_in02 = reg_0411;
    60: op2_02_in02 = reg_0411;
    66: op2_02_in02 = reg_0411;
    68: op2_02_in02 = reg_0411;
    74: op2_02_in02 = reg_0411;
    86: op2_02_in02 = reg_0411;
    92: op2_02_in02 = reg_0411;
    63: op2_02_in02 = reg_1008;
    71: op2_02_in02 = reg_0847;
    75: op2_02_in02 = reg_0847;
    81: op2_02_in02 = reg_0847;
    91: op2_02_in02 = reg_0847;
    85: op2_02_in02 = reg_0593;
    88: op2_02_in02 = reg_0687;
    89: op2_02_in02 = reg_1006;
    93: op2_02_in02 = reg_0612;
    95: op2_02_in02 = reg_0575;
    default: op2_02_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の3番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_02_in03 = reg_0939;
    7: op2_02_in03 = reg_1005;
    13: op2_02_in03 = reg_1005;
    8: op2_02_in03 = reg_0938;
    12: op2_02_in03 = reg_0938;
    54: op2_02_in03 = reg_0938;
    78: op2_02_in03 = reg_0938;
    9: op2_02_in03 = reg_1006;
    15: op2_02_in03 = reg_1006;
    83: op2_02_in03 = reg_1006;
    91: op2_02_in03 = reg_1006;
    93: op2_02_in03 = reg_1006;
    10: op2_02_in03 = reg_0934;
    11: op2_02_in03 = reg_1022;
    14: op2_02_in03 = reg_0937;
    18: op2_02_in03 = reg_0937;
    20: op2_02_in03 = reg_0937;
    22: op2_02_in03 = reg_0937;
    16: op2_02_in03 = reg_0940;
    17: op2_02_in03 = reg_1008;
    26: op2_02_in03 = reg_1008;
    28: op2_02_in03 = reg_1008;
    19: op2_02_in03 = reg_0846;
    21: op2_02_in03 = reg_0846;
    23: op2_02_in03 = reg_0846;
    30: op2_02_in03 = reg_0846;
    90: op2_02_in03 = reg_0846;
    24: op2_02_in03 = reg_0907;
    63: op2_02_in03 = reg_0907;
    25: op2_02_in03 = reg_0935;
    33: op2_02_in03 = reg_0935;
    27: op2_02_in03 = reg_0848;
    37: op2_02_in03 = reg_0848;
    29: op2_02_in03 = reg_0574;
    46: op2_02_in03 = reg_0574;
    56: op2_02_in03 = reg_0574;
    64: op2_02_in03 = reg_0574;
    80: op2_02_in03 = reg_0574;
    31: op2_02_in03 = reg_0575;
    41: op2_02_in03 = reg_0575;
    97: op2_02_in03 = reg_0575;
    32: op2_02_in03 = reg_0849;
    84: op2_02_in03 = reg_0849;
    34: op2_02_in03 = reg_0852;
    35: op2_02_in03 = reg_0414;
    42: op2_02_in03 = reg_0414;
    55: op2_02_in03 = reg_0414;
    70: op2_02_in03 = reg_0414;
    79: op2_02_in03 = reg_0414;
    36: op2_02_in03 = reg_0411;
    38: op2_02_in03 = reg_0411;
    44: op2_02_in03 = reg_0411;
    62: op2_02_in03 = reg_0411;
    72: op2_02_in03 = reg_0411;
    76: op2_02_in03 = reg_0411;
    82: op2_02_in03 = reg_0411;
    39: op2_02_in03 = reg_0853;
    40: op2_02_in03 = reg_0415;
    77: op2_02_in03 = reg_0415;
    85: op2_02_in03 = reg_0415;
    95: op2_02_in03 = reg_0415;
    43: op2_02_in03 = reg_0567;
    67: op2_02_in03 = reg_0567;
    45: op2_02_in03 = reg_0851;
    48: op2_02_in03 = reg_0851;
    53: op2_02_in03 = reg_0851;
    47: op2_02_in03 = reg_0550;
    71: op2_02_in03 = reg_0550;
    75: op2_02_in03 = reg_0550;
    81: op2_02_in03 = reg_0550;
    49: op2_02_in03 = reg_0413;
    51: op2_02_in03 = reg_0413;
    57: op2_02_in03 = reg_0413;
    65: op2_02_in03 = reg_0413;
    73: op2_02_in03 = reg_0413;
    50: op2_02_in03 = reg_0412;
    58: op2_02_in03 = reg_0412;
    60: op2_02_in03 = reg_0412;
    66: op2_02_in03 = reg_0412;
    68: op2_02_in03 = reg_0412;
    74: op2_02_in03 = reg_0412;
    86: op2_02_in03 = reg_0412;
    92: op2_02_in03 = reg_0412;
    52: op2_02_in03 = reg_0873;
    88: op2_02_in03 = reg_0873;
    59: op2_02_in03 = reg_0566;
    87: op2_02_in03 = reg_0566;
    69: op2_02_in03 = reg_0958;
    89: op2_02_in03 = reg_1007;
    94: op2_02_in03 = reg_0170;
    96: op2_02_in03 = reg_0170;
    default: op2_02_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の4番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_02_in04 = reg_0497;
    7: op2_02_in04 = reg_0838;
    9: op2_02_in04 = reg_1007;
    15: op2_02_in04 = reg_1007;
    10: op2_02_in04 = reg_0935;
    23: op2_02_in04 = reg_0935;
    11: op2_02_in04 = reg_0527;
    13: op2_02_in04 = reg_1006;
    87: op2_02_in04 = reg_1006;
    14: op2_02_in04 = reg_0938;
    18: op2_02_in04 = reg_0938;
    20: op2_02_in04 = reg_0938;
    65: op2_02_in04 = reg_0938;
    16: op2_02_in04 = reg_0941;
    17: op2_02_in04 = reg_0889;
    19: op2_02_in04 = reg_0848;
    33: op2_02_in04 = reg_0848;
    21: op2_02_in04 = reg_0316;
    24: op2_02_in04 = reg_0340;
    26: op2_02_in04 = reg_0907;
    31: op2_02_in04 = reg_0907;
    27: op2_02_in04 = reg_0574;
    50: op2_02_in04 = reg_0574;
    58: op2_02_in04 = reg_0574;
    60: op2_02_in04 = reg_0574;
    66: op2_02_in04 = reg_0574;
    68: op2_02_in04 = reg_0574;
    74: op2_02_in04 = reg_0574;
    91: op2_02_in04 = reg_0574;
    29: op2_02_in04 = reg_0575;
    30: op2_02_in04 = reg_0603;
    41: op2_02_in04 = reg_0603;
    55: op2_02_in04 = reg_0603;
    78: op2_02_in04 = reg_0603;
    32: op2_02_in04 = reg_0412;
    36: op2_02_in04 = reg_0412;
    38: op2_02_in04 = reg_0412;
    44: op2_02_in04 = reg_0412;
    62: op2_02_in04 = reg_0412;
    72: op2_02_in04 = reg_0412;
    76: op2_02_in04 = reg_0412;
    82: op2_02_in04 = reg_0412;
    34: op2_02_in04 = reg_1023;
    35: op2_02_in04 = reg_0634;
    40: op2_02_in04 = reg_0634;
    45: op2_02_in04 = reg_0634;
    77: op2_02_in04 = reg_0634;
    96: op2_02_in04 = reg_0634;
    37: op2_02_in04 = reg_0413;
    43: op2_02_in04 = reg_0413;
    47: op2_02_in04 = reg_0413;
    67: op2_02_in04 = reg_0413;
    71: op2_02_in04 = reg_0413;
    75: op2_02_in04 = reg_0413;
    81: op2_02_in04 = reg_0413;
    83: op2_02_in04 = reg_0413;
    92: op2_02_in04 = reg_0413;
    42: op2_02_in04 = reg_0415;
    52: op2_02_in04 = reg_0415;
    54: op2_02_in04 = reg_0415;
    70: op2_02_in04 = reg_0415;
    97: op2_02_in04 = reg_0415;
    46: op2_02_in04 = reg_0414;
    64: op2_02_in04 = reg_0414;
    84: op2_02_in04 = reg_0414;
    48: op2_02_in04 = reg_0852;
    53: op2_02_in04 = reg_0852;
    85: op2_02_in04 = reg_0852;
    49: op2_02_in04 = reg_0572;
    51: op2_02_in04 = reg_0572;
    56: op2_02_in04 = reg_0873;
    59: op2_02_in04 = reg_0550;
    63: op2_02_in04 = reg_1022;
    73: op2_02_in04 = reg_0593;
    80: op2_02_in04 = reg_0593;
    86: op2_02_in04 = reg_0849;
    88: op2_02_in04 = reg_0170;
    94: op2_02_in04 = reg_0940;
    95: op2_02_in04 = reg_0416;
    default: op2_02_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の5番目の入力
  always @ ( * ) begin
    case ( state )
    14: op2_02_in05 = reg_0280;
    26: op2_02_in05 = reg_0567;
    29: op2_02_in05 = reg_0852;
    31: op2_02_in05 = reg_0853;
    33: op2_02_in05 = reg_0414;
    66: op2_02_in05 = reg_0414;
    68: op2_02_in05 = reg_0414;
    92: op2_02_in05 = reg_0414;
    36: op2_02_in05 = reg_0849;
    41: op2_02_in05 = reg_0416;
    97: op2_02_in05 = reg_0416;
    59: op2_02_in05 = reg_0413;
    77: op2_02_in05 = reg_0635;
    84: op2_02_in05 = reg_0711;
    91: op2_02_in05 = reg_1008;
    96: op2_02_in05 = reg_0417;
    default: op2_02_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の6番目の入力
  always @ ( * ) begin
    case ( state )
    59: op2_02_in06 = reg_0938;
    97: op2_02_in06 = reg_0853;
    default: op2_02_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#2のバイアス入力
  always @ ( * ) begin
    case ( state )
    6: op2_02_bias = 64;
    7: op2_02_bias = 66;
    8: op2_02_bias = 55;
    9: op2_02_bias = 68;
    10: op2_02_bias = 84;
    11: op2_02_bias = 57;
    12: op2_02_bias = 59;
    13: op2_02_bias = 85;
    14: op2_02_bias = 84;
    15: op2_02_bias = 79;
    16: op2_02_bias = 70;
    17: op2_02_bias = 84;
    18: op2_02_bias = 83;
    19: op2_02_bias = 79;
    20: op2_02_bias = 78;
    21: op2_02_bias = 61;
    22: op2_02_bias = 62;
    23: op2_02_bias = 71;
    24: op2_02_bias = 48;
    25: op2_02_bias = 73;
    26: op2_02_bias = 93;
    27: op2_02_bias = 65;
    28: op2_02_bias = 61;
    29: op2_02_bias = 84;
    30: op2_02_bias = 70;
    31: op2_02_bias = 69;
    32: op2_02_bias = 63;
    33: op2_02_bias = 76;
    34: op2_02_bias = 68;
    35: op2_02_bias = 69;
    36: op2_02_bias = 83;
    37: op2_02_bias = 69;
    38: op2_02_bias = 71;
    39: op2_02_bias = 63;
    40: op2_02_bias = 56;
    41: op2_02_bias = 87;
    42: op2_02_bias = 73;
    43: op2_02_bias = 62;
    44: op2_02_bias = 70;
    45: op2_02_bias = 69;
    46: op2_02_bias = 75;
    47: op2_02_bias = 70;
    48: op2_02_bias = 78;
    49: op2_02_bias = 56;
    50: op2_02_bias = 63;
    51: op2_02_bias = 79;
    52: op2_02_bias = 71;
    53: op2_02_bias = 66;
    54: op2_02_bias = 70;
    55: op2_02_bias = 78;
    56: op2_02_bias = 67;
    57: op2_02_bias = 45;
    58: op2_02_bias = 70;
    59: op2_02_bias = 85;
    60: op2_02_bias = 64;
    62: op2_02_bias = 66;
    63: op2_02_bias = 71;
    64: op2_02_bias = 70;
    65: op2_02_bias = 64;
    66: op2_02_bias = 80;
    67: op2_02_bias = 72;
    68: op2_02_bias = 86;
    69: op2_02_bias = 50;
    70: op2_02_bias = 74;
    71: op2_02_bias = 61;
    72: op2_02_bias = 65;
    73: op2_02_bias = 67;
    74: op2_02_bias = 63;
    75: op2_02_bias = 62;
    76: op2_02_bias = 63;
    77: op2_02_bias = 64;
    78: op2_02_bias = 72;
    79: op2_02_bias = 69;
    80: op2_02_bias = 73;
    81: op2_02_bias = 67;
    82: op2_02_bias = 80;
    83: op2_02_bias = 69;
    84: op2_02_bias = 97;
    85: op2_02_bias = 60;
    86: op2_02_bias = 78;
    87: op2_02_bias = 56;
    88: op2_02_bias = 61;
    89: op2_02_bias = 66;
    90: op2_02_bias = 51;
    91: op2_02_bias = 86;
    92: op2_02_bias = 69;
    93: op2_02_bias = 54;
    94: op2_02_bias = 68;
    95: op2_02_bias = 68;
    96: op2_02_bias = 83;
    97: op2_02_bias = 76;
    default: op2_02_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#3の0番目の入力
  always @ ( * ) begin
    case ( state )
    7: op2_03_in00 = reg_1006;
    10: op2_03_in00 = reg_0936;
    13: op2_03_in00 = reg_1007;
    27: op2_03_in00 = reg_1007;
    15: op2_03_in00 = reg_1008;
    19: op2_03_in00 = reg_1005;
    21: op2_03_in00 = reg_0935;
    23: op2_03_in00 = reg_0848;
    25: op2_03_in00 = reg_0848;
    30: op2_03_in00 = reg_0566;
    33: op2_03_in00 = reg_0574;
    38: op2_03_in00 = reg_0574;
    44: op2_03_in00 = reg_0574;
    62: op2_03_in00 = reg_0574;
    72: op2_03_in00 = reg_0574;
    93: op2_03_in00 = reg_0574;
    47: op2_03_in00 = reg_0593;
    60: op2_03_in00 = reg_0414;
    69: op2_03_in00 = reg_0567;
    76: op2_03_in00 = reg_0849;
    90: op2_03_in00 = reg_0411;
    default: op2_03_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の1番目の入力
  always @ ( * ) begin
    case ( state )
    7: op2_03_in01 = reg_1007;
    23: op2_03_in01 = reg_1007;
    25: op2_03_in01 = reg_1007;
    10: op2_03_in01 = reg_0937;
    13: op2_03_in01 = reg_1008;
    15: op2_03_in01 = reg_0939;
    19: op2_03_in01 = reg_1006;
    21: op2_03_in01 = reg_0848;
    27: op2_03_in01 = reg_0938;
    30: op2_03_in01 = reg_0567;
    33: op2_03_in01 = reg_0575;
    38: op2_03_in01 = reg_0575;
    44: op2_03_in01 = reg_0414;
    62: op2_03_in01 = reg_0414;
    72: op2_03_in01 = reg_0414;
    47: op2_03_in01 = reg_0603;
    60: op2_03_in01 = reg_0907;
    69: op2_03_in01 = reg_0413;
    76: op2_03_in01 = reg_0873;
    93: op2_03_in01 = reg_0873;
    90: op2_03_in01 = reg_0412;
    default: op2_03_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の2番目の入力
  always @ ( * ) begin
    case ( state )
    7: op2_03_in02 = reg_1008;
    23: op2_03_in02 = reg_1008;
    10: op2_03_in02 = reg_0938;
    25: op2_03_in02 = reg_0938;
    13: op2_03_in02 = reg_0939;
    27: op2_03_in02 = reg_0939;
    15: op2_03_in02 = reg_0909;
    19: op2_03_in02 = reg_1007;
    21: op2_03_in02 = reg_1007;
    30: op2_03_in02 = reg_0849;
    33: op2_03_in02 = reg_0851;
    38: op2_03_in02 = reg_0415;
    44: op2_03_in02 = reg_0415;
    62: op2_03_in02 = reg_0415;
    72: op2_03_in02 = reg_0415;
    47: op2_03_in02 = reg_0634;
    60: op2_03_in02 = reg_0634;
    69: op2_03_in02 = reg_0959;
    76: op2_03_in02 = reg_0603;
    93: op2_03_in02 = reg_0603;
    90: op2_03_in02 = reg_0413;
    default: op2_03_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の3番目の入力
  always @ ( * ) begin
    case ( state )
    7: op2_03_in03 = reg_1009;
    10: op2_03_in03 = reg_0907;
    69: op2_03_in03 = reg_0907;
    13: op2_03_in03 = reg_0909;
    27: op2_03_in03 = reg_0909;
    15: op2_03_in03 = reg_0917;
    19: op2_03_in03 = reg_1008;
    21: op2_03_in03 = reg_1008;
    23: op2_03_in03 = reg_0889;
    25: op2_03_in03 = reg_0889;
    30: op2_03_in03 = reg_0850;
    33: op2_03_in03 = reg_1022;
    38: op2_03_in03 = reg_0852;
    44: op2_03_in03 = reg_0852;
    62: op2_03_in03 = reg_0852;
    72: op2_03_in03 = reg_0852;
    47: op2_03_in03 = reg_0635;
    60: op2_03_in03 = reg_0853;
    76: op2_03_in03 = reg_0416;
    93: op2_03_in03 = reg_0416;
    90: op2_03_in03 = reg_0873;
    default: op2_03_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の4番目の入力
  always @ ( * ) begin
    case ( state )
    7: op2_03_in04 = reg_1010;
    10: op2_03_in04 = reg_0525;
    13: op2_03_in04 = reg_0917;
    15: op2_03_in04 = reg_0845;
    19: op2_03_in04 = reg_0889;
    21: op2_03_in04 = reg_0889;
    23: op2_03_in04 = reg_0909;
    25: op2_03_in04 = reg_0909;
    27: op2_03_in04 = reg_0941;
    30: op2_03_in04 = reg_0851;
    33: op2_03_in04 = reg_0853;
    38: op2_03_in04 = reg_0635;
    44: op2_03_in04 = reg_0635;
    62: op2_03_in04 = reg_0635;
    69: op2_03_in04 = reg_0852;
    76: op2_03_in04 = reg_0417;
    90: op2_03_in04 = reg_0170;
    default: op2_03_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の5番目の入力
  always @ ( * ) begin
    case ( state )
    7: op2_03_in05 = reg_1011;
    13: op2_03_in05 = reg_0843;
    23: op2_03_in05 = reg_0917;
    25: op2_03_in05 = reg_0366;
    27: op2_03_in05 = reg_0575;
    30: op2_03_in05 = reg_1022;
    33: op2_03_in05 = reg_0415;
    default: op2_03_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の6番目の入力
  always @ ( * ) begin
    case ( state )
    30: op2_03_in06 = reg_0501;
    default: op2_03_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#3のバイアス入力
  always @ ( * ) begin
    case ( state )
    7: op2_03_bias = 86;
    10: op2_03_bias = 73;
    13: op2_03_bias = 94;
    15: op2_03_bias = 65;
    19: op2_03_bias = 83;
    21: op2_03_bias = 70;
    23: op2_03_bias = 92;
    25: op2_03_bias = 85;
    27: op2_03_bias = 87;
    30: op2_03_bias = 107;
    33: op2_03_bias = 78;
    38: op2_03_bias = 72;
    44: op2_03_bias = 60;
    47: op2_03_bias = 64;
    60: op2_03_bias = 54;
    62: op2_03_bias = 70;
    69: op2_03_bias = 84;
    72: op2_03_bias = 51;
    76: op2_03_bias = 72;
    90: op2_03_bias = 65;
    93: op2_03_bias = 53;
    default: op2_03_bias = 0;
    endcase
  end // always @ ( * )

  // REG#0の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0000 <= imem03_in[3:0];
    7: reg_0000 <= imem03_in[3:0];
    9: reg_0000 <= imem07_in[95:92];
    11: reg_0000 <= imem03_in[3:0];
    13: reg_0000 <= imem00_in[67:64];
    15: reg_0000 <= imem07_in[95:92];
    17: reg_0000 <= imem03_in[3:0];
    19: reg_0000 <= imem06_in[127:124];
    21: reg_0000 <= imem06_in[127:124];
    23: reg_0000 <= imem00_in[67:64];
    25: reg_0000 <= imem03_in[3:0];
    27: reg_0000 <= imem07_in[95:92];
    29: reg_0000 <= imem06_in[127:124];
    54: reg_0000 <= imem03_in[3:0];
    56: reg_0000 <= imem06_in[127:124];
    60: reg_0000 <= imem00_in[67:64];
    62: reg_0000 <= imem00_in[67:64];
    64: reg_0000 <= imem06_in[127:124];
    66: reg_0000 <= imem06_in[127:124];
    68: reg_0000 <= imem00_in[67:64];
    70: reg_0000 <= imem07_in[95:92];
    72: reg_0000 <= imem00_in[67:64];
    74: reg_0000 <= imem06_in[127:124];
    76: reg_0000 <= imem07_in[95:92];
    78: reg_0000 <= imem00_in[67:64];
    80: reg_0000 <= imem07_in[95:92];
    83: reg_0000 <= imem06_in[127:124];
    85: reg_0000 <= imem03_in[3:0];
    87: reg_0000 <= imem07_in[95:92];
    89: reg_0000 <= imem03_in[3:0];
    92: reg_0000 <= imem00_in[55:52];
    94: reg_0000 <= imem04_in[19:16];
    96: reg_0000 <= imem06_in[127:124];
    endcase
  end

  // REG#1の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0001 <= imem03_in[23:20];
    7: reg_0001 <= imem03_in[23:20];
    9: reg_0001 <= imem07_in[107:104];
    11: reg_0001 <= imem07_in[107:104];
    13: reg_0001 <= imem07_in[107:104];
    15: reg_0001 <= imem07_in[107:104];
    17: reg_0001 <= imem07_in[107:104];
    19: reg_0001 <= imem00_in[3:0];
    21: reg_0001 <= imem07_in[107:104];
    23: reg_0001 <= imem07_in[107:104];
    25: reg_0001 <= imem07_in[107:104];
    27: reg_0001 <= imem00_in[3:0];
    29: reg_0001 <= imem04_in[55:52];
    31: reg_0001 <= imem07_in[107:104];
    33: reg_0001 <= imem00_in[3:0];
    35: reg_0001 <= imem06_in[111:108];
    37: reg_0001 <= imem04_in[55:52];
    39: reg_0001 <= imem04_in[55:52];
    41: reg_0001 <= imem07_in[107:104];
    43: reg_0001 <= imem00_in[3:0];
    45: reg_0001 <= imem00_in[3:0];
    47: reg_0001 <= imem03_in[23:20];
    49: reg_0001 <= imem06_in[111:108];
    51: reg_0001 <= imem00_in[3:0];
    53: reg_0001 <= imem00_in[3:0];
    55: reg_0001 <= imem00_in[3:0];
    91: reg_0001 <= imem03_in[23:20];
    93: reg_0001 <= imem04_in[55:52];
    95: reg_0001 <= imem05_in[127:124];
    97: reg_0001 <= imem06_in[111:108];
    endcase
  end

  // REG#2の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0002 <= imem03_in[27:24];
    7: reg_0002 <= imem00_in[23:20];
    9: reg_0002 <= imem00_in[19:16];
    11: reg_0002 <= imem00_in[23:20];
    13: reg_0002 <= imem03_in[27:24];
    15: reg_0002 <= imem00_in[51:48];
    17: reg_0002 <= imem04_in[99:96];
    19: reg_0002 <= imem00_in[23:20];
    21: reg_0002 <= imem04_in[99:96];
    23: reg_0002 <= imem04_in[99:96];
    25: reg_0002 <= imem03_in[27:24];
    27: reg_0002 <= imem00_in[23:20];
    29: reg_0002 <= imem00_in[51:48];
    31: reg_0002 <= imem00_in[51:48];
    33: reg_0002 <= imem00_in[19:16];
    35: reg_0002 <= imem00_in[23:20];
    37: reg_0002 <= imem07_in[15:12];
    39: reg_0002 <= imem00_in[23:20];
    41: reg_0002 <= imem07_in[15:12];
    43: reg_0002 <= imem07_in[15:12];
    endcase
  end

  // REG#3の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0003 <= imem03_in[35:32];
    7: reg_0003 <= imem03_in[35:32];
    9: reg_0003 <= imem00_in[75:72];
    11: reg_0003 <= imem00_in[75:72];
    13: reg_0003 <= imem00_in[75:72];
    15: reg_0003 <= imem01_in[31:28];
    17: reg_0003 <= imem03_in[35:32];
    19: reg_0003 <= imem01_in[31:28];
    21: reg_0003 <= imem00_in[75:72];
    23: reg_0003 <= imem00_in[111:108];
    25: reg_0003 <= imem01_in[31:28];
    49: reg_0003 <= imem00_in[111:108];
    51: reg_0003 <= imem07_in[39:36];
    53: reg_0003 <= imem01_in[31:28];
    endcase
  end

  // REG#4の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0004 <= imem03_in[115:112];
    7: reg_0004 <= imem03_in[115:112];
    9: reg_0004 <= imem02_in[15:12];
    11: reg_0004 <= imem03_in[115:112];
    13: reg_0004 <= imem03_in[115:112];
    15: reg_0004 <= imem01_in[83:80];
    17: reg_0004 <= imem01_in[83:80];
    19: reg_0004 <= imem01_in[79:76];
    21: reg_0004 <= imem01_in[79:76];
    23: reg_0004 <= imem01_in[79:76];
    25: reg_0004 <= imem02_in[15:12];
    27: reg_0004 <= imem01_in[79:76];
    29: reg_0004 <= imem01_in[79:76];
    31: reg_0004 <= imem03_in[115:112];
    54: reg_0004 <= imem01_in[79:76];
    56: reg_0004 <= imem03_in[115:112];
    58: reg_0004 <= imem02_in[15:12];
    60: reg_0004 <= imem02_in[15:12];
    62: reg_0004 <= imem03_in[115:112];
    64: reg_0004 <= imem05_in[91:88];
    66: reg_0004 <= imem05_in[91:88];
    79: reg_0004 <= imem01_in[79:76];
    81: reg_0004 <= imem01_in[83:80];
    83: reg_0004 <= imem05_in[43:40];
    85: reg_0004 <= imem01_in[79:76];
    87: reg_0004 <= imem02_in[15:12];
    89: reg_0004 <= imem03_in[115:112];
    92: reg_0004 <= imem05_in[43:40];
    94: reg_0004 <= imem02_in[15:12];
    96: reg_0004 <= imem05_in[91:88];
    endcase
  end

  // REG#5の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0005 <= imem06_in[103:100];
    7: reg_0005 <= imem06_in[103:100];
    9: reg_0005 <= imem06_in[103:100];
    32: reg_0005 <= imem06_in[103:100];
    37: reg_0005 <= imem06_in[103:100];
    62: reg_0005 <= imem00_in[127:124];
    64: reg_0005 <= imem00_in[127:124];
    66: reg_0005 <= imem06_in[107:104];
    68: reg_0005 <= imem06_in[107:104];
    70: reg_0005 <= imem06_in[107:104];
    73: reg_0005 <= imem07_in[63:60];
    75: reg_0005 <= imem06_in[103:100];
    77: reg_0005 <= imem00_in[127:124];
    79: reg_0005 <= imem06_in[103:100];
    81: reg_0005 <= imem06_in[107:104];
    83: reg_0005 <= imem00_in[127:124];
    85: reg_0005 <= imem06_in[107:104];
    88: reg_0005 <= imem00_in[127:124];
    90: reg_0005 <= imem06_in[107:104];
    92: reg_0005 <= imem00_in[127:124];
    94: reg_0005 <= imem06_in[103:100];
    96: reg_0005 <= imem06_in[103:100];
    endcase
  end

  // REG#6の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0006 <= imem03_in[7:4];
    7: reg_0006 <= imem00_in[27:24];
    9: reg_0006 <= imem03_in[7:4];
    11: reg_0006 <= imem02_in[91:88];
    13: reg_0006 <= imem00_in[27:24];
    15: reg_0006 <= imem00_in[27:24];
    17: reg_0006 <= imem00_in[27:24];
    19: reg_0006 <= imem02_in[91:88];
    21: reg_0006 <= imem03_in[7:4];
    23: reg_0006 <= imem03_in[7:4];
    25: reg_0006 <= imem02_in[75:72];
    27: reg_0006 <= imem02_in[91:88];
    29: reg_0006 <= imem00_in[27:24];
    31: reg_0006 <= imem03_in[7:4];
    55: reg_0006 <= imem03_in[7:4];
    88: reg_0006 <= imem02_in[75:72];
    90: reg_0006 <= imem02_in[91:88];
    92: reg_0006 <= imem03_in[7:4];
    94: reg_0006 <= imem02_in[75:72];
    96: reg_0006 <= imem02_in[63:60];
    endcase
  end

  // REG#7の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0007 <= imem03_in[47:44];
    7: reg_0007 <= imem03_in[47:44];
    9: reg_0007 <= imem03_in[47:44];
    11: reg_0007 <= imem03_in[47:44];
    13: reg_0007 <= imem03_in[71:68];
    15: reg_0007 <= imem03_in[47:44];
    17: reg_0007 <= imem06_in[83:80];
    19: reg_0007 <= imem02_in[7:4];
    21: reg_0007 <= imem02_in[7:4];
    86: reg_0007 <= imem03_in[71:68];
    88: reg_0007 <= imem03_in[71:68];
    96: reg_0007 <= imem06_in[83:80];
    endcase
  end

  // REG#8の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0008 <= imem03_in[75:72];
    7: reg_0008 <= imem03_in[75:72];
    9: reg_0008 <= imem02_in[83:80];
    11: reg_0008 <= imem02_in[83:80];
    13: reg_0008 <= imem04_in[103:100];
    15: reg_0008 <= imem03_in[75:72];
    17: reg_0008 <= imem06_in[91:88];
    19: reg_0008 <= imem06_in[91:88];
    21: reg_0008 <= imem04_in[103:100];
    23: reg_0008 <= imem06_in[91:88];
    25: reg_0008 <= imem03_in[75:72];
    27: reg_0008 <= imem04_in[103:100];
    29: reg_0008 <= imem04_in[103:100];
    31: reg_0008 <= imem06_in[91:88];
    33: reg_0008 <= imem00_in[111:108];
    35: reg_0008 <= imem03_in[75:72];
    37: reg_0008 <= imem06_in[91:88];
    58: reg_0008 <= imem06_in[91:88];
    83: reg_0008 <= imem04_in[103:100];
    endcase
  end

  // REG#9の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0009 <= imem03_in[103:100];
    7: reg_0009 <= imem00_in[63:60];
    9: reg_0009 <= imem03_in[103:100];
    11: reg_0009 <= imem03_in[111:108];
    13: reg_0009 <= imem04_in[115:112];
    15: reg_0009 <= imem00_in[63:60];
    17: reg_0009 <= imem03_in[103:100];
    19: reg_0009 <= imem04_in[115:112];
    43: reg_0009 <= imem03_in[103:100];
    45: reg_0009 <= imem03_in[103:100];
    47: reg_0009 <= imem03_in[3:0];
    49: reg_0009 <= imem03_in[111:108];
    51: reg_0009 <= imem03_in[111:108];
    53: reg_0009 <= imem03_in[3:0];
    56: reg_0009 <= imem00_in[63:60];
    58: reg_0009 <= imem00_in[63:60];
    60: reg_0009 <= imem00_in[95:92];
    62: reg_0009 <= imem04_in[115:112];
    64: reg_0009 <= imem04_in[115:112];
    66: reg_0009 <= imem00_in[95:92];
    68: reg_0009 <= imem03_in[3:0];
    70: reg_0009 <= imem00_in[95:92];
    72: reg_0009 <= imem03_in[103:100];
    74: reg_0009 <= imem00_in[95:92];
    76: reg_0009 <= imem03_in[103:100];
    78: reg_0009 <= imem03_in[103:100];
    80: reg_0009 <= imem00_in[63:60];
    82: reg_0009 <= imem00_in[63:60];
    84: reg_0009 <= imem00_in[63:60];
    86: reg_0009 <= imem03_in[3:0];
    88: reg_0009 <= imem03_in[3:0];
    91: reg_0009 <= imem00_in[63:60];
    endcase
  end

  // REG#10の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0010 <= imem03_in[107:104];
    7: reg_0010 <= imem03_in[107:104];
    9: reg_0010 <= imem03_in[107:104];
    11: reg_0010 <= imem04_in[43:40];
    13: reg_0010 <= imem05_in[15:12];
    15: reg_0010 <= imem04_in[43:40];
    17: reg_0010 <= imem04_in[43:40];
    19: reg_0010 <= imem03_in[107:104];
    21: reg_0010 <= imem03_in[107:104];
    23: reg_0010 <= imem04_in[43:40];
    25: reg_0010 <= imem05_in[15:12];
    27: reg_0010 <= imem03_in[107:104];
    29: reg_0010 <= imem04_in[43:40];
    31: reg_0010 <= imem05_in[15:12];
    33: reg_0010 <= imem04_in[43:40];
    35: reg_0010 <= imem03_in[107:104];
    37: reg_0010 <= imem03_in[107:104];
    39: reg_0010 <= imem05_in[15:12];
    41: reg_0010 <= imem04_in[43:40];
    43: reg_0010 <= imem03_in[107:104];
    45: reg_0010 <= imem07_in[43:40];
    47: reg_0010 <= imem06_in[7:4];
    49: reg_0010 <= imem06_in[7:4];
    51: reg_0010 <= imem03_in[107:104];
    53: reg_0010 <= imem07_in[43:40];
    55: reg_0010 <= imem06_in[7:4];
    57: reg_0010 <= imem06_in[7:4];
    96: reg_0010 <= imem07_in[43:40];
    endcase
  end

  // REG#11の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0011 <= imem06_in[107:104];
    7: reg_0011 <= imem00_in[95:92];
    9: reg_0011 <= imem06_in[107:104];
    32: reg_0011 <= imem06_in[107:104];
    38: reg_0011 <= imem06_in[107:104];
    40: reg_0011 <= imem06_in[107:104];
    42: reg_0011 <= imem07_in[83:80];
    44: reg_0011 <= imem00_in[63:60];
    46: reg_0011 <= imem00_in[63:60];
    48: reg_0011 <= imem07_in[83:80];
    50: reg_0011 <= imem00_in[63:60];
    52: reg_0011 <= imem07_in[83:80];
    54: reg_0011 <= imem00_in[63:60];
    56: reg_0011 <= imem00_in[95:92];
    58: reg_0011 <= imem06_in[107:104];
    86: reg_0011 <= imem06_in[107:104];
    endcase
  end

  // REG#12の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0012 <= imem03_in[19:16];
    7: reg_0012 <= imem00_in[123:120];
    9: reg_0012 <= imem00_in[123:120];
    11: reg_0012 <= imem00_in[123:120];
    13: reg_0012 <= imem00_in[123:120];
    15: reg_0012 <= imem03_in[19:16];
    17: reg_0012 <= imem03_in[19:16];
    19: reg_0012 <= imem00_in[123:120];
    21: reg_0012 <= imem04_in[59:56];
    23: reg_0012 <= imem03_in[19:16];
    25: reg_0012 <= imem03_in[19:16];
    27: reg_0012 <= imem03_in[19:16];
    30: reg_0012 <= imem00_in[27:24];
    32: reg_0012 <= imem00_in[27:24];
    34: reg_0012 <= imem04_in[59:56];
    36: reg_0012 <= imem07_in[47:44];
    38: reg_0012 <= imem00_in[27:24];
    40: reg_0012 <= imem00_in[27:24];
    42: reg_0012 <= imem00_in[27:24];
    44: reg_0012 <= imem00_in[123:120];
    46: reg_0012 <= imem00_in[123:120];
    48: reg_0012 <= imem04_in[59:56];
    51: reg_0012 <= imem04_in[59:56];
    53: reg_0012 <= imem07_in[47:44];
    55: reg_0012 <= imem03_in[19:16];
    88: reg_0012 <= imem00_in[123:120];
    90: reg_0012 <= imem04_in[59:56];
    92: reg_0012 <= imem04_in[59:56];
    94: reg_0012 <= imem07_in[47:44];
    96: reg_0012 <= imem04_in[59:56];
    endcase
  end

  // REG#13の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0013 <= imem03_in[43:40];
    7: reg_0013 <= imem01_in[3:0];
    9: reg_0013 <= imem03_in[43:40];
    11: reg_0013 <= imem01_in[3:0];
    25: reg_0013 <= imem01_in[3:0];
    48: reg_0013 <= imem03_in[43:40];
    50: reg_0013 <= imem01_in[3:0];
    52: reg_0013 <= imem01_in[3:0];
    54: reg_0013 <= imem03_in[43:40];
    56: reg_0013 <= imem03_in[43:40];
    58: reg_0013 <= imem01_in[3:0];
    60: reg_0013 <= imem01_in[3:0];
    62: reg_0013 <= imem03_in[43:40];
    64: reg_0013 <= imem05_in[99:96];
    66: reg_0013 <= imem01_in[3:0];
    68: reg_0013 <= imem05_in[99:96];
    73: reg_0013 <= imem05_in[99:96];
    endcase
  end

  // REG#14の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0014 <= imem03_in[67:64];
    7: reg_0014 <= imem02_in[39:36];
    9: reg_0014 <= imem02_in[39:36];
    11: reg_0014 <= imem04_in[59:56];
    13: reg_0014 <= imem02_in[39:36];
    15: reg_0014 <= imem02_in[39:36];
    17: reg_0014 <= imem02_in[39:36];
    19: reg_0014 <= imem04_in[59:56];
    42: reg_0014 <= imem04_in[59:56];
    endcase
  end

  // REG#15の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0015 <= imem03_in[83:80];
    7: reg_0015 <= imem04_in[123:120];
    9: reg_0015 <= imem03_in[83:80];
    11: reg_0015 <= imem04_in[83:80];
    13: reg_0015 <= imem03_in[83:80];
    15: reg_0015 <= imem03_in[83:80];
    17: reg_0015 <= imem03_in[83:80];
    19: reg_0015 <= imem04_in[123:120];
    38: reg_0015 <= imem04_in[123:120];
    40: reg_0015 <= imem03_in[83:80];
    42: reg_0015 <= imem04_in[83:80];
    97: reg_0015 <= imem03_in[83:80];
    endcase
  end

  // REG#16の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0016 <= imem03_in[91:88];
    7: reg_0016 <= imem03_in[91:88];
    9: reg_0016 <= imem02_in[95:92];
    11: reg_0016 <= imem04_in[119:116];
    13: reg_0016 <= imem04_in[119:116];
    15: reg_0016 <= imem03_in[11:8];
    17: reg_0016 <= imem03_in[91:88];
    19: reg_0016 <= imem03_in[11:8];
    21: reg_0016 <= imem02_in[95:92];
    81: reg_0016 <= imem03_in[11:8];
    83: reg_0016 <= imem04_in[119:116];
    97: reg_0016 <= imem02_in[95:92];
    endcase
  end

  // REG#17の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0017 <= imem06_in[55:52];
    7: reg_0017 <= imem06_in[55:52];
    9: reg_0017 <= imem06_in[55:52];
    33: reg_0017 <= imem06_in[55:52];
    35: reg_0017 <= imem07_in[67:64];
    37: reg_0017 <= imem06_in[55:52];
    61: reg_0017 <= imem07_in[67:64];
    63: reg_0017 <= imem07_in[67:64];
    65: reg_0017 <= imem06_in[55:52];
    67: reg_0017 <= imem06_in[55:52];
    69: reg_0017 <= imem07_in[67:64];
    71: reg_0017 <= imem06_in[55:52];
    89: reg_0017 <= imem07_in[67:64];
    91: reg_0017 <= imem07_in[67:64];
    93: reg_0017 <= imem06_in[55:52];
    95: reg_0017 <= imem04_in[79:76];
    endcase
  end

  // REG#18の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0018 <= imem06_in[75:72];
    7: reg_0018 <= imem06_in[75:72];
    9: reg_0018 <= imem06_in[75:72];
    30: reg_0018 <= imem01_in[87:84];
    32: reg_0018 <= imem06_in[75:72];
    38: reg_0018 <= imem01_in[87:84];
    40: reg_0018 <= imem03_in[7:4];
    42: reg_0018 <= imem00_in[79:76];
    44: reg_0018 <= imem03_in[7:4];
    46: reg_0018 <= imem01_in[87:84];
    48: reg_0018 <= imem01_in[99:96];
    50: reg_0018 <= imem06_in[75:72];
    52: reg_0018 <= imem01_in[87:84];
    55: reg_0018 <= imem01_in[99:96];
    57: reg_0018 <= imem01_in[99:96];
    59: reg_0018 <= imem06_in[75:72];
    61: reg_0018 <= imem01_in[87:84];
    63: reg_0018 <= imem01_in[87:84];
    65: reg_0018 <= imem01_in[87:84];
    67: reg_0018 <= imem00_in[79:76];
    69: reg_0018 <= imem03_in[7:4];
    71: reg_0018 <= imem06_in[75:72];
    87: reg_0018 <= imem00_in[79:76];
    89: reg_0018 <= imem06_in[75:72];
    endcase
  end

  // REG#19の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0019 <= imem03_in[11:8];
    7: reg_0019 <= imem05_in[7:4];
    9: reg_0019 <= imem03_in[11:8];
    11: reg_0019 <= imem05_in[7:4];
    14: reg_0019 <= imem03_in[11:8];
    16: reg_0019 <= imem05_in[7:4];
    18: reg_0019 <= imem03_in[11:8];
    20: reg_0019 <= imem03_in[11:8];
    22: reg_0019 <= imem05_in[7:4];
    24: reg_0019 <= imem03_in[11:8];
    26: reg_0019 <= imem03_in[51:48];
    28: reg_0019 <= imem05_in[7:4];
    30: reg_0019 <= imem03_in[51:48];
    32: reg_0019 <= imem03_in[51:48];
    34: reg_0019 <= imem03_in[51:48];
    36: reg_0019 <= imem03_in[51:48];
    38: reg_0019 <= imem05_in[7:4];
    40: reg_0019 <= imem05_in[7:4];
    42: reg_0019 <= imem03_in[11:8];
    44: reg_0019 <= imem03_in[51:48];
    46: reg_0019 <= imem05_in[7:4];
    48: reg_0019 <= imem05_in[7:4];
    50: reg_0019 <= imem05_in[7:4];
    65: reg_0019 <= imem03_in[11:8];
    67: reg_0019 <= imem03_in[51:48];
    69: reg_0019 <= imem03_in[11:8];
    72: reg_0019 <= imem05_in[7:4];
    74: reg_0019 <= imem05_in[7:4];
    endcase
  end

  // REG#20の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0020 <= imem06_in[59:56];
    8: reg_0020 <= imem06_in[59:56];
    11: reg_0020 <= imem06_in[59:56];
    13: reg_0020 <= imem05_in[39:36];
    15: reg_0020 <= imem05_in[39:36];
    17: reg_0020 <= imem05_in[39:36];
    19: reg_0020 <= imem03_in[15:12];
    21: reg_0020 <= imem05_in[7:4];
    23: reg_0020 <= imem03_in[15:12];
    25: reg_0020 <= imem05_in[39:36];
    27: reg_0020 <= imem06_in[59:56];
    29: reg_0020 <= imem05_in[39:36];
    31: reg_0020 <= imem05_in[7:4];
    33: reg_0020 <= imem05_in[7:4];
    35: reg_0020 <= imem05_in[7:4];
    37: reg_0020 <= imem05_in[7:4];
    39: reg_0020 <= imem06_in[59:56];
    57: reg_0020 <= imem03_in[15:12];
    59: reg_0020 <= imem05_in[39:36];
    61: reg_0020 <= imem05_in[39:36];
    64: reg_0020 <= imem05_in[39:36];
    66: reg_0020 <= imem05_in[39:36];
    76: reg_0020 <= imem05_in[39:36];
    78: reg_0020 <= imem05_in[7:4];
    80: reg_0020 <= imem05_in[7:4];
    82: reg_0020 <= imem05_in[39:36];
    84: reg_0020 <= imem05_in[7:4];
    86: reg_0020 <= imem05_in[7:4];
    89: reg_0020 <= imem06_in[59:56];
    endcase
  end

  // REG#21の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0021 <= imem06_in[83:80];
    8: reg_0021 <= imem04_in[115:112];
    10: reg_0021 <= imem04_in[115:112];
    12: reg_0021 <= imem06_in[83:80];
    14: reg_0021 <= imem07_in[3:0];
    16: reg_0021 <= imem04_in[115:112];
    18: reg_0021 <= imem04_in[115:112];
    43: reg_0021 <= imem06_in[83:80];
    45: reg_0021 <= imem06_in[83:80];
    47: reg_0021 <= imem06_in[83:80];
    49: reg_0021 <= imem06_in[83:80];
    51: reg_0021 <= imem04_in[115:112];
    53: reg_0021 <= imem06_in[83:80];
    55: reg_0021 <= imem07_in[3:0];
    57: reg_0021 <= imem06_in[83:80];
    endcase
  end

  // REG#22の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0022 <= imem06_in[99:96];
    8: reg_0022 <= imem05_in[23:20];
    10: reg_0022 <= imem06_in[99:96];
    12: reg_0022 <= imem06_in[99:96];
    14: reg_0022 <= imem06_in[99:96];
    16: reg_0022 <= imem05_in[23:20];
    18: reg_0022 <= imem05_in[23:20];
    20: reg_0022 <= imem05_in[23:20];
    48: reg_0022 <= imem06_in[99:96];
    50: reg_0022 <= imem05_in[23:20];
    65: reg_0022 <= imem05_in[23:20];
    69: reg_0022 <= imem05_in[23:20];
    71: reg_0022 <= imem06_in[99:96];
    89: reg_0022 <= imem04_in[39:36];
    91: reg_0022 <= imem06_in[99:96];
    93: reg_0022 <= imem06_in[99:96];
    95: reg_0022 <= imem05_in[23:20];
    endcase
  end

  // REG#23の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0023 <= imem06_in[115:112];
    8: reg_0023 <= imem05_in[63:60];
    10: reg_0023 <= imem05_in[63:60];
    12: reg_0023 <= imem06_in[115:112];
    14: reg_0023 <= imem06_in[115:112];
    16: reg_0023 <= imem06_in[115:112];
    18: reg_0023 <= imem05_in[63:60];
    20: reg_0023 <= imem06_in[115:112];
    22: reg_0023 <= imem06_in[123:120];
    24: reg_0023 <= imem05_in[63:60];
    26: reg_0023 <= imem06_in[115:112];
    28: reg_0023 <= imem05_in[63:60];
    30: reg_0023 <= imem02_in[43:40];
    32: reg_0023 <= imem05_in[63:60];
    34: reg_0023 <= imem00_in[127:124];
    36: reg_0023 <= imem05_in[63:60];
    38: reg_0023 <= imem02_in[43:40];
    40: reg_0023 <= imem00_in[127:124];
    42: reg_0023 <= imem00_in[127:124];
    44: reg_0023 <= imem02_in[43:40];
    46: reg_0023 <= imem06_in[115:112];
    48: reg_0023 <= imem06_in[115:112];
    50: reg_0023 <= imem05_in[63:60];
    65: reg_0023 <= imem06_in[115:112];
    67: reg_0023 <= imem00_in[127:124];
    69: reg_0023 <= imem02_in[43:40];
    71: reg_0023 <= imem00_in[127:124];
    73: reg_0023 <= imem06_in[123:120];
    75: reg_0023 <= imem06_in[115:112];
    77: reg_0023 <= imem06_in[115:112];
    79: reg_0023 <= imem06_in[115:112];
    81: reg_0023 <= imem05_in[63:60];
    83: reg_0023 <= imem06_in[115:112];
    85: reg_0023 <= imem05_in[63:60];
    87: reg_0023 <= imem05_in[63:60];
    endcase
  end

  // REG#24の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0024 <= imem06_in[87:84];
    8: reg_0024 <= imem05_in[75:72];
    10: reg_0024 <= imem05_in[75:72];
    12: reg_0024 <= imem05_in[75:72];
    17: reg_0024 <= imem07_in[115:112];
    19: reg_0024 <= imem07_in[115:112];
    21: reg_0024 <= imem05_in[75:72];
    23: reg_0024 <= imem01_in[63:60];
    25: reg_0024 <= imem05_in[75:72];
    27: reg_0024 <= imem05_in[75:72];
    29: reg_0024 <= imem05_in[75:72];
    31: reg_0024 <= imem05_in[75:72];
    33: reg_0024 <= imem06_in[87:84];
    35: reg_0024 <= imem05_in[75:72];
    37: reg_0024 <= imem05_in[75:72];
    39: reg_0024 <= imem05_in[75:72];
    41: reg_0024 <= imem06_in[87:84];
    43: reg_0024 <= imem07_in[115:112];
    endcase
  end

  // REG#25の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0025 <= imem06_in[67:64];
    9: reg_0025 <= imem06_in[67:64];
    32: reg_0025 <= imem06_in[67:64];
    37: reg_0025 <= imem06_in[67:64];
    57: reg_0025 <= imem06_in[67:64];
    endcase
  end

  // REG#26の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0026 <= imem06_in[23:20];
    9: reg_0026 <= imem06_in[23:20];
    32: reg_0026 <= imem06_in[23:20];
    35: reg_0026 <= imem06_in[23:20];
    38: reg_0026 <= imem06_in[23:20];
    41: reg_0026 <= imem02_in[79:76];
    43: reg_0026 <= imem02_in[79:76];
    45: reg_0026 <= imem02_in[79:76];
    60: reg_0026 <= imem02_in[79:76];
    62: reg_0026 <= imem02_in[79:76];
    65: reg_0026 <= imem06_in[23:20];
    67: reg_0026 <= imem07_in[103:100];
    69: reg_0026 <= imem07_in[103:100];
    71: reg_0026 <= imem06_in[23:20];
    90: reg_0026 <= imem06_in[23:20];
    92: reg_0026 <= imem02_in[79:76];
    94: reg_0026 <= imem02_in[79:76];
    96: reg_0026 <= imem02_in[79:76];
    endcase
  end

  // REG#27の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0027 <= imem06_in[19:16];
    9: reg_0027 <= imem06_in[19:16];
    32: reg_0027 <= imem07_in[39:36];
    34: reg_0027 <= imem07_in[39:36];
    36: reg_0027 <= imem06_in[19:16];
    40: reg_0027 <= imem04_in[47:44];
    42: reg_0027 <= imem07_in[39:36];
    45: reg_0027 <= imem06_in[19:16];
    47: reg_0027 <= imem06_in[19:16];
    49: reg_0027 <= imem04_in[47:44];
    59: reg_0027 <= imem04_in[47:44];
    endcase
  end

  // REG#28の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0028 <= imem06_in[7:4];
    10: reg_0028 <= imem06_in[7:4];
    12: reg_0028 <= imem06_in[7:4];
    14: reg_0028 <= imem00_in[15:12];
    16: reg_0028 <= imem06_in[7:4];
    18: reg_0028 <= imem00_in[15:12];
    20: reg_0028 <= imem06_in[7:4];
    22: reg_0028 <= imem07_in[15:12];
    24: reg_0028 <= imem06_in[7:4];
    26: reg_0028 <= imem06_in[7:4];
    28: reg_0028 <= imem00_in[15:12];
    30: reg_0028 <= imem06_in[7:4];
    32: reg_0028 <= imem07_in[15:12];
    34: reg_0028 <= imem06_in[7:4];
    36: reg_0028 <= imem07_in[15:12];
    38: reg_0028 <= imem00_in[3:0];
    40: reg_0028 <= imem07_in[99:96];
    42: reg_0028 <= imem07_in[15:12];
    44: reg_0028 <= imem00_in[3:0];
    46: reg_0028 <= imem06_in[7:4];
    48: reg_0028 <= imem06_in[7:4];
    50: reg_0028 <= imem00_in[87:84];
    52: reg_0028 <= imem06_in[7:4];
    54: reg_0028 <= imem00_in[15:12];
    56: reg_0028 <= imem07_in[99:96];
    58: reg_0028 <= imem06_in[7:4];
    87: reg_0028 <= imem07_in[15:12];
    89: reg_0028 <= imem00_in[15:12];
    91: reg_0028 <= imem00_in[87:84];
    endcase
  end

  // REG#29の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0029 <= imem06_in[95:92];
    10: reg_0029 <= imem06_in[95:92];
    12: reg_0029 <= imem06_in[119:116];
    14: reg_0029 <= imem00_in[51:48];
    16: reg_0029 <= imem06_in[95:92];
    18: reg_0029 <= imem06_in[119:116];
    20: reg_0029 <= imem06_in[119:116];
    22: reg_0029 <= imem06_in[95:92];
    24: reg_0029 <= imem06_in[95:92];
    26: reg_0029 <= imem06_in[119:116];
    28: reg_0029 <= imem06_in[95:92];
    30: reg_0029 <= imem06_in[95:92];
    32: reg_0029 <= imem06_in[95:92];
    37: reg_0029 <= imem06_in[95:92];
    62: reg_0029 <= imem06_in[119:116];
    64: reg_0029 <= imem07_in[63:60];
    66: reg_0029 <= imem06_in[119:116];
    68: reg_0029 <= imem06_in[119:116];
    70: reg_0029 <= imem00_in[51:48];
    72: reg_0029 <= imem06_in[95:92];
    74: reg_0029 <= imem06_in[95:92];
    76: reg_0029 <= imem06_in[95:92];
    78: reg_0029 <= imem06_in[119:116];
    80: reg_0029 <= imem00_in[7:4];
    82: reg_0029 <= imem06_in[119:116];
    84: reg_0029 <= imem00_in[7:4];
    86: reg_0029 <= imem06_in[95:92];
    endcase
  end

  // REG#30の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0030 <= imem06_in[91:88];
    10: reg_0030 <= imem02_in[3:0];
    12: reg_0030 <= imem02_in[3:0];
    14: reg_0030 <= imem02_in[3:0];
    16: reg_0030 <= imem00_in[107:104];
    18: reg_0030 <= imem05_in[59:56];
    20: reg_0030 <= imem06_in[91:88];
    22: reg_0030 <= imem02_in[3:0];
    24: reg_0030 <= imem05_in[59:56];
    26: reg_0030 <= imem05_in[59:56];
    28: reg_0030 <= imem05_in[59:56];
    30: reg_0030 <= imem00_in[107:104];
    32: reg_0030 <= imem06_in[91:88];
    35: reg_0030 <= imem02_in[3:0];
    37: reg_0030 <= imem00_in[107:104];
    39: reg_0030 <= imem02_in[3:0];
    41: reg_0030 <= imem06_in[91:88];
    43: reg_0030 <= imem02_in[3:0];
    45: reg_0030 <= imem00_in[107:104];
    47: reg_0030 <= imem00_in[107:104];
    49: reg_0030 <= imem06_in[51:48];
    51: reg_0030 <= imem05_in[71:68];
    53: reg_0030 <= imem00_in[107:104];
    55: reg_0030 <= imem02_in[3:0];
    57: reg_0030 <= imem02_in[3:0];
    59: reg_0030 <= imem00_in[107:104];
    61: reg_0030 <= imem05_in[71:68];
    66: reg_0030 <= imem06_in[91:88];
    68: reg_0030 <= imem05_in[71:68];
    73: reg_0030 <= imem06_in[51:48];
    75: reg_0030 <= imem05_in[59:56];
    77: reg_0030 <= imem02_in[3:0];
    79: reg_0030 <= imem06_in[91:88];
    81: reg_0030 <= imem05_in[59:56];
    83: reg_0030 <= imem06_in[91:88];
    85: reg_0030 <= imem06_in[91:88];
    87: reg_0030 <= imem02_in[3:0];
    89: reg_0030 <= imem02_in[3:0];
    91: reg_0030 <= imem00_in[107:104];
    endcase
  end

  // REG#31の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0031 <= imem06_in[15:12];
    10: reg_0031 <= imem06_in[15:12];
    12: reg_0031 <= imem07_in[99:96];
    14: reg_0031 <= imem07_in[99:96];
    16: reg_0031 <= imem06_in[15:12];
    18: reg_0031 <= imem07_in[99:96];
    20: reg_0031 <= imem06_in[15:12];
    22: reg_0031 <= imem02_in[95:92];
    24: reg_0031 <= imem07_in[99:96];
    26: reg_0031 <= imem07_in[99:96];
    28: reg_0031 <= imem04_in[107:104];
    30: reg_0031 <= imem07_in[99:96];
    32: reg_0031 <= imem06_in[15:12];
    36: reg_0031 <= imem02_in[95:92];
    38: reg_0031 <= imem07_in[99:96];
    40: reg_0031 <= imem02_in[95:92];
    42: reg_0031 <= imem06_in[15:12];
    44: reg_0031 <= imem02_in[95:92];
    46: reg_0031 <= imem04_in[107:104];
    49: reg_0031 <= imem04_in[107:104];
    60: reg_0031 <= imem04_in[119:116];
    62: reg_0031 <= imem04_in[119:116];
    64: reg_0031 <= imem07_in[95:92];
    66: reg_0031 <= imem02_in[95:92];
    68: reg_0031 <= imem07_in[95:92];
    70: reg_0031 <= imem04_in[119:116];
    72: reg_0031 <= imem07_in[99:96];
    74: reg_0031 <= imem04_in[119:116];
    76: reg_0031 <= imem04_in[107:104];
    78: reg_0031 <= imem04_in[107:104];
    80: reg_0031 <= imem07_in[99:96];
    83: reg_0031 <= imem04_in[107:104];
    endcase
  end

  // REG#32の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0032 <= imem06_in[35:32];
    10: reg_0032 <= imem02_in[19:16];
    12: reg_0032 <= imem02_in[19:16];
    14: reg_0032 <= imem00_in[91:88];
    16: reg_0032 <= imem00_in[91:88];
    18: reg_0032 <= imem02_in[19:16];
    20: reg_0032 <= imem00_in[91:88];
    22: reg_0032 <= imem06_in[35:32];
    24: reg_0032 <= imem05_in[31:28];
    26: reg_0032 <= imem05_in[31:28];
    28: reg_0032 <= imem05_in[31:28];
    30: reg_0032 <= imem06_in[35:32];
    32: reg_0032 <= imem06_in[35:32];
    38: reg_0032 <= imem02_in[19:16];
    40: reg_0032 <= imem02_in[19:16];
    42: reg_0032 <= imem02_in[19:16];
    44: reg_0032 <= imem00_in[91:88];
    46: reg_0032 <= imem00_in[91:88];
    48: reg_0032 <= imem05_in[31:28];
    50: reg_0032 <= imem05_in[31:28];
    67: reg_0032 <= imem05_in[31:28];
    69: reg_0032 <= imem05_in[31:28];
    71: reg_0032 <= imem06_in[35:32];
    88: reg_0032 <= imem06_in[35:32];
    90: reg_0032 <= imem00_in[91:88];
    92: reg_0032 <= imem02_in[19:16];
    94: reg_0032 <= imem06_in[35:32];
    96: reg_0032 <= imem05_in[31:28];
    endcase
  end

  // REG#33の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0033 <= imem06_in[3:0];
    10: reg_0033 <= imem06_in[3:0];
    12: reg_0033 <= imem06_in[3:0];
    14: reg_0033 <= imem00_in[111:108];
    16: reg_0033 <= imem00_in[115:112];
    18: reg_0033 <= imem00_in[51:48];
    20: reg_0033 <= imem07_in[83:80];
    22: reg_0033 <= imem00_in[51:48];
    24: reg_0033 <= imem00_in[51:48];
    26: reg_0033 <= imem03_in[79:76];
    28: reg_0033 <= imem07_in[83:80];
    30: reg_0033 <= imem02_in[123:120];
    32: reg_0033 <= imem00_in[111:108];
    34: reg_0033 <= imem02_in[123:120];
    36: reg_0033 <= imem00_in[115:112];
    38: reg_0033 <= imem00_in[51:48];
    40: reg_0033 <= imem00_in[51:48];
    42: reg_0033 <= imem06_in[3:0];
    44: reg_0033 <= imem00_in[51:48];
    46: reg_0033 <= imem00_in[111:108];
    48: reg_0033 <= imem03_in[67:64];
    50: reg_0033 <= imem00_in[51:48];
    52: reg_0033 <= imem00_in[51:48];
    54: reg_0033 <= imem00_in[111:108];
    56: reg_0033 <= imem02_in[123:120];
    58: reg_0033 <= imem02_in[123:120];
    60: reg_0033 <= imem00_in[51:48];
    62: reg_0033 <= imem00_in[115:112];
    64: reg_0033 <= imem03_in[79:76];
    66: reg_0033 <= imem00_in[115:112];
    68: reg_0033 <= imem00_in[115:112];
    70: reg_0033 <= imem00_in[111:108];
    72: reg_0033 <= imem03_in[79:76];
    74: reg_0033 <= imem00_in[51:48];
    76: reg_0033 <= imem02_in[123:120];
    78: reg_0033 <= imem00_in[115:112];
    80: reg_0033 <= imem02_in[123:120];
    82: reg_0033 <= imem03_in[79:76];
    84: reg_0033 <= imem07_in[83:80];
    86: reg_0033 <= imem00_in[111:108];
    88: reg_0033 <= imem03_in[79:76];
    endcase
  end

  // REG#34の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0034 <= imem06_in[39:36];
    10: reg_0034 <= imem06_in[39:36];
    12: reg_0034 <= imem01_in[31:28];
    14: reg_0034 <= imem06_in[39:36];
    16: reg_0034 <= imem06_in[39:36];
    18: reg_0034 <= imem06_in[39:36];
    20: reg_0034 <= imem06_in[39:36];
    22: reg_0034 <= imem01_in[31:28];
    24: reg_0034 <= imem05_in[95:92];
    26: reg_0034 <= imem01_in[31:28];
    28: reg_0034 <= imem01_in[31:28];
    30: reg_0034 <= imem01_in[31:28];
    32: reg_0034 <= imem01_in[31:28];
    34: reg_0034 <= imem06_in[39:36];
    36: reg_0034 <= imem06_in[39:36];
    40: reg_0034 <= imem01_in[55:52];
    42: reg_0034 <= imem01_in[55:52];
    44: reg_0034 <= imem02_in[91:88];
    46: reg_0034 <= imem06_in[39:36];
    48: reg_0034 <= imem01_in[55:52];
    50: reg_0034 <= imem01_in[55:52];
    52: reg_0034 <= imem05_in[95:92];
    54: reg_0034 <= imem01_in[55:52];
    56: reg_0034 <= imem02_in[91:88];
    58: reg_0034 <= imem01_in[31:28];
    60: reg_0034 <= imem01_in[55:52];
    62: reg_0034 <= imem02_in[91:88];
    64: reg_0034 <= imem06_in[39:36];
    66: reg_0034 <= imem02_in[91:88];
    68: reg_0034 <= imem06_in[39:36];
    70: reg_0034 <= imem01_in[55:52];
    72: reg_0034 <= imem02_in[91:88];
    83: reg_0034 <= imem06_in[39:36];
    85: reg_0034 <= imem06_in[39:36];
    87: reg_0034 <= imem02_in[91:88];
    89: reg_0034 <= imem06_in[39:36];
    94: reg_0034 <= imem01_in[31:28];
    96: reg_0034 <= imem06_in[39:36];
    endcase
  end

  // REG#35の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0035 <= imem06_in[43:40];
    10: reg_0035 <= imem02_in[59:56];
    12: reg_0035 <= imem06_in[43:40];
    14: reg_0035 <= imem02_in[27:24];
    16: reg_0035 <= imem02_in[59:56];
    18: reg_0035 <= imem02_in[27:24];
    20: reg_0035 <= imem06_in[43:40];
    22: reg_0035 <= imem03_in[43:40];
    24: reg_0035 <= imem02_in[27:24];
    26: reg_0035 <= imem03_in[43:40];
    28: reg_0035 <= imem06_in[43:40];
    30: reg_0035 <= imem02_in[27:24];
    32: reg_0035 <= imem03_in[43:40];
    34: reg_0035 <= imem06_in[43:40];
    36: reg_0035 <= imem03_in[43:40];
    38: reg_0035 <= imem03_in[43:40];
    40: reg_0035 <= imem03_in[43:40];
    42: reg_0035 <= imem05_in[79:76];
    44: reg_0035 <= imem02_in[27:24];
    47: reg_0035 <= imem02_in[59:56];
    49: reg_0035 <= imem03_in[43:40];
    51: reg_0035 <= imem02_in[59:56];
    54: reg_0035 <= imem04_in[31:28];
    56: reg_0035 <= imem05_in[79:76];
    62: reg_0035 <= imem02_in[27:24];
    65: reg_0035 <= imem03_in[43:40];
    67: reg_0035 <= imem03_in[43:40];
    69: reg_0035 <= imem02_in[59:56];
    71: reg_0035 <= imem04_in[31:28];
    73: reg_0035 <= imem02_in[59:56];
    75: reg_0035 <= imem02_in[59:56];
    77: reg_0035 <= imem04_in[31:28];
    79: reg_0035 <= imem02_in[27:24];
    81: reg_0035 <= imem02_in[59:56];
    83: reg_0035 <= imem03_in[43:40];
    85: reg_0035 <= imem03_in[43:40];
    87: reg_0035 <= imem02_in[59:56];
    89: reg_0035 <= imem02_in[59:56];
    91: reg_0035 <= imem07_in[3:0];
    93: reg_0035 <= imem03_in[43:40];
    95: reg_0035 <= imem07_in[23:20];
    97: reg_0035 <= imem04_in[31:28];
    endcase
  end

  // REG#36の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0036 <= imem06_in[71:68];
    10: reg_0036 <= imem06_in[71:68];
    12: reg_0036 <= imem06_in[71:68];
    14: reg_0036 <= imem06_in[71:68];
    16: reg_0036 <= imem02_in[79:76];
    18: reg_0036 <= imem06_in[71:68];
    20: reg_0036 <= imem06_in[71:68];
    22: reg_0036 <= imem02_in[79:76];
    24: reg_0036 <= imem02_in[79:76];
    26: reg_0036 <= imem06_in[71:68];
    28: reg_0036 <= imem06_in[71:68];
    31: reg_0036 <= imem02_in[79:76];
    33: reg_0036 <= imem02_in[75:72];
    35: reg_0036 <= imem06_in[71:68];
    38: reg_0036 <= imem00_in[31:28];
    40: reg_0036 <= imem06_in[71:68];
    42: reg_0036 <= imem06_in[71:68];
    44: reg_0036 <= imem02_in[79:76];
    47: reg_0036 <= imem00_in[31:28];
    49: reg_0036 <= imem06_in[71:68];
    51: reg_0036 <= imem06_in[71:68];
    53: reg_0036 <= imem00_in[31:28];
    55: reg_0036 <= imem02_in[79:76];
    57: reg_0036 <= imem02_in[75:72];
    59: reg_0036 <= imem00_in[31:28];
    61: reg_0036 <= imem02_in[79:76];
    63: reg_0036 <= imem02_in[75:72];
    73: reg_0036 <= imem00_in[31:28];
    75: reg_0036 <= imem00_in[31:28];
    77: reg_0036 <= imem02_in[75:72];
    79: reg_0036 <= imem02_in[75:72];
    81: reg_0036 <= imem00_in[31:28];
    83: reg_0036 <= imem00_in[31:28];
    85: reg_0036 <= imem00_in[31:28];
    87: reg_0036 <= imem02_in[75:72];
    89: reg_0036 <= imem06_in[71:68];
    endcase
  end

  // REG#37の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0037 <= imem06_in[79:76];
    10: reg_0037 <= imem02_in[103:100];
    12: reg_0037 <= imem06_in[79:76];
    14: reg_0037 <= imem02_in[103:100];
    16: reg_0037 <= imem06_in[79:76];
    18: reg_0037 <= imem02_in[103:100];
    20: reg_0037 <= imem00_in[55:52];
    22: reg_0037 <= imem00_in[55:52];
    24: reg_0037 <= imem02_in[103:100];
    26: reg_0037 <= imem02_in[103:100];
    43: reg_0037 <= imem01_in[31:28];
    45: reg_0037 <= imem06_in[79:76];
    47: reg_0037 <= imem01_in[31:28];
    50: reg_0037 <= imem06_in[79:76];
    52: reg_0037 <= imem02_in[103:100];
    endcase
  end

  // REG#38の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0038 <= imem06_in[111:108];
    10: reg_0038 <= imem03_in[39:36];
    12: reg_0038 <= imem06_in[111:108];
    14: reg_0038 <= imem06_in[111:108];
    16: reg_0038 <= imem03_in[39:36];
    18: reg_0038 <= imem03_in[39:36];
    20: reg_0038 <= imem03_in[39:36];
    22: reg_0038 <= imem06_in[111:108];
    24: reg_0038 <= imem07_in[11:8];
    26: reg_0038 <= imem03_in[39:36];
    28: reg_0038 <= imem03_in[39:36];
    70: reg_0038 <= imem03_in[39:36];
    97: reg_0038 <= imem03_in[39:36];
    endcase
  end

  // REG#39の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0039 <= imem06_in[11:8];
    10: reg_0039 <= imem06_in[11:8];
    12: reg_0039 <= imem02_in[39:36];
    14: reg_0039 <= imem06_in[11:8];
    16: reg_0039 <= imem02_in[39:36];
    18: reg_0039 <= imem01_in[75:72];
    20: reg_0039 <= imem01_in[75:72];
    22: reg_0039 <= imem01_in[75:72];
    24: reg_0039 <= imem02_in[39:36];
    26: reg_0039 <= imem02_in[39:36];
    52: reg_0039 <= imem02_in[39:36];
    endcase
  end

  // REG#40の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0040 <= imem06_in[51:48];
    10: reg_0040 <= imem03_in[47:44];
    12: reg_0040 <= imem06_in[51:48];
    14: reg_0040 <= imem06_in[51:48];
    16: reg_0040 <= imem05_in[19:16];
    18: reg_0040 <= imem02_in[119:116];
    20: reg_0040 <= imem03_in[47:44];
    22: reg_0040 <= imem03_in[47:44];
    24: reg_0040 <= imem05_in[19:16];
    26: reg_0040 <= imem03_in[47:44];
    28: reg_0040 <= imem03_in[47:44];
    70: reg_0040 <= imem03_in[47:44];
    89: reg_0040 <= imem06_in[51:48];
    endcase
  end

  // REG#41の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0041 <= imem04_in[31:28];
    11: reg_0041 <= imem04_in[127:124];
    13: reg_0041 <= imem04_in[127:124];
    15: reg_0041 <= imem04_in[83:80];
    17: reg_0041 <= imem04_in[83:80];
    21: reg_0041 <= imem04_in[83:80];
    23: reg_0041 <= imem04_in[127:124];
    25: reg_0041 <= imem04_in[83:80];
    27: reg_0041 <= imem04_in[127:124];
    29: reg_0041 <= imem04_in[31:28];
    31: reg_0041 <= imem04_in[83:80];
    33: reg_0041 <= imem04_in[31:28];
    35: reg_0041 <= imem04_in[83:80];
    37: reg_0041 <= imem04_in[31:28];
    39: reg_0041 <= imem04_in[127:124];
    41: reg_0041 <= imem04_in[83:80];
    43: reg_0041 <= imem04_in[127:124];
    45: reg_0041 <= imem04_in[31:28];
    47: reg_0041 <= imem04_in[127:124];
    49: reg_0041 <= imem04_in[83:80];
    57: reg_0041 <= imem04_in[127:124];
    59: reg_0041 <= imem04_in[31:28];
    endcase
  end

  // REG#42の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0042 <= imem02_in[15:12];
    13: reg_0042 <= imem06_in[39:36];
    15: reg_0042 <= imem06_in[39:36];
    17: reg_0042 <= imem01_in[11:8];
    19: reg_0042 <= imem01_in[11:8];
    21: reg_0042 <= imem06_in[39:36];
    23: reg_0042 <= imem02_in[127:124];
    25: reg_0042 <= imem06_in[39:36];
    27: reg_0042 <= imem06_in[39:36];
    29: reg_0042 <= imem06_in[39:36];
    57: reg_0042 <= imem01_in[11:8];
    59: reg_0042 <= imem05_in[3:0];
    61: reg_0042 <= imem05_in[3:0];
    66: reg_0042 <= imem02_in[15:12];
    68: reg_0042 <= imem02_in[15:12];
    70: reg_0042 <= imem01_in[11:8];
    72: reg_0042 <= imem05_in[3:0];
    76: reg_0042 <= imem05_in[3:0];
    78: reg_0042 <= imem06_in[39:36];
    80: reg_0042 <= imem06_in[39:36];
    82: reg_0042 <= imem02_in[127:124];
    84: reg_0042 <= imem01_in[11:8];
    86: reg_0042 <= imem01_in[11:8];
    88: reg_0042 <= imem06_in[39:36];
    91: reg_0042 <= imem04_in[91:88];
    93: reg_0042 <= imem04_in[91:88];
    95: reg_0042 <= imem01_in[11:8];
    97: reg_0042 <= imem06_in[39:36];
    endcase
  end

  // REG#43の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0043 <= imem04_in[59:56];
    14: reg_0043 <= imem03_in[55:52];
    16: reg_0043 <= imem03_in[55:52];
    18: reg_0043 <= imem04_in[59:56];
    47: reg_0043 <= imem03_in[55:52];
    49: reg_0043 <= imem04_in[59:56];
    56: reg_0043 <= imem03_in[55:52];
    58: reg_0043 <= imem04_in[59:56];
    60: reg_0043 <= imem04_in[59:56];
    62: reg_0043 <= imem04_in[59:56];
    64: reg_0043 <= imem02_in[47:44];
    66: reg_0043 <= imem04_in[79:76];
    68: reg_0043 <= imem02_in[47:44];
    70: reg_0043 <= imem04_in[59:56];
    72: reg_0043 <= imem04_in[59:56];
    74: reg_0043 <= imem02_in[47:44];
    76: reg_0043 <= imem01_in[63:60];
    78: reg_0043 <= imem02_in[47:44];
    80: reg_0043 <= imem02_in[47:44];
    82: reg_0043 <= imem01_in[63:60];
    84: reg_0043 <= imem01_in[63:60];
    86: reg_0043 <= imem07_in[47:44];
    88: reg_0043 <= imem04_in[79:76];
    90: reg_0043 <= imem04_in[79:76];
    92: reg_0043 <= imem07_in[47:44];
    94: reg_0043 <= imem02_in[47:44];
    96: reg_0043 <= imem04_in[79:76];
    endcase
  end

  // REG#44の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0044 <= imem04_in[111:108];
    14: reg_0044 <= imem04_in[111:108];
    16: reg_0044 <= imem05_in[87:84];
    18: reg_0044 <= imem04_in[111:108];
    47: reg_0044 <= imem07_in[75:72];
    49: reg_0044 <= imem07_in[75:72];
    51: reg_0044 <= imem05_in[87:84];
    53: reg_0044 <= imem04_in[111:108];
    55: reg_0044 <= imem05_in[87:84];
    57: reg_0044 <= imem04_in[111:108];
    59: reg_0044 <= imem04_in[111:108];
    97: reg_0044 <= imem04_in[111:108];
    endcase
  end

  // REG#45の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0045 <= imem02_in[11:8];
    14: reg_0045 <= imem02_in[11:8];
    16: reg_0045 <= imem02_in[11:8];
    18: reg_0045 <= imem03_in[63:60];
    20: reg_0045 <= imem01_in[51:48];
    22: reg_0045 <= imem02_in[11:8];
    24: reg_0045 <= imem02_in[11:8];
    26: reg_0045 <= imem02_in[11:8];
    52: reg_0045 <= imem03_in[63:60];
    54: reg_0045 <= imem02_in[11:8];
    56: reg_0045 <= imem05_in[19:16];
    58: reg_0045 <= imem01_in[119:116];
    60: reg_0045 <= imem01_in[119:116];
    62: reg_0045 <= imem03_in[63:60];
    64: reg_0045 <= imem05_in[19:16];
    66: reg_0045 <= imem02_in[11:8];
    68: reg_0045 <= imem01_in[119:116];
    71: reg_0045 <= imem01_in[51:48];
    73: reg_0045 <= imem01_in[119:116];
    75: reg_0045 <= imem01_in[119:116];
    77: reg_0045 <= imem01_in[119:116];
    79: reg_0045 <= imem02_in[11:8];
    81: reg_0045 <= imem01_in[51:48];
    83: reg_0045 <= imem01_in[51:48];
    85: reg_0045 <= imem02_in[11:8];
    97: reg_0045 <= imem01_in[119:116];
    endcase
  end

  // REG#46の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0046 <= imem04_in[11:8];
    15: reg_0046 <= imem06_in[7:4];
    17: reg_0046 <= imem04_in[11:8];
    20: reg_0046 <= imem04_in[11:8];
    22: reg_0046 <= imem04_in[11:8];
    25: reg_0046 <= imem03_in[91:88];
    27: reg_0046 <= imem03_in[91:88];
    29: reg_0046 <= imem04_in[11:8];
    31: reg_0046 <= imem03_in[91:88];
    55: reg_0046 <= imem03_in[91:88];
    88: reg_0046 <= imem06_in[7:4];
    91: reg_0046 <= imem03_in[91:88];
    93: reg_0046 <= imem04_in[11:8];
    95: reg_0046 <= imem03_in[91:88];
    97: reg_0046 <= imem06_in[7:4];
    endcase
  end

  // REG#47の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0047 <= imem04_in[19:16];
    16: reg_0047 <= imem07_in[47:44];
    18: reg_0047 <= imem04_in[19:16];
    43: reg_0047 <= imem07_in[47:44];
    endcase
  end

  // REG#48の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0048 <= imem04_in[71:68];
    17: reg_0048 <= imem04_in[71:68];
    21: reg_0048 <= imem04_in[71:68];
    24: reg_0048 <= imem04_in[71:68];
    83: reg_0048 <= imem04_in[71:68];
    endcase
  end

  // REG#49の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0049 <= imem02_in[75:72];
    17: reg_0049 <= imem02_in[75:72];
    19: reg_0049 <= imem03_in[59:56];
    21: reg_0049 <= imem02_in[75:72];
    86: reg_0049 <= imem03_in[23:20];
    88: reg_0049 <= imem03_in[59:56];
    endcase
  end

  // REG#50の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0050 <= imem04_in[115:112];
    17: reg_0050 <= imem04_in[115:112];
    20: reg_0050 <= imem04_in[115:112];
    22: reg_0050 <= imem03_in[51:48];
    24: reg_0050 <= imem04_in[115:112];
    81: reg_0050 <= imem05_in[123:120];
    83: reg_0050 <= imem05_in[123:120];
    85: reg_0050 <= imem04_in[115:112];
    87: reg_0050 <= imem03_in[51:48];
    90: reg_0050 <= imem03_in[51:48];
    94: reg_0050 <= imem04_in[127:124];
    96: reg_0050 <= imem04_in[71:68];
    endcase
  end

  // REG#51の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0051 <= imem02_in[63:60];
    18: reg_0051 <= imem02_in[67:64];
    20: reg_0051 <= imem03_in[71:68];
    22: reg_0051 <= imem02_in[63:60];
    24: reg_0051 <= imem02_in[67:64];
    26: reg_0051 <= imem03_in[71:68];
    28: reg_0051 <= imem03_in[71:68];
    68: reg_0051 <= imem03_in[71:68];
    70: reg_0051 <= imem03_in[71:68];
    endcase
  end

  // REG#52の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0052 <= imem02_in[51:48];
    18: reg_0052 <= imem02_in[51:48];
    20: reg_0052 <= imem02_in[51:48];
    23: reg_0052 <= imem02_in[51:48];
    25: reg_0052 <= imem02_in[51:48];
    28: reg_0052 <= imem02_in[51:48];
    30: reg_0052 <= imem07_in[27:24];
    32: reg_0052 <= imem02_in[51:48];
    34: reg_0052 <= imem07_in[27:24];
    36: reg_0052 <= imem00_in[119:116];
    38: reg_0052 <= imem02_in[51:48];
    40: reg_0052 <= imem02_in[51:48];
    42: reg_0052 <= imem07_in[27:24];
    44: reg_0052 <= imem02_in[51:48];
    46: reg_0052 <= imem03_in[99:96];
    48: reg_0052 <= imem03_in[99:96];
    50: reg_0052 <= imem02_in[51:48];
    52: reg_0052 <= imem02_in[51:48];
    endcase
  end

  // REG#53の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0053 <= imem04_in[63:60];
    18: reg_0053 <= imem04_in[63:60];
    45: reg_0053 <= imem04_in[63:60];
    47: reg_0053 <= imem07_in[119:116];
    49: reg_0053 <= imem04_in[63:60];
    60: reg_0053 <= imem07_in[119:116];
    62: reg_0053 <= imem04_in[63:60];
    64: reg_0053 <= imem04_in[55:52];
    66: reg_0053 <= imem06_in[75:72];
    68: reg_0053 <= imem06_in[75:72];
    70: reg_0053 <= imem04_in[63:60];
    72: reg_0053 <= imem04_in[55:52];
    74: reg_0053 <= imem07_in[119:116];
    76: reg_0053 <= imem07_in[119:116];
    78: reg_0053 <= imem03_in[23:20];
    80: reg_0053 <= imem06_in[75:72];
    82: reg_0053 <= imem04_in[55:52];
    85: reg_0053 <= imem06_in[75:72];
    88: reg_0053 <= imem06_in[75:72];
    90: reg_0053 <= imem06_in[75:72];
    92: reg_0053 <= imem07_in[119:116];
    94: reg_0053 <= imem07_in[119:116];
    96: reg_0053 <= imem04_in[55:52];
    endcase
  end

  // REG#54の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0054 <= imem04_in[15:12];
    18: reg_0054 <= imem04_in[15:12];
    46: reg_0054 <= imem04_in[15:12];
    50: reg_0054 <= imem02_in[119:116];
    52: reg_0054 <= imem02_in[119:116];
    endcase
  end

  // REG#55の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0055 <= imem02_in[87:84];
    18: reg_0055 <= imem02_in[87:84];
    20: reg_0055 <= imem04_in[67:64];
    22: reg_0055 <= imem04_in[67:64];
    24: reg_0055 <= imem04_in[67:64];
    84: reg_0055 <= imem02_in[87:84];
    96: reg_0055 <= imem02_in[87:84];
    endcase
  end

  // REG#56の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0056 <= imem04_in[55:52];
    18: reg_0056 <= imem04_in[55:52];
    40: reg_0056 <= imem04_in[55:52];
    42: reg_0056 <= imem04_in[55:52];
    endcase
  end

  // REG#57の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0057 <= imem04_in[87:84];
    18: reg_0057 <= imem04_in[87:84];
    46: reg_0057 <= imem04_in[87:84];
    50: reg_0057 <= imem04_in[87:84];
    52: reg_0057 <= imem04_in[87:84];
    54: reg_0057 <= imem05_in[127:124];
    56: reg_0057 <= imem05_in[127:124];
    61: reg_0057 <= imem04_in[87:84];
    63: reg_0057 <= imem04_in[87:84];
    65: reg_0057 <= imem04_in[87:84];
    67: reg_0057 <= imem04_in[87:84];
    69: reg_0057 <= imem04_in[87:84];
    71: reg_0057 <= imem05_in[127:124];
    73: reg_0057 <= imem05_in[127:124];
    endcase
  end

  // REG#58の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0058 <= imem04_in[39:36];
    18: reg_0058 <= imem04_in[39:36];
    40: reg_0058 <= imem04_in[39:36];
    42: reg_0058 <= imem04_in[39:36];
    endcase
  end

  // REG#59の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0059 <= imem04_in[3:0];
    18: reg_0059 <= imem04_in[3:0];
    47: reg_0059 <= imem04_in[3:0];
    49: reg_0059 <= imem04_in[3:0];
    56: reg_0059 <= imem01_in[87:84];
    58: reg_0059 <= imem01_in[87:84];
    60: reg_0059 <= imem01_in[87:84];
    62: reg_0059 <= imem04_in[99:96];
    64: reg_0059 <= imem04_in[111:108];
    66: reg_0059 <= imem04_in[3:0];
    68: reg_0059 <= imem04_in[3:0];
    70: reg_0059 <= imem04_in[3:0];
    72: reg_0059 <= imem01_in[87:84];
    74: reg_0059 <= imem04_in[99:96];
    76: reg_0059 <= imem02_in[107:104];
    78: reg_0059 <= imem04_in[3:0];
    80: reg_0059 <= imem04_in[99:96];
    82: reg_0059 <= imem04_in[3:0];
    84: reg_0059 <= imem04_in[111:108];
    86: reg_0059 <= imem04_in[99:96];
    88: reg_0059 <= imem01_in[87:84];
    90: reg_0059 <= imem04_in[3:0];
    92: reg_0059 <= imem02_in[107:104];
    94: reg_0059 <= imem01_in[87:84];
    97: reg_0059 <= imem01_in[87:84];
    endcase
  end

  // REG#60の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0060 <= imem02_in[91:88];
    18: reg_0060 <= imem02_in[91:88];
    20: reg_0060 <= imem04_in[91:88];
    22: reg_0060 <= imem04_in[91:88];
    25: reg_0060 <= imem04_in[91:88];
    27: reg_0060 <= imem00_in[31:28];
    29: reg_0060 <= imem02_in[91:88];
    31: reg_0060 <= imem02_in[91:88];
    33: reg_0060 <= imem03_in[3:0];
    35: reg_0060 <= imem00_in[31:28];
    37: reg_0060 <= imem00_in[59:56];
    39: reg_0060 <= imem00_in[59:56];
    41: reg_0060 <= imem03_in[3:0];
    43: reg_0060 <= imem00_in[59:56];
    45: reg_0060 <= imem00_in[59:56];
    47: reg_0060 <= imem00_in[59:56];
    49: reg_0060 <= imem03_in[3:0];
    51: reg_0060 <= imem06_in[3:0];
    53: reg_0060 <= imem02_in[91:88];
    55: reg_0060 <= imem03_in[3:0];
    88: reg_0060 <= imem04_in[91:88];
    90: reg_0060 <= imem03_in[3:0];
    endcase
  end

  // REG#61の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0061 <= imem04_in[7:4];
    19: reg_0061 <= imem04_in[7:4];
    43: reg_0061 <= imem01_in[71:68];
    45: reg_0061 <= imem01_in[71:68];
    47: reg_0061 <= imem04_in[7:4];
    49: reg_0061 <= imem04_in[7:4];
    59: reg_0061 <= imem04_in[7:4];
    endcase
  end

  // REG#62の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0062 <= imem04_in[27:24];
    19: reg_0062 <= imem04_in[27:24];
    43: reg_0062 <= imem04_in[27:24];
    45: reg_0062 <= imem04_in[27:24];
    48: reg_0062 <= imem03_in[91:88];
    50: reg_0062 <= imem03_in[91:88];
    52: reg_0062 <= imem04_in[27:24];
    54: reg_0062 <= imem03_in[91:88];
    56: reg_0062 <= imem04_in[27:24];
    58: reg_0062 <= imem03_in[51:48];
    60: reg_0062 <= imem03_in[51:48];
    62: reg_0062 <= imem03_in[91:88];
    64: reg_0062 <= imem07_in[7:4];
    66: reg_0062 <= imem07_in[7:4];
    68: reg_0062 <= imem03_in[91:88];
    70: reg_0062 <= imem07_in[7:4];
    72: reg_0062 <= imem03_in[59:56];
    74: reg_0062 <= imem03_in[91:88];
    76: reg_0062 <= imem03_in[59:56];
    78: reg_0062 <= imem04_in[27:24];
    80: reg_0062 <= imem03_in[59:56];
    82: reg_0062 <= imem03_in[59:56];
    84: reg_0062 <= imem03_in[59:56];
    86: reg_0062 <= imem04_in[27:24];
    88: reg_0062 <= imem03_in[91:88];
    endcase
  end

  // REG#63の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0063 <= imem04_in[79:76];
    19: reg_0063 <= imem04_in[79:76];
    39: reg_0063 <= imem02_in[31:28];
    41: reg_0063 <= imem04_in[79:76];
    44: reg_0063 <= imem02_in[31:28];
    46: reg_0063 <= imem05_in[15:12];
    48: reg_0063 <= imem04_in[79:76];
    50: reg_0063 <= imem05_in[15:12];
    67: reg_0063 <= imem04_in[79:76];
    69: reg_0063 <= imem02_in[31:28];
    71: reg_0063 <= imem02_in[31:28];
    74: reg_0063 <= imem04_in[79:76];
    76: reg_0063 <= imem05_in[15:12];
    78: reg_0063 <= imem02_in[31:28];
    80: reg_0063 <= imem05_in[15:12];
    82: reg_0063 <= imem04_in[79:76];
    85: reg_0063 <= imem04_in[79:76];
    87: reg_0063 <= imem05_in[15:12];
    endcase
  end

  // REG#64の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0064 <= imem04_in[103:100];
    19: reg_0064 <= imem04_in[103:100];
    36: reg_0064 <= imem01_in[39:36];
    38: reg_0064 <= imem04_in[103:100];
    40: reg_0064 <= imem04_in[31:28];
    42: reg_0064 <= imem04_in[103:100];
    96: reg_0064 <= imem01_in[39:36];
    endcase
  end

  // REG#65の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0065 <= imem04_in[35:32];
    19: reg_0065 <= imem04_in[35:32];
    43: reg_0065 <= imem04_in[35:32];
    45: reg_0065 <= imem04_in[35:32];
    48: reg_0065 <= imem04_in[35:32];
    51: reg_0065 <= imem00_in[43:40];
    53: reg_0065 <= imem04_in[35:32];
    55: reg_0065 <= imem04_in[35:32];
    57: reg_0065 <= imem07_in[111:108];
    59: reg_0065 <= imem04_in[35:32];
    endcase
  end

  // REG#66の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0066 <= imem04_in[43:40];
    19: reg_0066 <= imem04_in[43:40];
    42: reg_0066 <= imem04_in[43:40];
    endcase
  end

  // REG#67の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0067 <= imem04_in[51:48];
    19: reg_0067 <= imem04_in[51:48];
    36: reg_0067 <= imem04_in[51:48];
    38: reg_0067 <= imem02_in[111:108];
    40: reg_0067 <= imem02_in[111:108];
    42: reg_0067 <= imem04_in[51:48];
    endcase
  end

  // REG#68の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0068 <= imem04_in[67:64];
    19: reg_0068 <= imem04_in[67:64];
    36: reg_0068 <= imem01_in[95:92];
    38: reg_0068 <= imem05_in[27:24];
    40: reg_0068 <= imem01_in[95:92];
    42: reg_0068 <= imem04_in[67:64];
    93: reg_0068 <= imem04_in[67:64];
    95: reg_0068 <= imem01_in[95:92];
    97: reg_0068 <= imem04_in[67:64];
    endcase
  end

  // REG#69の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0069 <= imem04_in[83:80];
    19: reg_0069 <= imem04_in[83:80];
    41: reg_0069 <= imem05_in[123:120];
    43: reg_0069 <= imem05_in[123:120];
    45: reg_0069 <= imem00_in[91:88];
    47: reg_0069 <= imem05_in[123:120];
    49: reg_0069 <= imem05_in[123:120];
    51: reg_0069 <= imem00_in[91:88];
    53: reg_0069 <= imem02_in[43:40];
    55: reg_0069 <= imem00_in[91:88];
    84: reg_0069 <= imem02_in[43:40];
    endcase
  end

  // REG#70の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0070 <= imem04_in[95:92];
    19: reg_0070 <= imem04_in[95:92];
    43: reg_0070 <= imem04_in[95:92];
    45: reg_0070 <= imem04_in[95:92];
    47: reg_0070 <= imem01_in[111:108];
    49: reg_0070 <= imem04_in[95:92];
    55: reg_0070 <= imem04_in[95:92];
    57: reg_0070 <= imem01_in[111:108];
    59: reg_0070 <= imem04_in[95:92];
    96: reg_0070 <= imem01_in[111:108];
    endcase
  end

  // REG#71の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0071 <= imem04_in[75:72];
    19: reg_0071 <= imem04_in[75:72];
    41: reg_0071 <= imem06_in[3:0];
    43: reg_0071 <= imem06_in[3:0];
    45: reg_0071 <= imem04_in[75:72];
    48: reg_0071 <= imem06_in[59:56];
    50: reg_0071 <= imem06_in[59:56];
    52: reg_0071 <= imem04_in[75:72];
    54: reg_0071 <= imem04_in[75:72];
    56: reg_0071 <= imem06_in[3:0];
    59: reg_0071 <= imem04_in[75:72];
    97: reg_0071 <= imem06_in[3:0];
    endcase
  end

  // REG#72の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0072 <= imem04_in[107:104];
    19: reg_0072 <= imem04_in[107:104];
    40: reg_0072 <= imem04_in[107:104];
    42: reg_0072 <= imem04_in[107:104];
    endcase
  end

  // REG#73の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0073 <= imem02_in[111:108];
    19: reg_0073 <= imem06_in[15:12];
    21: reg_0073 <= imem06_in[15:12];
    23: reg_0073 <= imem06_in[15:12];
    25: reg_0073 <= imem02_in[111:108];
    28: reg_0073 <= imem05_in[123:120];
    30: reg_0073 <= imem02_in[111:108];
    32: reg_0073 <= imem02_in[111:108];
    34: reg_0073 <= imem05_in[123:120];
    36: reg_0073 <= imem06_in[15:12];
    39: reg_0073 <= imem06_in[15:12];
    58: reg_0073 <= imem02_in[111:108];
    60: reg_0073 <= imem02_in[111:108];
    62: reg_0073 <= imem06_in[15:12];
    64: reg_0073 <= imem02_in[111:108];
    66: reg_0073 <= imem06_in[15:12];
    68: reg_0073 <= imem06_in[15:12];
    70: reg_0073 <= imem04_in[55:52];
    72: reg_0073 <= imem06_in[15:12];
    74: reg_0073 <= imem02_in[111:108];
    76: reg_0073 <= imem06_in[15:12];
    78: reg_0073 <= imem02_in[111:108];
    80: reg_0073 <= imem02_in[111:108];
    82: reg_0073 <= imem00_in[3:0];
    84: reg_0073 <= imem02_in[111:108];
    endcase
  end

  // REG#74の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0074 <= imem04_in[99:96];
    19: reg_0074 <= imem04_in[99:96];
    42: reg_0074 <= imem04_in[99:96];
    endcase
  end

  // REG#75の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0075 <= imem04_in[91:88];
    19: reg_0075 <= imem04_in[91:88];
    43: reg_0075 <= imem02_in[31:28];
    45: reg_0075 <= imem04_in[91:88];
    47: reg_0075 <= imem04_in[91:88];
    49: reg_0075 <= imem04_in[91:88];
    60: reg_0075 <= imem07_in[3:0];
    62: reg_0075 <= imem07_in[3:0];
    64: reg_0075 <= imem00_in[71:68];
    66: reg_0075 <= imem00_in[71:68];
    68: reg_0075 <= imem04_in[91:88];
    70: reg_0075 <= imem05_in[127:124];
    72: reg_0075 <= imem00_in[71:68];
    74: reg_0075 <= imem03_in[123:120];
    76: reg_0075 <= imem04_in[91:88];
    78: reg_0075 <= imem07_in[3:0];
    80: reg_0075 <= imem00_in[71:68];
    82: reg_0075 <= imem00_in[71:68];
    84: reg_0075 <= imem02_in[31:28];
    endcase
  end

  // REG#76の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0076 <= imem04_in[47:44];
    19: reg_0076 <= imem04_in[47:44];
    42: reg_0076 <= imem04_in[47:44];
    96: reg_0076 <= imem04_in[47:44];
    endcase
  end

  // REG#77の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0077 <= imem02_in[99:96];
    19: reg_0077 <= imem02_in[99:96];
    21: reg_0077 <= imem02_in[99:96];
    84: reg_0077 <= imem02_in[99:96];
    96: reg_0077 <= imem03_in[127:124];
    endcase
  end

  // REG#78の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0078 <= imem04_in[23:20];
    19: reg_0078 <= imem04_in[23:20];
    43: reg_0078 <= imem04_in[59:56];
    45: reg_0078 <= imem04_in[59:56];
    47: reg_0078 <= imem04_in[59:56];
    49: reg_0078 <= imem04_in[23:20];
    60: reg_0078 <= imem00_in[83:80];
    62: reg_0078 <= imem04_in[23:20];
    64: reg_0078 <= imem04_in[23:20];
    66: reg_0078 <= imem00_in[83:80];
    68: reg_0078 <= imem04_in[59:56];
    70: reg_0078 <= imem06_in[47:44];
    72: reg_0078 <= imem04_in[23:20];
    74: reg_0078 <= imem06_in[11:8];
    76: reg_0078 <= imem06_in[11:8];
    78: reg_0078 <= imem00_in[83:80];
    80: reg_0078 <= imem04_in[59:56];
    82: reg_0078 <= imem04_in[59:56];
    85: reg_0078 <= imem00_in[83:80];
    87: reg_0078 <= imem00_in[83:80];
    89: reg_0078 <= imem00_in[83:80];
    91: reg_0078 <= imem00_in[83:80];
    97: reg_0078 <= imem04_in[23:20];
    endcase
  end

  // REG#79の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0079 <= imem02_in[115:112];
    19: reg_0079 <= imem02_in[115:112];
    21: reg_0079 <= imem02_in[115:112];
    83: reg_0079 <= imem02_in[115:112];
    86: reg_0079 <= imem04_in[15:12];
    88: reg_0079 <= imem04_in[15:12];
    90: reg_0079 <= imem05_in[111:108];
    92: reg_0079 <= imem02_in[115:112];
    94: reg_0079 <= imem02_in[115:112];
    96: reg_0079 <= imem02_in[115:112];
    endcase
  end

  // REG#80の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0080 <= imem02_in[31:28];
    20: reg_0080 <= imem06_in[11:8];
    22: reg_0080 <= imem02_in[31:28];
    24: reg_0080 <= imem02_in[31:28];
    26: reg_0080 <= imem02_in[31:28];
    53: reg_0080 <= imem02_in[31:28];
    55: reg_0080 <= imem02_in[31:28];
    57: reg_0080 <= imem06_in[11:8];
    endcase
  end

  // REG#81の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0081 <= imem02_in[27:24];
    20: reg_0081 <= imem00_in[99:96];
    22: reg_0081 <= imem04_in[39:36];
    24: reg_0081 <= imem00_in[99:96];
    26: reg_0081 <= imem02_in[27:24];
    52: reg_0081 <= imem02_in[27:24];
    93: reg_0081 <= imem06_in[91:88];
    95: reg_0081 <= imem06_in[91:88];
    97: reg_0081 <= imem00_in[99:96];
    endcase
  end

  // REG#82の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0082 <= imem02_in[67:64];
    20: reg_0082 <= imem02_in[75:72];
    22: reg_0082 <= imem02_in[67:64];
    24: reg_0082 <= imem02_in[75:72];
    26: reg_0082 <= imem02_in[75:72];
    45: reg_0082 <= imem02_in[75:72];
    58: reg_0082 <= imem04_in[31:28];
    60: reg_0082 <= imem02_in[75:72];
    62: reg_0082 <= imem02_in[75:72];
    64: reg_0082 <= imem02_in[67:64];
    66: reg_0082 <= imem07_in[123:120];
    68: reg_0082 <= imem06_in[111:108];
    70: reg_0082 <= imem04_in[31:28];
    72: reg_0082 <= imem02_in[75:72];
    85: reg_0082 <= imem02_in[75:72];
    endcase
  end

  // REG#83の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0083 <= imem02_in[3:0];
    21: reg_0083 <= imem02_in[3:0];
    81: reg_0083 <= imem07_in[31:28];
    83: reg_0083 <= imem07_in[31:28];
    85: reg_0083 <= imem02_in[3:0];
    endcase
  end

  // REG#84の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0084 <= imem02_in[79:76];
    21: reg_0084 <= imem02_in[79:76];
    83: reg_0084 <= imem02_in[79:76];
    87: reg_0084 <= imem06_in[107:104];
    89: reg_0084 <= imem06_in[107:104];
    endcase
  end

  // REG#85の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0085 <= imem02_in[39:36];
    21: reg_0085 <= imem02_in[39:36];
    81: reg_0085 <= imem00_in[27:24];
    83: reg_0085 <= imem00_in[27:24];
    85: reg_0085 <= imem02_in[39:36];
    endcase
  end

  // REG#86の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0086 <= imem02_in[55:52];
    21: reg_0086 <= imem02_in[55:52];
    85: reg_0086 <= imem02_in[55:52];
    endcase
  end

  // REG#87の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0087 <= imem02_in[95:92];
    21: reg_0087 <= imem01_in[107:104];
    23: reg_0087 <= imem01_in[107:104];
    25: reg_0087 <= imem01_in[107:104];
    46: reg_0087 <= imem05_in[19:16];
    48: reg_0087 <= imem02_in[95:92];
    50: reg_0087 <= imem02_in[95:92];
    52: reg_0087 <= imem02_in[95:92];
    97: reg_0087 <= imem01_in[107:104];
    endcase
  end

  // REG#88の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0088 <= imem02_in[19:16];
    21: reg_0088 <= imem02_in[19:16];
    86: reg_0088 <= imem00_in[19:16];
    88: reg_0088 <= imem02_in[19:16];
    90: reg_0088 <= imem02_in[19:16];
    92: reg_0088 <= imem00_in[103:100];
    94: reg_0088 <= imem00_in[19:16];
    96: reg_0088 <= imem00_in[103:100];
    endcase
  end

  // REG#89の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0089 <= imem02_in[23:20];
    21: reg_0089 <= imem02_in[23:20];
    83: reg_0089 <= imem02_in[23:20];
    87: reg_0089 <= imem01_in[35:32];
    89: reg_0089 <= imem01_in[35:32];
    91: reg_0089 <= imem01_in[35:32];
    93: reg_0089 <= imem02_in[23:20];
    95: reg_0089 <= imem01_in[35:32];
    endcase
  end

  // REG#90の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0090 <= imem02_in[59:56];
    21: reg_0090 <= imem02_in[59:56];
    84: reg_0090 <= imem02_in[59:56];
    endcase
  end

  // REG#91の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0091 <= imem02_in[71:68];
    21: reg_0091 <= imem02_in[71:68];
    84: reg_0091 <= imem02_in[71:68];
    endcase
  end

  // REG#92の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0092 <= imem02_in[7:4];
    22: reg_0092 <= imem02_in[7:4];
    24: reg_0092 <= imem07_in[35:32];
    26: reg_0092 <= imem07_in[35:32];
    28: reg_0092 <= imem02_in[91:88];
    30: reg_0092 <= imem02_in[7:4];
    32: reg_0092 <= imem02_in[7:4];
    34: reg_0092 <= imem02_in[7:4];
    36: reg_0092 <= imem02_in[7:4];
    38: reg_0092 <= imem07_in[35:32];
    40: reg_0092 <= imem04_in[91:88];
    42: reg_0092 <= imem02_in[91:88];
    44: reg_0092 <= imem02_in[7:4];
    46: reg_0092 <= imem04_in[91:88];
    48: reg_0092 <= imem02_in[7:4];
    50: reg_0092 <= imem07_in[35:32];
    52: reg_0092 <= imem04_in[91:88];
    54: reg_0092 <= imem04_in[91:88];
    56: reg_0092 <= imem02_in[7:4];
    58: reg_0092 <= imem07_in[35:32];
    60: reg_0092 <= imem02_in[7:4];
    62: reg_0092 <= imem02_in[7:4];
    64: reg_0092 <= imem01_in[67:64];
    66: reg_0092 <= imem02_in[7:4];
    68: reg_0092 <= imem02_in[91:88];
    70: reg_0092 <= imem07_in[35:32];
    72: reg_0092 <= imem07_in[35:32];
    74: reg_0092 <= imem07_in[35:32];
    77: reg_0092 <= imem01_in[67:64];
    79: reg_0092 <= imem01_in[67:64];
    81: reg_0092 <= imem03_in[87:84];
    83: reg_0092 <= imem02_in[7:4];
    85: reg_0092 <= imem04_in[91:88];
    87: reg_0092 <= imem07_in[35:32];
    89: reg_0092 <= imem03_in[87:84];
    92: reg_0092 <= imem03_in[87:84];
    94: reg_0092 <= imem01_in[67:64];
    96: reg_0092 <= imem01_in[67:64];
    endcase
  end

  // REG#93の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0093 <= imem02_in[107:104];
    22: reg_0093 <= imem02_in[107:104];
    24: reg_0093 <= imem07_in[47:44];
    26: reg_0093 <= imem02_in[107:104];
    50: reg_0093 <= imem06_in[107:104];
    52: reg_0093 <= imem07_in[47:44];
    54: reg_0093 <= imem06_in[67:64];
    56: reg_0093 <= imem06_in[67:64];
    60: reg_0093 <= imem06_in[107:104];
    62: reg_0093 <= imem06_in[107:104];
    64: reg_0093 <= imem07_in[47:44];
    66: reg_0093 <= imem06_in[67:64];
    68: reg_0093 <= imem02_in[107:104];
    70: reg_0093 <= imem06_in[67:64];
    73: reg_0093 <= imem02_in[107:104];
    75: reg_0093 <= imem06_in[67:64];
    77: reg_0093 <= imem06_in[67:64];
    79: reg_0093 <= imem02_in[107:104];
    81: reg_0093 <= imem07_in[47:44];
    83: reg_0093 <= imem06_in[67:64];
    85: reg_0093 <= imem06_in[67:64];
    88: reg_0093 <= imem06_in[107:104];
    91: reg_0093 <= imem05_in[7:4];
    93: reg_0093 <= imem02_in[107:104];
    95: reg_0093 <= imem06_in[107:104];
    endcase
  end

  // REG#94の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0094 <= imem02_in[103:100];
    22: reg_0094 <= imem05_in[83:80];
    24: reg_0094 <= imem07_in[91:88];
    26: reg_0094 <= imem05_in[83:80];
    28: reg_0094 <= imem02_in[103:100];
    30: reg_0094 <= imem02_in[103:100];
    32: reg_0094 <= imem07_in[43:40];
    34: reg_0094 <= imem02_in[103:100];
    36: reg_0094 <= imem02_in[103:100];
    38: reg_0094 <= imem02_in[103:100];
    40: reg_0094 <= imem05_in[83:80];
    42: reg_0094 <= imem07_in[43:40];
    44: reg_0094 <= imem05_in[83:80];
    46: reg_0094 <= imem07_in[43:40];
    48: reg_0094 <= imem02_in[103:100];
    50: reg_0094 <= imem05_in[83:80];
    67: reg_0094 <= imem02_in[103:100];
    69: reg_0094 <= imem02_in[103:100];
    71: reg_0094 <= imem02_in[103:100];
    74: reg_0094 <= imem07_in[43:40];
    76: reg_0094 <= imem02_in[103:100];
    78: reg_0094 <= imem05_in[83:80];
    81: reg_0094 <= imem02_in[103:100];
    83: reg_0094 <= imem02_in[103:100];
    85: reg_0094 <= imem07_in[91:88];
    87: reg_0094 <= imem02_in[103:100];
    89: reg_0094 <= imem02_in[127:124];
    91: reg_0094 <= imem06_in[31:28];
    93: reg_0094 <= imem05_in[83:80];
    95: reg_0094 <= imem02_in[103:100];
    97: reg_0094 <= imem06_in[31:28];
    endcase
  end

  // REG#95の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0095 <= imem02_in[35:32];
    22: reg_0095 <= imem06_in[119:116];
    24: reg_0095 <= imem06_in[119:116];
    26: reg_0095 <= imem02_in[35:32];
    47: reg_0095 <= imem02_in[51:48];
    49: reg_0095 <= imem02_in[51:48];
    51: reg_0095 <= imem02_in[35:32];
    54: reg_0095 <= imem02_in[35:32];
    56: reg_0095 <= imem06_in[119:116];
    58: reg_0095 <= imem02_in[51:48];
    60: reg_0095 <= imem02_in[35:32];
    62: reg_0095 <= imem02_in[51:48];
    64: reg_0095 <= imem02_in[123:120];
    66: reg_0095 <= imem07_in[3:0];
    68: reg_0095 <= imem02_in[51:48];
    70: reg_0095 <= imem02_in[51:48];
    72: reg_0095 <= imem02_in[123:120];
    80: reg_0095 <= imem07_in[3:0];
    84: reg_0095 <= imem02_in[123:120];
    endcase
  end

  // REG#96の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0096 <= imem02_in[43:40];
    22: reg_0096 <= imem00_in[91:88];
    24: reg_0096 <= imem02_in[43:40];
    26: reg_0096 <= imem02_in[43:40];
    52: reg_0096 <= imem00_in[91:88];
    54: reg_0096 <= imem07_in[19:16];
    56: reg_0096 <= imem00_in[91:88];
    58: reg_0096 <= imem07_in[19:16];
    60: reg_0096 <= imem01_in[111:108];
    62: reg_0096 <= imem07_in[19:16];
    64: reg_0096 <= imem04_in[15:12];
    66: reg_0096 <= imem02_in[43:40];
    68: reg_0096 <= imem00_in[91:88];
    70: reg_0096 <= imem07_in[19:16];
    72: reg_0096 <= imem02_in[43:40];
    83: reg_0096 <= imem00_in[91:88];
    85: reg_0096 <= imem07_in[19:16];
    87: reg_0096 <= imem00_in[91:88];
    89: reg_0096 <= imem00_in[91:88];
    91: reg_0096 <= imem07_in[19:16];
    93: reg_0096 <= imem04_in[15:12];
    95: reg_0096 <= imem01_in[111:108];
    endcase
  end

  // REG#97の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0097 <= imem02_in[47:44];
    22: reg_0097 <= imem00_in[111:108];
    24: reg_0097 <= imem00_in[111:108];
    26: reg_0097 <= imem02_in[47:44];
    53: reg_0097 <= imem00_in[111:108];
    55: reg_0097 <= imem02_in[47:44];
    57: reg_0097 <= imem02_in[47:44];
    59: reg_0097 <= imem01_in[39:36];
    61: reg_0097 <= imem01_in[39:36];
    63: reg_0097 <= imem01_in[39:36];
    65: reg_0097 <= imem00_in[111:108];
    67: reg_0097 <= imem07_in[115:112];
    69: reg_0097 <= imem00_in[111:108];
    71: reg_0097 <= imem00_in[111:108];
    73: reg_0097 <= imem00_in[111:108];
    75: reg_0097 <= imem07_in[115:112];
    77: reg_0097 <= imem01_in[39:36];
    79: reg_0097 <= imem01_in[39:36];
    81: reg_0097 <= imem07_in[115:112];
    83: reg_0097 <= imem02_in[47:44];
    85: reg_0097 <= imem00_in[111:108];
    87: reg_0097 <= imem01_in[39:36];
    89: reg_0097 <= imem01_in[39:36];
    91: reg_0097 <= imem01_in[39:36];
    93: reg_0097 <= imem01_in[39:36];
    96: reg_0097 <= imem07_in[115:112];
    endcase
  end

  // REG#98の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0098 <= imem02_in[83:80];
    22: reg_0098 <= imem02_in[83:80];
    24: reg_0098 <= imem00_in[119:116];
    26: reg_0098 <= imem02_in[83:80];
    47: reg_0098 <= imem00_in[119:116];
    49: reg_0098 <= imem07_in[51:48];
    51: reg_0098 <= imem02_in[83:80];
    53: reg_0098 <= imem02_in[83:80];
    55: reg_0098 <= imem07_in[51:48];
    57: reg_0098 <= imem00_in[119:116];
    59: reg_0098 <= imem00_in[119:116];
    61: reg_0098 <= imem07_in[51:48];
    63: reg_0098 <= imem02_in[83:80];
    72: reg_0098 <= imem02_in[83:80];
    84: reg_0098 <= imem00_in[119:116];
    86: reg_0098 <= imem07_in[51:48];
    88: reg_0098 <= imem07_in[3:0];
    90: reg_0098 <= imem07_in[3:0];
    92: reg_0098 <= imem07_in[3:0];
    94: reg_0098 <= imem07_in[3:0];
    96: reg_0098 <= imem07_in[51:48];
    endcase
  end

  // REG#99の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0099 <= imem01_in[43:40];
    48: reg_0099 <= imem03_in[31:28];
    50: reg_0099 <= imem01_in[43:40];
    52: reg_0099 <= imem01_in[43:40];
    55: reg_0099 <= imem03_in[31:28];
    88: reg_0099 <= imem01_in[43:40];
    90: reg_0099 <= imem01_in[43:40];
    92: reg_0099 <= imem07_in[43:40];
    94: reg_0099 <= imem07_in[43:40];
    96: reg_0099 <= imem03_in[31:28];
    endcase
  end

  // REG#100の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0100 <= imem01_in[71:68];
    50: reg_0100 <= imem07_in[83:80];
    52: reg_0100 <= imem01_in[71:68];
    54: reg_0100 <= imem07_in[59:56];
    56: reg_0100 <= imem07_in[59:56];
    58: reg_0100 <= imem07_in[59:56];
    60: reg_0100 <= imem07_in[59:56];
    62: reg_0100 <= imem01_in[71:68];
    64: reg_0100 <= imem01_in[71:68];
    66: reg_0100 <= imem07_in[59:56];
    68: reg_0100 <= imem01_in[71:68];
    71: reg_0100 <= imem07_in[59:56];
    73: reg_0100 <= imem07_in[83:80];
    75: reg_0100 <= imem01_in[71:68];
    77: reg_0100 <= imem07_in[59:56];
    79: reg_0100 <= imem07_in[59:56];
    88: reg_0100 <= imem07_in[19:16];
    90: reg_0100 <= imem07_in[59:56];
    92: reg_0100 <= imem07_in[19:16];
    94: reg_0100 <= imem07_in[59:56];
    96: reg_0100 <= imem01_in[71:68];
    endcase
  end

  // REG#101の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0101 <= imem01_in[79:76];
    51: reg_0101 <= imem01_in[79:76];
    53: reg_0101 <= imem01_in[79:76];
    endcase
  end

  // REG#102の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0102 <= imem01_in[63:60];
    51: reg_0102 <= imem00_in[99:96];
    53: reg_0102 <= imem00_in[99:96];
    55: reg_0102 <= imem00_in[99:96];
    89: reg_0102 <= imem07_in[27:24];
    91: reg_0102 <= imem07_in[27:24];
    93: reg_0102 <= imem07_in[27:24];
    95: reg_0102 <= imem07_in[27:24];
    endcase
  end

  // REG#103の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0103 <= imem01_in[19:16];
    51: reg_0103 <= imem01_in[95:92];
    53: reg_0103 <= imem01_in[95:92];
    endcase
  end

  // REG#104の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0104 <= imem01_in[39:36];
    52: reg_0104 <= imem01_in[39:36];
    54: reg_0104 <= imem00_in[123:120];
    56: reg_0104 <= imem01_in[39:36];
    58: reg_0104 <= imem01_in[39:36];
    60: reg_0104 <= imem00_in[123:120];
    62: reg_0104 <= imem01_in[39:36];
    64: reg_0104 <= imem00_in[123:120];
    66: reg_0104 <= imem01_in[39:36];
    68: reg_0104 <= imem01_in[39:36];
    70: reg_0104 <= imem00_in[123:120];
    72: reg_0104 <= imem04_in[67:64];
    74: reg_0104 <= imem00_in[123:120];
    76: reg_0104 <= imem04_in[67:64];
    78: reg_0104 <= imem01_in[39:36];
    80: reg_0104 <= imem04_in[67:64];
    82: reg_0104 <= imem00_in[123:120];
    84: reg_0104 <= imem04_in[67:64];
    86: reg_0104 <= imem00_in[27:24];
    88: reg_0104 <= imem01_in[39:36];
    90: reg_0104 <= imem00_in[123:120];
    93: reg_0104 <= imem00_in[27:24];
    95: reg_0104 <= imem01_in[39:36];
    endcase
  end

  // REG#105の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0105 <= imem01_in[7:4];
    52: reg_0105 <= imem01_in[7:4];
    55: reg_0105 <= imem07_in[71:68];
    57: reg_0105 <= imem03_in[3:0];
    59: reg_0105 <= imem03_in[3:0];
    61: reg_0105 <= imem07_in[71:68];
    63: reg_0105 <= imem07_in[71:68];
    65: reg_0105 <= imem07_in[71:68];
    67: reg_0105 <= imem03_in[99:96];
    69: reg_0105 <= imem01_in[7:4];
    95: reg_0105 <= imem03_in[99:96];
    endcase
  end

  // REG#106の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0106 <= imem01_in[75:72];
    52: reg_0106 <= imem01_in[75:72];
    55: reg_0106 <= imem01_in[19:16];
    57: reg_0106 <= imem01_in[75:72];
    59: reg_0106 <= imem01_in[75:72];
    61: reg_0106 <= imem01_in[75:72];
    63: reg_0106 <= imem01_in[19:16];
    65: reg_0106 <= imem01_in[19:16];
    67: reg_0106 <= imem06_in[3:0];
    69: reg_0106 <= imem01_in[19:16];
    95: reg_0106 <= imem01_in[19:16];
    endcase
  end

  // REG#107の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0107 <= imem01_in[91:88];
    52: reg_0107 <= imem01_in[91:88];
    55: reg_0107 <= imem01_in[95:92];
    57: reg_0107 <= imem03_in[79:76];
    59: reg_0107 <= imem03_in[79:76];
    61: reg_0107 <= imem03_in[79:76];
    63: reg_0107 <= imem05_in[27:24];
    65: reg_0107 <= imem01_in[95:92];
    67: reg_0107 <= imem01_in[91:88];
    69: reg_0107 <= imem05_in[27:24];
    71: reg_0107 <= imem03_in[79:76];
    73: reg_0107 <= imem03_in[79:76];
    75: reg_0107 <= imem05_in[27:24];
    77: reg_0107 <= imem01_in[91:88];
    79: reg_0107 <= imem05_in[27:24];
    87: reg_0107 <= imem01_in[91:88];
    89: reg_0107 <= imem03_in[79:76];
    91: reg_0107 <= imem01_in[91:88];
    93: reg_0107 <= imem03_in[79:76];
    95: reg_0107 <= imem03_in[79:76];
    endcase
  end

  // REG#108の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0108 <= imem01_in[59:56];
    52: reg_0108 <= imem01_in[59:56];
    55: reg_0108 <= imem01_in[59:56];
    57: reg_0108 <= imem04_in[71:68];
    59: reg_0108 <= imem04_in[71:68];
    97: reg_0108 <= imem04_in[71:68];
    endcase
  end

  // REG#109の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0109 <= imem01_in[87:84];
    53: reg_0109 <= imem01_in[87:84];
    endcase
  end

  // REG#110の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0110 <= imem01_in[115:112];
    53: reg_0110 <= imem01_in[115:112];
    endcase
  end

  // REG#111の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0111 <= imem01_in[23:20];
    53: reg_0111 <= imem01_in[23:20];
    endcase
  end

  // REG#112の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0112 <= imem01_in[55:52];
    53: reg_0112 <= imem01_in[55:52];
    endcase
  end

  // REG#113の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0113 <= imem01_in[103:100];
    53: reg_0113 <= imem01_in[103:100];
    endcase
  end

  // REG#114の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0114 <= imem01_in[67:64];
    53: reg_0114 <= imem01_in[67:64];
    endcase
  end

  // REG#115の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0115 <= imem01_in[83:80];
    53: reg_0115 <= imem01_in[83:80];
    endcase
  end

  // REG#116の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0116 <= imem01_in[35:32];
    53: reg_0116 <= imem01_in[35:32];
    endcase
  end

  // REG#117の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0117 <= imem01_in[99:96];
    53: reg_0117 <= imem01_in[99:96];
    endcase
  end

  // REG#118の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0118 <= imem01_in[27:24];
    54: reg_0118 <= imem02_in[75:72];
    56: reg_0118 <= imem02_in[75:72];
    58: reg_0118 <= imem00_in[31:28];
    60: reg_0118 <= imem01_in[27:24];
    62: reg_0118 <= imem06_in[11:8];
    64: reg_0118 <= imem01_in[27:24];
    66: reg_0118 <= imem01_in[95:92];
    68: reg_0118 <= imem06_in[11:8];
    70: reg_0118 <= imem06_in[11:8];
    73: reg_0118 <= imem02_in[75:72];
    75: reg_0118 <= imem00_in[35:32];
    77: reg_0118 <= imem00_in[35:32];
    79: reg_0118 <= imem00_in[35:32];
    81: reg_0118 <= imem00_in[35:32];
    83: reg_0118 <= imem00_in[35:32];
    85: reg_0118 <= imem01_in[27:24];
    87: reg_0118 <= imem00_in[35:32];
    89: reg_0118 <= imem00_in[35:32];
    91: reg_0118 <= imem00_in[31:28];
    endcase
  end

  // REG#119の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0119 <= imem01_in[47:44];
    54: reg_0119 <= imem01_in[47:44];
    56: reg_0119 <= imem01_in[47:44];
    58: reg_0119 <= imem03_in[3:0];
    60: reg_0119 <= imem06_in[119:116];
    62: reg_0119 <= imem01_in[47:44];
    64: reg_0119 <= imem03_in[3:0];
    66: reg_0119 <= imem01_in[47:44];
    68: reg_0119 <= imem01_in[47:44];
    70: reg_0119 <= imem06_in[119:116];
    73: reg_0119 <= imem06_in[119:116];
    75: reg_0119 <= imem03_in[3:0];
    77: reg_0119 <= imem07_in[123:120];
    79: reg_0119 <= imem06_in[119:116];
    81: reg_0119 <= imem05_in[11:8];
    83: reg_0119 <= imem05_in[11:8];
    85: reg_0119 <= imem06_in[119:116];
    87: reg_0119 <= imem07_in[123:120];
    89: reg_0119 <= imem01_in[47:44];
    91: reg_0119 <= imem06_in[119:116];
    93: reg_0119 <= imem03_in[3:0];
    95: reg_0119 <= imem01_in[47:44];
    endcase
  end

  // REG#120の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0120 <= imem01_in[51:48];
    54: reg_0120 <= imem03_in[79:76];
    56: reg_0120 <= imem02_in[19:16];
    58: reg_0120 <= imem04_in[19:16];
    60: reg_0120 <= imem01_in[51:48];
    62: reg_0120 <= imem02_in[19:16];
    65: reg_0120 <= imem06_in[35:32];
    67: reg_0120 <= imem01_in[51:48];
    69: reg_0120 <= imem01_in[51:48];
    92: reg_0120 <= imem01_in[51:48];
    95: reg_0120 <= imem01_in[51:48];
    endcase
  end

  // REG#121の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0121 <= imem01_in[107:104];
    54: reg_0121 <= imem01_in[99:96];
    56: reg_0121 <= imem01_in[99:96];
    58: reg_0121 <= imem01_in[99:96];
    60: reg_0121 <= imem01_in[99:96];
    62: reg_0121 <= imem06_in[91:88];
    64: reg_0121 <= imem06_in[91:88];
    66: reg_0121 <= imem01_in[107:104];
    68: reg_0121 <= imem06_in[91:88];
    70: reg_0121 <= imem01_in[107:104];
    72: reg_0121 <= imem01_in[99:96];
    74: reg_0121 <= imem01_in[107:104];
    76: reg_0121 <= imem01_in[99:96];
    78: reg_0121 <= imem01_in[99:96];
    80: reg_0121 <= imem01_in[99:96];
    82: reg_0121 <= imem01_in[99:96];
    84: reg_0121 <= imem01_in[99:96];
    86: reg_0121 <= imem06_in[91:88];
    97: reg_0121 <= imem06_in[91:88];
    endcase
  end

  // REG#122の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0122 <= imem01_in[11:8];
    54: reg_0122 <= imem01_in[11:8];
    56: reg_0122 <= imem04_in[23:20];
    58: reg_0122 <= imem04_in[23:20];
    61: reg_0122 <= imem04_in[23:20];
    63: reg_0122 <= imem04_in[23:20];
    65: reg_0122 <= imem01_in[11:8];
    67: reg_0122 <= imem00_in[99:96];
    69: reg_0122 <= imem01_in[11:8];
    94: reg_0122 <= imem01_in[11:8];
    97: reg_0122 <= imem01_in[11:8];
    endcase
  end

  // REG#123の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0123 <= imem01_in[3:0];
    54: reg_0123 <= imem01_in[3:0];
    56: reg_0123 <= imem04_in[127:124];
    58: reg_0123 <= imem04_in[127:124];
    61: reg_0123 <= imem01_in[107:104];
    63: reg_0123 <= imem01_in[107:104];
    65: reg_0123 <= imem07_in[119:116];
    67: reg_0123 <= imem01_in[107:104];
    69: reg_0123 <= imem07_in[119:116];
    71: reg_0123 <= imem00_in[67:64];
    73: reg_0123 <= imem07_in[119:116];
    75: reg_0123 <= imem07_in[119:116];
    80: reg_0123 <= imem07_in[119:116];
    83: reg_0123 <= imem04_in[127:124];
    endcase
  end

  // REG#124の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0124 <= imem01_in[15:12];
    54: reg_0124 <= imem03_in[7:4];
    56: reg_0124 <= imem01_in[23:20];
    58: reg_0124 <= imem01_in[15:12];
    60: reg_0124 <= imem01_in[23:20];
    62: reg_0124 <= imem01_in[15:12];
    64: reg_0124 <= imem01_in[15:12];
    66: reg_0124 <= imem01_in[23:20];
    68: reg_0124 <= imem01_in[15:12];
    71: reg_0124 <= imem01_in[15:12];
    73: reg_0124 <= imem01_in[23:20];
    75: reg_0124 <= imem01_in[15:12];
    77: reg_0124 <= imem01_in[23:20];
    79: reg_0124 <= imem01_in[23:20];
    81: reg_0124 <= imem01_in[23:20];
    83: reg_0124 <= imem03_in[7:4];
    85: reg_0124 <= imem01_in[23:20];
    87: reg_0124 <= imem06_in[55:52];
    89: reg_0124 <= imem06_in[55:52];
    endcase
  end

  // REG#125の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0125 <= imem01_in[31:28];
    54: reg_0125 <= imem01_in[31:28];
    56: reg_0125 <= imem01_in[31:28];
    58: reg_0125 <= imem05_in[67:64];
    60: reg_0125 <= imem07_in[67:64];
    62: reg_0125 <= imem07_in[67:64];
    64: reg_0125 <= imem07_in[67:64];
    66: reg_0125 <= imem05_in[67:64];
    76: reg_0125 <= imem07_in[67:64];
    78: reg_0125 <= imem07_in[67:64];
    80: reg_0125 <= imem03_in[83:80];
    82: reg_0125 <= imem03_in[83:80];
    84: reg_0125 <= imem06_in[87:84];
    86: reg_0125 <= imem07_in[67:64];
    88: reg_0125 <= imem05_in[67:64];
    90: reg_0125 <= imem07_in[67:64];
    92: reg_0125 <= imem03_in[83:80];
    94: reg_0125 <= imem03_in[83:80];
    96: reg_0125 <= imem05_in[67:64];
    endcase
  end

  // REG#126の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0126 <= imem01_in[111:108];
    54: reg_0126 <= imem04_in[15:12];
    56: reg_0126 <= imem01_in[111:108];
    58: reg_0126 <= imem04_in[15:12];
    61: reg_0126 <= imem01_in[111:108];
    63: reg_0126 <= imem04_in[15:12];
    65: reg_0126 <= imem04_in[15:12];
    67: reg_0126 <= imem01_in[111:108];
    69: reg_0126 <= imem04_in[15:12];
    71: reg_0126 <= imem01_in[111:108];
    73: reg_0126 <= imem04_in[15:12];
    75: reg_0126 <= imem04_in[15:12];
    77: reg_0126 <= imem00_in[59:56];
    79: reg_0126 <= imem00_in[59:56];
    81: reg_0126 <= imem04_in[15:12];
    83: reg_0126 <= imem04_in[15:12];
    96: reg_0126 <= imem04_in[15:12];
    endcase
  end

  // REG#127の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0127 <= imem01_in[95:92];
    54: reg_0127 <= imem07_in[79:76];
    56: reg_0127 <= imem01_in[95:92];
    58: reg_0127 <= imem01_in[95:92];
    60: reg_0127 <= imem07_in[87:84];
    62: reg_0127 <= imem07_in[11:8];
    64: reg_0127 <= imem07_in[11:8];
    66: reg_0127 <= imem07_in[87:84];
    68: reg_0127 <= imem07_in[11:8];
    70: reg_0127 <= imem01_in[95:92];
    72: reg_0127 <= imem07_in[11:8];
    74: reg_0127 <= imem07_in[79:76];
    76: reg_0127 <= imem07_in[87:84];
    78: reg_0127 <= imem07_in[11:8];
    80: reg_0127 <= imem07_in[79:76];
    83: reg_0127 <= imem07_in[87:84];
    85: reg_0127 <= imem07_in[79:76];
    87: reg_0127 <= imem07_in[87:84];
    89: reg_0127 <= imem07_in[79:76];
    91: reg_0127 <= imem07_in[87:84];
    93: reg_0127 <= imem07_in[79:76];
    95: reg_0127 <= imem06_in[123:120];
    97: reg_0127 <= imem07_in[87:84];
    endcase
  end

  // REG#128の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0128 <= imem05_in[43:40];
    67: reg_0128 <= imem05_in[43:40];
    70: reg_0128 <= imem06_in[35:32];
    73: reg_0128 <= imem05_in[43:40];
    endcase
  end

  // REG#129の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0129 <= imem05_in[79:76];
    70: reg_0129 <= imem05_in[79:76];
    72: reg_0129 <= imem05_in[79:76];
    76: reg_0129 <= imem05_in[55:52];
    78: reg_0129 <= imem05_in[55:52];
    81: reg_0129 <= imem05_in[55:52];
    83: reg_0129 <= imem05_in[55:52];
    85: reg_0129 <= imem05_in[79:76];
    87: reg_0129 <= imem05_in[55:52];
    endcase
  end

  // REG#130の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0130 <= imem05_in[91:88];
    70: reg_0130 <= imem05_in[91:88];
    72: reg_0130 <= imem05_in[91:88];
    76: reg_0130 <= imem05_in[59:56];
    78: reg_0130 <= imem05_in[91:88];
    81: reg_0130 <= imem05_in[91:88];
    83: reg_0130 <= imem05_in[59:56];
    85: reg_0130 <= imem05_in[91:88];
    87: reg_0130 <= imem05_in[91:88];
    94: reg_0130 <= imem05_in[59:56];
    96: reg_0130 <= imem05_in[59:56];
    endcase
  end

  // REG#131の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0131 <= imem05_in[107:104];
    70: reg_0131 <= imem05_in[107:104];
    72: reg_0131 <= imem05_in[107:104];
    76: reg_0131 <= imem06_in[99:96];
    78: reg_0131 <= imem00_in[127:124];
    80: reg_0131 <= imem06_in[99:96];
    82: reg_0131 <= imem05_in[107:104];
    84: reg_0131 <= imem05_in[107:104];
    86: reg_0131 <= imem00_in[127:124];
    88: reg_0131 <= imem06_in[99:96];
    90: reg_0131 <= imem06_in[43:40];
    92: reg_0131 <= imem06_in[43:40];
    94: reg_0131 <= imem06_in[43:40];
    97: reg_0131 <= imem05_in[107:104];
    endcase
  end

  // REG#132の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0132 <= imem05_in[3:0];
    71: reg_0132 <= imem00_in[99:96];
    73: reg_0132 <= imem00_in[99:96];
    75: reg_0132 <= imem01_in[31:28];
    77: reg_0132 <= imem00_in[99:96];
    79: reg_0132 <= imem01_in[31:28];
    81: reg_0132 <= imem01_in[31:28];
    83: reg_0132 <= imem05_in[3:0];
    85: reg_0132 <= imem01_in[31:28];
    87: reg_0132 <= imem00_in[99:96];
    89: reg_0132 <= imem05_in[3:0];
    91: reg_0132 <= imem00_in[99:96];
    endcase
  end

  // REG#133の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0133 <= imem05_in[31:28];
    72: reg_0133 <= imem05_in[31:28];
    75: reg_0133 <= imem05_in[31:28];
    77: reg_0133 <= imem02_in[123:120];
    79: reg_0133 <= imem02_in[123:120];
    81: reg_0133 <= imem06_in[15:12];
    83: reg_0133 <= imem02_in[123:120];
    85: reg_0133 <= imem05_in[31:28];
    87: reg_0133 <= imem02_in[123:120];
    89: reg_0133 <= imem06_in[15:12];
    endcase
  end

  // REG#134の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0134 <= imem05_in[111:108];
    72: reg_0134 <= imem05_in[111:108];
    76: reg_0134 <= imem01_in[51:48];
    78: reg_0134 <= imem05_in[111:108];
    80: reg_0134 <= imem05_in[111:108];
    82: reg_0134 <= imem01_in[51:48];
    84: reg_0134 <= imem07_in[71:68];
    86: reg_0134 <= imem05_in[111:108];
    89: reg_0134 <= imem05_in[111:108];
    91: reg_0134 <= imem05_in[111:108];
    93: reg_0134 <= imem01_in[51:48];
    endcase
  end

  // REG#135の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0135 <= imem05_in[23:20];
    72: reg_0135 <= imem05_in[23:20];
    74: reg_0135 <= imem05_in[23:20];
    endcase
  end

  // REG#136の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0136 <= imem05_in[27:24];
    73: reg_0136 <= imem05_in[27:24];
    endcase
  end

  // REG#137の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0137 <= imem05_in[103:100];
    73: reg_0137 <= imem05_in[103:100];
    95: reg_0137 <= imem05_in[103:100];
    endcase
  end

  // REG#138の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0138 <= imem05_in[75:72];
    73: reg_0138 <= imem05_in[75:72];
    endcase
  end

  // REG#139の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0139 <= imem05_in[71:68];
    73: reg_0139 <= imem05_in[71:68];
    endcase
  end

  // REG#140の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0140 <= imem05_in[95:92];
    73: reg_0140 <= imem05_in[95:92];
    endcase
  end

  // REG#141の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0141 <= imem05_in[87:84];
    73: reg_0141 <= imem05_in[87:84];
    97: reg_0141 <= imem05_in[87:84];
    endcase
  end

  // REG#142の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0142 <= imem05_in[51:48];
    73: reg_0142 <= imem05_in[51:48];
    92: reg_0142 <= imem05_in[51:48];
    94: reg_0142 <= imem02_in[99:96];
    endcase
  end

  // REG#143の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0143 <= imem05_in[67:64];
    73: reg_0143 <= imem05_in[67:64];
    97: reg_0143 <= imem05_in[67:64];
    endcase
  end

  // REG#144の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0144 <= imem05_in[115:112];
    74: reg_0144 <= imem05_in[115:112];
    endcase
  end

  // REG#145の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0145 <= imem05_in[19:16];
    74: reg_0145 <= imem05_in[19:16];
    endcase
  end

  // REG#146の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0146 <= imem05_in[55:52];
    74: reg_0146 <= imem05_in[55:52];
    endcase
  end

  // REG#147の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0147 <= imem05_in[7:4];
    75: reg_0147 <= imem04_in[3:0];
    77: reg_0147 <= imem04_in[3:0];
    79: reg_0147 <= imem04_in[3:0];
    81: reg_0147 <= imem04_in[3:0];
    83: reg_0147 <= imem04_in[3:0];
    endcase
  end

  // REG#148の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0148 <= imem05_in[11:8];
    75: reg_0148 <= imem05_in[87:84];
    77: reg_0148 <= imem05_in[87:84];
    79: reg_0148 <= imem05_in[87:84];
    88: reg_0148 <= imem05_in[87:84];
    90: reg_0148 <= imem05_in[87:84];
    92: reg_0148 <= imem03_in[47:44];
    94: reg_0148 <= imem03_in[47:44];
    96: reg_0148 <= imem03_in[47:44];
    endcase
  end

  // REG#149の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0149 <= imem05_in[15:12];
    75: reg_0149 <= imem05_in[15:12];
    77: reg_0149 <= imem03_in[71:68];
    79: reg_0149 <= imem05_in[15:12];
    82: reg_0149 <= imem03_in[71:68];
    84: reg_0149 <= imem03_in[99:96];
    86: reg_0149 <= imem03_in[99:96];
    88: reg_0149 <= imem03_in[99:96];
    95: reg_0149 <= imem05_in[15:12];
    endcase
  end

  // REG#150の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0150 <= imem05_in[35:32];
    75: reg_0150 <= imem05_in[35:32];
    77: reg_0150 <= imem07_in[31:28];
    79: reg_0150 <= imem05_in[35:32];
    88: reg_0150 <= imem07_in[31:28];
    90: reg_0150 <= imem07_in[31:28];
    92: reg_0150 <= imem05_in[35:32];
    94: reg_0150 <= imem05_in[35:32];
    endcase
  end

  // REG#151の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0151 <= imem05_in[39:36];
    75: reg_0151 <= imem06_in[23:20];
    77: reg_0151 <= imem05_in[39:36];
    79: reg_0151 <= imem06_in[23:20];
    81: reg_0151 <= imem06_in[87:84];
    83: reg_0151 <= imem06_in[87:84];
    85: reg_0151 <= imem06_in[23:20];
    88: reg_0151 <= imem00_in[99:96];
    90: reg_0151 <= imem00_in[99:96];
    92: reg_0151 <= imem00_in[99:96];
    94: reg_0151 <= imem06_in[23:20];
    96: reg_0151 <= imem05_in[39:36];
    endcase
  end

  // REG#152の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0152 <= imem05_in[47:44];
    75: reg_0152 <= imem06_in[87:84];
    77: reg_0152 <= imem07_in[67:64];
    79: reg_0152 <= imem06_in[87:84];
    81: reg_0152 <= imem07_in[67:64];
    83: reg_0152 <= imem07_in[67:64];
    85: reg_0152 <= imem06_in[87:84];
    87: reg_0152 <= imem05_in[47:44];
    endcase
  end

  // REG#153の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0153 <= imem05_in[83:80];
    75: reg_0153 <= imem00_in[123:120];
    77: reg_0153 <= imem00_in[3:0];
    79: reg_0153 <= imem05_in[83:80];
    88: reg_0153 <= imem01_in[95:92];
    90: reg_0153 <= imem05_in[83:80];
    92: reg_0153 <= imem00_in[3:0];
    94: reg_0153 <= imem05_in[83:80];
    96: reg_0153 <= imem01_in[95:92];
    endcase
  end

  // REG#154の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0154 <= imem05_in[63:60];
    75: reg_0154 <= imem02_in[7:4];
    77: reg_0154 <= imem02_in[7:4];
    79: reg_0154 <= imem05_in[63:60];
    88: reg_0154 <= imem07_in[35:32];
    90: reg_0154 <= imem05_in[63:60];
    92: reg_0154 <= imem07_in[35:32];
    94: reg_0154 <= imem01_in[103:100];
    97: reg_0154 <= imem05_in[63:60];
    endcase
  end

  // REG#155の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0155 <= imem05_in[99:96];
    75: reg_0155 <= imem02_in[31:28];
    77: reg_0155 <= imem02_in[19:16];
    79: reg_0155 <= imem02_in[19:16];
    81: reg_0155 <= imem02_in[31:28];
    83: reg_0155 <= imem05_in[99:96];
    85: reg_0155 <= imem02_in[31:28];
    97: reg_0155 <= imem02_in[31:28];
    endcase
  end

  // REG#156の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0156 <= imem05_in[59:56];
    75: reg_0156 <= imem04_in[51:48];
    77: reg_0156 <= imem04_in[51:48];
    79: reg_0156 <= imem04_in[51:48];
    81: reg_0156 <= imem04_in[51:48];
    83: reg_0156 <= imem04_in[51:48];
    endcase
  end

  // REG#157の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0157 <= imem07_in[95:92];
    76: reg_0157 <= imem01_in[67:64];
    78: reg_0157 <= imem07_in[95:92];
    80: reg_0157 <= imem01_in[67:64];
    82: reg_0157 <= imem07_in[95:92];
    endcase
  end

  // REG#158の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0158 <= imem07_in[103:100];
    76: reg_0158 <= imem07_in[103:100];
    78: reg_0158 <= imem07_in[103:100];
    81: reg_0158 <= imem05_in[47:44];
    83: reg_0158 <= imem07_in[103:100];
    85: reg_0158 <= imem05_in[47:44];
    87: reg_0158 <= imem07_in[31:28];
    89: reg_0158 <= imem07_in[31:28];
    91: reg_0158 <= imem07_in[31:28];
    93: reg_0158 <= imem07_in[31:28];
    95: reg_0158 <= imem07_in[31:28];
    97: reg_0158 <= imem07_in[103:100];
    endcase
  end

  // REG#159の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0159 <= imem07_in[43:40];
    77: reg_0159 <= imem02_in[119:116];
    79: reg_0159 <= imem07_in[43:40];
    96: reg_0159 <= imem02_in[119:116];
    endcase
  end

  // REG#160の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0160 <= imem07_in[55:52];
    78: reg_0160 <= imem00_in[47:44];
    80: reg_0160 <= imem07_in[55:52];
    83: reg_0160 <= imem07_in[55:52];
    85: reg_0160 <= imem00_in[47:44];
    87: reg_0160 <= imem00_in[47:44];
    89: reg_0160 <= imem00_in[115:112];
    91: reg_0160 <= imem00_in[115:112];
    endcase
  end

  // REG#161の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0161 <= imem07_in[31:28];
    78: reg_0161 <= imem07_in[31:28];
    80: reg_0161 <= imem03_in[99:96];
    82: reg_0161 <= imem07_in[31:28];
    endcase
  end

  // REG#162の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0162 <= imem07_in[35:32];
    79: reg_0162 <= imem07_in[35:32];
    endcase
  end

  // REG#163の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0163 <= imem07_in[59:56];
    79: reg_0163 <= imem00_in[75:72];
    81: reg_0163 <= imem07_in[59:56];
    83: reg_0163 <= imem07_in[59:56];
    85: reg_0163 <= imem07_in[59:56];
    87: reg_0163 <= imem07_in[59:56];
    89: reg_0163 <= imem00_in[75:72];
    91: reg_0163 <= imem07_in[59:56];
    93: reg_0163 <= imem00_in[75:72];
    97: reg_0163 <= imem00_in[75:72];
    endcase
  end

  // REG#164の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0164 <= imem07_in[75:72];
    79: reg_0164 <= imem07_in[75:72];
    endcase
  end

  // REG#165の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0165 <= imem07_in[19:16];
    79: reg_0165 <= imem07_in[19:16];
    endcase
  end

  // REG#166の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0166 <= imem07_in[67:64];
    80: reg_0166 <= imem04_in[71:68];
    82: reg_0166 <= imem04_in[71:68];
    85: reg_0166 <= imem00_in[59:56];
    87: reg_0166 <= imem00_in[15:12];
    89: reg_0166 <= imem04_in[71:68];
    91: reg_0166 <= imem00_in[15:12];
    95: reg_0166 <= imem04_in[71:68];
    97: reg_0166 <= imem00_in[15:12];
    endcase
  end

  // REG#167の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0167 <= imem07_in[39:36];
    80: reg_0167 <= imem07_in[39:36];
    84: reg_0167 <= imem00_in[35:32];
    86: reg_0167 <= imem00_in[35:32];
    88: reg_0167 <= imem04_in[47:44];
    90: reg_0167 <= imem07_in[43:40];
    92: reg_0167 <= imem00_in[35:32];
    94: reg_0167 <= imem04_in[47:44];
    96: reg_0167 <= imem00_in[35:32];
    endcase
  end

  // REG#168の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0168 <= imem07_in[83:80];
    81: reg_0168 <= imem07_in[83:80];
    83: reg_0168 <= imem05_in[103:100];
    85: reg_0168 <= imem07_in[83:80];
    87: reg_0168 <= imem07_in[83:80];
    89: reg_0168 <= imem02_in[31:28];
    91: reg_0168 <= imem07_in[83:80];
    93: reg_0168 <= imem05_in[103:100];
    95: reg_0168 <= imem02_in[31:28];
    endcase
  end

  // REG#169の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0169 <= imem07_in[47:44];
    81: reg_0169 <= imem06_in[27:24];
    83: reg_0169 <= imem00_in[15:12];
    85: reg_0169 <= imem04_in[15:12];
    87: reg_0169 <= imem06_in[27:24];
    89: reg_0169 <= imem06_in[27:24];
    endcase
  end

  // REG#170の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0170 <= imem07_in[91:88];
    80: reg_0170 <= op1_13_out;
    84: reg_0170 <= imem07_in[91:88];
    86: reg_0170 <= imem07_in[91:88];
    87: reg_0170 <= op1_13_out;
    89: reg_0170 <= op1_13_out;
    92: reg_0170 <= imem07_in[91:88];
    93: reg_0170 <= op1_13_out;
    95: reg_0170 <= op1_13_out;
    endcase
  end

  // REG#171の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0171 <= imem07_in[111:108];
    82: reg_0171 <= imem07_in[111:108];
    endcase
  end

  // REG#172の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0172 <= imem07_in[15:12];
    82: reg_0172 <= imem07_in[15:12];
    endcase
  end

  // REG#173の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0173 <= imem07_in[107:104];
    81: reg_0173 <= imem07_in[107:104];
    83: reg_0173 <= imem01_in[71:68];
    85: reg_0173 <= imem01_in[71:68];
    87: reg_0173 <= imem01_in[71:68];
    89: reg_0173 <= imem01_in[71:68];
    91: reg_0173 <= imem07_in[107:104];
    93: reg_0173 <= imem01_in[71:68];
    97: reg_0173 <= imem01_in[71:68];
    endcase
  end

  // REG#174の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0174 <= imem07_in[3:0];
    82: reg_0174 <= imem07_in[3:0];
    endcase
  end

  // REG#175の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0175 <= imem07_in[7:4];
    82: reg_0175 <= imem07_in[7:4];
    endcase
  end

  // REG#176の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0176 <= imem07_in[99:96];
    81: reg_0176 <= imem07_in[99:96];
    83: reg_0176 <= imem06_in[43:40];
    85: reg_0176 <= imem06_in[43:40];
    87: reg_0176 <= imem07_in[99:96];
    89: reg_0176 <= imem07_in[99:96];
    91: reg_0176 <= imem01_in[75:72];
    93: reg_0176 <= imem07_in[99:96];
    95: reg_0176 <= imem01_in[75:72];
    endcase
  end

  // REG#177の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0177 <= imem07_in[71:68];
    81: reg_0177 <= imem07_in[71:68];
    83: reg_0177 <= imem07_in[71:68];
    85: reg_0177 <= imem07_in[71:68];
    87: reg_0177 <= imem07_in[71:68];
    89: reg_0177 <= imem06_in[63:60];
    endcase
  end

  // REG#178の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0178 <= imem07_in[87:84];
    81: reg_0178 <= imem07_in[87:84];
    83: reg_0178 <= imem03_in[107:104];
    85: reg_0178 <= imem05_in[11:8];
    87: reg_0178 <= imem05_in[11:8];
    95: reg_0178 <= imem03_in[107:104];
    endcase
  end

  // REG#179の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0179 <= imem07_in[27:24];
    82: reg_0179 <= imem07_in[27:24];
    endcase
  end

  // REG#180の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0180 <= imem07_in[11:8];
    82: reg_0180 <= imem07_in[11:8];
    endcase
  end

  // REG#181の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0181 <= imem07_in[23:20];
    82: reg_0181 <= imem07_in[23:20];
    endcase
  end

  // REG#182の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0182 <= imem07_in[51:48];
    82: reg_0182 <= imem07_in[51:48];
    endcase
  end

  // REG#183の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0183 <= imem07_in[63:60];
    82: reg_0183 <= imem07_in[63:60];
    endcase
  end

  // REG#184の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0184 <= imem07_in[115:112];
    82: reg_0184 <= imem07_in[115:112];
    endcase
  end

  // REG#185の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0185 <= imem07_in[79:76];
    82: reg_0185 <= imem07_in[79:76];
    96: reg_0185 <= imem07_in[79:76];
    endcase
  end

  // REG#186の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0186 <= imem00_in[59:56];
    89: reg_0186 <= imem00_in[59:56];
    91: reg_0186 <= imem00_in[59:56];
    endcase
  end

  // REG#187の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0187 <= imem00_in[27:24];
    90: reg_0187 <= imem00_in[27:24];
    93: reg_0187 <= imem00_in[83:80];
    95: reg_0187 <= imem00_in[83:80];
    endcase
  end

  // REG#188の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0188 <= imem00_in[39:36];
    91: reg_0188 <= imem00_in[39:36];
    93: reg_0188 <= imem02_in[11:8];
    96: reg_0188 <= imem02_in[11:8];
    endcase
  end

  // REG#189の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0189 <= imem00_in[23:20];
    92: reg_0189 <= imem00_in[23:20];
    93: reg_0189 <= op2_00_out;
    endcase
  end

  // REG#190の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0190 <= imem00_in[91:88];
    endcase
  end

  // REG#191の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0191 <= imem00_in[15:12];
    94: reg_0191 <= imem00_in[15:12];
    endcase
  end

  // REG#192の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0192 <= imem00_in[111:108];
    97: reg_0192 <= imem00_in[111:108];
    endcase
  end

  // REG#193の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0193 <= imem00_in[47:44];
    96: reg_0193 <= imem00_in[47:44];
    endcase
  end

  // REG#194の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0194 <= imem00_in[63:60];
    96: reg_0194 <= imem00_in[63:60];
    endcase
  end

  // REG#195の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0195 <= imem00_in[99:96];
    endcase
  end

  // REG#196の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0196 <= imem00_in[79:76];
    96: reg_0196 <= imem00_in[79:76];
    endcase
  end

  // REG#197の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0197 <= imem00_in[115:112];
    endcase
  end

  // REG#198の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0198 <= imem00_in[67:64];
    97: reg_0198 <= imem00_in[67:64];
    endcase
  end

  // REG#199の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0199 <= imem00_in[107:104];
    endcase
  end

  // REG#200の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0200 <= imem00_in[7:4];
    97: reg_0200 <= imem00_in[7:4];
    endcase
  end

  // REG#201の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0201 <= imem00_in[71:68];
    endcase
  end

  // REG#202の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0202 <= imem00_in[95:92];
    endcase
  end

  // REG#203の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0203 <= imem00_in[43:40];
    endcase
  end

  // REG#204の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0204 <= imem00_in[35:32];
    endcase
  end

  // REG#205の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0205 <= imem00_in[87:84];
    endcase
  end

  // REG#206の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0206 <= imem00_in[103:100];
    endcase
  end

  // REG#207の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0207 <= imem00_in[51:48];
    endcase
  end

  // REG#208の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0208 <= imem00_in[11:8];
    endcase
  end

  // REG#209の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0209 <= imem00_in[31:28];
    endcase
  end

  // REG#210の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0210 <= imem00_in[19:16];
    endcase
  end

  // REG#211の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0211 <= imem00_in[55:52];
    endcase
  end

  // REG#212の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0212 <= imem00_in[83:80];
    endcase
  end

  // REG#213の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0213 <= imem00_in[75:72];
    endcase
  end

  // REG#214の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0214 <= imem00_in[3:0];
    endcase
  end

  // REG#215の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0215 <= imem05_in[11:8];
    8: reg_0215 <= imem05_in[99:96];
    10: reg_0215 <= imem05_in[99:96];
    12: reg_0215 <= imem05_in[11:8];
    20: reg_0215 <= imem05_in[11:8];
    50: reg_0215 <= imem05_in[11:8];
    67: reg_0215 <= imem05_in[11:8];
    70: reg_0215 <= imem06_in[91:88];
    73: reg_0215 <= imem05_in[11:8];
    endcase
  end

  // REG#216の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0216 <= imem01_in[67:64];
    8: reg_0216 <= imem05_in[107:104];
    10: reg_0216 <= imem01_in[67:64];
    41: reg_0216 <= imem01_in[67:64];
    91: reg_0216 <= imem04_in[83:80];
    93: reg_0216 <= imem04_in[83:80];
    95: reg_0216 <= imem01_in[67:64];
    endcase
  end

  // REG#217の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0217 <= imem05_in[15:12];
    8: reg_0217 <= imem05_in[15:12];
    10: reg_0217 <= imem03_in[71:68];
    12: reg_0217 <= imem05_in[15:12];
    17: reg_0217 <= imem05_in[15:12];
    19: reg_0217 <= imem05_in[15:12];
    21: reg_0217 <= imem04_in[127:124];
    23: reg_0217 <= imem05_in[15:12];
    25: reg_0217 <= imem04_in[127:124];
    27: reg_0217 <= imem03_in[71:68];
    30: reg_0217 <= imem04_in[127:124];
    32: reg_0217 <= imem05_in[15:12];
    34: reg_0217 <= imem04_in[127:124];
    36: reg_0217 <= imem01_in[107:104];
    38: reg_0217 <= imem03_in[71:68];
    40: reg_0217 <= imem05_in[35:32];
    42: reg_0217 <= imem05_in[15:12];
    44: reg_0217 <= imem03_in[71:68];
    46: reg_0217 <= imem03_in[71:68];
    48: reg_0217 <= imem03_in[71:68];
    50: reg_0217 <= imem03_in[71:68];
    52: reg_0217 <= imem05_in[15:12];
    54: reg_0217 <= imem03_in[71:68];
    56: reg_0217 <= imem03_in[71:68];
    58: reg_0217 <= imem03_in[71:68];
    60: reg_0217 <= imem01_in[107:104];
    62: reg_0217 <= imem05_in[35:32];
    64: reg_0217 <= imem01_in[107:104];
    66: reg_0217 <= imem04_in[127:124];
    68: reg_0217 <= imem05_in[35:32];
    73: reg_0217 <= imem05_in[35:32];
    endcase
  end

  // REG#218の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0218 <= imem01_in[35:32];
    9: reg_0218 <= imem01_in[35:32];
    13: reg_0218 <= imem06_in[79:76];
    15: reg_0218 <= imem01_in[35:32];
    17: reg_0218 <= imem06_in[79:76];
    19: reg_0218 <= imem06_in[99:96];
    21: reg_0218 <= imem06_in[79:76];
    23: reg_0218 <= imem06_in[79:76];
    25: reg_0218 <= imem01_in[35:32];
    47: reg_0218 <= imem06_in[99:96];
    49: reg_0218 <= imem01_in[35:32];
    68: reg_0218 <= imem06_in[99:96];
    70: reg_0218 <= imem06_in[79:76];
    73: reg_0218 <= imem02_in[19:16];
    75: reg_0218 <= imem02_in[19:16];
    77: reg_0218 <= imem06_in[79:76];
    79: reg_0218 <= imem02_in[71:68];
    81: reg_0218 <= imem06_in[99:96];
    83: reg_0218 <= imem02_in[71:68];
    85: reg_0218 <= imem02_in[71:68];
    endcase
  end

  // REG#219の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0219 <= imem01_in[119:116];
    9: reg_0219 <= imem01_in[119:116];
    13: reg_0219 <= imem01_in[119:116];
    15: reg_0219 <= imem01_in[119:116];
    17: reg_0219 <= imem01_in[119:116];
    19: reg_0219 <= imem06_in[103:100];
    21: reg_0219 <= imem07_in[11:8];
    23: reg_0219 <= imem06_in[103:100];
    25: reg_0219 <= imem01_in[119:116];
    49: reg_0219 <= imem06_in[103:100];
    51: reg_0219 <= imem06_in[103:100];
    53: reg_0219 <= imem04_in[123:120];
    55: reg_0219 <= imem06_in[103:100];
    57: reg_0219 <= imem01_in[119:116];
    59: reg_0219 <= imem06_in[103:100];
    61: reg_0219 <= imem06_in[103:100];
    72: reg_0219 <= imem06_in[103:100];
    74: reg_0219 <= imem06_in[103:100];
    76: reg_0219 <= imem07_in[11:8];
    78: reg_0219 <= imem04_in[39:36];
    80: reg_0219 <= imem06_in[23:20];
    82: reg_0219 <= imem06_in[23:20];
    84: reg_0219 <= imem01_in[119:116];
    86: reg_0219 <= imem07_in[11:8];
    88: reg_0219 <= imem01_in[119:116];
    90: reg_0219 <= imem02_in[3:0];
    92: reg_0219 <= imem04_in[39:36];
    94: reg_0219 <= imem02_in[3:0];
    96: reg_0219 <= imem01_in[119:116];
    endcase
  end

  // REG#220の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0220 <= imem01_in[71:68];
    9: reg_0220 <= imem01_in[71:68];
    11: reg_0220 <= imem01_in[71:68];
    24: reg_0220 <= imem01_in[71:68];
    27: reg_0220 <= imem01_in[71:68];
    29: reg_0220 <= imem05_in[91:88];
    31: reg_0220 <= imem04_in[67:64];
    33: reg_0220 <= imem06_in[39:36];
    35: reg_0220 <= imem01_in[71:68];
    37: reg_0220 <= imem05_in[91:88];
    39: reg_0220 <= imem06_in[39:36];
    58: reg_0220 <= imem04_in[67:64];
    61: reg_0220 <= imem04_in[67:64];
    63: reg_0220 <= imem04_in[67:64];
    65: reg_0220 <= imem01_in[71:68];
    67: reg_0220 <= imem04_in[67:64];
    69: reg_0220 <= imem04_in[67:64];
    71: reg_0220 <= imem06_in[39:36];
    90: reg_0220 <= imem06_in[39:36];
    92: reg_0220 <= imem04_in[67:64];
    94: reg_0220 <= imem06_in[39:36];
    endcase
  end

  // REG#221の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0221 <= imem01_in[115:112];
    9: reg_0221 <= imem01_in[115:112];
    13: reg_0221 <= imem01_in[115:112];
    15: reg_0221 <= imem06_in[31:28];
    17: reg_0221 <= imem06_in[31:28];
    19: reg_0221 <= imem07_in[27:24];
    21: reg_0221 <= imem07_in[27:24];
    23: reg_0221 <= imem06_in[31:28];
    25: reg_0221 <= imem01_in[115:112];
    48: reg_0221 <= imem01_in[115:112];
    50: reg_0221 <= imem01_in[99:96];
    52: reg_0221 <= imem05_in[71:68];
    54: reg_0221 <= imem05_in[71:68];
    56: reg_0221 <= imem05_in[71:68];
    62: reg_0221 <= imem06_in[31:28];
    64: reg_0221 <= imem05_in[71:68];
    66: reg_0221 <= imem05_in[71:68];
    79: reg_0221 <= imem07_in[27:24];
    95: reg_0221 <= imem01_in[99:96];
    endcase
  end

  // REG#222の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0222 <= imem01_in[23:20];
    9: reg_0222 <= imem01_in[23:20];
    13: reg_0222 <= imem06_in[111:108];
    15: reg_0222 <= imem07_in[79:76];
    17: reg_0222 <= imem01_in[47:44];
    19: reg_0222 <= imem06_in[111:108];
    21: reg_0222 <= imem07_in[79:76];
    23: reg_0222 <= imem01_in[23:20];
    25: reg_0222 <= imem07_in[79:76];
    27: reg_0222 <= imem06_in[111:108];
    29: reg_0222 <= imem06_in[111:108];
    58: reg_0222 <= imem06_in[111:108];
    85: reg_0222 <= imem07_in[39:36];
    87: reg_0222 <= imem01_in[47:44];
    89: reg_0222 <= imem06_in[111:108];
    95: reg_0222 <= imem01_in[23:20];
    endcase
  end

  // REG#223の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0223 <= imem05_in[127:124];
    9: reg_0223 <= imem05_in[127:124];
    11: reg_0223 <= imem05_in[79:76];
    13: reg_0223 <= imem01_in[19:16];
    15: reg_0223 <= imem05_in[127:124];
    17: reg_0223 <= imem02_in[3:0];
    19: reg_0223 <= imem05_in[79:76];
    21: reg_0223 <= imem00_in[27:24];
    23: reg_0223 <= imem01_in[19:16];
    25: reg_0223 <= imem01_in[19:16];
    49: reg_0223 <= imem01_in[19:16];
    67: reg_0223 <= imem00_in[27:24];
    69: reg_0223 <= imem05_in[127:124];
    71: reg_0223 <= imem00_in[27:24];
    73: reg_0223 <= imem02_in[3:0];
    75: reg_0223 <= imem00_in[27:24];
    77: reg_0223 <= imem00_in[27:24];
    79: reg_0223 <= imem05_in[79:76];
    87: reg_0223 <= imem01_in[19:16];
    89: reg_0223 <= imem05_in[127:124];
    91: reg_0223 <= imem00_in[27:24];
    endcase
  end

  // REG#224の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0224 <= imem01_in[59:56];
    9: reg_0224 <= imem01_in[59:56];
    13: reg_0224 <= imem01_in[59:56];
    15: reg_0224 <= imem01_in[59:56];
    17: reg_0224 <= imem02_in[95:92];
    19: reg_0224 <= imem01_in[59:56];
    21: reg_0224 <= imem01_in[59:56];
    23: reg_0224 <= imem01_in[59:56];
    25: reg_0224 <= imem01_in[59:56];
    47: reg_0224 <= imem01_in[59:56];
    51: reg_0224 <= imem04_in[63:60];
    53: reg_0224 <= imem02_in[95:92];
    55: reg_0224 <= imem04_in[63:60];
    57: reg_0224 <= imem07_in[119:116];
    59: reg_0224 <= imem07_in[119:116];
    61: reg_0224 <= imem04_in[63:60];
    63: reg_0224 <= imem02_in[95:92];
    73: reg_0224 <= imem01_in[59:56];
    75: reg_0224 <= imem02_in[95:92];
    77: reg_0224 <= imem03_in[23:20];
    79: reg_0224 <= imem04_in[63:60];
    81: reg_0224 <= imem04_in[63:60];
    83: reg_0224 <= imem04_in[63:60];
    endcase
  end

  // REG#225の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0225 <= imem01_in[127:124];
    9: reg_0225 <= imem01_in[127:124];
    12: reg_0225 <= imem01_in[127:124];
    14: reg_0225 <= imem05_in[43:40];
    16: reg_0225 <= imem01_in[127:124];
    18: reg_0225 <= imem01_in[127:124];
    20: reg_0225 <= imem01_in[127:124];
    22: reg_0225 <= imem05_in[43:40];
    24: reg_0225 <= imem02_in[55:52];
    26: reg_0225 <= imem02_in[55:52];
    52: reg_0225 <= imem05_in[43:40];
    54: reg_0225 <= imem05_in[43:40];
    56: reg_0225 <= imem05_in[43:40];
    59: reg_0225 <= imem01_in[127:124];
    61: reg_0225 <= imem02_in[55:52];
    63: reg_0225 <= imem02_in[55:52];
    69: reg_0225 <= imem01_in[127:124];
    92: reg_0225 <= imem01_in[127:124];
    95: reg_0225 <= imem01_in[127:124];
    endcase
  end

  // REG#226の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0226 <= imem01_in[11:8];
    10: reg_0226 <= imem01_in[11:8];
    40: reg_0226 <= imem01_in[11:8];
    42: reg_0226 <= imem05_in[115:112];
    44: reg_0226 <= imem03_in[27:24];
    46: reg_0226 <= imem06_in[87:84];
    48: reg_0226 <= imem06_in[87:84];
    50: reg_0226 <= imem03_in[27:24];
    52: reg_0226 <= imem03_in[27:24];
    54: reg_0226 <= imem07_in[119:116];
    56: reg_0226 <= imem03_in[27:24];
    58: reg_0226 <= imem01_in[11:8];
    60: reg_0226 <= imem06_in[87:84];
    62: reg_0226 <= imem01_in[91:88];
    64: reg_0226 <= imem06_in[87:84];
    66: reg_0226 <= imem06_in[87:84];
    68: reg_0226 <= imem01_in[91:88];
    71: reg_0226 <= imem01_in[11:8];
    73: reg_0226 <= imem05_in[115:112];
    endcase
  end

  // REG#227の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0227 <= imem01_in[63:60];
    10: reg_0227 <= imem01_in[63:60];
    41: reg_0227 <= imem01_in[63:60];
    91: reg_0227 <= imem05_in[91:88];
    93: reg_0227 <= imem01_in[63:60];
    96: reg_0227 <= imem01_in[63:60];
    endcase
  end

  // REG#228の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0228 <= imem01_in[107:104];
    10: reg_0228 <= imem01_in[107:104];
    39: reg_0228 <= imem01_in[107:104];
    43: reg_0228 <= imem05_in[39:36];
    45: reg_0228 <= imem03_in[43:40];
    47: reg_0228 <= imem02_in[115:112];
    49: reg_0228 <= imem05_in[39:36];
    51: reg_0228 <= imem01_in[107:104];
    53: reg_0228 <= imem02_in[115:112];
    55: reg_0228 <= imem03_in[43:40];
    89: reg_0228 <= imem03_in[43:40];
    92: reg_0228 <= imem05_in[39:36];
    94: reg_0228 <= imem03_in[43:40];
    97: reg_0228 <= imem05_in[39:36];
    endcase
  end

  // REG#229の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0229 <= imem05_in[63:60];
    10: reg_0229 <= imem03_in[123:120];
    12: reg_0229 <= imem05_in[63:60];
    18: reg_0229 <= imem06_in[107:104];
    20: reg_0229 <= imem05_in[63:60];
    51: reg_0229 <= imem05_in[63:60];
    53: reg_0229 <= imem05_in[63:60];
    55: reg_0229 <= imem06_in[107:104];
    57: reg_0229 <= imem06_in[107:104];
    endcase
  end

  // REG#230の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0230 <= imem01_in[31:28];
    10: reg_0230 <= imem01_in[31:28];
    38: reg_0230 <= imem07_in[75:72];
    40: reg_0230 <= imem00_in[47:44];
    42: reg_0230 <= imem07_in[115:112];
    44: reg_0230 <= imem00_in[47:44];
    46: reg_0230 <= imem07_in[75:72];
    48: reg_0230 <= imem07_in[115:112];
    50: reg_0230 <= imem07_in[75:72];
    52: reg_0230 <= imem07_in[75:72];
    54: reg_0230 <= imem00_in[47:44];
    56: reg_0230 <= imem00_in[47:44];
    58: reg_0230 <= imem05_in[103:100];
    60: reg_0230 <= imem05_in[103:100];
    62: reg_0230 <= imem07_in[115:112];
    64: reg_0230 <= imem05_in[103:100];
    66: reg_0230 <= imem00_in[47:44];
    68: reg_0230 <= imem07_in[115:112];
    70: reg_0230 <= imem03_in[51:48];
    97: reg_0230 <= imem00_in[47:44];
    endcase
  end

  // REG#231の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0231 <= op1_00_out;
    9: reg_0231 <= op1_00_out;
    11: reg_0231 <= op1_00_out;
    13: reg_0231 <= op1_00_out;
    15: reg_0231 <= op1_00_out;
    17: reg_0231 <= op1_00_out;
    19: reg_0231 <= op1_00_out;
    21: reg_0231 <= op1_00_out;
    23: reg_0231 <= op1_00_out;
    25: reg_0231 <= op1_00_out;
    27: reg_0231 <= op1_00_out;
    29: reg_0231 <= op1_00_out;
    31: reg_0231 <= op1_00_out;
    33: reg_0231 <= op1_00_out;
    35: reg_0231 <= op1_00_out;
    37: reg_0231 <= op1_00_out;
    39: reg_0231 <= op1_00_out;
    41: reg_0231 <= op1_00_out;
    43: reg_0231 <= op1_00_out;
    45: reg_0231 <= op1_00_out;
    47: reg_0231 <= op1_00_out;
    49: reg_0231 <= op1_00_out;
    51: reg_0231 <= op1_00_out;
    53: reg_0231 <= op1_00_out;
    55: reg_0231 <= op1_00_out;
    57: reg_0231 <= op1_00_out;
    59: reg_0231 <= op1_00_out;
    61: reg_0231 <= op1_00_out;
    63: reg_0231 <= op1_00_out;
    65: reg_0231 <= op1_00_out;
    67: reg_0231 <= op1_00_out;
    69: reg_0231 <= op1_00_out;
    71: reg_0231 <= op1_00_out;
    73: reg_0231 <= op1_00_out;
    75: reg_0231 <= op1_00_out;
    77: reg_0231 <= op1_00_out;
    79: reg_0231 <= op1_00_out;
    81: reg_0231 <= op1_00_out;
    83: reg_0231 <= op1_00_out;
    85: reg_0231 <= op1_00_out;
    87: reg_0231 <= op1_00_out;
    89: reg_0231 <= op1_00_out;
    91: reg_0231 <= op1_00_out;
    93: reg_0231 <= op1_00_out;
    95: reg_0231 <= op1_00_out;
    97: reg_0231 <= op1_00_out;
    endcase
  end

  // REG#232の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0232 <= imem01_in[3:0];
    11: reg_0232 <= imem06_in[19:16];
    13: reg_0232 <= imem01_in[99:96];
    15: reg_0232 <= imem01_in[99:96];
    17: reg_0232 <= imem06_in[19:16];
    19: reg_0232 <= imem06_in[19:16];
    21: reg_0232 <= imem00_in[99:96];
    23: reg_0232 <= imem06_in[19:16];
    25: reg_0232 <= imem00_in[99:96];
    27: reg_0232 <= imem01_in[3:0];
    29: reg_0232 <= imem01_in[99:96];
    31: reg_0232 <= imem01_in[99:96];
    33: reg_0232 <= imem06_in[103:100];
    35: reg_0232 <= imem06_in[103:100];
    37: reg_0232 <= imem01_in[3:0];
    39: reg_0232 <= imem00_in[99:96];
    41: reg_0232 <= imem06_in[103:100];
    43: reg_0232 <= imem00_in[99:96];
    45: reg_0232 <= imem01_in[99:96];
    47: reg_0232 <= imem01_in[3:0];
    51: reg_0232 <= imem01_in[99:96];
    53: reg_0232 <= imem01_in[3:0];
    endcase
  end

  // REG#233の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0233 <= imem01_in[19:16];
    11: reg_0233 <= imem01_in[19:16];
    26: reg_0233 <= imem01_in[19:16];
    28: reg_0233 <= imem05_in[3:0];
    30: reg_0233 <= imem01_in[19:16];
    32: reg_0233 <= imem05_in[3:0];
    34: reg_0233 <= imem05_in[3:0];
    36: reg_0233 <= imem01_in[19:16];
    38: reg_0233 <= imem01_in[19:16];
    40: reg_0233 <= imem02_in[123:120];
    42: reg_0233 <= imem01_in[19:16];
    44: reg_0233 <= imem05_in[3:0];
    46: reg_0233 <= imem05_in[3:0];
    48: reg_0233 <= imem05_in[3:0];
    50: reg_0233 <= imem05_in[3:0];
    63: reg_0233 <= imem02_in[123:120];
    70: reg_0233 <= imem03_in[119:116];
    endcase
  end

  // REG#234の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0234 <= imem01_in[95:92];
    11: reg_0234 <= imem01_in[95:92];
    24: reg_0234 <= imem03_in[123:120];
    26: reg_0234 <= imem01_in[95:92];
    28: reg_0234 <= imem03_in[123:120];
    67: reg_0234 <= imem03_in[123:120];
    69: reg_0234 <= imem01_in[95:92];
    94: reg_0234 <= imem03_in[123:120];
    endcase
  end

  // REG#235の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0235 <= imem01_in[7:4];
    11: reg_0235 <= imem01_in[7:4];
    23: reg_0235 <= imem03_in[83:80];
    25: reg_0235 <= imem01_in[7:4];
    46: reg_0235 <= imem00_in[35:32];
    48: reg_0235 <= imem05_in[83:80];
    50: reg_0235 <= imem00_in[35:32];
    52: reg_0235 <= imem00_in[35:32];
    54: reg_0235 <= imem00_in[35:32];
    56: reg_0235 <= imem05_in[83:80];
    60: reg_0235 <= imem03_in[83:80];
    62: reg_0235 <= imem03_in[83:80];
    64: reg_0235 <= imem05_in[83:80];
    67: reg_0235 <= imem03_in[83:80];
    69: reg_0235 <= imem00_in[35:32];
    71: reg_0235 <= imem01_in[31:28];
    73: reg_0235 <= imem05_in[83:80];
    95: reg_0235 <= imem01_in[7:4];
    endcase
  end

  // REG#236の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0236 <= imem01_in[83:80];
    11: reg_0236 <= imem01_in[83:80];
    25: reg_0236 <= imem01_in[83:80];
    49: reg_0236 <= imem01_in[83:80];
    70: reg_0236 <= imem01_in[83:80];
    72: reg_0236 <= imem01_in[83:80];
    74: reg_0236 <= imem01_in[83:80];
    76: reg_0236 <= imem01_in[71:68];
    78: reg_0236 <= imem01_in[75:72];
    80: reg_0236 <= imem00_in[59:56];
    82: reg_0236 <= imem01_in[75:72];
    84: reg_0236 <= imem01_in[83:80];
    86: reg_0236 <= imem01_in[83:80];
    88: reg_0236 <= imem01_in[75:72];
    90: reg_0236 <= imem01_in[75:72];
    92: reg_0236 <= imem01_in[75:72];
    endcase
  end

  // REG#237の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0237 <= imem01_in[91:88];
    11: reg_0237 <= imem01_in[91:88];
    22: reg_0237 <= imem01_in[91:88];
    24: reg_0237 <= imem05_in[75:72];
    26: reg_0237 <= imem01_in[91:88];
    28: reg_0237 <= imem05_in[75:72];
    30: reg_0237 <= imem01_in[91:88];
    32: reg_0237 <= imem05_in[75:72];
    34: reg_0237 <= imem01_in[91:88];
    36: reg_0237 <= imem05_in[87:84];
    38: reg_0237 <= imem05_in[87:84];
    40: reg_0237 <= imem05_in[75:72];
    42: reg_0237 <= imem05_in[87:84];
    44: reg_0237 <= imem05_in[87:84];
    46: reg_0237 <= imem05_in[87:84];
    48: reg_0237 <= imem05_in[75:72];
    50: reg_0237 <= imem05_in[87:84];
    61: reg_0237 <= imem05_in[75:72];
    66: reg_0237 <= imem05_in[87:84];
    80: reg_0237 <= imem01_in[103:100];
    82: reg_0237 <= imem00_in[67:64];
    84: reg_0237 <= imem05_in[75:72];
    86: reg_0237 <= imem05_in[87:84];
    88: reg_0237 <= imem05_in[75:72];
    90: reg_0237 <= imem05_in[75:72];
    92: reg_0237 <= imem01_in[91:88];
    endcase
  end

  // REG#238の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0238 <= imem01_in[111:108];
    11: reg_0238 <= imem01_in[111:108];
    25: reg_0238 <= imem01_in[111:108];
    49: reg_0238 <= imem01_in[111:108];
    70: reg_0238 <= imem03_in[7:4];
    endcase
  end

  // REG#239の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0239 <= imem01_in[43:40];
    11: reg_0239 <= imem01_in[43:40];
    25: reg_0239 <= imem01_in[43:40];
    46: reg_0239 <= imem00_in[59:56];
    48: reg_0239 <= imem00_in[59:56];
    50: reg_0239 <= imem03_in[43:40];
    52: reg_0239 <= imem06_in[71:68];
    54: reg_0239 <= imem00_in[87:84];
    56: reg_0239 <= imem06_in[71:68];
    58: reg_0239 <= imem00_in[59:56];
    60: reg_0239 <= imem00_in[87:84];
    62: reg_0239 <= imem01_in[43:40];
    64: reg_0239 <= imem00_in[59:56];
    66: reg_0239 <= imem06_in[71:68];
    68: reg_0239 <= imem00_in[59:56];
    70: reg_0239 <= imem03_in[43:40];
    97: reg_0239 <= imem01_in[43:40];
    endcase
  end

  // REG#240の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0240 <= imem01_in[55:52];
    11: reg_0240 <= imem01_in[55:52];
    25: reg_0240 <= imem01_in[55:52];
    44: reg_0240 <= imem03_in[107:104];
    46: reg_0240 <= imem01_in[111:108];
    48: reg_0240 <= imem03_in[107:104];
    50: reg_0240 <= imem01_in[111:108];
    52: reg_0240 <= imem01_in[111:108];
    55: reg_0240 <= imem03_in[107:104];
    87: reg_0240 <= imem03_in[107:104];
    89: reg_0240 <= imem03_in[107:104];
    92: reg_0240 <= imem01_in[55:52];
    97: reg_0240 <= imem01_in[55:52];
    endcase
  end

  // REG#241の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0241 <= imem05_in[47:44];
    11: reg_0241 <= imem06_in[43:40];
    13: reg_0241 <= imem05_in[47:44];
    15: reg_0241 <= imem05_in[47:44];
    17: reg_0241 <= imem06_in[43:40];
    19: reg_0241 <= imem06_in[43:40];
    21: reg_0241 <= imem01_in[51:48];
    23: reg_0241 <= imem05_in[47:44];
    25: reg_0241 <= imem06_in[43:40];
    27: reg_0241 <= imem05_in[47:44];
    29: reg_0241 <= imem01_in[51:48];
    31: reg_0241 <= imem05_in[123:120];
    33: reg_0241 <= imem01_in[51:48];
    35: reg_0241 <= imem05_in[123:120];
    37: reg_0241 <= imem06_in[43:40];
    61: reg_0241 <= imem06_in[43:40];
    72: reg_0241 <= imem01_in[51:48];
    74: reg_0241 <= imem01_in[51:48];
    76: reg_0241 <= imem06_in[43:40];
    78: reg_0241 <= imem05_in[47:44];
    80: reg_0241 <= imem06_in[43:40];
    82: reg_0241 <= imem05_in[47:44];
    84: reg_0241 <= imem00_in[47:44];
    86: reg_0241 <= imem05_in[47:44];
    89: reg_0241 <= imem05_in[47:44];
    91: reg_0241 <= imem05_in[123:120];
    93: reg_0241 <= imem00_in[47:44];
    95: reg_0241 <= imem05_in[123:120];
    97: reg_0241 <= imem05_in[123:120];
    endcase
  end

  // REG#242の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0242 <= imem01_in[51:48];
    11: reg_0242 <= imem01_in[51:48];
    25: reg_0242 <= imem01_in[51:48];
    49: reg_0242 <= imem01_in[51:48];
    68: reg_0242 <= imem01_in[51:48];
    71: reg_0242 <= imem01_in[63:60];
    73: reg_0242 <= imem01_in[51:48];
    75: reg_0242 <= imem01_in[63:60];
    77: reg_0242 <= imem03_in[31:28];
    79: reg_0242 <= imem03_in[31:28];
    81: reg_0242 <= imem01_in[63:60];
    83: reg_0242 <= imem03_in[31:28];
    85: reg_0242 <= imem01_in[63:60];
    87: reg_0242 <= imem01_in[51:48];
    90: reg_0242 <= imem03_in[31:28];
    endcase
  end

  // REG#243の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0243 <= imem05_in[71:68];
    11: reg_0243 <= imem06_in[87:84];
    13: reg_0243 <= imem05_in[71:68];
    15: reg_0243 <= imem06_in[87:84];
    17: reg_0243 <= imem05_in[71:68];
    19: reg_0243 <= imem05_in[71:68];
    21: reg_0243 <= imem01_in[55:52];
    23: reg_0243 <= imem05_in[71:68];
    25: reg_0243 <= imem04_in[19:16];
    27: reg_0243 <= imem04_in[19:16];
    29: reg_0243 <= imem06_in[87:84];
    59: reg_0243 <= imem04_in[19:16];
    endcase
  end

  // REG#244の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0244 <= imem05_in[95:92];
    11: reg_0244 <= imem05_in[95:92];
    14: reg_0244 <= imem05_in[95:92];
    16: reg_0244 <= imem05_in[95:92];
    18: reg_0244 <= imem05_in[95:92];
    20: reg_0244 <= imem05_in[95:92];
    41: reg_0244 <= imem06_in[39:36];
    43: reg_0244 <= imem06_in[39:36];
    45: reg_0244 <= imem06_in[39:36];
    47: reg_0244 <= imem06_in[39:36];
    49: reg_0244 <= imem05_in[95:92];
    51: reg_0244 <= imem06_in[39:36];
    53: reg_0244 <= imem05_in[95:92];
    55: reg_0244 <= imem04_in[103:100];
    57: reg_0244 <= imem06_in[39:36];
    endcase
  end

  // REG#245の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0245 <= imem01_in[103:100];
    11: reg_0245 <= imem01_in[103:100];
    24: reg_0245 <= imem01_in[103:100];
    27: reg_0245 <= imem03_in[67:64];
    29: reg_0245 <= imem03_in[67:64];
    31: reg_0245 <= imem03_in[67:64];
    55: reg_0245 <= imem03_in[67:64];
    83: reg_0245 <= imem01_in[91:88];
    85: reg_0245 <= imem01_in[91:88];
    87: reg_0245 <= imem03_in[67:64];
    89: reg_0245 <= imem03_in[67:64];
    92: reg_0245 <= imem01_in[103:100];
    endcase
  end

  // REG#246の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0246 <= imem01_in[27:24];
    11: reg_0246 <= imem01_in[27:24];
    26: reg_0246 <= imem03_in[115:112];
    28: reg_0246 <= imem03_in[115:112];
    67: reg_0246 <= imem01_in[27:24];
    69: reg_0246 <= imem01_in[27:24];
    94: reg_0246 <= imem01_in[27:24];
    96: reg_0246 <= imem01_in[27:24];
    endcase
  end

  // REG#247の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0247 <= imem01_in[75:72];
    11: reg_0247 <= imem01_in[75:72];
    25: reg_0247 <= imem01_in[75:72];
    48: reg_0247 <= imem01_in[75:72];
    50: reg_0247 <= imem01_in[75:72];
    52: reg_0247 <= imem07_in[91:88];
    54: reg_0247 <= imem01_in[19:16];
    56: reg_0247 <= imem01_in[75:72];
    58: reg_0247 <= imem01_in[19:16];
    60: reg_0247 <= imem01_in[75:72];
    62: reg_0247 <= imem01_in[75:72];
    64: reg_0247 <= imem07_in[91:88];
    66: reg_0247 <= imem07_in[91:88];
    68: reg_0247 <= imem01_in[19:16];
    71: reg_0247 <= imem01_in[19:16];
    73: reg_0247 <= imem01_in[75:72];
    75: reg_0247 <= imem07_in[91:88];
    77: reg_0247 <= imem01_in[19:16];
    79: reg_0247 <= imem07_in[91:88];
    endcase
  end

  // REG#248の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0248 <= imem01_in[87:84];
    11: reg_0248 <= imem01_in[87:84];
    25: reg_0248 <= imem01_in[87:84];
    44: reg_0248 <= imem02_in[83:80];
    46: reg_0248 <= imem02_in[115:112];
    48: reg_0248 <= imem02_in[83:80];
    50: reg_0248 <= imem03_in[111:108];
    52: reg_0248 <= imem02_in[83:80];
    endcase
  end

  // REG#249の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0249 <= imem01_in[123:120];
    11: reg_0249 <= imem01_in[123:120];
    25: reg_0249 <= imem01_in[123:120];
    49: reg_0249 <= imem01_in[123:120];
    68: reg_0249 <= imem01_in[123:120];
    71: reg_0249 <= imem01_in[83:80];
    73: reg_0249 <= imem04_in[19:16];
    75: reg_0249 <= imem04_in[19:16];
    77: reg_0249 <= imem01_in[83:80];
    79: reg_0249 <= imem01_in[83:80];
    82: reg_0249 <= imem02_in[19:16];
    84: reg_0249 <= imem01_in[123:120];
    86: reg_0249 <= imem00_in[83:80];
    88: reg_0249 <= imem04_in[19:16];
    90: reg_0249 <= imem01_in[83:80];
    92: reg_0249 <= imem01_in[123:120];
    endcase
  end

  // REG#250の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0250 <= imem05_in[35:32];
    12: reg_0250 <= imem05_in[35:32];
    21: reg_0250 <= imem01_in[123:120];
    23: reg_0250 <= imem05_in[35:32];
    25: reg_0250 <= imem00_in[67:64];
    27: reg_0250 <= imem01_in[123:120];
    29: reg_0250 <= imem00_in[67:64];
    31: reg_0250 <= imem00_in[67:64];
    33: reg_0250 <= imem07_in[23:20];
    35: reg_0250 <= imem00_in[79:76];
    37: reg_0250 <= imem05_in[35:32];
    39: reg_0250 <= imem01_in[123:120];
    43: reg_0250 <= imem07_in[23:20];
    endcase
  end

  // REG#251の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0251 <= imem05_in[67:64];
    12: reg_0251 <= imem05_in[67:64];
    20: reg_0251 <= imem05_in[67:64];
    51: reg_0251 <= imem04_in[87:84];
    53: reg_0251 <= imem05_in[67:64];
    55: reg_0251 <= imem05_in[67:64];
    57: reg_0251 <= imem05_in[67:64];
    59: reg_0251 <= imem04_in[87:84];
    95: reg_0251 <= imem05_in[67:64];
    endcase
  end

  // REG#252の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0252 <= imem05_in[51:48];
    12: reg_0252 <= imem05_in[51:48];
    20: reg_0252 <= imem05_in[51:48];
    48: reg_0252 <= imem06_in[43:40];
    50: reg_0252 <= imem05_in[51:48];
    65: reg_0252 <= imem05_in[51:48];
    67: reg_0252 <= imem05_in[51:48];
    70: reg_0252 <= imem05_in[51:48];
    72: reg_0252 <= imem06_in[67:64];
    74: reg_0252 <= imem05_in[51:48];
    endcase
  end

  // REG#253の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0253 <= imem05_in[115:112];
    12: reg_0253 <= imem05_in[115:112];
    21: reg_0253 <= imem04_in[23:20];
    23: reg_0253 <= imem05_in[115:112];
    25: reg_0253 <= imem00_in[87:84];
    27: reg_0253 <= imem00_in[87:84];
    29: reg_0253 <= imem00_in[87:84];
    31: reg_0253 <= imem04_in[23:20];
    33: reg_0253 <= imem00_in[87:84];
    35: reg_0253 <= imem00_in[87:84];
    37: reg_0253 <= imem01_in[119:116];
    39: reg_0253 <= imem00_in[87:84];
    41: reg_0253 <= imem00_in[87:84];
    43: reg_0253 <= imem05_in[115:112];
    45: reg_0253 <= imem03_in[55:52];
    47: reg_0253 <= imem00_in[87:84];
    49: reg_0253 <= imem01_in[119:116];
    69: reg_0253 <= imem04_in[23:20];
    71: reg_0253 <= imem05_in[115:112];
    73: reg_0253 <= imem03_in[55:52];
    75: reg_0253 <= imem05_in[115:112];
    77: reg_0253 <= imem00_in[87:84];
    79: reg_0253 <= imem00_in[87:84];
    81: reg_0253 <= imem03_in[55:52];
    83: reg_0253 <= imem00_in[87:84];
    85: reg_0253 <= imem03_in[55:52];
    87: reg_0253 <= imem04_in[23:20];
    89: reg_0253 <= imem03_in[55:52];
    91: reg_0253 <= imem01_in[119:116];
    93: reg_0253 <= imem01_in[119:116];
    95: reg_0253 <= imem03_in[55:52];
    endcase
  end

  // REG#254の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0254 <= imem05_in[103:100];
    12: reg_0254 <= imem05_in[103:100];
    20: reg_0254 <= imem05_in[103:100];
    51: reg_0254 <= imem05_in[103:100];
    53: reg_0254 <= imem05_in[103:100];
    55: reg_0254 <= imem05_in[103:100];
    57: reg_0254 <= imem00_in[95:92];
    59: reg_0254 <= imem00_in[95:92];
    61: reg_0254 <= imem05_in[103:100];
    65: reg_0254 <= imem00_in[31:28];
    67: reg_0254 <= imem02_in[15:12];
    69: reg_0254 <= imem00_in[31:28];
    71: reg_0254 <= imem07_in[107:104];
    73: reg_0254 <= imem00_in[95:92];
    75: reg_0254 <= imem02_in[15:12];
    77: reg_0254 <= imem02_in[15:12];
    79: reg_0254 <= imem00_in[31:28];
    82: reg_0254 <= imem00_in[31:28];
    84: reg_0254 <= imem00_in[31:28];
    86: reg_0254 <= imem05_in[103:100];
    88: reg_0254 <= imem05_in[103:100];
    90: reg_0254 <= imem02_in[15:12];
    92: reg_0254 <= imem05_in[103:100];
    94: reg_0254 <= imem05_in[103:100];
    96: reg_0254 <= imem05_in[103:100];
    endcase
  end

  // REG#255の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0255 <= imem05_in[111:108];
    12: reg_0255 <= imem05_in[111:108];
    21: reg_0255 <= imem05_in[11:8];
    23: reg_0255 <= imem05_in[111:108];
    25: reg_0255 <= imem05_in[11:8];
    27: reg_0255 <= imem05_in[11:8];
    29: reg_0255 <= imem07_in[111:108];
    31: reg_0255 <= imem05_in[11:8];
    33: reg_0255 <= imem05_in[11:8];
    35: reg_0255 <= imem07_in[111:108];
    37: reg_0255 <= imem07_in[111:108];
    39: reg_0255 <= imem05_in[111:108];
    41: reg_0255 <= imem05_in[11:8];
    43: reg_0255 <= imem05_in[11:8];
    45: reg_0255 <= imem07_in[111:108];
    47: reg_0255 <= imem05_in[11:8];
    49: reg_0255 <= imem05_in[111:108];
    52: reg_0255 <= imem05_in[11:8];
    54: reg_0255 <= imem05_in[11:8];
    56: reg_0255 <= imem05_in[11:8];
    62: reg_0255 <= imem05_in[111:108];
    64: reg_0255 <= imem05_in[111:108];
    66: reg_0255 <= imem05_in[11:8];
    78: reg_0255 <= imem02_in[127:124];
    80: reg_0255 <= imem02_in[127:124];
    82: reg_0255 <= imem02_in[51:48];
    84: reg_0255 <= imem02_in[51:48];
    endcase
  end

  // REG#256の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0256 <= imem05_in[39:36];
    12: reg_0256 <= imem05_in[39:36];
    16: reg_0256 <= imem07_in[91:88];
    18: reg_0256 <= imem07_in[19:16];
    20: reg_0256 <= imem05_in[39:36];
    51: reg_0256 <= imem07_in[19:16];
    53: reg_0256 <= imem05_in[39:36];
    55: reg_0256 <= imem07_in[19:16];
    57: reg_0256 <= imem07_in[91:88];
    59: reg_0256 <= imem07_in[19:16];
    61: reg_0256 <= imem07_in[91:88];
    63: reg_0256 <= imem05_in[123:120];
    65: reg_0256 <= imem05_in[123:120];
    69: reg_0256 <= imem07_in[19:16];
    71: reg_0256 <= imem07_in[91:88];
    73: reg_0256 <= imem05_in[123:120];
    endcase
  end

  // REG#257の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0257 <= imem05_in[75:72];
    12: reg_0257 <= imem03_in[91:88];
    14: reg_0257 <= imem05_in[67:64];
    16: reg_0257 <= imem03_in[91:88];
    18: reg_0257 <= imem05_in[67:64];
    20: reg_0257 <= imem05_in[75:72];
    49: reg_0257 <= imem05_in[67:64];
    51: reg_0257 <= imem06_in[27:24];
    53: reg_0257 <= imem03_in[91:88];
    55: reg_0257 <= imem06_in[27:24];
    57: reg_0257 <= imem03_in[91:88];
    59: reg_0257 <= imem06_in[27:24];
    61: reg_0257 <= imem06_in[27:24];
    69: reg_0257 <= imem05_in[75:72];
    71: reg_0257 <= imem05_in[75:72];
    73: reg_0257 <= imem00_in[91:88];
    75: reg_0257 <= imem03_in[91:88];
    77: reg_0257 <= imem00_in[91:88];
    79: reg_0257 <= imem00_in[91:88];
    81: reg_0257 <= imem05_in[67:64];
    83: reg_0257 <= imem03_in[91:88];
    85: reg_0257 <= imem05_in[67:64];
    87: reg_0257 <= imem05_in[75:72];
    endcase
  end

  // REG#258の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0258 <= imem05_in[79:76];
    12: reg_0258 <= imem05_in[79:76];
    19: reg_0258 <= imem07_in[123:120];
    21: reg_0258 <= imem00_in[7:4];
    23: reg_0258 <= imem07_in[123:120];
    25: reg_0258 <= imem07_in[123:120];
    27: reg_0258 <= imem05_in[79:76];
    29: reg_0258 <= imem05_in[79:76];
    31: reg_0258 <= imem05_in[79:76];
    33: reg_0258 <= imem07_in[123:120];
    35: reg_0258 <= imem00_in[7:4];
    37: reg_0258 <= imem05_in[51:48];
    39: reg_0258 <= imem05_in[79:76];
    41: reg_0258 <= imem05_in[51:48];
    43: reg_0258 <= imem05_in[51:48];
    45: reg_0258 <= imem05_in[51:48];
    47: reg_0258 <= imem05_in[79:76];
    49: reg_0258 <= imem05_in[51:48];
    52: reg_0258 <= imem00_in[7:4];
    54: reg_0258 <= imem07_in[123:120];
    56: reg_0258 <= imem07_in[123:120];
    58: reg_0258 <= imem00_in[7:4];
    60: reg_0258 <= imem05_in[79:76];
    62: reg_0258 <= imem00_in[7:4];
    64: reg_0258 <= imem07_in[123:120];
    66: reg_0258 <= imem00_in[7:4];
    68: reg_0258 <= imem00_in[7:4];
    70: reg_0258 <= imem00_in[7:4];
    72: reg_0258 <= imem00_in[7:4];
    74: reg_0258 <= imem05_in[79:76];
    96: reg_0258 <= imem00_in[7:4];
    endcase
  end

  // REG#259の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0259 <= imem05_in[27:24];
    13: reg_0259 <= imem04_in[55:52];
    15: reg_0259 <= imem05_in[27:24];
    17: reg_0259 <= imem05_in[27:24];
    19: reg_0259 <= imem04_in[55:52];
    43: reg_0259 <= imem04_in[55:52];
    45: reg_0259 <= imem04_in[55:52];
    48: reg_0259 <= imem04_in[55:52];
    50: reg_0259 <= imem05_in[27:24];
    66: reg_0259 <= imem05_in[27:24];
    79: reg_0259 <= imem03_in[75:72];
    81: reg_0259 <= imem03_in[75:72];
    83: reg_0259 <= imem03_in[75:72];
    85: reg_0259 <= imem05_in[27:24];
    87: reg_0259 <= imem05_in[27:24];
    endcase
  end

  // REG#260の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0260 <= imem05_in[83:80];
    13: reg_0260 <= imem04_in[59:56];
    15: reg_0260 <= imem04_in[59:56];
    17: reg_0260 <= imem04_in[59:56];
    20: reg_0260 <= imem05_in[83:80];
    50: reg_0260 <= imem00_in[47:44];
    52: reg_0260 <= imem04_in[59:56];
    54: reg_0260 <= imem04_in[59:56];
    56: reg_0260 <= imem02_in[67:64];
    58: reg_0260 <= imem05_in[83:80];
    60: reg_0260 <= imem05_in[83:80];
    63: reg_0260 <= imem02_in[67:64];
    72: reg_0260 <= imem02_in[67:64];
    85: reg_0260 <= imem05_in[83:80];
    87: reg_0260 <= imem05_in[83:80];
    endcase
  end

  // REG#261の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0261 <= imem05_in[107:104];
    13: reg_0261 <= imem04_in[111:108];
    15: reg_0261 <= imem02_in[67:64];
    17: reg_0261 <= imem05_in[107:104];
    19: reg_0261 <= imem05_in[107:104];
    21: reg_0261 <= imem02_in[67:64];
    77: reg_0261 <= imem07_in[39:36];
    79: reg_0261 <= imem02_in[67:64];
    81: reg_0261 <= imem02_in[67:64];
    83: reg_0261 <= imem02_in[67:64];
    86: reg_0261 <= imem02_in[67:64];
    88: reg_0261 <= imem05_in[107:104];
    90: reg_0261 <= imem04_in[31:28];
    92: reg_0261 <= imem02_in[67:64];
    94: reg_0261 <= imem04_in[31:28];
    96: reg_0261 <= imem07_in[39:36];
    endcase
  end

  // REG#262の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0262 <= imem05_in[19:16];
    13: reg_0262 <= imem06_in[71:68];
    15: reg_0262 <= imem02_in[91:88];
    17: reg_0262 <= imem02_in[91:88];
    19: reg_0262 <= imem00_in[91:88];
    21: reg_0262 <= imem05_in[19:16];
    23: reg_0262 <= imem00_in[91:88];
    25: reg_0262 <= imem06_in[71:68];
    27: reg_0262 <= imem00_in[91:88];
    29: reg_0262 <= imem05_in[19:16];
    31: reg_0262 <= imem00_in[91:88];
    33: reg_0262 <= imem00_in[91:88];
    35: reg_0262 <= imem02_in[55:52];
    37: reg_0262 <= imem05_in[19:16];
    39: reg_0262 <= imem00_in[91:88];
    41: reg_0262 <= imem06_in[51:48];
    43: reg_0262 <= imem02_in[55:52];
    45: reg_0262 <= imem06_in[71:68];
    47: reg_0262 <= imem02_in[55:52];
    49: reg_0262 <= imem05_in[19:16];
    51: reg_0262 <= imem05_in[19:16];
    53: reg_0262 <= imem02_in[55:52];
    55: reg_0262 <= imem02_in[55:52];
    57: reg_0262 <= imem06_in[71:68];
    90: reg_0262 <= imem06_in[71:68];
    92: reg_0262 <= imem06_in[71:68];
    94: reg_0262 <= imem05_in[19:16];
    96: reg_0262 <= imem06_in[51:48];
    endcase
  end

  // REG#263の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0263 <= imem05_in[119:116];
    13: reg_0263 <= imem06_in[115:112];
    15: reg_0263 <= imem06_in[115:112];
    17: reg_0263 <= imem02_in[123:120];
    19: reg_0263 <= imem05_in[119:116];
    21: reg_0263 <= imem00_in[63:60];
    23: reg_0263 <= imem00_in[63:60];
    25: reg_0263 <= imem05_in[119:116];
    27: reg_0263 <= imem05_in[119:116];
    29: reg_0263 <= imem02_in[123:120];
    31: reg_0263 <= imem05_in[119:116];
    33: reg_0263 <= imem05_in[119:116];
    35: reg_0263 <= imem05_in[119:116];
    37: reg_0263 <= imem06_in[115:112];
    61: reg_0263 <= imem06_in[115:112];
    70: reg_0263 <= imem05_in[119:116];
    72: reg_0263 <= imem00_in[63:60];
    74: reg_0263 <= imem06_in[115:112];
    76: reg_0263 <= imem00_in[63:60];
    78: reg_0263 <= imem05_in[119:116];
    81: reg_0263 <= imem05_in[119:116];
    83: reg_0263 <= imem05_in[119:116];
    85: reg_0263 <= imem06_in[115:112];
    88: reg_0263 <= imem02_in[123:120];
    90: reg_0263 <= imem06_in[115:112];
    92: reg_0263 <= imem02_in[123:120];
    94: reg_0263 <= imem06_in[115:112];
    97: reg_0263 <= imem02_in[123:120];
    endcase
  end

  // REG#264の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0264 <= imem05_in[59:56];
    13: reg_0264 <= imem07_in[51:48];
    15: reg_0264 <= imem03_in[71:68];
    17: reg_0264 <= imem07_in[51:48];
    19: reg_0264 <= imem05_in[59:56];
    21: reg_0264 <= imem07_in[51:48];
    23: reg_0264 <= imem03_in[71:68];
    25: reg_0264 <= imem07_in[51:48];
    27: reg_0264 <= imem06_in[71:68];
    29: reg_0264 <= imem06_in[71:68];
    59: reg_0264 <= imem05_in[59:56];
    61: reg_0264 <= imem06_in[71:68];
    71: reg_0264 <= imem05_in[59:56];
    73: reg_0264 <= imem07_in[51:48];
    75: reg_0264 <= imem07_in[51:48];
    78: reg_0264 <= imem03_in[71:68];
    80: reg_0264 <= imem06_in[71:68];
    82: reg_0264 <= imem05_in[59:56];
    84: reg_0264 <= imem06_in[71:68];
    86: reg_0264 <= imem06_in[71:68];
    94: reg_0264 <= imem07_in[51:48];
    97: reg_0264 <= imem06_in[71:68];
    endcase
  end

  // REG#265の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0265 <= imem05_in[91:88];
    13: reg_0265 <= imem07_in[111:108];
    15: reg_0265 <= imem04_in[35:32];
    17: reg_0265 <= imem04_in[35:32];
    20: reg_0265 <= imem07_in[111:108];
    22: reg_0265 <= imem07_in[111:108];
    24: reg_0265 <= imem04_in[35:32];
    75: reg_0265 <= imem07_in[111:108];
    79: reg_0265 <= imem05_in[91:88];
    87: reg_0265 <= imem07_in[111:108];
    90: reg_0265 <= imem07_in[111:108];
    92: reg_0265 <= imem04_in[35:32];
    94: reg_0265 <= imem07_in[111:108];
    96: reg_0265 <= imem04_in[35:32];
    endcase
  end

  // REG#266の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0266 <= imem05_in[123:120];
    13: reg_0266 <= imem00_in[15:12];
    15: reg_0266 <= imem00_in[15:12];
    17: reg_0266 <= imem03_in[55:52];
    19: reg_0266 <= imem05_in[123:120];
    21: reg_0266 <= imem00_in[15:12];
    23: reg_0266 <= imem03_in[123:120];
    25: reg_0266 <= imem03_in[55:52];
    27: reg_0266 <= imem03_in[123:120];
    30: reg_0266 <= imem03_in[123:120];
    32: reg_0266 <= imem07_in[71:68];
    34: reg_0266 <= imem07_in[71:68];
    36: reg_0266 <= imem07_in[71:68];
    38: reg_0266 <= imem07_in[71:68];
    40: reg_0266 <= imem03_in[55:52];
    42: reg_0266 <= imem05_in[123:120];
    44: reg_0266 <= imem05_in[123:120];
    46: reg_0266 <= imem05_in[123:120];
    48: reg_0266 <= imem00_in[15:12];
    50: reg_0266 <= imem07_in[71:68];
    52: reg_0266 <= imem03_in[55:52];
    54: reg_0266 <= imem07_in[71:68];
    56: reg_0266 <= imem03_in[123:120];
    58: reg_0266 <= imem07_in[71:68];
    60: reg_0266 <= imem07_in[71:68];
    62: reg_0266 <= imem03_in[123:120];
    64: reg_0266 <= imem05_in[123:120];
    68: reg_0266 <= imem07_in[71:68];
    70: reg_0266 <= imem03_in[123:120];
    endcase
  end

  // REG#267の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0267 <= imem05_in[3:0];
    13: reg_0267 <= imem00_in[43:40];
    15: reg_0267 <= imem06_in[59:56];
    17: reg_0267 <= imem05_in[3:0];
    19: reg_0267 <= imem00_in[43:40];
    21: reg_0267 <= imem04_in[27:24];
    23: reg_0267 <= imem00_in[43:40];
    25: reg_0267 <= imem03_in[47:44];
    27: reg_0267 <= imem03_in[47:44];
    29: reg_0267 <= imem05_in[3:0];
    31: reg_0267 <= imem00_in[43:40];
    33: reg_0267 <= imem03_in[47:44];
    35: reg_0267 <= imem00_in[43:40];
    37: reg_0267 <= imem05_in[3:0];
    39: reg_0267 <= imem03_in[47:44];
    41: reg_0267 <= imem03_in[47:44];
    43: reg_0267 <= imem03_in[47:44];
    45: reg_0267 <= imem05_in[3:0];
    47: reg_0267 <= imem05_in[3:0];
    49: reg_0267 <= imem03_in[47:44];
    51: reg_0267 <= imem06_in[59:56];
    53: reg_0267 <= imem04_in[27:24];
    55: reg_0267 <= imem06_in[59:56];
    57: reg_0267 <= imem06_in[59:56];
    endcase
  end

  // REG#268の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0268 <= imem05_in[7:4];
    13: reg_0268 <= imem05_in[7:4];
    15: reg_0268 <= imem07_in[15:12];
    17: reg_0268 <= imem04_in[39:36];
    19: reg_0268 <= imem04_in[39:36];
    42: reg_0268 <= imem00_in[119:116];
    44: reg_0268 <= imem05_in[7:4];
    46: reg_0268 <= imem04_in[39:36];
    48: reg_0268 <= imem07_in[15:12];
    50: reg_0268 <= imem04_in[39:36];
    52: reg_0268 <= imem05_in[7:4];
    54: reg_0268 <= imem05_in[7:4];
    56: reg_0268 <= imem07_in[15:12];
    58: reg_0268 <= imem04_in[39:36];
    60: reg_0268 <= imem00_in[119:116];
    62: reg_0268 <= imem00_in[119:116];
    64: reg_0268 <= imem07_in[15:12];
    66: reg_0268 <= imem00_in[119:116];
    68: reg_0268 <= imem07_in[15:12];
    70: reg_0268 <= imem05_in[7:4];
    72: reg_0268 <= imem07_in[47:44];
    74: reg_0268 <= imem04_in[39:36];
    76: reg_0268 <= imem07_in[47:44];
    78: reg_0268 <= imem00_in[119:116];
    80: reg_0268 <= imem07_in[47:44];
    82: reg_0268 <= imem04_in[39:36];
    85: reg_0268 <= imem00_in[119:116];
    87: reg_0268 <= imem05_in[7:4];
    endcase
  end

  // REG#269の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0269 <= imem05_in[87:84];
    13: reg_0269 <= imem05_in[87:84];
    15: reg_0269 <= imem05_in[87:84];
    17: reg_0269 <= imem05_in[111:108];
    19: reg_0269 <= imem05_in[111:108];
    22: reg_0269 <= imem05_in[111:108];
    24: reg_0269 <= imem05_in[87:84];
    26: reg_0269 <= imem04_in[59:56];
    28: reg_0269 <= imem05_in[87:84];
    30: reg_0269 <= imem07_in[75:72];
    32: reg_0269 <= imem04_in[59:56];
    34: reg_0269 <= imem05_in[87:84];
    36: reg_0269 <= imem05_in[111:108];
    38: reg_0269 <= imem04_in[59:56];
    40: reg_0269 <= imem05_in[87:84];
    42: reg_0269 <= imem01_in[51:48];
    44: reg_0269 <= imem01_in[51:48];
    46: reg_0269 <= imem04_in[59:56];
    50: reg_0269 <= imem05_in[111:108];
    56: reg_0269 <= imem05_in[87:84];
    62: reg_0269 <= imem05_in[87:84];
    64: reg_0269 <= imem05_in[87:84];
    67: reg_0269 <= imem05_in[87:84];
    69: reg_0269 <= imem05_in[87:84];
    71: reg_0269 <= imem05_in[87:84];
    73: reg_0269 <= imem05_in[111:108];
    endcase
  end

  // REG#270の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0270 <= imem05_in[43:40];
    13: reg_0270 <= imem05_in[43:40];
    15: reg_0270 <= imem05_in[43:40];
    17: reg_0270 <= imem07_in[59:56];
    19: reg_0270 <= imem05_in[43:40];
    22: reg_0270 <= imem07_in[59:56];
    24: reg_0270 <= imem07_in[59:56];
    26: reg_0270 <= imem04_in[71:68];
    28: reg_0270 <= imem07_in[59:56];
    30: reg_0270 <= imem00_in[7:4];
    32: reg_0270 <= imem00_in[7:4];
    34: reg_0270 <= imem05_in[43:40];
    36: reg_0270 <= imem07_in[59:56];
    38: reg_0270 <= imem04_in[71:68];
    40: reg_0270 <= imem04_in[71:68];
    42: reg_0270 <= imem07_in[59:56];
    45: reg_0270 <= imem01_in[35:32];
    47: reg_0270 <= imem00_in[7:4];
    49: reg_0270 <= imem05_in[43:40];
    51: reg_0270 <= imem04_in[71:68];
    53: reg_0270 <= imem06_in[47:44];
    55: reg_0270 <= imem05_in[43:40];
    58: reg_0270 <= imem01_in[35:32];
    60: reg_0270 <= imem05_in[43:40];
    63: reg_0270 <= imem04_in[71:68];
    65: reg_0270 <= imem06_in[47:44];
    67: reg_0270 <= imem04_in[71:68];
    69: reg_0270 <= imem00_in[7:4];
    71: reg_0270 <= imem06_in[47:44];
    90: reg_0270 <= imem04_in[71:68];
    92: reg_0270 <= imem01_in[35:32];
    endcase
  end

  // REG#271の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0271 <= imem05_in[23:20];
    13: reg_0271 <= imem01_in[15:12];
    15: reg_0271 <= imem01_in[43:40];
    17: reg_0271 <= imem05_in[23:20];
    19: reg_0271 <= imem01_in[15:12];
    21: reg_0271 <= imem01_in[43:40];
    23: reg_0271 <= imem01_in[15:12];
    25: reg_0271 <= imem05_in[23:20];
    27: reg_0271 <= imem05_in[23:20];
    29: reg_0271 <= imem01_in[15:12];
    31: reg_0271 <= imem01_in[15:12];
    33: reg_0271 <= imem01_in[43:40];
    35: reg_0271 <= imem01_in[15:12];
    37: reg_0271 <= imem00_in[3:0];
    39: reg_0271 <= imem01_in[43:40];
    42: reg_0271 <= imem01_in[43:40];
    44: reg_0271 <= imem01_in[43:40];
    46: reg_0271 <= imem03_in[115:112];
    48: reg_0271 <= imem03_in[115:112];
    50: reg_0271 <= imem01_in[35:32];
    52: reg_0271 <= imem05_in[23:20];
    54: reg_0271 <= imem05_in[23:20];
    56: reg_0271 <= imem01_in[43:40];
    58: reg_0271 <= imem00_in[3:0];
    60: reg_0271 <= imem01_in[43:40];
    62: reg_0271 <= imem05_in[23:20];
    64: reg_0271 <= imem01_in[35:32];
    66: reg_0271 <= imem01_in[35:32];
    68: reg_0271 <= imem00_in[3:0];
    70: reg_0271 <= imem01_in[35:32];
    72: reg_0271 <= imem01_in[119:116];
    74: reg_0271 <= imem00_in[3:0];
    76: reg_0271 <= imem03_in[115:112];
    78: reg_0271 <= imem01_in[35:32];
    80: reg_0271 <= imem05_in[23:20];
    82: reg_0271 <= imem03_in[115:112];
    84: reg_0271 <= imem03_in[115:112];
    86: reg_0271 <= imem01_in[119:116];
    88: reg_0271 <= imem05_in[23:20];
    90: reg_0271 <= imem03_in[115:112];
    endcase
  end

  // REG#272の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0272 <= imem05_in[99:96];
    13: reg_0272 <= imem01_in[55:52];
    15: reg_0272 <= imem01_in[55:52];
    17: reg_0272 <= imem05_in[99:96];
    19: reg_0272 <= imem05_in[99:96];
    22: reg_0272 <= imem01_in[55:52];
    24: reg_0272 <= imem06_in[127:124];
    26: reg_0272 <= imem06_in[127:124];
    28: reg_0272 <= imem06_in[127:124];
    30: reg_0272 <= imem02_in[127:124];
    32: reg_0272 <= imem02_in[127:124];
    34: reg_0272 <= imem01_in[103:100];
    36: reg_0272 <= imem02_in[127:124];
    38: reg_0272 <= imem02_in[127:124];
    40: reg_0272 <= imem02_in[127:124];
    42: reg_0272 <= imem02_in[127:124];
    44: reg_0272 <= imem02_in[127:124];
    47: reg_0272 <= imem01_in[55:52];
    51: reg_0272 <= imem07_in[7:4];
    53: reg_0272 <= imem06_in[123:120];
    55: reg_0272 <= imem06_in[123:120];
    57: reg_0272 <= imem02_in[127:124];
    59: reg_0272 <= imem01_in[55:52];
    61: reg_0272 <= imem05_in[99:96];
    65: reg_0272 <= imem05_in[99:96];
    67: reg_0272 <= imem02_in[127:124];
    69: reg_0272 <= imem05_in[99:96];
    71: reg_0272 <= imem02_in[99:96];
    73: reg_0272 <= imem01_in[103:100];
    75: reg_0272 <= imem02_in[127:124];
    77: reg_0272 <= imem02_in[127:124];
    79: reg_0272 <= imem01_in[103:100];
    81: reg_0272 <= imem06_in[127:124];
    83: reg_0272 <= imem02_in[127:124];
    85: reg_0272 <= imem07_in[7:4];
    87: reg_0272 <= imem05_in[99:96];
    endcase
  end

  // REG#273の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0273 <= imem05_in[31:28];
    13: reg_0273 <= imem01_in[87:84];
    15: reg_0273 <= imem01_in[51:48];
    17: reg_0273 <= imem01_in[51:48];
    19: reg_0273 <= imem00_in[127:124];
    21: reg_0273 <= imem05_in[31:28];
    23: reg_0273 <= imem05_in[31:28];
    25: reg_0273 <= imem03_in[51:48];
    27: reg_0273 <= imem00_in[127:124];
    29: reg_0273 <= imem03_in[51:48];
    31: reg_0273 <= imem01_in[87:84];
    33: reg_0273 <= imem03_in[51:48];
    35: reg_0273 <= imem01_in[87:84];
    37: reg_0273 <= imem05_in[31:28];
    39: reg_0273 <= imem05_in[31:28];
    41: reg_0273 <= imem03_in[51:48];
    43: reg_0273 <= imem01_in[51:48];
    45: reg_0273 <= imem03_in[51:48];
    47: reg_0273 <= imem05_in[31:28];
    49: reg_0273 <= imem05_in[31:28];
    51: reg_0273 <= imem00_in[127:124];
    53: reg_0273 <= imem01_in[51:48];
    endcase
  end

  // REG#274の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0274 <= imem05_in[55:52];
    13: reg_0274 <= imem01_in[91:88];
    15: reg_0274 <= imem01_in[91:88];
    17: reg_0274 <= imem05_in[55:52];
    19: reg_0274 <= imem05_in[55:52];
    21: reg_0274 <= imem05_in[55:52];
    23: reg_0274 <= imem05_in[55:52];
    25: reg_0274 <= imem01_in[91:88];
    49: reg_0274 <= imem01_in[91:88];
    64: reg_0274 <= imem01_in[91:88];
    66: reg_0274 <= imem05_in[55:52];
    80: reg_0274 <= imem05_in[55:52];
    82: reg_0274 <= imem00_in[7:4];
    84: reg_0274 <= imem01_in[91:88];
    86: reg_0274 <= imem00_in[7:4];
    88: reg_0274 <= imem00_in[7:4];
    90: reg_0274 <= imem05_in[55:52];
    92: reg_0274 <= imem04_in[55:52];
    94: reg_0274 <= imem05_in[55:52];
    96: reg_0274 <= imem05_in[55:52];
    endcase
  end

  // REG#275の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0275 <= imem04_in[111:108];
    14: reg_0275 <= imem05_in[79:76];
    16: reg_0275 <= imem00_in[79:76];
    18: reg_0275 <= imem00_in[79:76];
    20: reg_0275 <= imem05_in[79:76];
    51: reg_0275 <= imem07_in[99:96];
    53: reg_0275 <= imem07_in[99:96];
    55: reg_0275 <= imem04_in[111:108];
    57: reg_0275 <= imem05_in[79:76];
    59: reg_0275 <= imem02_in[43:40];
    61: reg_0275 <= imem02_in[43:40];
    63: reg_0275 <= imem00_in[79:76];
    65: reg_0275 <= imem02_in[43:40];
    67: reg_0275 <= imem07_in[99:96];
    69: reg_0275 <= imem07_in[99:96];
    71: reg_0275 <= imem07_in[99:96];
    73: reg_0275 <= imem05_in[79:76];
    endcase
  end

  // REG#276の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0276 <= imem04_in[71:68];
    15: reg_0276 <= imem04_in[71:68];
    17: reg_0276 <= imem01_in[87:84];
    19: reg_0276 <= imem04_in[71:68];
    39: reg_0276 <= imem01_in[87:84];
    42: reg_0276 <= imem04_in[71:68];
    92: reg_0276 <= imem01_in[87:84];
    endcase
  end

  // REG#277の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0277 <= imem04_in[47:44];
    15: reg_0277 <= imem04_in[47:44];
    17: reg_0277 <= imem04_in[47:44];
    21: reg_0277 <= imem04_in[47:44];
    24: reg_0277 <= imem04_in[47:44];
    84: reg_0277 <= imem02_in[55:52];
    97: reg_0277 <= imem04_in[47:44];
    endcase
  end

  // REG#278の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0278 <= imem04_in[127:124];
    15: reg_0278 <= imem01_in[71:68];
    17: reg_0278 <= imem01_in[71:68];
    19: reg_0278 <= imem04_in[127:124];
    40: reg_0278 <= imem05_in[55:52];
    42: reg_0278 <= imem05_in[55:52];
    44: reg_0278 <= imem03_in[11:8];
    46: reg_0278 <= imem04_in[51:48];
    48: reg_0278 <= imem01_in[71:68];
    50: reg_0278 <= imem04_in[127:124];
    52: reg_0278 <= imem03_in[11:8];
    54: reg_0278 <= imem04_in[51:48];
    56: reg_0278 <= imem03_in[11:8];
    58: reg_0278 <= imem03_in[11:8];
    60: reg_0278 <= imem03_in[11:8];
    62: reg_0278 <= imem04_in[51:48];
    64: reg_0278 <= imem04_in[127:124];
    66: reg_0278 <= imem02_in[127:124];
    68: reg_0278 <= imem03_in[11:8];
    70: reg_0278 <= imem03_in[11:8];
    endcase
  end

  // REG#279の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0279 <= imem04_in[31:28];
    16: reg_0279 <= imem00_in[127:124];
    18: reg_0279 <= imem04_in[31:28];
    44: reg_0279 <= imem00_in[127:124];
    46: reg_0279 <= imem04_in[31:28];
    50: reg_0279 <= imem02_in[7:4];
    52: reg_0279 <= imem02_in[7:4];
    endcase
  end

  // REG#280の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0280 <= op1_01_out;
    15: reg_0280 <= op1_01_out;
    17: reg_0280 <= op1_01_out;
    19: reg_0280 <= op1_01_out;
    21: reg_0280 <= op1_01_out;
    23: reg_0280 <= op1_01_out;
    25: reg_0280 <= op1_01_out;
    27: reg_0280 <= op1_01_out;
    29: reg_0280 <= op1_01_out;
    31: reg_0280 <= op1_01_out;
    33: reg_0280 <= op1_01_out;
    35: reg_0280 <= op1_01_out;
    37: reg_0280 <= op1_01_out;
    39: reg_0280 <= op1_01_out;
    41: reg_0280 <= op1_01_out;
    43: reg_0280 <= op1_01_out;
    45: reg_0280 <= op1_01_out;
    47: reg_0280 <= op1_01_out;
    49: reg_0280 <= op1_01_out;
    51: reg_0280 <= op1_01_out;
    53: reg_0280 <= op1_01_out;
    55: reg_0280 <= op1_01_out;
    57: reg_0280 <= op1_01_out;
    59: reg_0280 <= op1_01_out;
    61: reg_0280 <= op1_01_out;
    63: reg_0280 <= op1_01_out;
    65: reg_0280 <= op1_01_out;
    67: reg_0280 <= op1_01_out;
    69: reg_0280 <= op1_01_out;
    71: reg_0280 <= op1_01_out;
    73: reg_0280 <= op1_01_out;
    75: reg_0280 <= op1_01_out;
    77: reg_0280 <= op1_01_out;
    79: reg_0280 <= op1_01_out;
    81: reg_0280 <= op1_01_out;
    83: reg_0280 <= op1_01_out;
    85: reg_0280 <= op1_01_out;
    87: reg_0280 <= op1_01_out;
    89: reg_0280 <= op1_01_out;
    91: reg_0280 <= op1_01_out;
    93: reg_0280 <= op1_01_out;
    95: reg_0280 <= op1_01_out;
    97: reg_0280 <= op1_01_out;
    endcase
  end

  // REG#281の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0281 <= imem04_in[15:12];
    17: reg_0281 <= imem04_in[15:12];
    20: reg_0281 <= imem04_in[15:12];
    22: reg_0281 <= imem04_in[15:12];
    25: reg_0281 <= imem04_in[15:12];
    27: reg_0281 <= imem04_in[15:12];
    29: reg_0281 <= imem00_in[103:100];
    31: reg_0281 <= imem04_in[15:12];
    33: reg_0281 <= imem04_in[15:12];
    35: reg_0281 <= imem04_in[15:12];
    37: reg_0281 <= imem02_in[119:116];
    39: reg_0281 <= imem03_in[31:28];
    41: reg_0281 <= imem05_in[55:52];
    43: reg_0281 <= imem02_in[119:116];
    45: reg_0281 <= imem00_in[103:100];
    47: reg_0281 <= imem04_in[15:12];
    49: reg_0281 <= imem04_in[15:12];
    58: reg_0281 <= imem00_in[103:100];
    60: reg_0281 <= imem02_in[119:116];
    62: reg_0281 <= imem02_in[119:116];
    65: reg_0281 <= imem00_in[103:100];
    67: reg_0281 <= imem05_in[55:52];
    70: reg_0281 <= imem03_in[31:28];
    97: reg_0281 <= imem02_in[119:116];
    endcase
  end

  // REG#282の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0282 <= imem04_in[51:48];
    17: reg_0282 <= imem04_in[51:48];
    21: reg_0282 <= imem04_in[51:48];
    24: reg_0282 <= imem04_in[51:48];
    84: reg_0282 <= imem04_in[51:48];
    86: reg_0282 <= imem04_in[51:48];
    88: reg_0282 <= imem04_in[51:48];
    90: reg_0282 <= imem04_in[51:48];
    92: reg_0282 <= imem01_in[59:56];
    94: reg_0282 <= imem04_in[51:48];
    endcase
  end

  // REG#283の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0283 <= imem04_in[23:20];
    18: reg_0283 <= imem04_in[23:20];
    47: reg_0283 <= imem04_in[23:20];
    49: reg_0283 <= imem02_in[71:68];
    51: reg_0283 <= imem01_in[43:40];
    53: reg_0283 <= imem01_in[43:40];
    endcase
  end

  // REG#284の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0284 <= imem04_in[123:120];
    18: reg_0284 <= imem07_in[23:20];
    20: reg_0284 <= imem07_in[23:20];
    22: reg_0284 <= imem00_in[115:112];
    24: reg_0284 <= imem07_in[23:20];
    26: reg_0284 <= imem07_in[23:20];
    28: reg_0284 <= imem07_in[23:20];
    30: reg_0284 <= imem04_in[123:120];
    32: reg_0284 <= imem00_in[115:112];
    34: reg_0284 <= imem07_in[23:20];
    36: reg_0284 <= imem06_in[71:68];
    38: reg_0284 <= imem07_in[23:20];
    40: reg_0284 <= imem07_in[23:20];
    42: reg_0284 <= imem04_in[123:120];
    endcase
  end

  // REG#285の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0285 <= imem04_in[83:80];
    18: reg_0285 <= imem04_in[83:80];
    45: reg_0285 <= imem01_in[115:112];
    47: reg_0285 <= imem04_in[83:80];
    49: reg_0285 <= imem01_in[115:112];
    69: reg_0285 <= imem04_in[83:80];
    71: reg_0285 <= imem01_in[115:112];
    73: reg_0285 <= imem04_in[83:80];
    75: reg_0285 <= imem07_in[75:72];
    77: reg_0285 <= imem04_in[83:80];
    79: reg_0285 <= imem01_in[115:112];
    82: reg_0285 <= imem04_in[83:80];
    84: reg_0285 <= imem02_in[23:20];
    97: reg_0285 <= imem01_in[115:112];
    endcase
  end

  // REG#286の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0286 <= imem04_in[103:100];
    18: reg_0286 <= imem04_in[103:100];
    44: reg_0286 <= imem03_in[75:72];
    46: reg_0286 <= imem04_in[103:100];
    50: reg_0286 <= imem02_in[27:24];
    52: reg_0286 <= imem03_in[75:72];
    54: reg_0286 <= imem01_in[127:124];
    56: reg_0286 <= imem03_in[95:92];
    58: reg_0286 <= imem02_in[27:24];
    60: reg_0286 <= imem02_in[27:24];
    62: reg_0286 <= imem04_in[103:100];
    64: reg_0286 <= imem02_in[27:24];
    66: reg_0286 <= imem02_in[27:24];
    68: reg_0286 <= imem03_in[95:92];
    70: reg_0286 <= imem02_in[27:24];
    72: reg_0286 <= imem04_in[103:100];
    74: reg_0286 <= imem03_in[95:92];
    76: reg_0286 <= imem03_in[95:92];
    78: reg_0286 <= imem03_in[95:92];
    80: reg_0286 <= imem05_in[43:40];
    82: reg_0286 <= imem03_in[75:72];
    84: reg_0286 <= imem03_in[75:72];
    86: reg_0286 <= imem04_in[103:100];
    88: reg_0286 <= imem01_in[127:124];
    90: reg_0286 <= imem03_in[75:72];
    endcase
  end

  // REG#287の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0287 <= op1_02_out;
    17: reg_0287 <= op1_02_out;
    19: reg_0287 <= op1_02_out;
    21: reg_0287 <= op1_02_out;
    23: reg_0287 <= op1_02_out;
    25: reg_0287 <= op1_02_out;
    27: reg_0287 <= op1_02_out;
    29: reg_0287 <= op1_02_out;
    31: reg_0287 <= op1_02_out;
    33: reg_0287 <= op1_02_out;
    35: reg_0287 <= op1_02_out;
    37: reg_0287 <= op1_02_out;
    39: reg_0287 <= op1_02_out;
    41: reg_0287 <= op1_02_out;
    43: reg_0287 <= op1_02_out;
    45: reg_0287 <= op1_02_out;
    47: reg_0287 <= op1_02_out;
    49: reg_0287 <= op1_02_out;
    51: reg_0287 <= op1_02_out;
    53: reg_0287 <= op1_02_out;
    55: reg_0287 <= op1_02_out;
    57: reg_0287 <= op1_02_out;
    59: reg_0287 <= op1_02_out;
    61: reg_0287 <= op1_02_out;
    63: reg_0287 <= op1_02_out;
    65: reg_0287 <= op1_02_out;
    67: reg_0287 <= op1_02_out;
    69: reg_0287 <= op1_02_out;
    71: reg_0287 <= op1_02_out;
    73: reg_0287 <= op1_02_out;
    75: reg_0287 <= op1_02_out;
    77: reg_0287 <= op1_02_out;
    79: reg_0287 <= op1_02_out;
    81: reg_0287 <= op1_02_out;
    83: reg_0287 <= op1_02_out;
    85: reg_0287 <= op1_02_out;
    87: reg_0287 <= op1_02_out;
    89: reg_0287 <= op1_02_out;
    91: reg_0287 <= op1_02_out;
    93: reg_0287 <= op1_02_out;
    95: reg_0287 <= op1_02_out;
    97: reg_0287 <= op1_02_out;
    endcase
  end

  // REG#288の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0288 <= imem04_in[115:112];
    19: reg_0288 <= imem01_in[7:4];
    21: reg_0288 <= imem04_in[115:112];
    23: reg_0288 <= imem04_in[115:112];
    26: reg_0288 <= imem05_in[19:16];
    28: reg_0288 <= imem05_in[19:16];
    30: reg_0288 <= imem06_in[59:56];
    32: reg_0288 <= imem01_in[7:4];
    34: reg_0288 <= imem04_in[115:112];
    36: reg_0288 <= imem07_in[87:84];
    38: reg_0288 <= imem05_in[19:16];
    40: reg_0288 <= imem07_in[87:84];
    42: reg_0288 <= imem04_in[115:112];
    96: reg_0288 <= imem06_in[59:56];
    endcase
  end

  // REG#289の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0289 <= imem04_in[55:52];
    19: reg_0289 <= imem01_in[23:20];
    21: reg_0289 <= imem01_in[23:20];
    23: reg_0289 <= imem04_in[55:52];
    26: reg_0289 <= imem05_in[119:116];
    28: reg_0289 <= imem07_in[47:44];
    30: reg_0289 <= imem04_in[55:52];
    32: reg_0289 <= imem05_in[119:116];
    34: reg_0289 <= imem07_in[47:44];
    36: reg_0289 <= imem05_in[119:116];
    38: reg_0289 <= imem04_in[55:52];
    40: reg_0289 <= imem06_in[11:8];
    42: reg_0289 <= imem07_in[47:44];
    45: reg_0289 <= imem07_in[47:44];
    47: reg_0289 <= imem04_in[55:52];
    49: reg_0289 <= imem06_in[11:8];
    51: reg_0289 <= imem05_in[119:116];
    53: reg_0289 <= imem06_in[11:8];
    55: reg_0289 <= imem07_in[47:44];
    57: reg_0289 <= imem01_in[43:40];
    59: reg_0289 <= imem05_in[119:116];
    61: reg_0289 <= imem01_in[43:40];
    63: reg_0289 <= imem06_in[3:0];
    65: reg_0289 <= imem07_in[47:44];
    67: reg_0289 <= imem04_in[55:52];
    69: reg_0289 <= imem04_in[55:52];
    71: reg_0289 <= imem06_in[11:8];
    87: reg_0289 <= imem06_in[3:0];
    89: reg_0289 <= imem06_in[11:8];
    endcase
  end

  // REG#290の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0290 <= imem04_in[75:72];
    19: reg_0290 <= imem02_in[51:48];
    21: reg_0290 <= imem04_in[75:72];
    23: reg_0290 <= imem04_in[75:72];
    26: reg_0290 <= imem02_in[51:48];
    51: reg_0290 <= imem02_in[51:48];
    53: reg_0290 <= imem02_in[51:48];
    55: reg_0290 <= imem04_in[75:72];
    57: reg_0290 <= imem04_in[75:72];
    59: reg_0290 <= imem03_in[43:40];
    61: reg_0290 <= imem02_in[51:48];
    63: reg_0290 <= imem02_in[51:48];
    71: reg_0290 <= imem04_in[39:36];
    73: reg_0290 <= imem04_in[75:72];
    75: reg_0290 <= imem07_in[83:80];
    77: reg_0290 <= imem07_in[83:80];
    79: reg_0290 <= imem03_in[43:40];
    81: reg_0290 <= imem02_in[51:48];
    83: reg_0290 <= imem02_in[51:48];
    86: reg_0290 <= imem04_in[75:72];
    88: reg_0290 <= imem02_in[51:48];
    90: reg_0290 <= imem03_in[43:40];
    95: reg_0290 <= imem07_in[83:80];
    endcase
  end

  // REG#291の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0291 <= imem04_in[79:76];
    19: reg_0291 <= imem02_in[103:100];
    21: reg_0291 <= imem02_in[103:100];
    86: reg_0291 <= imem02_in[27:24];
    88: reg_0291 <= imem05_in[123:120];
    90: reg_0291 <= imem05_in[123:120];
    92: reg_0291 <= imem01_in[63:60];
    94: reg_0291 <= imem01_in[63:60];
    96: reg_0291 <= imem02_in[27:24];
    endcase
  end

  // REG#292の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0292 <= imem04_in[95:92];
    19: reg_0292 <= imem03_in[91:88];
    21: reg_0292 <= imem04_in[87:84];
    24: reg_0292 <= imem04_in[87:84];
    81: reg_0292 <= imem04_in[95:92];
    83: reg_0292 <= imem04_in[87:84];
    endcase
  end

  // REG#293の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0293 <= imem04_in[67:64];
    19: reg_0293 <= imem06_in[7:4];
    21: reg_0293 <= imem04_in[67:64];
    23: reg_0293 <= imem06_in[7:4];
    25: reg_0293 <= imem04_in[67:64];
    27: reg_0293 <= imem06_in[7:4];
    29: reg_0293 <= imem06_in[7:4];
    59: reg_0293 <= imem06_in[7:4];
    61: reg_0293 <= imem06_in[7:4];
    69: reg_0293 <= imem02_in[75:72];
    71: reg_0293 <= imem06_in[7:4];
    89: reg_0293 <= imem06_in[7:4];
    92: reg_0293 <= imem06_in[7:4];
    94: reg_0293 <= imem04_in[67:64];
    endcase
  end

  // REG#294の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0294 <= imem04_in[43:40];
    19: reg_0294 <= imem06_in[47:44];
    21: reg_0294 <= imem04_in[43:40];
    23: reg_0294 <= imem04_in[15:12];
    25: reg_0294 <= imem06_in[47:44];
    27: reg_0294 <= imem04_in[43:40];
    29: reg_0294 <= imem06_in[47:44];
    55: reg_0294 <= imem06_in[47:44];
    57: reg_0294 <= imem06_in[47:44];
    91: reg_0294 <= imem01_in[111:108];
    93: reg_0294 <= imem01_in[111:108];
    96: reg_0294 <= imem04_in[43:40];
    endcase
  end

  // REG#295の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0295 <= imem04_in[99:96];
    19: reg_0295 <= imem07_in[99:96];
    21: reg_0295 <= imem07_in[99:96];
    23: reg_0295 <= imem05_in[67:64];
    25: reg_0295 <= imem05_in[67:64];
    27: reg_0295 <= imem06_in[75:72];
    29: reg_0295 <= imem06_in[75:72];
    59: reg_0295 <= imem04_in[99:96];
    endcase
  end

  // REG#296の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0296 <= imem04_in[87:84];
    19: reg_0296 <= imem04_in[87:84];
    42: reg_0296 <= imem04_in[87:84];
    endcase
  end

  // REG#297の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0297 <= imem04_in[91:88];
    19: reg_0297 <= imem07_in[119:116];
    21: reg_0297 <= imem04_in[91:88];
    23: reg_0297 <= imem04_in[91:88];
    26: reg_0297 <= imem06_in[23:20];
    28: reg_0297 <= imem04_in[91:88];
    30: reg_0297 <= imem04_in[91:88];
    32: reg_0297 <= imem07_in[79:76];
    34: reg_0297 <= imem04_in[91:88];
    36: reg_0297 <= imem07_in[79:76];
    38: reg_0297 <= imem07_in[79:76];
    40: reg_0297 <= imem07_in[119:116];
    42: reg_0297 <= imem06_in[23:20];
    44: reg_0297 <= imem07_in[79:76];
    46: reg_0297 <= imem06_in[27:24];
    48: reg_0297 <= imem07_in[79:76];
    50: reg_0297 <= imem06_in[27:24];
    52: reg_0297 <= imem07_in[79:76];
    54: reg_0297 <= imem06_in[23:20];
    56: reg_0297 <= imem06_in[27:24];
    58: reg_0297 <= imem06_in[23:20];
    86: reg_0297 <= imem06_in[23:20];
    95: reg_0297 <= imem06_in[27:24];
    endcase
  end

  // REG#298の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0298 <= imem04_in[107:104];
    19: reg_0298 <= imem00_in[115:112];
    21: reg_0298 <= imem00_in[115:112];
    23: reg_0298 <= imem04_in[107:104];
    25: reg_0298 <= imem04_in[107:104];
    27: reg_0298 <= imem00_in[115:112];
    29: reg_0298 <= imem00_in[115:112];
    31: reg_0298 <= imem04_in[107:104];
    33: reg_0298 <= imem04_in[107:104];
    35: reg_0298 <= imem02_in[59:56];
    37: reg_0298 <= imem03_in[99:96];
    39: reg_0298 <= imem02_in[59:56];
    41: reg_0298 <= imem04_in[107:104];
    43: reg_0298 <= imem02_in[59:56];
    45: reg_0298 <= imem03_in[99:96];
    47: reg_0298 <= imem00_in[115:112];
    49: reg_0298 <= imem05_in[99:96];
    51: reg_0298 <= imem04_in[107:104];
    53: reg_0298 <= imem03_in[99:96];
    55: reg_0298 <= imem03_in[99:96];
    88: reg_0298 <= imem05_in[99:96];
    90: reg_0298 <= imem03_in[99:96];
    92: reg_0298 <= imem00_in[115:112];
    95: reg_0298 <= imem05_in[99:96];
    endcase
  end

  // REG#299の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0299 <= imem04_in[39:36];
    19: reg_0299 <= imem01_in[47:44];
    21: reg_0299 <= imem01_in[47:44];
    23: reg_0299 <= imem01_in[47:44];
    25: reg_0299 <= imem01_in[47:44];
    48: reg_0299 <= imem04_in[39:36];
    50: reg_0299 <= imem01_in[47:44];
    52: reg_0299 <= imem07_in[111:108];
    54: reg_0299 <= imem07_in[111:108];
    56: reg_0299 <= imem07_in[111:108];
    58: reg_0299 <= imem07_in[39:36];
    60: reg_0299 <= imem04_in[39:36];
    62: reg_0299 <= imem04_in[39:36];
    64: reg_0299 <= imem04_in[39:36];
    66: reg_0299 <= imem04_in[39:36];
    68: reg_0299 <= imem07_in[111:108];
    70: reg_0299 <= imem07_in[111:108];
    72: reg_0299 <= imem07_in[39:36];
    74: reg_0299 <= imem07_in[39:36];
    77: reg_0299 <= imem07_in[111:108];
    79: reg_0299 <= imem07_in[111:108];
    94: reg_0299 <= imem04_in[39:36];
    96: reg_0299 <= imem04_in[39:36];
    endcase
  end

  // REG#300の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0300 <= imem04_in[35:32];
    19: reg_0300 <= imem02_in[23:20];
    21: reg_0300 <= imem04_in[35:32];
    23: reg_0300 <= imem02_in[23:20];
    25: reg_0300 <= imem02_in[23:20];
    27: reg_0300 <= imem02_in[71:68];
    29: reg_0300 <= imem02_in[99:96];
    31: reg_0300 <= imem02_in[71:68];
    33: reg_0300 <= imem02_in[23:20];
    35: reg_0300 <= imem02_in[99:96];
    37: reg_0300 <= imem02_in[23:20];
    39: reg_0300 <= imem02_in[71:68];
    41: reg_0300 <= imem02_in[71:68];
    43: reg_0300 <= imem02_in[23:20];
    45: reg_0300 <= imem02_in[99:96];
    64: reg_0300 <= imem02_in[23:20];
    66: reg_0300 <= imem02_in[99:96];
    68: reg_0300 <= imem02_in[23:20];
    70: reg_0300 <= imem02_in[99:96];
    72: reg_0300 <= imem04_in[35:32];
    74: reg_0300 <= imem02_in[99:96];
    76: reg_0300 <= imem04_in[35:32];
    78: reg_0300 <= imem04_in[35:32];
    80: reg_0300 <= imem02_in[99:96];
    82: reg_0300 <= imem04_in[35:32];
    85: reg_0300 <= imem04_in[35:32];
    87: reg_0300 <= imem02_in[35:32];
    89: reg_0300 <= imem02_in[35:32];
    91: reg_0300 <= imem02_in[99:96];
    93: reg_0300 <= imem04_in[35:32];
    95: reg_0300 <= imem02_in[71:68];
    endcase
  end

  // REG#301の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0301 <= imem04_in[19:16];
    20: reg_0301 <= imem04_in[19:16];
    22: reg_0301 <= imem04_in[19:16];
    24: reg_0301 <= imem04_in[19:16];
    84: reg_0301 <= imem04_in[19:16];
    86: reg_0301 <= imem03_in[87:84];
    88: reg_0301 <= imem03_in[87:84];
    endcase
  end

  // REG#302の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0302 <= imem04_in[63:60];
    20: reg_0302 <= imem03_in[55:52];
    22: reg_0302 <= imem04_in[63:60];
    25: reg_0302 <= imem03_in[59:56];
    27: reg_0302 <= imem03_in[59:56];
    30: reg_0302 <= imem04_in[63:60];
    32: reg_0302 <= imem04_in[63:60];
    34: reg_0302 <= imem03_in[59:56];
    36: reg_0302 <= imem03_in[59:56];
    38: reg_0302 <= imem03_in[59:56];
    40: reg_0302 <= imem03_in[59:56];
    42: reg_0302 <= imem04_in[63:60];
    96: reg_0302 <= imem04_in[63:60];
    endcase
  end

  // REG#303の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0303 <= imem04_in[3:0];
    20: reg_0303 <= imem04_in[3:0];
    22: reg_0303 <= imem04_in[3:0];
    25: reg_0303 <= imem04_in[3:0];
    27: reg_0303 <= imem04_in[3:0];
    29: reg_0303 <= imem03_in[39:36];
    31: reg_0303 <= imem04_in[3:0];
    33: reg_0303 <= imem03_in[39:36];
    35: reg_0303 <= imem03_in[39:36];
    37: reg_0303 <= imem07_in[19:16];
    39: reg_0303 <= imem03_in[39:36];
    41: reg_0303 <= imem04_in[3:0];
    43: reg_0303 <= imem07_in[19:16];
    endcase
  end

  // REG#304の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0304 <= imem04_in[11:8];
    20: reg_0304 <= imem06_in[63:60];
    22: reg_0304 <= imem01_in[115:112];
    24: reg_0304 <= imem01_in[115:112];
    27: reg_0304 <= imem04_in[79:76];
    29: reg_0304 <= imem04_in[79:76];
    31: reg_0304 <= imem06_in[63:60];
    33: reg_0304 <= imem04_in[11:8];
    35: reg_0304 <= imem04_in[79:76];
    37: reg_0304 <= imem01_in[115:112];
    39: reg_0304 <= imem04_in[11:8];
    41: reg_0304 <= imem01_in[115:112];
    92: reg_0304 <= imem01_in[115:112];
    endcase
  end

  // REG#305の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0305 <= imem04_in[27:24];
    20: reg_0305 <= imem04_in[27:24];
    22: reg_0305 <= imem04_in[27:24];
    25: reg_0305 <= imem07_in[63:60];
    27: reg_0305 <= imem04_in[27:24];
    29: reg_0305 <= imem07_in[63:60];
    31: reg_0305 <= imem07_in[63:60];
    33: reg_0305 <= imem07_in[63:60];
    35: reg_0305 <= imem07_in[63:60];
    37: reg_0305 <= imem07_in[63:60];
    39: reg_0305 <= imem04_in[27:24];
    41: reg_0305 <= imem04_in[27:24];
    44: reg_0305 <= imem07_in[63:60];
    46: reg_0305 <= imem07_in[63:60];
    48: reg_0305 <= imem07_in[31:28];
    50: reg_0305 <= imem07_in[63:60];
    52: reg_0305 <= imem07_in[63:60];
    54: reg_0305 <= imem02_in[47:44];
    56: reg_0305 <= imem04_in[15:12];
    58: reg_0305 <= imem07_in[63:60];
    60: reg_0305 <= imem02_in[47:44];
    62: reg_0305 <= imem02_in[47:44];
    64: reg_0305 <= imem07_in[31:28];
    66: reg_0305 <= imem07_in[31:28];
    68: reg_0305 <= imem07_in[31:28];
    70: reg_0305 <= imem07_in[31:28];
    72: reg_0305 <= imem04_in[15:12];
    74: reg_0305 <= imem04_in[15:12];
    76: reg_0305 <= imem03_in[7:4];
    78: reg_0305 <= imem04_in[7:4];
    80: reg_0305 <= imem04_in[27:24];
    82: reg_0305 <= imem04_in[15:12];
    84: reg_0305 <= imem02_in[47:44];
    endcase
  end

  // REG#306の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0306 <= imem04_in[59:56];
    20: reg_0306 <= imem00_in[39:36];
    22: reg_0306 <= imem04_in[59:56];
    24: reg_0306 <= imem04_in[59:56];
    83: reg_0306 <= imem04_in[59:56];
    97: reg_0306 <= imem00_in[39:36];
    endcase
  end

  // REG#307の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0307 <= imem04_in[119:116];
    20: reg_0307 <= imem01_in[27:24];
    22: reg_0307 <= imem04_in[119:116];
    24: reg_0307 <= imem01_in[27:24];
    27: reg_0307 <= imem04_in[119:116];
    29: reg_0307 <= imem03_in[63:60];
    31: reg_0307 <= imem01_in[27:24];
    33: reg_0307 <= imem04_in[119:116];
    35: reg_0307 <= imem04_in[119:116];
    37: reg_0307 <= imem07_in[119:116];
    39: reg_0307 <= imem03_in[63:60];
    41: reg_0307 <= imem04_in[119:116];
    44: reg_0307 <= imem01_in[27:24];
    46: reg_0307 <= imem03_in[63:60];
    48: reg_0307 <= imem01_in[27:24];
    50: reg_0307 <= imem04_in[119:116];
    52: reg_0307 <= imem01_in[27:24];
    55: reg_0307 <= imem03_in[63:60];
    88: reg_0307 <= imem03_in[63:60];
    96: reg_0307 <= imem03_in[63:60];
    endcase
  end

  // REG#308の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0308 <= imem04_in[7:4];
    20: reg_0308 <= imem01_in[107:104];
    22: reg_0308 <= imem01_in[107:104];
    24: reg_0308 <= imem01_in[107:104];
    26: reg_0308 <= imem04_in[7:4];
    28: reg_0308 <= imem04_in[7:4];
    30: reg_0308 <= imem07_in[19:16];
    32: reg_0308 <= imem01_in[107:104];
    34: reg_0308 <= imem04_in[7:4];
    36: reg_0308 <= imem07_in[19:16];
    38: reg_0308 <= imem00_in[67:64];
    40: reg_0308 <= imem04_in[7:4];
    42: reg_0308 <= imem01_in[107:104];
    44: reg_0308 <= imem07_in[19:16];
    46: reg_0308 <= imem04_in[7:4];
    50: reg_0308 <= imem02_in[99:96];
    52: reg_0308 <= imem07_in[19:16];
    54: reg_0308 <= imem04_in[7:4];
    56: reg_0308 <= imem01_in[107:104];
    58: reg_0308 <= imem00_in[67:64];
    60: reg_0308 <= imem04_in[7:4];
    62: reg_0308 <= imem04_in[7:4];
    64: reg_0308 <= imem04_in[7:4];
    66: reg_0308 <= imem04_in[7:4];
    68: reg_0308 <= imem04_in[7:4];
    70: reg_0308 <= imem04_in[7:4];
    72: reg_0308 <= imem04_in[7:4];
    74: reg_0308 <= imem07_in[19:16];
    77: reg_0308 <= imem00_in[67:64];
    79: reg_0308 <= imem02_in[99:96];
    81: reg_0308 <= imem01_in[107:104];
    83: reg_0308 <= imem02_in[99:96];
    87: reg_0308 <= imem01_in[107:104];
    90: reg_0308 <= imem07_in[19:16];
    92: reg_0308 <= imem02_in[99:96];
    94: reg_0308 <= imem04_in[7:4];
    96: reg_0308 <= imem04_in[7:4];
    endcase
  end

  // REG#309の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0309 <= imem03_in[115:112];
    20: reg_0309 <= imem04_in[43:40];
    22: reg_0309 <= imem04_in[43:40];
    25: reg_0309 <= imem03_in[115:112];
    27: reg_0309 <= imem03_in[115:112];
    29: reg_0309 <= imem04_in[47:44];
    31: reg_0309 <= imem06_in[35:32];
    33: reg_0309 <= imem04_in[47:44];
    35: reg_0309 <= imem04_in[43:40];
    37: reg_0309 <= imem06_in[35:32];
    50: reg_0309 <= imem06_in[35:32];
    52: reg_0309 <= imem04_in[11:8];
    54: reg_0309 <= imem04_in[47:44];
    56: reg_0309 <= imem06_in[35:32];
    58: reg_0309 <= imem04_in[11:8];
    60: reg_0309 <= imem04_in[11:8];
    62: reg_0309 <= imem03_in[127:124];
    64: reg_0309 <= imem04_in[11:8];
    66: reg_0309 <= imem04_in[11:8];
    68: reg_0309 <= imem03_in[127:124];
    70: reg_0309 <= imem04_in[11:8];
    72: reg_0309 <= imem04_in[43:40];
    74: reg_0309 <= imem01_in[7:4];
    76: reg_0309 <= imem04_in[11:8];
    78: reg_0309 <= imem04_in[11:8];
    80: reg_0309 <= imem06_in[35:32];
    82: reg_0309 <= imem04_in[11:8];
    85: reg_0309 <= imem03_in[115:112];
    87: reg_0309 <= imem04_in[11:8];
    89: reg_0309 <= imem03_in[127:124];
    91: reg_0309 <= imem06_in[35:32];
    93: reg_0309 <= imem03_in[119:116];
    95: reg_0309 <= imem04_in[47:44];
    97: reg_0309 <= imem04_in[43:40];
    endcase
  end

  // REG#310の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0310 <= imem02_in[87:84];
    21: reg_0310 <= imem02_in[87:84];
    81: reg_0310 <= imem02_in[87:84];
    83: reg_0310 <= imem01_in[99:96];
    85: reg_0310 <= imem01_in[99:96];
    87: reg_0310 <= imem02_in[107:104];
    89: reg_0310 <= imem02_in[87:84];
    91: reg_0310 <= imem00_in[67:64];
    endcase
  end

  // REG#311の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0311 <= imem03_in[35:32];
    22: reg_0311 <= imem03_in[59:56];
    24: reg_0311 <= imem03_in[59:56];
    26: reg_0311 <= imem03_in[35:32];
    28: reg_0311 <= imem03_in[59:56];
    69: reg_0311 <= imem03_in[35:32];
    71: reg_0311 <= imem03_in[35:32];
    73: reg_0311 <= imem06_in[71:68];
    75: reg_0311 <= imem03_in[59:56];
    77: reg_0311 <= imem00_in[7:4];
    79: reg_0311 <= imem00_in[7:4];
    81: reg_0311 <= imem06_in[71:68];
    83: reg_0311 <= imem00_in[7:4];
    85: reg_0311 <= imem03_in[59:56];
    87: reg_0311 <= imem03_in[59:56];
    89: reg_0311 <= imem03_in[35:32];
    92: reg_0311 <= imem03_in[59:56];
    97: reg_0311 <= imem03_in[59:56];
    endcase
  end

  // REG#312の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0312 <= imem03_in[95:92];
    22: reg_0312 <= imem04_in[87:84];
    24: reg_0312 <= imem07_in[87:84];
    26: reg_0312 <= imem03_in[95:92];
    28: reg_0312 <= imem03_in[95:92];
    68: reg_0312 <= imem07_in[87:84];
    70: reg_0312 <= imem03_in[95:92];
    95: reg_0312 <= imem03_in[95:92];
    endcase
  end

  // REG#313の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0313 <= imem06_in[71:68];
    22: reg_0313 <= imem04_in[127:124];
    24: reg_0313 <= imem04_in[127:124];
    82: reg_0313 <= imem04_in[127:124];
    85: reg_0313 <= imem01_in[67:64];
    87: reg_0313 <= imem06_in[71:68];
    89: reg_0313 <= imem04_in[127:124];
    91: reg_0313 <= imem06_in[71:68];
    93: reg_0313 <= imem04_in[127:124];
    95: reg_0313 <= imem04_in[127:124];
    97: reg_0313 <= imem01_in[67:64];
    endcase
  end

  // REG#314の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0314 <= imem02_in[119:116];
    22: reg_0314 <= imem05_in[55:52];
    24: reg_0314 <= imem07_in[95:92];
    26: reg_0314 <= imem05_in[55:52];
    28: reg_0314 <= imem07_in[95:92];
    30: reg_0314 <= imem07_in[31:28];
    32: reg_0314 <= imem05_in[55:52];
    34: reg_0314 <= imem02_in[119:116];
    36: reg_0314 <= imem07_in[31:28];
    38: reg_0314 <= imem02_in[119:116];
    40: reg_0314 <= imem02_in[119:116];
    42: reg_0314 <= imem07_in[31:28];
    44: reg_0314 <= imem02_in[119:116];
    47: reg_0314 <= imem00_in[3:0];
    49: reg_0314 <= imem07_in[95:92];
    51: reg_0314 <= imem02_in[39:36];
    54: reg_0314 <= imem05_in[55:52];
    56: reg_0314 <= imem02_in[119:116];
    58: reg_0314 <= imem02_in[39:36];
    60: reg_0314 <= imem05_in[55:52];
    62: reg_0314 <= imem02_in[39:36];
    65: reg_0314 <= imem05_in[55:52];
    68: reg_0314 <= imem05_in[55:52];
    71: reg_0314 <= imem07_in[31:28];
    73: reg_0314 <= imem07_in[31:28];
    75: reg_0314 <= imem05_in[55:52];
    77: reg_0314 <= imem07_in[95:92];
    79: reg_0314 <= imem05_in[55:52];
    88: reg_0314 <= imem05_in[55:52];
    90: reg_0314 <= imem02_in[39:36];
    92: reg_0314 <= imem02_in[39:36];
    94: reg_0314 <= imem02_in[119:116];
    96: reg_0314 <= imem02_in[39:36];
    endcase
  end

  // REG#315の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0315 <= imem06_in[99:96];
    23: reg_0315 <= imem07_in[59:56];
    25: reg_0315 <= imem07_in[59:56];
    27: reg_0315 <= imem04_in[111:108];
    29: reg_0315 <= imem07_in[59:56];
    31: reg_0315 <= imem04_in[111:108];
    33: reg_0315 <= imem04_in[111:108];
    35: reg_0315 <= imem07_in[59:56];
    37: reg_0315 <= imem07_in[59:56];
    39: reg_0315 <= imem07_in[59:56];
    41: reg_0315 <= imem07_in[59:56];
    43: reg_0315 <= imem07_in[59:56];
    endcase
  end

  // REG#316の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0316 <= op1_03_out;
    22: reg_0316 <= op1_03_out;
    24: reg_0316 <= op1_03_out;
    26: reg_0316 <= op1_03_out;
    28: reg_0316 <= op1_03_out;
    30: reg_0316 <= op1_03_out;
    32: reg_0316 <= op1_03_out;
    34: reg_0316 <= op1_03_out;
    36: reg_0316 <= op1_03_out;
    38: reg_0316 <= op1_03_out;
    40: reg_0316 <= op1_03_out;
    42: reg_0316 <= op1_03_out;
    44: reg_0316 <= op1_03_out;
    46: reg_0316 <= op1_03_out;
    48: reg_0316 <= op1_03_out;
    50: reg_0316 <= op1_03_out;
    52: reg_0316 <= op1_03_out;
    54: reg_0316 <= op1_03_out;
    56: reg_0316 <= op1_03_out;
    58: reg_0316 <= op1_03_out;
    60: reg_0316 <= op1_03_out;
    62: reg_0316 <= op1_03_out;
    64: reg_0316 <= op1_03_out;
    66: reg_0316 <= op1_03_out;
    68: reg_0316 <= op1_03_out;
    70: reg_0316 <= op1_03_out;
    72: reg_0316 <= op1_03_out;
    74: reg_0316 <= op1_03_out;
    76: reg_0316 <= op1_03_out;
    78: reg_0316 <= op1_03_out;
    80: reg_0316 <= op1_03_out;
    82: reg_0316 <= op1_03_out;
    84: reg_0316 <= op1_03_out;
    86: reg_0316 <= op1_03_out;
    88: reg_0316 <= op1_03_out;
    90: reg_0316 <= op1_03_out;
    92: reg_0316 <= op1_03_out;
    94: reg_0316 <= op1_03_out;
    96: reg_0316 <= op1_03_out;
    endcase
  end

  // REG#317の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0317 <= imem03_in[39:36];
    24: reg_0317 <= imem03_in[19:16];
    26: reg_0317 <= imem06_in[59:56];
    28: reg_0317 <= imem06_in[59:56];
    31: reg_0317 <= imem03_in[39:36];
    54: reg_0317 <= imem06_in[59:56];
    56: reg_0317 <= imem06_in[59:56];
    60: reg_0317 <= imem06_in[59:56];
    62: reg_0317 <= imem03_in[39:36];
    64: reg_0317 <= imem03_in[19:16];
    66: reg_0317 <= imem03_in[39:36];
    68: reg_0317 <= imem07_in[39:36];
    70: reg_0317 <= imem06_in[59:56];
    72: reg_0317 <= imem06_in[59:56];
    74: reg_0317 <= imem06_in[59:56];
    76: reg_0317 <= imem03_in[19:16];
    78: reg_0317 <= imem03_in[19:16];
    80: reg_0317 <= imem03_in[39:36];
    82: reg_0317 <= imem06_in[59:56];
    84: reg_0317 <= imem03_in[39:36];
    86: reg_0317 <= imem07_in[39:36];
    88: reg_0317 <= imem03_in[39:36];
    endcase
  end

  // REG#318の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0318 <= imem02_in[59:56];
    24: reg_0318 <= imem03_in[47:44];
    26: reg_0318 <= imem02_in[59:56];
    53: reg_0318 <= imem03_in[47:44];
    57: reg_0318 <= imem02_in[59:56];
    59: reg_0318 <= imem03_in[107:104];
    61: reg_0318 <= imem03_in[47:44];
    63: reg_0318 <= imem03_in[107:104];
    65: reg_0318 <= imem02_in[59:56];
    67: reg_0318 <= imem02_in[87:84];
    69: reg_0318 <= imem03_in[107:104];
    71: reg_0318 <= imem03_in[47:44];
    73: reg_0318 <= imem03_in[47:44];
    75: reg_0318 <= imem02_in[87:84];
    77: reg_0318 <= imem02_in[87:84];
    79: reg_0318 <= imem03_in[47:44];
    82: reg_0318 <= imem03_in[107:104];
    84: reg_0318 <= imem03_in[107:104];
    86: reg_0318 <= imem02_in[87:84];
    88: reg_0318 <= imem02_in[87:84];
    90: reg_0318 <= imem03_in[107:104];
    endcase
  end

  // REG#319の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0319 <= imem03_in[59:56];
    24: reg_0319 <= imem05_in[15:12];
    26: reg_0319 <= imem00_in[19:16];
    28: reg_0319 <= imem05_in[15:12];
    30: reg_0319 <= imem03_in[59:56];
    33: reg_0319 <= imem03_in[59:56];
    35: reg_0319 <= imem05_in[15:12];
    37: reg_0319 <= imem03_in[59:56];
    39: reg_0319 <= imem03_in[59:56];
    41: reg_0319 <= imem00_in[19:16];
    43: reg_0319 <= imem05_in[55:52];
    45: reg_0319 <= imem03_in[15:12];
    47: reg_0319 <= imem03_in[59:56];
    49: reg_0319 <= imem03_in[59:56];
    51: reg_0319 <= imem00_in[19:16];
    53: reg_0319 <= imem00_in[19:16];
    55: reg_0319 <= imem05_in[55:52];
    58: reg_0319 <= imem03_in[59:56];
    60: reg_0319 <= imem03_in[59:56];
    62: reg_0319 <= imem03_in[59:56];
    64: reg_0319 <= imem05_in[15:12];
    67: reg_0319 <= imem02_in[7:4];
    69: reg_0319 <= imem05_in[15:12];
    71: reg_0319 <= imem00_in[19:16];
    73: reg_0319 <= imem05_in[55:52];
    95: reg_0319 <= imem05_in[55:52];
    endcase
  end

  // REG#320の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0320 <= imem02_in[31:28];
    25: reg_0320 <= imem02_in[31:28];
    28: reg_0320 <= imem07_in[111:108];
    30: reg_0320 <= imem07_in[111:108];
    32: reg_0320 <= imem02_in[31:28];
    34: reg_0320 <= imem07_in[35:32];
    36: reg_0320 <= imem00_in[7:4];
    38: reg_0320 <= imem07_in[111:108];
    40: reg_0320 <= imem07_in[111:108];
    42: reg_0320 <= imem07_in[35:32];
    44: reg_0320 <= imem07_in[111:108];
    46: reg_0320 <= imem06_in[103:100];
    48: reg_0320 <= imem07_in[51:48];
    50: reg_0320 <= imem00_in[7:4];
    52: reg_0320 <= imem07_in[51:48];
    54: reg_0320 <= imem07_in[51:48];
    56: reg_0320 <= imem07_in[51:48];
    58: reg_0320 <= imem07_in[51:48];
    60: reg_0320 <= imem06_in[103:100];
    63: reg_0320 <= imem07_in[35:32];
    65: reg_0320 <= imem06_in[103:100];
    67: reg_0320 <= imem07_in[111:108];
    69: reg_0320 <= imem07_in[111:108];
    71: reg_0320 <= imem06_in[103:100];
    82: reg_0320 <= imem06_in[103:100];
    84: reg_0320 <= imem06_in[103:100];
    86: reg_0320 <= imem06_in[103:100];
    92: reg_0320 <= imem02_in[31:28];
    94: reg_0320 <= imem02_in[31:28];
    96: reg_0320 <= imem07_in[111:108];
    endcase
  end

  // REG#321の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0321 <= imem03_in[23:20];
    25: reg_0321 <= imem07_in[91:88];
    27: reg_0321 <= imem03_in[23:20];
    30: reg_0321 <= imem03_in[23:20];
    33: reg_0321 <= imem07_in[51:48];
    35: reg_0321 <= imem02_in[111:108];
    37: reg_0321 <= imem07_in[91:88];
    39: reg_0321 <= imem07_in[51:48];
    41: reg_0321 <= imem03_in[23:20];
    43: reg_0321 <= imem07_in[51:48];
    endcase
  end

  // REG#322の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0322 <= imem03_in[79:76];
    25: reg_0322 <= imem07_in[103:100];
    27: reg_0322 <= imem05_in[83:80];
    29: reg_0322 <= imem05_in[83:80];
    31: reg_0322 <= imem03_in[79:76];
    45: reg_0322 <= imem03_in[79:76];
    47: reg_0322 <= imem00_in[51:48];
    49: reg_0322 <= imem00_in[51:48];
    51: reg_0322 <= imem03_in[79:76];
    53: reg_0322 <= imem07_in[119:116];
    55: reg_0322 <= imem03_in[79:76];
    89: reg_0322 <= imem07_in[103:100];
    91: reg_0322 <= imem07_in[103:100];
    93: reg_0322 <= imem00_in[51:48];
    95: reg_0322 <= imem07_in[119:116];
    endcase
  end

  // REG#323の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0323 <= imem03_in[83:80];
    25: reg_0323 <= imem00_in[123:120];
    27: reg_0323 <= imem03_in[83:80];
    30: reg_0323 <= imem00_in[75:72];
    32: reg_0323 <= imem02_in[15:12];
    34: reg_0323 <= imem00_in[75:72];
    36: reg_0323 <= imem01_in[123:120];
    38: reg_0323 <= imem02_in[15:12];
    40: reg_0323 <= imem00_in[123:120];
    42: reg_0323 <= imem00_in[123:120];
    44: reg_0323 <= imem03_in[91:88];
    46: reg_0323 <= imem00_in[75:72];
    48: reg_0323 <= imem02_in[15:12];
    50: reg_0323 <= imem00_in[123:120];
    52: reg_0323 <= imem02_in[15:12];
    endcase
  end

  // REG#324の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0324 <= imem02_in[79:76];
    25: reg_0324 <= imem02_in[79:76];
    28: reg_0324 <= imem00_in[59:56];
    30: reg_0324 <= imem00_in[59:56];
    32: reg_0324 <= imem02_in[79:76];
    34: reg_0324 <= imem00_in[19:16];
    36: reg_0324 <= imem00_in[59:56];
    38: reg_0324 <= imem00_in[59:56];
    40: reg_0324 <= imem02_in[79:76];
    42: reg_0324 <= imem00_in[59:56];
    44: reg_0324 <= imem00_in[19:16];
    46: reg_0324 <= imem02_in[79:76];
    48: reg_0324 <= imem00_in[19:16];
    50: reg_0324 <= imem00_in[19:16];
    52: reg_0324 <= imem00_in[19:16];
    54: reg_0324 <= imem02_in[91:88];
    56: reg_0324 <= imem00_in[59:56];
    58: reg_0324 <= imem02_in[79:76];
    60: reg_0324 <= imem00_in[79:76];
    62: reg_0324 <= imem00_in[79:76];
    64: reg_0324 <= imem06_in[11:8];
    66: reg_0324 <= imem04_in[47:44];
    68: reg_0324 <= imem00_in[79:76];
    70: reg_0324 <= imem00_in[19:16];
    72: reg_0324 <= imem00_in[19:16];
    74: reg_0324 <= imem00_in[59:56];
    76: reg_0324 <= imem04_in[7:4];
    78: reg_0324 <= imem00_in[19:16];
    80: reg_0324 <= imem00_in[79:76];
    82: reg_0324 <= imem04_in[7:4];
    84: reg_0324 <= imem00_in[19:16];
    86: reg_0324 <= imem00_in[79:76];
    88: reg_0324 <= imem02_in[79:76];
    90: reg_0324 <= imem00_in[79:76];
    93: reg_0324 <= imem02_in[91:88];
    95: reg_0324 <= imem02_in[91:88];
    97: reg_0324 <= imem02_in[79:76];
    endcase
  end

  // REG#325の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0325 <= imem02_in[23:20];
    25: reg_0325 <= imem05_in[59:56];
    27: reg_0325 <= imem07_in[27:24];
    29: reg_0325 <= imem07_in[27:24];
    31: reg_0325 <= imem05_in[59:56];
    33: reg_0325 <= imem05_in[59:56];
    35: reg_0325 <= imem05_in[59:56];
    37: reg_0325 <= imem07_in[27:24];
    39: reg_0325 <= imem05_in[59:56];
    41: reg_0325 <= imem05_in[59:56];
    43: reg_0325 <= imem07_in[27:24];
    endcase
  end

  // REG#326の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0326 <= imem02_in[35:32];
    25: reg_0326 <= imem07_in[119:116];
    27: reg_0326 <= imem07_in[119:116];
    29: reg_0326 <= imem07_in[119:116];
    31: reg_0326 <= imem02_in[35:32];
    33: reg_0326 <= imem02_in[35:32];
    35: reg_0326 <= imem02_in[35:32];
    37: reg_0326 <= imem02_in[35:32];
    39: reg_0326 <= imem07_in[119:116];
    41: reg_0326 <= imem05_in[87:84];
    43: reg_0326 <= imem05_in[87:84];
    45: reg_0326 <= imem02_in[35:32];
    64: reg_0326 <= imem06_in[35:32];
    66: reg_0326 <= imem06_in[35:32];
    68: reg_0326 <= imem05_in[87:84];
    74: reg_0326 <= imem05_in[87:84];
    96: reg_0326 <= imem07_in[119:116];
    endcase
  end

  // REG#327の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0327 <= imem03_in[71:68];
    25: reg_0327 <= imem00_in[59:56];
    27: reg_0327 <= imem00_in[59:56];
    29: reg_0327 <= imem07_in[19:16];
    31: reg_0327 <= imem03_in[71:68];
    55: reg_0327 <= imem03_in[71:68];
    89: reg_0327 <= imem03_in[71:68];
    92: reg_0327 <= imem00_in[59:56];
    94: reg_0327 <= imem03_in[71:68];
    endcase
  end

  // REG#328の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0328 <= imem02_in[115:112];
    25: reg_0328 <= imem02_in[115:112];
    28: reg_0328 <= imem01_in[123:120];
    30: reg_0328 <= imem00_in[99:96];
    32: reg_0328 <= imem01_in[123:120];
    34: reg_0328 <= imem02_in[115:112];
    36: reg_0328 <= imem00_in[99:96];
    38: reg_0328 <= imem02_in[115:112];
    40: reg_0328 <= imem06_in[103:100];
    42: reg_0328 <= imem00_in[99:96];
    44: reg_0328 <= imem00_in[99:96];
    46: reg_0328 <= imem00_in[99:96];
    48: reg_0328 <= imem07_in[55:52];
    50: reg_0328 <= imem00_in[99:96];
    52: reg_0328 <= imem07_in[55:52];
    54: reg_0328 <= imem00_in[99:96];
    57: reg_0328 <= imem06_in[103:100];
    endcase
  end

  // REG#329の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0329 <= imem02_in[55:52];
    26: reg_0329 <= imem00_in[39:36];
    28: reg_0329 <= imem02_in[55:52];
    30: reg_0329 <= imem00_in[39:36];
    32: reg_0329 <= imem00_in[39:36];
    34: reg_0329 <= imem00_in[91:88];
    36: reg_0329 <= imem02_in[55:52];
    38: reg_0329 <= imem02_in[55:52];
    40: reg_0329 <= imem07_in[127:124];
    42: reg_0329 <= imem00_in[39:36];
    44: reg_0329 <= imem07_in[127:124];
    46: reg_0329 <= imem00_in[39:36];
    48: reg_0329 <= imem07_in[127:124];
    50: reg_0329 <= imem03_in[67:64];
    52: reg_0329 <= imem02_in[55:52];
    endcase
  end

  // REG#330の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0330 <= imem02_in[63:60];
    26: reg_0330 <= imem02_in[63:60];
    53: reg_0330 <= imem00_in[55:52];
    55: reg_0330 <= imem02_in[63:60];
    57: reg_0330 <= imem02_in[63:60];
    59: reg_0330 <= imem07_in[59:56];
    61: reg_0330 <= imem07_in[59:56];
    63: reg_0330 <= imem07_in[59:56];
    65: reg_0330 <= imem02_in[55:52];
    67: reg_0330 <= imem02_in[63:60];
    69: reg_0330 <= imem00_in[55:52];
    71: reg_0330 <= imem02_in[63:60];
    74: reg_0330 <= imem02_in[63:60];
    76: reg_0330 <= imem02_in[55:52];
    78: reg_0330 <= imem05_in[87:84];
    81: reg_0330 <= imem02_in[63:60];
    83: reg_0330 <= imem02_in[55:52];
    85: reg_0330 <= imem05_in[87:84];
    87: reg_0330 <= imem05_in[87:84];
    endcase
  end

  // REG#331の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0331 <= imem03_in[127:124];
    26: reg_0331 <= imem04_in[15:12];
    28: reg_0331 <= imem04_in[15:12];
    30: reg_0331 <= imem03_in[127:124];
    32: reg_0331 <= imem04_in[15:12];
    34: reg_0331 <= imem03_in[127:124];
    36: reg_0331 <= imem03_in[127:124];
    38: reg_0331 <= imem04_in[15:12];
    40: reg_0331 <= imem03_in[127:124];
    42: reg_0331 <= imem03_in[127:124];
    44: reg_0331 <= imem03_in[127:124];
    46: reg_0331 <= imem02_in[87:84];
    48: reg_0331 <= imem02_in[87:84];
    50: reg_0331 <= imem03_in[127:124];
    52: reg_0331 <= imem02_in[87:84];
    88: reg_0331 <= imem03_in[127:124];
    endcase
  end

  // REG#332の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0332 <= imem06_in[11:8];
    26: reg_0332 <= imem04_in[103:100];
    28: reg_0332 <= imem04_in[103:100];
    30: reg_0332 <= imem06_in[11:8];
    32: reg_0332 <= imem06_in[11:8];
    37: reg_0332 <= imem06_in[11:8];
    59: reg_0332 <= imem04_in[103:100];
    endcase
  end

  // REG#333の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0333 <= imem02_in[11:8];
    26: reg_0333 <= imem05_in[107:104];
    28: reg_0333 <= imem02_in[19:16];
    30: reg_0333 <= imem02_in[11:8];
    32: reg_0333 <= imem03_in[19:16];
    34: reg_0333 <= imem02_in[11:8];
    36: reg_0333 <= imem02_in[19:16];
    38: reg_0333 <= imem00_in[119:116];
    40: reg_0333 <= imem00_in[119:116];
    42: reg_0333 <= imem05_in[107:104];
    44: reg_0333 <= imem00_in[119:116];
    46: reg_0333 <= imem02_in[19:16];
    48: reg_0333 <= imem03_in[19:16];
    50: reg_0333 <= imem05_in[107:104];
    66: reg_0333 <= imem05_in[107:104];
    79: reg_0333 <= imem03_in[19:16];
    81: reg_0333 <= imem02_in[11:8];
    83: reg_0333 <= imem05_in[107:104];
    85: reg_0333 <= imem03_in[19:16];
    87: reg_0333 <= imem02_in[11:8];
    89: reg_0333 <= imem02_in[19:16];
    91: reg_0333 <= imem00_in[119:116];
    endcase
  end

  // REG#334の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0334 <= imem02_in[7:4];
    26: reg_0334 <= imem02_in[7:4];
    52: reg_0334 <= imem04_in[107:104];
    54: reg_0334 <= imem04_in[107:104];
    56: reg_0334 <= imem04_in[107:104];
    58: reg_0334 <= imem02_in[63:60];
    60: reg_0334 <= imem01_in[39:36];
    62: reg_0334 <= imem04_in[107:104];
    64: reg_0334 <= imem01_in[39:36];
    66: reg_0334 <= imem04_in[107:104];
    68: reg_0334 <= imem02_in[7:4];
    70: reg_0334 <= imem02_in[7:4];
    72: reg_0334 <= imem04_in[107:104];
    74: reg_0334 <= imem04_in[51:48];
    76: reg_0334 <= imem04_in[51:48];
    78: reg_0334 <= imem05_in[23:20];
    82: reg_0334 <= imem04_in[51:48];
    84: reg_0334 <= imem02_in[7:4];
    endcase
  end

  // REG#335の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0335 <= imem02_in[111:108];
    26: reg_0335 <= imem02_in[111:108];
    52: reg_0335 <= imem02_in[111:108];
    endcase
  end

  // REG#336の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0336 <= imem02_in[127:124];
    26: reg_0336 <= imem02_in[127:124];
    50: reg_0336 <= imem05_in[75:72];
    63: reg_0336 <= imem02_in[127:124];
    71: reg_0336 <= imem00_in[43:40];
    73: reg_0336 <= imem00_in[43:40];
    75: reg_0336 <= imem00_in[43:40];
    77: reg_0336 <= imem00_in[43:40];
    79: reg_0336 <= imem05_in[75:72];
    88: reg_0336 <= imem06_in[19:16];
    90: reg_0336 <= imem02_in[127:124];
    92: reg_0336 <= imem02_in[119:116];
    94: reg_0336 <= imem00_in[43:40];
    96: reg_0336 <= imem00_in[43:40];
    endcase
  end

  // REG#337の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0337 <= imem06_in[119:116];
    26: reg_0337 <= imem05_in[127:124];
    28: reg_0337 <= imem05_in[127:124];
    30: reg_0337 <= imem01_in[47:44];
    32: reg_0337 <= imem04_in[11:8];
    34: reg_0337 <= imem04_in[11:8];
    36: reg_0337 <= imem04_in[11:8];
    38: reg_0337 <= imem04_in[11:8];
    40: reg_0337 <= imem01_in[47:44];
    42: reg_0337 <= imem05_in[127:124];
    44: reg_0337 <= imem05_in[127:124];
    46: reg_0337 <= imem05_in[127:124];
    48: reg_0337 <= imem04_in[11:8];
    51: reg_0337 <= imem01_in[47:44];
    53: reg_0337 <= imem04_in[11:8];
    55: reg_0337 <= imem01_in[47:44];
    57: reg_0337 <= imem01_in[47:44];
    59: reg_0337 <= imem01_in[47:44];
    61: reg_0337 <= imem05_in[127:124];
    65: reg_0337 <= imem04_in[11:8];
    67: reg_0337 <= imem04_in[11:8];
    69: reg_0337 <= imem01_in[47:44];
    94: reg_0337 <= imem04_in[11:8];
    96: reg_0337 <= imem04_in[11:8];
    endcase
  end

  // REG#338の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0338 <= imem02_in[99:96];
    26: reg_0338 <= imem02_in[99:96];
    49: reg_0338 <= imem06_in[87:84];
    51: reg_0338 <= imem06_in[87:84];
    53: reg_0338 <= imem02_in[99:96];
    55: reg_0338 <= imem06_in[99:96];
    57: reg_0338 <= imem06_in[87:84];
    endcase
  end

  // REG#339の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0339 <= imem02_in[71:68];
    26: reg_0339 <= imem02_in[71:68];
    53: reg_0339 <= imem02_in[71:68];
    55: reg_0339 <= imem07_in[55:52];
    57: reg_0339 <= imem01_in[107:104];
    59: reg_0339 <= imem00_in[87:84];
    61: reg_0339 <= imem00_in[87:84];
    63: reg_0339 <= imem00_in[87:84];
    65: reg_0339 <= imem02_in[91:88];
    67: reg_0339 <= imem00_in[87:84];
    69: reg_0339 <= imem02_in[91:88];
    71: reg_0339 <= imem07_in[55:52];
    73: reg_0339 <= imem00_in[87:84];
    75: reg_0339 <= imem07_in[55:52];
    78: reg_0339 <= imem01_in[107:104];
    80: reg_0339 <= imem02_in[91:88];
    82: reg_0339 <= imem07_in[55:52];
    endcase
  end

  // REG#340の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0340 <= op1_04_out;
    25: reg_0340 <= op1_04_out;
    27: reg_0340 <= op1_04_out;
    29: reg_0340 <= op1_04_out;
    31: reg_0340 <= op1_04_out;
    33: reg_0340 <= op1_04_out;
    35: reg_0340 <= op1_04_out;
    37: reg_0340 <= op1_04_out;
    39: reg_0340 <= op1_04_out;
    41: reg_0340 <= op1_04_out;
    43: reg_0340 <= op1_04_out;
    45: reg_0340 <= op1_04_out;
    47: reg_0340 <= op1_04_out;
    49: reg_0340 <= op1_04_out;
    51: reg_0340 <= op1_04_out;
    53: reg_0340 <= op1_04_out;
    55: reg_0340 <= op1_04_out;
    57: reg_0340 <= op1_04_out;
    59: reg_0340 <= op1_04_out;
    61: reg_0340 <= op1_04_out;
    63: reg_0340 <= op1_04_out;
    65: reg_0340 <= op1_04_out;
    67: reg_0340 <= op1_04_out;
    69: reg_0340 <= op1_04_out;
    71: reg_0340 <= op1_04_out;
    73: reg_0340 <= op1_04_out;
    75: reg_0340 <= op1_04_out;
    77: reg_0340 <= op1_04_out;
    79: reg_0340 <= op1_04_out;
    81: reg_0340 <= op1_04_out;
    83: reg_0340 <= op1_04_out;
    85: reg_0340 <= op1_04_out;
    87: reg_0340 <= op1_04_out;
    89: reg_0340 <= op1_04_out;
    91: reg_0340 <= op1_04_out;
    93: reg_0340 <= op1_04_out;
    95: reg_0340 <= op1_04_out;
    97: reg_0340 <= op1_04_out;
    endcase
  end

  // REG#341の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0341 <= imem02_in[43:40];
    27: reg_0341 <= imem02_in[43:40];
    29: reg_0341 <= imem02_in[43:40];
    31: reg_0341 <= imem02_in[43:40];
    33: reg_0341 <= imem02_in[43:40];
    35: reg_0341 <= imem02_in[43:40];
    37: reg_0341 <= imem02_in[107:104];
    39: reg_0341 <= imem02_in[43:40];
    41: reg_0341 <= imem02_in[107:104];
    43: reg_0341 <= imem02_in[43:40];
    45: reg_0341 <= imem02_in[43:40];
    63: reg_0341 <= imem02_in[43:40];
    72: reg_0341 <= imem02_in[107:104];
    83: reg_0341 <= imem02_in[107:104];
    85: reg_0341 <= imem02_in[107:104];
    endcase
  end

  // REG#342の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0342 <= imem02_in[95:92];
    27: reg_0342 <= imem07_in[71:68];
    29: reg_0342 <= imem07_in[71:68];
    31: reg_0342 <= imem02_in[95:92];
    33: reg_0342 <= imem02_in[95:92];
    35: reg_0342 <= imem03_in[91:88];
    37: reg_0342 <= imem07_in[71:68];
    39: reg_0342 <= imem03_in[115:112];
    41: reg_0342 <= imem02_in[95:92];
    43: reg_0342 <= imem03_in[91:88];
    45: reg_0342 <= imem03_in[91:88];
    47: reg_0342 <= imem03_in[91:88];
    49: reg_0342 <= imem07_in[83:80];
    51: reg_0342 <= imem07_in[71:68];
    53: reg_0342 <= imem03_in[115:112];
    56: reg_0342 <= imem07_in[83:80];
    58: reg_0342 <= imem07_in[83:80];
    60: reg_0342 <= imem03_in[91:88];
    62: reg_0342 <= imem07_in[83:80];
    64: reg_0342 <= imem07_in[83:80];
    66: reg_0342 <= imem07_in[83:80];
    68: reg_0342 <= imem02_in[95:92];
    70: reg_0342 <= imem07_in[83:80];
    72: reg_0342 <= imem07_in[71:68];
    74: reg_0342 <= imem07_in[71:68];
    76: reg_0342 <= imem02_in[95:92];
    78: reg_0342 <= imem07_in[71:68];
    80: reg_0342 <= imem07_in[71:68];
    84: reg_0342 <= imem03_in[91:88];
    86: reg_0342 <= imem04_in[35:32];
    88: reg_0342 <= imem03_in[115:112];
    endcase
  end

  // REG#343の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0343 <= imem03_in[43:40];
    27: reg_0343 <= imem03_in[43:40];
    29: reg_0343 <= imem07_in[103:100];
    31: reg_0343 <= imem03_in[43:40];
    51: reg_0343 <= imem03_in[43:40];
    53: reg_0343 <= imem03_in[43:40];
    56: reg_0343 <= imem05_in[123:120];
    58: reg_0343 <= imem03_in[43:40];
    60: reg_0343 <= imem03_in[43:40];
    62: reg_0343 <= imem07_in[103:100];
    64: reg_0343 <= imem06_in[83:80];
    66: reg_0343 <= imem06_in[83:80];
    68: reg_0343 <= imem05_in[123:120];
    74: reg_0343 <= imem06_in[83:80];
    76: reg_0343 <= imem06_in[83:80];
    78: reg_0343 <= imem05_in[123:120];
    80: reg_0343 <= imem06_in[83:80];
    82: reg_0343 <= imem06_in[83:80];
    84: reg_0343 <= imem03_in[43:40];
    86: reg_0343 <= imem06_in[83:80];
    93: reg_0343 <= imem07_in[103:100];
    95: reg_0343 <= imem06_in[83:80];
    endcase
  end

  // REG#344の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0344 <= imem06_in[23:20];
    27: reg_0344 <= imem00_in[75:72];
    29: reg_0344 <= imem06_in[23:20];
    57: reg_0344 <= imem06_in[23:20];
    91: reg_0344 <= imem00_in[75:72];
    endcase
  end

  // REG#345の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0345 <= imem02_in[51:48];
    27: reg_0345 <= imem02_in[51:48];
    29: reg_0345 <= imem00_in[35:32];
    31: reg_0345 <= imem00_in[35:32];
    33: reg_0345 <= imem00_in[35:32];
    35: reg_0345 <= imem00_in[35:32];
    37: reg_0345 <= imem03_in[23:20];
    39: reg_0345 <= imem03_in[123:120];
    41: reg_0345 <= imem00_in[35:32];
    43: reg_0345 <= imem03_in[23:20];
    45: reg_0345 <= imem03_in[123:120];
    47: reg_0345 <= imem00_in[35:32];
    49: reg_0345 <= imem03_in[123:120];
    51: reg_0345 <= imem00_in[35:32];
    53: reg_0345 <= imem00_in[35:32];
    55: reg_0345 <= imem03_in[23:20];
    89: reg_0345 <= imem03_in[123:120];
    91: reg_0345 <= imem00_in[35:32];
    endcase
  end

  // REG#346の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0346 <= imem02_in[75:72];
    27: reg_0346 <= imem03_in[103:100];
    29: reg_0346 <= imem02_in[75:72];
    31: reg_0346 <= imem03_in[103:100];
    55: reg_0346 <= imem03_in[103:100];
    86: reg_0346 <= imem03_in[103:100];
    88: reg_0346 <= imem03_in[103:100];
    endcase
  end

  // REG#347の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0347 <= imem02_in[123:120];
    27: reg_0347 <= imem05_in[63:60];
    29: reg_0347 <= imem05_in[63:60];
    31: reg_0347 <= imem05_in[63:60];
    33: reg_0347 <= imem02_in[123:120];
    35: reg_0347 <= imem02_in[123:120];
    37: reg_0347 <= imem05_in[63:60];
    39: reg_0347 <= imem04_in[99:96];
    41: reg_0347 <= imem04_in[99:96];
    44: reg_0347 <= imem05_in[63:60];
    46: reg_0347 <= imem05_in[63:60];
    48: reg_0347 <= imem05_in[63:60];
    50: reg_0347 <= imem02_in[123:120];
    52: reg_0347 <= imem02_in[123:120];
    endcase
  end

  // REG#348の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0348 <= imem06_in[7:4];
    27: reg_0348 <= imem06_in[15:12];
    29: reg_0348 <= imem06_in[15:12];
    59: reg_0348 <= imem02_in[75:72];
    61: reg_0348 <= imem06_in[15:12];
    70: reg_0348 <= imem06_in[7:4];
    72: reg_0348 <= imem06_in[7:4];
    74: reg_0348 <= imem06_in[7:4];
    76: reg_0348 <= imem06_in[7:4];
    78: reg_0348 <= imem02_in[75:72];
    80: reg_0348 <= imem02_in[75:72];
    82: reg_0348 <= imem06_in[7:4];
    84: reg_0348 <= imem02_in[75:72];
    endcase
  end

  // REG#349の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0349 <= imem06_in[39:36];
    27: reg_0349 <= imem06_in[107:104];
    29: reg_0349 <= imem06_in[107:104];
    53: reg_0349 <= imem02_in[103:100];
    55: reg_0349 <= imem05_in[111:108];
    57: reg_0349 <= imem02_in[103:100];
    59: reg_0349 <= imem05_in[111:108];
    61: reg_0349 <= imem06_in[107:104];
    67: reg_0349 <= imem05_in[111:108];
    70: reg_0349 <= imem06_in[39:36];
    73: reg_0349 <= imem06_in[39:36];
    75: reg_0349 <= imem00_in[79:76];
    77: reg_0349 <= imem00_in[79:76];
    79: reg_0349 <= imem06_in[107:104];
    82: reg_0349 <= imem06_in[107:104];
    84: reg_0349 <= imem02_in[103:100];
    endcase
  end

  // REG#350の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0350 <= imem02_in[107:104];
    27: reg_0350 <= imem02_in[107:104];
    29: reg_0350 <= imem02_in[107:104];
    31: reg_0350 <= imem07_in[91:88];
    33: reg_0350 <= imem02_in[107:104];
    35: reg_0350 <= imem04_in[63:60];
    37: reg_0350 <= imem04_in[63:60];
    39: reg_0350 <= imem04_in[63:60];
    41: reg_0350 <= imem04_in[63:60];
    43: reg_0350 <= imem07_in[91:88];
    endcase
  end

  // REG#351の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0351 <= imem06_in[51:48];
    27: reg_0351 <= imem06_in[51:48];
    29: reg_0351 <= imem06_in[51:48];
    57: reg_0351 <= imem06_in[51:48];
    endcase
  end

  // REG#352の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0352 <= imem02_in[3:0];
    27: reg_0352 <= imem06_in[127:124];
    29: reg_0352 <= imem02_in[3:0];
    31: reg_0352 <= imem00_in[11:8];
    33: reg_0352 <= imem00_in[51:48];
    35: reg_0352 <= imem00_in[51:48];
    37: reg_0352 <= imem04_in[7:4];
    39: reg_0352 <= imem00_in[11:8];
    41: reg_0352 <= imem06_in[127:124];
    43: reg_0352 <= imem00_in[39:36];
    45: reg_0352 <= imem04_in[7:4];
    48: reg_0352 <= imem02_in[3:0];
    50: reg_0352 <= imem02_in[3:0];
    52: reg_0352 <= imem06_in[127:124];
    54: reg_0352 <= imem00_in[51:48];
    57: reg_0352 <= imem00_in[51:48];
    59: reg_0352 <= imem03_in[91:88];
    61: reg_0352 <= imem00_in[11:8];
    63: reg_0352 <= imem00_in[39:36];
    65: reg_0352 <= imem00_in[51:48];
    67: reg_0352 <= imem00_in[51:48];
    69: reg_0352 <= imem00_in[51:48];
    71: reg_0352 <= imem00_in[51:48];
    73: reg_0352 <= imem04_in[7:4];
    75: reg_0352 <= imem00_in[39:36];
    77: reg_0352 <= imem00_in[51:48];
    79: reg_0352 <= imem00_in[11:8];
    81: reg_0352 <= imem00_in[51:48];
    83: reg_0352 <= imem02_in[3:0];
    87: reg_0352 <= imem00_in[39:36];
    89: reg_0352 <= imem03_in[91:88];
    92: reg_0352 <= imem00_in[39:36];
    94: reg_0352 <= imem03_in[91:88];
    96: reg_0352 <= imem02_in[3:0];
    endcase
  end

  // REG#353の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0353 <= imem02_in[83:80];
    27: reg_0353 <= imem07_in[79:76];
    29: reg_0353 <= imem00_in[99:96];
    31: reg_0353 <= imem02_in[83:80];
    33: reg_0353 <= imem00_in[123:120];
    35: reg_0353 <= imem00_in[99:96];
    37: reg_0353 <= imem07_in[79:76];
    39: reg_0353 <= imem02_in[83:80];
    41: reg_0353 <= imem07_in[79:76];
    43: reg_0353 <= imem07_in[79:76];
    97: reg_0353 <= imem00_in[123:120];
    endcase
  end

  // REG#354の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0354 <= imem02_in[39:36];
    27: reg_0354 <= imem00_in[63:60];
    29: reg_0354 <= imem01_in[95:92];
    31: reg_0354 <= imem02_in[39:36];
    33: reg_0354 <= imem01_in[95:92];
    35: reg_0354 <= imem02_in[39:36];
    37: reg_0354 <= imem02_in[39:36];
    39: reg_0354 <= imem02_in[39:36];
    41: reg_0354 <= imem01_in[95:92];
    93: reg_0354 <= imem02_in[39:36];
    95: reg_0354 <= imem02_in[39:36];
    endcase
  end

  // REG#355の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0355 <= imem02_in[103:100];
    27: reg_0355 <= imem02_in[103:100];
    29: reg_0355 <= imem02_in[115:112];
    31: reg_0355 <= imem02_in[103:100];
    33: reg_0355 <= imem02_in[103:100];
    35: reg_0355 <= imem05_in[99:96];
    37: reg_0355 <= imem02_in[115:112];
    39: reg_0355 <= imem07_in[15:12];
    41: reg_0355 <= imem00_in[31:28];
    43: reg_0355 <= imem02_in[15:12];
    45: reg_0355 <= imem02_in[15:12];
    55: reg_0355 <= imem02_in[115:112];
    57: reg_0355 <= imem07_in[15:12];
    59: reg_0355 <= imem02_in[115:112];
    61: reg_0355 <= imem02_in[115:112];
    63: reg_0355 <= imem02_in[15:12];
    71: reg_0355 <= imem07_in[15:12];
    73: reg_0355 <= imem02_in[15:12];
    75: reg_0355 <= imem02_in[115:112];
    77: reg_0355 <= imem00_in[119:116];
    79: reg_0355 <= imem02_in[115:112];
    81: reg_0355 <= imem05_in[99:96];
    83: reg_0355 <= imem00_in[119:116];
    85: reg_0355 <= imem02_in[15:12];
    94: reg_0355 <= imem02_in[103:100];
    96: reg_0355 <= imem02_in[103:100];
    endcase
  end

  // REG#356の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0356 <= imem06_in[19:16];
    27: reg_0356 <= imem00_in[79:76];
    29: reg_0356 <= imem06_in[19:16];
    55: reg_0356 <= imem00_in[79:76];
    92: reg_0356 <= imem00_in[79:76];
    94: reg_0356 <= imem00_in[79:76];
    97: reg_0356 <= imem06_in[19:16];
    endcase
  end

  // REG#357の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0357 <= imem02_in[15:12];
    27: reg_0357 <= imem02_in[15:12];
    29: reg_0357 <= imem03_in[35:32];
    31: reg_0357 <= imem03_in[35:32];
    55: reg_0357 <= imem03_in[35:32];
    88: reg_0357 <= imem03_in[35:32];
    endcase
  end

  // REG#358の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0358 <= imem02_in[19:16];
    27: reg_0358 <= imem00_in[111:108];
    29: reg_0358 <= imem03_in[75:72];
    31: reg_0358 <= imem03_in[75:72];
    52: reg_0358 <= imem02_in[19:16];
    endcase
  end

  // REG#359の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0359 <= imem02_in[47:44];
    27: reg_0359 <= imem02_in[47:44];
    29: reg_0359 <= imem04_in[27:24];
    31: reg_0359 <= imem00_in[71:68];
    33: reg_0359 <= imem00_in[71:68];
    35: reg_0359 <= imem07_in[103:100];
    37: reg_0359 <= imem07_in[103:100];
    39: reg_0359 <= imem02_in[47:44];
    41: reg_0359 <= imem02_in[47:44];
    43: reg_0359 <= imem00_in[71:68];
    45: reg_0359 <= imem02_in[47:44];
    52: reg_0359 <= imem02_in[47:44];
    96: reg_0359 <= imem04_in[27:24];
    endcase
  end

  // REG#360の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0360 <= imem03_in[27:24];
    27: reg_0360 <= imem03_in[27:24];
    30: reg_0360 <= imem03_in[27:24];
    33: reg_0360 <= imem03_in[27:24];
    35: reg_0360 <= imem00_in[39:36];
    37: reg_0360 <= imem00_in[39:36];
    39: reg_0360 <= imem01_in[103:100];
    41: reg_0360 <= imem00_in[39:36];
    43: reg_0360 <= imem01_in[103:100];
    45: reg_0360 <= imem03_in[27:24];
    47: reg_0360 <= imem00_in[39:36];
    49: reg_0360 <= imem00_in[39:36];
    51: reg_0360 <= imem02_in[115:112];
    54: reg_0360 <= imem00_in[39:36];
    56: reg_0360 <= imem01_in[103:100];
    58: reg_0360 <= imem00_in[39:36];
    60: reg_0360 <= imem00_in[39:36];
    62: reg_0360 <= imem02_in[115:112];
    64: reg_0360 <= imem00_in[39:36];
    66: reg_0360 <= imem00_in[39:36];
    68: reg_0360 <= imem01_in[103:100];
    71: reg_0360 <= imem02_in[115:112];
    74: reg_0360 <= imem00_in[39:36];
    76: reg_0360 <= imem00_in[39:36];
    78: reg_0360 <= imem05_in[3:0];
    81: reg_0360 <= imem03_in[27:24];
    83: reg_0360 <= imem02_in[119:116];
    87: reg_0360 <= imem02_in[119:116];
    89: reg_0360 <= imem02_in[115:112];
    91: reg_0360 <= imem01_in[103:100];
    93: reg_0360 <= imem02_in[119:116];
    95: reg_0360 <= imem02_in[119:116];
    97: reg_0360 <= imem03_in[27:24];
    endcase
  end

  // REG#361の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0361 <= imem03_in[107:104];
    27: reg_0361 <= imem00_in[119:116];
    29: reg_0361 <= imem07_in[7:4];
    31: reg_0361 <= imem00_in[119:116];
    33: reg_0361 <= imem01_in[19:16];
    35: reg_0361 <= imem07_in[7:4];
    37: reg_0361 <= imem00_in[119:116];
    39: reg_0361 <= imem03_in[35:32];
    41: reg_0361 <= imem03_in[35:32];
    43: reg_0361 <= imem07_in[7:4];
    endcase
  end

  // REG#362の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0362 <= imem03_in[51:48];
    27: reg_0362 <= imem03_in[51:48];
    28: reg_0362 <= op2_00_out;
    40: reg_0362 <= op2_00_out;
    79: reg_0362 <= op2_00_out;
    endcase
  end

  // REG#363の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0363 <= imem02_in[67:64];
    27: reg_0363 <= imem01_in[7:4];
    29: reg_0363 <= imem02_in[67:64];
    31: reg_0363 <= imem01_in[7:4];
    33: reg_0363 <= imem02_in[11:8];
    35: reg_0363 <= imem02_in[11:8];
    37: reg_0363 <= imem02_in[11:8];
    39: reg_0363 <= imem01_in[7:4];
    41: reg_0363 <= imem02_in[11:8];
    43: reg_0363 <= imem03_in[3:0];
    45: reg_0363 <= imem02_in[11:8];
    62: reg_0363 <= imem02_in[11:8];
    65: reg_0363 <= imem03_in[75:72];
    67: reg_0363 <= imem02_in[11:8];
    69: reg_0363 <= imem03_in[75:72];
    71: reg_0363 <= imem03_in[75:72];
    73: reg_0363 <= imem01_in[7:4];
    75: reg_0363 <= imem02_in[67:64];
    78: reg_0363 <= imem03_in[3:0];
    80: reg_0363 <= imem01_in[7:4];
    82: reg_0363 <= imem03_in[3:0];
    84: reg_0363 <= imem01_in[7:4];
    86: reg_0363 <= imem01_in[7:4];
    88: reg_0363 <= imem03_in[75:72];
    endcase
  end

  // REG#364の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0364 <= imem02_in[27:24];
    27: reg_0364 <= imem02_in[27:24];
    29: reg_0364 <= imem02_in[27:24];
    31: reg_0364 <= imem00_in[107:104];
    33: reg_0364 <= imem02_in[27:24];
    35: reg_0364 <= imem02_in[27:24];
    37: reg_0364 <= imem04_in[111:108];
    39: reg_0364 <= imem00_in[107:104];
    41: reg_0364 <= imem04_in[111:108];
    43: reg_0364 <= imem02_in[27:24];
    45: reg_0364 <= imem04_in[111:108];
    48: reg_0364 <= imem04_in[111:108];
    52: reg_0364 <= imem04_in[111:108];
    54: reg_0364 <= imem00_in[107:104];
    56: reg_0364 <= imem02_in[23:20];
    58: reg_0364 <= imem00_in[107:104];
    60: reg_0364 <= imem00_in[107:104];
    62: reg_0364 <= imem02_in[23:20];
    65: reg_0364 <= imem02_in[23:20];
    67: reg_0364 <= imem00_in[107:104];
    69: reg_0364 <= imem03_in[63:60];
    71: reg_0364 <= imem02_in[27:24];
    74: reg_0364 <= imem02_in[23:20];
    76: reg_0364 <= imem02_in[23:20];
    78: reg_0364 <= imem03_in[63:60];
    80: reg_0364 <= imem04_in[111:108];
    82: reg_0364 <= imem00_in[107:104];
    84: reg_0364 <= imem03_in[63:60];
    86: reg_0364 <= imem03_in[63:60];
    88: reg_0364 <= imem07_in[27:24];
    90: reg_0364 <= imem07_in[27:24];
    92: reg_0364 <= imem01_in[7:4];
    95: reg_0364 <= imem02_in[23:20];
    97: reg_0364 <= imem02_in[27:24];
    endcase
  end

  // REG#365の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0365 <= imem02_in[91:88];
    27: reg_0365 <= imem01_in[111:108];
    29: reg_0365 <= imem01_in[111:108];
    31: reg_0365 <= imem01_in[111:108];
    33: reg_0365 <= imem02_in[63:60];
    35: reg_0365 <= imem02_in[63:60];
    37: reg_0365 <= imem01_in[111:108];
    39: reg_0365 <= imem05_in[3:0];
    41: reg_0365 <= imem02_in[63:60];
    43: reg_0365 <= imem01_in[111:108];
    45: reg_0365 <= imem02_in[91:88];
    64: reg_0365 <= imem07_in[127:124];
    66: reg_0365 <= imem01_in[111:108];
    68: reg_0365 <= imem05_in[3:0];
    71: reg_0365 <= imem02_in[91:88];
    74: reg_0365 <= imem07_in[127:124];
    77: reg_0365 <= imem02_in[91:88];
    79: reg_0365 <= imem05_in[3:0];
    85: reg_0365 <= imem02_in[91:88];
    endcase
  end

  // REG#366の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0366 <= op1_05_out;
    26: reg_0366 <= op1_05_out;
    28: reg_0366 <= op1_05_out;
    30: reg_0366 <= op1_05_out;
    32: reg_0366 <= op1_05_out;
    34: reg_0366 <= op1_05_out;
    36: reg_0366 <= op1_05_out;
    38: reg_0366 <= op1_05_out;
    40: reg_0366 <= op1_05_out;
    42: reg_0366 <= op1_05_out;
    44: reg_0366 <= op1_05_out;
    46: reg_0366 <= op1_05_out;
    48: reg_0366 <= op1_05_out;
    50: reg_0366 <= op1_05_out;
    52: reg_0366 <= op1_05_out;
    54: reg_0366 <= op1_05_out;
    56: reg_0366 <= op1_05_out;
    58: reg_0366 <= op1_05_out;
    60: reg_0366 <= op1_05_out;
    62: reg_0366 <= op1_05_out;
    64: reg_0366 <= op1_05_out;
    66: reg_0366 <= op1_05_out;
    68: reg_0366 <= op1_05_out;
    70: reg_0366 <= op1_05_out;
    72: reg_0366 <= op1_05_out;
    74: reg_0366 <= op1_05_out;
    76: reg_0366 <= op1_05_out;
    78: reg_0366 <= op1_05_out;
    80: reg_0366 <= op1_05_out;
    82: reg_0366 <= op1_05_out;
    84: reg_0366 <= op1_05_out;
    86: reg_0366 <= op1_05_out;
    88: reg_0366 <= op1_05_out;
    90: reg_0366 <= op1_05_out;
    92: reg_0366 <= op1_05_out;
    94: reg_0366 <= op1_05_out;
    96: reg_0366 <= op1_05_out;
    endcase
  end

  // REG#367の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0367 <= imem06_in[111:108];
    28: reg_0367 <= imem06_in[111:108];
    30: reg_0367 <= imem01_in[75:72];
    32: reg_0367 <= imem06_in[111:108];
    38: reg_0367 <= imem01_in[11:8];
    40: reg_0367 <= imem01_in[75:72];
    42: reg_0367 <= imem01_in[75:72];
    44: reg_0367 <= imem04_in[35:32];
    46: reg_0367 <= imem04_in[35:32];
    50: reg_0367 <= imem04_in[35:32];
    52: reg_0367 <= imem05_in[47:44];
    54: reg_0367 <= imem06_in[111:108];
    56: reg_0367 <= imem04_in[35:32];
    58: reg_0367 <= imem04_in[35:32];
    61: reg_0367 <= imem04_in[35:32];
    63: reg_0367 <= imem01_in[11:8];
    65: reg_0367 <= imem01_in[75:72];
    67: reg_0367 <= imem02_in[111:108];
    69: reg_0367 <= imem02_in[111:108];
    71: reg_0367 <= imem01_in[75:72];
    73: reg_0367 <= imem02_in[111:108];
    75: reg_0367 <= imem00_in[83:80];
    77: reg_0367 <= imem01_in[75:72];
    79: reg_0367 <= imem06_in[111:108];
    81: reg_0367 <= imem01_in[11:8];
    83: reg_0367 <= imem00_in[83:80];
    85: reg_0367 <= imem02_in[111:108];
    endcase
  end

  // REG#368の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0368 <= imem06_in[127:124];
    28: reg_0368 <= imem06_in[55:52];
    30: reg_0368 <= imem01_in[111:108];
    32: reg_0368 <= imem01_in[111:108];
    34: reg_0368 <= imem02_in[67:64];
    36: reg_0368 <= imem01_in[111:108];
    38: reg_0368 <= imem02_in[67:64];
    40: reg_0368 <= imem01_in[111:108];
    42: reg_0368 <= imem02_in[43:40];
    44: reg_0368 <= imem01_in[111:108];
    46: reg_0368 <= imem02_in[67:64];
    48: reg_0368 <= imem02_in[67:64];
    50: reg_0368 <= imem02_in[67:64];
    52: reg_0368 <= imem02_in[67:64];
    92: reg_0368 <= imem01_in[111:108];
    endcase
  end

  // REG#369の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0369 <= imem03_in[63:60];
    28: reg_0369 <= imem03_in[63:60];
    71: reg_0369 <= imem06_in[95:92];
    90: reg_0369 <= imem06_in[95:92];
    92: reg_0369 <= imem01_in[19:16];
    endcase
  end

  // REG#370の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0370 <= imem03_in[31:28];
    28: reg_0370 <= imem03_in[31:28];
    69: reg_0370 <= imem06_in[31:28];
    71: reg_0370 <= imem06_in[31:28];
    89: reg_0370 <= imem06_in[31:28];
    endcase
  end

  // REG#371の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0371 <= imem06_in[67:64];
    28: reg_0371 <= imem06_in[67:64];
    31: reg_0371 <= imem06_in[67:64];
    33: reg_0371 <= imem06_in[67:64];
    35: reg_0371 <= imem06_in[67:64];
    37: reg_0371 <= imem05_in[83:80];
    39: reg_0371 <= imem06_in[67:64];
    57: reg_0371 <= imem05_in[83:80];
    59: reg_0371 <= imem07_in[103:100];
    61: reg_0371 <= imem06_in[67:64];
    71: reg_0371 <= imem07_in[103:100];
    73: reg_0371 <= imem07_in[103:100];
    75: reg_0371 <= imem07_in[103:100];
    80: reg_0371 <= imem07_in[103:100];
    82: reg_0371 <= imem07_in[103:100];
    endcase
  end

  // REG#372の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0372 <= imem06_in[31:28];
    28: reg_0372 <= imem06_in[31:28];
    31: reg_0372 <= imem06_in[31:28];
    34: reg_0372 <= imem05_in[23:20];
    36: reg_0372 <= imem06_in[31:28];
    40: reg_0372 <= imem00_in[23:20];
    42: reg_0372 <= imem06_in[31:28];
    44: reg_0372 <= imem06_in[31:28];
    46: reg_0372 <= imem06_in[31:28];
    48: reg_0372 <= imem00_in[55:52];
    50: reg_0372 <= imem00_in[23:20];
    52: reg_0372 <= imem02_in[79:76];
    endcase
  end

  // REG#373の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0373 <= imem03_in[55:52];
    28: reg_0373 <= imem03_in[55:52];
    72: reg_0373 <= imem03_in[15:12];
    74: reg_0373 <= imem03_in[15:12];
    76: reg_0373 <= imem04_in[95:92];
    79: reg_0373 <= imem03_in[15:12];
    82: reg_0373 <= imem03_in[15:12];
    84: reg_0373 <= imem03_in[55:52];
    86: reg_0373 <= imem03_in[15:12];
    88: reg_0373 <= imem04_in[95:92];
    90: reg_0373 <= imem03_in[15:12];
    endcase
  end

  // REG#374の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0374 <= imem03_in[119:116];
    28: reg_0374 <= imem03_in[119:116];
    69: reg_0374 <= imem07_in[63:60];
    72: reg_0374 <= imem03_in[119:116];
    74: reg_0374 <= imem07_in[63:60];
    76: reg_0374 <= imem03_in[119:116];
    79: reg_0374 <= imem07_in[63:60];
    endcase
  end

  // REG#375の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0375 <= imem06_in[75:72];
    28: reg_0375 <= imem07_in[123:120];
    30: reg_0375 <= imem02_in[23:20];
    32: reg_0375 <= imem04_in[43:40];
    34: reg_0375 <= imem04_in[43:40];
    36: reg_0375 <= imem04_in[43:40];
    38: reg_0375 <= imem07_in[123:120];
    40: reg_0375 <= imem04_in[43:40];
    42: reg_0375 <= imem03_in[71:68];
    44: reg_0375 <= imem02_in[23:20];
    46: reg_0375 <= imem02_in[23:20];
    48: reg_0375 <= imem04_in[63:60];
    50: reg_0375 <= imem02_in[23:20];
    52: reg_0375 <= imem04_in[63:60];
    54: reg_0375 <= imem00_in[115:112];
    57: reg_0375 <= imem07_in[123:120];
    59: reg_0375 <= imem07_in[123:120];
    61: reg_0375 <= imem02_in[23:20];
    63: reg_0375 <= imem00_in[115:112];
    65: reg_0375 <= imem04_in[43:40];
    67: reg_0375 <= imem04_in[63:60];
    69: reg_0375 <= imem04_in[43:40];
    71: reg_0375 <= imem02_in[23:20];
    73: reg_0375 <= imem07_in[123:120];
    75: reg_0375 <= imem02_in[23:20];
    77: reg_0375 <= imem00_in[115:112];
    79: reg_0375 <= imem03_in[71:68];
    81: reg_0375 <= imem02_in[23:20];
    83: reg_0375 <= imem03_in[71:68];
    85: reg_0375 <= imem04_in[43:40];
    87: reg_0375 <= imem04_in[43:40];
    89: reg_0375 <= imem04_in[43:40];
    91: reg_0375 <= imem03_in[71:68];
    93: reg_0375 <= imem00_in[115:112];
    95: reg_0375 <= imem06_in[75:72];
    endcase
  end

  // REG#376の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0376 <= imem03_in[91:88];
    28: reg_0376 <= imem03_in[91:88];
    70: reg_0376 <= imem03_in[91:88];
    endcase
  end

  // REG#377の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0377 <= imem03_in[75:72];
    28: reg_0377 <= imem03_in[75:72];
    70: reg_0377 <= imem03_in[75:72];
    endcase
  end

  // REG#378の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0378 <= op1_06_out;
    27: reg_0378 <= op1_06_out;
    29: reg_0378 <= op1_06_out;
    31: reg_0378 <= op1_06_out;
    33: reg_0378 <= op1_06_out;
    35: reg_0378 <= op1_06_out;
    37: reg_0378 <= op1_06_out;
    39: reg_0378 <= op1_06_out;
    41: reg_0378 <= op1_06_out;
    43: reg_0378 <= op1_06_out;
    45: reg_0378 <= op1_06_out;
    47: reg_0378 <= op1_06_out;
    49: reg_0378 <= op1_06_out;
    51: reg_0378 <= op1_06_out;
    53: reg_0378 <= op1_06_out;
    55: reg_0378 <= op1_06_out;
    57: reg_0378 <= op1_06_out;
    59: reg_0378 <= op1_06_out;
    61: reg_0378 <= op1_06_out;
    63: reg_0378 <= op1_06_out;
    65: reg_0378 <= op1_06_out;
    67: reg_0378 <= op1_06_out;
    69: reg_0378 <= op1_06_out;
    71: reg_0378 <= op1_06_out;
    73: reg_0378 <= op1_06_out;
    75: reg_0378 <= op1_06_out;
    77: reg_0378 <= op1_06_out;
    79: reg_0378 <= op1_06_out;
    81: reg_0378 <= op1_06_out;
    83: reg_0378 <= op1_06_out;
    85: reg_0378 <= op1_06_out;
    87: reg_0378 <= op1_06_out;
    89: reg_0378 <= op1_06_out;
    91: reg_0378 <= op1_06_out;
    93: reg_0378 <= op1_06_out;
    95: reg_0378 <= op1_06_out;
    97: reg_0378 <= op1_06_out;
    endcase
  end

  // REG#379の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0379 <= imem06_in[15:12];
    28: reg_0379 <= op2_01_out;
    41: reg_0379 <= op2_01_out;
    84: reg_0379 <= imem06_in[15:12];
    86: reg_0379 <= imem06_in[15:12];
    94: reg_0379 <= op2_01_out;
    endcase
  end

  // REG#380の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0380 <= imem06_in[115:112];
    29: reg_0380 <= imem06_in[115:112];
    58: reg_0380 <= imem06_in[115:112];
    86: reg_0380 <= imem06_in[115:112];
    endcase
  end

  // REG#381の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0381 <= imem06_in[27:24];
    29: reg_0381 <= imem06_in[27:24];
    56: reg_0381 <= imem02_in[43:40];
    58: reg_0381 <= imem02_in[43:40];
    60: reg_0381 <= imem02_in[127:124];
    62: reg_0381 <= imem02_in[127:124];
    65: reg_0381 <= imem04_in[31:28];
    67: reg_0381 <= imem04_in[47:44];
    69: reg_0381 <= imem04_in[47:44];
    71: reg_0381 <= imem06_in[27:24];
    85: reg_0381 <= imem02_in[43:40];
    endcase
  end

  // REG#382の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0382 <= imem06_in[79:76];
    29: reg_0382 <= imem06_in[79:76];
    58: reg_0382 <= imem06_in[79:76];
    86: reg_0382 <= imem06_in[79:76];
    endcase
  end

  // REG#383の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0383 <= imem06_in[83:80];
    29: reg_0383 <= imem06_in[83:80];
    54: reg_0383 <= imem00_in[119:116];
    57: reg_0383 <= imem03_in[23:20];
    59: reg_0383 <= imem03_in[23:20];
    61: reg_0383 <= imem00_in[119:116];
    63: reg_0383 <= imem06_in[119:116];
    65: reg_0383 <= imem02_in[35:32];
    67: reg_0383 <= imem06_in[83:80];
    69: reg_0383 <= imem00_in[119:116];
    71: reg_0383 <= imem06_in[83:80];
    89: reg_0383 <= imem00_in[119:116];
    91: reg_0383 <= imem02_in[35:32];
    93: reg_0383 <= imem02_in[35:32];
    endcase
  end

  // REG#384の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0384 <= imem03_in[11:8];
    29: reg_0384 <= imem06_in[123:120];
    54: reg_0384 <= imem00_in[27:24];
    57: reg_0384 <= imem06_in[123:120];
    endcase
  end

  // REG#385の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0385 <= imem03_in[67:64];
    29: reg_0385 <= imem06_in[3:0];
    54: reg_0385 <= imem06_in[3:0];
    56: reg_0385 <= imem03_in[111:108];
    58: reg_0385 <= imem03_in[111:108];
    60: reg_0385 <= imem03_in[67:64];
    62: reg_0385 <= imem03_in[111:108];
    64: reg_0385 <= imem06_in[3:0];
    66: reg_0385 <= imem03_in[67:64];
    68: reg_0385 <= imem03_in[111:108];
    70: reg_0385 <= imem03_in[111:108];
    endcase
  end

  // REG#386の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0386 <= imem06_in[59:56];
    29: reg_0386 <= imem06_in[59:56];
    59: reg_0386 <= imem00_in[23:20];
    61: reg_0386 <= imem06_in[59:56];
    72: reg_0386 <= imem04_in[63:60];
    74: reg_0386 <= imem04_in[63:60];
    76: reg_0386 <= imem00_in[23:20];
    79: reg_0386 <= imem06_in[59:56];
    81: reg_0386 <= imem00_in[23:20];
    83: reg_0386 <= imem00_in[23:20];
    85: reg_0386 <= imem00_in[23:20];
    87: reg_0386 <= imem07_in[119:116];
    89: reg_0386 <= imem04_in[63:60];
    91: reg_0386 <= imem00_in[23:20];
    endcase
  end

  // REG#387の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0387 <= imem03_in[15:12];
    29: reg_0387 <= imem06_in[11:8];
    56: reg_0387 <= imem06_in[11:8];
    60: reg_0387 <= imem06_in[11:8];
    63: reg_0387 <= imem03_in[15:12];
    65: reg_0387 <= imem06_in[11:8];
    67: reg_0387 <= imem04_in[123:120];
    69: reg_0387 <= imem02_in[107:104];
    71: reg_0387 <= imem04_in[123:120];
    73: reg_0387 <= imem06_in[11:8];
    75: reg_0387 <= imem01_in[7:4];
    77: reg_0387 <= imem02_in[107:104];
    79: reg_0387 <= imem04_in[123:120];
    81: reg_0387 <= imem01_in[7:4];
    83: reg_0387 <= imem01_in[7:4];
    85: reg_0387 <= imem05_in[111:108];
    87: reg_0387 <= imem04_in[123:120];
    89: reg_0387 <= imem01_in[7:4];
    91: reg_0387 <= imem03_in[15:12];
    93: reg_0387 <= imem04_in[71:68];
    95: reg_0387 <= imem04_in[123:120];
    97: reg_0387 <= imem04_in[123:120];
    endcase
  end

  // REG#388の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0388 <= imem03_in[47:44];
    29: reg_0388 <= imem06_in[99:96];
    56: reg_0388 <= imem04_in[51:48];
    58: reg_0388 <= imem03_in[47:44];
    60: reg_0388 <= imem03_in[47:44];
    62: reg_0388 <= imem06_in[99:96];
    64: reg_0388 <= imem06_in[99:96];
    65: reg_0388 <= op2_02_out;
    77: reg_0388 <= op2_02_out;
    endcase
  end

  // REG#389の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0389 <= imem03_in[123:120];
    29: reg_0389 <= imem03_in[123:120];
    31: reg_0389 <= imem03_in[123:120];
    52: reg_0389 <= imem02_in[71:68];
    endcase
  end

  // REG#390の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0390 <= imem06_in[103:100];
    29: reg_0390 <= imem06_in[103:100];
    56: reg_0390 <= imem06_in[103:100];
    60: reg_0390 <= imem04_in[67:64];
    62: reg_0390 <= imem04_in[67:64];
    64: reg_0390 <= imem04_in[67:64];
    67: reg_0390 <= imem05_in[75:72];
    70: reg_0390 <= imem06_in[103:100];
    73: reg_0390 <= imem04_in[67:64];
    75: reg_0390 <= imem05_in[75:72];
    77: reg_0390 <= imem04_in[67:64];
    79: reg_0390 <= imem04_in[67:64];
    81: reg_0390 <= imem06_in[103:100];
    83: reg_0390 <= imem04_in[67:64];
    endcase
  end

  // REG#391の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0391 <= imem03_in[19:16];
    29: reg_0391 <= imem06_in[55:52];
    57: reg_0391 <= imem06_in[55:52];
    endcase
  end

  // REG#392の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0392 <= imem06_in[43:40];
    29: reg_0392 <= imem06_in[43:40];
    58: reg_0392 <= imem06_in[43:40];
    87: reg_0392 <= imem01_in[27:24];
    89: reg_0392 <= imem06_in[43:40];
    endcase
  end

  // REG#393の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0393 <= imem03_in[103:100];
    29: reg_0393 <= imem06_in[63:60];
    57: reg_0393 <= imem06_in[63:60];
    endcase
  end

  // REG#394の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0394 <= imem03_in[3:0];
    29: reg_0394 <= imem03_in[3:0];
    31: reg_0394 <= imem03_in[3:0];
    50: reg_0394 <= imem03_in[3:0];
    52: reg_0394 <= imem02_in[63:60];
    endcase
  end

  // REG#395の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0395 <= imem03_in[7:4];
    29: reg_0395 <= imem06_in[31:28];
    58: reg_0395 <= imem06_in[31:28];
    83: reg_0395 <= imem04_in[27:24];
    endcase
  end

  // REG#396の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0396 <= imem03_in[111:108];
    29: reg_0396 <= imem03_in[111:108];
    31: reg_0396 <= imem03_in[111:108];
    55: reg_0396 <= imem03_in[111:108];
    87: reg_0396 <= imem03_in[111:108];
    90: reg_0396 <= imem03_in[111:108];
    endcase
  end

  // REG#397の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0397 <= imem03_in[99:96];
    29: reg_0397 <= imem03_in[99:96];
    31: reg_0397 <= imem03_in[99:96];
    54: reg_0397 <= imem03_in[99:96];
    56: reg_0397 <= imem03_in[99:96];
    58: reg_0397 <= imem03_in[23:20];
    60: reg_0397 <= imem04_in[95:92];
    62: reg_0397 <= imem03_in[23:20];
    64: reg_0397 <= imem03_in[99:96];
    66: reg_0397 <= imem03_in[23:20];
    68: reg_0397 <= imem00_in[47:44];
    70: reg_0397 <= imem03_in[23:20];
    endcase
  end

  // REG#398の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0398 <= imem03_in[87:84];
    29: reg_0398 <= imem03_in[87:84];
    31: reg_0398 <= imem03_in[87:84];
    54: reg_0398 <= imem03_in[87:84];
    56: reg_0398 <= imem04_in[83:80];
    58: reg_0398 <= imem04_in[83:80];
    60: reg_0398 <= imem03_in[87:84];
    62: reg_0398 <= imem04_in[95:92];
    64: reg_0398 <= imem04_in[83:80];
    67: reg_0398 <= imem03_in[87:84];
    69: reg_0398 <= imem03_in[87:84];
    71: reg_0398 <= imem04_in[95:92];
    73: reg_0398 <= imem04_in[95:92];
    75: reg_0398 <= imem01_in[43:40];
    77: reg_0398 <= imem01_in[43:40];
    79: reg_0398 <= imem03_in[103:100];
    81: reg_0398 <= imem03_in[103:100];
    83: reg_0398 <= imem01_in[43:40];
    85: reg_0398 <= imem03_in[87:84];
    87: reg_0398 <= imem04_in[83:80];
    89: reg_0398 <= imem04_in[95:92];
    91: reg_0398 <= imem03_in[87:84];
    93: reg_0398 <= imem03_in[87:84];
    95: reg_0398 <= imem01_in[43:40];
    endcase
  end

  // REG#399の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0399 <= imem06_in[91:88];
    29: reg_0399 <= imem06_in[91:88];
    59: reg_0399 <= imem03_in[35:32];
    61: reg_0399 <= imem06_in[91:88];
    72: reg_0399 <= imem06_in[91:88];
    74: reg_0399 <= imem06_in[91:88];
    76: reg_0399 <= imem03_in[35:32];
    78: reg_0399 <= imem06_in[91:88];
    80: reg_0399 <= imem03_in[35:32];
    82: reg_0399 <= imem00_in[47:44];
    84: reg_0399 <= imem06_in[91:88];
    86: reg_0399 <= imem03_in[35:32];
    88: reg_0399 <= imem00_in[39:36];
    90: reg_0399 <= imem06_in[91:88];
    92: reg_0399 <= imem01_in[119:116];
    endcase
  end

  // REG#400の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0400 <= op1_07_out;
    28: reg_0400 <= op1_07_out;
    30: reg_0400 <= op1_07_out;
    32: reg_0400 <= op1_07_out;
    34: reg_0400 <= op1_07_out;
    36: reg_0400 <= op1_07_out;
    38: reg_0400 <= op1_07_out;
    40: reg_0400 <= op1_07_out;
    42: reg_0400 <= op1_07_out;
    44: reg_0400 <= op1_07_out;
    46: reg_0400 <= op1_07_out;
    48: reg_0400 <= op1_07_out;
    50: reg_0400 <= op1_07_out;
    52: reg_0400 <= op1_07_out;
    54: reg_0400 <= op1_07_out;
    56: reg_0400 <= op1_07_out;
    58: reg_0400 <= op1_07_out;
    60: reg_0400 <= op1_07_out;
    62: reg_0400 <= op1_07_out;
    64: reg_0400 <= op1_07_out;
    66: reg_0400 <= op1_07_out;
    68: reg_0400 <= op1_07_out;
    70: reg_0400 <= op1_07_out;
    72: reg_0400 <= op1_07_out;
    74: reg_0400 <= op1_07_out;
    76: reg_0400 <= op1_07_out;
    78: reg_0400 <= op1_07_out;
    80: reg_0400 <= op1_07_out;
    82: reg_0400 <= op1_07_out;
    84: reg_0400 <= op1_07_out;
    86: reg_0400 <= op1_07_out;
    88: reg_0400 <= op1_07_out;
    90: reg_0400 <= op1_07_out;
    92: reg_0400 <= op1_07_out;
    94: reg_0400 <= op1_07_out;
    96: reg_0400 <= op1_07_out;
    endcase
  end

  // REG#401の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0401 <= imem06_in[123:120];
    30: reg_0401 <= imem04_in[79:76];
    32: reg_0401 <= imem04_in[79:76];
    34: reg_0401 <= imem04_in[79:76];
    36: reg_0401 <= imem06_in[123:120];
    38: reg_0401 <= imem04_in[79:76];
    40: reg_0401 <= imem06_in[123:120];
    42: reg_0401 <= imem04_in[79:76];
    endcase
  end

  // REG#402の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0402 <= imem06_in[3:0];
    30: reg_0402 <= imem05_in[3:0];
    32: reg_0402 <= imem06_in[3:0];
    38: reg_0402 <= imem06_in[3:0];
    39: reg_0402 <= op2_02_out;
    79: reg_0402 <= imem06_in[3:0];
    81: reg_0402 <= imem05_in[3:0];
    82: reg_0402 <= op2_02_out;
    90: reg_0402 <= op2_02_out;
    endcase
  end

  // REG#403の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0403 <= imem06_in[87:84];
    30: reg_0403 <= imem05_in[35:32];
    32: reg_0403 <= imem05_in[35:32];
    34: reg_0403 <= imem05_in[115:112];
    36: reg_0403 <= imem06_in[87:84];
    39: reg_0403 <= imem06_in[87:84];
    55: reg_0403 <= imem07_in[7:4];
    57: reg_0403 <= imem05_in[115:112];
    59: reg_0403 <= imem07_in[7:4];
    61: reg_0403 <= imem05_in[115:112];
    63: reg_0403 <= imem05_in[35:32];
    65: reg_0403 <= imem06_in[87:84];
    67: reg_0403 <= imem06_in[87:84];
    69: reg_0403 <= imem05_in[115:112];
    71: reg_0403 <= imem06_in[87:84];
    89: reg_0403 <= imem06_in[87:84];
    endcase
  end

  // REG#404の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0404 <= imem06_in[95:92];
    30: reg_0404 <= imem06_in[71:68];
    32: reg_0404 <= imem06_in[71:68];
    38: reg_0404 <= imem01_in[67:64];
    40: reg_0404 <= imem01_in[67:64];
    42: reg_0404 <= imem03_in[119:116];
    44: reg_0404 <= imem01_in[67:64];
    46: reg_0404 <= imem06_in[95:92];
    48: reg_0404 <= imem06_in[95:92];
    50: reg_0404 <= imem05_in[95:92];
    65: reg_0404 <= imem01_in[67:64];
    67: reg_0404 <= imem06_in[95:92];
    69: reg_0404 <= imem06_in[71:68];
    71: reg_0404 <= imem01_in[67:64];
    73: reg_0404 <= imem01_in[67:64];
    75: reg_0404 <= imem05_in[95:92];
    77: reg_0404 <= imem03_in[119:116];
    79: reg_0404 <= imem05_in[95:92];
    86: reg_0404 <= imem01_in[67:64];
    88: reg_0404 <= imem06_in[71:68];
    90: reg_0404 <= imem05_in[95:92];
    92: reg_0404 <= imem03_in[119:116];
    94: reg_0404 <= imem05_in[95:92];
    endcase
  end

  // REG#405の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0405 <= imem06_in[55:52];
    30: reg_0405 <= imem07_in[47:44];
    32: reg_0405 <= imem06_in[55:52];
    38: reg_0405 <= imem07_in[47:44];
    41: reg_0405 <= imem06_in[55:52];
    43: reg_0405 <= imem03_in[7:4];
    45: reg_0405 <= imem03_in[7:4];
    47: reg_0405 <= imem06_in[55:52];
    49: reg_0405 <= imem03_in[7:4];
    51: reg_0405 <= imem06_in[55:52];
    53: reg_0405 <= imem03_in[7:4];
    57: reg_0405 <= imem03_in[51:48];
    59: reg_0405 <= imem03_in[7:4];
    61: reg_0405 <= imem06_in[55:52];
    71: reg_0405 <= imem03_in[51:48];
    73: reg_0405 <= imem03_in[7:4];
    75: reg_0405 <= imem07_in[47:44];
    79: reg_0405 <= imem06_in[55:52];
    81: reg_0405 <= imem03_in[7:4];
    83: reg_0405 <= imem04_in[19:16];
    endcase
  end

  // REG#406の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0406 <= imem06_in[107:104];
    30: reg_0406 <= imem07_in[55:52];
    32: reg_0406 <= imem07_in[63:60];
    34: reg_0406 <= imem01_in[51:48];
    36: reg_0406 <= imem06_in[107:104];
    41: reg_0406 <= imem07_in[55:52];
    43: reg_0406 <= imem07_in[63:60];
    endcase
  end

  // REG#407の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0407 <= imem06_in[47:44];
    30: reg_0407 <= imem00_in[79:76];
    32: reg_0407 <= imem00_in[79:76];
    34: reg_0407 <= imem00_in[79:76];
    36: reg_0407 <= imem06_in[47:44];
    39: reg_0407 <= imem06_in[47:44];
    57: reg_0407 <= imem00_in[79:76];
    59: reg_0407 <= imem04_in[15:12];
    90: reg_0407 <= imem06_in[47:44];
    92: reg_0407 <= imem04_in[15:12];
    94: reg_0407 <= imem06_in[47:44];
    96: reg_0407 <= imem06_in[47:44];
    endcase
  end

  // REG#408の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0408 <= imem06_in[35:32];
    30: reg_0408 <= imem02_in[35:32];
    32: reg_0408 <= imem00_in[55:52];
    34: reg_0408 <= imem02_in[35:32];
    36: reg_0408 <= imem06_in[35:32];
    41: reg_0408 <= imem00_in[55:52];
    43: reg_0408 <= imem03_in[115:112];
    45: reg_0408 <= imem00_in[55:52];
    47: reg_0408 <= imem00_in[55:52];
    49: reg_0408 <= imem02_in[35:32];
    51: reg_0408 <= imem06_in[35:32];
    53: reg_0408 <= imem02_in[35:32];
    55: reg_0408 <= imem06_in[35:32];
    57: reg_0408 <= imem02_in[35:32];
    59: reg_0408 <= imem06_in[35:32];
    61: reg_0408 <= imem06_in[35:32];
    69: reg_0408 <= imem02_in[35:32];
    71: reg_0408 <= imem00_in[55:52];
    73: reg_0408 <= imem07_in[35:32];
    75: reg_0408 <= imem03_in[115:112];
    77: reg_0408 <= imem00_in[55:52];
    79: reg_0408 <= imem03_in[115:112];
    81: reg_0408 <= imem00_in[55:52];
    83: reg_0408 <= imem02_in[35:32];
    85: reg_0408 <= imem02_in[35:32];
    endcase
  end

  // REG#409の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0409 <= imem06_in[63:60];
    30: reg_0409 <= imem03_in[99:96];
    32: reg_0409 <= imem03_in[99:96];
    34: reg_0409 <= imem01_in[79:76];
    36: reg_0409 <= imem01_in[79:76];
    38: reg_0409 <= imem03_in[99:96];
    40: reg_0409 <= imem06_in[63:60];
    42: reg_0409 <= imem03_in[99:96];
    44: reg_0409 <= imem03_in[99:96];
    46: reg_0409 <= imem06_in[63:60];
    48: reg_0409 <= imem01_in[79:76];
    50: reg_0409 <= imem03_in[99:96];
    52: reg_0409 <= imem06_in[63:60];
    54: reg_0409 <= imem00_in[3:0];
    57: reg_0409 <= imem01_in[79:76];
    59: reg_0409 <= imem04_in[55:52];
    95: reg_0409 <= imem01_in[79:76];
    endcase
  end

  // REG#410の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0410 <= op1_08_out;
    30: reg_0410 <= op1_08_out;
    32: reg_0410 <= op1_08_out;
    34: reg_0410 <= op1_08_out;
    36: reg_0410 <= op1_08_out;
    38: reg_0410 <= op1_08_out;
    40: reg_0410 <= op1_08_out;
    42: reg_0410 <= op1_08_out;
    44: reg_0410 <= op1_08_out;
    46: reg_0410 <= op1_08_out;
    48: reg_0410 <= op1_08_out;
    50: reg_0410 <= op1_08_out;
    52: reg_0410 <= op1_08_out;
    54: reg_0410 <= op1_08_out;
    56: reg_0410 <= op1_08_out;
    58: reg_0410 <= op1_08_out;
    60: reg_0410 <= op1_08_out;
    62: reg_0410 <= op1_08_out;
    64: reg_0410 <= op1_08_out;
    66: reg_0410 <= op1_08_out;
    68: reg_0410 <= op1_08_out;
    70: reg_0410 <= op1_08_out;
    72: reg_0410 <= op1_08_out;
    74: reg_0410 <= op1_08_out;
    76: reg_0410 <= op1_08_out;
    78: reg_0410 <= op1_08_out;
    80: reg_0410 <= op1_08_out;
    82: reg_0410 <= op1_08_out;
    84: reg_0410 <= op1_08_out;
    86: reg_0410 <= op1_08_out;
    88: reg_0410 <= op1_08_out;
    90: reg_0410 <= op1_08_out;
    92: reg_0410 <= op1_08_out;
    94: reg_0410 <= op1_08_out;
    96: reg_0410 <= op1_08_out;
    endcase
  end

  // REG#411の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0411 <= op1_09_out;
    31: reg_0411 <= op1_09_out;
    33: reg_0411 <= op1_09_out;
    35: reg_0411 <= op1_09_out;
    37: reg_0411 <= op1_09_out;
    39: reg_0411 <= op1_09_out;
    41: reg_0411 <= op1_09_out;
    43: reg_0411 <= op1_09_out;
    45: reg_0411 <= op1_09_out;
    47: reg_0411 <= op1_09_out;
    49: reg_0411 <= op1_09_out;
    51: reg_0411 <= op1_09_out;
    53: reg_0411 <= op1_09_out;
    55: reg_0411 <= op1_09_out;
    57: reg_0411 <= op1_09_out;
    59: reg_0411 <= op1_09_out;
    61: reg_0411 <= op1_09_out;
    63: reg_0411 <= op1_09_out;
    65: reg_0411 <= op1_09_out;
    67: reg_0411 <= op1_09_out;
    69: reg_0411 <= op1_09_out;
    71: reg_0411 <= op1_09_out;
    73: reg_0411 <= op1_09_out;
    75: reg_0411 <= op1_09_out;
    77: reg_0411 <= op1_09_out;
    79: reg_0411 <= op1_09_out;
    81: reg_0411 <= op1_09_out;
    83: reg_0411 <= op1_09_out;
    85: reg_0411 <= op1_09_out;
    87: reg_0411 <= op1_09_out;
    89: reg_0411 <= op1_09_out;
    91: reg_0411 <= op1_09_out;
    93: reg_0411 <= op1_09_out;
    95: reg_0411 <= op1_09_out;
    97: reg_0411 <= op1_09_out;
    endcase
  end

  // REG#412の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0412 <= op1_10_out;
    33: reg_0412 <= op1_10_out;
    35: reg_0412 <= op1_10_out;
    37: reg_0412 <= op1_10_out;
    39: reg_0412 <= op1_10_out;
    41: reg_0412 <= op1_10_out;
    43: reg_0412 <= op1_10_out;
    45: reg_0412 <= op1_10_out;
    47: reg_0412 <= op1_10_out;
    49: reg_0412 <= op1_10_out;
    51: reg_0412 <= op1_10_out;
    53: reg_0412 <= op1_10_out;
    55: reg_0412 <= op1_10_out;
    57: reg_0412 <= op1_10_out;
    59: reg_0412 <= op1_10_out;
    61: reg_0412 <= op1_10_out;
    63: reg_0412 <= op1_10_out;
    65: reg_0412 <= op1_10_out;
    67: reg_0412 <= op1_10_out;
    69: reg_0412 <= op1_10_out;
    71: reg_0412 <= op1_10_out;
    73: reg_0412 <= op1_10_out;
    75: reg_0412 <= op1_10_out;
    77: reg_0412 <= op1_10_out;
    79: reg_0412 <= op1_10_out;
    81: reg_0412 <= op1_10_out;
    83: reg_0412 <= op1_10_out;
    85: reg_0412 <= op1_10_out;
    87: reg_0412 <= op1_10_out;
    89: reg_0412 <= op1_10_out;
    91: reg_0412 <= op1_10_out;
    93: reg_0412 <= op1_10_out;
    95: reg_0412 <= op1_10_out;
    97: reg_0412 <= op1_10_out;
    endcase
  end

  // REG#413の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0413 <= op1_11_out;
    34: reg_0413 <= op1_11_out;
    36: reg_0413 <= op1_11_out;
    38: reg_0413 <= op1_11_out;
    40: reg_0413 <= op1_11_out;
    42: reg_0413 <= op1_11_out;
    44: reg_0413 <= op1_11_out;
    46: reg_0413 <= op1_11_out;
    48: reg_0413 <= op1_11_out;
    50: reg_0413 <= op1_11_out;
    52: reg_0413 <= op1_11_out;
    54: reg_0413 <= op1_11_out;
    56: reg_0413 <= op1_11_out;
    58: reg_0413 <= op1_11_out;
    60: reg_0413 <= op1_11_out;
    62: reg_0413 <= op1_11_out;
    64: reg_0413 <= op1_11_out;
    66: reg_0413 <= op1_11_out;
    68: reg_0413 <= op1_11_out;
    70: reg_0413 <= op1_11_out;
    72: reg_0413 <= op1_11_out;
    74: reg_0413 <= op1_11_out;
    76: reg_0413 <= op1_11_out;
    78: reg_0413 <= op1_11_out;
    80: reg_0413 <= op1_11_out;
    82: reg_0413 <= op1_11_out;
    84: reg_0413 <= op1_11_out;
    86: reg_0413 <= op1_11_out;
    89: reg_0413 <= op1_11_out;
    91: reg_0413 <= op1_11_out;
    93: reg_0413 <= op1_11_out;
    95: reg_0413 <= op1_11_out;
    endcase
  end

  // REG#414の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0414 <= op1_12_out;
    34: reg_0414 <= op1_12_out;
    36: reg_0414 <= op1_12_out;
    39: reg_0414 <= op1_12_out;
    41: reg_0414 <= op1_12_out;
    43: reg_0414 <= op1_12_out;
    45: reg_0414 <= op1_12_out;
    47: reg_0414 <= op1_12_out;
    49: reg_0414 <= op1_12_out;
    52: reg_0414 <= op1_12_out;
    54: reg_0414 <= op1_12_out;
    56: reg_0414 <= op1_12_out;
    59: reg_0414 <= op1_12_out;
    61: reg_0414 <= op1_12_out;
    63: reg_0414 <= op1_12_out;
    65: reg_0414 <= op1_12_out;
    67: reg_0414 <= op1_12_out;
    69: reg_0414 <= op1_12_out;
    71: reg_0414 <= op1_12_out;
    73: reg_0414 <= op1_12_out;
    76: reg_0414 <= op1_12_out;
    78: reg_0414 <= op1_12_out;
    80: reg_0414 <= op1_12_out;
    83: reg_0414 <= op1_12_out;
    85: reg_0414 <= op1_12_out;
    88: reg_0414 <= op1_12_out;
    91: reg_0414 <= op1_12_out;
    93: reg_0414 <= op1_12_out;
    95: reg_0414 <= op1_12_out;
    endcase
  end

  // REG#415の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0415 <= op1_13_out;
    34: reg_0415 <= op1_13_out;
    37: reg_0415 <= op1_13_out;
    39: reg_0415 <= op1_13_out;
    41: reg_0415 <= op1_13_out;
    43: reg_0415 <= op1_13_out;
    45: reg_0415 <= op1_13_out;
    48: reg_0415 <= op1_13_out;
    51: reg_0415 <= op1_13_out;
    53: reg_0415 <= op1_13_out;
    55: reg_0415 <= op1_13_out;
    58: reg_0415 <= op1_13_out;
    61: reg_0415 <= op1_13_out;
    63: reg_0415 <= op1_13_out;
    66: reg_0415 <= op1_13_out;
    69: reg_0415 <= op1_13_out;
    71: reg_0415 <= op1_13_out;
    73: reg_0415 <= op1_13_out;
    76: reg_0415 <= op1_13_out;
    78: reg_0415 <= op1_13_out;
    81: reg_0415 <= op1_13_out;
    84: reg_0415 <= op1_13_out;
    86: reg_0415 <= op1_13_out;
    90: reg_0415 <= imem07_in[35:32];
    91: reg_0415 <= op1_13_out;
    94: reg_0415 <= op1_13_out;
    96: reg_0415 <= op1_13_out;
    endcase
  end

  // REG#416の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0416 <= op1_14_out;
    35: reg_0416 <= op1_14_out;
    38: reg_0416 <= op1_14_out;
    40: reg_0416 <= op1_14_out;
    42: reg_0416 <= op1_14_out;
    45: reg_0416 <= op1_14_out;
    48: reg_0416 <= op1_14_out;
    51: reg_0416 <= op1_14_out;
    54: reg_0416 <= op1_14_out;
    57: reg_0416 <= op1_14_out;
    60: reg_0416 <= op1_14_out;
    63: reg_0416 <= op1_14_out;
    66: reg_0416 <= op1_14_out;
    69: reg_0416 <= op1_14_out;
    72: reg_0416 <= op1_14_out;
    75: reg_0416 <= op1_14_out;
    77: reg_0416 <= op1_14_out;
    80: reg_0416 <= op1_14_out;
    83: reg_0416 <= op1_14_out;
    86: reg_0416 <= op1_14_out;
    89: reg_0416 <= op1_14_out;
    92: reg_0416 <= op1_14_out;
    94: reg_0416 <= op1_14_out;
    96: reg_0416 <= op1_14_out;
    endcase
  end

  // REG#417の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0417 <= op1_15_out;
    36: reg_0417 <= op1_15_out;
    39: reg_0417 <= op1_15_out;
    42: reg_0417 <= op1_15_out;
    45: reg_0417 <= op1_15_out;
    48: reg_0417 <= op1_15_out;
    51: reg_0417 <= op1_15_out;
    54: reg_0417 <= op1_15_out;
    57: reg_0417 <= op1_15_out;
    60: reg_0417 <= op1_15_out;
    63: reg_0417 <= op1_15_out;
    66: reg_0417 <= op1_15_out;
    69: reg_0417 <= op1_15_out;
    72: reg_0417 <= op1_15_out;
    75: reg_0417 <= op1_15_out;
    77: reg_0417 <= op1_15_out;
    80: reg_0417 <= op1_15_out;
    83: reg_0417 <= op1_15_out;
    86: reg_0417 <= op1_15_out;
    89: reg_0417 <= op1_15_out;
    92: reg_0417 <= op1_15_out;
    95: reg_0417 <= op1_15_out;
    endcase
  end

  // REG#418の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0418 <= imem07_in[51:48];
    38: reg_0418 <= imem07_in[51:48];
    41: reg_0418 <= imem02_in[127:124];
    43: reg_0418 <= imem02_in[127:124];
    45: reg_0418 <= imem02_in[127:124];
    61: reg_0418 <= imem04_in[51:48];
    63: reg_0418 <= imem04_in[51:48];
    65: reg_0418 <= imem04_in[51:48];
    67: reg_0418 <= imem04_in[51:48];
    69: reg_0418 <= imem04_in[51:48];
    72: reg_0418 <= imem02_in[127:124];
    84: reg_0418 <= imem02_in[127:124];
    endcase
  end

  // REG#419の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0419 <= imem07_in[55:52];
    39: reg_0419 <= imem07_in[67:64];
    41: reg_0419 <= imem05_in[43:40];
    43: reg_0419 <= imem07_in[67:64];
    endcase
  end

  // REG#420の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0420 <= imem07_in[111:108];
    39: reg_0420 <= imem07_in[99:96];
    41: reg_0420 <= imem07_in[111:108];
    43: reg_0420 <= imem07_in[99:96];
    endcase
  end

  // REG#421の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0421 <= imem07_in[39:36];
    39: reg_0421 <= imem07_in[39:36];
    41: reg_0421 <= imem07_in[39:36];
    43: reg_0421 <= imem07_in[39:36];
    97: reg_0421 <= imem07_in[39:36];
    endcase
  end

  // REG#422の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0422 <= imem07_in[31:28];
    41: reg_0422 <= imem05_in[83:80];
    43: reg_0422 <= imem07_in[31:28];
    endcase
  end

  // REG#423の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0423 <= imem07_in[59:56];
    42: reg_0423 <= imem05_in[63:60];
    44: reg_0423 <= imem04_in[83:80];
    46: reg_0423 <= imem04_in[83:80];
    49: reg_0423 <= imem00_in[71:68];
    52: reg_0423 <= imem02_in[59:56];
    endcase
  end

  // REG#424の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0424 <= imem07_in[11:8];
    42: reg_0424 <= imem07_in[119:116];
    44: reg_0424 <= imem05_in[27:24];
    46: reg_0424 <= imem05_in[27:24];
    48: reg_0424 <= imem07_in[11:8];
    50: reg_0424 <= imem07_in[11:8];
    52: reg_0424 <= imem02_in[35:32];
    endcase
  end

  // REG#425の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0425 <= imem07_in[3:0];
    42: reg_0425 <= imem07_in[3:0];
    45: reg_0425 <= imem07_in[3:0];
    47: reg_0425 <= imem00_in[75:72];
    49: reg_0425 <= imem00_in[75:72];
    52: reg_0425 <= imem02_in[75:72];
    endcase
  end

  // REG#426の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0426 <= imem07_in[43:40];
    43: reg_0426 <= imem07_in[43:40];
    97: reg_0426 <= imem07_in[43:40];
    endcase
  end

  // REG#427の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0427 <= imem07_in[103:100];
    43: reg_0427 <= imem07_in[103:100];
    endcase
  end

  // REG#428の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0428 <= imem07_in[71:68];
    43: reg_0428 <= imem07_in[71:68];
    endcase
  end

  // REG#429の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0429 <= imem07_in[19:16];
    43: reg_0429 <= imem04_in[67:64];
    45: reg_0429 <= imem04_in[67:64];
    47: reg_0429 <= imem04_in[67:64];
    49: reg_0429 <= imem04_in[67:64];
    57: reg_0429 <= imem03_in[95:92];
    59: reg_0429 <= imem03_in[95:92];
    61: reg_0429 <= imem07_in[19:16];
    63: reg_0429 <= imem07_in[3:0];
    65: reg_0429 <= imem02_in[103:100];
    68: reg_0429 <= imem02_in[103:100];
    71: reg_0429 <= imem04_in[67:64];
    73: reg_0429 <= imem07_in[3:0];
    75: reg_0429 <= imem07_in[19:16];
    78: reg_0429 <= imem02_in[103:100];
    80: reg_0429 <= imem07_in[19:16];
    82: reg_0429 <= imem07_in[19:16];
    endcase
  end

  // REG#430の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0430 <= imem07_in[15:12];
    43: reg_0430 <= imem04_in[79:76];
    45: reg_0430 <= imem04_in[79:76];
    47: reg_0430 <= imem03_in[127:124];
    49: reg_0430 <= imem03_in[127:124];
    51: reg_0430 <= imem03_in[127:124];
    53: reg_0430 <= imem03_in[127:124];
    55: reg_0430 <= imem07_in[15:12];
    57: reg_0430 <= imem04_in[79:76];
    59: reg_0430 <= imem07_in[15:12];
    61: reg_0430 <= imem03_in[127:124];
    63: reg_0430 <= imem04_in[79:76];
    65: reg_0430 <= imem04_in[79:76];
    67: reg_0430 <= imem03_in[127:124];
    69: reg_0430 <= imem05_in[51:48];
    71: reg_0430 <= imem05_in[51:48];
    73: reg_0430 <= imem04_in[79:76];
    75: reg_0430 <= imem04_in[79:76];
    77: reg_0430 <= imem04_in[79:76];
    79: reg_0430 <= imem04_in[79:76];
    81: reg_0430 <= imem04_in[79:76];
    83: reg_0430 <= imem04_in[79:76];
    endcase
  end

  // REG#431の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0431 <= imem07_in[127:124];
    43: reg_0431 <= imem07_in[127:124];
    endcase
  end

  // REG#432の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0432 <= imem07_in[23:20];
    43: reg_0432 <= imem05_in[27:24];
    45: reg_0432 <= imem06_in[7:4];
    47: reg_0432 <= imem05_in[27:24];
    49: reg_0432 <= imem05_in[27:24];
    51: reg_0432 <= imem07_in[23:20];
    53: reg_0432 <= imem05_in[27:24];
    55: reg_0432 <= imem01_in[71:68];
    57: reg_0432 <= imem07_in[23:20];
    59: reg_0432 <= imem04_in[11:8];
    endcase
  end

  // REG#433の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0433 <= imem07_in[35:32];
    43: reg_0433 <= imem07_in[35:32];
    endcase
  end

  // REG#434の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0434 <= imem07_in[75:72];
    44: reg_0434 <= imem05_in[119:116];
    46: reg_0434 <= imem03_in[87:84];
    48: reg_0434 <= imem03_in[87:84];
    50: reg_0434 <= imem03_in[87:84];
    52: reg_0434 <= imem03_in[87:84];
    55: reg_0434 <= imem03_in[87:84];
    88: reg_0434 <= imem00_in[75:72];
    90: reg_0434 <= imem00_in[75:72];
    92: reg_0434 <= imem07_in[75:72];
    94: reg_0434 <= imem05_in[119:116];
    endcase
  end

  // REG#435の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0435 <= imem07_in[123:120];
    44: reg_0435 <= imem07_in[51:48];
    46: reg_0435 <= imem05_in[71:68];
    48: reg_0435 <= imem05_in[71:68];
    50: reg_0435 <= imem05_in[71:68];
    67: reg_0435 <= imem05_in[71:68];
    72: reg_0435 <= imem07_in[123:120];
    74: reg_0435 <= imem07_in[51:48];
    76: reg_0435 <= imem07_in[123:120];
    78: reg_0435 <= imem07_in[51:48];
    81: reg_0435 <= imem07_in[51:48];
    83: reg_0435 <= imem05_in[71:68];
    85: reg_0435 <= imem07_in[51:48];
    87: reg_0435 <= imem07_in[51:48];
    89: reg_0435 <= imem07_in[51:48];
    91: reg_0435 <= imem05_in[71:68];
    93: reg_0435 <= imem07_in[51:48];
    96: reg_0435 <= imem05_in[71:68];
    endcase
  end

  // REG#436の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0436 <= imem07_in[27:24];
    44: reg_0436 <= imem01_in[19:16];
    46: reg_0436 <= imem05_in[79:76];
    48: reg_0436 <= imem05_in[79:76];
    50: reg_0436 <= imem05_in[79:76];
    66: reg_0436 <= imem05_in[79:76];
    76: reg_0436 <= imem07_in[91:88];
    78: reg_0436 <= imem01_in[19:16];
    80: reg_0436 <= imem07_in[91:88];
    83: reg_0436 <= imem01_in[19:16];
    85: reg_0436 <= imem01_in[19:16];
    87: reg_0436 <= imem05_in[79:76];
    97: reg_0436 <= imem05_in[79:76];
    endcase
  end

  // REG#437の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0437 <= imem07_in[107:104];
    44: reg_0437 <= imem07_in[107:104];
    46: reg_0437 <= imem05_in[95:92];
    48: reg_0437 <= imem05_in[95:92];
    50: reg_0437 <= imem07_in[107:104];
    52: reg_0437 <= imem07_in[107:104];
    55: reg_0437 <= imem05_in[7:4];
    57: reg_0437 <= imem07_in[107:104];
    59: reg_0437 <= imem05_in[95:92];
    61: reg_0437 <= imem05_in[7:4];
    65: reg_0437 <= imem05_in[95:92];
    68: reg_0437 <= imem07_in[107:104];
    70: reg_0437 <= imem07_in[107:104];
    72: reg_0437 <= imem04_in[119:116];
    74: reg_0437 <= imem07_in[107:104];
    77: reg_0437 <= imem05_in[95:92];
    79: reg_0437 <= imem04_in[119:116];
    81: reg_0437 <= imem05_in[7:4];
    83: reg_0437 <= imem05_in[95:92];
    85: reg_0437 <= imem07_in[107:104];
    87: reg_0437 <= imem05_in[95:92];
    96: reg_0437 <= imem05_in[7:4];
    endcase
  end

  // REG#438の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0438 <= imem07_in[115:112];
    44: reg_0438 <= imem01_in[23:20];
    46: reg_0438 <= imem07_in[115:112];
    48: reg_0438 <= imem04_in[83:80];
    50: reg_0438 <= imem05_in[119:116];
    66: reg_0438 <= imem05_in[119:116];
    80: reg_0438 <= imem07_in[115:112];
    84: reg_0438 <= imem07_in[115:112];
    86: reg_0438 <= imem01_in[23:20];
    88: reg_0438 <= imem01_in[15:12];
    90: reg_0438 <= imem04_in[83:80];
    92: reg_0438 <= imem07_in[115:112];
    95: reg_0438 <= imem04_in[83:80];
    endcase
  end

  // REG#439の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0439 <= imem07_in[67:64];
    44: reg_0439 <= imem02_in[111:108];
    46: reg_0439 <= imem02_in[111:108];
    48: reg_0439 <= imem06_in[55:52];
    50: reg_0439 <= imem06_in[55:52];
    52: reg_0439 <= imem07_in[67:64];
    54: reg_0439 <= imem07_in[67:64];
    56: reg_0439 <= imem02_in[111:108];
    58: reg_0439 <= imem06_in[55:52];
    86: reg_0439 <= imem06_in[55:52];
    94: reg_0439 <= imem06_in[55:52];
    96: reg_0439 <= imem06_in[55:52];
    endcase
  end

  // REG#440の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0440 <= imem07_in[87:84];
    44: reg_0440 <= imem07_in[87:84];
    46: reg_0440 <= imem06_in[19:16];
    48: reg_0440 <= imem07_in[87:84];
    50: reg_0440 <= imem07_in[87:84];
    52: reg_0440 <= imem07_in[87:84];
    54: reg_0440 <= imem07_in[87:84];
    56: reg_0440 <= imem07_in[3:0];
    58: reg_0440 <= imem06_in[19:16];
    86: reg_0440 <= imem06_in[19:16];
    endcase
  end

  // REG#441の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0441 <= imem07_in[7:4];
    44: reg_0441 <= imem04_in[67:64];
    46: reg_0441 <= imem04_in[67:64];
    48: reg_0441 <= imem07_in[7:4];
    50: reg_0441 <= imem04_in[67:64];
    52: reg_0441 <= imem02_in[31:28];
    endcase
  end

  // REG#442の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0442 <= imem07_in[95:92];
    44: reg_0442 <= imem07_in[95:92];
    46: reg_0442 <= imem07_in[11:8];
    48: reg_0442 <= imem04_in[19:16];
    50: reg_0442 <= imem04_in[19:16];
    52: reg_0442 <= imem07_in[95:92];
    55: reg_0442 <= imem07_in[11:8];
    57: reg_0442 <= imem04_in[23:20];
    59: reg_0442 <= imem07_in[11:8];
    61: reg_0442 <= imem04_in[19:16];
    63: reg_0442 <= imem07_in[11:8];
    65: reg_0442 <= imem03_in[59:56];
    67: reg_0442 <= imem04_in[19:16];
    69: reg_0442 <= imem07_in[11:8];
    71: reg_0442 <= imem07_in[11:8];
    73: reg_0442 <= imem07_in[11:8];
    75: reg_0442 <= imem07_in[11:8];
    77: reg_0442 <= imem07_in[11:8];
    79: reg_0442 <= imem07_in[95:92];
    endcase
  end

  // REG#443の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0443 <= imem07_in[99:96];
    44: reg_0443 <= imem04_in[87:84];
    46: reg_0443 <= imem07_in[99:96];
    47: reg_0443 <= op1_03_out;
    49: reg_0443 <= op1_03_out;
    52: reg_0443 <= imem07_in[99:96];
    53: reg_0443 <= op1_03_out;
    55: reg_0443 <= op1_03_out;
    57: reg_0443 <= op1_03_out;
    59: reg_0443 <= op1_03_out;
    61: reg_0443 <= op1_03_out;
    63: reg_0443 <= op1_03_out;
    66: reg_0443 <= imem04_in[87:84];
    67: reg_0443 <= op1_03_out;
    69: reg_0443 <= op1_03_out;
    71: reg_0443 <= op1_03_out;
    73: reg_0443 <= op1_03_out;
    76: reg_0443 <= imem04_in[87:84];
    78: reg_0443 <= imem04_in[87:84];
    79: reg_0443 <= op1_03_out;
    81: reg_0443 <= op1_03_out;
    84: reg_0443 <= imem04_in[87:84];
    85: reg_0443 <= op1_03_out;
    87: reg_0443 <= op1_03_out;
    89: reg_0443 <= op1_03_out;
    91: reg_0443 <= op1_03_out;
    94: reg_0443 <= imem07_in[99:96];
    96: reg_0443 <= imem04_in[87:84];
    97: reg_0443 <= op1_03_out;
    endcase
  end

  // REG#444の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0444 <= imem07_in[91:88];
    44: reg_0444 <= imem07_in[91:88];
    46: reg_0444 <= imem04_in[27:24];
    49: reg_0444 <= imem04_in[27:24];
    57: reg_0444 <= imem04_in[27:24];
    59: reg_0444 <= imem04_in[27:24];
    endcase
  end

  // REG#445の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0445 <= imem07_in[63:60];
    44: reg_0445 <= imem04_in[95:92];
    46: reg_0445 <= imem04_in[95:92];
    49: reg_0445 <= imem07_in[63:60];
    51: reg_0445 <= imem04_in[95:92];
    53: reg_0445 <= imem03_in[59:56];
    55: reg_0445 <= imem03_in[59:56];
    90: reg_0445 <= imem03_in[59:56];
    endcase
  end

  // REG#446の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0446 <= imem07_in[79:76];
    44: reg_0446 <= imem06_in[3:0];
    46: reg_0446 <= imem04_in[23:20];
    50: reg_0446 <= imem05_in[55:52];
    66: reg_0446 <= imem07_in[79:76];
    68: reg_0446 <= imem04_in[23:20];
    71: reg_0446 <= imem05_in[55:52];
    73: reg_0446 <= imem04_in[23:20];
    75: reg_0446 <= imem07_in[79:76];
    79: reg_0446 <= imem04_in[23:20];
    81: reg_0446 <= imem07_in[79:76];
    83: reg_0446 <= imem04_in[23:20];
    92: reg_0446 <= imem06_in[3:0];
    96: reg_0446 <= imem06_in[3:0];
    endcase
  end

  // REG#447の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0447 <= imem07_in[47:44];
    44: reg_0447 <= imem07_in[47:44];
    46: reg_0447 <= imem07_in[47:44];
    48: reg_0447 <= imem07_in[47:44];
    50: reg_0447 <= imem05_in[103:100];
    66: reg_0447 <= imem05_in[103:100];
    78: reg_0447 <= imem05_in[103:100];
    82: reg_0447 <= imem07_in[47:44];
    endcase
  end

  // REG#448の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0448 <= imem07_in[119:116];
    44: reg_0448 <= imem06_in[123:120];
    46: reg_0448 <= imem04_in[115:112];
    50: reg_0448 <= imem05_in[91:88];
    67: reg_0448 <= imem04_in[115:112];
    69: reg_0448 <= imem04_in[115:112];
    71: reg_0448 <= imem05_in[91:88];
    73: reg_0448 <= imem05_in[91:88];
    endcase
  end

  // REG#449の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0449 <= imem07_in[83:80];
    44: reg_0449 <= imem02_in[87:84];
    47: reg_0449 <= imem02_in[87:84];
    49: reg_0449 <= imem02_in[87:84];
    53: reg_0449 <= imem06_in[63:60];
    55: reg_0449 <= imem07_in[83:80];
    57: reg_0449 <= imem07_in[83:80];
    59: reg_0449 <= imem07_in[83:80];
    61: reg_0449 <= imem06_in[63:60];
    70: reg_0449 <= imem02_in[87:84];
    72: reg_0449 <= imem06_in[63:60];
    74: reg_0449 <= imem02_in[87:84];
    76: reg_0449 <= imem02_in[87:84];
    78: reg_0449 <= imem02_in[87:84];
    80: reg_0449 <= imem06_in[63:60];
    82: reg_0449 <= imem07_in[83:80];
    endcase
  end

  // REG#450の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0450 <= imem00_in[19:16];
    93: reg_0450 <= imem00_in[19:16];
    96: reg_0450 <= imem00_in[19:16];
    endcase
  end

  // REG#451の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0451 <= imem00_in[23:20];
    endcase
  end

  // REG#452の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0452 <= imem00_in[115:112];
    95: reg_0452 <= imem00_in[115:112];
    endcase
  end

  // REG#453の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0453 <= imem00_in[11:8];
    endcase
  end

  // REG#454の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0454 <= imem00_in[15:12];
    endcase
  end

  // REG#455の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0455 <= imem00_in[27:24];
    endcase
  end

  // REG#456の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0456 <= imem00_in[119:116];
    endcase
  end

  // REG#457の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0457 <= imem00_in[31:28];
    endcase
  end

  // REG#458の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0458 <= imem00_in[127:124];
    endcase
  end

  // REG#459の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0459 <= imem00_in[111:108];
    endcase
  end

  // REG#460の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0460 <= imem00_in[63:60];
    endcase
  end

  // REG#461の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0461 <= imem00_in[39:36];
    endcase
  end

  // REG#462の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0462 <= imem00_in[67:64];
    endcase
  end

  // REG#463の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0463 <= imem00_in[3:0];
    endcase
  end

  // REG#464の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0464 <= imem00_in[35:32];
    endcase
  end

  // REG#465の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0465 <= imem00_in[7:4];
    endcase
  end

  // REG#466の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0466 <= imem00_in[55:52];
    endcase
  end

  // REG#467の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0467 <= imem00_in[87:84];
    endcase
  end

  // REG#468の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0468 <= imem00_in[103:100];
    endcase
  end

  // REG#469の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0469 <= imem00_in[47:44];
    endcase
  end

  // REG#470の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0470 <= imem00_in[91:88];
    endcase
  end

  // REG#471の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0471 <= imem00_in[99:96];
    endcase
  end

  // REG#472の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0472 <= imem00_in[75:72];
    endcase
  end

  // REG#473の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0473 <= imem00_in[83:80];
    endcase
  end

  // REG#474の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0474 <= imem00_in[95:92];
    endcase
  end

  // REG#475の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0475 <= imem00_in[59:56];
    endcase
  end

  // REG#476の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0476 <= imem00_in[51:48];
    endcase
  end

  // REG#477の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0477 <= imem00_in[43:40];
    endcase
  end

  // REG#478の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0478 <= imem00_in[123:120];
    endcase
  end

  // REG#479の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0479 <= imem00_in[107:104];
    endcase
  end

  // REG#480の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0480 <= imem00_in[79:76];
    endcase
  end

  // REG#481の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0481 <= imem00_in[71:68];
    endcase
  end

  // REG#482の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0482 <= imem05_in[19:16];
    7: reg_0482 <= imem05_in[47:44];
    9: reg_0482 <= imem05_in[19:16];
    11: reg_0482 <= imem06_in[103:100];
    13: reg_0482 <= imem06_in[103:100];
    15: reg_0482 <= imem02_in[11:8];
    17: reg_0482 <= imem05_in[19:16];
    19: reg_0482 <= imem02_in[11:8];
    21: reg_0482 <= imem02_in[11:8];
    85: reg_0482 <= imem06_in[103:100];
    88: reg_0482 <= imem05_in[47:44];
    90: reg_0482 <= imem05_in[47:44];
    92: reg_0482 <= imem05_in[47:44];
    94: reg_0482 <= imem02_in[11:8];
    96: reg_0482 <= imem05_in[47:44];
    endcase
  end

  // REG#483の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0483 <= imem05_in[23:20];
    7: reg_0483 <= imem05_in[23:20];
    9: reg_0483 <= imem04_in[7:4];
    11: reg_0483 <= imem04_in[7:4];
    13: reg_0483 <= imem04_in[7:4];
    15: reg_0483 <= imem03_in[127:124];
    17: reg_0483 <= imem04_in[7:4];
    19: reg_0483 <= imem05_in[23:20];
    22: reg_0483 <= imem03_in[127:124];
    24: reg_0483 <= imem04_in[7:4];
    84: reg_0483 <= imem02_in[79:76];
    endcase
  end

  // REG#484の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0484 <= imem05_in[43:40];
    7: reg_0484 <= imem05_in[43:40];
    9: reg_0484 <= imem04_in[91:88];
    11: reg_0484 <= imem04_in[91:88];
    13: reg_0484 <= imem02_in[91:88];
    15: reg_0484 <= imem04_in[91:88];
    17: reg_0484 <= imem04_in[91:88];
    21: reg_0484 <= imem02_in[91:88];
    86: reg_0484 <= imem02_in[91:88];
    88: reg_0484 <= imem05_in[43:40];
    90: reg_0484 <= imem07_in[127:124];
    92: reg_0484 <= imem07_in[127:124];
    94: reg_0484 <= imem05_in[43:40];
    96: reg_0484 <= imem04_in[91:88];
    endcase
  end

  // REG#485の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0485 <= imem05_in[115:112];
    7: reg_0485 <= imem05_in[115:112];
    9: reg_0485 <= imem04_in[107:104];
    11: reg_0485 <= imem05_in[115:112];
    13: reg_0485 <= imem05_in[115:112];
    15: reg_0485 <= imem05_in[51:48];
    17: reg_0485 <= imem04_in[107:104];
    21: reg_0485 <= imem04_in[107:104];
    23: reg_0485 <= imem05_in[51:48];
    25: reg_0485 <= imem02_in[83:80];
    27: reg_0485 <= imem05_in[115:112];
    30: reg_0485 <= imem02_in[83:80];
    32: reg_0485 <= imem02_in[83:80];
    34: reg_0485 <= imem02_in[83:80];
    36: reg_0485 <= imem04_in[107:104];
    38: reg_0485 <= imem05_in[115:112];
    41: reg_0485 <= imem05_in[115:112];
    43: reg_0485 <= imem02_in[83:80];
    45: reg_0485 <= imem04_in[107:104];
    47: reg_0485 <= imem05_in[51:48];
    49: reg_0485 <= imem05_in[115:112];
    51: reg_0485 <= imem05_in[51:48];
    53: reg_0485 <= imem04_in[107:104];
    55: reg_0485 <= imem05_in[51:48];
    58: reg_0485 <= imem05_in[51:48];
    60: reg_0485 <= imem02_in[83:80];
    62: reg_0485 <= imem02_in[83:80];
    65: reg_0485 <= imem06_in[71:68];
    67: reg_0485 <= imem04_in[107:104];
    69: reg_0485 <= imem04_in[107:104];
    71: reg_0485 <= imem06_in[71:68];
    87: reg_0485 <= imem02_in[83:80];
    89: reg_0485 <= imem02_in[83:80];
    91: reg_0485 <= imem04_in[107:104];
    93: reg_0485 <= imem02_in[83:80];
    95: reg_0485 <= imem05_in[51:48];
    endcase
  end

  // REG#486の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0486 <= imem05_in[127:124];
    7: reg_0486 <= imem06_in[43:40];
    9: reg_0486 <= imem06_in[43:40];
    32: reg_0486 <= imem06_in[43:40];
    35: reg_0486 <= imem06_in[43:40];
    39: reg_0486 <= imem06_in[43:40];
    56: reg_0486 <= imem06_in[43:40];
    60: reg_0486 <= imem05_in[31:28];
    62: reg_0486 <= imem05_in[127:124];
    64: reg_0486 <= imem06_in[43:40];
    66: reg_0486 <= imem06_in[43:40];
    68: reg_0486 <= imem05_in[127:124];
    74: reg_0486 <= imem05_in[31:28];
    endcase
  end

  // REG#487の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0487 <= imem01_in[99:96];
    7: reg_0487 <= imem01_in[99:96];
    9: reg_0487 <= imem04_in[111:108];
    11: reg_0487 <= imem01_in[99:96];
    25: reg_0487 <= imem01_in[99:96];
    47: reg_0487 <= imem06_in[3:0];
    49: reg_0487 <= imem01_in[99:96];
    69: reg_0487 <= imem01_in[99:96];
    90: reg_0487 <= imem01_in[99:96];
    92: reg_0487 <= imem01_in[99:96];
    95: reg_0487 <= imem04_in[111:108];
    endcase
  end

  // REG#488の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0488 <= imem05_in[39:36];
    7: reg_0488 <= imem06_in[79:76];
    9: reg_0488 <= imem05_in[39:36];
    11: reg_0488 <= imem05_in[39:36];
    14: reg_0488 <= imem05_in[39:36];
    16: reg_0488 <= imem01_in[83:80];
    18: reg_0488 <= imem01_in[83:80];
    20: reg_0488 <= imem01_in[83:80];
    22: reg_0488 <= imem05_in[39:36];
    24: reg_0488 <= imem05_in[39:36];
    26: reg_0488 <= imem05_in[39:36];
    28: reg_0488 <= imem05_in[39:36];
    30: reg_0488 <= imem01_in[83:80];
    32: reg_0488 <= imem05_in[39:36];
    34: reg_0488 <= imem05_in[39:36];
    36: reg_0488 <= imem01_in[83:80];
    38: reg_0488 <= imem01_in[115:112];
    40: reg_0488 <= imem06_in[79:76];
    42: reg_0488 <= imem05_in[39:36];
    44: reg_0488 <= imem05_in[39:36];
    46: reg_0488 <= imem06_in[79:76];
    48: reg_0488 <= imem05_in[39:36];
    50: reg_0488 <= imem05_in[39:36];
    65: reg_0488 <= imem05_in[39:36];
    69: reg_0488 <= imem01_in[83:80];
    95: reg_0488 <= imem05_in[39:36];
    endcase
  end

  // REG#489の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0489 <= imem05_in[123:120];
    7: reg_0489 <= imem05_in[123:120];
    9: reg_0489 <= imem04_in[115:112];
    11: reg_0489 <= imem05_in[123:120];
    14: reg_0489 <= imem05_in[123:120];
    16: reg_0489 <= imem05_in[123:120];
    18: reg_0489 <= imem05_in[123:120];
    20: reg_0489 <= imem05_in[123:120];
    48: reg_0489 <= imem05_in[123:120];
    50: reg_0489 <= imem05_in[123:120];
    68: reg_0489 <= imem03_in[107:104];
    70: reg_0489 <= imem04_in[115:112];
    72: reg_0489 <= imem03_in[107:104];
    74: reg_0489 <= imem03_in[107:104];
    76: reg_0489 <= imem05_in[123:120];
    78: reg_0489 <= imem04_in[115:112];
    80: reg_0489 <= imem05_in[115:112];
    82: reg_0489 <= imem01_in[19:16];
    84: reg_0489 <= imem04_in[115:112];
    86: reg_0489 <= imem05_in[115:112];
    89: reg_0489 <= imem01_in[19:16];
    91: reg_0489 <= imem04_in[115:112];
    93: reg_0489 <= imem03_in[107:104];
    95: reg_0489 <= imem04_in[115:112];
    endcase
  end

  // REG#490の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0490 <= imem05_in[35:32];
    7: reg_0490 <= imem07_in[11:8];
    9: reg_0490 <= imem05_in[63:60];
    11: reg_0490 <= imem05_in[63:60];
    13: reg_0490 <= imem05_in[35:32];
    15: reg_0490 <= imem05_in[103:100];
    17: reg_0490 <= imem05_in[63:60];
    19: reg_0490 <= imem05_in[103:100];
    21: reg_0490 <= imem05_in[63:60];
    23: reg_0490 <= imem07_in[11:8];
    25: reg_0490 <= imem07_in[11:8];
    27: reg_0490 <= imem07_in[11:8];
    29: reg_0490 <= imem07_in[11:8];
    31: reg_0490 <= imem01_in[55:52];
    33: reg_0490 <= imem03_in[111:108];
    35: reg_0490 <= imem01_in[55:52];
    37: reg_0490 <= imem05_in[103:100];
    39: reg_0490 <= imem05_in[35:32];
    41: reg_0490 <= imem05_in[35:32];
    43: reg_0490 <= imem05_in[63:60];
    45: reg_0490 <= imem05_in[63:60];
    47: reg_0490 <= imem05_in[103:100];
    49: reg_0490 <= imem05_in[103:100];
    52: reg_0490 <= imem01_in[55:52];
    54: reg_0490 <= imem05_in[103:100];
    56: reg_0490 <= imem07_in[11:8];
    58: reg_0490 <= imem07_in[11:8];
    60: reg_0490 <= imem05_in[63:60];
    63: reg_0490 <= imem01_in[55:52];
    65: reg_0490 <= imem05_in[35:32];
    68: reg_0490 <= imem01_in[55:52];
    72: reg_0490 <= imem05_in[63:60];
    74: reg_0490 <= imem05_in[103:100];
    96: reg_0490 <= imem05_in[63:60];
    endcase
  end

  // REG#491の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0491 <= imem05_in[55:52];
    7: reg_0491 <= imem07_in[23:20];
    9: reg_0491 <= imem05_in[55:52];
    11: reg_0491 <= imem05_in[55:52];
    14: reg_0491 <= imem05_in[55:52];
    16: reg_0491 <= imem02_in[35:32];
    18: reg_0491 <= imem02_in[35:32];
    20: reg_0491 <= imem05_in[55:52];
    50: reg_0491 <= imem07_in[23:20];
    52: reg_0491 <= imem07_in[23:20];
    54: reg_0491 <= imem07_in[23:20];
    56: reg_0491 <= imem02_in[35:32];
    58: reg_0491 <= imem04_in[43:40];
    61: reg_0491 <= imem05_in[55:52];
    66: reg_0491 <= imem07_in[23:20];
    68: reg_0491 <= imem02_in[35:32];
    71: reg_0491 <= imem04_in[43:40];
    73: reg_0491 <= imem04_in[99:96];
    75: reg_0491 <= imem04_in[99:96];
    77: reg_0491 <= imem07_in[23:20];
    79: reg_0491 <= imem02_in[35:32];
    82: reg_0491 <= imem04_in[43:40];
    84: reg_0491 <= imem05_in[55:52];
    86: reg_0491 <= imem04_in[43:40];
    88: reg_0491 <= imem07_in[23:20];
    90: reg_0491 <= imem02_in[35:32];
    92: reg_0491 <= imem04_in[99:96];
    94: reg_0491 <= imem04_in[43:40];
    96: reg_0491 <= imem07_in[23:20];
    endcase
  end

  // REG#492の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0492 <= imem05_in[59:56];
    7: reg_0492 <= imem05_in[59:56];
    9: reg_0492 <= imem07_in[39:36];
    11: reg_0492 <= imem07_in[39:36];
    13: reg_0492 <= imem07_in[39:36];
    15: reg_0492 <= imem07_in[39:36];
    17: reg_0492 <= imem05_in[59:56];
    19: reg_0492 <= imem03_in[27:24];
    21: reg_0492 <= imem03_in[27:24];
    23: reg_0492 <= imem00_in[47:44];
    25: reg_0492 <= imem07_in[39:36];
    27: reg_0492 <= imem07_in[39:36];
    29: reg_0492 <= imem07_in[39:36];
    31: reg_0492 <= imem03_in[27:24];
    52: reg_0492 <= imem00_in[47:44];
    54: reg_0492 <= imem07_in[39:36];
    56: reg_0492 <= imem05_in[59:56];
    61: reg_0492 <= imem05_in[23:20];
    63: reg_0492 <= imem03_in[27:24];
    65: reg_0492 <= imem00_in[47:44];
    67: reg_0492 <= imem03_in[27:24];
    69: reg_0492 <= imem07_in[39:36];
    71: reg_0492 <= imem07_in[39:36];
    73: reg_0492 <= imem05_in[23:20];
    endcase
  end

  // REG#493の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0493 <= imem05_in[67:64];
    7: reg_0493 <= imem05_in[67:64];
    9: reg_0493 <= imem05_in[67:64];
    11: reg_0493 <= imem07_in[3:0];
    13: reg_0493 <= imem05_in[67:64];
    15: reg_0493 <= imem07_in[3:0];
    17: reg_0493 <= imem02_in[35:32];
    19: reg_0493 <= imem07_in[3:0];
    21: reg_0493 <= imem05_in[67:64];
    23: reg_0493 <= imem02_in[35:32];
    25: reg_0493 <= imem07_in[3:0];
    27: reg_0493 <= imem03_in[3:0];
    30: reg_0493 <= imem05_in[67:64];
    32: reg_0493 <= imem07_in[3:0];
    34: reg_0493 <= imem05_in[67:64];
    36: reg_0493 <= imem02_in[115:112];
    38: reg_0493 <= imem07_in[3:0];
    40: reg_0493 <= imem03_in[3:0];
    42: reg_0493 <= imem05_in[67:64];
    44: reg_0493 <= imem07_in[3:0];
    46: reg_0493 <= imem03_in[3:0];
    48: reg_0493 <= imem05_in[67:64];
    50: reg_0493 <= imem05_in[67:64];
    67: reg_0493 <= imem02_in[35:32];
    69: reg_0493 <= imem07_in[3:0];
    71: reg_0493 <= imem07_in[3:0];
    72: reg_0493 <= op1_00_out;
    74: reg_0493 <= op1_00_out;
    76: reg_0493 <= op1_00_out;
    78: reg_0493 <= op1_00_out;
    80: reg_0493 <= op1_00_out;
    83: reg_0493 <= imem07_in[3:0];
    85: reg_0493 <= imem02_in[115:112];
    endcase
  end

  // REG#494の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0494 <= imem05_in[75:72];
    7: reg_0494 <= imem07_in[47:44];
    9: reg_0494 <= imem07_in[47:44];
    11: reg_0494 <= imem05_in[75:72];
    13: reg_0494 <= imem05_in[75:72];
    15: reg_0494 <= imem05_in[75:72];
    17: reg_0494 <= imem07_in[47:44];
    19: reg_0494 <= imem03_in[99:96];
    21: reg_0494 <= imem03_in[99:96];
    23: reg_0494 <= imem03_in[99:96];
    25: reg_0494 <= imem03_in[99:96];
    27: reg_0494 <= imem07_in[47:44];
    29: reg_0494 <= imem07_in[47:44];
    31: reg_0494 <= imem07_in[47:44];
    33: reg_0494 <= imem05_in[75:72];
    35: reg_0494 <= imem00_in[103:100];
    37: reg_0494 <= imem07_in[47:44];
    39: reg_0494 <= imem01_in[35:32];
    41: reg_0494 <= imem03_in[99:96];
    43: reg_0494 <= imem03_in[99:96];
    45: reg_0494 <= imem05_in[75:72];
    47: reg_0494 <= imem07_in[47:44];
    49: reg_0494 <= imem05_in[75:72];
    53: reg_0494 <= imem05_in[75:72];
    55: reg_0494 <= imem01_in[35:32];
    57: reg_0494 <= imem05_in[75:72];
    59: reg_0494 <= imem04_in[43:40];
    endcase
  end

  // REG#495の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0495 <= imem05_in[87:84];
    7: reg_0495 <= imem05_in[87:84];
    9: reg_0495 <= imem02_in[107:104];
    11: reg_0495 <= imem05_in[87:84];
    13: reg_0495 <= imem02_in[107:104];
    15: reg_0495 <= imem06_in[123:120];
    17: reg_0495 <= imem06_in[123:120];
    19: reg_0495 <= imem05_in[87:84];
    21: reg_0495 <= imem06_in[123:120];
    23: reg_0495 <= imem00_in[55:52];
    25: reg_0495 <= imem06_in[123:120];
    27: reg_0495 <= imem00_in[55:52];
    29: reg_0495 <= imem05_in[87:84];
    31: reg_0495 <= imem05_in[87:84];
    33: reg_0495 <= imem06_in[123:120];
    35: reg_0495 <= imem00_in[55:52];
    37: reg_0495 <= imem00_in[55:52];
    39: reg_0495 <= imem06_in[123:120];
    57: reg_0495 <= imem00_in[55:52];
    59: reg_0495 <= imem04_in[59:56];
    endcase
  end

  // REG#496の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0496 <= imem01_in[19:16];
    8: reg_0496 <= imem01_in[19:16];
    10: reg_0496 <= imem01_in[19:16];
    41: reg_0496 <= imem01_in[19:16];
    93: reg_0496 <= imem06_in[23:20];
    endcase
  end

  // REG#497の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0497 <= op1_00_out;
    7: reg_0497 <= op1_00_out;
    10: reg_0497 <= imem04_in[87:84];
    12: reg_0497 <= imem04_in[87:84];
    14: reg_0497 <= imem05_in[127:124];
    16: reg_0497 <= imem02_in[51:48];
    18: reg_0497 <= imem07_in[27:24];
    20: reg_0497 <= imem05_in[127:124];
    48: reg_0497 <= imem02_in[51:48];
    50: reg_0497 <= imem05_in[127:124];
    64: reg_0497 <= imem05_in[127:124];
    67: reg_0497 <= imem05_in[127:124];
    68: reg_0497 <= op1_00_out;
    70: reg_0497 <= op1_00_out;
    73: reg_0497 <= imem07_in[27:24];
    75: reg_0497 <= imem04_in[87:84];
    78: reg_0497 <= imem02_in[51:48];
    80: reg_0497 <= imem07_in[27:24];
    84: reg_0497 <= imem05_in[127:124];
    86: reg_0497 <= imem04_in[87:84];
    88: reg_0497 <= imem05_in[127:124];
    90: reg_0497 <= imem01_in[19:16];
    92: reg_0497 <= imem05_in[127:124];
    94: reg_0497 <= imem02_in[51:48];
    96: reg_0497 <= imem05_in[127:124];
    endcase
  end

  // REG#498の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0498 <= imem01_in[115:112];
    9: reg_0498 <= imem03_in[55:52];
    11: reg_0498 <= imem03_in[55:52];
    13: reg_0498 <= imem02_in[95:92];
    14: reg_0498 <= op2_00_out;
    35: reg_0498 <= op2_00_out;
    64: reg_0498 <= imem01_in[115:112];
    65: reg_0498 <= op2_00_out;
    75: reg_0498 <= op2_00_out;
    endcase
  end

  // REG#499の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0499 <= imem01_in[75:72];
    9: reg_0499 <= imem01_in[75:72];
    11: reg_0499 <= imem07_in[87:84];
    13: reg_0499 <= imem01_in[75:72];
    15: reg_0499 <= imem07_in[87:84];
    17: reg_0499 <= imem01_in[75:72];
    19: reg_0499 <= imem07_in[87:84];
    21: reg_0499 <= imem07_in[87:84];
    23: reg_0499 <= imem00_in[87:84];
    25: reg_0499 <= imem07_in[87:84];
    27: reg_0499 <= imem07_in[87:84];
    30: reg_0499 <= imem00_in[87:84];
    32: reg_0499 <= imem02_in[75:72];
    34: reg_0499 <= imem07_in[87:84];
    36: reg_0499 <= imem00_in[87:84];
    38: reg_0499 <= imem00_in[87:84];
    40: reg_0499 <= imem00_in[87:84];
    42: reg_0499 <= imem00_in[51:48];
    44: reg_0499 <= imem02_in[75:72];
    46: reg_0499 <= imem02_in[75:72];
    48: reg_0499 <= imem04_in[99:96];
    51: reg_0499 <= imem02_in[75:72];
    53: reg_0499 <= imem07_in[87:84];
    55: reg_0499 <= imem00_in[87:84];
    86: reg_0499 <= imem07_in[87:84];
    88: reg_0499 <= imem07_in[87:84];
    90: reg_0499 <= imem00_in[51:48];
    92: reg_0499 <= imem07_in[87:84];
    94: reg_0499 <= imem07_in[87:84];
    96: reg_0499 <= imem01_in[75:72];
    endcase
  end

  // REG#500の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0500 <= imem01_in[55:52];
    10: reg_0500 <= imem01_in[55:52];
    41: reg_0500 <= imem01_in[55:52];
    94: reg_0500 <= imem01_in[55:52];
    endcase
  end

  // REG#501の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0501 <= imem01_in[11:8];
    10: reg_0501 <= imem04_in[111:108];
    12: reg_0501 <= imem01_in[11:8];
    14: reg_0501 <= imem01_in[11:8];
    16: reg_0501 <= imem01_in[11:8];
    18: reg_0501 <= imem07_in[67:64];
    20: reg_0501 <= imem04_in[111:108];
    22: reg_0501 <= imem01_in[11:8];
    24: reg_0501 <= imem07_in[67:64];
    26: reg_0501 <= imem04_in[111:108];
    28: reg_0501 <= imem01_in[11:8];
    29: reg_0501 <= op1_15_out;
    32: reg_0501 <= imem04_in[111:108];
    34: reg_0501 <= imem01_in[11:8];
    36: reg_0501 <= imem04_in[111:108];
    38: reg_0501 <= imem04_in[111:108];
    41: reg_0501 <= imem01_in[11:8];
    93: reg_0501 <= imem01_in[11:8];
    96: reg_0501 <= imem07_in[67:64];
    endcase
  end

  // REG#502の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0502 <= imem01_in[59:56];
    11: reg_0502 <= imem01_in[59:56];
    26: reg_0502 <= imem07_in[107:104];
    28: reg_0502 <= imem00_in[95:92];
    30: reg_0502 <= imem03_in[15:12];
    33: reg_0502 <= imem01_in[59:56];
    35: reg_0502 <= imem01_in[59:56];
    37: reg_0502 <= imem00_in[95:92];
    39: reg_0502 <= imem00_in[95:92];
    41: reg_0502 <= imem00_in[95:92];
    43: reg_0502 <= imem07_in[107:104];
    94: reg_0502 <= imem00_in[95:92];
    96: reg_0502 <= imem00_in[95:92];
    endcase
  end

  // REG#503の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0503 <= imem01_in[79:76];
    11: reg_0503 <= imem01_in[79:76];
    26: reg_0503 <= imem00_in[43:40];
    28: reg_0503 <= imem00_in[43:40];
    30: reg_0503 <= imem03_in[111:108];
    33: reg_0503 <= imem00_in[43:40];
    35: reg_0503 <= imem03_in[111:108];
    37: reg_0503 <= imem01_in[79:76];
    39: reg_0503 <= imem01_in[79:76];
    43: reg_0503 <= imem05_in[79:76];
    45: reg_0503 <= imem03_in[111:108];
    47: reg_0503 <= imem00_in[43:40];
    49: reg_0503 <= imem01_in[79:76];
    67: reg_0503 <= imem01_in[79:76];
    69: reg_0503 <= imem01_in[79:76];
    94: reg_0503 <= imem01_in[79:76];
    97: reg_0503 <= imem00_in[43:40];
    endcase
  end

  // REG#504の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0504 <= imem01_in[7:4];
    11: reg_0504 <= imem00_in[99:96];
    13: reg_0504 <= imem01_in[7:4];
    14: reg_0504 <= op2_01_out;
    36: reg_0504 <= op2_01_out;
    68: reg_0504 <= imem01_in[7:4];
    69: reg_0504 <= op2_01_out;
    88: reg_0504 <= op2_01_out;
    endcase
  end

  // REG#505の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0505 <= imem01_in[123:120];
    11: reg_0505 <= imem02_in[55:52];
    13: reg_0505 <= imem01_in[123:120];
    14: reg_0505 <= op2_02_out;
    37: reg_0505 <= op2_02_out;
    71: reg_0505 <= op2_02_out;
    97: reg_0505 <= imem01_in[123:120];
    endcase
  end

  // REG#506の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0506 <= imem01_in[103:100];
    11: reg_0506 <= imem02_in[63:60];
    13: reg_0506 <= imem02_in[127:124];
    15: reg_0506 <= imem01_in[103:100];
    17: reg_0506 <= imem01_in[103:100];
    19: reg_0506 <= imem02_in[63:60];
    21: reg_0506 <= imem02_in[63:60];
    86: reg_0506 <= imem02_in[63:60];
    88: reg_0506 <= imem02_in[115:112];
    90: reg_0506 <= imem00_in[55:52];
    93: reg_0506 <= imem00_in[55:52];
    95: reg_0506 <= imem02_in[127:124];
    endcase
  end

  // REG#507の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0507 <= imem01_in[119:116];
    11: reg_0507 <= imem01_in[119:116];
    26: reg_0507 <= imem00_in[95:92];
    28: reg_0507 <= imem01_in[119:116];
    30: reg_0507 <= imem01_in[119:116];
    32: reg_0507 <= imem01_in[119:116];
    34: reg_0507 <= imem02_in[27:24];
    36: reg_0507 <= imem04_in[3:0];
    38: reg_0507 <= imem01_in[119:116];
    40: reg_0507 <= imem01_in[119:116];
    42: reg_0507 <= imem04_in[3:0];
    endcase
  end

  // REG#508の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0508 <= imem01_in[127:124];
    11: reg_0508 <= imem01_in[127:124];
    21: reg_0508 <= imem04_in[7:4];
    24: reg_0508 <= imem05_in[67:64];
    26: reg_0508 <= imem05_in[67:64];
    28: reg_0508 <= imem02_in[35:32];
    30: reg_0508 <= imem01_in[127:124];
    32: reg_0508 <= imem01_in[127:124];
    34: reg_0508 <= imem03_in[35:32];
    36: reg_0508 <= imem05_in[43:40];
    38: reg_0508 <= imem02_in[107:104];
    40: reg_0508 <= imem03_in[35:32];
    42: reg_0508 <= imem01_in[127:124];
    44: reg_0508 <= imem04_in[7:4];
    46: reg_0508 <= imem02_in[35:32];
    48: reg_0508 <= imem04_in[7:4];
    50: reg_0508 <= imem05_in[43:40];
    66: reg_0508 <= imem05_in[43:40];
    72: reg_0508 <= imem05_in[43:40];
    74: reg_0508 <= imem05_in[43:40];
    endcase
  end

  // REG#509の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0509 <= imem01_in[43:40];
    11: reg_0509 <= imem05_in[51:48];
    13: reg_0509 <= imem03_in[67:64];
    15: reg_0509 <= imem03_in[67:64];
    17: reg_0509 <= imem05_in[51:48];
    19: reg_0509 <= imem05_in[47:44];
    22: reg_0509 <= imem03_in[67:64];
    24: reg_0509 <= imem05_in[71:68];
    26: reg_0509 <= imem04_in[27:24];
    28: reg_0509 <= imem03_in[67:64];
    70: reg_0509 <= imem01_in[43:40];
    72: reg_0509 <= imem05_in[47:44];
    76: reg_0509 <= imem05_in[71:68];
    78: reg_0509 <= imem03_in[67:64];
    80: reg_0509 <= imem05_in[47:44];
    82: reg_0509 <= imem01_in[43:40];
    84: reg_0509 <= imem01_in[43:40];
    86: reg_0509 <= imem03_in[67:64];
    88: reg_0509 <= imem05_in[51:48];
    90: reg_0509 <= imem03_in[103:100];
    93: reg_0509 <= imem05_in[71:68];
    95: reg_0509 <= imem03_in[67:64];
    97: reg_0509 <= imem05_in[71:68];
    endcase
  end

  // REG#510の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0510 <= imem01_in[111:108];
    11: reg_0510 <= imem05_in[83:80];
    13: reg_0510 <= imem06_in[43:40];
    15: reg_0510 <= imem06_in[43:40];
    17: reg_0510 <= imem05_in[83:80];
    19: reg_0510 <= imem01_in[111:108];
    21: reg_0510 <= imem05_in[83:80];
    23: reg_0510 <= imem01_in[39:36];
    25: reg_0510 <= imem01_in[39:36];
    49: reg_0510 <= imem01_in[39:36];
    65: reg_0510 <= imem01_in[39:36];
    67: reg_0510 <= imem05_in[83:80];
    70: reg_0510 <= imem06_in[43:40];
    73: reg_0510 <= imem01_in[111:108];
    75: reg_0510 <= imem01_in[39:36];
    78: reg_0510 <= imem01_in[111:108];
    80: reg_0510 <= imem01_in[39:36];
    82: reg_0510 <= imem01_in[39:36];
    84: reg_0510 <= imem05_in[83:80];
    86: reg_0510 <= imem06_in[43:40];
    endcase
  end

  // REG#511の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0511 <= imem01_in[31:28];
    11: reg_0511 <= imem01_in[31:28];
    21: reg_0511 <= imem04_in[31:28];
    24: reg_0511 <= imem04_in[31:28];
    83: reg_0511 <= imem04_in[31:28];
    96: reg_0511 <= imem01_in[31:28];
    endcase
  end

  // REG#512の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0512 <= imem01_in[27:24];
    11: reg_0512 <= imem05_in[103:100];
    13: reg_0512 <= imem06_in[51:48];
    15: reg_0512 <= imem01_in[27:24];
    17: reg_0512 <= imem05_in[103:100];
    19: reg_0512 <= imem05_in[11:8];
    22: reg_0512 <= imem05_in[103:100];
    24: reg_0512 <= imem05_in[11:8];
    26: reg_0512 <= imem05_in[11:8];
    28: reg_0512 <= imem01_in[27:24];
    30: reg_0512 <= imem05_in[103:100];
    32: reg_0512 <= imem01_in[27:24];
    34: reg_0512 <= imem05_in[11:8];
    36: reg_0512 <= imem05_in[11:8];
    38: reg_0512 <= imem05_in[11:8];
    40: reg_0512 <= imem06_in[51:48];
    42: reg_0512 <= imem05_in[11:8];
    44: reg_0512 <= imem05_in[103:100];
    46: reg_0512 <= imem05_in[11:8];
    48: reg_0512 <= imem04_in[107:104];
    51: reg_0512 <= imem01_in[27:24];
    53: reg_0512 <= imem01_in[27:24];
    endcase
  end

  // REG#513の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0513 <= imem01_in[23:20];
    12: reg_0513 <= imem03_in[107:104];
    14: reg_0513 <= imem03_in[107:104];
    16: reg_0513 <= imem01_in[23:20];
    18: reg_0513 <= imem01_in[87:84];
    20: reg_0513 <= imem01_in[23:20];
    22: reg_0513 <= imem06_in[3:0];
    24: reg_0513 <= imem03_in[107:104];
    26: reg_0513 <= imem00_in[15:12];
    28: reg_0513 <= imem03_in[107:104];
    71: reg_0513 <= imem00_in[15:12];
    73: reg_0513 <= imem03_in[107:104];
    75: reg_0513 <= imem01_in[87:84];
    77: reg_0513 <= imem03_in[107:104];
    79: reg_0513 <= imem03_in[107:104];
    82: reg_0513 <= imem00_in[15:12];
    84: reg_0513 <= imem00_in[15:12];
    86: reg_0513 <= imem03_in[107:104];
    88: reg_0513 <= imem00_in[15:12];
    90: reg_0513 <= imem00_in[15:12];
    93: reg_0513 <= imem06_in[3:0];
    95: reg_0513 <= imem01_in[87:84];
    endcase
  end

  // REG#514の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0514 <= imem01_in[47:44];
    12: reg_0514 <= imem01_in[47:44];
    14: reg_0514 <= imem01_in[47:44];
    16: reg_0514 <= imem01_in[47:44];
    18: reg_0514 <= imem01_in[99:96];
    20: reg_0514 <= imem01_in[99:96];
    22: reg_0514 <= imem01_in[47:44];
    24: reg_0514 <= imem01_in[47:44];
    26: reg_0514 <= imem01_in[47:44];
    28: reg_0514 <= imem01_in[99:96];
    30: reg_0514 <= imem01_in[99:96];
    32: reg_0514 <= imem02_in[91:88];
    34: reg_0514 <= imem03_in[39:36];
    36: reg_0514 <= imem01_in[99:96];
    38: reg_0514 <= imem02_in[91:88];
    41: reg_0514 <= imem01_in[47:44];
    92: reg_0514 <= imem01_in[47:44];
    95: reg_0514 <= imem03_in[39:36];
    endcase
  end

  // REG#515の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0515 <= imem01_in[95:92];
    12: reg_0515 <= imem01_in[95:92];
    14: reg_0515 <= imem01_in[95:92];
    16: reg_0515 <= imem03_in[71:68];
    18: reg_0515 <= imem01_in[95:92];
    20: reg_0515 <= imem01_in[95:92];
    22: reg_0515 <= imem01_in[95:92];
    24: reg_0515 <= imem07_in[71:68];
    26: reg_0515 <= imem07_in[71:68];
    28: reg_0515 <= imem07_in[71:68];
    30: reg_0515 <= imem03_in[71:68];
    33: reg_0515 <= imem07_in[71:68];
    35: reg_0515 <= imem02_in[51:48];
    37: reg_0515 <= imem07_in[51:48];
    39: reg_0515 <= imem01_in[95:92];
    41: reg_0515 <= imem03_in[71:68];
    43: reg_0515 <= imem03_in[71:68];
    45: reg_0515 <= imem02_in[51:48];
    64: reg_0515 <= imem07_in[51:48];
    66: reg_0515 <= imem07_in[51:48];
    68: reg_0515 <= imem07_in[51:48];
    71: reg_0515 <= imem01_in[95:92];
    73: reg_0515 <= imem07_in[71:68];
    75: reg_0515 <= imem07_in[71:68];
    79: reg_0515 <= imem07_in[71:68];
    94: reg_0515 <= imem01_in[95:92];
    endcase
  end

  // REG#516の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0516 <= imem01_in[107:104];
    12: reg_0516 <= imem03_in[127:124];
    14: reg_0516 <= imem06_in[103:100];
    16: reg_0516 <= imem01_in[107:104];
    18: reg_0516 <= imem02_in[115:112];
    20: reg_0516 <= imem03_in[127:124];
    22: reg_0516 <= imem06_in[103:100];
    24: reg_0516 <= imem06_in[103:100];
    26: reg_0516 <= imem02_in[115:112];
    50: reg_0516 <= imem06_in[103:100];
    52: reg_0516 <= imem02_in[115:112];
    endcase
  end

  // REG#517の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0517 <= imem01_in[83:80];
    12: reg_0517 <= imem04_in[51:48];
    14: reg_0517 <= imem07_in[79:76];
    16: reg_0517 <= imem04_in[51:48];
    18: reg_0517 <= imem04_in[51:48];
    44: reg_0517 <= imem02_in[39:36];
    47: reg_0517 <= imem01_in[83:80];
    49: reg_0517 <= imem04_in[51:48];
    59: reg_0517 <= imem04_in[51:48];
    endcase
  end

  // REG#518の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0518 <= imem01_in[91:88];
    12: reg_0518 <= imem06_in[47:44];
    14: reg_0518 <= imem06_in[47:44];
    16: reg_0518 <= imem06_in[47:44];
    18: reg_0518 <= imem03_in[103:100];
    20: reg_0518 <= imem03_in[103:100];
    22: reg_0518 <= imem06_in[47:44];
    24: reg_0518 <= imem00_in[35:32];
    26: reg_0518 <= imem03_in[103:100];
    28: reg_0518 <= imem03_in[103:100];
    67: reg_0518 <= imem00_in[35:32];
    69: reg_0518 <= imem01_in[91:88];
    93: reg_0518 <= imem07_in[63:60];
    95: reg_0518 <= imem07_in[63:60];
    97: reg_0518 <= imem06_in[47:44];
    endcase
  end

  // REG#519の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0519 <= imem01_in[67:64];
    12: reg_0519 <= imem01_in[67:64];
    14: reg_0519 <= imem00_in[11:8];
    16: reg_0519 <= imem00_in[11:8];
    18: reg_0519 <= imem01_in[67:64];
    20: reg_0519 <= imem04_in[99:96];
    22: reg_0519 <= imem06_in[55:52];
    24: reg_0519 <= imem00_in[11:8];
    26: reg_0519 <= imem04_in[99:96];
    28: reg_0519 <= imem00_in[11:8];
    30: reg_0519 <= imem01_in[67:64];
    32: reg_0519 <= imem04_in[99:96];
    34: reg_0519 <= imem00_in[11:8];
    36: reg_0519 <= imem06_in[55:52];
    38: reg_0519 <= imem00_in[11:8];
    41: reg_0519 <= imem00_in[11:8];
    43: reg_0519 <= imem06_in[19:16];
    45: reg_0519 <= imem00_in[15:12];
    47: reg_0519 <= imem04_in[99:96];
    49: reg_0519 <= imem00_in[15:12];
    51: reg_0519 <= imem00_in[11:8];
    53: reg_0519 <= imem04_in[99:96];
    55: reg_0519 <= imem00_in[15:12];
    92: reg_0519 <= imem01_in[67:64];
    endcase
  end

  // REG#520の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0520 <= imem01_in[35:32];
    12: reg_0520 <= imem01_in[35:32];
    14: reg_0520 <= imem01_in[35:32];
    16: reg_0520 <= imem03_in[107:104];
    18: reg_0520 <= imem06_in[15:12];
    20: reg_0520 <= imem03_in[107:104];
    22: reg_0520 <= imem01_in[35:32];
    24: reg_0520 <= imem06_in[15:12];
    26: reg_0520 <= imem06_in[15:12];
    28: reg_0520 <= imem02_in[99:96];
    30: reg_0520 <= imem01_in[35:32];
    32: reg_0520 <= imem01_in[35:32];
    34: reg_0520 <= imem02_in[99:96];
    36: reg_0520 <= imem02_in[99:96];
    38: reg_0520 <= imem06_in[15:12];
    41: reg_0520 <= imem01_in[35:32];
    93: reg_0520 <= imem01_in[35:32];
    96: reg_0520 <= imem01_in[35:32];
    endcase
  end

  // REG#521の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0521 <= imem01_in[71:68];
    12: reg_0521 <= imem01_in[71:68];
    14: reg_0521 <= imem01_in[87:84];
    16: reg_0521 <= imem05_in[27:24];
    18: reg_0521 <= imem01_in[71:68];
    20: reg_0521 <= imem01_in[71:68];
    22: reg_0521 <= imem06_in[59:56];
    24: reg_0521 <= imem01_in[87:84];
    27: reg_0521 <= imem01_in[87:84];
    29: reg_0521 <= imem05_in[27:24];
    31: reg_0521 <= imem05_in[27:24];
    33: reg_0521 <= imem05_in[27:24];
    35: reg_0521 <= imem06_in[59:56];
    39: reg_0521 <= imem01_in[71:68];
    41: reg_0521 <= imem01_in[87:84];
    91: reg_0521 <= imem00_in[91:88];
    endcase
  end

  // REG#522の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0522 <= imem01_in[15:12];
    12: reg_0522 <= imem00_in[103:100];
    14: reg_0522 <= imem01_in[15:12];
    16: reg_0522 <= imem00_in[103:100];
    18: reg_0522 <= imem06_in[99:96];
    20: reg_0522 <= imem00_in[103:100];
    22: reg_0522 <= imem06_in[99:96];
    24: reg_0522 <= imem00_in[103:100];
    26: reg_0522 <= imem01_in[15:12];
    28: reg_0522 <= imem00_in[103:100];
    30: reg_0522 <= imem01_in[15:12];
    32: reg_0522 <= imem00_in[103:100];
    34: reg_0522 <= imem06_in[99:96];
    36: reg_0522 <= imem00_in[103:100];
    38: reg_0522 <= imem00_in[103:100];
    41: reg_0522 <= imem01_in[15:12];
    95: reg_0522 <= imem01_in[15:12];
    endcase
  end

  // REG#523の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0523 <= imem01_in[3:0];
    12: reg_0523 <= imem02_in[63:60];
    14: reg_0523 <= imem01_in[103:100];
    16: reg_0523 <= imem01_in[103:100];
    18: reg_0523 <= imem01_in[3:0];
    20: reg_0523 <= imem01_in[3:0];
    22: reg_0523 <= imem01_in[103:100];
    24: reg_0523 <= imem00_in[43:40];
    26: reg_0523 <= imem01_in[103:100];
    28: reg_0523 <= imem01_in[3:0];
    30: reg_0523 <= imem01_in[3:0];
    32: reg_0523 <= imem01_in[3:0];
    34: reg_0523 <= imem00_in[43:40];
    36: reg_0523 <= imem00_in[43:40];
    38: reg_0523 <= imem00_in[43:40];
    40: reg_0523 <= imem00_in[43:40];
    42: reg_0523 <= imem01_in[3:0];
    44: reg_0523 <= imem01_in[103:100];
    46: reg_0523 <= imem02_in[63:60];
    48: reg_0523 <= imem01_in[3:0];
    50: reg_0523 <= imem02_in[63:60];
    52: reg_0523 <= imem01_in[103:100];
    55: reg_0523 <= imem00_in[43:40];
    90: reg_0523 <= imem03_in[39:36];
    endcase
  end

  // REG#524の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0524 <= imem01_in[63:60];
    12: reg_0524 <= imem02_in[87:84];
    14: reg_0524 <= imem01_in[63:60];
    16: reg_0524 <= imem02_in[87:84];
    18: reg_0524 <= imem03_in[91:88];
    20: reg_0524 <= imem07_in[55:52];
    22: reg_0524 <= imem03_in[91:88];
    24: reg_0524 <= imem07_in[55:52];
    26: reg_0524 <= imem03_in[91:88];
    28: reg_0524 <= imem01_in[63:60];
    30: reg_0524 <= imem01_in[63:60];
    32: reg_0524 <= imem04_in[31:28];
    34: reg_0524 <= imem02_in[87:84];
    36: reg_0524 <= imem05_in[71:68];
    38: reg_0524 <= imem03_in[91:88];
    40: reg_0524 <= imem02_in[87:84];
    42: reg_0524 <= imem04_in[31:28];
    95: reg_0524 <= imem01_in[63:60];
    endcase
  end

  // REG#525の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0525 <= op1_01_out;
    11: reg_0525 <= op1_01_out;
    13: reg_0525 <= op1_01_out;
    16: reg_0525 <= imem05_in[31:28];
    18: reg_0525 <= imem04_in[7:4];
    44: reg_0525 <= imem05_in[31:28];
    46: reg_0525 <= imem04_in[55:52];
    50: reg_0525 <= imem04_in[55:52];
    53: reg_0525 <= imem04_in[55:52];
    55: reg_0525 <= imem04_in[7:4];
    57: reg_0525 <= imem05_in[31:28];
    59: reg_0525 <= imem05_in[31:28];
    61: reg_0525 <= imem04_in[55:52];
    62: reg_0525 <= op1_01_out;
    65: reg_0525 <= imem04_in[7:4];
    67: reg_0525 <= imem04_in[7:4];
    69: reg_0525 <= imem04_in[7:4];
    70: reg_0525 <= op1_01_out;
    72: reg_0525 <= op1_01_out;
    74: reg_0525 <= op1_01_out;
    77: reg_0525 <= imem04_in[55:52];
    79: reg_0525 <= imem05_in[31:28];
    88: reg_0525 <= imem05_in[31:28];
    91: reg_0525 <= imem04_in[55:52];
    92: reg_0525 <= op1_01_out;
    95: reg_0525 <= imem05_in[31:28];
    96: reg_0525 <= op1_01_out;
    endcase
  end

  // REG#526の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0526 <= op1_02_out;
    12: reg_0526 <= op1_02_out;
    14: reg_0526 <= op1_02_out;
    16: reg_0526 <= op1_02_out;
    18: reg_0526 <= op1_02_out;
    20: reg_0526 <= op1_02_out;
    22: reg_0526 <= op1_02_out;
    24: reg_0526 <= op1_02_out;
    26: reg_0526 <= op1_02_out;
    28: reg_0526 <= op1_02_out;
    30: reg_0526 <= op1_02_out;
    32: reg_0526 <= op1_02_out;
    34: reg_0526 <= op1_02_out;
    36: reg_0526 <= op1_02_out;
    38: reg_0526 <= op1_02_out;
    40: reg_0526 <= op1_02_out;
    42: reg_0526 <= op1_02_out;
    44: reg_0526 <= op1_02_out;
    46: reg_0526 <= op1_02_out;
    48: reg_0526 <= op1_02_out;
    50: reg_0526 <= op1_02_out;
    52: reg_0526 <= op1_02_out;
    54: reg_0526 <= op1_02_out;
    56: reg_0526 <= op1_02_out;
    58: reg_0526 <= op1_02_out;
    60: reg_0526 <= op1_02_out;
    62: reg_0526 <= op1_02_out;
    64: reg_0526 <= op1_02_out;
    66: reg_0526 <= op1_02_out;
    68: reg_0526 <= op1_02_out;
    70: reg_0526 <= op1_02_out;
    72: reg_0526 <= op1_02_out;
    74: reg_0526 <= op1_02_out;
    76: reg_0526 <= op1_02_out;
    78: reg_0526 <= op1_02_out;
    80: reg_0526 <= op1_02_out;
    82: reg_0526 <= op1_02_out;
    84: reg_0526 <= op1_02_out;
    86: reg_0526 <= op1_02_out;
    88: reg_0526 <= op1_02_out;
    90: reg_0526 <= op1_02_out;
    92: reg_0526 <= op1_02_out;
    94: reg_0526 <= op1_02_out;
    96: reg_0526 <= op1_02_out;
    endcase
  end

  // REG#527の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0527 <= op1_03_out;
    12: reg_0527 <= op1_03_out;
    14: reg_0527 <= op1_03_out;
    16: reg_0527 <= op1_03_out;
    18: reg_0527 <= op1_03_out;
    20: reg_0527 <= op1_03_out;
    23: reg_0527 <= imem01_in[83:80];
    24: reg_0527 <= op2_00_out;
    26: reg_0527 <= op2_00_out;
    33: reg_0527 <= op2_00_out;
    56: reg_0527 <= op2_00_out;
    88: reg_0527 <= op2_00_out;
    endcase
  end

  // REG#528の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0528 <= imem04_in[43:40];
    16: reg_0528 <= imem05_in[63:60];
    18: reg_0528 <= imem04_in[43:40];
    47: reg_0528 <= imem06_in[27:24];
    49: reg_0528 <= imem04_in[43:40];
    60: reg_0528 <= imem04_in[43:40];
    62: reg_0528 <= imem07_in[107:104];
    64: reg_0528 <= imem04_in[43:40];
    66: reg_0528 <= imem04_in[43:40];
    68: reg_0528 <= imem05_in[63:60];
    74: reg_0528 <= imem05_in[63:60];
    97: reg_0528 <= imem07_in[107:104];
    endcase
  end

  // REG#529の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0529 <= imem04_in[55:52];
    19: reg_0529 <= imem05_in[67:64];
    22: reg_0529 <= imem04_in[55:52];
    25: reg_0529 <= imem02_in[67:64];
    28: reg_0529 <= imem04_in[99:96];
    30: reg_0529 <= imem02_in[67:64];
    32: reg_0529 <= imem05_in[71:68];
    34: reg_0529 <= imem05_in[71:68];
    36: reg_0529 <= imem04_in[55:52];
    38: reg_0529 <= imem05_in[71:68];
    41: reg_0529 <= imem07_in[87:84];
    43: reg_0529 <= imem05_in[71:68];
    45: reg_0529 <= imem05_in[71:68];
    47: reg_0529 <= imem05_in[71:68];
    49: reg_0529 <= imem04_in[55:52];
    59: reg_0529 <= imem07_in[87:84];
    61: reg_0529 <= imem07_in[87:84];
    63: reg_0529 <= imem05_in[71:68];
    65: reg_0529 <= imem04_in[55:52];
    67: reg_0529 <= imem07_in[87:84];
    69: reg_0529 <= imem07_in[87:84];
    71: reg_0529 <= imem04_in[99:96];
    73: reg_0529 <= imem07_in[87:84];
    75: reg_0529 <= imem07_in[87:84];
    80: reg_0529 <= imem05_in[71:68];
    82: reg_0529 <= imem07_in[87:84];
    endcase
  end

  // REG#530の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0530 <= imem04_in[23:20];
    19: reg_0530 <= imem05_in[115:112];
    22: reg_0530 <= imem05_in[115:112];
    24: reg_0530 <= imem04_in[23:20];
    78: reg_0530 <= imem05_in[115:112];
    82: reg_0530 <= imem04_in[23:20];
    85: reg_0530 <= imem04_in[23:20];
    87: reg_0530 <= imem05_in[115:112];
    endcase
  end

  // REG#531の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0531 <= imem04_in[115:112];
    20: reg_0531 <= imem01_in[55:52];
    22: reg_0531 <= imem06_in[83:80];
    24: reg_0531 <= imem00_in[47:44];
    26: reg_0531 <= imem06_in[83:80];
    28: reg_0531 <= imem00_in[47:44];
    30: reg_0531 <= imem03_in[7:4];
    33: reg_0531 <= imem00_in[47:44];
    35: reg_0531 <= imem00_in[47:44];
    37: reg_0531 <= imem06_in[83:80];
    57: reg_0531 <= imem01_in[55:52];
    59: reg_0531 <= imem04_in[115:112];
    86: reg_0531 <= imem01_in[55:52];
    88: reg_0531 <= imem06_in[83:80];
    90: reg_0531 <= imem06_in[83:80];
    92: reg_0531 <= imem06_in[83:80];
    94: reg_0531 <= imem06_in[83:80];
    endcase
  end

  // REG#532の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0532 <= imem04_in[95:92];
    20: reg_0532 <= imem01_in[59:56];
    22: reg_0532 <= imem04_in[95:92];
    24: reg_0532 <= imem01_in[59:56];
    27: reg_0532 <= imem03_in[11:8];
    30: reg_0532 <= imem03_in[103:100];
    33: reg_0532 <= imem03_in[103:100];
    35: reg_0532 <= imem03_in[103:100];
    37: reg_0532 <= imem07_in[83:80];
    39: reg_0532 <= imem07_in[83:80];
    41: reg_0532 <= imem03_in[103:100];
    43: reg_0532 <= imem07_in[83:80];
    93: reg_0532 <= imem07_in[83:80];
    95: reg_0532 <= imem03_in[11:8];
    endcase
  end

  // REG#533の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0533 <= imem04_in[107:104];
    20: reg_0533 <= imem02_in[55:52];
    22: reg_0533 <= imem04_in[107:104];
    25: reg_0533 <= imem02_in[55:52];
    27: reg_0533 <= imem02_in[55:52];
    30: reg_0533 <= imem04_in[107:104];
    32: reg_0533 <= imem02_in[55:52];
    34: reg_0533 <= imem03_in[91:88];
    36: reg_0533 <= imem06_in[51:48];
    39: reg_0533 <= imem06_in[51:48];
    58: reg_0533 <= imem06_in[51:48];
    82: reg_0533 <= imem03_in[91:88];
    84: reg_0533 <= imem06_in[51:48];
    86: reg_0533 <= imem06_in[51:48];
    endcase
  end

  // REG#534の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0534 <= imem04_in[51:48];
    20: reg_0534 <= imem04_in[51:48];
    22: reg_0534 <= imem04_in[51:48];
    25: reg_0534 <= imem04_in[51:48];
    27: reg_0534 <= imem04_in[51:48];
    30: reg_0534 <= imem04_in[51:48];
    32: reg_0534 <= imem00_in[59:56];
    34: reg_0534 <= imem03_in[107:104];
    36: reg_0534 <= imem06_in[11:8];
    39: reg_0534 <= imem06_in[11:8];
    58: reg_0534 <= imem06_in[11:8];
    87: reg_0534 <= imem02_in[95:92];
    89: reg_0534 <= imem04_in[51:48];
    91: reg_0534 <= imem04_in[51:48];
    93: reg_0534 <= imem04_in[51:48];
    95: reg_0534 <= imem00_in[59:56];
    endcase
  end

  // REG#535の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0535 <= imem04_in[59:56];
    20: reg_0535 <= imem02_in[107:104];
    23: reg_0535 <= imem04_in[59:56];
    25: reg_0535 <= imem04_in[59:56];
    27: reg_0535 <= imem03_in[15:12];
    29: reg_0535 <= imem04_in[59:56];
    31: reg_0535 <= imem03_in[15:12];
    55: reg_0535 <= imem03_in[15:12];
    89: reg_0535 <= imem04_in[59:56];
    91: reg_0535 <= imem04_in[59:56];
    93: reg_0535 <= imem04_in[59:56];
    endcase
  end

  // REG#536の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0536 <= imem04_in[15:12];
    21: reg_0536 <= imem04_in[15:12];
    24: reg_0536 <= imem04_in[15:12];
    84: reg_0536 <= imem02_in[27:24];
    endcase
  end

  // REG#537の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0537 <= imem04_in[71:68];
    21: reg_0537 <= imem04_in[123:120];
    24: reg_0537 <= imem04_in[123:120];
    83: reg_0537 <= imem04_in[123:120];
    endcase
  end

  // REG#538の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0538 <= op1_04_out;
    20: reg_0538 <= op1_04_out;
    22: reg_0538 <= op1_04_out;
    24: reg_0538 <= op1_04_out;
    26: reg_0538 <= op1_04_out;
    28: reg_0538 <= op1_04_out;
    30: reg_0538 <= op1_04_out;
    32: reg_0538 <= op1_04_out;
    34: reg_0538 <= op1_04_out;
    36: reg_0538 <= op1_04_out;
    38: reg_0538 <= op1_04_out;
    40: reg_0538 <= op1_04_out;
    42: reg_0538 <= op1_04_out;
    44: reg_0538 <= op1_04_out;
    46: reg_0538 <= op1_04_out;
    48: reg_0538 <= op1_04_out;
    50: reg_0538 <= op1_04_out;
    52: reg_0538 <= op1_04_out;
    54: reg_0538 <= op1_04_out;
    56: reg_0538 <= op1_04_out;
    58: reg_0538 <= op1_04_out;
    60: reg_0538 <= op1_04_out;
    62: reg_0538 <= op1_04_out;
    64: reg_0538 <= op1_04_out;
    66: reg_0538 <= op1_04_out;
    68: reg_0538 <= op1_04_out;
    70: reg_0538 <= op1_04_out;
    72: reg_0538 <= op1_04_out;
    74: reg_0538 <= op1_04_out;
    76: reg_0538 <= op1_04_out;
    78: reg_0538 <= op1_04_out;
    80: reg_0538 <= op1_04_out;
    82: reg_0538 <= op1_04_out;
    84: reg_0538 <= op1_04_out;
    86: reg_0538 <= op1_04_out;
    88: reg_0538 <= op1_04_out;
    90: reg_0538 <= op1_04_out;
    92: reg_0538 <= op1_04_out;
    94: reg_0538 <= op1_04_out;
    96: reg_0538 <= op1_04_out;
    endcase
  end

  // REG#539の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0539 <= imem04_in[63:60];
    22: reg_0539 <= imem07_in[67:64];
    24: reg_0539 <= imem04_in[63:60];
    82: reg_0539 <= imem07_in[67:64];
    endcase
  end

  // REG#540の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0540 <= imem04_in[91:88];
    22: reg_0540 <= imem01_in[111:108];
    24: reg_0540 <= imem04_in[91:88];
    83: reg_0540 <= imem04_in[91:88];
    97: reg_0540 <= imem01_in[111:108];
    endcase
  end

  // REG#541の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0541 <= imem04_in[119:116];
    22: reg_0541 <= imem01_in[127:124];
    24: reg_0541 <= imem04_in[119:116];
    80: reg_0541 <= imem01_in[11:8];
    82: reg_0541 <= imem04_in[119:116];
    85: reg_0541 <= imem04_in[119:116];
    87: reg_0541 <= imem04_in[119:116];
    89: reg_0541 <= imem01_in[127:124];
    92: reg_0541 <= imem01_in[11:8];
    endcase
  end

  // REG#542の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0542 <= imem04_in[47:44];
    22: reg_0542 <= imem04_in[47:44];
    24: reg_0542 <= imem00_in[71:68];
    26: reg_0542 <= imem00_in[67:64];
    28: reg_0542 <= imem00_in[71:68];
    30: reg_0542 <= imem00_in[71:68];
    32: reg_0542 <= imem01_in[51:48];
    34: reg_0542 <= imem04_in[47:44];
    36: reg_0542 <= imem06_in[23:20];
    39: reg_0542 <= imem04_in[47:44];
    41: reg_0542 <= imem04_in[47:44];
    43: reg_0542 <= imem04_in[47:44];
    45: reg_0542 <= imem04_in[47:44];
    48: reg_0542 <= imem06_in[23:20];
    50: reg_0542 <= imem01_in[51:48];
    53: reg_0542 <= imem04_in[47:44];
    55: reg_0542 <= imem04_in[47:44];
    57: reg_0542 <= imem04_in[91:88];
    59: reg_0542 <= imem04_in[91:88];
    endcase
  end

  // REG#543の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0543 <= imem04_in[3:0];
    23: reg_0543 <= imem04_in[3:0];
    26: reg_0543 <= imem03_in[27:24];
    28: reg_0543 <= imem03_in[27:24];
    72: reg_0543 <= imem04_in[3:0];
    74: reg_0543 <= imem03_in[27:24];
    76: reg_0543 <= imem02_in[35:32];
    78: reg_0543 <= imem02_in[35:32];
    80: reg_0543 <= imem04_in[3:0];
    82: reg_0543 <= imem02_in[35:32];
    84: reg_0543 <= imem02_in[35:32];
    endcase
  end

  // REG#544の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0544 <= imem04_in[7:4];
    23: reg_0544 <= imem01_in[95:92];
    25: reg_0544 <= imem01_in[95:92];
    48: reg_0544 <= imem01_in[95:92];
    49: reg_0544 <= op2_00_out;
    68: reg_0544 <= imem01_in[95:92];
    70: reg_0544 <= op2_00_out;
    92: reg_0544 <= imem01_in[95:92];
    97: reg_0544 <= op2_00_out;
    endcase
  end

  // REG#545の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0545 <= imem04_in[11:8];
    23: reg_0545 <= imem04_in[11:8];
    25: reg_0545 <= imem02_in[71:68];
    28: reg_0545 <= imem06_in[107:104];
    31: reg_0545 <= imem06_in[107:104];
    33: reg_0545 <= imem04_in[99:96];
    35: reg_0545 <= imem04_in[99:96];
    37: reg_0545 <= imem06_in[107:104];
    61: reg_0545 <= imem02_in[71:68];
    63: reg_0545 <= imem04_in[11:8];
    65: reg_0545 <= imem04_in[99:96];
    67: reg_0545 <= imem04_in[99:96];
    69: reg_0545 <= imem02_in[71:68];
    71: reg_0545 <= imem06_in[107:104];
    89: reg_0545 <= imem02_in[71:68];
    91: reg_0545 <= imem04_in[99:96];
    93: reg_0545 <= imem07_in[87:84];
    95: reg_0545 <= imem04_in[99:96];
    endcase
  end

  // REG#546の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0546 <= imem04_in[87:84];
    23: reg_0546 <= imem04_in[87:84];
    26: reg_0546 <= imem04_in[87:84];
    28: reg_0546 <= imem04_in[87:84];
    30: reg_0546 <= imem04_in[87:84];
    32: reg_0546 <= imem01_in[59:56];
    34: reg_0546 <= imem01_in[59:56];
    36: reg_0546 <= imem04_in[87:84];
    38: reg_0546 <= imem01_in[59:56];
    41: reg_0546 <= imem04_in[87:84];
    43: reg_0546 <= imem01_in[59:56];
    45: reg_0546 <= imem04_in[87:84];
    48: reg_0546 <= imem01_in[59:56];
    49: reg_0546 <= op2_01_out;
    69: reg_0546 <= imem01_in[59:56];
    89: reg_0546 <= op2_01_out;
    endcase
  end

  // REG#547の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0547 <= imem04_in[127:124];
    23: reg_0547 <= imem03_in[95:92];
    25: reg_0547 <= imem02_in[99:96];
    28: reg_0547 <= imem04_in[127:124];
    30: reg_0547 <= imem02_in[99:96];
    32: reg_0547 <= imem03_in[95:92];
    34: reg_0547 <= imem03_in[95:92];
    36: reg_0547 <= imem03_in[95:92];
    38: reg_0547 <= imem02_in[99:96];
    41: reg_0547 <= imem03_in[95:92];
    43: reg_0547 <= imem06_in[103:100];
    45: reg_0547 <= imem04_in[127:124];
    48: reg_0547 <= imem04_in[127:124];
    51: reg_0547 <= imem02_in[99:96];
    55: reg_0547 <= imem03_in[95:92];
    88: reg_0547 <= imem04_in[127:124];
    90: reg_0547 <= imem03_in[95:92];
    endcase
  end

  // REG#548の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0548 <= imem04_in[67:64];
    23: reg_0548 <= imem04_in[67:64];
    26: reg_0548 <= imem04_in[43:40];
    28: reg_0548 <= imem04_in[43:40];
    29: reg_0548 <= op2_02_out;
    46: reg_0548 <= imem04_in[43:40];
    47: reg_0548 <= op2_02_out;
    62: reg_0548 <= op2_02_out;
    67: reg_0548 <= op2_02_out;
    83: reg_0548 <= op2_02_out;
    93: reg_0548 <= op2_02_out;
    endcase
  end

  // REG#549の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0549 <= imem04_in[79:76];
    23: reg_0549 <= imem04_in[79:76];
    24: reg_0549 <= op2_01_out;
    27: reg_0549 <= op2_01_out;
    37: reg_0549 <= op2_01_out;
    70: reg_0549 <= op2_01_out;
    92: reg_0549 <= op2_01_out;
    endcase
  end

  // REG#550の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0550 <= imem04_in[35:32];
    23: reg_0550 <= imem04_in[35:32];
    26: reg_0550 <= imem04_in[95:92];
    28: reg_0550 <= imem04_in[35:32];
    30: reg_0550 <= imem04_in[35:32];
    32: reg_0550 <= imem04_in[35:32];
    34: reg_0550 <= imem04_in[35:32];
    36: reg_0550 <= imem04_in[95:92];
    38: reg_0550 <= imem04_in[95:92];
    41: reg_0550 <= imem04_in[35:32];
    43: reg_0550 <= imem06_in[119:116];
    44: reg_0550 <= op1_10_out;
    46: reg_0550 <= op1_10_out;
    48: reg_0550 <= op1_10_out;
    50: reg_0550 <= op1_10_out;
    52: reg_0550 <= op1_10_out;
    54: reg_0550 <= op1_10_out;
    56: reg_0550 <= op1_10_out;
    58: reg_0550 <= op1_10_out;
    60: reg_0550 <= op1_10_out;
    63: reg_0550 <= imem04_in[95:92];
    65: reg_0550 <= imem04_in[95:92];
    67: reg_0550 <= imem04_in[95:92];
    69: reg_0550 <= imem04_in[95:92];
    70: reg_0550 <= op1_10_out;
    72: reg_0550 <= op1_10_out;
    74: reg_0550 <= op1_10_out;
    76: reg_0550 <= op1_10_out;
    78: reg_0550 <= op1_10_out;
    80: reg_0550 <= op1_10_out;
    83: reg_0550 <= imem04_in[35:32];
    endcase
  end

  // REG#551の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0551 <= imem04_in[103:100];
    23: reg_0551 <= imem03_in[127:124];
    25: reg_0551 <= imem03_in[127:124];
    27: reg_0551 <= imem03_in[127:124];
    31: reg_0551 <= imem04_in[103:100];
    33: reg_0551 <= imem03_in[127:124];
    35: reg_0551 <= imem03_in[119:116];
    37: reg_0551 <= imem03_in[119:116];
    39: reg_0551 <= imem04_in[103:100];
    41: reg_0551 <= imem03_in[127:124];
    43: reg_0551 <= imem02_in[39:36];
    45: reg_0551 <= imem04_in[103:100];
    48: reg_0551 <= imem03_in[127:124];
    49: reg_0551 <= op2_02_out;
    70: reg_0551 <= imem03_in[127:124];
    95: reg_0551 <= imem03_in[119:116];
    96: reg_0551 <= op2_02_out;
    endcase
  end

  // REG#552の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0552 <= imem04_in[39:36];
    23: reg_0552 <= imem04_in[119:116];
    25: reg_0552 <= imem04_in[39:36];
    27: reg_0552 <= imem03_in[95:92];
    30: reg_0552 <= imem03_in[95:92];
    32: reg_0552 <= imem04_in[39:36];
    34: reg_0552 <= imem04_in[39:36];
    36: reg_0552 <= imem04_in[39:36];
    38: reg_0552 <= imem04_in[39:36];
    41: reg_0552 <= imem04_in[39:36];
    43: reg_0552 <= imem04_in[39:36];
    45: reg_0552 <= imem04_in[39:36];
    47: reg_0552 <= imem07_in[63:60];
    49: reg_0552 <= imem03_in[95:92];
    51: reg_0552 <= imem04_in[39:36];
    53: reg_0552 <= imem03_in[95:92];
    57: reg_0552 <= imem04_in[119:116];
    59: reg_0552 <= imem04_in[39:36];
    endcase
  end

  // REG#553の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0553 <= imem04_in[31:28];
    23: reg_0553 <= imem05_in[119:116];
    24: reg_0553 <= op2_02_out;
    28: reg_0553 <= op2_02_out;
    42: reg_0553 <= op2_02_out;
    46: reg_0553 <= op2_02_out;
    60: reg_0553 <= imem04_in[31:28];
    62: reg_0553 <= imem00_in[83:80];
    63: reg_0553 <= op2_02_out;
    72: reg_0553 <= imem04_in[31:28];
    73: reg_0553 <= op2_02_out;
    endcase
  end

  // REG#554の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0554 <= imem04_in[83:80];
    23: reg_0554 <= imem04_in[83:80];
    26: reg_0554 <= imem04_in[83:80];
    28: reg_0554 <= imem06_in[123:120];
    31: reg_0554 <= imem02_in[67:64];
    33: reg_0554 <= imem04_in[123:120];
    35: reg_0554 <= imem04_in[35:32];
    37: reg_0554 <= imem07_in[107:104];
    39: reg_0554 <= imem04_in[123:120];
    41: reg_0554 <= imem04_in[123:120];
    43: reg_0554 <= imem04_in[123:120];
    45: reg_0554 <= imem04_in[123:120];
    47: reg_0554 <= imem04_in[123:120];
    49: reg_0554 <= imem04_in[35:32];
    60: reg_0554 <= imem04_in[35:32];
    62: reg_0554 <= imem04_in[123:120];
    64: reg_0554 <= imem04_in[35:32];
    66: reg_0554 <= imem07_in[107:104];
    68: reg_0554 <= imem06_in[123:120];
    70: reg_0554 <= imem04_in[123:120];
    72: reg_0554 <= imem04_in[123:120];
    74: reg_0554 <= imem06_in[123:120];
    76: reg_0554 <= imem02_in[67:64];
    78: reg_0554 <= imem04_in[83:80];
    80: reg_0554 <= imem04_in[35:32];
    82: reg_0554 <= imem02_in[67:64];
    84: reg_0554 <= imem02_in[67:64];
    94: reg_0554 <= imem02_in[67:64];
    96: reg_0554 <= imem04_in[123:120];
    endcase
  end

  // REG#555の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0555 <= imem04_in[75:72];
    23: reg_0555 <= imem06_in[127:124];
    25: reg_0555 <= imem01_in[63:60];
    46: reg_0555 <= imem01_in[63:60];
    48: reg_0555 <= imem04_in[95:92];
    51: reg_0555 <= imem04_in[75:72];
    53: reg_0555 <= imem01_in[63:60];
    endcase
  end

  // REG#556の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0556 <= imem04_in[123:120];
    23: reg_0556 <= imem04_in[123:120];
    26: reg_0556 <= imem04_in[119:116];
    28: reg_0556 <= imem06_in[103:100];
    31: reg_0556 <= imem06_in[103:100];
    34: reg_0556 <= imem04_in[119:116];
    36: reg_0556 <= imem06_in[75:72];
    39: reg_0556 <= imem06_in[75:72];
    58: reg_0556 <= imem06_in[75:72];
    86: reg_0556 <= imem04_in[119:116];
    88: reg_0556 <= imem06_in[103:100];
    91: reg_0556 <= imem06_in[103:100];
    93: reg_0556 <= imem06_in[103:100];
    95: reg_0556 <= imem04_in[119:116];
    97: reg_0556 <= imem04_in[119:116];
    endcase
  end

  // REG#557の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0557 <= imem04_in[19:16];
    23: reg_0557 <= imem04_in[19:16];
    26: reg_0557 <= imem04_in[19:16];
    28: reg_0557 <= imem06_in[91:88];
    31: reg_0557 <= imem04_in[19:16];
    33: reg_0557 <= imem07_in[39:36];
    35: reg_0557 <= imem04_in[19:16];
    37: reg_0557 <= imem07_in[115:112];
    39: reg_0557 <= imem04_in[19:16];
    41: reg_0557 <= imem04_in[19:16];
    43: reg_0557 <= op2_02_out;
    50: reg_0557 <= imem07_in[39:36];
    51: reg_0557 <= op2_02_out;
    75: reg_0557 <= op2_02_out;
    endcase
  end

  // REG#558の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0558 <= imem04_in[99:96];
    23: reg_0558 <= imem07_in[23:20];
    25: reg_0558 <= imem07_in[23:20];
    27: reg_0558 <= imem03_in[111:108];
    30: reg_0558 <= imem07_in[23:20];
    32: reg_0558 <= imem07_in[23:20];
    34: reg_0558 <= imem03_in[111:108];
    36: reg_0558 <= imem06_in[63:60];
    41: reg_0558 <= imem07_in[23:20];
    43: reg_0558 <= imem02_in[123:120];
    45: reg_0558 <= imem02_in[123:120];
    61: reg_0558 <= imem04_in[99:96];
    63: reg_0558 <= imem06_in[63:60];
    65: reg_0558 <= imem07_in[23:20];
    67: reg_0558 <= imem07_in[23:20];
    69: reg_0558 <= imem06_in[63:60];
    71: reg_0558 <= imem02_in[123:120];
    74: reg_0558 <= imem06_in[63:60];
    76: reg_0558 <= imem03_in[111:108];
    78: reg_0558 <= imem03_in[111:108];
    80: reg_0558 <= imem03_in[111:108];
    82: reg_0558 <= imem01_in[35:32];
    84: reg_0558 <= imem07_in[23:20];
    86: reg_0558 <= imem07_in[23:20];
    88: reg_0558 <= imem03_in[111:108];
    endcase
  end

  // REG#559の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0559 <= imem04_in[111:108];
    23: reg_0559 <= imem04_in[111:108];
    25: reg_0559 <= op2_01_out;
    30: reg_0559 <= op2_01_out;
    47: reg_0559 <= op2_01_out;
    61: reg_0559 <= op2_01_out;
    65: reg_0559 <= imem04_in[111:108];
    66: reg_0559 <= op2_01_out;
    79: reg_0559 <= op2_01_out;
    endcase
  end

  // REG#560の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0560 <= imem04_in[27:24];
    23: reg_0560 <= imem04_in[27:24];
    25: reg_0560 <= imem01_in[23:20];
    47: reg_0560 <= imem01_in[23:20];
    52: reg_0560 <= imem01_in[23:20];
    55: reg_0560 <= imem04_in[27:24];
    57: reg_0560 <= imem07_in[67:64];
    59: reg_0560 <= imem07_in[67:64];
    61: reg_0560 <= imem01_in[23:20];
    63: reg_0560 <= imem04_in[27:24];
    65: reg_0560 <= imem07_in[67:64];
    68: reg_0560 <= imem07_in[67:64];
    70: reg_0560 <= imem07_in[67:64];
    72: reg_0560 <= imem07_in[67:64];
    74: reg_0560 <= imem01_in[23:20];
    76: reg_0560 <= imem01_in[23:20];
    79: reg_0560 <= imem07_in[67:64];
    endcase
  end

  // REG#561の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0561 <= op1_05_out;
    22: reg_0561 <= op1_05_out;
    24: reg_0561 <= op1_05_out;
    27: reg_0561 <= imem03_in[31:28];
    30: reg_0561 <= imem03_in[31:28];
    33: reg_0561 <= imem03_in[31:28];
    35: reg_0561 <= imem05_in[3:0];
    36: reg_0561 <= op2_02_out;
    68: reg_0561 <= op2_02_out;
    86: reg_0561 <= op2_02_out;
    endcase
  end

  // REG#562の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0562 <= op1_06_out;
    22: reg_0562 <= op1_06_out;
    24: reg_0562 <= op1_06_out;
    26: reg_0562 <= op1_06_out;
    28: reg_0562 <= op1_06_out;
    30: reg_0562 <= op1_06_out;
    32: reg_0562 <= op1_06_out;
    34: reg_0562 <= op1_06_out;
    36: reg_0562 <= op1_06_out;
    38: reg_0562 <= op1_06_out;
    40: reg_0562 <= op1_06_out;
    42: reg_0562 <= op1_06_out;
    44: reg_0562 <= op1_06_out;
    46: reg_0562 <= op1_06_out;
    48: reg_0562 <= op1_06_out;
    50: reg_0562 <= op1_06_out;
    52: reg_0562 <= op1_06_out;
    54: reg_0562 <= op1_06_out;
    56: reg_0562 <= op1_06_out;
    58: reg_0562 <= op1_06_out;
    60: reg_0562 <= op1_06_out;
    62: reg_0562 <= op1_06_out;
    64: reg_0562 <= op1_06_out;
    66: reg_0562 <= op1_06_out;
    68: reg_0562 <= op1_06_out;
    70: reg_0562 <= op1_06_out;
    72: reg_0562 <= op1_06_out;
    74: reg_0562 <= op1_06_out;
    76: reg_0562 <= op1_06_out;
    78: reg_0562 <= op1_06_out;
    80: reg_0562 <= op1_06_out;
    82: reg_0562 <= op1_06_out;
    84: reg_0562 <= op1_06_out;
    86: reg_0562 <= op1_06_out;
    88: reg_0562 <= op1_06_out;
    90: reg_0562 <= op1_06_out;
    92: reg_0562 <= op1_06_out;
    94: reg_0562 <= op1_06_out;
    96: reg_0562 <= op1_06_out;
    endcase
  end

  // REG#563の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0563 <= imem03_in[67:64];
    25: reg_0563 <= imem01_in[27:24];
    47: reg_0563 <= imem03_in[67:64];
    49: reg_0563 <= imem03_in[67:64];
    51: reg_0563 <= imem03_in[67:64];
    53: reg_0563 <= imem07_in[107:104];
    55: reg_0563 <= imem05_in[11:8];
    57: reg_0563 <= imem00_in[7:4];
    59: reg_0563 <= imem05_in[11:8];
    61: reg_0563 <= imem00_in[7:4];
    63: reg_0563 <= imem07_in[107:104];
    65: reg_0563 <= imem03_in[67:64];
    67: reg_0563 <= imem00_in[7:4];
    69: reg_0563 <= imem03_in[67:64];
    71: reg_0563 <= imem05_in[11:8];
    73: reg_0563 <= imem01_in[27:24];
    75: reg_0563 <= imem07_in[107:104];
    79: reg_0563 <= imem07_in[107:104];
    endcase
  end

  // REG#564の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0564 <= op1_07_out;
    24: reg_0564 <= op1_07_out;
    26: reg_0564 <= op1_07_out;
    29: reg_0564 <= op1_07_out;
    31: reg_0564 <= op1_07_out;
    33: reg_0564 <= op1_07_out;
    35: reg_0564 <= op1_07_out;
    37: reg_0564 <= op1_07_out;
    39: reg_0564 <= op1_07_out;
    41: reg_0564 <= op1_07_out;
    43: reg_0564 <= op1_07_out;
    45: reg_0564 <= op1_07_out;
    47: reg_0564 <= op1_07_out;
    49: reg_0564 <= op1_07_out;
    51: reg_0564 <= op1_07_out;
    53: reg_0564 <= op1_07_out;
    55: reg_0564 <= op1_07_out;
    57: reg_0564 <= op1_07_out;
    59: reg_0564 <= op1_07_out;
    61: reg_0564 <= op1_07_out;
    63: reg_0564 <= op1_07_out;
    65: reg_0564 <= op1_07_out;
    67: reg_0564 <= op1_07_out;
    69: reg_0564 <= op1_07_out;
    71: reg_0564 <= op1_07_out;
    73: reg_0564 <= op1_07_out;
    75: reg_0564 <= op1_07_out;
    77: reg_0564 <= op1_07_out;
    79: reg_0564 <= op1_07_out;
    81: reg_0564 <= op1_07_out;
    83: reg_0564 <= op1_07_out;
    85: reg_0564 <= op1_07_out;
    87: reg_0564 <= op1_07_out;
    89: reg_0564 <= op1_07_out;
    91: reg_0564 <= op1_07_out;
    93: reg_0564 <= op1_07_out;
    95: reg_0564 <= op1_07_out;
    97: reg_0564 <= op1_07_out;
    endcase
  end

  // REG#565の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0565 <= op1_08_out;
    24: reg_0565 <= op1_08_out;
    26: reg_0565 <= op1_08_out;
    28: reg_0565 <= op1_08_out;
    31: reg_0565 <= imem02_in[87:84];
    33: reg_0565 <= imem07_in[75:72];
    35: reg_0565 <= imem05_in[23:20];
    37: reg_0565 <= imem07_in[75:72];
    39: reg_0565 <= imem07_in[75:72];
    41: reg_0565 <= imem05_in[23:20];
    43: reg_0565 <= imem02_in[87:84];
    45: reg_0565 <= imem02_in[87:84];
    63: reg_0565 <= imem02_in[87:84];
    71: reg_0565 <= op1_08_out;
    73: reg_0565 <= op1_08_out;
    75: reg_0565 <= op1_08_out;
    77: reg_0565 <= op1_08_out;
    79: reg_0565 <= op1_08_out;
    82: reg_0565 <= imem07_in[75:72];
    endcase
  end

  // REG#566の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0566 <= op1_09_out;
    27: reg_0566 <= op1_09_out;
    29: reg_0566 <= op1_09_out;
    32: reg_0566 <= imem02_in[63:60];
    34: reg_0566 <= imem02_in[63:60];
    36: reg_0566 <= imem06_in[115:112];
    40: reg_0566 <= imem02_in[63:60];
    42: reg_0566 <= imem02_in[63:60];
    45: reg_0566 <= imem06_in[115:112];
    46: reg_0566 <= op1_09_out;
    49: reg_0566 <= imem06_in[115:112];
    51: reg_0566 <= imem02_in[63:60];
    54: reg_0566 <= imem06_in[115:112];
    56: reg_0566 <= imem06_in[115:112];
    58: reg_0566 <= op1_09_out;
    60: reg_0566 <= op1_09_out;
    62: reg_0566 <= op1_09_out;
    64: reg_0566 <= op1_09_out;
    66: reg_0566 <= op1_09_out;
    69: reg_0566 <= imem02_in[63:60];
    71: reg_0566 <= imem06_in[115:112];
    82: reg_0566 <= op1_09_out;
    84: reg_0566 <= op1_09_out;
    86: reg_0566 <= op1_09_out;
    89: reg_0566 <= imem06_in[115:112];
    96: reg_0566 <= op1_09_out;
    endcase
  end

  // REG#567の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0567 <= op1_10_out;
    27: reg_0567 <= op1_10_out;
    29: reg_0567 <= op1_10_out;
    31: reg_0567 <= op1_10_out;
    34: reg_0567 <= imem07_in[11:8];
    36: reg_0567 <= imem07_in[11:8];
    38: reg_0567 <= imem03_in[87:84];
    40: reg_0567 <= op1_10_out;
    42: reg_0567 <= op1_10_out;
    45: reg_0567 <= imem07_in[11:8];
    47: reg_0567 <= imem00_in[79:76];
    49: reg_0567 <= imem07_in[11:8];
    53: reg_0567 <= imem03_in[87:84];
    57: reg_0567 <= imem03_in[87:84];
    59: reg_0567 <= imem03_in[87:84];
    61: reg_0567 <= imem03_in[87:84];
    62: reg_0567 <= op1_10_out;
    64: reg_0567 <= op1_10_out;
    66: reg_0567 <= op1_10_out;
    68: reg_0567 <= op1_10_out;
    72: reg_0567 <= imem00_in[79:76];
    74: reg_0567 <= imem07_in[11:8];
    77: reg_0567 <= imem03_in[87:84];
    79: reg_0567 <= imem07_in[11:8];
    96: reg_0567 <= op1_10_out;
    endcase
  end

  // REG#568の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0568 <= imem03_in[43:40];
    30: reg_0568 <= imem03_in[43:40];
    33: reg_0568 <= imem07_in[87:84];
    35: reg_0568 <= imem07_in[87:84];
    38: reg_0568 <= imem04_in[27:24];
    40: reg_0568 <= imem04_in[27:24];
    42: reg_0568 <= imem04_in[27:24];
    endcase
  end

  // REG#569の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0569 <= imem03_in[55:52];
    30: reg_0569 <= imem03_in[55:52];
    33: reg_0569 <= imem03_in[55:52];
    35: reg_0569 <= imem03_in[55:52];
    38: reg_0569 <= imem04_in[115:112];
    40: reg_0569 <= imem04_in[115:112];
    42: reg_0569 <= imem00_in[107:104];
    44: reg_0569 <= imem03_in[55:52];
    46: reg_0569 <= imem00_in[107:104];
    48: reg_0569 <= imem04_in[115:112];
    52: reg_0569 <= imem00_in[107:104];
    54: reg_0569 <= imem04_in[115:112];
    56: reg_0569 <= imem05_in[7:4];
    59: reg_0569 <= imem03_in[55:52];
    61: reg_0569 <= imem07_in[55:52];
    63: reg_0569 <= imem04_in[115:112];
    65: reg_0569 <= imem00_in[107:104];
    68: reg_0569 <= imem00_in[107:104];
    70: reg_0569 <= imem00_in[107:104];
    72: reg_0569 <= imem07_in[55:52];
    74: reg_0569 <= imem07_in[55:52];
    77: reg_0569 <= imem07_in[55:52];
    79: reg_0569 <= imem07_in[55:52];
    95: reg_0569 <= imem05_in[7:4];
    endcase
  end

  // REG#570の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0570 <= imem03_in[119:116];
    30: reg_0570 <= imem03_in[119:116];
    32: reg_0570 <= imem03_in[119:116];
    34: reg_0570 <= imem00_in[63:60];
    36: reg_0570 <= imem00_in[63:60];
    38: reg_0570 <= imem00_in[63:60];
    41: reg_0570 <= imem00_in[75:72];
    43: reg_0570 <= imem04_in[11:8];
    45: reg_0570 <= imem00_in[63:60];
    47: reg_0570 <= imem04_in[11:8];
    49: reg_0570 <= imem03_in[119:116];
    51: reg_0570 <= imem04_in[11:8];
    53: reg_0570 <= imem03_in[119:116];
    57: reg_0570 <= imem04_in[11:8];
    59: reg_0570 <= imem00_in[63:60];
    61: reg_0570 <= imem03_in[119:116];
    63: reg_0570 <= imem00_in[63:60];
    65: reg_0570 <= imem07_in[51:48];
    67: reg_0570 <= imem07_in[51:48];
    69: reg_0570 <= imem07_in[51:48];
    71: reg_0570 <= imem00_in[63:60];
    73: reg_0570 <= imem03_in[119:116];
    75: reg_0570 <= imem00_in[75:72];
    77: reg_0570 <= imem00_in[75:72];
    79: reg_0570 <= imem00_in[63:60];
    81: reg_0570 <= imem00_in[63:60];
    83: reg_0570 <= imem00_in[63:60];
    85: reg_0570 <= imem00_in[75:72];
    87: reg_0570 <= imem03_in[119:116];
    89: reg_0570 <= imem03_in[119:116];
    92: reg_0570 <= imem00_in[63:60];
    94: reg_0570 <= imem00_in[63:60];
    endcase
  end

  // REG#571の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0571 <= imem03_in[19:16];
    31: reg_0571 <= imem03_in[19:16];
    54: reg_0571 <= imem03_in[19:16];
    56: reg_0571 <= imem06_in[75:72];
    59: reg_0571 <= imem03_in[19:16];
    61: reg_0571 <= imem06_in[75:72];
    68: reg_0571 <= imem06_in[103:100];
    70: reg_0571 <= imem03_in[19:16];
    94: reg_0571 <= imem06_in[75:72];
    96: reg_0571 <= imem06_in[75:72];
    endcase
  end

  // REG#572の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0572 <= imem03_in[47:44];
    30: reg_0572 <= imem03_in[47:44];
    32: reg_0572 <= imem03_in[23:20];
    34: reg_0572 <= imem00_in[107:104];
    36: reg_0572 <= imem00_in[107:104];
    38: reg_0572 <= imem07_in[115:112];
    40: reg_0572 <= imem03_in[47:44];
    42: reg_0572 <= imem03_in[23:20];
    44: reg_0572 <= op1_12_out;
    47: reg_0572 <= imem03_in[47:44];
    48: reg_0572 <= op1_12_out;
    50: reg_0572 <= op1_12_out;
    53: reg_0572 <= imem00_in[11:8];
    55: reg_0572 <= imem03_in[47:44];
    89: reg_0572 <= imem07_in[115:112];
    91: reg_0572 <= imem00_in[11:8];
    endcase
  end

  // REG#573の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0573 <= imem03_in[23:20];
    31: reg_0573 <= imem03_in[23:20];
    52: reg_0573 <= imem03_in[23:20];
    54: reg_0573 <= imem03_in[23:20];
    56: reg_0573 <= imem06_in[111:108];
    60: reg_0573 <= imem06_in[111:108];
    63: reg_0573 <= imem07_in[83:80];
    65: reg_0573 <= imem07_in[83:80];
    67: reg_0573 <= imem03_in[23:20];
    69: reg_0573 <= imem06_in[111:108];
    71: reg_0573 <= imem06_in[111:108];
    89: reg_0573 <= imem03_in[23:20];
    92: reg_0573 <= imem07_in[83:80];
    94: reg_0573 <= imem07_in[83:80];
    endcase
  end

  // REG#574の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0574 <= op1_11_out;
    28: reg_0574 <= op1_11_out;
    30: reg_0574 <= op1_11_out;
    32: reg_0574 <= op1_11_out;
    35: reg_0574 <= imem05_in[87:84];
    37: reg_0574 <= op1_11_out;
    39: reg_0574 <= op1_11_out;
    41: reg_0574 <= op1_11_out;
    43: reg_0574 <= op1_11_out;
    45: reg_0574 <= op1_11_out;
    47: reg_0574 <= op1_11_out;
    49: reg_0574 <= op1_11_out;
    52: reg_0574 <= imem05_in[87:84];
    54: reg_0574 <= imem05_in[87:84];
    55: reg_0574 <= op1_11_out;
    57: reg_0574 <= op1_11_out;
    59: reg_0574 <= op1_11_out;
    61: reg_0574 <= op1_11_out;
    63: reg_0574 <= op1_11_out;
    65: reg_0574 <= op1_11_out;
    67: reg_0574 <= op1_11_out;
    69: reg_0574 <= op1_11_out;
    71: reg_0574 <= op1_11_out;
    73: reg_0574 <= op1_11_out;
    76: reg_0574 <= imem05_in[87:84];
    77: reg_0574 <= op1_11_out;
    79: reg_0574 <= op1_11_out;
    81: reg_0574 <= op1_11_out;
    85: reg_0574 <= imem00_in[19:16];
    87: reg_0574 <= imem03_in[123:120];
    90: reg_0574 <= op1_11_out;
    92: reg_0574 <= op1_11_out;
    95: reg_0574 <= imem03_in[123:120];
    96: reg_0574 <= op1_11_out;
    endcase
  end

  // REG#575の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0575 <= op1_12_out;
    28: reg_0575 <= op1_12_out;
    30: reg_0575 <= op1_12_out;
    32: reg_0575 <= op1_12_out;
    35: reg_0575 <= imem07_in[11:8];
    37: reg_0575 <= op1_12_out;
    40: reg_0575 <= op1_12_out;
    43: reg_0575 <= imem07_in[11:8];
    94: reg_0575 <= op1_12_out;
    96: reg_0575 <= op1_12_out;
    endcase
  end

  // REG#576の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0576 <= imem03_in[127:124];
    31: reg_0576 <= imem03_in[127:124];
    55: reg_0576 <= imem03_in[127:124];
    85: reg_0576 <= imem00_in[39:36];
    87: reg_0576 <= imem03_in[127:124];
    91: reg_0576 <= op2_01_out;
    endcase
  end

  // REG#577の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0577 <= imem06_in[95:92];
    31: reg_0577 <= imem04_in[7:4];
    33: reg_0577 <= imem04_in[7:4];
    35: reg_0577 <= imem06_in[95:92];
    39: reg_0577 <= imem06_in[95:92];
    53: reg_0577 <= imem06_in[95:92];
    55: reg_0577 <= imem03_in[75:72];
    83: reg_0577 <= imem04_in[7:4];
    96: reg_0577 <= imem03_in[75:72];
    endcase
  end

  // REG#578の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0578 <= imem03_in[99:96];
    31: reg_0578 <= imem04_in[87:84];
    33: reg_0578 <= imem04_in[87:84];
    35: reg_0578 <= imem00_in[27:24];
    37: reg_0578 <= imem04_in[87:84];
    39: reg_0578 <= imem03_in[67:64];
    41: reg_0578 <= imem00_in[123:120];
    43: reg_0578 <= imem00_in[123:120];
    45: reg_0578 <= imem03_in[67:64];
    47: reg_0578 <= imem03_in[99:96];
    49: reg_0578 <= imem04_in[87:84];
    60: reg_0578 <= imem00_in[27:24];
    62: reg_0578 <= imem01_in[3:0];
    64: reg_0578 <= imem00_in[27:24];
    66: reg_0578 <= imem00_in[27:24];
    68: reg_0578 <= imem00_in[27:24];
    70: reg_0578 <= imem00_in[27:24];
    72: reg_0578 <= imem04_in[87:84];
    74: reg_0578 <= imem03_in[67:64];
    76: reg_0578 <= imem00_in[27:24];
    78: reg_0578 <= imem03_in[99:96];
    80: reg_0578 <= imem00_in[27:24];
    82: reg_0578 <= imem00_in[27:24];
    84: reg_0578 <= imem00_in[27:24];
    86: reg_0578 <= imem01_in[3:0];
    88: reg_0578 <= imem03_in[67:64];
    endcase
  end

  // REG#579の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0579 <= imem03_in[35:32];
    31: reg_0579 <= imem05_in[107:104];
    33: reg_0579 <= imem03_in[35:32];
    35: reg_0579 <= imem03_in[35:32];
    38: reg_0579 <= imem00_in[79:76];
    41: reg_0579 <= imem04_in[91:88];
    45: reg_0579 <= imem04_in[119:116];
    48: reg_0579 <= imem03_in[35:32];
    50: reg_0579 <= imem04_in[91:88];
    52: reg_0579 <= imem05_in[107:104];
    54: reg_0579 <= imem04_in[119:116];
    56: reg_0579 <= imem04_in[119:116];
    58: reg_0579 <= imem04_in[119:116];
    61: reg_0579 <= imem04_in[91:88];
    63: reg_0579 <= imem05_in[107:104];
    65: reg_0579 <= imem03_in[35:32];
    67: reg_0579 <= imem05_in[107:104];
    70: reg_0579 <= imem03_in[35:32];
    94: reg_0579 <= imem04_in[119:116];
    endcase
  end

  // REG#580の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0580 <= imem03_in[95:92];
    31: reg_0580 <= imem03_in[95:92];
    55: reg_0580 <= imem03_in[55:52];
    85: reg_0580 <= imem00_in[123:120];
    87: reg_0580 <= imem03_in[55:52];
    89: reg_0580 <= imem03_in[95:92];
    91: reg_0580 <= imem00_in[123:120];
    endcase
  end

  // REG#581の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0581 <= imem03_in[107:104];
    31: reg_0581 <= imem03_in[107:104];
    52: reg_0581 <= imem03_in[107:104];
    54: reg_0581 <= imem03_in[107:104];
    56: reg_0581 <= imem05_in[23:20];
    60: reg_0581 <= imem03_in[107:104];
    62: reg_0581 <= imem03_in[107:104];
    64: reg_0581 <= imem05_in[23:20];
    67: reg_0581 <= imem05_in[23:20];
    70: reg_0581 <= imem03_in[107:104];
    endcase
  end

  // REG#582の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0582 <= imem03_in[15:12];
    32: reg_0582 <= imem03_in[67:64];
    34: reg_0582 <= imem01_in[3:0];
    36: reg_0582 <= imem03_in[67:64];
    38: reg_0582 <= imem01_in[27:24];
    40: reg_0582 <= imem03_in[15:12];
    42: reg_0582 <= imem02_in[55:52];
    44: reg_0582 <= imem02_in[55:52];
    45: reg_0582 <= op2_02_out;
    57: reg_0582 <= imem02_in[55:52];
    58: reg_0582 <= op2_02_out;
    97: reg_0582 <= op2_02_out;
    endcase
  end

  // REG#583の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0583 <= imem03_in[39:36];
    32: reg_0583 <= imem04_in[19:16];
    34: reg_0583 <= imem04_in[19:16];
    36: reg_0583 <= imem03_in[39:36];
    38: reg_0583 <= imem03_in[119:116];
    41: reg_0583 <= imem03_in[39:36];
    43: reg_0583 <= imem05_in[3:0];
    45: reg_0583 <= imem03_in[39:36];
    47: reg_0583 <= imem03_in[39:36];
    49: reg_0583 <= imem03_in[39:36];
    52: reg_0583 <= imem03_in[119:116];
    54: reg_0583 <= imem03_in[39:36];
    56: reg_0583 <= imem03_in[119:116];
    58: reg_0583 <= imem03_in[39:36];
    60: reg_0583 <= imem03_in[39:36];
    62: reg_0583 <= imem03_in[119:116];
    64: reg_0583 <= imem03_in[39:36];
    66: reg_0583 <= imem05_in[3:0];
    80: reg_0583 <= imem03_in[119:116];
    82: reg_0583 <= imem02_in[7:4];
    85: reg_0583 <= imem04_in[19:16];
    87: reg_0583 <= imem05_in[3:0];
    endcase
  end

  // REG#584の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0584 <= imem03_in[79:76];
    32: reg_0584 <= imem04_in[75:72];
    34: reg_0584 <= imem03_in[79:76];
    36: reg_0584 <= imem03_in[79:76];
    38: reg_0584 <= imem03_in[79:76];
    40: reg_0584 <= imem04_in[75:72];
    42: reg_0584 <= imem04_in[75:72];
    endcase
  end

  // REG#585の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0585 <= imem03_in[83:80];
    32: reg_0585 <= imem04_in[115:112];
    34: reg_0585 <= imem03_in[83:80];
    36: reg_0585 <= imem06_in[119:116];
    40: reg_0585 <= imem06_in[119:116];
    42: reg_0585 <= imem06_in[119:116];
    45: reg_0585 <= imem04_in[115:112];
    48: reg_0585 <= imem06_in[119:116];
    50: reg_0585 <= imem03_in[83:80];
    52: reg_0585 <= imem06_in[119:116];
    55: reg_0585 <= imem03_in[83:80];
    87: reg_0585 <= imem03_in[83:80];
    89: reg_0585 <= imem03_in[83:80];
    92: reg_0585 <= imem06_in[119:116];
    endcase
  end

  // REG#586の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0586 <= imem03_in[11:8];
    32: reg_0586 <= imem05_in[19:16];
    34: reg_0586 <= imem01_in[7:4];
    36: reg_0586 <= imem03_in[11:8];
    38: reg_0586 <= imem01_in[7:4];
    41: reg_0586 <= imem03_in[11:8];
    43: reg_0586 <= imem06_in[59:56];
    45: reg_0586 <= imem01_in[7:4];
    47: reg_0586 <= imem03_in[11:8];
    49: reg_0586 <= imem01_in[7:4];
    71: reg_0586 <= imem05_in[19:16];
    73: reg_0586 <= imem03_in[11:8];
    75: reg_0586 <= imem06_in[59:56];
    78: reg_0586 <= imem05_in[19:16];
    81: reg_0586 <= imem05_in[19:16];
    83: reg_0586 <= imem04_in[115:112];
    endcase
  end

  // REG#587の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0587 <= imem03_in[51:48];
    32: reg_0587 <= imem05_in[103:100];
    34: reg_0587 <= imem05_in[103:100];
    36: reg_0587 <= imem05_in[103:100];
    38: reg_0587 <= imem07_in[27:24];
    41: reg_0587 <= imem07_in[27:24];
    42: reg_0587 <= op2_01_out;
    45: reg_0587 <= op2_01_out;
    55: reg_0587 <= op2_01_out;
    87: reg_0587 <= imem05_in[103:100];
    95: reg_0587 <= op2_01_out;
    endcase
  end

  // REG#588の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0588 <= imem03_in[115:112];
    32: reg_0588 <= imem07_in[27:24];
    34: reg_0588 <= imem03_in[115:112];
    36: reg_0588 <= imem06_in[127:124];
    41: reg_0588 <= imem04_in[115:112];
    45: reg_0588 <= imem06_in[127:124];
    47: reg_0588 <= imem03_in[115:112];
    49: reg_0588 <= imem06_in[127:124];
    52: reg_0588 <= imem04_in[115:112];
    54: reg_0588 <= imem06_in[127:124];
    56: reg_0588 <= imem07_in[27:24];
    58: reg_0588 <= imem04_in[115:112];
    61: reg_0588 <= imem07_in[27:24];
    63: reg_0588 <= imem07_in[27:24];
    65: reg_0588 <= imem03_in[115:112];
    68: reg_0588 <= imem06_in[127:124];
    70: reg_0588 <= imem03_in[115:112];
    endcase
  end

  // REG#589の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0589 <= imem03_in[71:68];
    32: reg_0589 <= imem07_in[95:92];
    34: reg_0589 <= imem01_in[35:32];
    36: reg_0589 <= imem01_in[35:32];
    38: reg_0589 <= imem07_in[95:92];
    41: reg_0589 <= imem07_in[95:92];
    43: reg_0589 <= imem07_in[95:92];
    endcase
  end

  // REG#590の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0590 <= imem03_in[123:120];
    31: reg_0590 <= op1_03_out;
    34: reg_0590 <= imem03_in[123:120];
    35: reg_0590 <= op1_03_out;
    37: reg_0590 <= op1_03_out;
    39: reg_0590 <= op1_03_out;
    41: reg_0590 <= op1_03_out;
    43: reg_0590 <= op1_03_out;
    45: reg_0590 <= op1_03_out;
    48: reg_0590 <= imem03_in[123:120];
    51: reg_0590 <= op1_03_out;
    55: reg_0590 <= imem03_in[123:120];
    92: reg_0590 <= imem03_in[123:120];
    93: reg_0590 <= op1_03_out;
    95: reg_0590 <= op1_03_out;
    endcase
  end

  // REG#591の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0591 <= imem03_in[63:60];
    32: reg_0591 <= imem06_in[83:80];
    38: reg_0591 <= imem03_in[63:60];
    40: reg_0591 <= imem06_in[83:80];
    42: reg_0591 <= imem03_in[115:112];
    45: reg_0591 <= imem03_in[63:60];
    47: reg_0591 <= imem01_in[123:120];
    49: reg_0591 <= imem03_in[63:60];
    52: reg_0591 <= imem01_in[123:120];
    54: reg_0591 <= imem01_in[123:120];
    56: reg_0591 <= imem06_in[83:80];
    58: reg_0591 <= imem06_in[83:80];
    87: reg_0591 <= imem06_in[83:80];
    89: reg_0591 <= imem01_in[123:120];
    91: reg_0591 <= imem01_in[123:120];
    93: reg_0591 <= imem06_in[83:80];
    95: reg_0591 <= imem01_in[123:120];
    endcase
  end

  // REG#592の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0592 <= imem03_in[59:56];
    32: reg_0592 <= imem03_in[59:56];
    34: reg_0592 <= imem01_in[71:68];
    36: reg_0592 <= imem01_in[71:68];
    38: reg_0592 <= imem07_in[107:104];
    40: reg_0592 <= imem07_in[107:104];
    42: reg_0592 <= imem05_in[35:32];
    44: reg_0592 <= imem05_in[35:32];
    47: reg_0592 <= imem07_in[107:104];
    49: reg_0592 <= imem01_in[71:68];
    69: reg_0592 <= imem01_in[71:68];
    92: reg_0592 <= imem01_in[71:68];
    endcase
  end

  // REG#593の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0593 <= imem03_in[87:84];
    32: reg_0593 <= imem03_in[87:84];
    34: reg_0593 <= imem03_in[87:84];
    36: reg_0593 <= imem06_in[67:64];
    41: reg_0593 <= imem04_in[103:100];
    45: reg_0593 <= imem06_in[67:64];
    46: reg_0593 <= op1_12_out;
    49: reg_0593 <= imem04_in[103:100];
    60: reg_0593 <= imem06_in[7:4];
    63: reg_0593 <= imem03_in[87:84];
    65: reg_0593 <= imem04_in[103:100];
    67: reg_0593 <= imem04_in[103:100];
    69: reg_0593 <= imem06_in[67:64];
    71: reg_0593 <= imem04_in[103:100];
    72: reg_0593 <= op1_12_out;
    74: reg_0593 <= op1_12_out;
    78: reg_0593 <= imem04_in[103:100];
    79: reg_0593 <= op1_12_out;
    81: reg_0593 <= op1_12_out;
    84: reg_0593 <= op1_12_out;
    86: reg_0593 <= op1_12_out;
    90: reg_0593 <= imem06_in[7:4];
    93: reg_0593 <= imem04_in[103:100];
    96: reg_0593 <= imem06_in[67:64];
    endcase
  end

  // REG#594の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0594 <= imem03_in[75:72];
    32: reg_0594 <= imem06_in[27:24];
    37: reg_0594 <= imem06_in[27:24];
    62: reg_0594 <= imem01_in[55:52];
    64: reg_0594 <= imem00_in[43:40];
    66: reg_0594 <= imem00_in[43:40];
    68: reg_0594 <= imem00_in[43:40];
    70: reg_0594 <= imem06_in[27:24];
    72: reg_0594 <= op1_13_out;
    76: reg_0594 <= imem06_in[27:24];
    78: reg_0594 <= imem01_in[55:52];
    80: reg_0594 <= imem01_in[55:52];
    82: reg_0594 <= imem00_in[43:40];
    84: reg_0594 <= imem01_in[55:52];
    85: reg_0594 <= op1_13_out;
    88: reg_0594 <= op1_13_out;
    93: reg_0594 <= imem03_in[75:72];
    95: reg_0594 <= imem01_in[55:52];
    endcase
  end

  // REG#595の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0595 <= imem03_in[111:108];
    32: reg_0595 <= imem06_in[115:112];
    37: reg_0595 <= imem03_in[111:108];
    39: reg_0595 <= imem06_in[115:112];
    58: reg_0595 <= imem06_in[59:56];
    81: reg_0595 <= imem06_in[115:112];
    84: reg_0595 <= imem06_in[59:56];
    86: reg_0595 <= imem06_in[59:56];
    91: reg_0595 <= imem06_in[115:112];
    93: reg_0595 <= imem06_in[59:56];
    endcase
  end

  // REG#596の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0596 <= imem03_in[27:24];
    32: reg_0596 <= imem06_in[59:56];
    37: reg_0596 <= imem06_in[59:56];
    62: reg_0596 <= imem02_in[55:52];
    64: reg_0596 <= imem02_in[55:52];
    66: reg_0596 <= imem03_in[27:24];
    68: reg_0596 <= imem02_in[111:108];
    70: reg_0596 <= imem03_in[27:24];
    endcase
  end

  // REG#597の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0597 <= imem03_in[103:100];
    32: reg_0597 <= imem06_in[87:84];
    38: reg_0597 <= imem06_in[87:84];
    40: reg_0597 <= imem03_in[103:100];
    42: reg_0597 <= imem06_in[87:84];
    45: reg_0597 <= imem06_in[87:84];
    47: reg_0597 <= imem01_in[7:4];
    50: reg_0597 <= imem03_in[103:100];
    52: reg_0597 <= imem06_in[87:84];
    54: reg_0597 <= imem03_in[103:100];
    56: reg_0597 <= imem06_in[87:84];
    59: reg_0597 <= imem03_in[103:100];
    61: reg_0597 <= imem01_in[7:4];
    63: reg_0597 <= imem03_in[103:100];
    65: reg_0597 <= imem07_in[63:60];
    68: reg_0597 <= imem03_in[103:100];
    70: reg_0597 <= imem03_in[103:100];
    endcase
  end

  // REG#598の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0598 <= imem03_in[3:0];
    32: reg_0598 <= imem03_in[3:0];
    34: reg_0598 <= imem02_in[51:48];
    35: reg_0598 <= op2_01_out;
    64: reg_0598 <= op2_01_out;
    74: reg_0598 <= imem02_in[51:48];
    75: reg_0598 <= op2_01_out;
    endcase
  end

  // REG#599の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0599 <= imem03_in[31:28];
    32: reg_0599 <= imem06_in[7:4];
    38: reg_0599 <= imem03_in[31:28];
    41: reg_0599 <= imem06_in[7:4];
    43: reg_0599 <= imem07_in[87:84];
    endcase
  end

  // REG#600の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0600 <= imem03_in[91:88];
    31: reg_0600 <= op2_00_out;
    50: reg_0600 <= op2_00_out;
    71: reg_0600 <= op2_00_out;
    94: reg_0600 <= op2_00_out;
    endcase
  end

  // REG#601の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0601 <= imem06_in[123:120];
    31: reg_0601 <= op2_01_out;
    51: reg_0601 <= op2_01_out;
    74: reg_0601 <= op2_01_out;
    endcase
  end

  // REG#602の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0602 <= imem03_in[7:4];
    33: reg_0602 <= imem03_in[7:4];
    35: reg_0602 <= imem03_in[3:0];
    37: reg_0602 <= op2_00_out;
    69: reg_0602 <= op2_00_out;
    87: reg_0602 <= op2_00_out;
    endcase
  end

  // REG#603の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0603 <= op1_13_out;
    31: reg_0603 <= op1_13_out;
    35: reg_0603 <= imem03_in[15:12];
    36: reg_0603 <= op1_13_out;
    40: reg_0603 <= op1_13_out;
    42: reg_0603 <= op1_13_out;
    46: reg_0603 <= op1_13_out;
    49: reg_0603 <= imem03_in[15:12];
    51: reg_0603 <= imem03_in[15:12];
    53: reg_0603 <= imem03_in[15:12];
    54: reg_0603 <= op1_13_out;
    56: reg_0603 <= op1_13_out;
    60: reg_0603 <= imem03_in[15:12];
    62: reg_0603 <= imem05_in[47:44];
    64: reg_0603 <= imem00_in[55:52];
    66: reg_0603 <= imem05_in[47:44];
    75: reg_0603 <= op1_13_out;
    77: reg_0603 <= op1_13_out;
    79: reg_0603 <= op1_13_out;
    83: reg_0603 <= imem00_in[55:52];
    85: reg_0603 <= imem00_in[55:52];
    87: reg_0603 <= imem03_in[15:12];
    89: reg_0603 <= imem00_in[55:52];
    91: reg_0603 <= imem05_in[47:44];
    92: reg_0603 <= op1_13_out;
    endcase
  end

  // REG#604の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0604 <= imem06_in[19:16];
    33: reg_0604 <= imem01_in[31:28];
    35: reg_0604 <= imem06_in[19:16];
    38: reg_0604 <= imem06_in[19:16];
    41: reg_0604 <= imem01_in[31:28];
    95: reg_0604 <= imem01_in[31:28];
    endcase
  end

  // REG#605の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0605 <= imem06_in[51:48];
    33: reg_0605 <= imem01_in[83:80];
    35: reg_0605 <= imem01_in[83:80];
    37: reg_0605 <= imem06_in[51:48];
    61: reg_0605 <= imem06_in[51:48];
    72: reg_0605 <= imem06_in[51:48];
    74: reg_0605 <= imem00_in[115:112];
    76: reg_0605 <= imem02_in[39:36];
    78: reg_0605 <= imem06_in[51:48];
    80: reg_0605 <= imem06_in[51:48];
    82: reg_0605 <= imem02_in[39:36];
    84: reg_0605 <= imem02_in[39:36];
    endcase
  end

  // REG#606の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0606 <= imem06_in[67:64];
    33: reg_0606 <= imem02_in[15:12];
    35: reg_0606 <= imem03_in[47:44];
    37: reg_0606 <= imem02_in[15:12];
    39: reg_0606 <= imem02_in[15:12];
    40: reg_0606 <= op2_01_out;
    80: reg_0606 <= op2_01_out;
    84: reg_0606 <= imem06_in[67:64];
    86: reg_0606 <= imem06_in[67:64];
    97: reg_0606 <= op2_01_out;
    endcase
  end

  // REG#607の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0607 <= imem06_in[27:24];
    34: reg_0607 <= imem06_in[27:24];
    36: reg_0607 <= imem06_in[27:24];
    38: reg_0607 <= imem06_in[27:24];
    41: reg_0607 <= imem01_in[3:0];
    92: reg_0607 <= imem01_in[3:0];
    endcase
  end

  // REG#608の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0608 <= imem06_in[91:88];
    34: reg_0608 <= imem02_in[107:104];
    36: reg_0608 <= imem06_in[91:88];
    38: reg_0608 <= imem06_in[91:88];
    40: reg_0608 <= imem06_in[91:88];
    42: reg_0608 <= imem07_in[71:68];
    44: reg_0608 <= imem07_in[71:68];
    46: reg_0608 <= imem07_in[71:68];
    48: reg_0608 <= imem02_in[107:104];
    52: reg_0608 <= imem02_in[107:104];
    endcase
  end

  // REG#609の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0609 <= imem06_in[71:68];
    35: reg_0609 <= imem03_in[67:64];
    37: reg_0609 <= imem06_in[71:68];
    62: reg_0609 <= imem06_in[71:68];
    64: reg_0609 <= imem06_in[71:68];
    68: reg_0609 <= imem03_in[67:64];
    70: reg_0609 <= imem03_in[67:64];
    endcase
  end

  // REG#610の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0610 <= imem06_in[11:8];
    35: reg_0610 <= imem06_in[11:8];
    38: reg_0610 <= imem06_in[11:8];
    41: reg_0610 <= imem01_in[103:100];
    93: reg_0610 <= imem01_in[103:100];
    96: reg_0610 <= imem01_in[103:100];
    endcase
  end

  // REG#611の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0611 <= imem06_in[79:76];
    35: reg_0611 <= imem06_in[79:76];
    39: reg_0611 <= imem06_in[79:76];
    58: reg_0611 <= imem06_in[67:64];
    84: reg_0611 <= imem06_in[79:76];
    86: reg_0611 <= imem05_in[27:24];
    89: reg_0611 <= imem06_in[79:76];
    endcase
  end

  // REG#612の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0612 <= imem06_in[127:124];
    35: reg_0612 <= imem06_in[51:48];
    39: reg_0612 <= imem06_in[127:124];
    56: reg_0612 <= imem06_in[51:48];
    59: reg_0612 <= imem06_in[51:48];
    61: reg_0612 <= imem07_in[127:124];
    63: reg_0612 <= imem07_in[127:124];
    65: reg_0612 <= imem06_in[127:124];
    67: reg_0612 <= imem06_in[51:48];
    69: reg_0612 <= imem06_in[127:124];
    71: reg_0612 <= imem06_in[51:48];
    89: reg_0612 <= imem07_in[127:124];
    92: reg_0612 <= op1_09_out;
    94: reg_0612 <= op1_09_out;
    endcase
  end

  // REG#613の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0613 <= imem06_in[39:36];
    35: reg_0613 <= imem06_in[7:4];
    39: reg_0613 <= imem06_in[7:4];
    58: reg_0613 <= imem06_in[39:36];
    87: reg_0613 <= imem03_in[23:20];
    90: reg_0613 <= imem03_in[23:20];
    endcase
  end

  // REG#614の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0614 <= imem06_in[3:0];
    35: reg_0614 <= imem06_in[3:0];
    39: reg_0614 <= imem06_in[3:0];
    58: reg_0614 <= imem06_in[3:0];
    86: reg_0614 <= imem06_in[3:0];
    endcase
  end

  // REG#615の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0615 <= imem06_in[119:116];
    35: reg_0615 <= imem06_in[119:116];
    38: reg_0615 <= imem06_in[119:116];
    41: reg_0615 <= imem01_in[127:124];
    93: reg_0615 <= imem01_in[127:124];
    endcase
  end

  // REG#616の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0616 <= imem06_in[59:56];
    38: reg_0616 <= imem06_in[59:56];
    41: reg_0616 <= imem01_in[91:88];
    94: reg_0616 <= imem01_in[91:88];
    endcase
  end

  // REG#617の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0617 <= imem06_in[47:44];
    37: reg_0617 <= imem06_in[47:44];
    58: reg_0617 <= imem06_in[47:44];
    87: reg_0617 <= imem05_in[107:104];
    endcase
  end

  // REG#618の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0618 <= imem06_in[99:96];
    36: reg_0618 <= imem06_in[99:96];
    42: reg_0618 <= imem06_in[99:96];
    44: reg_0618 <= op2_00_out;
    51: reg_0618 <= op2_00_out;
    73: reg_0618 <= op2_00_out;
    endcase
  end

  // REG#619の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0619 <= imem06_in[83:80];
    39: reg_0619 <= imem06_in[83:80];
    58: reg_0619 <= imem06_in[127:124];
    85: reg_0619 <= imem06_in[127:124];
    87: reg_0619 <= imem06_in[127:124];
    89: reg_0619 <= imem06_in[83:80];
    91: reg_0619 <= imem06_in[83:80];
    93: reg_0619 <= imem01_in[31:28];
    endcase
  end

  // REG#620の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0620 <= imem06_in[43:40];
    39: reg_0620 <= imem03_in[83:80];
    41: reg_0620 <= imem03_in[83:80];
    43: reg_0620 <= imem06_in[43:40];
    45: reg_0620 <= imem06_in[43:40];
    47: reg_0620 <= imem06_in[43:40];
    49: reg_0620 <= imem06_in[43:40];
    51: reg_0620 <= imem03_in[83:80];
    53: reg_0620 <= imem06_in[43:40];
    55: reg_0620 <= imem03_in[11:8];
    86: reg_0620 <= imem03_in[11:8];
    88: reg_0620 <= imem03_in[83:80];
    endcase
  end

  // REG#621の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0621 <= imem06_in[55:52];
    38: reg_0621 <= imem06_in[55:52];
    42: reg_0621 <= imem07_in[7:4];
    45: reg_0621 <= imem02_in[95:92];
    57: reg_0621 <= imem07_in[7:4];
    59: reg_0621 <= imem06_in[55:52];
    61: reg_0621 <= imem02_in[95:92];
    63: reg_0621 <= imem03_in[3:0];
    65: reg_0621 <= imem00_in[23:20];
    67: reg_0621 <= imem00_in[23:20];
    69: reg_0621 <= imem03_in[3:0];
    71: reg_0621 <= imem02_in[95:92];
    74: reg_0621 <= imem06_in[55:52];
    76: reg_0621 <= imem06_in[55:52];
    78: reg_0621 <= imem02_in[95:92];
    80: reg_0621 <= imem03_in[3:0];
    82: reg_0621 <= imem00_in[23:20];
    84: reg_0621 <= imem02_in[95:92];
    97: reg_0621 <= imem07_in[7:4];
    endcase
  end

  // REG#622の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0622 <= imem06_in[111:108];
    37: reg_0622 <= imem06_in[111:108];
    62: reg_0622 <= imem06_in[123:120];
    64: reg_0622 <= imem00_in[103:100];
    66: reg_0622 <= imem00_in[103:100];
    68: reg_0622 <= imem00_in[103:100];
    71: reg_0622 <= imem00_in[103:100];
    73: reg_0622 <= imem00_in[103:100];
    75: reg_0622 <= imem04_in[43:40];
    78: reg_0622 <= imem04_in[43:40];
    80: reg_0622 <= imem04_in[43:40];
    82: reg_0622 <= imem00_in[103:100];
    84: reg_0622 <= imem04_in[43:40];
    86: reg_0622 <= imem00_in[103:100];
    88: reg_0622 <= imem06_in[123:120];
    91: reg_0622 <= imem06_in[123:120];
    93: reg_0622 <= imem01_in[83:80];
    endcase
  end

  // REG#623の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0623 <= imem06_in[115:112];
    38: reg_0623 <= imem06_in[115:112];
    40: reg_0623 <= imem06_in[115:112];
    42: reg_0623 <= imem07_in[103:100];
    45: reg_0623 <= imem07_in[103:100];
    47: reg_0623 <= imem01_in[19:16];
    50: reg_0623 <= imem01_in[19:16];
    52: reg_0623 <= imem01_in[19:16];
    54: reg_0623 <= imem07_in[103:100];
    56: reg_0623 <= imem01_in[19:16];
    58: reg_0623 <= imem07_in[103:100];
    60: reg_0623 <= imem06_in[115:112];
    62: reg_0623 <= imem01_in[19:16];
    64: reg_0623 <= imem01_in[19:16];
    66: reg_0623 <= imem06_in[115:112];
    68: reg_0623 <= imem03_in[35:32];
    70: reg_0623 <= imem06_in[115:112];
    72: reg_0623 <= imem06_in[107:104];
    74: reg_0623 <= imem07_in[103:100];
    76: reg_0623 <= imem03_in[123:120];
    78: reg_0623 <= imem06_in[107:104];
    80: reg_0623 <= imem03_in[123:120];
    82: reg_0623 <= imem06_in[115:112];
    84: reg_0623 <= imem06_in[115:112];
    86: reg_0623 <= imem01_in[19:16];
    88: reg_0623 <= imem03_in[123:120];
    endcase
  end

  // REG#624の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0624 <= imem06_in[35:32];
    39: reg_0624 <= imem06_in[35:32];
    58: reg_0624 <= imem06_in[35:32];
    82: reg_0624 <= imem02_in[95:92];
    85: reg_0624 <= imem02_in[95:92];
    endcase
  end

  // REG#625の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0625 <= imem06_in[15:12];
    37: reg_0625 <= imem06_in[15:12];
    57: reg_0625 <= imem06_in[15:12];
    endcase
  end

  // REG#626の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0626 <= imem06_in[75:72];
    37: reg_0626 <= imem06_in[75:72];
    57: reg_0626 <= imem06_in[75:72];
    endcase
  end

  // REG#627の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0627 <= imem06_in[107:104];
    39: reg_0627 <= imem06_in[107:104];
    57: reg_0627 <= imem00_in[123:120];
    59: reg_0627 <= imem04_in[63:60];
    endcase
  end

  // REG#628の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0628 <= imem06_in[7:4];
    37: reg_0628 <= imem06_in[7:4];
    62: reg_0628 <= imem07_in[127:124];
    64: reg_0628 <= imem06_in[7:4];
    66: reg_0628 <= imem07_in[127:124];
    68: reg_0628 <= imem06_in[67:64];
    71: reg_0628 <= imem07_in[127:124];
    73: reg_0628 <= imem06_in[7:4];
    75: reg_0628 <= imem07_in[127:124];
    79: reg_0628 <= imem06_in[7:4];
    81: reg_0628 <= imem06_in[7:4];
    85: reg_0628 <= imem06_in[7:4];
    87: reg_0628 <= imem07_in[127:124];
    89: reg_0628 <= imem06_in[67:64];
    endcase
  end

  // REG#629の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0629 <= imem06_in[23:20];
    37: reg_0629 <= imem06_in[23:20];
    61: reg_0629 <= op2_00_out;
    63: reg_0629 <= op2_00_out;
    70: reg_0629 <= imem06_in[23:20];
    72: reg_0629 <= op2_00_out;
    98: reg_0629 <= op2_00_out;
    endcase
  end

  // REG#630の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0630 <= imem06_in[31:28];
    37: reg_0630 <= imem06_in[31:28];
    61: reg_0630 <= imem06_in[31:28];
    72: reg_0630 <= imem01_in[79:76];
    74: reg_0630 <= imem01_in[35:32];
    76: reg_0630 <= imem01_in[35:32];
    78: reg_0630 <= imem01_in[79:76];
    80: reg_0630 <= imem06_in[31:28];
    82: reg_0630 <= imem06_in[31:28];
    84: reg_0630 <= imem06_in[31:28];
    86: reg_0630 <= imem06_in[31:28];
    endcase
  end

  // REG#631の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0631 <= imem06_in[63:60];
    37: reg_0631 <= imem06_in[63:60];
    56: reg_0631 <= imem06_in[63:60];
    60: reg_0631 <= imem06_in[63:60];
    62: reg_0631 <= imem06_in[63:60];
    64: reg_0631 <= imem01_in[59:56];
    66: reg_0631 <= imem01_in[59:56];
    68: reg_0631 <= imem07_in[47:44];
    71: reg_0631 <= imem01_in[59:56];
    73: reg_0631 <= imem07_in[47:44];
    75: reg_0631 <= imem06_in[63:60];
    77: reg_0631 <= imem07_in[47:44];
    79: reg_0631 <= imem06_in[63:60];
    82: reg_0631 <= imem03_in[7:4];
    85: reg_0631 <= imem06_in[63:60];
    88: reg_0631 <= imem03_in[7:4];
    endcase
  end

  // REG#632の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0632 <= imem06_in[103:100];
    39: reg_0632 <= imem06_in[103:100];
    58: reg_0632 <= imem06_in[103:100];
    87: reg_0632 <= imem06_in[103:100];
    89: reg_0632 <= imem06_in[103:100];
    endcase
  end

  // REG#633の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0633 <= imem06_in[87:84];
    37: reg_0633 <= imem06_in[87:84];
    61: reg_0633 <= imem06_in[87:84];
    72: reg_0633 <= imem04_in[47:44];
    74: reg_0633 <= imem06_in[87:84];
    76: reg_0633 <= imem04_in[127:124];
    78: reg_0633 <= imem04_in[47:44];
    80: reg_0633 <= imem06_in[87:84];
    82: reg_0633 <= imem04_in[95:92];
    85: reg_0633 <= imem04_in[95:92];
    87: reg_0633 <= imem04_in[47:44];
    89: reg_0633 <= imem04_in[47:44];
    91: reg_0633 <= imem04_in[47:44];
    92: reg_0633 <= op2_02_out;
    endcase
  end

  // REG#634の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0634 <= op1_14_out;
    36: reg_0634 <= op1_14_out;
    39: reg_0634 <= op1_14_out;
    41: reg_0634 <= op1_14_out;
    44: reg_0634 <= op1_14_out;
    46: reg_0634 <= op1_14_out;
    49: reg_0634 <= imem02_in[43:40];
    50: reg_0634 <= op1_14_out;
    53: reg_0634 <= op1_14_out;
    56: reg_0634 <= op1_14_out;
    59: reg_0634 <= op1_14_out;
    62: reg_0634 <= imem02_in[43:40];
    64: reg_0634 <= op1_14_out;
    67: reg_0634 <= op1_14_out;
    70: reg_0634 <= op1_14_out;
    73: reg_0634 <= op1_14_out;
    76: reg_0634 <= op1_14_out;
    79: reg_0634 <= imem02_in[43:40];
    81: reg_0634 <= imem02_in[43:40];
    83: reg_0634 <= imem02_in[43:40];
    85: reg_0634 <= op1_14_out;
    89: reg_0634 <= imem02_in[43:40];
    90: reg_0634 <= op1_14_out;
    94: reg_0634 <= imem02_in[43:40];
    95: reg_0634 <= op1_14_out;
    endcase
  end

  // REG#635の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0635 <= op1_15_out;
    37: reg_0635 <= op1_15_out;
    40: reg_0635 <= op1_15_out;
    43: reg_0635 <= op1_15_out;
    46: reg_0635 <= op1_15_out;
    49: reg_0635 <= imem03_in[51:48];
    50: reg_0635 <= op1_15_out;
    54: reg_0635 <= imem03_in[51:48];
    55: reg_0635 <= op1_15_out;
    58: reg_0635 <= op1_15_out;
    61: reg_0635 <= op1_15_out;
    64: reg_0635 <= imem01_in[127:124];
    66: reg_0635 <= imem03_in[51:48];
    67: reg_0635 <= op1_15_out;
    70: reg_0635 <= op1_15_out;
    73: reg_0635 <= op1_15_out;
    76: reg_0635 <= op1_15_out;
    79: reg_0635 <= imem01_in[127:124];
    82: reg_0635 <= imem03_in[51:48];
    84: reg_0635 <= imem03_in[51:48];
    85: reg_0635 <= op1_15_out;
    89: reg_0635 <= imem03_in[51:48];
    91: reg_0635 <= op1_15_out;
    94: reg_0635 <= op1_15_out;
    endcase
  end

  // REG#636の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0636 <= imem02_in[115:112];
    42: reg_0636 <= imem07_in[111:108];
    45: reg_0636 <= imem02_in[115:112];
    63: reg_0636 <= imem02_in[115:112];
    73: reg_0636 <= imem05_in[7:4];
    endcase
  end

  // REG#637の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0637 <= imem02_in[35:32];
    42: reg_0637 <= imem07_in[63:60];
    45: reg_0637 <= imem02_in[83:80];
    59: reg_0637 <= imem07_in[63:60];
    61: reg_0637 <= imem07_in[63:60];
    63: reg_0637 <= imem02_in[35:32];
    72: reg_0637 <= imem02_in[35:32];
    84: reg_0637 <= imem02_in[83:80];
    endcase
  end

  // REG#638の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0638 <= imem02_in[83:80];
    41: reg_0638 <= op2_00_out;
    83: reg_0638 <= imem02_in[83:80];
    86: reg_0638 <= op2_00_out;
    endcase
  end

  // REG#639の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0639 <= imem02_in[63:60];
    43: reg_0639 <= imem02_in[63:60];
    45: reg_0639 <= imem02_in[63:60];
    64: reg_0639 <= imem03_in[127:124];
    66: reg_0639 <= imem03_in[127:124];
    68: reg_0639 <= imem00_in[75:72];
    70: reg_0639 <= imem00_in[75:72];
    72: reg_0639 <= imem00_in[75:72];
    74: reg_0639 <= imem00_in[75:72];
    76: reg_0639 <= imem00_in[75:72];
    78: reg_0639 <= imem00_in[75:72];
    80: reg_0639 <= imem00_in[75:72];
    82: reg_0639 <= imem02_in[63:60];
    84: reg_0639 <= imem02_in[63:60];
    endcase
  end

  // REG#640の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0640 <= imem02_in[75:72];
    43: reg_0640 <= imem07_in[119:116];
    endcase
  end

  // REG#641の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0641 <= imem02_in[91:88];
    43: reg_0641 <= imem07_in[75:72];
    endcase
  end

  // REG#642の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0642 <= imem02_in[3:0];
    45: reg_0642 <= imem02_in[3:0];
    62: reg_0642 <= imem02_in[107:104];
    65: reg_0642 <= imem02_in[3:0];
    68: reg_0642 <= imem02_in[3:0];
    71: reg_0642 <= imem02_in[107:104];
    74: reg_0642 <= imem01_in[71:68];
    76: reg_0642 <= imem02_in[3:0];
    78: reg_0642 <= imem02_in[107:104];
    80: reg_0642 <= imem02_in[3:0];
    82: reg_0642 <= imem01_in[71:68];
    84: reg_0642 <= imem02_in[107:104];
    endcase
  end

  // REG#643の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0643 <= imem02_in[103:100];
    45: reg_0643 <= imem02_in[103:100];
    63: reg_0643 <= imem02_in[103:100];
    72: reg_0643 <= imem02_in[103:100];
    85: reg_0643 <= imem02_in[103:100];
    endcase
  end

  // REG#644の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0644 <= imem02_in[99:96];
    44: reg_0644 <= imem02_in[99:96];
    47: reg_0644 <= imem02_in[99:96];
    49: reg_0644 <= imem03_in[71:68];
    52: reg_0644 <= imem02_in[99:96];
    endcase
  end

  // REG#645の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0645 <= imem02_in[11:8];
    44: reg_0645 <= imem02_in[11:8];
    47: reg_0645 <= imem01_in[63:60];
    50: reg_0645 <= imem01_in[63:60];
    52: reg_0645 <= imem02_in[11:8];
    97: reg_0645 <= imem02_in[11:8];
    endcase
  end

  // REG#646の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0646 <= imem02_in[39:36];
    45: reg_0646 <= imem02_in[39:36];
    64: reg_0646 <= imem02_in[39:36];
    68: reg_0646 <= imem01_in[87:84];
    71: reg_0646 <= imem02_in[39:36];
    73: reg_0646 <= imem02_in[39:36];
    75: reg_0646 <= imem07_in[43:40];
    79: reg_0646 <= imem01_in[87:84];
    81: reg_0646 <= imem07_in[43:40];
    83: reg_0646 <= imem01_in[87:84];
    85: reg_0646 <= imem07_in[43:40];
    87: reg_0646 <= imem05_in[23:20];
    endcase
  end

  // REG#647の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0647 <= imem02_in[71:68];
    45: reg_0647 <= imem02_in[71:68];
    63: reg_0647 <= imem02_in[71:68];
    73: reg_0647 <= imem05_in[63:60];
    endcase
  end

  // REG#648の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0648 <= imem02_in[79:76];
    45: reg_0648 <= imem02_in[107:104];
    63: reg_0648 <= imem02_in[107:104];
    71: reg_0648 <= imem02_in[79:76];
    73: reg_0648 <= imem05_in[119:116];
    endcase
  end

  // REG#649の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0649 <= imem02_in[87:84];
    45: reg_0649 <= imem02_in[55:52];
    64: reg_0649 <= imem02_in[87:84];
    66: reg_0649 <= imem02_in[87:84];
    68: reg_0649 <= imem02_in[87:84];
    70: reg_0649 <= imem02_in[55:52];
    72: reg_0649 <= imem02_in[55:52];
    80: reg_0649 <= imem01_in[47:44];
    81: reg_0649 <= op2_01_out;
    86: reg_0649 <= op2_01_out;
    endcase
  end

  // REG#650の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0650 <= imem02_in[7:4];
    45: reg_0650 <= imem02_in[7:4];
    64: reg_0650 <= imem05_in[7:4];
    68: reg_0650 <= imem05_in[7:4];
    72: reg_0650 <= imem02_in[7:4];
    85: reg_0650 <= imem02_in[7:4];
    endcase
  end

  // REG#651の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0651 <= imem02_in[67:64];
    45: reg_0651 <= imem02_in[67:64];
    63: reg_0651 <= imem03_in[7:4];
    65: reg_0651 <= imem01_in[63:60];
    68: reg_0651 <= imem05_in[39:36];
    72: reg_0651 <= imem05_in[39:36];
    74: reg_0651 <= imem05_in[39:36];
    endcase
  end

  // REG#652の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0652 <= imem02_in[119:116];
    45: reg_0652 <= imem02_in[119:116];
    64: reg_0652 <= imem05_in[51:48];
    68: reg_0652 <= imem05_in[51:48];
    73: reg_0652 <= imem05_in[39:36];
    endcase
  end

  // REG#653の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0653 <= imem02_in[27:24];
    45: reg_0653 <= imem02_in[27:24];
    53: reg_0653 <= imem05_in[55:52];
    55: reg_0653 <= imem02_in[27:24];
    57: reg_0653 <= imem03_in[31:28];
    59: reg_0653 <= imem05_in[55:52];
    61: reg_0653 <= imem03_in[31:28];
    63: reg_0653 <= imem02_in[27:24];
    73: reg_0653 <= imem02_in[27:24];
    75: reg_0653 <= imem07_in[123:120];
    79: reg_0653 <= imem07_in[123:120];
    94: reg_0653 <= imem07_in[123:120];
    96: reg_0653 <= imem07_in[123:120];
    endcase
  end

  // REG#654の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0654 <= imem02_in[31:28];
    45: reg_0654 <= imem02_in[31:28];
    59: reg_0654 <= imem02_in[31:28];
    61: reg_0654 <= imem01_in[123:120];
    63: reg_0654 <= imem02_in[31:28];
    74: reg_0654 <= imem02_in[75:72];
    76: reg_0654 <= imem02_in[31:28];
    79: reg_0654 <= imem04_in[87:84];
    82: reg_0654 <= imem04_in[87:84];
    85: reg_0654 <= imem01_in[123:120];
    88: reg_0654 <= imem04_in[23:20];
    91: reg_0654 <= imem04_in[23:20];
    94: reg_0654 <= imem04_in[87:84];
    endcase
  end

  // REG#655の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0655 <= imem02_in[23:20];
    45: reg_0655 <= imem02_in[23:20];
    64: reg_0655 <= imem05_in[59:56];
    68: reg_0655 <= imem05_in[59:56];
    73: reg_0655 <= imem05_in[59:56];
    endcase
  end

  // REG#656の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0656 <= imem02_in[59:56];
    45: reg_0656 <= imem02_in[59:56];
    62: reg_0656 <= imem02_in[59:56];
    65: reg_0656 <= imem04_in[91:88];
    68: reg_0656 <= imem05_in[95:92];
    73: reg_0656 <= imem04_in[91:88];
    75: reg_0656 <= imem04_in[91:88];
    77: reg_0656 <= imem02_in[59:56];
    79: reg_0656 <= imem04_in[91:88];
    82: reg_0656 <= imem04_in[91:88];
    85: reg_0656 <= imem02_in[59:56];
    endcase
  end

  // REG#657の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0657 <= imem02_in[51:48];
    45: reg_0657 <= imem02_in[19:16];
    65: reg_0657 <= imem05_in[111:108];
    68: reg_0657 <= imem02_in[19:16];
    71: reg_0657 <= imem02_in[19:16];
    74: reg_0657 <= imem05_in[111:108];
    endcase
  end

  // REG#658の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0658 <= imem02_in[15:12];
    47: reg_0658 <= imem02_in[15:12];
    49: reg_0658 <= imem06_in[23:20];
    51: reg_0658 <= imem06_in[23:20];
    53: reg_0658 <= imem06_in[23:20];
    55: reg_0658 <= imem02_in[15:12];
    57: reg_0658 <= imem02_in[15:12];
    59: reg_0658 <= imem04_in[23:20];
    endcase
  end

  // REG#659の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0659 <= imem02_in[111:108];
    46: reg_0659 <= op2_01_out;
    58: reg_0659 <= op2_01_out;
    96: reg_0659 <= op2_01_out;
    endcase
  end

  // REG#660の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0660 <= imem02_in[47:44];
    48: reg_0660 <= imem02_in[47:44];
    53: reg_0660 <= imem06_in[3:0];
    55: reg_0660 <= imem06_in[3:0];
    57: reg_0660 <= imem06_in[3:0];
    endcase
  end

  // REG#661の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0661 <= imem02_in[55:52];
    48: reg_0661 <= imem02_in[55:52];
    51: reg_0661 <= imem02_in[55:52];
    55: reg_0661 <= imem03_in[115:112];
    87: reg_0661 <= imem03_in[115:112];
    91: reg_0661 <= imem02_in[55:52];
    endcase
  end

  // REG#662の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0662 <= imem02_in[95:92];
    47: reg_0662 <= imem02_in[95:92];
    49: reg_0662 <= imem02_in[11:8];
    53: reg_0662 <= imem02_in[11:8];
    55: reg_0662 <= imem03_in[119:116];
    88: reg_0662 <= imem03_in[119:116];
    endcase
  end

  // REG#663の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0663 <= imem02_in[127:124];
    48: reg_0663 <= imem04_in[3:0];
    51: reg_0663 <= imem04_in[3:0];
    53: reg_0663 <= imem04_in[3:0];
    55: reg_0663 <= imem00_in[127:124];
    88: reg_0663 <= imem04_in[67:64];
    91: reg_0663 <= imem04_in[67:64];
    93: reg_0663 <= imem04_in[3:0];
    95: reg_0663 <= imem00_in[127:124];
    endcase
  end

  // REG#664の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0664 <= imem02_in[43:40];
    48: reg_0664 <= imem02_in[43:40];
    52: reg_0664 <= imem02_in[43:40];
    endcase
  end

  // REG#665の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0665 <= imem02_in[107:104];
    46: reg_0665 <= imem02_in[107:104];
    49: reg_0665 <= imem02_in[107:104];
    53: reg_0665 <= imem02_in[107:104];
    55: reg_0665 <= imem02_in[107:104];
    56: reg_0665 <= op2_02_out;
    91: reg_0665 <= op2_02_out;
    endcase
  end

  // REG#666の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0666 <= imem02_in[19:16];
    48: reg_0666 <= imem02_in[19:16];
    53: reg_0666 <= imem02_in[19:16];
    55: reg_0666 <= imem02_in[19:16];
    57: reg_0666 <= imem02_in[19:16];
    59: reg_0666 <= imem02_in[19:16];
    61: reg_0666 <= imem02_in[19:16];
    63: reg_0666 <= imem02_in[19:16];
    72: reg_0666 <= imem02_in[19:16];
    84: reg_0666 <= imem02_in[19:16];
    endcase
  end

  // REG#667の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0667 <= imem02_in[123:120];
    49: reg_0667 <= imem02_in[123:120];
    51: reg_0667 <= imem02_in[123:120];
    55: reg_0667 <= imem02_in[123:120];
    57: reg_0667 <= imem02_in[123:120];
    60: reg_0667 <= imem02_in[123:120];
    62: reg_0667 <= imem02_in[123:120];
    65: reg_0667 <= imem05_in[11:8];
    68: reg_0667 <= imem05_in[115:112];
    73: reg_0667 <= imem02_in[123:120];
    75: reg_0667 <= imem07_in[39:36];
    79: reg_0667 <= imem05_in[11:8];
    87: reg_0667 <= imem07_in[39:36];
    89: reg_0667 <= imem05_in[115:112];
    91: reg_0667 <= imem07_in[39:36];
    93: reg_0667 <= imem05_in[11:8];
    endcase
  end

  // REG#668の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0668 <= imem00_in[95:92];
    51: reg_0668 <= imem00_in[95:92];
    53: reg_0668 <= imem06_in[59:56];
    55: reg_0668 <= imem00_in[95:92];
    88: reg_0668 <= imem06_in[59:56];
    90: reg_0668 <= imem00_in[95:92];
    92: reg_0668 <= imem06_in[59:56];
    endcase
  end

  // REG#669の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0669 <= imem00_in[123:120];
    53: reg_0669 <= imem07_in[91:88];
    55: reg_0669 <= imem00_in[123:120];
    92: reg_0669 <= imem00_in[123:120];
    endcase
  end

  // REG#670の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0670 <= imem00_in[63:60];
    53: reg_0670 <= imem00_in[63:60];
    55: reg_0670 <= imem00_in[63:60];
    endcase
  end

  // REG#671の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0671 <= imem00_in[87:84];
    53: reg_0671 <= imem00_in[23:20];
    55: reg_0671 <= imem00_in[23:20];
    90: reg_0671 <= imem00_in[23:20];
    94: reg_0671 <= imem00_in[87:84];
    endcase
  end

  // REG#672の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0672 <= imem00_in[35:32];
    53: reg_0672 <= imem02_in[119:116];
    55: reg_0672 <= imem02_in[119:116];
    57: reg_0672 <= imem02_in[119:116];
    59: reg_0672 <= imem00_in[35:32];
    61: reg_0672 <= imem03_in[83:80];
    63: reg_0672 <= imem03_in[83:80];
    65: reg_0672 <= imem03_in[83:80];
    68: reg_0672 <= imem00_in[35:32];
    70: reg_0672 <= imem03_in[83:80];
    endcase
  end

  // REG#673の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0673 <= imem00_in[111:108];
    53: reg_0673 <= imem03_in[103:100];
    56: reg_0673 <= imem06_in[79:76];
    60: reg_0673 <= imem00_in[111:108];
    62: reg_0673 <= imem02_in[99:96];
    66: reg_0673 <= imem00_in[111:108];
    68: reg_0673 <= imem05_in[79:76];
    74: reg_0673 <= imem03_in[103:100];
    76: reg_0673 <= imem00_in[111:108];
    78: reg_0673 <= imem06_in[79:76];
    80: reg_0673 <= imem05_in[3:0];
    82: reg_0673 <= imem00_in[111:108];
    84: reg_0673 <= imem03_in[103:100];
    86: reg_0673 <= imem05_in[79:76];
    89: reg_0673 <= imem05_in[79:76];
    91: reg_0673 <= imem03_in[103:100];
    93: reg_0673 <= imem02_in[99:96];
    96: reg_0673 <= imem05_in[3:0];
    endcase
  end

  // REG#674の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0674 <= imem00_in[83:80];
    53: reg_0674 <= imem00_in[83:80];
    55: reg_0674 <= imem00_in[83:80];
    92: reg_0674 <= imem00_in[83:80];
    endcase
  end

  // REG#675の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0675 <= imem00_in[99:96];
    53: reg_0675 <= imem03_in[55:52];
    56: reg_0675 <= imem05_in[35:32];
    63: reg_0675 <= imem06_in[123:120];
    66: reg_0675 <= imem05_in[35:32];
    79: reg_0675 <= imem06_in[123:120];
    82: reg_0675 <= imem03_in[55:52];
    85: reg_0675 <= imem00_in[99:96];
    87: reg_0675 <= imem05_in[35:32];
    endcase
  end

  // REG#676の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0676 <= imem00_in[43:40];
    53: reg_0676 <= imem03_in[71:68];
    57: reg_0676 <= imem03_in[71:68];
    60: reg_0676 <= imem00_in[43:40];
    63: reg_0676 <= imem01_in[111:108];
    65: reg_0676 <= imem01_in[111:108];
    67: reg_0676 <= imem03_in[71:68];
    69: reg_0676 <= imem03_in[71:68];
    72: reg_0676 <= imem06_in[71:68];
    74: reg_0676 <= imem04_in[19:16];
    76: reg_0676 <= imem05_in[27:24];
    78: reg_0676 <= imem05_in[27:24];
    81: reg_0676 <= imem05_in[27:24];
    83: reg_0676 <= imem00_in[43:40];
    85: reg_0676 <= imem01_in[111:108];
    87: reg_0676 <= imem00_in[43:40];
    90: reg_0676 <= imem05_in[27:24];
    93: reg_0676 <= imem00_in[43:40];
    endcase
  end

  // REG#677の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0677 <= imem00_in[75:72];
    53: reg_0677 <= imem03_in[111:108];
    57: reg_0677 <= imem03_in[111:108];
    60: reg_0677 <= imem00_in[75:72];
    63: reg_0677 <= imem04_in[119:116];
    67: reg_0677 <= imem00_in[75:72];
    69: reg_0677 <= imem03_in[111:108];
    71: reg_0677 <= imem00_in[75:72];
    73: reg_0677 <= imem04_in[119:116];
    75: reg_0677 <= imem07_in[67:64];
    78: reg_0677 <= imem04_in[119:116];
    80: reg_0677 <= imem07_in[15:12];
    83: reg_0677 <= imem07_in[15:12];
    85: reg_0677 <= imem03_in[99:96];
    87: reg_0677 <= imem03_in[99:96];
    89: reg_0677 <= imem03_in[111:108];
    92: reg_0677 <= imem07_in[67:64];
    95: reg_0677 <= imem07_in[15:12];
    endcase
  end

  // REG#678の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0678 <= imem00_in[91:88];
    53: reg_0678 <= imem03_in[75:72];
    57: reg_0678 <= imem00_in[91:88];
    60: reg_0678 <= imem03_in[75:72];
    62: reg_0678 <= imem00_in[91:88];
    65: reg_0678 <= imem00_in[91:88];
    67: reg_0678 <= imem03_in[75:72];
    69: reg_0678 <= imem07_in[23:20];
    72: reg_0678 <= imem03_in[75:72];
    74: reg_0678 <= imem07_in[23:20];
    78: reg_0678 <= imem07_in[23:20];
    80: reg_0678 <= imem07_in[23:20];
    83: reg_0678 <= imem07_in[23:20];
    85: reg_0678 <= imem04_in[51:48];
    87: reg_0678 <= imem03_in[75:72];
    90: reg_0678 <= imem07_in[23:20];
    94: reg_0678 <= imem03_in[75:72];
    endcase
  end

  // REG#679の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0679 <= imem00_in[67:64];
    54: reg_0679 <= imem00_in[67:64];
    57: reg_0679 <= imem06_in[79:76];
    94: reg_0679 <= imem06_in[79:76];
    endcase
  end

  // REG#680の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0680 <= imem00_in[103:100];
    55: reg_0680 <= imem00_in[103:100];
    91: reg_0680 <= imem00_in[103:100];
    endcase
  end

  // REG#681の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0681 <= imem00_in[23:20];
    55: reg_0681 <= imem03_in[27:24];
    89: reg_0681 <= imem03_in[27:24];
    93: reg_0681 <= imem03_in[27:24];
    95: reg_0681 <= imem03_in[27:24];
    endcase
  end

  // REG#682の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0682 <= imem00_in[7:4];
    55: reg_0682 <= imem00_in[7:4];
    91: reg_0682 <= imem00_in[7:4];
    endcase
  end

  // REG#683の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0683 <= imem00_in[19:16];
    55: reg_0683 <= imem00_in[19:16];
    91: reg_0683 <= imem00_in[19:16];
    endcase
  end

  // REG#684の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0684 <= imem00_in[55:52];
    55: reg_0684 <= imem00_in[55:52];
    91: reg_0684 <= imem00_in[55:52];
    endcase
  end

  // REG#685の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0685 <= imem00_in[31:28];
    55: reg_0685 <= imem00_in[31:28];
    93: reg_0685 <= imem00_in[31:28];
    95: reg_0685 <= imem00_in[31:28];
    endcase
  end

  // REG#686の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0686 <= imem00_in[59:56];
    55: reg_0686 <= imem00_in[59:56];
    endcase
  end

  // REG#687の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0687 <= imem00_in[115:112];
    55: reg_0687 <= imem00_in[115:112];
    85: reg_0687 <= imem00_in[115:112];
    87: reg_0687 <= op1_11_out;
    90: reg_0687 <= imem00_in[115:112];
    94: reg_0687 <= op1_11_out;
    endcase
  end

  // REG#688の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0688 <= imem00_in[107:104];
    56: reg_0688 <= imem05_in[63:60];
    62: reg_0688 <= imem00_in[107:104];
    64: reg_0688 <= imem05_in[63:60];
    66: reg_0688 <= imem05_in[63:60];
    78: reg_0688 <= imem05_in[63:60];
    80: reg_0688 <= imem07_in[123:120];
    84: reg_0688 <= imem05_in[63:60];
    86: reg_0688 <= imem00_in[107:104];
    88: reg_0688 <= imem06_in[27:24];
    91: reg_0688 <= imem06_in[27:24];
    93: reg_0688 <= imem05_in[63:60];
    endcase
  end

  // REG#689の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0689 <= imem00_in[51:48];
    56: reg_0689 <= imem05_in[107:104];
    62: reg_0689 <= imem00_in[51:48];
    64: reg_0689 <= imem05_in[107:104];
    68: reg_0689 <= imem05_in[107:104];
    73: reg_0689 <= imem05_in[107:104];
    endcase
  end

  // REG#690の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0690 <= imem00_in[71:68];
    56: reg_0690 <= imem00_in[71:68];
    58: reg_0690 <= imem00_in[71:68];
    60: reg_0690 <= imem06_in[71:68];
    63: reg_0690 <= imem00_in[71:68];
    65: reg_0690 <= imem00_in[71:68];
    68: reg_0690 <= imem05_in[19:16];
    74: reg_0690 <= imem04_in[67:64];
    76: reg_0690 <= imem05_in[19:16];
    78: reg_0690 <= imem06_in[71:68];
    80: reg_0690 <= imem05_in[19:16];
    82: reg_0690 <= imem07_in[91:88];
    95: reg_0690 <= imem00_in[71:68];
    97: reg_0690 <= imem05_in[19:16];
    endcase
  end

  // REG#691の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0691 <= imem00_in[79:76];
    57: reg_0691 <= imem06_in[35:32];
    95: reg_0691 <= imem00_in[79:76];
    endcase
  end

  // REG#692の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0692 <= imem00_in[119:116];
    57: reg_0692 <= imem06_in[127:124];
    endcase
  end

  // REG#693の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0693 <= imem00_in[11:8];
    57: reg_0693 <= imem00_in[11:8];
    60: reg_0693 <= imem06_in[79:76];
    63: reg_0693 <= imem00_in[11:8];
    68: reg_0693 <= imem05_in[23:20];
    74: reg_0693 <= imem00_in[11:8];
    76: reg_0693 <= imem05_in[31:28];
    78: reg_0693 <= imem05_in[31:28];
    80: reg_0693 <= imem07_in[51:48];
    84: reg_0693 <= imem00_in[11:8];
    86: reg_0693 <= imem00_in[11:8];
    88: reg_0693 <= imem00_in[11:8];
    90: reg_0693 <= imem07_in[51:48];
    92: reg_0693 <= imem05_in[23:20];
    94: reg_0693 <= imem05_in[23:20];
    endcase
  end

  // REG#694の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0694 <= imem00_in[39:36];
    57: reg_0694 <= imem06_in[19:16];
    endcase
  end

  // REG#695の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0695 <= imem00_in[3:0];
    56: reg_0695 <= imem00_in[3:0];
    58: reg_0695 <= imem06_in[123:120];
    85: reg_0695 <= imem05_in[43:40];
    87: reg_0695 <= imem05_in[43:40];
    endcase
  end

  // REG#696の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0696 <= imem00_in[27:24];
    57: reg_0696 <= imem06_in[31:28];
    endcase
  end

  // REG#697の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0697 <= imem00_in[15:12];
    57: reg_0697 <= imem00_in[15:12];
    60: reg_0697 <= imem06_in[19:16];
    63: reg_0697 <= imem06_in[43:40];
    68: reg_0697 <= imem06_in[43:40];
    70: reg_0697 <= imem00_in[15:12];
    72: reg_0697 <= imem06_in[79:76];
    74: reg_0697 <= imem06_in[43:40];
    76: reg_0697 <= imem00_in[15:12];
    78: reg_0697 <= imem06_in[43:40];
    80: reg_0697 <= imem06_in[19:16];
    82: reg_0697 <= imem07_in[99:96];
    97: reg_0697 <= imem07_in[99:96];
    endcase
  end

  // REG#698の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0698 <= imem00_in[47:44];
    58: reg_0698 <= imem06_in[63:60];
    86: reg_0698 <= imem06_in[63:60];
    endcase
  end

  // REG#699の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0699 <= imem00_in[127:124];
    56: reg_0699 <= imem00_in[127:124];
    58: reg_0699 <= imem06_in[99:96];
    87: reg_0699 <= imem06_in[99:96];
    91: reg_0699 <= imem00_in[127:124];
    endcase
  end

  // REG#700の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0700 <= imem07_in[123:120];
    63: reg_0700 <= imem07_in[123:120];
    65: reg_0700 <= imem07_in[123:120];
    67: reg_0700 <= imem07_in[123:120];
    69: reg_0700 <= imem02_in[47:44];
    72: reg_0700 <= imem02_in[47:44];
    85: reg_0700 <= imem02_in[47:44];
    endcase
  end

  // REG#701の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0701 <= imem07_in[115:112];
    72: reg_0701 <= imem00_in[35:32];
    74: reg_0701 <= imem07_in[31:28];
    76: reg_0701 <= imem05_in[75:72];
    78: reg_0701 <= imem00_in[35:32];
    80: reg_0701 <= imem00_in[35:32];
    82: reg_0701 <= imem07_in[71:68];
    endcase
  end

  // REG#702の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0702 <= imem07_in[63:60];
    72: reg_0702 <= imem07_in[63:60];
    73: reg_0702 <= op1_05_out;
    75: reg_0702 <= op1_05_out;
    77: reg_0702 <= op1_05_out;
    79: reg_0702 <= op1_05_out;
    81: reg_0702 <= op1_05_out;
    83: reg_0702 <= op1_05_out;
    85: reg_0702 <= op1_05_out;
    87: reg_0702 <= op1_05_out;
    89: reg_0702 <= op1_05_out;
    91: reg_0702 <= op1_05_out;
    93: reg_0702 <= op1_05_out;
    95: reg_0702 <= op1_05_out;
    97: reg_0702 <= op1_05_out;
    endcase
  end

  // REG#703の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0703 <= imem07_in[67:64];
    72: reg_0703 <= imem00_in[99:96];
    74: reg_0703 <= imem00_in[99:96];
    76: reg_0703 <= imem05_in[83:80];
    78: reg_0703 <= imem00_in[99:96];
    80: reg_0703 <= imem05_in[83:80];
    82: reg_0703 <= imem07_in[39:36];
    endcase
  end

  // REG#704の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0704 <= imem07_in[15:12];
    74: reg_0704 <= imem07_in[15:12];
    78: reg_0704 <= imem07_in[15:12];
    85: reg_0704 <= imem06_in[59:56];
    88: reg_0704 <= imem07_in[15:12];
    91: reg_0704 <= imem07_in[15:12];
    endcase
  end

  // REG#705の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0705 <= imem07_in[91:88];
    74: reg_0705 <= imem07_in[91:88];
    78: reg_0705 <= imem07_in[91:88];
    80: reg_0705 <= imem07_in[111:108];
    85: reg_0705 <= imem07_in[111:108];
    88: reg_0705 <= imem06_in[79:76];
    93: reg_0705 <= imem07_in[111:108];
    endcase
  end

  // REG#706の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0706 <= imem07_in[119:116];
    74: reg_0706 <= imem05_in[47:44];
    endcase
  end

  // REG#707の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0707 <= imem07_in[111:108];
    74: reg_0707 <= imem05_in[3:0];
    endcase
  end

  // REG#708の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0708 <= imem07_in[83:80];
    74: reg_0708 <= imem07_in[83:80];
    79: reg_0708 <= imem07_in[83:80];
    endcase
  end

  // REG#709の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0709 <= imem07_in[87:84];
    74: reg_0709 <= imem05_in[27:24];
    endcase
  end

  // REG#710の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0710 <= imem07_in[31:28];
    75: reg_0710 <= imem07_in[31:28];
    79: reg_0710 <= imem07_in[31:28];
    endcase
  end

  // REG#711の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0711 <= imem07_in[107:104];
    74: reg_0711 <= op1_13_out;
    78: reg_0711 <= imem07_in[107:104];
    80: reg_0711 <= imem07_in[107:104];
    83: reg_0711 <= op1_13_out;
    86: reg_0711 <= imem05_in[63:60];
    89: reg_0711 <= imem07_in[107:104];
    91: reg_0711 <= imem05_in[63:60];
    endcase
  end

  // REG#712の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0712 <= imem07_in[71:68];
    75: reg_0712 <= imem07_in[15:12];
    79: reg_0712 <= imem07_in[15:12];
    93: reg_0712 <= imem07_in[71:68];
    endcase
  end

  // REG#713の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0713 <= imem07_in[95:92];
    75: reg_0713 <= imem07_in[35:32];
    80: reg_0713 <= imem07_in[35:32];
    85: reg_0713 <= imem02_in[83:80];
    93: reg_0713 <= imem07_in[95:92];
    95: reg_0713 <= imem07_in[95:92];
    endcase
  end

  // REG#714の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0714 <= imem07_in[59:56];
    75: reg_0714 <= imem07_in[59:56];
    79: reg_0714 <= imem04_in[127:124];
    82: reg_0714 <= imem07_in[59:56];
    endcase
  end

  // REG#715の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0715 <= imem07_in[99:96];
    75: reg_0715 <= imem07_in[99:96];
    79: reg_0715 <= imem07_in[99:96];
    endcase
  end

  // REG#716の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0716 <= imem07_in[11:8];
    75: reg_0716 <= imem07_in[7:4];
    80: reg_0716 <= imem07_in[7:4];
    83: reg_0716 <= imem07_in[7:4];
    85: reg_0716 <= imem07_in[11:8];
    88: reg_0716 <= imem07_in[7:4];
    90: reg_0716 <= imem07_in[7:4];
    92: reg_0716 <= imem07_in[7:4];
    94: reg_0716 <= imem07_in[11:8];
    endcase
  end

  // REG#717の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0717 <= imem07_in[51:48];
    76: reg_0717 <= imem07_in[51:48];
    79: reg_0717 <= imem07_in[51:48];
    endcase
  end

  // REG#718の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0718 <= imem07_in[103:100];
    76: reg_0718 <= imem06_in[23:20];
    79: reg_0718 <= imem07_in[103:100];
    endcase
  end

  // REG#719の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0719 <= imem07_in[19:16];
    76: reg_0719 <= imem07_in[19:16];
    78: reg_0719 <= imem07_in[19:16];
    84: reg_0719 <= imem07_in[19:16];
    86: reg_0719 <= imem06_in[111:108];
    94: reg_0719 <= imem06_in[111:108];
    endcase
  end

  // REG#720の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0720 <= imem07_in[23:20];
    76: reg_0720 <= imem07_in[23:20];
    79: reg_0720 <= imem07_in[23:20];
    endcase
  end

  // REG#721の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0721 <= imem07_in[39:36];
    76: reg_0721 <= imem07_in[39:36];
    79: reg_0721 <= imem07_in[39:36];
    endcase
  end

  // REG#722の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0722 <= imem07_in[3:0];
    76: reg_0722 <= imem07_in[3:0];
    79: reg_0722 <= imem07_in[3:0];
    endcase
  end

  // REG#723の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0723 <= imem07_in[43:40];
    76: reg_0723 <= imem06_in[63:60];
    79: reg_0723 <= imem01_in[15:12];
    82: reg_0723 <= imem07_in[43:40];
    endcase
  end

  // REG#724の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0724 <= imem07_in[75:72];
    76: reg_0724 <= imem07_in[107:104];
    78: reg_0724 <= imem07_in[75:72];
    82: reg_0724 <= imem07_in[107:104];
    endcase
  end

  // REG#725の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0725 <= imem07_in[55:52];
    75: reg_0725 <= op1_03_out;
    77: reg_0725 <= op1_03_out;
    80: reg_0725 <= imem07_in[127:124];
    83: reg_0725 <= op1_03_out;
    86: reg_0725 <= imem07_in[55:52];
    88: reg_0725 <= imem06_in[127:124];
    92: reg_0725 <= imem07_in[55:52];
    endcase
  end

  // REG#726の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0726 <= imem07_in[47:44];
    79: reg_0726 <= imem07_in[47:44];
    endcase
  end

  // REG#727の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0727 <= imem07_in[127:124];
    77: reg_0727 <= imem07_in[127:124];
    79: reg_0727 <= imem07_in[127:124];
    endcase
  end

  // REG#728の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0728 <= imem07_in[7:4];
    79: reg_0728 <= imem07_in[7:4];
    endcase
  end

  // REG#729の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0729 <= imem07_in[79:76];
    76: reg_0729 <= imem07_in[79:76];
    78: reg_0729 <= imem07_in[79:76];
    84: reg_0729 <= imem07_in[79:76];
    86: reg_0729 <= imem06_in[39:36];
    endcase
  end

  // REG#730の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0730 <= imem07_in[27:24];
    78: reg_0730 <= imem07_in[27:24];
    85: reg_0730 <= imem02_in[87:84];
    endcase
  end

  // REG#731の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0731 <= imem07_in[35:32];
    79: reg_0731 <= imem04_in[103:100];
    82: reg_0731 <= imem07_in[35:32];
    endcase
  end

  // REG#732の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0732 <= imem00_in[59:56];
    7: reg_0732 <= imem07_in[51:48];
    9: reg_0732 <= imem00_in[59:56];
    11: reg_0732 <= imem00_in[59:56];
    13: reg_0732 <= imem00_in[59:56];
    15: reg_0732 <= imem00_in[59:56];
    17: reg_0732 <= imem00_in[59:56];
    19: reg_0732 <= imem04_in[119:116];
    39: reg_0732 <= imem04_in[119:116];
    42: reg_0732 <= imem04_in[119:116];
    endcase
  end

  // REG#733の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0733 <= imem00_in[111:108];
    7: reg_0733 <= imem07_in[67:64];
    9: reg_0733 <= imem00_in[111:108];
    11: reg_0733 <= imem00_in[111:108];
    13: reg_0733 <= imem07_in[23:20];
    15: reg_0733 <= imem07_in[23:20];
    17: reg_0733 <= imem00_in[111:108];
    19: reg_0733 <= imem04_in[15:12];
    42: reg_0733 <= imem00_in[111:108];
    44: reg_0733 <= imem04_in[15:12];
    46: reg_0733 <= imem07_in[23:20];
    48: reg_0733 <= imem04_in[15:12];
    51: reg_0733 <= imem07_in[67:64];
    53: reg_0733 <= imem01_in[59:56];
    endcase
  end

  // REG#734の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0734 <= imem00_in[115:112];
    7: reg_0734 <= imem07_in[71:68];
    9: reg_0734 <= imem00_in[115:112];
    11: reg_0734 <= imem00_in[115:112];
    13: reg_0734 <= imem07_in[35:32];
    15: reg_0734 <= imem00_in[115:112];
    17: reg_0734 <= imem00_in[115:112];
    19: reg_0734 <= imem07_in[35:32];
    21: reg_0734 <= imem07_in[35:32];
    23: reg_0734 <= imem07_in[35:32];
    25: reg_0734 <= imem07_in[71:68];
    27: reg_0734 <= imem07_in[35:32];
    29: reg_0734 <= imem07_in[35:32];
    31: reg_0734 <= imem07_in[71:68];
    33: reg_0734 <= imem03_in[123:120];
    35: reg_0734 <= imem03_in[123:120];
    38: reg_0734 <= imem00_in[115:112];
    41: reg_0734 <= imem00_in[115:112];
    44: reg_0734 <= imem07_in[35:32];
    47: reg_0734 <= imem07_in[35:32];
    49: reg_0734 <= imem02_in[19:16];
    53: reg_0734 <= imem03_in[123:120];
    57: reg_0734 <= imem00_in[115:112];
    60: reg_0734 <= imem06_in[95:92];
    63: reg_0734 <= imem03_in[123:120];
    66: reg_0734 <= imem07_in[71:68];
    68: reg_0734 <= imem06_in[95:92];
    70: reg_0734 <= imem06_in[95:92];
    72: reg_0734 <= imem05_in[127:124];
    75: reg_0734 <= imem03_in[123:120];
    77: reg_0734 <= imem03_in[123:120];
    79: reg_0734 <= imem06_in[95:92];
    81: reg_0734 <= imem05_in[127:124];
    83: reg_0734 <= imem05_in[127:124];
    85: reg_0734 <= imem02_in[19:16];
    endcase
  end

  // REG#735の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0735 <= imem01_in[47:44];
    7: reg_0735 <= imem07_in[79:76];
    9: reg_0735 <= imem07_in[79:76];
    11: reg_0735 <= imem01_in[47:44];
    26: reg_0735 <= imem07_in[79:76];
    28: reg_0735 <= imem06_in[115:112];
    31: reg_0735 <= imem06_in[115:112];
    33: reg_0735 <= imem06_in[115:112];
    35: reg_0735 <= imem06_in[115:112];
    39: reg_0735 <= imem01_in[47:44];
    42: reg_0735 <= imem07_in[79:76];
    45: reg_0735 <= imem01_in[47:44];
    47: reg_0735 <= imem01_in[47:44];
    51: reg_0735 <= imem07_in[79:76];
    53: reg_0735 <= imem06_in[115:112];
    55: reg_0735 <= imem07_in[79:76];
    57: reg_0735 <= imem06_in[115:112];
    endcase
  end

  // REG#736の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0736 <= imem01_in[59:56];
    7: reg_0736 <= imem00_in[11:8];
    9: reg_0736 <= imem04_in[27:24];
    11: reg_0736 <= imem05_in[111:108];
    13: reg_0736 <= imem00_in[11:8];
    16: reg_0736 <= imem04_in[27:24];
    18: reg_0736 <= imem04_in[27:24];
    46: reg_0736 <= imem00_in[11:8];
    48: reg_0736 <= imem05_in[111:108];
    50: reg_0736 <= imem04_in[27:24];
    52: reg_0736 <= imem05_in[111:108];
    54: reg_0736 <= imem00_in[11:8];
    56: reg_0736 <= imem01_in[59:56];
    58: reg_0736 <= imem01_in[59:56];
    60: reg_0736 <= imem01_in[59:56];
    63: reg_0736 <= imem05_in[111:108];
    65: reg_0736 <= imem01_in[59:56];
    67: reg_0736 <= imem01_in[59:56];
    69: reg_0736 <= imem05_in[111:108];
    72: reg_0736 <= imem05_in[11:8];
    77: reg_0736 <= imem05_in[111:108];
    79: reg_0736 <= imem05_in[111:108];
    87: reg_0736 <= imem05_in[111:108];
    93: reg_0736 <= imem00_in[11:8];
    endcase
  end

  // REG#737の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0737 <= imem01_in[83:80];
    7: reg_0737 <= imem00_in[39:36];
    9: reg_0737 <= imem01_in[83:80];
    13: reg_0737 <= imem00_in[39:36];
    15: reg_0737 <= imem00_in[39:36];
    17: reg_0737 <= imem02_in[59:56];
    19: reg_0737 <= imem00_in[39:36];
    21: reg_0737 <= imem00_in[39:36];
    23: reg_0737 <= imem00_in[39:36];
    25: reg_0737 <= imem02_in[59:56];
    28: reg_0737 <= imem02_in[59:56];
    30: reg_0737 <= imem02_in[59:56];
    32: reg_0737 <= imem02_in[59:56];
    34: reg_0737 <= imem02_in[59:56];
    39: reg_0737 <= imem04_in[95:92];
    41: reg_0737 <= imem01_in[83:80];
    95: reg_0737 <= imem01_in[83:80];
    endcase
  end

  // REG#738の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0738 <= imem01_in[91:88];
    7: reg_0738 <= imem00_in[71:68];
    9: reg_0738 <= imem01_in[91:88];
    11: reg_0738 <= imem06_in[51:48];
    13: reg_0738 <= imem00_in[71:68];
    16: reg_0738 <= imem00_in[71:68];
    18: reg_0738 <= imem04_in[35:32];
    45: reg_0738 <= imem00_in[71:68];
    47: reg_0738 <= imem01_in[91:88];
    50: reg_0738 <= imem01_in[91:88];
    52: reg_0738 <= imem06_in[51:48];
    55: reg_0738 <= imem00_in[71:68];
    91: reg_0738 <= imem00_in[71:68];
    endcase
  end

  // REG#739の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0739 <= imem02_in[23:20];
    7: reg_0739 <= imem00_in[83:80];
    9: reg_0739 <= imem02_in[23:20];
    11: reg_0739 <= imem00_in[83:80];
    13: reg_0739 <= imem02_in[23:20];
    15: reg_0739 <= imem00_in[83:80];
    17: reg_0739 <= imem00_in[83:80];
    19: reg_0739 <= imem00_in[83:80];
    21: reg_0739 <= imem00_in[83:80];
    23: reg_0739 <= imem07_in[103:100];
    25: reg_0739 <= imem00_in[83:80];
    27: reg_0739 <= imem00_in[83:80];
    29: reg_0739 <= imem00_in[83:80];
    31: reg_0739 <= imem00_in[123:120];
    33: reg_0739 <= imem00_in[83:80];
    35: reg_0739 <= imem00_in[83:80];
    37: reg_0739 <= imem00_in[123:120];
    39: reg_0739 <= imem07_in[103:100];
    41: reg_0739 <= imem00_in[83:80];
    43: reg_0739 <= imem00_in[83:80];
    46: reg_0739 <= imem07_in[103:100];
    49: reg_0739 <= imem05_in[23:20];
    52: reg_0739 <= imem02_in[23:20];
    endcase
  end

  // REG#740の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0740 <= imem02_in[43:40];
    7: reg_0740 <= imem01_in[107:104];
    9: reg_0740 <= imem01_in[107:104];
    13: reg_0740 <= imem02_in[43:40];
    15: reg_0740 <= imem01_in[107:104];
    17: reg_0740 <= imem02_in[43:40];
    19: reg_0740 <= imem04_in[11:8];
    41: reg_0740 <= imem01_in[107:104];
    93: reg_0740 <= imem01_in[107:104];
    95: reg_0740 <= imem01_in[107:104];
    endcase
  end

  // REG#741の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0741 <= imem02_in[71:68];
    7: reg_0741 <= imem02_in[11:8];
    9: reg_0741 <= imem02_in[71:68];
    11: reg_0741 <= imem06_in[67:64];
    13: reg_0741 <= imem07_in[91:88];
    15: reg_0741 <= imem02_in[71:68];
    17: reg_0741 <= imem06_in[67:64];
    19: reg_0741 <= imem06_in[67:64];
    21: reg_0741 <= imem07_in[91:88];
    23: reg_0741 <= imem02_in[11:8];
    25: reg_0741 <= imem06_in[67:64];
    27: reg_0741 <= imem02_in[11:8];
    29: reg_0741 <= imem06_in[67:64];
    60: reg_0741 <= imem07_in[91:88];
    63: reg_0741 <= imem02_in[11:8];
    74: reg_0741 <= imem05_in[107:104];
    endcase
  end

  // REG#742の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0742 <= imem02_in[75:72];
    7: reg_0742 <= imem02_in[75:72];
    9: reg_0742 <= imem04_in[95:92];
    11: reg_0742 <= imem06_in[107:104];
    13: reg_0742 <= imem00_in[47:44];
    15: reg_0742 <= imem00_in[47:44];
    17: reg_0742 <= imem04_in[95:92];
    20: reg_0742 <= op2_00_out;
    55: reg_0742 <= op2_00_out;
    85: reg_0742 <= op2_00_out;
    endcase
  end

  // REG#743の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0743 <= imem03_in[39:36];
    7: reg_0743 <= imem02_in[19:16];
    9: reg_0743 <= imem03_in[39:36];
    11: reg_0743 <= imem02_in[19:16];
    13: reg_0743 <= imem00_in[83:80];
    16: reg_0743 <= imem05_in[115:112];
    18: reg_0743 <= imem05_in[115:112];
    20: reg_0743 <= imem02_in[19:16];
    23: reg_0743 <= imem02_in[19:16];
    25: reg_0743 <= imem02_in[19:16];
    28: reg_0743 <= imem05_in[115:112];
    30: reg_0743 <= imem05_in[115:112];
    33: reg_0743 <= imem05_in[115:112];
    35: reg_0743 <= imem02_in[19:16];
    39: reg_0743 <= imem00_in[83:80];
    41: reg_0743 <= imem02_in[19:16];
    44: reg_0743 <= imem00_in[83:80];
    46: reg_0743 <= imem00_in[83:80];
    48: reg_0743 <= imem03_in[39:36];
    50: reg_0743 <= imem03_in[39:36];
    53: reg_0743 <= imem03_in[39:36];
    57: reg_0743 <= imem03_in[39:36];
    59: reg_0743 <= imem03_in[39:36];
    61: reg_0743 <= imem00_in[83:80];
    63: reg_0743 <= imem03_in[47:44];
    65: reg_0743 <= imem00_in[83:80];
    67: reg_0743 <= imem00_in[83:80];
    69: reg_0743 <= imem03_in[47:44];
    72: reg_0743 <= imem03_in[47:44];
    74: reg_0743 <= imem03_in[39:36];
    76: reg_0743 <= imem03_in[39:36];
    79: reg_0743 <= imem03_in[39:36];
    81: reg_0743 <= imem03_in[39:36];
    83: reg_0743 <= imem03_in[39:36];
    85: reg_0743 <= imem03_in[39:36];
    88: reg_0743 <= imem03_in[47:44];
    endcase
  end

  // REG#744の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0744 <= imem03_in[43:40];
    7: reg_0744 <= imem02_in[115:112];
    9: reg_0744 <= imem02_in[115:112];
    11: reg_0744 <= imem07_in[55:52];
    13: reg_0744 <= imem03_in[43:40];
    15: reg_0744 <= imem03_in[43:40];
    17: reg_0744 <= imem02_in[115:112];
    19: reg_0744 <= imem03_in[43:40];
    21: reg_0744 <= imem03_in[43:40];
    23: reg_0744 <= imem02_in[115:112];
    25: reg_0744 <= imem03_in[43:40];
    27: reg_0744 <= imem03_in[87:84];
    30: reg_0744 <= imem03_in[87:84];
    33: reg_0744 <= imem03_in[87:84];
    35: reg_0744 <= imem03_in[43:40];
    37: reg_0744 <= imem03_in[87:84];
    39: reg_0744 <= imem04_in[115:112];
    41: reg_0744 <= imem03_in[43:40];
    43: reg_0744 <= imem07_in[55:52];
    endcase
  end

  // REG#745の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0745 <= imem03_in[79:76];
    7: reg_0745 <= imem03_in[79:76];
    9: reg_0745 <= imem07_in[123:120];
    11: reg_0745 <= imem07_in[95:92];
    13: reg_0745 <= imem00_in[95:92];
    15: reg_0745 <= imem03_in[79:76];
    17: reg_0745 <= imem03_in[79:76];
    19: reg_0745 <= imem03_in[79:76];
    21: reg_0745 <= imem07_in[95:92];
    23: reg_0745 <= imem07_in[95:92];
    25: reg_0745 <= imem07_in[95:92];
    27: reg_0745 <= imem00_in[95:92];
    29: reg_0745 <= imem00_in[95:92];
    31: reg_0745 <= imem07_in[95:92];
    33: reg_0745 <= imem00_in[95:92];
    35: reg_0745 <= imem06_in[107:104];
    38: reg_0745 <= imem00_in[95:92];
    41: reg_0745 <= imem06_in[107:104];
    43: reg_0745 <= imem03_in[79:76];
    45: reg_0745 <= imem06_in[107:104];
    47: reg_0745 <= imem06_in[107:104];
    49: reg_0745 <= imem00_in[95:92];
    51: reg_0745 <= imem06_in[107:104];
    53: reg_0745 <= imem01_in[111:108];
    endcase
  end

  // REG#746の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0746 <= imem03_in[99:96];
    7: reg_0746 <= imem02_in[119:116];
    9: reg_0746 <= imem02_in[119:116];
    11: reg_0746 <= imem03_in[99:96];
    13: reg_0746 <= imem01_in[63:60];
    15: reg_0746 <= imem03_in[99:96];
    17: reg_0746 <= imem03_in[99:96];
    19: reg_0746 <= imem01_in[63:60];
    20: reg_0746 <= op2_01_out;
    57: reg_0746 <= imem01_in[63:60];
    59: reg_0746 <= imem02_in[119:116];
    60: reg_0746 <= op2_01_out;
    endcase
  end

  // REG#747の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0747 <= imem04_in[7:4];
    7: reg_0747 <= imem03_in[31:28];
    9: reg_0747 <= imem03_in[31:28];
    11: reg_0747 <= imem03_in[31:28];
    13: reg_0747 <= imem03_in[31:28];
    16: reg_0747 <= imem03_in[31:28];
    18: reg_0747 <= imem03_in[31:28];
    20: reg_0747 <= imem03_in[31:28];
    22: reg_0747 <= imem03_in[31:28];
    24: reg_0747 <= imem00_in[87:84];
    25: reg_0747 <= op2_02_out;
    31: reg_0747 <= op2_02_out;
    53: reg_0747 <= imem04_in[7:4];
    54: reg_0747 <= op2_02_out;
    85: reg_0747 <= imem00_in[87:84];
    87: reg_0747 <= imem00_in[87:84];
    88: reg_0747 <= op2_02_out;
    endcase
  end

  // REG#748の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0748 <= imem04_in[11:8];
    7: reg_0748 <= imem04_in[11:8];
    9: reg_0748 <= imem00_in[47:44];
    11: reg_0748 <= imem00_in[47:44];
    13: reg_0748 <= imem04_in[11:8];
    16: reg_0748 <= imem04_in[11:8];
    18: reg_0748 <= imem04_in[11:8];
    47: reg_0748 <= imem00_in[47:44];
    49: reg_0748 <= imem04_in[11:8];
    53: reg_0748 <= imem00_in[47:44];
    55: reg_0748 <= imem00_in[47:44];
    90: reg_0748 <= imem00_in[47:44];
    endcase
  end

  // REG#749の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0749 <= imem04_in[23:20];
    7: reg_0749 <= imem03_in[63:60];
    9: reg_0749 <= imem00_in[71:68];
    11: reg_0749 <= imem07_in[127:124];
    13: reg_0749 <= imem03_in[63:60];
    15: reg_0749 <= imem07_in[127:124];
    17: reg_0749 <= imem04_in[23:20];
    20: reg_0749 <= imem04_in[23:20];
    22: reg_0749 <= imem04_in[23:20];
    25: reg_0749 <= imem03_in[63:60];
    27: reg_0749 <= imem03_in[63:60];
    30: reg_0749 <= imem04_in[23:20];
    32: reg_0749 <= imem07_in[127:124];
    34: reg_0749 <= imem04_in[23:20];
    36: reg_0749 <= imem03_in[63:60];
    38: reg_0749 <= imem00_in[71:68];
    40: reg_0749 <= imem00_in[71:68];
    42: reg_0749 <= imem07_in[127:124];
    44: reg_0749 <= imem00_in[71:68];
    46: reg_0749 <= imem00_in[71:68];
    48: reg_0749 <= imem04_in[23:20];
    50: reg_0749 <= imem03_in[63:60];
    53: reg_0749 <= imem07_in[127:124];
    55: reg_0749 <= imem00_in[119:116];
    89: reg_0749 <= imem04_in[23:20];
    93: reg_0749 <= imem00_in[71:68];
    95: reg_0749 <= imem03_in[63:60];
    endcase
  end

  // REG#750の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0750 <= imem04_in[71:68];
    7: reg_0750 <= imem04_in[71:68];
    9: reg_0750 <= imem04_in[71:68];
    11: reg_0750 <= imem02_in[3:0];
    13: reg_0750 <= imem02_in[3:0];
    16: reg_0750 <= imem00_in[39:36];
    18: reg_0750 <= imem00_in[39:36];
    20: reg_0750 <= imem04_in[71:68];
    22: reg_0750 <= imem04_in[71:68];
    25: reg_0750 <= imem00_in[39:36];
    27: reg_0750 <= imem04_in[71:68];
    30: reg_0750 <= imem02_in[3:0];
    32: reg_0750 <= imem04_in[71:68];
    34: reg_0750 <= imem02_in[3:0];
    36: reg_0750 <= imem02_in[3:0];
    39: reg_0750 <= imem04_in[71:68];
    41: reg_0750 <= imem04_in[71:68];
    47: reg_0750 <= imem04_in[71:68];
    49: reg_0750 <= imem05_in[107:104];
    52: reg_0750 <= imem04_in[71:68];
    54: reg_0750 <= imem02_in[3:0];
    56: reg_0750 <= imem02_in[3:0];
    58: reg_0750 <= imem04_in[71:68];
    61: reg_0750 <= imem05_in[107:104];
    67: reg_0750 <= imem00_in[39:36];
    69: reg_0750 <= imem00_in[39:36];
    72: reg_0750 <= imem02_in[3:0];
    84: reg_0750 <= imem02_in[3:0];
    endcase
  end

  // REG#751の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0751 <= imem05_in[23:20];
    7: reg_0751 <= imem04_in[87:84];
    9: reg_0751 <= imem04_in[47:44];
    11: reg_0751 <= imem04_in[87:84];
    13: reg_0751 <= imem04_in[87:84];
    16: reg_0751 <= imem00_in[87:84];
    18: reg_0751 <= imem04_in[47:44];
    43: reg_0751 <= imem05_in[23:20];
    46: reg_0751 <= imem04_in[47:44];
    49: reg_0751 <= imem00_in[87:84];
    51: reg_0751 <= imem05_in[23:20];
    53: reg_0751 <= imem05_in[23:20];
    55: reg_0751 <= imem05_in[23:20];
    57: reg_0751 <= op2_00_out;
    91: reg_0751 <= op2_00_out;
    endcase
  end

  // REG#752の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0752 <= imem06_in[35:32];
    7: reg_0752 <= imem06_in[35:32];
    9: reg_0752 <= imem06_in[35:32];
    33: reg_0752 <= imem04_in[23:20];
    35: reg_0752 <= imem06_in[35:32];
    39: reg_0752 <= imem04_in[23:20];
    42: reg_0752 <= imem04_in[23:20];
    endcase
  end

  // REG#753の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0753 <= imem06_in[63:60];
    7: reg_0753 <= imem05_in[99:96];
    9: reg_0753 <= imem06_in[63:60];
    32: reg_0753 <= imem06_in[63:60];
    38: reg_0753 <= imem05_in[99:96];
    42: reg_0753 <= imem06_in[63:60];
    46: reg_0753 <= imem05_in[99:96];
    49: reg_0753 <= imem06_in[63:60];
    52: reg_0753 <= imem05_in[99:96];
    55: reg_0753 <= imem00_in[111:108];
    90: reg_0753 <= imem00_in[111:108];
    endcase
  end

  // REG#754の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0754 <= imem06_in[111:108];
    7: reg_0754 <= imem06_in[111:108];
    9: reg_0754 <= imem06_in[111:108];
    28: reg_0754 <= imem06_in[87:84];
    31: reg_0754 <= imem06_in[111:108];
    34: reg_0754 <= imem03_in[7:4];
    36: reg_0754 <= imem03_in[7:4];
    39: reg_0754 <= imem06_in[111:108];
    57: reg_0754 <= imem06_in[111:108];
    endcase
  end

  // REG#755の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0755 <= imem07_in[7:4];
    7: reg_0755 <= imem06_in[67:64];
    9: reg_0755 <= imem04_in[63:60];
    11: reg_0755 <= imem07_in[7:4];
    13: reg_0755 <= imem07_in[7:4];
    15: reg_0755 <= imem07_in[7:4];
    17: reg_0755 <= imem07_in[7:4];
    19: reg_0755 <= imem04_in[63:60];
    43: reg_0755 <= imem04_in[63:60];
    46: reg_0755 <= imem06_in[67:64];
    48: reg_0755 <= imem06_in[67:64];
    50: reg_0755 <= imem06_in[67:64];
    53: reg_0755 <= imem06_in[67:64];
    55: reg_0755 <= imem06_in[67:64];
    58: reg_0755 <= imem07_in[7:4];
    60: reg_0755 <= imem05_in[115:112];
    63: reg_0755 <= imem06_in[67:64];
    65: reg_0755 <= imem04_in[63:60];
    67: reg_0755 <= imem06_in[67:64];
    69: reg_0755 <= imem04_in[63:60];
    71: reg_0755 <= imem06_in[67:64];
    90: reg_0755 <= imem06_in[67:64];
    92: reg_0755 <= imem04_in[63:60];
    95: reg_0755 <= imem04_in[63:60];
    endcase
  end

  // REG#756の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0756 <= imem07_in[31:28];
    7: reg_0756 <= imem07_in[19:16];
    9: reg_0756 <= imem04_in[75:72];
    11: reg_0756 <= imem03_in[15:12];
    13: reg_0756 <= imem07_in[31:28];
    15: reg_0756 <= imem07_in[31:28];
    17: reg_0756 <= imem04_in[75:72];
    21: reg_0756 <= imem07_in[19:16];
    23: reg_0756 <= imem00_in[103:100];
    25: reg_0756 <= imem07_in[19:16];
    27: reg_0756 <= imem00_in[103:100];
    29: reg_0756 <= imem07_in[31:28];
    31: reg_0756 <= imem04_in[75:72];
    33: reg_0756 <= imem03_in[15:12];
    35: reg_0756 <= imem07_in[19:16];
    37: reg_0756 <= imem07_in[31:28];
    39: reg_0756 <= imem07_in[31:28];
    42: reg_0756 <= imem00_in[103:100];
    44: reg_0756 <= imem00_in[103:100];
    47: reg_0756 <= imem07_in[19:16];
    49: reg_0756 <= imem04_in[75:72];
    59: reg_0756 <= imem07_in[31:28];
    61: reg_0756 <= imem07_in[95:92];
    63: reg_0756 <= imem00_in[103:100];
    66: reg_0756 <= imem07_in[95:92];
    68: reg_0756 <= imem03_in[15:12];
    70: reg_0756 <= imem03_in[15:12];
    endcase
  end

  // REG#757の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0757 <= imem07_in[99:96];
    7: reg_0757 <= imem07_in[59:56];
    9: reg_0757 <= imem05_in[47:44];
    11: reg_0757 <= imem03_in[19:16];
    13: reg_0757 <= imem03_in[19:16];
    16: reg_0757 <= imem05_in[47:44];
    18: reg_0757 <= imem05_in[47:44];
    20: reg_0757 <= imem05_in[47:44];
    42: reg_0757 <= imem05_in[47:44];
    46: reg_0757 <= imem05_in[47:44];
    48: reg_0757 <= imem07_in[59:56];
    50: reg_0757 <= imem05_in[47:44];
    67: reg_0757 <= imem07_in[59:56];
    69: reg_0757 <= imem03_in[19:16];
    71: reg_0757 <= imem03_in[19:16];
    73: reg_0757 <= imem07_in[59:56];
    76: reg_0757 <= imem07_in[59:56];
    78: reg_0757 <= imem07_in[99:96];
    80: reg_0757 <= imem07_in[59:56];
    84: reg_0757 <= imem07_in[59:56];
    86: reg_0757 <= imem07_in[99:96];
    88: reg_0757 <= imem03_in[19:16];
    endcase
  end

  // REG#758の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0758 <= imem07_in[103:100];
    7: reg_0758 <= imem07_in[83:80];
    9: reg_0758 <= imem07_in[83:80];
    11: reg_0758 <= imem07_in[103:100];
    13: reg_0758 <= imem07_in[83:80];
    15: reg_0758 <= imem07_in[103:100];
    17: reg_0758 <= imem07_in[103:100];
    19: reg_0758 <= imem07_in[103:100];
    21: reg_0758 <= imem02_in[15:12];
    78: reg_0758 <= imem02_in[15:12];
    80: reg_0758 <= imem07_in[43:40];
    84: reg_0758 <= imem07_in[103:100];
    86: reg_0758 <= imem07_in[43:40];
    88: reg_0758 <= imem03_in[27:24];
    endcase
  end

  // REG#759の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0759 <= imem07_in[115:112];
    7: reg_0759 <= imem07_in[119:116];
    9: reg_0759 <= imem07_in[115:112];
    11: reg_0759 <= imem07_in[115:112];
    13: reg_0759 <= imem02_in[7:4];
    16: reg_0759 <= imem02_in[7:4];
    18: reg_0759 <= imem07_in[115:112];
    20: reg_0759 <= imem07_in[119:116];
    22: reg_0759 <= imem02_in[115:112];
    24: reg_0759 <= imem07_in[119:116];
    26: reg_0759 <= imem07_in[115:112];
    28: reg_0759 <= imem07_in[119:116];
    31: reg_0759 <= imem02_in[7:4];
    33: reg_0759 <= imem07_in[119:116];
    35: reg_0759 <= imem06_in[31:28];
    39: reg_0759 <= imem06_in[31:28];
    58: reg_0759 <= imem02_in[115:112];
    60: reg_0759 <= imem06_in[31:28];
    63: reg_0759 <= imem02_in[7:4];
    74: reg_0759 <= imem02_in[115:112];
    79: reg_0759 <= imem07_in[115:112];
    endcase
  end

  // REG#760の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0760 <= imem00_in[31:28];
    7: reg_0760 <= imem00_in[79:76];
    9: reg_0760 <= imem00_in[79:76];
    11: reg_0760 <= imem00_in[31:28];
    13: reg_0760 <= imem00_in[79:76];
    15: reg_0760 <= imem00_in[31:28];
    17: reg_0760 <= imem03_in[39:36];
    19: reg_0760 <= imem04_in[31:28];
    46: reg_0760 <= imem00_in[31:28];
    48: reg_0760 <= imem00_in[31:28];
    50: reg_0760 <= imem00_in[31:28];
    53: reg_0760 <= imem04_in[31:28];
    55: reg_0760 <= imem03_in[39:36];
    89: reg_0760 <= imem00_in[79:76];
    91: reg_0760 <= imem00_in[79:76];
    endcase
  end

  // REG#761の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0761 <= imem00_in[35:32];
    7: reg_0761 <= imem00_in[87:84];
    9: reg_0761 <= imem07_in[23:20];
    11: reg_0761 <= imem00_in[35:32];
    13: reg_0761 <= imem00_in[87:84];
    15: reg_0761 <= imem00_in[35:32];
    17: reg_0761 <= imem07_in[23:20];
    19: reg_0761 <= imem00_in[87:84];
    21: reg_0761 <= imem02_in[31:28];
    83: reg_0761 <= imem02_in[31:28];
    86: reg_0761 <= imem02_in[31:28];
    88: reg_0761 <= imem03_in[43:40];
    endcase
  end

  // REG#762の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0762 <= imem00_in[51:48];
    7: reg_0762 <= imem01_in[23:20];
    9: reg_0762 <= imem00_in[51:48];
    11: reg_0762 <= imem01_in[23:20];
    26: reg_0762 <= imem02_in[119:116];
    49: reg_0762 <= imem01_in[23:20];
    70: reg_0762 <= imem01_in[23:20];
    72: reg_0762 <= imem02_in[119:116];
    82: reg_0762 <= imem00_in[51:48];
    84: reg_0762 <= imem00_in[51:48];
    86: reg_0762 <= imem00_in[51:48];
    88: reg_0762 <= imem00_in[51:48];
    91: reg_0762 <= imem00_in[51:48];
    endcase
  end

  // REG#763の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0763 <= imem00_in[55:52];
    7: reg_0763 <= imem00_in[55:52];
    9: reg_0763 <= imem00_in[55:52];
    11: reg_0763 <= imem03_in[95:92];
    13: reg_0763 <= imem03_in[95:92];
    15: reg_0763 <= imem03_in[95:92];
    17: reg_0763 <= imem00_in[55:52];
    19: reg_0763 <= imem04_in[19:16];
    44: reg_0763 <= imem00_in[55:52];
    46: reg_0763 <= imem04_in[19:16];
    50: reg_0763 <= imem00_in[55:52];
    52: reg_0763 <= imem04_in[19:16];
    54: reg_0763 <= imem00_in[55:52];
    56: reg_0763 <= imem00_in[55:52];
    58: reg_0763 <= imem00_in[55:52];
    60: reg_0763 <= imem03_in[95:92];
    62: reg_0763 <= imem03_in[95:92];
    64: reg_0763 <= imem03_in[95:92];
    66: reg_0763 <= imem04_in[19:16];
    68: reg_0763 <= imem00_in[55:52];
    70: reg_0763 <= imem00_in[55:52];
    72: reg_0763 <= imem02_in[99:96];
    82: reg_0763 <= imem00_in[55:52];
    84: reg_0763 <= imem00_in[55:52];
    86: reg_0763 <= imem03_in[95:92];
    88: reg_0763 <= imem03_in[95:92];
    endcase
  end

  // REG#764の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0764 <= imem00_in[107:104];
    7: reg_0764 <= imem00_in[107:104];
    9: reg_0764 <= imem07_in[71:68];
    11: reg_0764 <= imem03_in[119:116];
    13: reg_0764 <= imem00_in[107:104];
    15: reg_0764 <= imem00_in[107:104];
    17: reg_0764 <= imem03_in[119:116];
    19: reg_0764 <= imem04_in[3:0];
    46: reg_0764 <= imem04_in[3:0];
    49: reg_0764 <= imem04_in[115:112];
    57: reg_0764 <= imem00_in[107:104];
    59: reg_0764 <= imem04_in[3:0];
    endcase
  end

  // REG#765の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0765 <= imem01_in[19:16];
    7: reg_0765 <= imem01_in[27:24];
    9: reg_0765 <= imem01_in[27:24];
    12: reg_0765 <= imem01_in[27:24];
    14: reg_0765 <= imem01_in[27:24];
    16: reg_0765 <= imem01_in[27:24];
    18: reg_0765 <= imem01_in[27:24];
    20: reg_0765 <= imem01_in[19:16];
    22: reg_0765 <= imem03_in[23:20];
    24: reg_0765 <= imem01_in[99:96];
    26: reg_0765 <= imem03_in[23:20];
    28: reg_0765 <= imem03_in[23:20];
    66: reg_0765 <= imem01_in[99:96];
    69: reg_0765 <= imem03_in[23:20];
    72: reg_0765 <= imem02_in[115:112];
    82: reg_0765 <= imem02_in[115:112];
    84: reg_0765 <= imem02_in[115:112];
    endcase
  end

  // REG#766の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0766 <= imem01_in[63:60];
    7: reg_0766 <= imem01_in[87:84];
    9: reg_0766 <= imem01_in[87:84];
    11: reg_0766 <= imem01_in[63:60];
    26: reg_0766 <= imem01_in[63:60];
    27: reg_0766 <= op2_00_out;
    36: reg_0766 <= op2_00_out;
    66: reg_0766 <= op2_00_out;
    78: reg_0766 <= op2_00_out;
    endcase
  end

  // REG#767の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0767 <= imem02_in[3:0];
    7: reg_0767 <= imem02_in[3:0];
    9: reg_0767 <= imem07_in[75:72];
    11: reg_0767 <= imem07_in[75:72];
    13: reg_0767 <= imem07_in[75:72];
    16: reg_0767 <= imem07_in[75:72];
    18: reg_0767 <= imem07_in[75:72];
    20: reg_0767 <= imem07_in[75:72];
    22: reg_0767 <= imem03_in[87:84];
    24: reg_0767 <= imem07_in[75:72];
    26: reg_0767 <= imem03_in[87:84];
    28: reg_0767 <= imem03_in[87:84];
    70: reg_0767 <= imem03_in[87:84];
    endcase
  end

  // REG#768の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0768 <= imem02_in[7:4];
    7: reg_0768 <= imem02_in[7:4];
    9: reg_0768 <= imem00_in[7:4];
    11: reg_0768 <= imem04_in[11:8];
    13: reg_0768 <= imem00_in[7:4];
    16: reg_0768 <= imem00_in[7:4];
    18: reg_0768 <= imem00_in[7:4];
    20: reg_0768 <= imem02_in[7:4];
    23: reg_0768 <= imem00_in[7:4];
    25: reg_0768 <= imem02_in[7:4];
    27: reg_0768 <= imem02_in[7:4];
    29: reg_0768 <= imem00_in[7:4];
    31: reg_0768 <= imem04_in[11:8];
    33: reg_0768 <= imem00_in[7:4];
    35: reg_0768 <= imem04_in[11:8];
    38: reg_0768 <= imem02_in[7:4];
    41: reg_0768 <= imem02_in[7:4];
    43: reg_0768 <= imem02_in[7:4];
    47: reg_0768 <= imem02_in[7:4];
    49: reg_0768 <= imem00_in[7:4];
    51: reg_0768 <= imem02_in[7:4];
    55: reg_0768 <= imem00_in[27:24];
    96: reg_0768 <= imem02_in[7:4];
    endcase
  end

  // REG#769の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0769 <= imem02_in[47:44];
    7: reg_0769 <= imem01_in[127:124];
    9: reg_0769 <= imem00_in[119:116];
    11: reg_0769 <= imem02_in[47:44];
    13: reg_0769 <= imem03_in[35:32];
    15: reg_0769 <= imem02_in[47:44];
    17: reg_0769 <= imem01_in[127:124];
    19: reg_0769 <= imem02_in[47:44];
    21: reg_0769 <= imem00_in[119:116];
    23: reg_0769 <= imem02_in[47:44];
    25: reg_0769 <= imem01_in[127:124];
    48: reg_0769 <= imem00_in[119:116];
    51: reg_0769 <= imem01_in[127:124];
    53: reg_0769 <= imem01_in[19:16];
    endcase
  end

  // REG#770の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0770 <= imem02_in[103:100];
    7: reg_0770 <= imem02_in[123:120];
    9: reg_0770 <= imem02_in[123:120];
    11: reg_0770 <= imem04_in[15:12];
    13: reg_0770 <= imem04_in[3:0];
    16: reg_0770 <= imem04_in[15:12];
    17: reg_0770 <= op2_00_out;
    45: reg_0770 <= op2_00_out;
    54: reg_0770 <= op2_00_out;
    82: reg_0770 <= op2_00_out;
    89: reg_0770 <= imem04_in[15:12];
    90: reg_0770 <= op2_00_out;
    endcase
  end

  // REG#771の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0771 <= imem02_in[111:108];
    7: reg_0771 <= imem02_in[111:108];
    9: reg_0771 <= imem02_in[111:108];
    11: reg_0771 <= imem04_in[51:48];
    13: reg_0771 <= imem04_in[71:68];
    15: reg_0771 <= imem02_in[111:108];
    17: reg_0771 <= imem02_in[111:108];
    18: reg_0771 <= op2_00_out;
    49: reg_0771 <= imem02_in[111:108];
    52: reg_0771 <= op2_00_out;
    76: reg_0771 <= op2_00_out;
    endcase
  end

  // REG#772の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0772 <= imem02_in[127:124];
    7: reg_0772 <= imem02_in[127:124];
    9: reg_0772 <= imem01_in[43:40];
    12: reg_0772 <= imem02_in[123:120];
    14: reg_0772 <= imem02_in[123:120];
    16: reg_0772 <= imem02_in[123:120];
    18: reg_0772 <= imem02_in[127:124];
    20: reg_0772 <= imem02_in[127:124];
    22: reg_0772 <= imem02_in[123:120];
    24: reg_0772 <= imem02_in[123:120];
    26: reg_0772 <= imem02_in[123:120];
    52: reg_0772 <= imem02_in[127:124];
    endcase
  end

  // REG#773の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0773 <= imem03_in[59:56];
    7: reg_0773 <= imem04_in[3:0];
    9: reg_0773 <= imem03_in[59:56];
    11: reg_0773 <= imem03_in[59:56];
    13: reg_0773 <= imem03_in[59:56];
    16: reg_0773 <= imem04_in[3:0];
    18: reg_0773 <= imem04_in[95:92];
    48: reg_0773 <= imem03_in[59:56];
    50: reg_0773 <= imem04_in[95:92];
    52: reg_0773 <= imem03_in[59:56];
    54: reg_0773 <= imem04_in[95:92];
    56: reg_0773 <= imem03_in[59:56];
    58: reg_0773 <= imem04_in[95:92];
    61: reg_0773 <= imem00_in[27:24];
    63: reg_0773 <= imem04_in[3:0];
    65: reg_0773 <= imem00_in[27:24];
    68: reg_0773 <= imem03_in[59:56];
    70: reg_0773 <= imem03_in[59:56];
    endcase
  end

  // REG#774の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0774 <= imem04_in[31:28];
    7: reg_0774 <= imem04_in[75:72];
    9: reg_0774 <= imem04_in[31:28];
    11: reg_0774 <= imem05_in[35:32];
    13: reg_0774 <= imem04_in[75:72];
    16: reg_0774 <= imem04_in[75:72];
    18: reg_0774 <= imem04_in[75:72];
    44: reg_0774 <= imem04_in[75:72];
    48: reg_0774 <= imem04_in[31:28];
    50: reg_0774 <= imem05_in[35:32];
    67: reg_0774 <= imem05_in[35:32];
    70: reg_0774 <= imem05_in[35:32];
    72: reg_0774 <= imem04_in[75:72];
    74: reg_0774 <= imem04_in[31:28];
    76: reg_0774 <= imem04_in[31:28];
    78: reg_0774 <= imem05_in[35:32];
    80: reg_0774 <= imem04_in[31:28];
    82: reg_0774 <= imem04_in[75:72];
    85: reg_0774 <= imem05_in[35:32];
    87: reg_0774 <= imem04_in[75:72];
    89: reg_0774 <= imem05_in[35:32];
    91: reg_0774 <= imem05_in[35:32];
    93: reg_0774 <= imem04_in[75:72];
    endcase
  end

  // REG#775の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0775 <= imem04_in[59:56];
    7: reg_0775 <= imem04_in[59:56];
    9: reg_0775 <= imem01_in[63:60];
    12: reg_0775 <= imem04_in[59:56];
    14: reg_0775 <= imem02_in[23:20];
    16: reg_0775 <= imem01_in[63:60];
    18: reg_0775 <= imem02_in[23:20];
    20: reg_0775 <= imem02_in[23:20];
    22: reg_0775 <= imem01_in[63:60];
    24: reg_0775 <= imem01_in[63:60];
    27: reg_0775 <= imem01_in[63:60];
    29: reg_0775 <= imem01_in[63:60];
    31: reg_0775 <= imem04_in[59:56];
    33: reg_0775 <= imem01_in[63:60];
    35: reg_0775 <= imem04_in[59:56];
    38: reg_0775 <= imem01_in[63:60];
    41: reg_0775 <= op2_02_out;
    85: reg_0775 <= imem02_in[23:20];
    endcase
  end

  // REG#776の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0776 <= imem04_in[67:64];
    7: reg_0776 <= imem04_in[107:104];
    9: reg_0776 <= imem04_in[67:64];
    11: reg_0776 <= imem04_in[107:104];
    13: reg_0776 <= imem04_in[67:64];
    15: reg_0776 <= imem04_in[67:64];
    17: reg_0776 <= imem04_in[67:64];
    21: reg_0776 <= imem02_in[27:24];
    85: reg_0776 <= imem02_in[27:24];
    endcase
  end

  // REG#777の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0777 <= imem04_in[79:76];
    7: reg_0777 <= imem04_in[79:76];
    9: reg_0777 <= imem01_in[55:52];
    12: reg_0777 <= imem03_in[59:56];
    14: reg_0777 <= imem02_in[107:104];
    16: reg_0777 <= imem01_in[7:4];
    18: reg_0777 <= imem04_in[79:76];
    45: reg_0777 <= imem01_in[55:52];
    47: reg_0777 <= imem02_in[107:104];
    49: reg_0777 <= imem04_in[79:76];
    57: reg_0777 <= imem03_in[59:56];
    59: reg_0777 <= imem04_in[79:76];
    endcase
  end

  // REG#778の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0778 <= imem04_in[99:96];
    7: reg_0778 <= imem05_in[107:104];
    9: reg_0778 <= imem01_in[47:44];
    12: reg_0778 <= imem04_in[99:96];
    14: reg_0778 <= imem05_in[107:104];
    16: reg_0778 <= imem05_in[107:104];
    18: reg_0778 <= imem05_in[107:104];
    20: reg_0778 <= imem01_in[47:44];
    22: reg_0778 <= imem05_in[107:104];
    24: reg_0778 <= imem04_in[99:96];
    85: reg_0778 <= imem02_in[51:48];
    endcase
  end

  // REG#779の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0779 <= imem04_in[103:100];
    7: reg_0779 <= imem05_in[111:108];
    9: reg_0779 <= imem01_in[15:12];
    12: reg_0779 <= imem03_in[79:76];
    14: reg_0779 <= imem05_in[111:108];
    16: reg_0779 <= imem03_in[79:76];
    18: reg_0779 <= imem03_in[79:76];
    20: reg_0779 <= imem03_in[79:76];
    22: reg_0779 <= imem04_in[103:100];
    25: reg_0779 <= imem01_in[15:12];
    49: reg_0779 <= imem01_in[15:12];
    70: reg_0779 <= imem03_in[79:76];
    endcase
  end

  // REG#780の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0780 <= imem04_in[127:124];
    7: reg_0780 <= imem06_in[39:36];
    9: reg_0780 <= imem06_in[39:36];
    26: reg_0780 <= imem04_in[127:124];
    28: reg_0780 <= imem06_in[39:36];
    30: reg_0780 <= imem06_in[39:36];
    32: reg_0780 <= imem06_in[39:36];
    37: reg_0780 <= imem06_in[39:36];
    61: reg_0780 <= imem06_in[39:36];
    72: reg_0780 <= imem04_in[127:124];
    74: reg_0780 <= imem05_in[11:8];
    endcase
  end

  // REG#781の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0781 <= imem05_in[31:28];
    7: reg_0781 <= imem06_in[71:68];
    9: reg_0781 <= imem06_in[71:68];
    33: reg_0781 <= imem05_in[31:28];
    35: reg_0781 <= imem05_in[31:28];
    39: reg_0781 <= imem06_in[71:68];
    58: reg_0781 <= imem06_in[71:68];
    83: reg_0781 <= imem06_in[71:68];
    86: reg_0781 <= imem06_in[127:124];
    endcase
  end

  // REG#782の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0782 <= imem05_in[35:32];
    7: reg_0782 <= imem06_in[91:88];
    9: reg_0782 <= imem06_in[91:88];
    33: reg_0782 <= imem05_in[83:80];
    35: reg_0782 <= imem06_in[91:88];
    39: reg_0782 <= imem06_in[91:88];
    60: reg_0782 <= imem05_in[35:32];
    63: reg_0782 <= imem06_in[91:88];
    65: reg_0782 <= imem05_in[83:80];
    69: reg_0782 <= imem02_in[79:76];
    71: reg_0782 <= imem06_in[91:88];
    89: reg_0782 <= imem06_in[91:88];
    endcase
  end

  // REG#783の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0783 <= imem05_in[39:36];
    7: reg_0783 <= imem06_in[99:96];
    9: reg_0783 <= imem06_in[99:96];
    33: reg_0783 <= imem06_in[47:44];
    35: reg_0783 <= imem06_in[47:44];
    37: reg_0783 <= imem05_in[39:36];
    39: reg_0783 <= imem06_in[99:96];
    57: reg_0783 <= imem05_in[39:36];
    60: reg_0783 <= imem06_in[99:96];
    63: reg_0783 <= imem03_in[51:48];
    65: reg_0783 <= imem03_in[51:48];
    67: reg_0783 <= imem06_in[47:44];
    69: reg_0783 <= imem02_in[87:84];
    72: reg_0783 <= imem02_in[87:84];
    82: reg_0783 <= imem06_in[99:96];
    84: reg_0783 <= imem06_in[47:44];
    86: reg_0783 <= imem06_in[99:96];
    endcase
  end

  // REG#784の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0784 <= imem05_in[75:72];
    7: reg_0784 <= imem07_in[63:60];
    9: reg_0784 <= imem05_in[75:72];
    11: reg_0784 <= imem07_in[63:60];
    13: reg_0784 <= imem07_in[63:60];
    16: reg_0784 <= imem07_in[63:60];
    18: reg_0784 <= imem07_in[63:60];
    20: reg_0784 <= imem07_in[63:60];
    22: reg_0784 <= imem05_in[35:32];
    24: reg_0784 <= imem07_in[63:60];
    26: reg_0784 <= imem07_in[63:60];
    28: reg_0784 <= imem03_in[51:48];
    66: reg_0784 <= imem05_in[75:72];
    75: reg_0784 <= imem07_in[63:60];
    80: reg_0784 <= imem05_in[35:32];
    86: reg_0784 <= imem05_in[35:32];
    88: reg_0784 <= imem03_in[51:48];
    endcase
  end

  // REG#785の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0785 <= imem05_in[91:88];
    7: reg_0785 <= imem05_in[91:88];
    9: reg_0785 <= imem05_in[91:88];
    11: reg_0785 <= imem05_in[91:88];
    14: reg_0785 <= imem03_in[39:36];
    16: reg_0785 <= imem03_in[11:8];
    18: reg_0785 <= imem05_in[91:88];
    20: reg_0785 <= imem05_in[91:88];
    52: reg_0785 <= imem05_in[91:88];
    54: reg_0785 <= imem05_in[91:88];
    56: reg_0785 <= imem05_in[91:88];
    61: reg_0785 <= imem03_in[11:8];
    63: reg_0785 <= imem03_in[11:8];
    65: reg_0785 <= imem03_in[39:36];
    67: reg_0785 <= imem03_in[39:36];
    69: reg_0785 <= imem05_in[91:88];
    71: reg_0785 <= imem03_in[39:36];
    73: reg_0785 <= imem03_in[39:36];
    75: reg_0785 <= imem03_in[39:36];
    77: reg_0785 <= imem03_in[39:36];
    79: reg_0785 <= imem03_in[11:8];
    84: reg_0785 <= imem03_in[11:8];
    86: reg_0785 <= imem03_in[39:36];
    88: reg_0785 <= imem03_in[11:8];
    endcase
  end

  // REG#786の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0786 <= imem05_in[95:92];
    7: reg_0786 <= imem07_in[111:108];
    9: reg_0786 <= imem01_in[11:8];
    13: reg_0786 <= imem01_in[11:8];
    15: reg_0786 <= imem05_in[95:92];
    17: reg_0786 <= imem05_in[95:92];
    19: reg_0786 <= imem07_in[111:108];
    21: reg_0786 <= imem01_in[11:8];
    23: reg_0786 <= imem05_in[95:92];
    25: reg_0786 <= imem01_in[11:8];
    49: reg_0786 <= imem01_in[11:8];
    66: reg_0786 <= imem05_in[95:92];
    78: reg_0786 <= imem01_in[11:8];
    80: reg_0786 <= imem05_in[95:92];
    84: reg_0786 <= imem05_in[95:92];
    86: reg_0786 <= imem07_in[111:108];
    88: reg_0786 <= imem01_in[11:8];
    90: reg_0786 <= imem01_in[11:8];
    92: reg_0786 <= imem05_in[95:92];
    96: reg_0786 <= imem01_in[11:8];
    endcase
  end

  // REG#787の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0787 <= imem06_in[11:8];
    7: reg_0787 <= imem00_in[15:12];
    9: reg_0787 <= imem06_in[11:8];
    33: reg_0787 <= imem06_in[11:8];
    35: reg_0787 <= imem06_in[83:80];
    39: reg_0787 <= imem00_in[15:12];
    42: reg_0787 <= imem06_in[11:8];
    44: reg_0787 <= imem00_in[15:12];
    48: reg_0787 <= imem06_in[11:8];
    50: reg_0787 <= imem06_in[11:8];
    52: reg_0787 <= imem00_in[15:12];
    54: reg_0787 <= imem06_in[11:8];
    58: reg_0787 <= imem00_in[15:12];
    60: reg_0787 <= imem06_in[83:80];
    63: reg_0787 <= imem04_in[39:36];
    68: reg_0787 <= imem00_in[15:12];
    70: reg_0787 <= imem06_in[83:80];
    73: reg_0787 <= imem00_in[15:12];
    75: reg_0787 <= imem06_in[83:80];
    77: reg_0787 <= imem06_in[11:8];
    79: reg_0787 <= imem00_in[15:12];
    81: reg_0787 <= imem06_in[83:80];
    83: reg_0787 <= imem06_in[83:80];
    86: reg_0787 <= imem06_in[11:8];
    endcase
  end

  // REG#788の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0788 <= imem07_in[43:40];
    7: reg_0788 <= imem02_in[79:76];
    9: reg_0788 <= imem01_in[3:0];
    13: reg_0788 <= imem02_in[79:76];
    15: reg_0788 <= imem02_in[79:76];
    17: reg_0788 <= imem01_in[3:0];
    19: reg_0788 <= imem01_in[3:0];
    21: reg_0788 <= imem07_in[43:40];
    23: reg_0788 <= imem01_in[3:0];
    25: reg_0788 <= imem07_in[43:40];
    26: reg_0788 <= op2_02_out;
    35: reg_0788 <= op2_02_out;
    66: reg_0788 <= imem07_in[43:40];
    68: reg_0788 <= imem02_in[79:76];
    70: reg_0788 <= imem07_in[43:40];
    72: reg_0788 <= imem07_in[43:40];
    74: reg_0788 <= imem02_in[79:76];
    77: reg_0788 <= imem02_in[79:76];
    79: reg_0788 <= imem01_in[3:0];
    80: reg_0788 <= op2_02_out;
    85: reg_0788 <= imem02_in[79:76];
    endcase
  end

  // REG#789の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0789 <= imem07_in[127:124];
    7: reg_0789 <= imem02_in[99:96];
    9: reg_0789 <= imem01_in[31:28];
    12: reg_0789 <= op2_00_out;
    29: reg_0789 <= imem07_in[127:124];
    31: reg_0789 <= imem07_in[127:124];
    33: reg_0789 <= imem07_in[127:124];
    34: reg_0789 <= op2_00_out;
    61: reg_0789 <= imem02_in[99:96];
    63: reg_0789 <= imem01_in[31:28];
    64: reg_0789 <= op2_00_out;
    74: reg_0789 <= imem01_in[31:28];
    76: reg_0789 <= imem02_in[99:96];
    78: reg_0789 <= imem07_in[127:124];
    80: reg_0789 <= op2_00_out;
    83: reg_0789 <= op2_00_out;
    92: reg_0789 <= imem01_in[31:28];
    endcase
  end

  // REG#790の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0790 <= imem00_in[103:100];
    7: reg_0790 <= imem00_in[103:100];
    9: reg_0790 <= imem01_in[7:4];
    12: reg_0790 <= op2_02_out;
    31: reg_0790 <= imem00_in[103:100];
    32: reg_0790 <= op2_02_out;
    55: reg_0790 <= op2_02_out;
    87: reg_0790 <= op2_02_out;
    endcase
  end

  // REG#791の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0791 <= imem01_in[51:48];
    7: reg_0791 <= imem01_in[51:48];
    9: reg_0791 <= imem01_in[51:48];
    14: reg_0791 <= imem01_in[51:48];
    16: reg_0791 <= imem01_in[51:48];
    17: reg_0791 <= op2_01_out;
    47: reg_0791 <= imem01_in[51:48];
    50: reg_0791 <= op2_01_out;
    71: reg_0791 <= op2_01_out;
    98: reg_0791 <= op2_01_out;
    endcase
  end

  // REG#792の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0792 <= imem01_in[95:92];
    7: reg_0792 <= imem03_in[51:48];
    9: reg_0792 <= imem01_in[95:92];
    13: reg_0792 <= imem03_in[51:48];
    15: reg_0792 <= imem03_in[51:48];
    17: reg_0792 <= imem01_in[95:92];
    19: reg_0792 <= imem03_in[51:48];
    21: reg_0792 <= imem02_in[47:44];
    86: reg_0792 <= imem06_in[35:32];
    endcase
  end

  // REG#793の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0793 <= imem01_in[111:108];
    7: reg_0793 <= imem01_in[111:108];
    9: reg_0793 <= imem01_in[111:108];
    14: reg_0793 <= imem01_in[111:108];
    16: reg_0793 <= imem01_in[111:108];
    18: reg_0793 <= imem01_in[111:108];
    20: reg_0793 <= imem02_in[123:120];
    23: reg_0793 <= imem02_in[123:120];
    25: reg_0793 <= imem02_in[123:120];
    28: reg_0793 <= imem03_in[19:16];
    69: reg_0793 <= imem01_in[111:108];
    94: reg_0793 <= imem01_in[111:108];
    endcase
  end

  // REG#794の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0794 <= imem03_in[47:44];
    7: reg_0794 <= imem03_in[95:92];
    9: reg_0794 <= imem01_in[39:36];
    13: reg_0794 <= imem01_in[39:36];
    15: reg_0794 <= imem01_in[39:36];
    17: reg_0794 <= imem07_in[95:92];
    18: reg_0794 <= op2_01_out;
    50: reg_0794 <= imem03_in[95:92];
    52: reg_0794 <= imem03_in[47:44];
    53: reg_0794 <= op2_01_out;
    81: reg_0794 <= imem03_in[95:92];
    83: reg_0794 <= imem07_in[95:92];
    84: reg_0794 <= op2_01_out;
    endcase
  end

  // REG#795の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0795 <= imem03_in[111:108];
    7: reg_0795 <= imem04_in[35:32];
    9: reg_0795 <= imem01_in[67:64];
    14: reg_0795 <= imem03_in[111:108];
    16: reg_0795 <= imem03_in[43:40];
    18: reg_0795 <= imem03_in[43:40];
    19: reg_0795 <= op1_15_out;
    23: reg_0795 <= imem03_in[43:40];
    24: reg_0795 <= op1_15_out;
    28: reg_0795 <= imem03_in[43:40];
    70: reg_0795 <= imem04_in[35:32];
    72: reg_0795 <= imem03_in[43:40];
    74: reg_0795 <= imem05_in[59:56];
    endcase
  end

  // REG#796の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0796 <= imem05_in[3:0];
    7: reg_0796 <= imem04_in[43:40];
    8: reg_0796 <= op2_01_out;
    16: reg_0796 <= op2_01_out;
    43: reg_0796 <= op2_01_out;
    48: reg_0796 <= op2_01_out;
    65: reg_0796 <= op2_01_out;
    76: reg_0796 <= op2_01_out;
    endcase
  end

  // REG#797の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0797 <= imem05_in[79:76];
    7: reg_0797 <= imem05_in[79:76];
    8: reg_0797 <= op2_02_out;
    17: reg_0797 <= op2_02_out;
    48: reg_0797 <= op2_02_out;
    66: reg_0797 <= op2_02_out;
    81: reg_0797 <= imem05_in[79:76];
    83: reg_0797 <= imem05_in[79:76];
    84: reg_0797 <= op2_02_out;
    endcase
  end

  // REG#798の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0798 <= imem05_in[119:116];
    7: reg_0798 <= imem05_in[119:116];
    9: reg_0798 <= imem06_in[115:112];
    31: reg_0798 <= imem01_in[23:20];
    33: reg_0798 <= imem01_in[23:20];
    35: reg_0798 <= imem01_in[23:20];
    37: reg_0798 <= imem01_in[23:20];
    39: reg_0798 <= imem01_in[23:20];
    41: reg_0798 <= imem01_in[23:20];
    93: reg_0798 <= imem01_in[23:20];
    96: reg_0798 <= imem01_in[23:20];
    endcase
  end

  // REG#799の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0799 <= imem06_in[19:16];
    7: reg_0799 <= imem04_in[51:48];
    9: reg_0799 <= imem06_in[7:4];
    31: reg_0799 <= imem06_in[7:4];
    34: reg_0799 <= imem03_in[103:100];
    36: reg_0799 <= imem06_in[7:4];
    40: reg_0799 <= imem04_in[51:48];
    42: reg_0799 <= imem04_in[11:8];
    96: reg_0799 <= imem03_in[103:100];
    endcase
  end

  // REG#800の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0800 <= imem06_in[27:24];
    7: reg_0800 <= imem06_in[27:24];
    9: reg_0800 <= imem06_in[27:24];
    28: reg_0800 <= imem06_in[27:24];
    31: reg_0800 <= imem05_in[43:40];
    33: reg_0800 <= imem07_in[95:92];
    34: reg_0800 <= op2_02_out;
    63: reg_0800 <= imem07_in[95:92];
    65: reg_0800 <= imem05_in[43:40];
    69: reg_0800 <= imem06_in[27:24];
    70: reg_0800 <= op2_02_out;
    94: reg_0800 <= op2_02_out;
    endcase
  end

  // REG#801の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0801 <= imem06_in[55:52];
    7: reg_0801 <= imem04_in[55:52];
    9: reg_0801 <= imem06_in[51:48];
    31: reg_0801 <= imem06_in[51:48];
    32: reg_0801 <= op2_00_out;
    53: reg_0801 <= op2_00_out;
    79: reg_0801 <= op2_02_out;
    endcase
  end

  // REG#802の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0802 <= imem06_in[59:56];
    7: reg_0802 <= imem04_in[83:80];
    9: reg_0802 <= imem06_in[59:56];
    34: reg_0802 <= imem04_in[15:12];
    36: reg_0802 <= imem04_in[83:80];
    38: reg_0802 <= imem04_in[83:80];
    40: reg_0802 <= imem06_in[59:56];
    42: reg_0802 <= imem04_in[15:12];
    endcase
  end

  // REG#803の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0803 <= imem06_in[83:80];
    6: reg_0803 <= op1_00_out;
    9: reg_0803 <= imem06_in[83:80];
    32: reg_0803 <= op1_00_out;
    34: reg_0803 <= op1_00_out;
    36: reg_0803 <= op1_00_out;
    38: reg_0803 <= op1_00_out;
    40: reg_0803 <= op1_00_out;
    42: reg_0803 <= op1_00_out;
    44: reg_0803 <= op1_00_out;
    46: reg_0803 <= op1_00_out;
    48: reg_0803 <= op1_00_out;
    50: reg_0803 <= op1_00_out;
    52: reg_0803 <= op1_00_out;
    54: reg_0803 <= op1_00_out;
    56: reg_0803 <= op1_00_out;
    58: reg_0803 <= op1_00_out;
    60: reg_0803 <= op1_00_out;
    62: reg_0803 <= op1_00_out;
    64: reg_0803 <= op1_00_out;
    66: reg_0803 <= op1_00_out;
    69: reg_0803 <= imem04_in[75:72];
    72: reg_0803 <= imem02_in[23:20];
    82: reg_0803 <= op1_00_out;
    84: reg_0803 <= op1_00_out;
    86: reg_0803 <= op1_00_out;
    88: reg_0803 <= op1_00_out;
    90: reg_0803 <= op1_00_out;
    92: reg_0803 <= op1_00_out;
    94: reg_0803 <= op1_00_out;
    96: reg_0803 <= op1_00_out;
    endcase
  end

  // REG#804の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0804 <= imem06_in[95:92];
    6: reg_0804 <= op1_01_out;
    8: reg_0804 <= op1_01_out;
    10: reg_0804 <= op1_01_out;
    13: reg_0804 <= imem06_in[95:92];
    15: reg_0804 <= imem06_in[95:92];
    17: reg_0804 <= imem06_in[95:92];
    18: reg_0804 <= op1_01_out;
    20: reg_0804 <= op1_01_out;
    23: reg_0804 <= imem06_in[95:92];
    24: reg_0804 <= op1_01_out;
    27: reg_0804 <= imem06_in[95:92];
    29: reg_0804 <= imem06_in[95:92];
    58: reg_0804 <= imem06_in[95:92];
    87: reg_0804 <= imem06_in[95:92];
    89: reg_0804 <= imem06_in[95:92];
    endcase
  end

  // REG#805の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0805 <= imem07_in[3:0];
    7: reg_0805 <= imem07_in[3:0];
    9: reg_0805 <= imem06_in[87:84];
    31: reg_0805 <= imem06_in[11:8];
    33: reg_0805 <= imem07_in[3:0];
    35: reg_0805 <= imem06_in[87:84];
    39: reg_0805 <= imem07_in[35:32];
    41: reg_0805 <= imem07_in[3:0];
    43: reg_0805 <= imem07_in[3:0];
    endcase
  end

  // REG#806の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0806 <= imem07_in[27:24];
    7: reg_0806 <= imem07_in[27:24];
    9: reg_0806 <= imem07_in[27:24];
    11: reg_0806 <= imem06_in[75:72];
    13: reg_0806 <= imem07_in[27:24];
    16: reg_0806 <= imem03_in[115:112];
    18: reg_0806 <= imem03_in[115:112];
    20: reg_0806 <= imem05_in[35:32];
    49: reg_0806 <= imem05_in[35:32];
    53: reg_0806 <= imem07_in[27:24];
    55: reg_0806 <= imem07_in[27:24];
    57: reg_0806 <= imem05_in[35:32];
    60: reg_0806 <= imem06_in[75:72];
    62: reg_0806 <= imem07_in[27:24];
    64: reg_0806 <= imem05_in[35:32];
    69: reg_0806 <= imem04_in[91:88];
    72: reg_0806 <= imem07_in[27:24];
    74: reg_0806 <= imem05_in[35:32];
    endcase
  end

  // REG#807の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0807 <= imem00_in[3:0];
    6: reg_0807 <= op1_02_out;
    8: reg_0807 <= op1_02_out;
    11: reg_0807 <= imem00_in[3:0];
    13: reg_0807 <= imem00_in[3:0];
    15: reg_0807 <= op1_02_out;
    18: reg_0807 <= imem00_in[3:0];
    20: reg_0807 <= imem00_in[3:0];
    22: reg_0807 <= imem05_in[79:76];
    24: reg_0807 <= imem00_in[3:0];
    26: reg_0807 <= imem00_in[3:0];
    28: reg_0807 <= imem03_in[79:76];
    69: reg_0807 <= imem06_in[19:16];
    71: reg_0807 <= imem06_in[19:16];
    89: reg_0807 <= imem06_in[19:16];
    93: reg_0807 <= imem00_in[3:0];
    endcase
  end

  // REG#808の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0808 <= imem00_in[91:88];
    7: reg_0808 <= imem00_in[91:88];
    9: reg_0808 <= imem06_in[31:28];
    32: reg_0808 <= imem06_in[31:28];
    38: reg_0808 <= imem06_in[31:28];
    42: reg_0808 <= imem04_in[91:88];
    endcase
  end

  // REG#809の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0809 <= imem01_in[43:40];
    6: reg_0809 <= op1_03_out;
    8: reg_0809 <= op1_03_out;
    10: reg_0809 <= op1_03_out;
    14: reg_0809 <= imem01_in[43:40];
    15: reg_0809 <= op1_03_out;
    18: reg_0809 <= imem01_in[43:40];
    19: reg_0809 <= op1_03_out;
    21: reg_0809 <= op1_03_out;
    23: reg_0809 <= op1_03_out;
    25: reg_0809 <= op1_03_out;
    27: reg_0809 <= op1_03_out;
    29: reg_0809 <= op1_03_out;
    32: reg_0809 <= imem01_in[43:40];
    33: reg_0809 <= op1_03_out;
    38: reg_0809 <= imem01_in[43:40];
    40: reg_0809 <= imem01_in[43:40];
    42: reg_0809 <= imem04_in[111:108];
    endcase
  end

  // REG#810の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0810 <= imem01_in[67:64];
    6: reg_0810 <= op1_04_out;
    8: reg_0810 <= op1_04_out;
    10: reg_0810 <= op1_04_out;
    12: reg_0810 <= op1_04_out;
    14: reg_0810 <= op1_04_out;
    17: reg_0810 <= imem01_in[67:64];
    19: reg_0810 <= imem01_in[67:64];
    21: reg_0810 <= imem01_in[67:64];
    23: reg_0810 <= imem02_in[27:24];
    25: reg_0810 <= imem01_in[67:64];
    47: reg_0810 <= imem01_in[67:64];
    52: reg_0810 <= imem01_in[67:64];
    54: reg_0810 <= imem01_in[67:64];
    59: reg_0810 <= imem01_in[67:64];
    61: reg_0810 <= imem00_in[111:108];
    63: reg_0810 <= imem02_in[3:0];
    72: reg_0810 <= imem02_in[27:24];
    83: reg_0810 <= imem02_in[27:24];
    87: reg_0810 <= imem02_in[27:24];
    89: reg_0810 <= imem02_in[27:24];
    91: reg_0810 <= imem00_in[111:108];
    endcase
  end

  // REG#811の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0811 <= imem01_in[75:72];
    6: reg_0811 <= op1_05_out;
    8: reg_0811 <= op1_05_out;
    10: reg_0811 <= op1_05_out;
    12: reg_0811 <= op1_05_out;
    15: reg_0811 <= imem01_in[75:72];
    16: reg_0811 <= op1_05_out;
    18: reg_0811 <= op1_05_out;
    20: reg_0811 <= op1_05_out;
    23: reg_0811 <= imem03_in[119:116];
    25: reg_0811 <= imem01_in[103:100];
    48: reg_0811 <= imem01_in[103:100];
    50: reg_0811 <= imem01_in[103:100];
    51: reg_0811 <= op1_05_out;
    53: reg_0811 <= op1_05_out;
    55: reg_0811 <= op1_05_out;
    57: reg_0811 <= op1_05_out;
    59: reg_0811 <= op1_05_out;
    61: reg_0811 <= op1_05_out;
    63: reg_0811 <= op1_05_out;
    65: reg_0811 <= op1_05_out;
    67: reg_0811 <= op1_05_out;
    69: reg_0811 <= op1_05_out;
    71: reg_0811 <= op1_05_out;
    74: reg_0811 <= imem01_in[75:72];
    77: reg_0811 <= imem01_in[103:100];
    79: reg_0811 <= imem01_in[75:72];
    81: reg_0811 <= imem03_in[119:116];
    84: reg_0811 <= imem01_in[103:100];
    86: reg_0811 <= imem06_in[119:116];
    endcase
  end

  // REG#812の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0812 <= imem01_in[123:120];
    7: reg_0812 <= imem01_in[123:120];
    9: reg_0812 <= imem01_in[123:120];
    14: reg_0812 <= imem03_in[95:92];
    16: reg_0812 <= imem03_in[95:92];
    18: reg_0812 <= op2_02_out;
    50: reg_0812 <= op2_02_out;
    72: reg_0812 <= op2_02_out;
    endcase
  end

  // REG#813の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0813 <= imem02_in[31:28];
    7: reg_0813 <= imem02_in[31:28];
    9: reg_0813 <= imem02_in[31:28];
    11: reg_0813 <= imem02_in[31:28];
    13: reg_0813 <= imem02_in[31:28];
    15: reg_0813 <= imem02_in[31:28];
    17: reg_0813 <= imem00_in[103:100];
    20: reg_0813 <= imem05_in[59:56];
    48: reg_0813 <= imem05_in[59:56];
    50: reg_0813 <= imem05_in[59:56];
    67: reg_0813 <= imem05_in[59:56];
    70: reg_0813 <= imem05_in[59:56];
    72: reg_0813 <= imem02_in[31:28];
    85: reg_0813 <= imem00_in[103:100];
    87: reg_0813 <= imem05_in[59:56];
    endcase
  end

  // REG#814の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0814 <= imem02_in[51:48];
    7: reg_0814 <= imem02_in[51:48];
    9: reg_0814 <= imem02_in[51:48];
    11: reg_0814 <= imem02_in[51:48];
    13: reg_0814 <= imem02_in[51:48];
    15: reg_0814 <= imem02_in[51:48];
    17: reg_0814 <= imem03_in[31:28];
    19: reg_0814 <= imem03_in[31:28];
    21: reg_0814 <= imem02_in[51:48];
    86: reg_0814 <= imem06_in[7:4];
    endcase
  end

  // REG#815の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0815 <= imem02_in[87:84];
    6: reg_0815 <= op1_06_out;
    8: reg_0815 <= op1_06_out;
    10: reg_0815 <= op1_06_out;
    12: reg_0815 <= op1_06_out;
    14: reg_0815 <= op1_06_out;
    17: reg_0815 <= imem02_in[87:84];
    18: reg_0815 <= op1_06_out;
    20: reg_0815 <= op1_06_out;
    23: reg_0815 <= imem04_in[95:92];
    25: reg_0815 <= imem02_in[87:84];
    28: reg_0815 <= imem04_in[95:92];
    30: reg_0815 <= imem02_in[87:84];
    33: reg_0815 <= imem04_in[95:92];
    35: reg_0815 <= imem04_in[95:92];
    37: reg_0815 <= imem02_in[87:84];
    39: reg_0815 <= imem02_in[87:84];
    42: reg_0815 <= imem04_in[95:92];
    endcase
  end

  // REG#816の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0816 <= imem03_in[87:84];
    7: reg_0816 <= imem03_in[87:84];
    9: reg_0816 <= imem03_in[87:84];
    11: reg_0816 <= imem03_in[87:84];
    14: reg_0816 <= imem06_in[19:16];
    16: reg_0816 <= imem03_in[119:116];
    18: reg_0816 <= imem06_in[19:16];
    20: reg_0816 <= imem05_in[71:68];
    49: reg_0816 <= imem04_in[39:36];
    57: reg_0816 <= imem04_in[39:36];
    59: reg_0816 <= imem03_in[119:116];
    61: reg_0816 <= imem06_in[19:16];
    72: reg_0816 <= imem03_in[87:84];
    74: reg_0816 <= imem05_in[71:68];
    endcase
  end

  // REG#817の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0817 <= imem03_in[7:4];
    8: reg_0817 <= imem06_in[91:88];
    10: reg_0817 <= imem03_in[7:4];
    12: reg_0817 <= imem03_in[7:4];
    14: reg_0817 <= imem03_in[7:4];
    16: reg_0817 <= imem03_in[7:4];
    18: reg_0817 <= imem03_in[7:4];
    20: reg_0817 <= imem03_in[7:4];
    22: reg_0817 <= imem06_in[39:36];
    24: reg_0817 <= imem03_in[7:4];
    26: reg_0817 <= imem02_in[95:92];
    52: reg_0817 <= imem03_in[7:4];
    54: reg_0817 <= imem02_in[95:92];
    57: reg_0817 <= imem06_in[91:88];
    endcase
  end

  // REG#818の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0818 <= imem03_in[95:92];
    8: reg_0818 <= imem07_in[43:40];
    10: reg_0818 <= imem07_in[43:40];
    12: reg_0818 <= imem07_in[43:40];
    14: reg_0818 <= imem07_in[43:40];
    16: reg_0818 <= imem07_in[43:40];
    18: reg_0818 <= imem07_in[43:40];
    20: reg_0818 <= imem03_in[95:92];
    22: reg_0818 <= imem07_in[43:40];
    24: reg_0818 <= imem03_in[119:116];
    26: reg_0818 <= imem02_in[91:88];
    52: reg_0818 <= imem02_in[91:88];
    endcase
  end

  // REG#819の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0819 <= imem05_in[115:112];
    8: reg_0819 <= imem05_in[115:112];
    10: reg_0819 <= imem05_in[119:116];
    12: reg_0819 <= imem05_in[119:116];
    17: reg_0819 <= imem04_in[119:116];
    20: reg_0819 <= imem05_in[115:112];
    50: reg_0819 <= imem05_in[115:112];
    66: reg_0819 <= imem05_in[115:112];
    79: reg_0819 <= imem05_in[119:116];
    88: reg_0819 <= imem03_in[15:12];
    endcase
  end

  // REG#820の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0820 <= imem03_in[27:24];
    8: reg_0820 <= imem03_in[27:24];
    10: reg_0820 <= imem07_in[27:24];
    12: reg_0820 <= imem03_in[99:96];
    14: reg_0820 <= imem00_in[7:4];
    16: reg_0820 <= imem03_in[27:24];
    18: reg_0820 <= imem03_in[99:96];
    20: reg_0820 <= imem03_in[99:96];
    22: reg_0820 <= imem07_in[27:24];
    24: reg_0820 <= imem03_in[27:24];
    26: reg_0820 <= imem03_in[99:96];
    28: reg_0820 <= imem03_in[99:96];
    70: reg_0820 <= imem03_in[99:96];
    endcase
  end

  // REG#821の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0821 <= imem05_in[15:12];
    8: reg_0821 <= imem07_in[59:56];
    10: reg_0821 <= imem07_in[59:56];
    12: reg_0821 <= imem07_in[59:56];
    14: reg_0821 <= imem05_in[15:12];
    16: reg_0821 <= imem05_in[15:12];
    20: reg_0821 <= imem05_in[15:12];
    49: reg_0821 <= imem05_in[15:12];
    53: reg_0821 <= imem01_in[107:104];
    endcase
  end

  // REG#822の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0822 <= imem05_in[55:52];
    8: reg_0822 <= imem07_in[75:72];
    10: reg_0822 <= imem05_in[55:52];
    12: reg_0822 <= imem05_in[55:52];
    16: reg_0822 <= imem04_in[23:20];
    19: reg_0822 <= imem07_in[75:72];
    21: reg_0822 <= imem07_in[75:72];
    23: reg_0822 <= imem05_in[107:104];
    25: reg_0822 <= imem05_in[55:52];
    28: reg_0822 <= imem03_in[127:124];
    72: reg_0822 <= imem05_in[55:52];
    74: reg_0822 <= imem07_in[75:72];
    78: reg_0822 <= imem03_in[127:124];
    80: reg_0822 <= imem07_in[75:72];
    83: reg_0822 <= imem07_in[75:72];
    86: reg_0822 <= imem06_in[87:84];
    endcase
  end

  // REG#823の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0823 <= imem03_in[3:0];
    8: reg_0823 <= imem00_in[27:24];
    10: reg_0823 <= imem00_in[27:24];
    12: reg_0823 <= imem00_in[27:24];
    14: reg_0823 <= imem03_in[3:0];
    16: reg_0823 <= imem00_in[27:24];
    18: reg_0823 <= imem00_in[27:24];
    20: reg_0823 <= imem00_in[27:24];
    22: reg_0823 <= imem00_in[27:24];
    24: reg_0823 <= imem03_in[3:0];
    26: reg_0823 <= imem03_in[3:0];
    28: reg_0823 <= imem03_in[3:0];
    70: reg_0823 <= imem03_in[3:0];
    endcase
  end

  // REG#824の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0824 <= imem03_in[119:116];
    8: reg_0824 <= imem03_in[119:116];
    10: reg_0824 <= imem07_in[31:28];
    12: reg_0824 <= imem07_in[31:28];
    14: reg_0824 <= imem07_in[31:28];
    16: reg_0824 <= imem07_in[31:28];
    18: reg_0824 <= imem07_in[31:28];
    20: reg_0824 <= imem07_in[31:28];
    22: reg_0824 <= imem04_in[83:80];
    25: reg_0824 <= imem07_in[31:28];
    27: reg_0824 <= imem03_in[119:116];
    29: reg_0824 <= imem04_in[83:80];
    31: reg_0824 <= imem03_in[119:116];
    55: reg_0824 <= imem07_in[31:28];
    57: reg_0824 <= imem07_in[31:28];
    59: reg_0824 <= imem04_in[83:80];
    endcase
  end

  // REG#825の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0825 <= imem03_in[83:80];
    8: reg_0825 <= imem00_in[71:68];
    10: reg_0825 <= imem03_in[83:80];
    12: reg_0825 <= imem04_in[7:4];
    14: reg_0825 <= imem00_in[35:32];
    16: reg_0825 <= imem04_in[7:4];
    18: reg_0825 <= imem03_in[83:80];
    20: reg_0825 <= imem05_in[87:84];
    53: reg_0825 <= imem03_in[83:80];
    55: reg_0825 <= imem00_in[35:32];
    88: reg_0825 <= imem00_in[71:68];
    90: reg_0825 <= imem03_in[83:80];
    endcase
  end

  // REG#826の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0826 <= imem05_in[19:16];
    8: reg_0826 <= imem00_in[79:76];
    10: reg_0826 <= imem00_in[3:0];
    12: reg_0826 <= imem05_in[19:16];
    20: reg_0826 <= imem05_in[19:16];
    50: reg_0826 <= imem05_in[19:16];
    67: reg_0826 <= imem05_in[19:16];
    69: reg_0826 <= imem05_in[19:16];
    71: reg_0826 <= imem00_in[3:0];
    73: reg_0826 <= imem05_in[19:16];
    90: reg_0826 <= imem00_in[3:0];
    endcase
  end

  // REG#827の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0827 <= imem05_in[43:40];
    8: reg_0827 <= imem00_in[83:80];
    10: reg_0827 <= imem00_in[83:80];
    12: reg_0827 <= imem05_in[43:40];
    20: reg_0827 <= imem05_in[43:40];
    51: reg_0827 <= imem00_in[83:80];
    53: reg_0827 <= imem01_in[75:72];
    endcase
  end

  // REG#828の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0828 <= imem05_in[87:84];
    8: reg_0828 <= imem00_in[107:104];
    10: reg_0828 <= imem00_in[107:104];
    12: reg_0828 <= imem05_in[87:84];
    21: reg_0828 <= imem00_in[107:104];
    23: reg_0828 <= imem00_in[107:104];
    25: reg_0828 <= imem01_in[79:76];
    49: reg_0828 <= imem05_in[87:84];
    52: reg_0828 <= imem01_in[79:76];
    55: reg_0828 <= imem00_in[107:104];
    90: reg_0828 <= imem01_in[79:76];
    93: reg_0828 <= imem00_in[107:104];
    95: reg_0828 <= imem05_in[87:84];
    endcase
  end

  // REG#829の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0829 <= imem05_in[111:108];
    8: reg_0829 <= imem01_in[43:40];
    10: reg_0829 <= imem05_in[111:108];
    12: reg_0829 <= imem04_in[75:72];
    14: reg_0829 <= imem01_in[31:28];
    16: reg_0829 <= imem04_in[119:116];
    18: reg_0829 <= imem05_in[111:108];
    20: reg_0829 <= imem04_in[75:72];
    22: reg_0829 <= imem04_in[75:72];
    25: reg_0829 <= imem05_in[111:108];
    27: reg_0829 <= imem05_in[111:108];
    30: reg_0829 <= imem04_in[119:116];
    32: reg_0829 <= imem05_in[111:108];
    34: reg_0829 <= imem01_in[31:28];
    36: reg_0829 <= imem01_in[31:28];
    39: reg_0829 <= imem04_in[75:72];
    41: reg_0829 <= imem01_in[43:40];
    94: reg_0829 <= imem01_in[43:40];
    endcase
  end

  // REG#830の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0830 <= imem03_in[11:8];
    8: reg_0830 <= imem01_in[51:48];
    10: reg_0830 <= imem01_in[51:48];
    39: reg_0830 <= imem01_in[51:48];
    41: reg_0830 <= imem01_in[51:48];
    94: reg_0830 <= imem01_in[51:48];
    endcase
  end

  // REG#831の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0831 <= imem03_in[103:100];
    8: reg_0831 <= imem03_in[103:100];
    10: reg_0831 <= imem03_in[103:100];
    12: reg_0831 <= imem03_in[103:100];
    14: reg_0831 <= imem01_in[115:112];
    16: reg_0831 <= imem04_in[127:124];
    18: reg_0831 <= imem01_in[115:112];
    20: reg_0831 <= imem05_in[119:116];
    51: reg_0831 <= imem03_in[103:100];
    53: reg_0831 <= imem04_in[127:124];
    55: reg_0831 <= imem05_in[119:116];
    58: reg_0831 <= imem03_in[103:100];
    60: reg_0831 <= imem01_in[115:112];
    63: reg_0831 <= imem01_in[115:112];
    65: reg_0831 <= imem01_in[115:112];
    67: reg_0831 <= imem01_in[115:112];
    69: reg_0831 <= imem01_in[115:112];
    82: reg_0831 <= imem03_in[103:100];
    85: reg_0831 <= imem01_in[115:112];
    87: reg_0831 <= imem05_in[119:116];
    endcase
  end

  // REG#832の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0832 <= imem05_in[123:120];
    8: reg_0832 <= imem02_in[27:24];
    10: reg_0832 <= imem02_in[27:24];
    12: reg_0832 <= imem05_in[123:120];
    20: reg_0832 <= imem05_in[111:108];
    51: reg_0832 <= imem05_in[111:108];
    53: reg_0832 <= imem01_in[7:4];
    endcase
  end

  // REG#833の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0833 <= imem03_in[35:32];
    8: reg_0833 <= imem02_in[51:48];
    10: reg_0833 <= imem00_in[39:36];
    12: reg_0833 <= imem02_in[51:48];
    14: reg_0833 <= imem02_in[43:40];
    16: reg_0833 <= imem02_in[43:40];
    18: reg_0833 <= imem03_in[35:32];
    20: reg_0833 <= imem03_in[35:32];
    22: reg_0833 <= imem04_in[7:4];
    25: reg_0833 <= imem02_in[43:40];
    28: reg_0833 <= imem03_in[35:32];
    72: reg_0833 <= imem02_in[51:48];
    85: reg_0833 <= imem03_in[35:32];
    87: reg_0833 <= imem02_in[43:40];
    89: reg_0833 <= imem00_in[39:36];
    93: reg_0833 <= imem02_in[43:40];
    endcase
  end

  // REG#834の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0834 <= imem05_in[7:4];
    8: reg_0834 <= imem05_in[7:4];
    10: reg_0834 <= imem05_in[7:4];
    12: reg_0834 <= imem05_in[7:4];
    20: reg_0834 <= imem05_in[7:4];
    49: reg_0834 <= imem04_in[19:16];
    60: reg_0834 <= imem04_in[19:16];
    63: reg_0834 <= imem04_in[19:16];
    65: reg_0834 <= imem05_in[7:4];
    69: reg_0834 <= imem06_in[43:40];
    71: reg_0834 <= imem06_in[43:40];
    89: reg_0834 <= imem05_in[7:4];
    91: reg_0834 <= imem04_in[19:16];
    93: reg_0834 <= imem04_in[19:16];
    endcase
  end

  // REG#835の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0835 <= imem05_in[27:24];
    8: reg_0835 <= imem05_in[27:24];
    10: reg_0835 <= imem05_in[27:24];
    12: reg_0835 <= imem05_in[27:24];
    20: reg_0835 <= imem05_in[27:24];
    54: reg_0835 <= imem05_in[27:24];
    56: reg_0835 <= imem05_in[27:24];
    61: reg_0835 <= imem05_in[27:24];
    65: reg_0835 <= imem05_in[27:24];
    69: reg_0835 <= imem06_in[59:56];
    71: reg_0835 <= imem06_in[59:56];
    87: reg_0835 <= op2_01_out;
    endcase
  end

  // REG#836の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0836 <= imem05_in[71:68];
    8: reg_0836 <= imem02_in[55:52];
    10: reg_0836 <= imem03_in[55:52];
    12: reg_0836 <= imem05_in[71:68];
    21: reg_0836 <= imem03_in[55:52];
    23: reg_0836 <= imem06_in[75:72];
    26: reg_0836 <= imem06_in[75:72];
    28: reg_0836 <= imem03_in[83:80];
    71: reg_0836 <= imem02_in[55:52];
    73: reg_0836 <= imem02_in[55:52];
    75: reg_0836 <= imem03_in[83:80];
    77: reg_0836 <= imem03_in[55:52];
    79: reg_0836 <= imem02_in[55:52];
    81: reg_0836 <= imem02_in[55:52];
    83: reg_0836 <= imem06_in[75:72];
    86: reg_0836 <= imem02_in[55:52];
    88: reg_0836 <= imem03_in[55:52];
    endcase
  end

  // REG#837の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0837 <= imem05_in[103:100];
    8: reg_0837 <= imem02_in[115:112];
    10: reg_0837 <= imem05_in[103:100];
    12: reg_0837 <= imem07_in[19:16];
    14: reg_0837 <= imem05_in[103:100];
    16: reg_0837 <= imem07_in[19:16];
    18: reg_0837 <= imem05_in[103:100];
    20: reg_0837 <= imem02_in[115:112];
    22: reg_0837 <= imem07_in[19:16];
    24: reg_0837 <= imem05_in[103:100];
    26: reg_0837 <= imem02_in[3:0];
    52: reg_0837 <= imem02_in[3:0];
    endcase
  end

  // REG#838の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0838 <= op1_00_out;
    8: reg_0838 <= op1_00_out;
    10: reg_0838 <= op1_00_out;
    12: reg_0838 <= op1_00_out;
    14: reg_0838 <= op1_00_out;
    16: reg_0838 <= op1_00_out;
    18: reg_0838 <= op1_00_out;
    20: reg_0838 <= op1_00_out;
    22: reg_0838 <= op1_00_out;
    24: reg_0838 <= op1_00_out;
    26: reg_0838 <= op1_00_out;
    28: reg_0838 <= op1_00_out;
    30: reg_0838 <= op1_00_out;
    34: reg_0838 <= imem05_in[7:4];
    39: reg_0838 <= imem07_in[123:120];
    41: reg_0838 <= imem07_in[123:120];
    43: reg_0838 <= imem07_in[123:120];
    endcase
  end

  // REG#839の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0839 <= op1_01_out;
    11: reg_0839 <= imem07_in[11:8];
    12: reg_0839 <= op1_01_out;
    14: reg_0839 <= op1_01_out;
    16: reg_0839 <= op1_01_out;
    20: reg_0839 <= imem07_in[11:8];
    21: reg_0839 <= op2_01_out;
    59: reg_0839 <= op2_01_out;
    endcase
  end

  // REG#840の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0840 <= op1_02_out;
    11: reg_0840 <= op1_02_out;
    13: reg_0840 <= op1_02_out;
    16: reg_0840 <= imem05_in[83:80];
    19: reg_0840 <= imem05_in[83:80];
    21: reg_0840 <= imem02_in[83:80];
    85: reg_0840 <= op2_02_out;
    endcase
  end

  // REG#841の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0841 <= op1_03_out;
    13: reg_0841 <= op1_03_out;
    16: reg_0841 <= imem06_in[103:100];
    17: reg_0841 <= op1_03_out;
    19: reg_0841 <= op2_00_out;
    52: reg_0841 <= imem06_in[103:100];
    55: reg_0841 <= imem00_in[11:8];
    92: reg_0841 <= op2_00_out;
    endcase
  end

  // REG#842の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0842 <= op1_04_out;
    13: reg_0842 <= op1_04_out;
    15: reg_0842 <= op1_04_out;
    17: reg_0842 <= op1_04_out;
    19: reg_0842 <= op1_04_out;
    21: reg_0842 <= op1_04_out;
    23: reg_0842 <= op1_04_out;
    26: reg_0842 <= imem02_in[19:16];
    55: reg_0842 <= imem00_in[67:64];
    95: reg_0842 <= imem00_in[67:64];
    endcase
  end

  // REG#843の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0843 <= op1_05_out;
    14: reg_0843 <= op1_05_out;
    17: reg_0843 <= imem04_in[123:120];
    20: reg_0843 <= imem04_in[123:120];
    21: reg_0843 <= op1_05_out;
    23: reg_0843 <= op1_05_out;
    25: reg_0843 <= op1_05_out;
    27: reg_0843 <= op1_05_out;
    29: reg_0843 <= op1_05_out;
    31: reg_0843 <= op1_05_out;
    33: reg_0843 <= op1_05_out;
    35: reg_0843 <= op1_05_out;
    37: reg_0843 <= op1_05_out;
    39: reg_0843 <= op1_05_out;
    41: reg_0843 <= op1_05_out;
    43: reg_0843 <= op1_05_out;
    45: reg_0843 <= op1_05_out;
    47: reg_0843 <= op1_05_out;
    49: reg_0843 <= op1_05_out;
    52: reg_0843 <= imem04_in[123:120];
    55: reg_0843 <= imem00_in[39:36];
    94: reg_0843 <= imem04_in[123:120];
    endcase
  end

  // REG#844の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0844 <= op1_06_out;
    15: reg_0844 <= op1_06_out;
    17: reg_0844 <= op1_06_out;
    19: reg_0844 <= op1_06_out;
    21: reg_0844 <= op1_06_out;
    23: reg_0844 <= op1_06_out;
    25: reg_0844 <= op1_06_out;
    28: reg_0844 <= imem03_in[111:108];
    72: reg_0844 <= imem02_in[11:8];
    84: reg_0844 <= imem02_in[11:8];
    endcase
  end

  // REG#845の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0845 <= op1_07_out;
    16: reg_0845 <= op1_07_out;
    18: reg_0845 <= op1_07_out;
    20: reg_0845 <= op1_07_out;
    22: reg_0845 <= op1_07_out;
    25: reg_0845 <= op1_07_out;
    27: reg_0845 <= op1_07_out;
    31: reg_0845 <= imem07_in[43:40];
    33: reg_0845 <= imem07_in[43:40];
    36: reg_0845 <= imem07_in[43:40];
    39: reg_0845 <= imem01_in[115:112];
    41: reg_0845 <= imem07_in[43:40];
    44: reg_0845 <= imem07_in[43:40];
    48: reg_0845 <= imem07_in[43:40];
    55: reg_0845 <= imem07_in[43:40];
    57: reg_0845 <= imem01_in[115:112];
    60: reg_0845 <= imem06_in[55:52];
    63: reg_0845 <= imem02_in[47:44];
    73: reg_0845 <= imem07_in[43:40];
    75: reg_0845 <= imem02_in[47:44];
    77: reg_0845 <= imem01_in[115:112];
    79: reg_0845 <= imem04_in[107:104];
    82: reg_0845 <= imem06_in[55:52];
    85: reg_0845 <= imem04_in[107:104];
    87: reg_0845 <= imem02_in[47:44];
    89: reg_0845 <= imem02_in[47:44];
    91: reg_0845 <= imem01_in[115:112];
    93: reg_0845 <= imem07_in[43:40];
    95: reg_0845 <= imem01_in[115:112];
    endcase
  end

  // REG#846の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0846 <= op1_08_out;
    18: reg_0846 <= op1_08_out;
    20: reg_0846 <= op1_08_out;
    22: reg_0846 <= op1_08_out;
    25: reg_0846 <= op1_08_out;
    27: reg_0846 <= op1_08_out;
    29: reg_0846 <= op1_08_out;
    31: reg_0846 <= op1_08_out;
    33: reg_0846 <= op1_08_out;
    35: reg_0846 <= op1_08_out;
    37: reg_0846 <= op1_08_out;
    39: reg_0846 <= op1_08_out;
    41: reg_0846 <= op1_08_out;
    43: reg_0846 <= op1_08_out;
    45: reg_0846 <= op1_08_out;
    47: reg_0846 <= op1_08_out;
    49: reg_0846 <= op1_08_out;
    51: reg_0846 <= op1_08_out;
    53: reg_0846 <= op1_08_out;
    55: reg_0846 <= op1_08_out;
    57: reg_0846 <= op1_08_out;
    59: reg_0846 <= op1_08_out;
    61: reg_0846 <= op1_08_out;
    63: reg_0846 <= op1_08_out;
    65: reg_0846 <= op1_08_out;
    67: reg_0846 <= op1_08_out;
    69: reg_0846 <= op1_08_out;
    72: reg_0846 <= imem02_in[59:56];
    83: reg_0846 <= op1_08_out;
    85: reg_0846 <= op1_08_out;
    87: reg_0846 <= op1_08_out;
    89: reg_0846 <= op1_08_out;
    91: reg_0846 <= op1_08_out;
    93: reg_0846 <= op1_08_out;
    95: reg_0846 <= op1_08_out;
    97: reg_0846 <= op1_08_out;
    endcase
  end

  // REG#847の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0847 <= op1_09_out;
    19: reg_0847 <= op1_09_out;
    21: reg_0847 <= op1_09_out;
    23: reg_0847 <= op1_09_out;
    25: reg_0847 <= op1_09_out;
    28: reg_0847 <= imem03_in[7:4];
    70: reg_0847 <= op1_09_out;
    72: reg_0847 <= op1_09_out;
    74: reg_0847 <= op1_09_out;
    77: reg_0847 <= imem03_in[7:4];
    78: reg_0847 <= op1_09_out;
    80: reg_0847 <= op1_09_out;
    85: reg_0847 <= imem03_in[7:4];
    88: reg_0847 <= op1_09_out;
    90: reg_0847 <= op1_09_out;
    93: reg_0847 <= imem03_in[7:4];
    95: reg_0847 <= imem03_in[7:4];
    endcase
  end

  // REG#848の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0848 <= op1_10_out;
    20: reg_0848 <= op1_10_out;
    22: reg_0848 <= op1_10_out;
    24: reg_0848 <= op1_10_out;
    26: reg_0848 <= op1_10_out;
    28: reg_0848 <= op1_10_out;
    30: reg_0848 <= op1_10_out;
    32: reg_0848 <= op1_10_out;
    34: reg_0848 <= op1_10_out;
    36: reg_0848 <= op1_10_out;
    38: reg_0848 <= op1_10_out;
    42: reg_0848 <= imem04_in[19:16];
    endcase
  end

  // REG#849の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0849 <= op1_11_out;
    23: reg_0849 <= op1_11_out;
    25: reg_0849 <= op1_11_out;
    27: reg_0849 <= op1_11_out;
    29: reg_0849 <= op1_11_out;
    31: reg_0849 <= op1_11_out;
    33: reg_0849 <= op1_11_out;
    35: reg_0849 <= op1_11_out;
    39: reg_0849 <= imem01_in[27:24];
    47: reg_0849 <= imem01_in[27:24];
    51: reg_0849 <= op1_11_out;
    53: reg_0849 <= op1_11_out;
    61: reg_0849 <= imem01_in[79:76];
    63: reg_0849 <= imem01_in[79:76];
    66: reg_0849 <= imem01_in[79:76];
    68: reg_0849 <= imem01_in[79:76];
    71: reg_0849 <= imem01_in[79:76];
    73: reg_0849 <= imem01_in[79:76];
    75: reg_0849 <= op1_11_out;
    78: reg_0849 <= imem01_in[27:24];
    82: reg_0849 <= imem01_in[79:76];
    83: reg_0849 <= op1_11_out;
    85: reg_0849 <= op1_11_out;
    88: reg_0849 <= imem01_in[79:76];
    92: reg_0849 <= imem01_in[27:24];
    endcase
  end

  // REG#850の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0850 <= op1_12_out;
    29: reg_0850 <= op1_12_out;
    31: reg_0850 <= op1_12_out;
    35: reg_0850 <= op1_12_out;
    38: reg_0850 <= op1_12_out;
    42: reg_0850 <= imem04_in[35:32];
    endcase
  end

  // REG#851の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0851 <= op1_13_out;
    29: reg_0851 <= op1_13_out;
    32: reg_0851 <= op1_13_out;
    35: reg_0851 <= op1_13_out;
    38: reg_0851 <= op1_13_out;
    44: reg_0851 <= op1_13_out;
    47: reg_0851 <= op1_13_out;
    49: reg_0851 <= op1_13_out;
    52: reg_0851 <= op1_13_out;
    57: reg_0851 <= op1_13_out;
    60: reg_0851 <= op1_13_out;
    64: reg_0851 <= op1_13_out;
    67: reg_0851 <= op1_13_out;
    70: reg_0851 <= op1_13_out;
    74: reg_0851 <= imem05_in[99:96];
    endcase
  end

  // REG#852の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0852 <= op1_14_out;
    30: reg_0852 <= op1_14_out;
    33: reg_0852 <= op1_14_out;
    37: reg_0852 <= op1_14_out;
    43: reg_0852 <= op1_14_out;
    47: reg_0852 <= op1_14_out;
    49: reg_0852 <= op1_14_out;
    52: reg_0852 <= op1_14_out;
    55: reg_0852 <= op1_14_out;
    58: reg_0852 <= op1_14_out;
    61: reg_0852 <= op1_14_out;
    65: reg_0852 <= op1_14_out;
    68: reg_0852 <= op1_14_out;
    71: reg_0852 <= op1_14_out;
    74: reg_0852 <= op1_14_out;
    78: reg_0852 <= op1_14_out;
    81: reg_0852 <= op1_14_out;
    84: reg_0852 <= op1_14_out;
    87: reg_0852 <= op1_14_out;
    91: reg_0852 <= op1_14_out;
    endcase
  end

  // REG#853の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0853 <= op1_15_out;
    32: reg_0853 <= op1_15_out;
    34: reg_0853 <= op1_15_out;
    38: reg_0853 <= op1_15_out;
    41: reg_0853 <= op1_15_out;
    44: reg_0853 <= op1_15_out;
    47: reg_0853 <= op1_15_out;
    52: reg_0853 <= op1_15_out;
    56: reg_0853 <= op1_15_out;
    59: reg_0853 <= op1_15_out;
    62: reg_0853 <= op1_15_out;
    65: reg_0853 <= op1_15_out;
    68: reg_0853 <= op1_15_out;
    71: reg_0853 <= op1_15_out;
    74: reg_0853 <= op1_15_out;
    78: reg_0853 <= op1_15_out;
    81: reg_0853 <= op1_15_out;
    84: reg_0853 <= op1_15_out;
    87: reg_0853 <= op1_15_out;
    90: reg_0853 <= op1_15_out;
    93: reg_0853 <= op1_15_out;
    96: reg_0853 <= op1_15_out;
    endcase
  end

  // REG#854の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0854 <= imem04_in[67:64];
    8: reg_0854 <= imem03_in[115:112];
    10: reg_0854 <= imem03_in[111:108];
    12: reg_0854 <= imem07_in[91:88];
    14: reg_0854 <= imem02_in[111:108];
    16: reg_0854 <= imem04_in[67:64];
    18: reg_0854 <= imem04_in[67:64];
    45: reg_0854 <= imem02_in[111:108];
    57: reg_0854 <= imem02_in[111:108];
    59: reg_0854 <= imem04_in[67:64];
    endcase
  end

  // REG#855の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0855 <= imem04_in[103:100];
    8: reg_0855 <= imem04_in[103:100];
    10: reg_0855 <= imem04_in[91:88];
    12: reg_0855 <= imem07_in[95:92];
    14: reg_0855 <= imem02_in[127:124];
    16: reg_0855 <= imem02_in[127:124];
    18: reg_0855 <= imem04_in[91:88];
    45: reg_0855 <= imem07_in[95:92];
    48: reg_0855 <= imem04_in[91:88];
    54: reg_0855 <= imem02_in[127:124];
    56: reg_0855 <= imem04_in[91:88];
    58: reg_0855 <= imem04_in[91:88];
    61: reg_0855 <= imem04_in[103:100];
    63: reg_0855 <= imem02_in[119:116];
    74: reg_0855 <= imem04_in[103:100];
    76: reg_0855 <= imem04_in[103:100];
    78: reg_0855 <= imem02_in[119:116];
    80: reg_0855 <= imem02_in[119:116];
    82: reg_0855 <= imem04_in[103:100];
    84: reg_0855 <= imem02_in[119:116];
    endcase
  end

  // REG#856の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0856 <= imem04_in[107:104];
    8: reg_0856 <= imem04_in[19:16];
    10: reg_0856 <= imem04_in[107:104];
    12: reg_0856 <= imem04_in[107:104];
    14: reg_0856 <= imem04_in[107:104];
    16: reg_0856 <= imem00_in[43:40];
    18: reg_0856 <= imem04_in[107:104];
    39: reg_0856 <= imem06_in[55:52];
    56: reg_0856 <= imem06_in[55:52];
    59: reg_0856 <= imem04_in[107:104];
    96: reg_0856 <= imem04_in[107:104];
    endcase
  end

  // REG#857の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0857 <= imem06_in[3:0];
    8: reg_0857 <= imem06_in[3:0];
    11: reg_0857 <= imem00_in[119:116];
    13: reg_0857 <= imem06_in[3:0];
    15: reg_0857 <= imem06_in[3:0];
    17: reg_0857 <= imem04_in[87:84];
    21: reg_0857 <= imem06_in[3:0];
    23: reg_0857 <= imem00_in[3:0];
    26: reg_0857 <= imem02_in[87:84];
    52: reg_0857 <= imem06_in[3:0];
    54: reg_0857 <= imem02_in[87:84];
    57: reg_0857 <= imem02_in[87:84];
    60: reg_0857 <= imem02_in[87:84];
    62: reg_0857 <= imem02_in[87:84];
    66: reg_0857 <= imem06_in[3:0];
    68: reg_0857 <= imem00_in[119:116];
    71: reg_0857 <= imem06_in[3:0];
    89: reg_0857 <= imem04_in[87:84];
    91: reg_0857 <= imem00_in[3:0];
    endcase
  end

  // REG#858の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0858 <= imem06_in[7:4];
    8: reg_0858 <= imem06_in[7:4];
    10: reg_0858 <= imem06_in[23:20];
    12: reg_0858 <= imem07_in[103:100];
    14: reg_0858 <= imem07_in[103:100];
    16: reg_0858 <= imem01_in[15:12];
    18: reg_0858 <= imem06_in[7:4];
    20: reg_0858 <= imem07_in[103:100];
    21: reg_0858 <= op2_02_out;
    60: reg_0858 <= op2_02_out;
    endcase
  end

  // REG#859の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0859 <= imem06_in[15:12];
    8: reg_0859 <= imem06_in[15:12];
    11: reg_0859 <= imem03_in[23:20];
    14: reg_0859 <= imem06_in[15:12];
    16: reg_0859 <= imem03_in[23:20];
    18: reg_0859 <= imem03_in[23:20];
    19: reg_0859 <= op2_02_out;
    53: reg_0859 <= op2_02_out;
    81: reg_0859 <= op2_02_out;
    88: reg_0859 <= imem03_in[23:20];
    endcase
  end

  // REG#860の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0860 <= imem06_in[71:68];
    8: reg_0860 <= imem06_in[71:68];
    10: reg_0860 <= imem06_in[55:52];
    12: reg_0860 <= imem07_in[127:124];
    14: reg_0860 <= imem07_in[127:124];
    16: reg_0860 <= imem06_in[55:52];
    19: reg_0860 <= imem07_in[127:124];
    21: reg_0860 <= imem06_in[71:68];
    23: reg_0860 <= imem01_in[71:68];
    25: reg_0860 <= imem01_in[71:68];
    47: reg_0860 <= imem01_in[71:68];
    51: reg_0860 <= imem07_in[127:124];
    53: reg_0860 <= imem01_in[71:68];
    endcase
  end

  // REG#861の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0861 <= imem06_in[75:72];
    8: reg_0861 <= imem04_in[59:56];
    10: reg_0861 <= imem06_in[75:72];
    12: reg_0861 <= imem00_in[19:16];
    14: reg_0861 <= imem03_in[19:16];
    16: reg_0861 <= imem01_in[59:56];
    20: reg_0861 <= imem00_in[19:16];
    21: reg_0861 <= op2_03_out;
    63: reg_0861 <= imem06_in[75:72];
    65: reg_0861 <= imem00_in[19:16];
    67: reg_0861 <= imem04_in[59:56];
    69: reg_0861 <= imem00_in[19:16];
    71: reg_0861 <= imem04_in[59:56];
    73: reg_0861 <= imem06_in[75:72];
    75: reg_0861 <= imem00_in[19:16];
    76: reg_0861 <= op2_03_out;
    endcase
  end

  // REG#862の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0862 <= imem06_in[79:76];
    8: reg_0862 <= imem06_in[79:76];
    10: reg_0862 <= imem07_in[75:72];
    12: reg_0862 <= imem07_in[75:72];
    14: reg_0862 <= imem07_in[75:72];
    16: reg_0862 <= imem01_in[119:116];
    18: reg_0862 <= imem06_in[79:76];
    19: reg_0862 <= op2_03_out;
    55: reg_0862 <= imem06_in[79:76];
    57: reg_0862 <= imem07_in[75:72];
    59: reg_0862 <= imem06_in[79:76];
    61: reg_0862 <= imem07_in[75:72];
    63: reg_0862 <= imem01_in[119:116];
    65: reg_0862 <= imem07_in[75:72];
    67: reg_0862 <= imem07_in[75:72];
    69: reg_0862 <= imem01_in[119:116];
    91: reg_0862 <= imem07_in[75:72];
    93: reg_0862 <= op2_03_out;
    endcase
  end

  // REG#863の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0863 <= imem06_in[87:84];
    8: reg_0863 <= imem05_in[3:0];
    10: reg_0863 <= imem06_in[87:84];
    12: reg_0863 <= imem05_in[3:0];
    20: reg_0863 <= imem06_in[87:84];
    22: reg_0863 <= imem05_in[3:0];
    24: reg_0863 <= imem06_in[87:84];
    26: reg_0863 <= imem02_in[23:20];
    55: reg_0863 <= imem05_in[3:0];
    58: reg_0863 <= imem06_in[87:84];
    85: reg_0863 <= imem05_in[3:0];
    88: reg_0863 <= imem05_in[3:0];
    91: reg_0863 <= imem06_in[87:84];
    94: reg_0863 <= imem05_in[3:0];
    endcase
  end

  // REG#864の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0864 <= imem06_in[127:124];
    8: reg_0864 <= imem06_in[127:124];
    11: reg_0864 <= imem04_in[99:96];
    14: reg_0864 <= imem04_in[99:96];
    16: reg_0864 <= imem04_in[99:96];
    18: reg_0864 <= imem04_in[99:96];
    46: reg_0864 <= imem04_in[99:96];
    49: reg_0864 <= imem04_in[99:96];
    60: reg_0864 <= imem06_in[127:124];
    63: reg_0864 <= imem04_in[99:96];
    69: reg_0864 <= imem00_in[71:68];
    71: reg_0864 <= imem00_in[71:68];
    73: reg_0864 <= imem00_in[71:68];
    75: reg_0864 <= imem00_in[71:68];
    77: reg_0864 <= imem04_in[99:96];
    79: reg_0864 <= imem00_in[71:68];
    81: reg_0864 <= imem00_in[71:68];
    83: reg_0864 <= imem04_in[99:96];
    endcase
  end

  // REG#865の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0865 <= imem07_in[47:44];
    8: reg_0865 <= imem05_in[83:80];
    10: reg_0865 <= imem05_in[83:80];
    12: reg_0865 <= imem05_in[83:80];
    21: reg_0865 <= imem07_in[47:44];
    23: reg_0865 <= imem03_in[67:64];
    26: reg_0865 <= imem02_in[79:76];
    54: reg_0865 <= imem03_in[67:64];
    58: reg_0865 <= imem07_in[47:44];
    60: reg_0865 <= imem07_in[47:44];
    63: reg_0865 <= imem02_in[79:76];
    66: reg_0865 <= imem05_in[83:80];
    79: reg_0865 <= imem06_in[51:48];
    81: reg_0865 <= imem05_in[83:80];
    83: reg_0865 <= imem06_in[51:48];
    85: reg_0865 <= imem06_in[51:48];
    88: reg_0865 <= imem06_in[51:48];
    91: reg_0865 <= imem03_in[67:64];
    93: reg_0865 <= imem03_in[67:64];
    endcase
  end

  // REG#866の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0866 <= imem07_in[123:120];
    8: reg_0866 <= imem07_in[67:64];
    10: reg_0866 <= imem00_in[59:56];
    12: reg_0866 <= imem07_in[123:120];
    14: reg_0866 <= imem07_in[123:120];
    16: reg_0866 <= imem00_in[59:56];
    18: reg_0866 <= imem00_in[59:56];
    21: reg_0866 <= imem00_in[59:56];
    23: reg_0866 <= imem00_in[59:56];
    25: reg_0866 <= imem07_in[67:64];
    27: reg_0866 <= imem07_in[123:120];
    29: reg_0866 <= imem07_in[67:64];
    31: reg_0866 <= imem07_in[67:64];
    34: reg_0866 <= imem05_in[15:12];
    36: reg_0866 <= imem07_in[67:64];
    38: reg_0866 <= imem05_in[15:12];
    40: reg_0866 <= imem00_in[59:56];
    42: reg_0866 <= imem07_in[67:64];
    45: reg_0866 <= imem07_in[123:120];
    47: reg_0866 <= imem07_in[123:120];
    49: reg_0866 <= imem07_in[67:64];
    53: reg_0866 <= imem00_in[59:56];
    56: reg_0866 <= imem05_in[15:12];
    63: reg_0866 <= imem05_in[15:12];
    65: reg_0866 <= imem00_in[59:56];
    67: reg_0866 <= imem00_in[59:56];
    69: reg_0866 <= imem00_in[59:56];
    71: reg_0866 <= imem00_in[59:56];
    73: reg_0866 <= imem05_in[15:12];
    endcase
  end

  // REG#867の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0867 <= imem00_in[43:40];
    8: reg_0867 <= imem07_in[95:92];
    10: reg_0867 <= imem07_in[95:92];
    12: reg_0867 <= imem00_in[43:40];
    14: reg_0867 <= imem03_in[123:120];
    16: reg_0867 <= imem03_in[123:120];
    21: reg_0867 <= imem02_in[35:32];
    86: reg_0867 <= imem07_in[95:92];
    91: reg_0867 <= imem00_in[43:40];
    endcase
  end

  // REG#868の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0868 <= imem00_in[127:124];
    8: reg_0868 <= imem07_in[111:108];
    10: reg_0868 <= imem00_in[63:60];
    12: reg_0868 <= imem00_in[67:64];
    14: reg_0868 <= imem07_in[111:108];
    16: reg_0868 <= imem00_in[63:60];
    18: reg_0868 <= imem00_in[127:124];
    20: reg_0868 <= imem00_in[127:124];
    22: reg_0868 <= imem00_in[127:124];
    24: reg_0868 <= imem07_in[111:108];
    26: reg_0868 <= imem00_in[127:124];
    28: reg_0868 <= imem00_in[127:124];
    30: reg_0868 <= imem00_in[127:124];
    33: reg_0868 <= imem07_in[111:108];
    35: reg_0868 <= imem00_in[127:124];
    37: reg_0868 <= imem00_in[67:64];
    39: reg_0868 <= imem00_in[67:64];
    41: reg_0868 <= imem00_in[67:64];
    43: reg_0868 <= imem07_in[111:108];
    endcase
  end

  // REG#869の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0869 <= imem01_in[27:24];
    8: reg_0869 <= imem01_in[27:24];
    10: reg_0869 <= imem01_in[27:24];
    41: reg_0869 <= imem01_in[27:24];
    95: reg_0869 <= imem01_in[27:24];
    endcase
  end

  // REG#870の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0870 <= imem01_in[59:56];
    8: reg_0870 <= imem00_in[23:20];
    10: reg_0870 <= imem00_in[23:20];
    12: reg_0870 <= imem00_in[23:20];
    14: reg_0870 <= imem04_in[47:44];
    16: reg_0870 <= imem00_in[23:20];
    18: reg_0870 <= imem00_in[23:20];
    20: reg_0870 <= imem04_in[47:44];
    23: reg_0870 <= imem04_in[71:68];
    25: reg_0870 <= imem04_in[71:68];
    28: reg_0870 <= imem04_in[71:68];
    31: reg_0870 <= imem00_in[23:20];
    33: reg_0870 <= imem04_in[71:68];
    35: reg_0870 <= imem04_in[71:68];
    39: reg_0870 <= imem01_in[59:56];
    44: reg_0870 <= imem01_in[59:56];
    47: reg_0870 <= imem00_in[23:20];
    49: reg_0870 <= imem01_in[59:56];
    71: reg_0870 <= imem00_in[23:20];
    73: reg_0870 <= imem00_in[23:20];
    75: reg_0870 <= imem01_in[59:56];
    77: reg_0870 <= imem04_in[47:44];
    79: reg_0870 <= imem04_in[71:68];
    81: reg_0870 <= imem04_in[47:44];
    83: reg_0870 <= imem04_in[47:44];
    endcase
  end

  // REG#871の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0871 <= imem01_in[103:100];
    8: reg_0871 <= imem00_in[95:92];
    10: reg_0871 <= imem01_in[103:100];
    40: reg_0871 <= imem01_in[103:100];
    42: reg_0871 <= imem01_in[103:100];
    47: reg_0871 <= imem01_in[103:100];
    49: reg_0871 <= imem01_in[103:100];
    66: reg_0871 <= imem01_in[103:100];
    68: reg_0871 <= imem00_in[95:92];
    70: reg_0871 <= imem01_in[103:100];
    72: reg_0871 <= imem00_in[95:92];
    79: reg_0871 <= imem00_in[95:92];
    89: reg_0871 <= imem01_in[103:100];
    91: reg_0871 <= imem00_in[95:92];
    endcase
  end

  // REG#872の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0872 <= imem02_in[7:4];
    8: reg_0872 <= imem02_in[7:4];
    10: reg_0872 <= imem02_in[7:4];
    12: reg_0872 <= imem00_in[95:92];
    14: reg_0872 <= imem00_in[95:92];
    16: reg_0872 <= imem02_in[111:108];
    18: reg_0872 <= imem00_in[95:92];
    21: reg_0872 <= imem02_in[111:108];
    86: reg_0872 <= imem02_in[7:4];
    89: reg_0872 <= imem00_in[95:92];
    93: reg_0872 <= imem02_in[111:108];
    95: reg_0872 <= imem02_in[111:108];
    endcase
  end

  // REG#873の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0873 <= imem04_in[3:0];
    8: reg_0873 <= imem04_in[3:0];
    10: reg_0873 <= imem00_in[71:68];
    12: reg_0873 <= imem02_in[59:56];
    14: reg_0873 <= imem04_in[63:60];
    16: reg_0873 <= imem04_in[63:60];
    19: reg_0873 <= imem00_in[71:68];
    21: reg_0873 <= imem00_in[71:68];
    23: reg_0873 <= imem04_in[63:60];
    25: reg_0873 <= imem00_in[71:68];
    27: reg_0873 <= imem00_in[71:68];
    29: reg_0873 <= imem04_in[63:60];
    31: reg_0873 <= imem04_in[63:60];
    33: reg_0873 <= op1_12_out;
    36: reg_0873 <= imem04_in[63:60];
    39: reg_0873 <= imem00_in[71:68];
    41: reg_0873 <= imem02_in[59:56];
    42: reg_0873 <= op1_12_out;
    46: reg_0873 <= imem04_in[63:60];
    50: reg_0873 <= imem00_in[71:68];
    51: reg_0873 <= op1_12_out;
    54: reg_0873 <= imem04_in[3:0];
    55: reg_0873 <= op1_12_out;
    58: reg_0873 <= imem04_in[3:0];
    61: reg_0873 <= imem00_in[71:68];
    63: reg_0873 <= imem02_in[59:56];
    71: reg_0873 <= imem02_in[59:56];
    74: reg_0873 <= imem04_in[3:0];
    75: reg_0873 <= op1_12_out;
    78: reg_0873 <= imem02_in[59:56];
    83: reg_0873 <= imem00_in[71:68];
    85: reg_0873 <= imem00_in[71:68];
    87: reg_0873 <= op1_12_out;
    89: reg_0873 <= op1_12_out;
    92: reg_0873 <= op1_12_out;
    95: reg_0873 <= imem04_in[3:0];
    endcase
  end

  // REG#874の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0874 <= imem04_in[23:20];
    8: reg_0874 <= imem04_in[23:20];
    10: reg_0874 <= imem00_in[87:84];
    12: reg_0874 <= imem03_in[3:0];
    14: reg_0874 <= imem05_in[119:116];
    16: reg_0874 <= imem05_in[119:116];
    18: reg_0874 <= imem05_in[119:116];
    20: reg_0874 <= imem00_in[87:84];
    22: reg_0874 <= imem05_in[119:116];
    24: reg_0874 <= imem05_in[119:116];
    26: reg_0874 <= imem04_in[23:20];
    28: reg_0874 <= imem03_in[11:8];
    72: reg_0874 <= imem03_in[3:0];
    74: reg_0874 <= imem00_in[87:84];
    76: reg_0874 <= imem05_in[119:116];
    78: reg_0874 <= imem03_in[11:8];
    80: reg_0874 <= imem03_in[11:8];
    82: reg_0874 <= imem05_in[119:116];
    85: reg_0874 <= imem03_in[11:8];
    87: reg_0874 <= imem03_in[3:0];
    90: reg_0874 <= imem03_in[11:8];
    94: reg_0874 <= imem03_in[11:8];
    endcase
  end

  // REG#875の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0875 <= imem04_in[71:68];
    8: reg_0875 <= imem01_in[47:44];
    10: reg_0875 <= imem04_in[71:68];
    12: reg_0875 <= imem03_in[35:32];
    14: reg_0875 <= imem06_in[31:28];
    16: reg_0875 <= imem03_in[35:32];
    18: reg_0875 <= imem04_in[71:68];
    43: reg_0875 <= imem01_in[47:44];
    45: reg_0875 <= imem06_in[31:28];
    48: reg_0875 <= imem04_in[71:68];
    51: reg_0875 <= imem06_in[31:28];
    53: reg_0875 <= imem06_in[31:28];
    56: reg_0875 <= imem04_in[71:68];
    58: reg_0875 <= imem03_in[35:32];
    60: reg_0875 <= imem04_in[71:68];
    62: reg_0875 <= imem04_in[71:68];
    64: reg_0875 <= imem04_in[71:68];
    66: reg_0875 <= imem06_in[31:28];
    68: reg_0875 <= imem06_in[31:28];
    71: reg_0875 <= imem01_in[47:44];
    73: reg_0875 <= imem01_in[47:44];
    75: reg_0875 <= imem04_in[71:68];
    79: reg_0875 <= imem01_in[47:44];
    81: reg_0875 <= imem04_in[71:68];
    84: reg_0875 <= imem04_in[71:68];
    86: reg_0875 <= imem04_in[71:68];
    88: reg_0875 <= imem04_in[71:68];
    90: reg_0875 <= imem01_in[47:44];
    92: reg_0875 <= imem04_in[71:68];
    94: reg_0875 <= imem01_in[47:44];
    endcase
  end

  // REG#876の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0876 <= imem06_in[47:44];
    8: reg_0876 <= imem06_in[47:44];
    11: reg_0876 <= imem05_in[43:40];
    13: reg_0876 <= imem06_in[47:44];
    15: reg_0876 <= imem06_in[47:44];
    17: reg_0876 <= imem04_in[111:108];
    21: reg_0876 <= imem02_in[43:40];
    86: reg_0876 <= imem05_in[43:40];
    88: reg_0876 <= imem06_in[47:44];
    endcase
  end

  // REG#877の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0877 <= imem06_in[67:64];
    8: reg_0877 <= imem01_in[91:88];
    10: reg_0877 <= imem06_in[67:64];
    12: reg_0877 <= imem06_in[67:64];
    14: reg_0877 <= imem06_in[67:64];
    16: reg_0877 <= imem01_in[91:88];
    19: reg_0877 <= imem01_in[91:88];
    21: reg_0877 <= imem01_in[91:88];
    23: reg_0877 <= imem04_in[51:48];
    28: reg_0877 <= imem04_in[51:48];
    31: reg_0877 <= imem04_in[51:48];
    33: reg_0877 <= imem04_in[51:48];
    35: reg_0877 <= imem01_in[91:88];
    38: reg_0877 <= imem06_in[67:64];
    41: reg_0877 <= imem04_in[51:48];
    43: reg_0877 <= imem06_in[67:64];
    45: reg_0877 <= imem04_in[51:48];
    48: reg_0877 <= imem04_in[51:48];
    51: reg_0877 <= imem06_in[67:64];
    53: reg_0877 <= imem01_in[91:88];
    95: reg_0877 <= imem01_in[91:88];
    endcase
  end

  // REG#878の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0878 <= imem06_in[95:92];
    8: reg_0878 <= imem06_in[95:92];
    11: reg_0878 <= imem05_in[59:56];
    14: reg_0878 <= imem05_in[59:56];
    15: reg_0878 <= op2_01_out;
    39: reg_0878 <= op2_01_out;
    77: reg_0878 <= op2_01_out;
    endcase
  end

  // REG#879の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0879 <= imem07_in[11:8];
    8: reg_0879 <= imem02_in[11:8];
    10: reg_0879 <= imem07_in[11:8];
    12: reg_0879 <= imem04_in[63:60];
    14: reg_0879 <= imem07_in[11:8];
    15: reg_0879 <= op2_02_out;
    40: reg_0879 <= op2_02_out;
    83: reg_0879 <= imem02_in[11:8];
    86: reg_0879 <= imem04_in[63:60];
    90: reg_0879 <= imem02_in[11:8];
    92: reg_0879 <= imem07_in[11:8];
    95: reg_0879 <= op2_02_out;
    endcase
  end

  // REG#880の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0880 <= imem07_in[15:12];
    8: reg_0880 <= imem07_in[15:12];
    10: reg_0880 <= imem02_in[31:28];
    12: reg_0880 <= imem07_in[15:12];
    14: reg_0880 <= imem07_in[15:12];
    16: reg_0880 <= imem02_in[31:28];
    21: reg_0880 <= imem07_in[15:12];
    23: reg_0880 <= imem02_in[31:28];
    27: reg_0880 <= imem02_in[31:28];
    31: reg_0880 <= imem02_in[59:56];
    33: reg_0880 <= op2_01_out;
    57: reg_0880 <= op2_01_out;
    93: reg_0880 <= op2_01_out;
    endcase
  end

  // REG#881の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0881 <= imem07_in[71:68];
    8: reg_0881 <= imem02_in[83:80];
    10: reg_0881 <= imem07_in[71:68];
    12: reg_0881 <= imem04_in[83:80];
    14: reg_0881 <= imem02_in[83:80];
    17: reg_0881 <= imem07_in[71:68];
    20: reg_0881 <= imem02_in[83:80];
    22: reg_0881 <= op2_02_out;
    64: reg_0881 <= op2_02_out;
    75: reg_0881 <= imem02_in[83:80];
    76: reg_0881 <= op2_02_out;
    endcase
  end

  // REG#882の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0882 <= imem00_in[55:52];
    8: reg_0882 <= imem03_in[19:16];
    10: reg_0882 <= imem00_in[55:52];
    12: reg_0882 <= imem04_in[111:108];
    14: reg_0882 <= imem00_in[55:52];
    16: reg_0882 <= imem00_in[55:52];
    19: reg_0882 <= imem04_in[111:108];
    42: reg_0882 <= imem00_in[55:52];
    46: reg_0882 <= imem04_in[111:108];
    49: reg_0882 <= imem04_in[111:108];
    60: reg_0882 <= imem03_in[19:16];
    63: reg_0882 <= imem00_in[55:52];
    66: reg_0882 <= imem00_in[55:52];
    68: reg_0882 <= imem04_in[111:108];
    71: reg_0882 <= imem04_in[111:108];
    75: reg_0882 <= imem04_in[111:108];
    78: reg_0882 <= imem04_in[111:108];
    81: reg_0882 <= imem04_in[111:108];
    83: reg_0882 <= imem04_in[111:108];
    endcase
  end

  // REG#883の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0883 <= imem00_in[75:72];
    8: reg_0883 <= imem03_in[23:20];
    10: reg_0883 <= imem03_in[23:20];
    12: reg_0883 <= imem00_in[75:72];
    14: reg_0883 <= imem03_in[23:20];
    17: reg_0883 <= imem00_in[75:72];
    19: reg_0883 <= imem00_in[75:72];
    21: reg_0883 <= imem03_in[23:20];
    23: reg_0883 <= imem03_in[23:20];
    26: reg_0883 <= imem00_in[75:72];
    29: reg_0883 <= imem00_in[75:72];
    31: reg_0883 <= imem00_in[75:72];
    33: reg_0883 <= imem00_in[75:72];
    36: reg_0883 <= imem03_in[23:20];
    39: reg_0883 <= imem06_in[19:16];
    55: reg_0883 <= imem00_in[75:72];
    91: reg_0883 <= imem06_in[19:16];
    93: reg_0883 <= imem03_in[23:20];
    endcase
  end

  // REG#884の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0884 <= imem00_in[123:120];
    8: reg_0884 <= imem03_in[51:48];
    10: reg_0884 <= imem03_in[51:48];
    12: reg_0884 <= imem04_in[119:116];
    14: reg_0884 <= imem07_in[71:68];
    16: reg_0884 <= imem03_in[51:48];
    18: reg_0884 <= imem07_in[71:68];
    21: reg_0884 <= imem02_in[107:104];
    86: reg_0884 <= imem02_in[107:104];
    90: reg_0884 <= imem04_in[119:116];
    92: reg_0884 <= imem04_in[119:116];
    94: reg_0884 <= imem07_in[71:68];
    endcase
  end

  // REG#885の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0885 <= imem01_in[35:32];
    8: reg_0885 <= imem01_in[35:32];
    10: reg_0885 <= imem01_in[35:32];
    42: reg_0885 <= imem01_in[35:32];
    44: reg_0885 <= imem01_in[35:32];
    47: reg_0885 <= imem01_in[35:32];
    57: reg_0885 <= imem01_in[35:32];
    60: reg_0885 <= imem01_in[35:32];
    62: reg_0885 <= imem01_in[35:32];
    68: reg_0885 <= imem01_in[35:32];
    72: reg_0885 <= imem02_in[63:60];
    85: reg_0885 <= imem02_in[63:60];
    endcase
  end

  // REG#886の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0886 <= imem02_in[67:64];
    8: reg_0886 <= imem03_in[63:60];
    10: reg_0886 <= imem02_in[67:64];
    12: reg_0886 <= imem03_in[63:60];
    14: reg_0886 <= imem03_in[63:60];
    17: reg_0886 <= imem03_in[63:60];
    19: reg_0886 <= imem03_in[63:60];
    21: reg_0886 <= imem03_in[63:60];
    24: reg_0886 <= imem06_in[19:16];
    26: reg_0886 <= imem02_in[67:64];
    53: reg_0886 <= imem02_in[67:64];
    55: reg_0886 <= imem06_in[19:16];
    57: reg_0886 <= imem02_in[67:64];
    59: reg_0886 <= imem06_in[19:16];
    61: reg_0886 <= imem03_in[63:60];
    63: reg_0886 <= imem03_in[63:60];
    68: reg_0886 <= imem06_in[19:16];
    70: reg_0886 <= imem06_in[19:16];
    72: reg_0886 <= imem02_in[79:76];
    85: reg_0886 <= imem02_in[67:64];
    endcase
  end

  // REG#887の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0887 <= imem02_in[91:88];
    8: reg_0887 <= imem02_in[91:88];
    10: reg_0887 <= imem02_in[95:92];
    12: reg_0887 <= imem02_in[95:92];
    14: reg_0887 <= imem07_in[115:112];
    16: reg_0887 <= imem02_in[91:88];
    18: reg_0887 <= imem02_in[95:92];
    20: reg_0887 <= imem02_in[95:92];
    23: reg_0887 <= imem02_in[91:88];
    25: reg_0887 <= imem07_in[115:112];
    27: reg_0887 <= imem07_in[115:112];
    30: reg_0887 <= imem02_in[95:92];
    32: reg_0887 <= imem07_in[115:112];
    33: reg_0887 <= op2_03_out;
    61: reg_0887 <= imem02_in[91:88];
    63: reg_0887 <= imem02_in[91:88];
    72: reg_0887 <= imem02_in[95:92];
    84: reg_0887 <= imem02_in[91:88];
    endcase
  end

  // REG#888の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0888 <= imem02_in[99:96];
    8: reg_0888 <= imem04_in[95:92];
    10: reg_0888 <= imem03_in[3:0];
    12: reg_0888 <= imem02_in[99:96];
    14: reg_0888 <= imem04_in[95:92];
    16: reg_0888 <= imem04_in[95:92];
    18: reg_0888 <= imem02_in[99:96];
    20: reg_0888 <= imem03_in[3:0];
    22: reg_0888 <= imem03_in[3:0];
    24: reg_0888 <= imem04_in[95:92];
    83: reg_0888 <= imem04_in[95:92];
    endcase
  end

  // REG#889の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0889 <= imem02_in[119:116];
    8: reg_0889 <= imem02_in[119:116];
    10: reg_0889 <= imem02_in[119:116];
    12: reg_0889 <= imem02_in[119:116];
    13: reg_0889 <= op1_13_out;
    16: reg_0889 <= op1_13_out;
    18: reg_0889 <= op1_13_out;
    20: reg_0889 <= op1_13_out;
    22: reg_0889 <= op1_13_out;
    24: reg_0889 <= op1_13_out;
    27: reg_0889 <= imem02_in[119:116];
    28: reg_0889 <= op1_13_out;
    33: reg_0889 <= op1_13_out;
    36: reg_0889 <= imem02_in[119:116];
    39: reg_0889 <= imem06_in[119:116];
    57: reg_0889 <= imem06_in[119:116];
    endcase
  end

  // REG#890の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0890 <= imem04_in[27:24];
    8: reg_0890 <= imem04_in[119:116];
    10: reg_0890 <= imem03_in[79:76];
    12: reg_0890 <= imem04_in[27:24];
    13: reg_0890 <= op2_00_out;
    32: reg_0890 <= imem04_in[119:116];
    34: reg_0890 <= imem04_in[27:24];
    37: reg_0890 <= imem03_in[79:76];
    38: reg_0890 <= op2_00_out;
    73: reg_0890 <= imem04_in[27:24];
    74: reg_0890 <= op2_00_out;
    endcase
  end

  // REG#891の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0891 <= imem04_in[43:40];
    8: reg_0891 <= imem05_in[39:36];
    10: reg_0891 <= imem04_in[59:56];
    12: reg_0891 <= imem05_in[59:56];
    13: reg_0891 <= op2_01_out;
    32: reg_0891 <= op2_01_out;
    55: reg_0891 <= imem04_in[59:56];
    56: reg_0891 <= op2_01_out;
    90: reg_0891 <= imem04_in[43:40];
    92: reg_0891 <= imem05_in[59:56];
    95: reg_0891 <= imem04_in[43:40];
    endcase
  end

  // REG#892の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0892 <= imem04_in[79:76];
    8: reg_0892 <= imem04_in[79:76];
    10: reg_0892 <= imem04_in[79:76];
    12: reg_0892 <= imem07_in[23:20];
    14: reg_0892 <= imem07_in[23:20];
    17: reg_0892 <= imem04_in[79:76];
    22: reg_0892 <= imem04_in[79:76];
    26: reg_0892 <= imem04_in[79:76];
    29: reg_0892 <= imem07_in[23:20];
    31: reg_0892 <= imem05_in[67:64];
    33: reg_0892 <= imem05_in[67:64];
    35: reg_0892 <= imem05_in[67:64];
    37: reg_0892 <= imem05_in[67:64];
    39: reg_0892 <= imem06_in[63:60];
    58: reg_0892 <= imem04_in[79:76];
    60: reg_0892 <= imem04_in[79:76];
    62: reg_0892 <= imem07_in[23:20];
    64: reg_0892 <= imem05_in[67:64];
    68: reg_0892 <= imem07_in[23:20];
    70: reg_0892 <= imem04_in[79:76];
    72: reg_0892 <= imem05_in[67:64];
    75: reg_0892 <= imem07_in[23:20];
    79: reg_0892 <= imem05_in[67:64];
    87: reg_0892 <= imem05_in[67:64];
    endcase
  end

  // REG#893の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0893 <= imem04_in[127:124];
    8: reg_0893 <= imem04_in[127:124];
    10: reg_0893 <= imem05_in[123:120];
    12: reg_0893 <= imem04_in[127:124];
    13: reg_0893 <= op2_03_out;
    38: reg_0893 <= imem04_in[127:124];
    40: reg_0893 <= imem05_in[123:120];
    42: reg_0893 <= imem04_in[127:124];
    endcase
  end

  // REG#894の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0894 <= imem06_in[19:16];
    8: reg_0894 <= imem06_in[19:16];
    10: reg_0894 <= imem05_in[127:124];
    12: reg_0894 <= imem05_in[127:124];
    19: reg_0894 <= imem05_in[127:124];
    23: reg_0894 <= imem05_in[127:124];
    25: reg_0894 <= imem05_in[127:124];
    31: reg_0894 <= imem06_in[19:16];
    37: reg_0894 <= imem06_in[19:16];
    61: reg_0894 <= imem03_in[67:64];
    63: reg_0894 <= imem02_in[99:96];
    73: reg_0894 <= imem06_in[19:16];
    75: reg_0894 <= imem05_in[127:124];
    77: reg_0894 <= imem03_in[67:64];
    79: reg_0894 <= imem02_in[103:100];
    83: reg_0894 <= imem06_in[19:16];
    85: reg_0894 <= imem02_in[99:96];
    endcase
  end

  // REG#895の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0895 <= imem07_in[51:48];
    8: reg_0895 <= imem07_in[51:48];
    10: reg_0895 <= imem07_in[51:48];
    12: reg_0895 <= imem07_in[55:52];
    14: reg_0895 <= imem07_in[51:48];
    17: reg_0895 <= imem07_in[55:52];
    19: reg_0895 <= imem07_in[55:52];
    22: reg_0895 <= imem07_in[55:52];
    24: reg_0895 <= imem07_in[127:124];
    26: reg_0895 <= imem07_in[55:52];
    28: reg_0895 <= imem07_in[127:124];
    30: reg_0895 <= imem07_in[51:48];
    32: reg_0895 <= imem07_in[51:48];
    36: reg_0895 <= imem07_in[127:124];
    39: reg_0895 <= imem06_in[27:24];
    58: reg_0895 <= imem06_in[27:24];
    86: reg_0895 <= imem06_in[27:24];
    endcase
  end

  // REG#896の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0896 <= imem07_in[115:112];
    8: reg_0896 <= imem05_in[79:76];
    10: reg_0896 <= imem00_in[47:44];
    12: reg_0896 <= imem05_in[107:104];
    16: reg_0896 <= imem00_in[47:44];
    18: reg_0896 <= imem00_in[47:44];
    20: reg_0896 <= imem05_in[107:104];
    51: reg_0896 <= imem07_in[115:112];
    55: reg_0896 <= imem05_in[107:104];
    57: reg_0896 <= imem07_in[115:112];
    59: reg_0896 <= imem05_in[107:104];
    61: reg_0896 <= imem07_in[115:112];
    63: reg_0896 <= imem05_in[79:76];
    65: reg_0896 <= imem05_in[107:104];
    69: reg_0896 <= imem05_in[107:104];
    72: reg_0896 <= imem02_in[39:36];
    86: reg_0896 <= imem07_in[115:112];
    89: reg_0896 <= imem02_in[39:36];
    91: reg_0896 <= imem07_in[115:112];
    93: reg_0896 <= imem05_in[107:104];
    endcase
  end

  // REG#897の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0897 <= imem00_in[31:28];
    8: reg_0897 <= imem06_in[111:108];
    10: reg_0897 <= imem00_in[31:28];
    12: reg_0897 <= imem05_in[91:88];
    16: reg_0897 <= imem00_in[31:28];
    18: reg_0897 <= imem00_in[31:28];
    21: reg_0897 <= imem05_in[91:88];
    24: reg_0897 <= imem00_in[83:80];
    26: reg_0897 <= imem05_in[91:88];
    28: reg_0897 <= imem05_in[91:88];
    30: reg_0897 <= imem05_in[91:88];
    32: reg_0897 <= imem00_in[31:28];
    34: reg_0897 <= imem00_in[83:80];
    36: reg_0897 <= imem06_in[111:108];
    40: reg_0897 <= imem00_in[83:80];
    47: reg_0897 <= imem00_in[83:80];
    49: reg_0897 <= imem05_in[91:88];
    51: reg_0897 <= imem06_in[111:108];
    54: reg_0897 <= imem00_in[83:80];
    57: reg_0897 <= imem00_in[83:80];
    59: reg_0897 <= imem06_in[111:108];
    61: reg_0897 <= imem06_in[111:108];
    72: reg_0897 <= imem00_in[83:80];
    74: reg_0897 <= imem00_in[31:28];
    78: reg_0897 <= imem06_in[111:108];
    80: reg_0897 <= imem06_in[111:108];
    82: reg_0897 <= imem06_in[111:108];
    84: reg_0897 <= imem05_in[91:88];
    86: reg_0897 <= imem00_in[31:28];
    88: reg_0897 <= imem00_in[31:28];
    90: reg_0897 <= imem05_in[91:88];
    92: reg_0897 <= imem06_in[111:108];
    endcase
  end

  // REG#898の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0898 <= imem00_in[35:32];
    8: reg_0898 <= imem00_in[35:32];
    10: reg_0898 <= imem00_in[35:32];
    12: reg_0898 <= imem05_in[95:92];
    19: reg_0898 <= imem00_in[35:32];
    23: reg_0898 <= imem00_in[35:32];
    26: reg_0898 <= imem00_in[35:32];
    28: reg_0898 <= imem05_in[95:92];
    30: reg_0898 <= imem05_in[95:92];
    32: reg_0898 <= imem05_in[95:92];
    34: reg_0898 <= imem05_in[95:92];
    36: reg_0898 <= imem05_in[95:92];
    38: reg_0898 <= op2_01_out;
    73: reg_0898 <= op2_01_out;
    endcase
  end

  // REG#899の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0899 <= imem00_in[47:44];
    8: reg_0899 <= imem07_in[7:4];
    10: reg_0899 <= imem07_in[7:4];
    12: reg_0899 <= imem07_in[7:4];
    17: reg_0899 <= imem04_in[31:28];
    21: reg_0899 <= imem07_in[7:4];
    23: reg_0899 <= imem07_in[7:4];
    26: reg_0899 <= imem00_in[47:44];
    28: reg_0899 <= imem04_in[31:28];
    31: reg_0899 <= imem07_in[7:4];
    34: reg_0899 <= imem00_in[47:44];
    39: reg_0899 <= imem00_in[47:44];
    41: reg_0899 <= imem00_in[47:44];
    47: reg_0899 <= imem07_in[7:4];
    49: reg_0899 <= imem04_in[31:28];
    61: reg_0899 <= imem03_in[75:72];
    63: reg_0899 <= imem02_in[39:36];
    73: reg_0899 <= imem07_in[7:4];
    75: reg_0899 <= imem03_in[75:72];
    77: reg_0899 <= imem00_in[47:44];
    79: reg_0899 <= imem00_in[47:44];
    81: reg_0899 <= imem00_in[47:44];
    83: reg_0899 <= imem00_in[47:44];
    89: reg_0899 <= imem07_in[7:4];
    91: reg_0899 <= imem00_in[47:44];
    endcase
  end

  // REG#900の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0900 <= imem00_in[51:48];
    8: reg_0900 <= imem00_in[51:48];
    10: reg_0900 <= imem00_in[51:48];
    12: reg_0900 <= imem05_in[31:28];
    20: reg_0900 <= imem05_in[31:28];
    51: reg_0900 <= imem00_in[51:48];
    53: reg_0900 <= imem05_in[31:28];
    55: reg_0900 <= imem00_in[51:48];
    89: reg_0900 <= imem00_in[51:48];
    92: reg_0900 <= imem00_in[51:48];
    94: reg_0900 <= imem05_in[31:28];
    endcase
  end

  // REG#901の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0901 <= imem00_in[99:96];
    8: reg_0901 <= imem07_in[55:52];
    10: reg_0901 <= imem07_in[55:52];
    12: reg_0901 <= imem00_in[99:96];
    16: reg_0901 <= op2_00_out;
    42: reg_0901 <= op2_00_out;
    45: reg_0901 <= imem07_in[55:52];
    46: reg_0901 <= op2_00_out;
    58: reg_0901 <= imem00_in[99:96];
    59: reg_0901 <= op2_00_out;
    endcase
  end

  // REG#902の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0902 <= imem01_in[75:72];
    8: reg_0902 <= imem07_in[83:80];
    10: reg_0902 <= imem07_in[83:80];
    12: reg_0902 <= imem05_in[99:96];
    21: reg_0902 <= imem01_in[75:72];
    24: reg_0902 <= imem01_in[15:12];
    27: reg_0902 <= imem05_in[99:96];
    29: reg_0902 <= imem05_in[99:96];
    31: reg_0902 <= imem05_in[99:96];
    34: reg_0902 <= imem07_in[83:80];
    36: reg_0902 <= imem01_in[75:72];
    38: reg_0902 <= imem01_in[15:12];
    41: reg_0902 <= imem01_in[75:72];
    90: reg_0902 <= imem07_in[83:80];
    92: reg_0902 <= imem01_in[15:12];
    endcase
  end

  // REG#903の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0903 <= imem01_in[87:84];
    8: reg_0903 <= imem07_in[119:116];
    10: reg_0903 <= imem07_in[119:116];
    12: reg_0903 <= imem05_in[23:20];
    21: reg_0903 <= imem07_in[119:116];
    23: reg_0903 <= op2_03_out;
    25: reg_0903 <= op2_03_out;
    34: reg_0903 <= imem01_in[87:84];
    36: reg_0903 <= imem05_in[23:20];
    38: reg_0903 <= op2_03_out;
    77: reg_0903 <= imem01_in[87:84];
    79: reg_0903 <= imem07_in[119:116];
    endcase
  end

  // REG#904の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0904 <= imem01_in[123:120];
    8: reg_0904 <= imem00_in[67:64];
    10: reg_0904 <= imem01_in[123:120];
    40: reg_0904 <= imem00_in[67:64];
    44: reg_0904 <= imem00_in[67:64];
    47: reg_0904 <= imem00_in[67:64];
    49: reg_0904 <= imem01_in[47:44];
    63: reg_0904 <= imem00_in[67:64];
    67: reg_0904 <= imem00_in[67:64];
    69: reg_0904 <= imem01_in[123:120];
    94: reg_0904 <= imem01_in[123:120];
    96: reg_0904 <= imem01_in[47:44];
    endcase
  end

  // REG#905の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0905 <= imem01_in[127:124];
    8: reg_0905 <= imem01_in[3:0];
    10: reg_0905 <= imem01_in[3:0];
    37: reg_0905 <= imem01_in[127:124];
    39: reg_0905 <= imem01_in[3:0];
    43: reg_0905 <= imem01_in[127:124];
    45: reg_0905 <= imem01_in[127:124];
    47: reg_0905 <= imem01_in[127:124];
    52: reg_0905 <= imem01_in[127:124];
    61: reg_0905 <= imem04_in[59:56];
    63: reg_0905 <= imem02_in[23:20];
    73: reg_0905 <= imem04_in[59:56];
    75: reg_0905 <= imem04_in[59:56];
    77: reg_0905 <= imem02_in[23:20];
    79: reg_0905 <= imem04_in[59:56];
    81: reg_0905 <= imem04_in[59:56];
    84: reg_0905 <= imem04_in[59:56];
    86: reg_0905 <= imem02_in[23:20];
    88: reg_0905 <= imem04_in[59:56];
    91: reg_0905 <= imem02_in[23:20];
    93: reg_0905 <= imem01_in[3:0];
    endcase
  end

  // REG#906の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0906 <= imem02_in[39:36];
    8: reg_0906 <= imem01_in[39:36];
    10: reg_0906 <= imem02_in[39:36];
    12: reg_0906 <= imem01_in[39:36];
    14: reg_0906 <= imem02_in[39:36];
    16: reg_0906 <= imem01_in[39:36];
    20: reg_0906 <= imem01_in[39:36];
    22: reg_0906 <= imem01_in[39:36];
    24: reg_0906 <= imem01_in[123:120];
    27: reg_0906 <= imem01_in[39:36];
    29: reg_0906 <= imem01_in[39:36];
    31: reg_0906 <= imem01_in[39:36];
    34: reg_0906 <= imem01_in[39:36];
    36: reg_0906 <= imem02_in[39:36];
    38: reg_0906 <= imem02_in[39:36];
    41: reg_0906 <= imem01_in[123:120];
    94: reg_0906 <= imem02_in[39:36];
    endcase
  end

  // REG#907の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0907 <= imem02_in[71:68];
    8: reg_0907 <= imem02_in[71:68];
    9: reg_0907 <= op1_13_out;
    12: reg_0907 <= imem02_in[71:68];
    14: reg_0907 <= imem02_in[71:68];
    15: reg_0907 <= op1_13_out;
    18: reg_0907 <= imem02_in[71:68];
    19: reg_0907 <= op1_13_out;
    23: reg_0907 <= op1_13_out;
    25: reg_0907 <= op1_13_out;
    27: reg_0907 <= op1_13_out;
    30: reg_0907 <= op1_13_out;
    42: reg_0907 <= imem02_in[71:68];
    44: reg_0907 <= imem02_in[71:68];
    48: reg_0907 <= imem02_in[71:68];
    50: reg_0907 <= op1_13_out;
    56: reg_0907 <= imem02_in[71:68];
    58: reg_0907 <= imem02_in[71:68];
    59: reg_0907 <= op1_13_out;
    62: reg_0907 <= op1_13_out;
    65: reg_0907 <= op1_13_out;
    68: reg_0907 <= op1_13_out;
    72: reg_0907 <= imem02_in[71:68];
    82: reg_0907 <= op1_13_out;
    86: reg_0907 <= imem02_in[71:68];
    88: reg_0907 <= imem02_in[71:68];
    90: reg_0907 <= op1_13_out;
    endcase
  end

  // REG#908の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0908 <= imem02_in[111:108];
    8: reg_0908 <= imem02_in[111:108];
    10: reg_0908 <= imem02_in[111:108];
    12: reg_0908 <= imem05_in[47:44];
    23: reg_0908 <= imem02_in[111:108];
    25: reg_0908 <= imem05_in[47:44];
    29: reg_0908 <= imem02_in[111:108];
    31: reg_0908 <= imem02_in[111:108];
    34: reg_0908 <= imem05_in[47:44];
    37: reg_0908 <= imem02_in[111:108];
    39: reg_0908 <= imem05_in[47:44];
    43: reg_0908 <= imem05_in[47:44];
    49: reg_0908 <= imem05_in[47:44];
    51: reg_0908 <= imem05_in[47:44];
    54: reg_0908 <= imem02_in[111:108];
    56: reg_0908 <= imem05_in[47:44];
    59: reg_0908 <= imem02_in[111:108];
    61: reg_0908 <= imem02_in[111:108];
    63: reg_0908 <= imem02_in[111:108];
    72: reg_0908 <= imem02_in[111:108];
    87: reg_0908 <= imem02_in[111:108];
    89: reg_0908 <= imem02_in[111:108];
    94: reg_0908 <= imem02_in[111:108];
    endcase
  end

  // REG#909の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0909 <= imem04_in[7:4];
    8: reg_0909 <= imem04_in[7:4];
    9: reg_0909 <= op1_14_out;
    12: reg_0909 <= op1_14_out;
    14: reg_0909 <= op1_14_out;
    16: reg_0909 <= op1_14_out;
    19: reg_0909 <= op1_14_out;
    22: reg_0909 <= op1_14_out;
    24: reg_0909 <= op1_14_out;
    26: reg_0909 <= op1_14_out;
    28: reg_0909 <= op1_14_out;
    31: reg_0909 <= op1_14_out;
    34: reg_0909 <= op1_14_out;
    42: reg_0909 <= imem04_in[7:4];
    endcase
  end

  // REG#910の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0910 <= imem04_in[11:8];
    8: reg_0910 <= imem04_in[11:8];
    10: reg_0910 <= imem04_in[11:8];
    11: reg_0910 <= op2_01_out;
    26: reg_0910 <= op2_01_out;
    34: reg_0910 <= op2_01_out;
    62: reg_0910 <= op2_01_out;
    67: reg_0910 <= op2_01_out;
    82: reg_0910 <= op2_01_out;
    90: reg_0910 <= op2_01_out;
    endcase
  end

  // REG#911の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0911 <= imem04_in[15:12];
    8: reg_0911 <= imem04_in[15:12];
    10: reg_0911 <= imem04_in[15:12];
    11: reg_0911 <= op2_02_out;
    27: reg_0911 <= op2_02_out;
    38: reg_0911 <= op2_02_out;
    74: reg_0911 <= op2_02_out;
    endcase
  end

  // REG#912の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0912 <= imem04_in[55:52];
    8: reg_0912 <= imem04_in[55:52];
    10: reg_0912 <= imem04_in[55:52];
    12: reg_0912 <= imem04_in[55:52];
    15: reg_0912 <= imem04_in[55:52];
    17: reg_0912 <= imem04_in[55:52];
    21: reg_0912 <= imem04_in[55:52];
    24: reg_0912 <= imem04_in[55:52];
    83: reg_0912 <= imem04_in[55:52];
    endcase
  end

  // REG#913の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0913 <= imem04_in[75:72];
    8: reg_0913 <= imem01_in[83:80];
    10: reg_0913 <= imem01_in[83:80];
    40: reg_0913 <= imem01_in[83:80];
    43: reg_0913 <= imem01_in[83:80];
    45: reg_0913 <= imem01_in[83:80];
    48: reg_0913 <= imem01_in[83:80];
    50: reg_0913 <= imem01_in[83:80];
    52: reg_0913 <= imem01_in[83:80];
    56: reg_0913 <= imem01_in[83:80];
    61: reg_0913 <= imem04_in[111:108];
    63: reg_0913 <= imem01_in[83:80];
    66: reg_0913 <= imem01_in[83:80];
    68: reg_0913 <= imem01_in[83:80];
    70: reg_0913 <= imem04_in[75:72];
    72: reg_0913 <= imem04_in[111:108];
    74: reg_0913 <= imem04_in[75:72];
    78: reg_0913 <= imem04_in[75:72];
    81: reg_0913 <= imem04_in[75:72];
    83: reg_0913 <= imem04_in[75:72];
    endcase
  end

  // REG#914の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0914 <= imem06_in[35:32];
    8: reg_0914 <= imem06_in[35:32];
    10: reg_0914 <= op1_02_out;
    16: reg_0914 <= imem06_in[35:32];
    18: reg_0914 <= imem06_in[35:32];
    21: reg_0914 <= imem06_in[35:32];
    23: reg_0914 <= imem06_in[35:32];
    25: reg_0914 <= imem06_in[35:32];
    29: reg_0914 <= imem06_in[35:32];
    61: reg_0914 <= imem07_in[79:76];
    63: reg_0914 <= imem02_in[63:60];
    73: reg_0914 <= imem07_in[79:76];
    79: reg_0914 <= imem02_in[63:60];
    83: reg_0914 <= imem02_in[63:60];
    87: reg_0914 <= imem06_in[35:32];
    89: reg_0914 <= imem06_in[35:32];
    endcase
  end

  // REG#915の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0915 <= imem06_in[63:60];
    8: reg_0915 <= imem06_in[63:60];
    10: reg_0915 <= imem06_in[63:60];
    12: reg_0915 <= imem06_in[63:60];
    17: reg_0915 <= imem06_in[63:60];
    19: reg_0915 <= imem06_in[63:60];
    24: reg_0915 <= imem06_in[63:60];
    28: reg_0915 <= imem06_in[63:60];
    31: reg_0915 <= imem06_in[23:20];
    33: reg_0915 <= imem06_in[63:60];
    35: reg_0915 <= imem06_in[63:60];
    39: reg_0915 <= imem06_in[23:20];
    56: reg_0915 <= imem06_in[23:20];
    61: reg_0915 <= imem06_in[23:20];
    71: reg_0915 <= imem06_in[63:60];
    90: reg_0915 <= imem06_in[63:60];
    92: reg_0915 <= imem06_in[23:20];
    endcase
  end

  // REG#916の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0916 <= imem06_in[83:80];
    8: reg_0916 <= imem02_in[15:12];
    10: reg_0916 <= imem02_in[15:12];
    16: reg_0916 <= imem02_in[15:12];
    18: reg_0916 <= imem06_in[83:80];
    20: reg_0916 <= imem06_in[83:80];
    22: reg_0916 <= imem02_in[15:12];
    24: reg_0916 <= imem02_in[15:12];
    26: reg_0916 <= imem02_in[15:12];
    51: reg_0916 <= imem02_in[15:12];
    55: reg_0916 <= imem06_in[83:80];
    61: reg_0916 <= imem06_in[83:80];
    69: reg_0916 <= imem00_in[123:120];
    72: reg_0916 <= imem02_in[15:12];
    84: reg_0916 <= imem02_in[15:12];
    endcase
  end

  // REG#917の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0917 <= imem06_in[119:116];
    8: reg_0917 <= imem02_in[43:40];
    9: reg_0917 <= op1_15_out;
    12: reg_0917 <= op1_15_out;
    14: reg_0917 <= op1_15_out;
    16: reg_0917 <= op1_15_out;
    20: reg_0917 <= imem02_in[43:40];
    22: reg_0917 <= op1_15_out;
    25: reg_0917 <= op1_15_out;
    29: reg_0917 <= imem06_in[119:116];
    58: reg_0917 <= imem06_in[119:116];
    88: reg_0917 <= op1_15_out;
    endcase
  end

  // REG#918の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0918 <= imem06_in[123:120];
    8: reg_0918 <= imem02_in[47:44];
    10: reg_0918 <= imem02_in[47:44];
    14: reg_0918 <= imem02_in[47:44];
    17: reg_0918 <= imem02_in[47:44];
    20: reg_0918 <= imem02_in[47:44];
    24: reg_0918 <= imem01_in[23:20];
    28: reg_0918 <= imem02_in[47:44];
    30: reg_0918 <= imem02_in[47:44];
    32: reg_0918 <= imem02_in[47:44];
    37: reg_0918 <= imem02_in[47:44];
    40: reg_0918 <= imem02_in[47:44];
    42: reg_0918 <= imem06_in[123:120];
    44: reg_0918 <= imem02_in[47:44];
    46: reg_0918 <= imem01_in[23:20];
    49: reg_0918 <= imem01_in[3:0];
    65: reg_0918 <= imem01_in[23:20];
    68: reg_0918 <= imem01_in[3:0];
    72: reg_0918 <= imem01_in[3:0];
    74: reg_0918 <= imem01_in[3:0];
    76: reg_0918 <= imem06_in[123:120];
    78: reg_0918 <= imem01_in[3:0];
    81: reg_0918 <= imem01_in[3:0];
    83: reg_0918 <= imem01_in[23:20];
    86: reg_0918 <= imem06_in[123:120];
    endcase
  end

  // REG#919の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0919 <= imem07_in[3:0];
    8: reg_0919 <= imem07_in[3:0];
    10: reg_0919 <= imem07_in[3:0];
    13: reg_0919 <= imem07_in[3:0];
    16: reg_0919 <= imem07_in[3:0];
    18: reg_0919 <= imem07_in[3:0];
    23: reg_0919 <= imem07_in[3:0];
    26: reg_0919 <= imem07_in[3:0];
    28: reg_0919 <= imem07_in[3:0];
    31: reg_0919 <= imem06_in[47:44];
    34: reg_0919 <= imem07_in[3:0];
    37: reg_0919 <= imem07_in[3:0];
    40: reg_0919 <= imem07_in[3:0];
    45: reg_0919 <= imem06_in[47:44];
    49: reg_0919 <= imem01_in[63:60];
    68: reg_0919 <= imem06_in[47:44];
    70: reg_0919 <= imem01_in[63:60];
    72: reg_0919 <= imem01_in[63:60];
    75: reg_0919 <= imem07_in[3:0];
    81: reg_0919 <= imem06_in[47:44];
    83: reg_0919 <= imem01_in[63:60];
    85: reg_0919 <= imem06_in[47:44];
    87: reg_0919 <= imem07_in[3:0];
    89: reg_0919 <= imem06_in[47:44];
    endcase
  end

  // REG#920の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0920 <= imem07_in[23:20];
    8: reg_0920 <= imem02_in[75:72];
    10: reg_0920 <= imem02_in[75:72];
    12: reg_0920 <= imem02_in[75:72];
    14: reg_0920 <= imem02_in[75:72];
    16: reg_0920 <= op2_02_out;
    44: reg_0920 <= op2_02_out;
    52: reg_0920 <= op2_02_out;
    78: reg_0920 <= op2_02_out;
    endcase
  end

  // REG#921の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0921 <= imem07_in[39:36];
    8: reg_0921 <= imem07_in[39:36];
    10: reg_0921 <= imem07_in[39:36];
    16: reg_0921 <= imem07_in[39:36];
    20: reg_0921 <= imem07_in[39:36];
    22: reg_0921 <= imem07_in[39:36];
    24: reg_0921 <= imem07_in[39:36];
    26: reg_0921 <= imem07_in[39:36];
    28: reg_0921 <= imem07_in[39:36];
    31: reg_0921 <= imem06_in[15:12];
    34: reg_0921 <= imem06_in[15:12];
    38: reg_0921 <= imem07_in[39:36];
    43: reg_0921 <= imem06_in[15:12];
    46: reg_0921 <= imem07_in[39:36];
    49: reg_0921 <= imem07_in[39:36];
    51: reg_0921 <= imem06_in[15:12];
    54: reg_0921 <= imem06_in[15:12];
    57: reg_0921 <= imem07_in[39:36];
    60: reg_0921 <= imem07_in[39:36];
    62: reg_0921 <= imem07_in[39:36];
    65: reg_0921 <= imem06_in[15:12];
    67: reg_0921 <= imem06_in[15:12];
    69: reg_0921 <= imem06_in[15:12];
    71: reg_0921 <= imem06_in[15:12];
    91: reg_0921 <= imem06_in[15:12];
    94: reg_0921 <= imem07_in[39:36];
    96: reg_0921 <= imem06_in[15:12];
    endcase
  end

  // REG#922の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0922 <= imem07_in[63:60];
    8: reg_0922 <= imem07_in[63:60];
    9: reg_0922 <= op2_00_out;
    19: reg_0922 <= imem07_in[63:60];
    21: reg_0922 <= imem07_in[63:60];
    22: reg_0922 <= op2_00_out;
    62: reg_0922 <= op2_00_out;
    67: reg_0922 <= op2_00_out;
    81: reg_0922 <= op2_00_out;
    89: reg_0922 <= op2_00_out;
    endcase
  end

  // REG#923の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0923 <= imem07_in[79:76];
    8: reg_0923 <= imem03_in[15:12];
    10: reg_0923 <= imem03_in[15:12];
    14: reg_0923 <= imem03_in[15:12];
    18: reg_0923 <= imem07_in[79:76];
    20: reg_0923 <= imem03_in[15:12];
    24: reg_0923 <= imem07_in[79:76];
    26: reg_0923 <= imem03_in[15:12];
    28: reg_0923 <= imem03_in[15:12];
    71: reg_0923 <= imem07_in[79:76];
    79: reg_0923 <= imem07_in[79:76];
    endcase
  end

  // REG#924の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0924 <= imem07_in[91:88];
    8: reg_0924 <= imem07_in[91:88];
    9: reg_0924 <= op2_02_out;
    20: reg_0924 <= op2_02_out;
    57: reg_0924 <= op2_02_out;
    endcase
  end

  // REG#925の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0925 <= imem07_in[107:104];
    8: reg_0925 <= imem03_in[75:72];
    10: reg_0925 <= imem03_in[75:72];
    12: reg_0925 <= imem07_in[107:104];
    14: reg_0925 <= imem07_in[107:104];
    16: reg_0925 <= imem07_in[107:104];
    18: reg_0925 <= imem07_in[107:104];
    20: reg_0925 <= imem07_in[107:104];
    22: reg_0925 <= imem07_in[107:104];
    24: reg_0925 <= imem01_in[119:116];
    27: reg_0925 <= imem03_in[75:72];
    31: reg_0925 <= imem06_in[79:76];
    34: reg_0925 <= imem06_in[79:76];
    36: reg_0925 <= imem06_in[79:76];
    41: reg_0925 <= imem01_in[119:116];
    95: reg_0925 <= imem01_in[119:116];
    endcase
  end

  // REG#926の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0926 <= op1_00_out;
    8: reg_0926 <= imem03_in[87:84];
    10: reg_0926 <= imem03_in[87:84];
    12: reg_0926 <= imem03_in[87:84];
    17: reg_0926 <= imem03_in[87:84];
    21: reg_0926 <= imem03_in[87:84];
    24: reg_0926 <= imem01_in[67:64];
    27: reg_0926 <= imem01_in[67:64];
    29: reg_0926 <= imem01_in[67:64];
    31: reg_0926 <= imem06_in[99:96];
    34: reg_0926 <= imem01_in[67:64];
    37: reg_0926 <= imem06_in[99:96];
    57: reg_0926 <= imem06_in[99:96];
    endcase
  end

  // REG#927の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0927 <= op1_01_out;
    7: reg_0927 <= op1_01_out;
    9: reg_0927 <= op1_01_out;
    22: reg_0927 <= op1_01_out;
    26: reg_0927 <= op1_01_out;
    28: reg_0927 <= op1_01_out;
    30: reg_0927 <= op1_01_out;
    32: reg_0927 <= op1_01_out;
    34: reg_0927 <= op1_01_out;
    36: reg_0927 <= op1_01_out;
    38: reg_0927 <= op1_01_out;
    40: reg_0927 <= op1_01_out;
    42: reg_0927 <= op1_01_out;
    44: reg_0927 <= op1_01_out;
    46: reg_0927 <= op1_01_out;
    48: reg_0927 <= op1_01_out;
    50: reg_0927 <= op1_01_out;
    52: reg_0927 <= op1_01_out;
    54: reg_0927 <= op1_01_out;
    56: reg_0927 <= op1_01_out;
    58: reg_0927 <= op1_01_out;
    60: reg_0927 <= op1_01_out;
    64: reg_0927 <= op1_01_out;
    66: reg_0927 <= op1_01_out;
    68: reg_0927 <= op1_01_out;
    76: reg_0927 <= op1_01_out;
    78: reg_0927 <= op1_01_out;
    80: reg_0927 <= op1_01_out;
    82: reg_0927 <= op1_01_out;
    84: reg_0927 <= op1_01_out;
    86: reg_0927 <= op1_01_out;
    88: reg_0927 <= op1_01_out;
    90: reg_0927 <= op1_01_out;
    94: reg_0927 <= op1_01_out;
    endcase
  end

  // REG#928の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0928 <= op1_02_out;
    7: reg_0928 <= op1_02_out;
    9: reg_0928 <= op1_02_out;
    24: reg_0928 <= imem01_in[83:80];
    28: reg_0928 <= imem01_in[83:80];
    31: reg_0928 <= imem06_in[75:72];
    35: reg_0928 <= imem06_in[75:72];
    38: reg_0928 <= imem06_in[75:72];
    41: reg_0928 <= imem06_in[75:72];
    45: reg_0928 <= imem06_in[75:72];
    47: reg_0928 <= imem06_in[75:72];
    49: reg_0928 <= imem01_in[27:24];
    70: reg_0928 <= imem01_in[27:24];
    72: reg_0928 <= imem06_in[75:72];
    77: reg_0928 <= imem01_in[27:24];
    79: reg_0928 <= imem01_in[27:24];
    81: reg_0928 <= imem06_in[75:72];
    83: reg_0928 <= imem01_in[27:24];
    86: reg_0928 <= imem06_in[75:72];
    endcase
  end

  // REG#929の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0929 <= op1_03_out;
    7: reg_0929 <= op1_03_out;
    9: reg_0929 <= op1_03_out;
    11: reg_0929 <= op1_03_out;
    23: reg_0929 <= op2_00_out;
    65: reg_0929 <= op1_03_out;
    68: reg_0929 <= op2_00_out;
    84: reg_0929 <= op2_00_out;
    95: reg_0929 <= op2_00_out;
    endcase
  end

  // REG#930の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0930 <= op1_04_out;
    7: reg_0930 <= op1_04_out;
    9: reg_0930 <= op1_04_out;
    11: reg_0930 <= op1_04_out;
    16: reg_0930 <= op1_04_out;
    18: reg_0930 <= op1_04_out;
    23: reg_0930 <= op2_01_out;
    68: reg_0930 <= op2_01_out;
    85: reg_0930 <= op2_01_out;
    endcase
  end

  // REG#931の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0931 <= op1_05_out;
    7: reg_0931 <= op1_05_out;
    9: reg_0931 <= op1_05_out;
    11: reg_0931 <= op1_05_out;
    13: reg_0931 <= op1_05_out;
    15: reg_0931 <= op1_05_out;
    17: reg_0931 <= op1_05_out;
    19: reg_0931 <= op1_05_out;
    24: reg_0931 <= imem04_in[107:104];
    82: reg_0931 <= imem04_in[107:104];
    93: reg_0931 <= imem04_in[107:104];
    endcase
  end

  // REG#932の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0932 <= op1_06_out;
    7: reg_0932 <= op1_06_out;
    9: reg_0932 <= op1_06_out;
    11: reg_0932 <= op1_06_out;
    13: reg_0932 <= op1_06_out;
    16: reg_0932 <= op1_06_out;
    24: reg_0932 <= imem04_in[111:108];
    82: reg_0932 <= imem04_in[111:108];
    endcase
  end

  // REG#933の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0933 <= op1_07_out;
    7: reg_0933 <= op1_07_out;
    9: reg_0933 <= op1_07_out;
    11: reg_0933 <= op1_07_out;
    13: reg_0933 <= op1_07_out;
    15: reg_0933 <= op1_07_out;
    17: reg_0933 <= op1_07_out;
    19: reg_0933 <= op1_07_out;
    21: reg_0933 <= op1_07_out;
    23: reg_0933 <= op1_07_out;
    31: reg_0933 <= imem03_in[83:80];
    47: reg_0933 <= imem03_in[83:80];
    49: reg_0933 <= imem01_in[55:52];
    72: reg_0933 <= imem03_in[83:80];
    74: reg_0933 <= imem03_in[83:80];
    77: reg_0933 <= imem01_in[55:52];
    79: reg_0933 <= imem03_in[83:80];
    81: reg_0933 <= imem01_in[55:52];
    83: reg_0933 <= imem01_in[55:52];
    91: reg_0933 <= imem01_in[55:52];
    93: reg_0933 <= imem01_in[55:52];
    endcase
  end

  // REG#934の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0934 <= op1_08_out;
    7: reg_0934 <= op1_08_out;
    9: reg_0934 <= op1_08_out;
    11: reg_0934 <= op1_08_out;
    13: reg_0934 <= op1_08_out;
    15: reg_0934 <= op1_08_out;
    17: reg_0934 <= op1_08_out;
    19: reg_0934 <= op1_08_out;
    21: reg_0934 <= op1_08_out;
    23: reg_0934 <= op1_08_out;
    30: reg_0934 <= op2_00_out;
    47: reg_0934 <= op2_00_out;
    60: reg_0934 <= op2_00_out;
    endcase
  end

  // REG#935の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0935 <= op1_09_out;
    7: reg_0935 <= op1_09_out;
    9: reg_0935 <= op1_09_out;
    11: reg_0935 <= op1_09_out;
    13: reg_0935 <= op1_09_out;
    15: reg_0935 <= op1_09_out;
    17: reg_0935 <= op1_09_out;
    20: reg_0935 <= op1_09_out;
    22: reg_0935 <= op1_09_out;
    24: reg_0935 <= op1_09_out;
    26: reg_0935 <= op1_09_out;
    28: reg_0935 <= op1_09_out;
    30: reg_0935 <= op1_09_out;
    32: reg_0935 <= op1_09_out;
    34: reg_0935 <= op1_09_out;
    36: reg_0935 <= op1_09_out;
    38: reg_0935 <= op1_09_out;
    40: reg_0935 <= op1_09_out;
    42: reg_0935 <= op1_09_out;
    44: reg_0935 <= op1_09_out;
    48: reg_0935 <= op1_09_out;
    50: reg_0935 <= op1_09_out;
    52: reg_0935 <= op1_09_out;
    54: reg_0935 <= op1_09_out;
    56: reg_0935 <= op1_09_out;
    61: reg_0935 <= imem05_in[31:28];
    66: reg_0935 <= imem05_in[31:28];
    84: reg_0935 <= imem05_in[31:28];
    87: reg_0935 <= imem05_in[31:28];
    endcase
  end

  // REG#936の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0936 <= op1_10_out;
    7: reg_0936 <= op1_10_out;
    9: reg_0936 <= op1_10_out;
    11: reg_0936 <= op1_10_out;
    13: reg_0936 <= op1_10_out;
    15: reg_0936 <= op1_10_out;
    17: reg_0936 <= op1_10_out;
    19: reg_0936 <= op1_10_out;
    21: reg_0936 <= op1_10_out;
    23: reg_0936 <= op1_10_out;
    25: reg_0936 <= op1_10_out;
    30: reg_0936 <= op2_02_out;
    49: reg_0936 <= imem01_in[31:28];
    69: reg_0936 <= op2_02_out;
    89: reg_0936 <= op2_02_out;
    endcase
  end

  // REG#937の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0937 <= op1_11_out;
    7: reg_0937 <= op1_11_out;
    9: reg_0937 <= op1_11_out;
    11: reg_0937 <= op1_11_out;
    13: reg_0937 <= op1_11_out;
    15: reg_0937 <= op1_11_out;
    17: reg_0937 <= op1_11_out;
    19: reg_0937 <= op1_11_out;
    21: reg_0937 <= op1_11_out;
    24: reg_0937 <= imem04_in[39:36];
    83: reg_0937 <= imem04_in[39:36];
    endcase
  end

  // REG#938の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0938 <= op1_12_out;
    7: reg_0938 <= op1_12_out;
    9: reg_0938 <= op1_12_out;
    11: reg_0938 <= op1_12_out;
    13: reg_0938 <= op1_12_out;
    15: reg_0938 <= op1_12_out;
    17: reg_0938 <= op1_12_out;
    19: reg_0938 <= op1_12_out;
    21: reg_0938 <= op1_12_out;
    24: reg_0938 <= op1_12_out;
    26: reg_0938 <= op1_12_out;
    31: reg_0938 <= imem03_in[47:44];
    51: reg_0938 <= imem03_in[47:44];
    53: reg_0938 <= op1_12_out;
    57: reg_0938 <= imem03_in[47:44];
    58: reg_0938 <= op1_12_out;
    60: reg_0938 <= op1_12_out;
    64: reg_0938 <= op1_12_out;
    66: reg_0938 <= op1_12_out;
    70: reg_0938 <= op1_12_out;
    75: reg_0938 <= imem03_in[47:44];
    77: reg_0938 <= op1_12_out;
    82: reg_0938 <= op1_12_out;
    90: reg_0938 <= imem03_in[47:44];
    endcase
  end

  // REG#939の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0939 <= op1_13_out;
    7: reg_0939 <= op1_13_out;
    10: reg_0939 <= op1_13_out;
    12: reg_0939 <= op1_13_out;
    14: reg_0939 <= op1_13_out;
    17: reg_0939 <= op1_13_out;
    21: reg_0939 <= op1_13_out;
    26: reg_0939 <= op1_13_out;
    30: reg_0939 <= op2_03_out;
    60: reg_0939 <= op2_03_out;
    endcase
  end

  // REG#940の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0940 <= op1_14_out;
    8: reg_0940 <= op1_14_out;
    11: reg_0940 <= op1_14_out;
    15: reg_0940 <= op1_14_out;
    17: reg_0940 <= op1_14_out;
    20: reg_0940 <= op1_14_out;
    23: reg_0940 <= op1_14_out;
    27: reg_0940 <= op1_14_out;
    31: reg_0940 <= imem03_in[11:8];
    53: reg_0940 <= imem03_in[11:8];
    57: reg_0940 <= imem03_in[11:8];
    61: reg_0940 <= imem05_in[19:16];
    66: reg_0940 <= imem05_in[19:16];
    79: reg_0940 <= op1_14_out;
    82: reg_0940 <= op1_14_out;
    86: reg_0940 <= imem05_in[19:16];
    89: reg_0940 <= imem05_in[19:16];
    91: reg_0940 <= imem05_in[19:16];
    93: reg_0940 <= op1_14_out;
    endcase
  end

  // REG#941の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0941 <= op1_15_out;
    8: reg_0941 <= op1_15_out;
    11: reg_0941 <= op1_15_out;
    15: reg_0941 <= op1_15_out;
    17: reg_0941 <= op1_15_out;
    20: reg_0941 <= op1_15_out;
    23: reg_0941 <= op1_15_out;
    26: reg_0941 <= op1_15_out;
    28: reg_0941 <= op1_15_out;
    31: reg_0941 <= op1_15_out;
    35: reg_0941 <= op1_15_out;
    49: reg_0941 <= op1_15_out;
    53: reg_0941 <= op1_15_out;
    61: reg_0941 <= imem05_in[15:12];
    66: reg_0941 <= imem05_in[15:12];
    79: reg_0941 <= op1_15_out;
    82: reg_0941 <= op1_15_out;
    endcase
  end

  // REG#942の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0942 <= imem05_in[79:76];
    55: reg_0942 <= imem05_in[79:76];
    61: reg_0942 <= imem05_in[79:76];
    67: reg_0942 <= imem05_in[79:76];
    75: reg_0942 <= imem05_in[79:76];
    77: reg_0942 <= imem05_in[79:76];
    79: reg_0942 <= imem04_in[11:8];
    81: reg_0942 <= imem04_in[11:8];
    83: reg_0942 <= imem04_in[11:8];
    endcase
  end

  // REG#943の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0943 <= imem05_in[115:112];
    53: reg_0943 <= imem05_in[115:112];
    56: reg_0943 <= imem05_in[115:112];
    67: reg_0943 <= imem05_in[115:112];
    70: reg_0943 <= imem05_in[115:112];
    72: reg_0943 <= imem05_in[115:112];
    79: reg_0943 <= imem05_in[115:112];
    90: reg_0943 <= imem05_in[115:112];
    92: reg_0943 <= imem05_in[115:112];
    endcase
  end

  // REG#944の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0944 <= imem05_in[31:28];
    56: reg_0944 <= imem05_in[31:28];
    62: reg_0944 <= imem05_in[31:28];
    68: reg_0944 <= imem05_in[31:28];
    73: reg_0944 <= imem05_in[31:28];
    endcase
  end

  // REG#945の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0945 <= imem05_in[91:88];
    55: reg_0945 <= imem05_in[91:88];
    59: reg_0945 <= imem05_in[91:88];
    61: reg_0945 <= imem05_in[91:88];
    65: reg_0945 <= imem05_in[91:88];
    68: reg_0945 <= imem05_in[91:88];
    74: reg_0945 <= imem05_in[91:88];
    endcase
  end

  // REG#946の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0946 <= imem05_in[99:96];
    59: reg_0946 <= imem05_in[99:96];
    61: reg_0946 <= imem06_in[11:8];
    72: reg_0946 <= imem05_in[99:96];
    78: reg_0946 <= imem05_in[99:96];
    80: reg_0946 <= imem06_in[11:8];
    82: reg_0946 <= imem06_in[11:8];
    86: reg_0946 <= imem05_in[99:96];
    91: reg_0946 <= imem05_in[99:96];
    96: reg_0946 <= imem06_in[11:8];
    endcase
  end

  // REG#947の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0947 <= imem05_in[111:108];
    54: reg_0947 <= imem05_in[111:108];
    61: reg_0947 <= imem05_in[111:108];
    66: reg_0947 <= imem05_in[111:108];
    79: reg_0947 <= imem05_in[39:36];
    87: reg_0947 <= imem05_in[39:36];
    endcase
  end

  // REG#948の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0948 <= imem05_in[59:56];
    60: reg_0948 <= imem05_in[59:56];
    63: reg_0948 <= imem05_in[59:56];
    66: reg_0948 <= imem05_in[59:56];
    79: reg_0948 <= imem05_in[59:56];
    91: reg_0948 <= imem05_in[59:56];
    95: reg_0948 <= imem05_in[59:56];
    endcase
  end

  // REG#949の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0949 <= imem05_in[83:80];
    55: reg_0949 <= imem05_in[83:80];
    61: reg_0949 <= imem05_in[83:80];
    68: reg_0949 <= imem05_in[83:80];
    74: reg_0949 <= imem05_in[83:80];
    endcase
  end

  // REG#950の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0950 <= imem05_in[67:64];
    56: reg_0950 <= imem05_in[67:64];
    63: reg_0950 <= imem05_in[67:64];
    65: reg_0950 <= imem05_in[67:64];
    68: reg_0950 <= imem05_in[67:64];
    74: reg_0950 <= imem05_in[67:64];
    endcase
  end

  // REG#951の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0951 <= imem05_in[75:72];
    56: reg_0951 <= imem05_in[75:72];
    62: reg_0951 <= imem05_in[75:72];
    64: reg_0951 <= imem05_in[75:72];
    68: reg_0951 <= imem05_in[75:72];
    74: reg_0951 <= imem05_in[75:72];
    endcase
  end

  // REG#952の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0952 <= imem05_in[103:100];
    56: reg_0952 <= imem05_in[103:100];
    68: reg_0952 <= imem05_in[103:100];
    72: reg_0952 <= imem05_in[103:100];
    75: reg_0952 <= imem05_in[103:100];
    79: reg_0952 <= imem05_in[103:100];
    90: reg_0952 <= imem05_in[103:100];
    endcase
  end

  // REG#953の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0953 <= imem05_in[119:116];
    56: reg_0953 <= imem05_in[119:116];
    64: reg_0953 <= imem05_in[119:116];
    68: reg_0953 <= imem05_in[119:116];
    72: reg_0953 <= imem05_in[119:116];
    79: reg_0953 <= imem05_in[51:48];
    90: reg_0953 <= imem05_in[119:116];
    95: reg_0953 <= imem05_in[119:116];
    endcase
  end

  // REG#954の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0954 <= imem05_in[47:44];
    58: reg_0954 <= imem05_in[47:44];
    60: reg_0954 <= imem05_in[47:44];
    63: reg_0954 <= imem05_in[47:44];
    65: reg_0954 <= imem05_in[47:44];
    69: reg_0954 <= imem02_in[119:116];
    71: reg_0954 <= imem02_in[119:116];
    73: reg_0954 <= imem05_in[47:44];
    endcase
  end

  // REG#955の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0955 <= imem05_in[39:36];
    56: reg_0955 <= imem05_in[39:36];
    61: reg_0955 <= imem06_in[95:92];
    73: reg_0955 <= imem06_in[95:92];
    78: reg_0955 <= imem05_in[39:36];
    82: reg_0955 <= imem06_in[95:92];
    85: reg_0955 <= imem05_in[39:36];
    88: reg_0955 <= imem06_in[95:92];
    endcase
  end

  // REG#956の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0956 <= imem05_in[51:48];
    56: reg_0956 <= imem05_in[51:48];
    61: reg_0956 <= imem05_in[51:48];
    66: reg_0956 <= imem05_in[51:48];
    81: reg_0956 <= imem05_in[51:48];
    84: reg_0956 <= imem05_in[51:48];
    87: reg_0956 <= imem05_in[51:48];
    endcase
  end

  // REG#957の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0957 <= imem05_in[55:52];
    56: reg_0957 <= imem05_in[55:52];
    61: reg_0957 <= imem06_in[99:96];
    75: reg_0957 <= imem06_in[99:96];
    77: reg_0957 <= imem06_in[99:96];
    79: reg_0957 <= imem05_in[107:104];
    89: reg_0957 <= imem05_in[107:104];
    94: reg_0957 <= imem05_in[107:104];
    endcase
  end

  // REG#958の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0958 <= imem05_in[19:16];
    57: reg_0958 <= imem05_in[19:16];
    60: reg_0958 <= imem05_in[19:16];
    62: reg_0958 <= imem05_in[19:16];
    65: reg_0958 <= imem05_in[19:16];
    68: reg_0958 <= op1_09_out;
    72: reg_0958 <= imem05_in[19:16];
    76: reg_0958 <= op1_09_out;
    79: reg_0958 <= imem05_in[19:16];
    87: reg_0958 <= imem05_in[19:16];
    endcase
  end

  // REG#959の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0959 <= imem05_in[35:32];
    68: reg_0959 <= op1_12_out;
    72: reg_0959 <= imem05_in[35:32];
    79: reg_0959 <= imem07_in[87:84];
    endcase
  end

  // REG#960の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0960 <= imem05_in[127:124];
    57: reg_0960 <= imem05_in[127:124];
    66: reg_0960 <= imem05_in[127:124];
    85: reg_0960 <= imem05_in[127:124];
    87: reg_0960 <= imem05_in[127:124];
    endcase
  end

  // REG#961の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0961 <= imem05_in[107:104];
    58: reg_0961 <= imem05_in[107:104];
    60: reg_0961 <= imem05_in[107:104];
    62: reg_0961 <= imem05_in[107:104];
    69: reg_0961 <= imem03_in[27:24];
    73: reg_0961 <= imem03_in[27:24];
    75: reg_0961 <= imem05_in[107:104];
    79: reg_0961 <= imem03_in[27:24];
    82: reg_0961 <= imem03_in[27:24];
    87: reg_0961 <= imem03_in[27:24];
    90: reg_0961 <= imem03_in[27:24];
    endcase
  end

  // REG#962の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0962 <= imem05_in[3:0];
    58: reg_0962 <= imem05_in[3:0];
    60: reg_0962 <= imem05_in[3:0];
    65: reg_0962 <= imem05_in[3:0];
    69: reg_0962 <= imem01_in[107:104];
    94: reg_0962 <= imem01_in[107:104];
    endcase
  end

  // REG#963の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0963 <= imem05_in[7:4];
    63: reg_0963 <= imem05_in[7:4];
    66: reg_0963 <= imem05_in[7:4];
    79: reg_0963 <= imem05_in[7:4];
    88: reg_0963 <= imem05_in[7:4];
    90: reg_0963 <= imem05_in[7:4];
    93: reg_0963 <= imem05_in[7:4];
    endcase
  end

  // REG#964の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0964 <= imem05_in[71:68];
    57: reg_0964 <= imem05_in[71:68];
    60: reg_0964 <= imem05_in[71:68];
    62: reg_0964 <= imem05_in[71:68];
    65: reg_0964 <= imem05_in[71:68];
    69: reg_0964 <= imem05_in[71:68];
    72: reg_0964 <= imem05_in[71:68];
    75: reg_0964 <= imem05_in[71:68];
    77: reg_0964 <= imem05_in[71:68];
    79: reg_0964 <= imem05_in[71:68];
    84: reg_0964 <= imem05_in[71:68];
    87: reg_0964 <= imem05_in[71:68];
    endcase
  end

  // REG#965の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0965 <= imem05_in[95:92];
    67: reg_0965 <= imem05_in[95:92];
    69: reg_0965 <= imem05_in[95:92];
    71: reg_0965 <= imem05_in[95:92];
    74: reg_0965 <= imem05_in[95:92];
    endcase
  end

  // REG#966の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0966 <= imem05_in[23:20];
    60: reg_0966 <= imem05_in[23:20];
    66: reg_0966 <= imem05_in[23:20];
    79: reg_0966 <= imem05_in[23:20];
    86: reg_0966 <= imem05_in[23:20];
    endcase
  end

  // REG#967の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0967 <= imem05_in[43:40];
    59: reg_0967 <= imem05_in[43:40];
    61: reg_0967 <= imem05_in[43:40];
    68: reg_0967 <= imem05_in[43:40];
    77: reg_0967 <= imem05_in[43:40];
    79: reg_0967 <= imem05_in[43:40];
    endcase
  end

  // REG#968の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0968 <= imem05_in[87:84];
    57: reg_0968 <= imem05_in[87:84];
    60: reg_0968 <= imem05_in[87:84];
    65: reg_0968 <= imem05_in[87:84];
    69: reg_0968 <= imem01_in[39:36];
    92: reg_0968 <= imem01_in[39:36];
    endcase
  end

  // REG#969の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0969 <= imem05_in[63:60];
    61: reg_0969 <= imem05_in[63:60];
    65: reg_0969 <= imem05_in[63:60];
    69: reg_0969 <= imem01_in[3:0];
    95: reg_0969 <= imem01_in[3:0];
    endcase
  end

  // REG#970の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0970 <= imem05_in[15:12];
    60: reg_0970 <= imem05_in[15:12];
    65: reg_0970 <= imem05_in[15:12];
    68: reg_0970 <= imem05_in[15:12];
    74: reg_0970 <= imem05_in[15:12];
    endcase
  end

  // REG#971の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0971 <= imem05_in[27:24];
    58: reg_0971 <= imem05_in[27:24];
    62: reg_0971 <= imem05_in[27:24];
    64: reg_0971 <= imem05_in[27:24];
    69: reg_0971 <= imem01_in[55:52];
    endcase
  end

  // REG#972の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0972 <= imem05_in[123:120];
    57: reg_0972 <= imem05_in[123:120];
    59: reg_0972 <= imem05_in[123:120];
    61: reg_0972 <= imem05_in[123:120];
    66: reg_0972 <= imem05_in[123:120];
    79: reg_0972 <= imem05_in[123:120];
    87: reg_0972 <= imem05_in[123:120];
    endcase
  end

  // REG#973の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0973 <= imem05_in[11:8];
    60: reg_0973 <= imem05_in[11:8];
    64: reg_0973 <= imem05_in[11:8];
    69: reg_0973 <= imem01_in[31:28];
    94: reg_0973 <= imem05_in[11:8];
    endcase
  end

  // REG#974の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0974 <= imem03_in[75:72];
    89: reg_0974 <= imem03_in[75:72];
    endcase
  end

  // REG#975の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0975 <= imem03_in[87:84];
    90: reg_0975 <= imem03_in[87:84];
    endcase
  end

  // REG#976の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0976 <= imem03_in[107:104];
    88: reg_0976 <= imem03_in[107:104];
    endcase
  end

  // REG#977の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0977 <= imem03_in[83:80];
    endcase
  end

  // REG#978の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0978 <= imem03_in[63:60];
    90: reg_0978 <= imem03_in[63:60];
    endcase
  end

  // REG#979の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0979 <= imem03_in[35:32];
    90: reg_0979 <= imem03_in[35:32];
    endcase
  end

  // REG#980の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0980 <= imem03_in[59:56];
    93: reg_0980 <= imem03_in[59:56];
    endcase
  end

  // REG#981の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0981 <= imem03_in[79:76];
    90: reg_0981 <= imem03_in[79:76];
    endcase
  end

  // REG#982の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0982 <= imem03_in[19:16];
    90: reg_0982 <= imem03_in[19:16];
    endcase
  end

  // REG#983の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0983 <= imem03_in[103:100];
    89: reg_0983 <= imem03_in[103:100];
    endcase
  end

  // REG#984の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0984 <= imem03_in[39:36];
    89: reg_0984 <= imem03_in[39:36];
    94: reg_0984 <= imem03_in[39:36];
    endcase
  end

  // REG#985の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0985 <= imem03_in[3:0];
    95: reg_0985 <= imem03_in[3:0];
    endcase
  end

  // REG#986の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0986 <= imem03_in[55:52];
    90: reg_0986 <= imem03_in[55:52];
    endcase
  end

  // REG#987の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0987 <= imem03_in[7:4];
    90: reg_0987 <= imem03_in[7:4];
    endcase
  end

  // REG#988の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0988 <= imem03_in[91:88];
    90: reg_0988 <= imem03_in[91:88];
    96: reg_0988 <= imem03_in[91:88];
    endcase
  end

  // REG#989の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0989 <= imem03_in[71:68];
    90: reg_0989 <= imem03_in[71:68];
    endcase
  end

  // REG#990の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0990 <= imem03_in[95:92];
    93: reg_0990 <= imem03_in[95:92];
    endcase
  end

  // REG#991の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0991 <= imem03_in[23:20];
    endcase
  end

  // REG#992の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0992 <= imem03_in[27:24];
    91: reg_0992 <= imem03_in[27:24];
    endcase
  end

  // REG#993の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0993 <= imem03_in[51:48];
    endcase
  end

  // REG#994の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0994 <= imem03_in[115:112];
    endcase
  end

  // REG#995の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0995 <= imem03_in[31:28];
    91: reg_0995 <= imem03_in[31:28];
    93: reg_0995 <= imem03_in[31:28];
    endcase
  end

  // REG#996の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0996 <= imem03_in[43:40];
    endcase
  end

  // REG#997の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0997 <= imem03_in[111:108];
    endcase
  end

  // REG#998の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0998 <= imem03_in[11:8];
    endcase
  end

  // REG#999の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0999 <= imem03_in[67:64];
    94: reg_0999 <= imem03_in[67:64];
    endcase
  end

  // REG#1000の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1000 <= imem03_in[99:96];
    endcase
  end

  // REG#1001の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1001 <= imem03_in[47:44];
    91: reg_1001 <= imem03_in[47:44];
    endcase
  end

  // REG#1002の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1002 <= imem03_in[15:12];
    92: reg_1002 <= imem03_in[15:12];
    endcase
  end

  // REG#1003の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1003 <= op1_07_out;
    8: reg_1003 <= op1_07_out;
    10: reg_1003 <= op1_07_out;
    12: reg_1003 <= op1_07_out;
    14: reg_1003 <= op1_07_out;
    24: reg_1003 <= imem04_in[27:24];
    82: reg_1003 <= imem04_in[27:24];
    94: reg_1003 <= imem04_in[27:24];
    endcase
  end

  // REG#1004の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1004 <= op1_08_out;
    8: reg_1004 <= op1_08_out;
    10: reg_1004 <= op1_08_out;
    12: reg_1004 <= op1_08_out;
    14: reg_1004 <= op1_08_out;
    16: reg_1004 <= op1_08_out;
    24: reg_1004 <= imem04_in[3:0];
    81: reg_1004 <= op1_08_out;
    84: reg_1004 <= imem04_in[3:0];
    89: reg_1004 <= imem04_in[3:0];
    91: reg_1004 <= imem04_in[3:0];
    endcase
  end

  // REG#1005の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1005 <= op1_09_out;
    8: reg_1005 <= op1_09_out;
    10: reg_1005 <= op1_09_out;
    12: reg_1005 <= op1_09_out;
    14: reg_1005 <= op1_09_out;
    16: reg_1005 <= op1_09_out;
    18: reg_1005 <= op1_09_out;
    24: reg_1005 <= imem04_in[83:80];
    83: reg_1005 <= imem04_in[83:80];
    endcase
  end

  // REG#1006の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1006 <= op1_10_out;
    8: reg_1006 <= op1_10_out;
    10: reg_1006 <= op1_10_out;
    12: reg_1006 <= op1_10_out;
    14: reg_1006 <= op1_10_out;
    16: reg_1006 <= op1_10_out;
    18: reg_1006 <= op1_10_out;
    24: reg_1006 <= imem04_in[11:8];
    82: reg_1006 <= op1_10_out;
    84: reg_1006 <= op1_10_out;
    86: reg_1006 <= op1_10_out;
    88: reg_1006 <= op1_10_out;
    90: reg_1006 <= op1_10_out;
    92: reg_1006 <= op1_10_out;
    94: reg_1006 <= op1_10_out;
    endcase
  end

  // REG#1007の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1007 <= op1_11_out;
    8: reg_1007 <= op1_11_out;
    10: reg_1007 <= op1_11_out;
    12: reg_1007 <= op1_11_out;
    14: reg_1007 <= op1_11_out;
    16: reg_1007 <= op1_11_out;
    18: reg_1007 <= op1_11_out;
    20: reg_1007 <= op1_11_out;
    22: reg_1007 <= op1_11_out;
    24: reg_1007 <= op1_11_out;
    26: reg_1007 <= op1_11_out;
    31: reg_1007 <= imem03_in[51:48];
    53: reg_1007 <= imem03_in[51:48];
    55: reg_1007 <= imem03_in[51:48];
    88: reg_1007 <= op1_11_out;
    endcase
  end

  // REG#1008の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1008 <= op1_12_out;
    8: reg_1008 <= op1_12_out;
    12: reg_1008 <= op1_12_out;
    14: reg_1008 <= op1_12_out;
    16: reg_1008 <= op1_12_out;
    18: reg_1008 <= op1_12_out;
    20: reg_1008 <= op1_12_out;
    22: reg_1008 <= op1_12_out;
    25: reg_1008 <= op1_12_out;
    27: reg_1008 <= op1_12_out;
    31: reg_1008 <= imem03_in[55:52];
    54: reg_1008 <= imem03_in[55:52];
    57: reg_1008 <= op1_12_out;
    62: reg_1008 <= op1_12_out;
    68: reg_1008 <= imem03_in[55:52];
    70: reg_1008 <= imem03_in[55:52];
    90: reg_1008 <= op1_12_out;
    endcase
  end

  // REG#1009の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1009 <= op1_13_out;
    8: reg_1009 <= op1_13_out;
    11: reg_1009 <= op1_13_out;
    24: reg_1009 <= imem04_in[43:40];
    83: reg_1009 <= imem04_in[43:40];
    endcase
  end

  // REG#1010の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1010 <= op1_14_out;
    9: reg_1010 <= imem06_in[79:76];
    32: reg_1010 <= imem06_in[79:76];
    37: reg_1010 <= imem06_in[79:76];
    61: reg_1010 <= imem06_in[79:76];
    71: reg_1010 <= imem06_in[79:76];
    88: reg_1010 <= op1_14_out;
    endcase
  end

  // REG#1011の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1011 <= op1_15_out;
    9: reg_1011 <= imem06_in[95:92];
    33: reg_1011 <= imem06_in[95:92];
    36: reg_1011 <= imem06_in[95:92];
    41: reg_1011 <= imem06_in[95:92];
    43: reg_1011 <= imem06_in[95:92];
    47: reg_1011 <= imem06_in[95:92];
    57: reg_1011 <= imem06_in[95:92];
    endcase
  end

  // REG#1012の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1012 <= op2_00_out;
    8: reg_1012 <= op2_00_out;
    15: reg_1012 <= op2_00_out;
    39: reg_1012 <= op2_00_out;
    77: reg_1012 <= op2_00_out;
    endcase
  end

  // REG#1013の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1013 <= op2_01_out;
    9: reg_1013 <= op2_01_out;
    19: reg_1013 <= op2_01_out;
    52: reg_1013 <= op2_01_out;
    78: reg_1013 <= op2_01_out;
    endcase
  end

  // REG#1014の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_1014 <= op2_02_out;
    10: reg_1014 <= op2_02_out;
    23: reg_1014 <= op2_02_out;
    69: reg_1014 <= imem01_in[35:32];
    94: reg_1014 <= imem01_in[35:32];
    endcase
  end

  // REG#1015の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_1015 <= imem05_in[47:44];
    10: reg_1015 <= imem01_in[91:88];
    40: reg_1015 <= imem01_in[91:88];
    51: reg_1015 <= imem01_in[91:88];
    59: reg_1015 <= imem05_in[47:44];
    61: reg_1015 <= imem01_in[91:88];
    65: reg_1015 <= imem01_in[91:88];
    68: reg_1015 <= imem05_in[47:44];
    73: reg_1015 <= imem01_in[91:88];
    76: reg_1015 <= imem05_in[47:44];
    79: reg_1015 <= imem05_in[47:44];
    86: reg_1015 <= imem01_in[91:88];
    90: reg_1015 <= imem01_in[91:88];
    96: reg_1015 <= imem01_in[91:88];
    endcase
  end

  // REG#1016の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_1016 <= imem05_in[51:48];
    10: reg_1016 <= imem05_in[51:48];
    14: reg_1016 <= imem05_in[51:48];
    16: reg_1016 <= imem05_in[51:48];
    24: reg_1016 <= imem04_in[103:100];
    85: reg_1016 <= imem04_in[103:100];
    94: reg_1016 <= imem04_in[103:100];
    endcase
  end

  // REG#1017の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_1017 <= imem05_in[67:64];
    10: reg_1017 <= imem01_in[111:108];
    38: reg_1017 <= imem01_in[111:108];
    41: reg_1017 <= imem01_in[111:108];
    endcase
  end

  // REG#1018の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_1018 <= imem06_in[43:40];
    10: reg_1018 <= imem01_in[119:116];
    39: reg_1018 <= imem01_in[119:116];
    44: reg_1018 <= imem06_in[43:40];
    46: reg_1018 <= imem06_in[43:40];
    48: reg_1018 <= imem01_in[119:116];
    52: reg_1018 <= imem01_in[119:116];
    55: reg_1018 <= imem01_in[119:116];
    57: reg_1018 <= imem06_in[43:40];
    endcase
  end

  // REG#1019の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_1019 <= imem06_in[27:24];
    10: reg_1019 <= op1_12_out;
    18: reg_1019 <= imem06_in[27:24];
    20: reg_1019 <= imem06_in[27:24];
    22: reg_1019 <= imem06_in[27:24];
    23: reg_1019 <= op1_12_out;
    31: reg_1019 <= imem03_in[59:56];
    54: reg_1019 <= imem03_in[59:56];
    57: reg_1019 <= imem06_in[27:24];
    endcase
  end

  // REG#1020の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_1020 <= imem06_in[23:20];
    11: reg_1020 <= imem05_in[11:8];
    14: reg_1020 <= imem05_in[11:8];
    18: reg_1020 <= imem05_in[11:8];
    20: reg_1020 <= imem06_in[23:20];
    24: reg_1020 <= imem04_in[79:76];
    84: reg_1020 <= imem04_in[79:76];
    86: reg_1020 <= imem05_in[11:8];
    89: reg_1020 <= imem06_in[23:20];
    endcase
  end

  // REG#1021の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_1021 <= imem06_in[55:52];
    11: reg_1021 <= imem05_in[3:0];
    14: reg_1021 <= imem05_in[3:0];
    16: reg_1021 <= imem05_in[3:0];
    20: reg_1021 <= imem05_in[3:0];
    49: reg_1021 <= imem06_in[55:52];
    52: reg_1021 <= imem05_in[3:0];
    56: reg_1021 <= imem05_in[3:0];
    66: reg_1021 <= imem06_in[55:52];
    68: reg_1021 <= imem06_in[55:52];
    70: reg_1021 <= imem06_in[55:52];
    73: reg_1021 <= imem05_in[3:0];
    endcase
  end

  // REG#1022の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_1022 <= op1_14_out;
    10: reg_1022 <= op1_14_out;
    13: reg_1022 <= op1_14_out;
    18: reg_1022 <= op1_14_out;
    21: reg_1022 <= op1_14_out;
    25: reg_1022 <= op1_14_out;
    29: reg_1022 <= op1_14_out;
    32: reg_1022 <= op1_14_out;
    62: reg_1022 <= op1_14_out;
    69: reg_1022 <= imem01_in[87:84];
    96: reg_1022 <= imem01_in[87:84];
    endcase
  end

  // REG#1023の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_1023 <= op1_15_out;
    10: reg_1023 <= op1_15_out;
    13: reg_1023 <= op1_15_out;
    18: reg_1023 <= op1_15_out;
    21: reg_1023 <= op1_15_out;
    27: reg_1023 <= op1_15_out;
    30: reg_1023 <= op1_15_out;
    33: reg_1023 <= op1_15_out;
    64: reg_1023 <= op1_15_out;
    69: reg_1023 <= imem01_in[63:60];
    endcase
  end

  // REG#1024の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_1024 <= op2_00_out;
    11: reg_1024 <= op2_00_out;
    25: reg_1024 <= op2_00_out;
    29: reg_1024 <= op2_00_out;
    43: reg_1024 <= op2_00_out;
    48: reg_1024 <= op2_00_out;
    69: reg_1024 <= imem01_in[103:100];
    96: reg_1024 <= op2_00_out;
    endcase
  end

  // REG#1025の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_1025 <= op2_01_out;
    12: reg_1025 <= op2_01_out;
    29: reg_1025 <= op2_01_out;
    44: reg_1025 <= op2_01_out;
    54: reg_1025 <= op2_01_out;
    83: reg_1025 <= op2_01_out;
    endcase
  end

  // REG#1026の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_1026 <= op2_02_out;
    13: reg_1026 <= op2_02_out;
    33: reg_1026 <= op2_02_out;
    59: reg_1026 <= op2_02_out;
    endcase
  end

  // REG#1027の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_1027 <= op2_03_out;
    15: reg_1027 <= op2_03_out;
    44: reg_1027 <= op2_03_out;
    62: reg_1027 <= op2_03_out;
    69: reg_1027 <= op2_03_out;
    90: reg_1027 <= op2_03_out;
    endcase
  end

  // REG#1028の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_1028 <= imem06_in[47:44];
    32: reg_1028 <= imem06_in[47:44];
    38: reg_1028 <= imem06_in[47:44];
    46: reg_1028 <= imem06_in[47:44];
    52: reg_1028 <= imem06_in[47:44];
    54: reg_1028 <= imem06_in[47:44];
    61: reg_1028 <= imem06_in[47:44];
    73: reg_1028 <= imem06_in[47:44];
    77: reg_1028 <= imem06_in[47:44];
    86: reg_1028 <= imem06_in[47:44];
    endcase
  end

  // REG#1029の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_1029 <= imem06_in[3:0];
    33: reg_1029 <= imem06_in[3:0];
    37: reg_1029 <= imem06_in[3:0];
    61: reg_1029 <= imem06_in[3:0];
    73: reg_1029 <= imem06_in[3:0];
    76: reg_1029 <= imem06_in[3:0];
    83: reg_1029 <= imem06_in[3:0];
    89: reg_1029 <= imem06_in[3:0];
    endcase
  end

  // REG#1030の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_1030 <= imem06_in[15:12];
    35: reg_1030 <= imem06_in[15:12];
    44: reg_1030 <= imem06_in[15:12];
    50: reg_1030 <= imem06_in[15:12];
    55: reg_1030 <= imem06_in[15:12];
    58: reg_1030 <= imem06_in[15:12];
    94: reg_1030 <= imem06_in[15:12];
    endcase
  end

  // REG#1031の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1031 <= imem01_in[79:76];
    41: reg_1031 <= imem01_in[79:76];
    93: reg_1031 <= imem01_in[79:76];
    endcase
  end

  // REG#1032の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1032 <= imem01_in[23:20];
    43: reg_1032 <= imem01_in[23:20];
    55: reg_1032 <= imem01_in[23:20];
    69: reg_1032 <= imem01_in[23:20];
    endcase
  end

  // REG#1033の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1033 <= imem01_in[47:44];
    48: reg_1033 <= imem01_in[47:44];
    53: reg_1033 <= imem01_in[47:44];
    endcase
  end

  // REG#1034の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1034 <= imem01_in[127:124];
    39: reg_1034 <= imem01_in[127:124];
    44: reg_1034 <= imem01_in[127:124];
    49: reg_1034 <= imem01_in[127:124];
    70: reg_1034 <= imem01_in[127:124];
    76: reg_1034 <= imem01_in[127:124];
    94: reg_1034 <= imem01_in[127:124];
    endcase
  end

  // REG#1035の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1035 <= imem01_in[75:72];
    47: reg_1035 <= imem01_in[75:72];
    49: reg_1035 <= imem01_in[75:72];
    69: reg_1035 <= imem01_in[75:72];
    endcase
  end

  // REG#1036の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1036 <= imem01_in[87:84];
    43: reg_1036 <= imem01_in[87:84];
    47: reg_1036 <= imem01_in[87:84];
    49: reg_1036 <= imem01_in[87:84];
    70: reg_1036 <= imem01_in[87:84];
    73: reg_1036 <= imem01_in[87:84];
    86: reg_1036 <= imem01_in[87:84];
    90: reg_1036 <= imem01_in[87:84];
    endcase
  end

  // REG#1037の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1037 <= imem01_in[59:56];
    41: reg_1037 <= imem01_in[59:56];
    endcase
  end

  // REG#1038の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1038 <= imem01_in[115:112];
    44: reg_1038 <= imem01_in[115:112];
    56: reg_1038 <= imem01_in[115:112];
    68: reg_1038 <= imem01_in[115:112];
    73: reg_1038 <= imem01_in[115:112];
    76: reg_1038 <= imem01_in[115:112];
    78: reg_1038 <= imem01_in[115:112];
    82: reg_1038 <= imem01_in[115:112];
    86: reg_1038 <= imem01_in[115:112];
    93: reg_1038 <= imem01_in[115:112];
    endcase
  end

  // REG#1039の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1039 <= imem01_in[7:4];
    41: reg_1039 <= imem01_in[7:4];
    94: reg_1039 <= imem01_in[7:4];
    endcase
  end

  // REG#1040の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1040 <= imem01_in[71:68];
    41: reg_1040 <= imem01_in[71:68];
    94: reg_1040 <= imem01_in[71:68];
    endcase
  end

  // REG#1041の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1041 <= imem01_in[99:96];
    41: reg_1041 <= imem01_in[99:96];
    94: reg_1041 <= imem01_in[99:96];
    endcase
  end

  // REG#1042の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1042 <= imem01_in[15:12];
    42: reg_1042 <= imem01_in[15:12];
    45: reg_1042 <= imem01_in[15:12];
    52: reg_1042 <= imem01_in[15:12];
    55: reg_1042 <= imem01_in[15:12];
    57: reg_1042 <= imem01_in[15:12];
    59: reg_1042 <= imem01_in[15:12];
    67: reg_1042 <= imem01_in[15:12];
    69: reg_1042 <= imem01_in[15:12];
    endcase
  end

  // REG#1043の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1043 <= imem01_in[39:36];
    41: reg_1043 <= imem01_in[39:36];
    endcase
  end

  // REG#1044の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1044 <= imem01_in[43:40];
    43: reg_1044 <= imem01_in[43:40];
    49: reg_1044 <= imem01_in[43:40];
    64: reg_1044 <= imem01_in[43:40];
    69: reg_1044 <= imem01_in[43:40];
    endcase
  end

  // REG#1045の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1045 <= imem01_in[95:92];
    43: reg_1045 <= imem01_in[95:92];
    49: reg_1045 <= imem01_in[95:92];
    72: reg_1045 <= imem01_in[95:92];
    78: reg_1045 <= imem01_in[95:92];
    80: reg_1045 <= imem01_in[95:92];
    83: reg_1045 <= imem01_in[95:92];
    87: reg_1045 <= imem01_in[95:92];
    93: reg_1045 <= imem01_in[95:92];
    endcase
  end

  // REG#1046の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_1046 <= imem05_in[99:96];
    18: reg_1046 <= imem05_in[99:96];
    20: reg_1046 <= imem05_in[99:96];
    50: reg_1046 <= imem05_in[99:96];
    66: reg_1046 <= imem05_in[99:96];
    79: reg_1046 <= imem05_in[99:96];
    92: reg_1046 <= imem05_in[99:96];
    endcase
  end

  // REG#1047の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1047 <= op2_00_out;
    21: reg_1047 <= op2_00_out;
    58: reg_1047 <= op2_00_out;
    endcase
  end

  // REG#1048の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1048 <= op2_01_out;
    22: reg_1048 <= op2_01_out;
    63: reg_1048 <= op2_01_out;
    72: reg_1048 <= op2_01_out;
    endcase
  end

  // REG#1049の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_1049 <= imem01_in[35:32];
    24: reg_1049 <= imem01_in[35:32];
    29: reg_1049 <= imem01_in[35:32];
    31: reg_1049 <= imem03_in[63:60];
    57: reg_1049 <= imem03_in[63:60];
    60: reg_1049 <= imem03_in[63:60];
    63: reg_1049 <= imem01_in[35:32];
    68: reg_1049 <= imem03_in[63:60];
    70: reg_1049 <= imem03_in[63:60];
    endcase
  end

  // REG#1050の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_1050 <= imem01_in[115:112];
    28: reg_1050 <= imem01_in[115:112];
    31: reg_1050 <= imem03_in[31:28];
    56: reg_1050 <= imem03_in[31:28];
    58: reg_1050 <= imem03_in[31:28];
    60: reg_1050 <= imem03_in[31:28];
    71: reg_1050 <= imem03_in[31:28];
    76: reg_1050 <= imem03_in[31:28];
    82: reg_1050 <= imem03_in[31:28];
    88: reg_1050 <= imem03_in[31:28];
    endcase
  end

  // REG#1051の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_1051 <= imem01_in[11:8];
    29: reg_1051 <= imem01_in[11:8];
    32: reg_1051 <= imem01_in[11:8];
    37: reg_1051 <= imem01_in[11:8];
    39: reg_1051 <= imem01_in[11:8];
    43: reg_1051 <= imem01_in[11:8];
    45: reg_1051 <= imem01_in[11:8];
    47: reg_1051 <= imem01_in[11:8];
    53: reg_1051 <= imem01_in[11:8];
    endcase
  end

  // REG#1052の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_1052 <= imem01_in[107:104];
    27: reg_1052 <= imem01_in[107:104];
    29: reg_1052 <= imem01_in[107:104];
    35: reg_1052 <= imem01_in[107:104];
    49: reg_1052 <= imem01_in[107:104];
    68: reg_1052 <= imem01_in[107:104];
    80: reg_1052 <= imem01_in[107:104];
    82: reg_1052 <= imem01_in[107:104];
    86: reg_1052 <= imem01_in[107:104];
    endcase
  end

  // REG#1053の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_1053 <= imem01_in[39:36];
    28: reg_1053 <= imem01_in[39:36];
    35: reg_1053 <= imem01_in[39:36];
    37: reg_1053 <= imem01_in[39:36];
    42: reg_1053 <= imem01_in[39:36];
    45: reg_1053 <= imem01_in[39:36];
    47: reg_1053 <= imem01_in[39:36];
    51: reg_1053 <= imem01_in[39:36];
    53: reg_1053 <= imem01_in[39:36];
    endcase
  end

  // REG#1054の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_1054 <= op2_03_out;
    27: reg_1054 <= op2_03_out;
    47: reg_1054 <= op2_03_out;
    72: reg_1054 <= op2_03_out;
    endcase
  end

  // REG#1055の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_1055 <= imem01_in[15:12];
    28: reg_1055 <= imem01_in[15:12];
    34: reg_1055 <= imem01_in[15:12];
    53: reg_1055 <= imem01_in[15:12];
    endcase
  end

  // REG#1056の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_1056 <= imem01_in[67:64];
    26: reg_1056 <= imem01_in[67:64];
    28: reg_1056 <= imem01_in[67:64];
    35: reg_1056 <= imem01_in[67:64];
    37: reg_1056 <= imem01_in[67:64];
    39: reg_1056 <= imem01_in[67:64];
    49: reg_1056 <= imem01_in[67:64];
    69: reg_1056 <= imem01_in[67:64];
    93: reg_1056 <= imem01_in[67:64];
    endcase
  end

  // REG#1057の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_1057 <= imem04_in[75:72];
    89: reg_1057 <= imem04_in[75:72];
    endcase
  end
endmodule
