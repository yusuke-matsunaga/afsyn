module affine2(
  input clock,
  input reset,
  input start,
  output busy,
  output [1:0] imem00_bank,
  output imem00_rd,
  input [127:0] imem00_in,
  output [1:0] imem01_bank,
  output imem01_rd,
  input [127:0] imem01_in,
  output [1:0] imem02_bank,
  output imem02_rd,
  input [127:0] imem02_in,
  output [1:0] imem03_bank,
  output imem03_rd,
  input [127:0] imem03_in,
  output [1:0] imem04_bank,
  output imem04_rd,
  input [127:0] imem04_in,
  output [1:0] imem05_bank,
  output imem05_rd,
  input [127:0] imem05_in,
  output [1:0] imem06_bank,
  output imem06_rd,
  input [127:0] imem06_in,
  output [1:0] imem07_bank,
  output imem07_rd,
  input [127:0] imem07_in,
  output [5:0] omem00_bank,
  output omem00_wr,
  output [8:0] omem00_out,
  output [5:0] omem01_bank,
  output omem01_wr,
  output [8:0] omem01_out,
  output [5:0] omem02_bank,
  output omem02_wr,
  output [8:0] omem02_out,
  output [5:0] omem03_bank,
  output omem03_wr,
  output [8:0] omem03_out,
  output [5:0] omem04_bank,
  output omem04_wr,
  output [8:0] omem04_out);


  // 0 番目の OP1
  reg [3:0] op1_00_in00;
  reg       op1_00_inv00;
  reg [3:0] op1_00_in01;
  reg       op1_00_inv01;
  reg [3:0] op1_00_in02;
  reg       op1_00_inv02;
  reg [3:0] op1_00_in03;
  reg       op1_00_inv03;
  reg [3:0] op1_00_in04;
  reg       op1_00_inv04;
  reg [3:0] op1_00_in05;
  reg       op1_00_inv05;
  reg [3:0] op1_00_in06;
  reg       op1_00_inv06;
  reg [3:0] op1_00_in07;
  reg       op1_00_inv07;
  reg [3:0] op1_00_in08;
  reg       op1_00_inv08;
  reg [3:0] op1_00_in09;
  reg       op1_00_inv09;
  reg [3:0] op1_00_in10;
  reg       op1_00_inv10;
  reg [3:0] op1_00_in11;
  reg       op1_00_inv11;
  reg [3:0] op1_00_in12;
  reg       op1_00_inv12;
  reg [3:0] op1_00_in13;
  reg       op1_00_inv13;
  reg [3:0] op1_00_in14;
  reg       op1_00_inv14;
  reg [3:0] op1_00_in15;
  reg       op1_00_inv15;
  reg [3:0] op1_00_in16;
  reg       op1_00_inv16;
  reg [3:0] op1_00_in17;
  reg       op1_00_inv17;
  reg [3:0] op1_00_in18;
  reg       op1_00_inv18;
  reg [3:0] op1_00_in19;
  reg       op1_00_inv19;
  reg [3:0] op1_00_in20;
  reg       op1_00_inv20;
  reg [3:0] op1_00_in21;
  reg       op1_00_inv21;
  reg [3:0] op1_00_in22;
  reg       op1_00_inv22;
  reg [3:0] op1_00_in23;
  reg       op1_00_inv23;
  reg [3:0] op1_00_in24;
  reg       op1_00_inv24;
  reg [3:0] op1_00_in25;
  reg       op1_00_inv25;
  reg [3:0] op1_00_in26;
  reg       op1_00_inv26;
  reg [3:0] op1_00_in27;
  reg       op1_00_inv27;
  reg [3:0] op1_00_in28;
  reg       op1_00_inv28;
  reg [3:0] op1_00_in29;
  reg       op1_00_inv29;
  reg [3:0] op1_00_in30;
  reg       op1_00_inv30;
  reg [3:0] op1_00_in31;
  reg       op1_00_inv31;
  wire [8:0] op1_00_out;
  op1 op1_00(
    .data0_in(op1_00_in00),
    .inv0_in(op1_00_inv00),
    .data1_in(op1_00_in01),
    .inv1_in(op1_00_inv01),
    .data2_in(op1_00_in02),
    .inv2_in(op1_00_inv02),
    .data3_in(op1_00_in03),
    .inv3_in(op1_00_inv03),
    .data4_in(op1_00_in04),
    .inv4_in(op1_00_inv04),
    .data5_in(op1_00_in05),
    .inv5_in(op1_00_inv05),
    .data6_in(op1_00_in06),
    .inv6_in(op1_00_inv06),
    .data7_in(op1_00_in07),
    .inv7_in(op1_00_inv07),
    .data8_in(op1_00_in08),
    .inv8_in(op1_00_inv08),
    .data9_in(op1_00_in09),
    .inv9_in(op1_00_inv09),
    .data10_in(op1_00_in10),
    .inv10_in(op1_00_inv10),
    .data11_in(op1_00_in11),
    .inv11_in(op1_00_inv11),
    .data12_in(op1_00_in12),
    .inv12_in(op1_00_inv12),
    .data13_in(op1_00_in13),
    .inv13_in(op1_00_inv13),
    .data14_in(op1_00_in14),
    .inv14_in(op1_00_inv14),
    .data15_in(op1_00_in15),
    .inv15_in(op1_00_inv15),
    .data16_in(op1_00_in16),
    .inv16_in(op1_00_inv16),
    .data17_in(op1_00_in17),
    .inv17_in(op1_00_inv17),
    .data18_in(op1_00_in18),
    .inv18_in(op1_00_inv18),
    .data19_in(op1_00_in19),
    .inv19_in(op1_00_inv19),
    .data20_in(op1_00_in20),
    .inv20_in(op1_00_inv20),
    .data21_in(op1_00_in21),
    .inv21_in(op1_00_inv21),
    .data22_in(op1_00_in22),
    .inv22_in(op1_00_inv22),
    .data23_in(op1_00_in23),
    .inv23_in(op1_00_inv23),
    .data24_in(op1_00_in24),
    .inv24_in(op1_00_inv24),
    .data25_in(op1_00_in25),
    .inv25_in(op1_00_inv25),
    .data26_in(op1_00_in26),
    .inv26_in(op1_00_inv26),
    .data27_in(op1_00_in27),
    .inv27_in(op1_00_inv27),
    .data28_in(op1_00_in28),
    .inv28_in(op1_00_inv28),
    .data29_in(op1_00_in29),
    .inv29_in(op1_00_inv29),
    .data30_in(op1_00_in30),
    .inv30_in(op1_00_inv30),
    .data31_in(op1_00_in31),
    .inv31_in(op1_00_inv31),
    .data_out(op1_00_out));

  // 1 番目の OP1
  reg [3:0] op1_01_in00;
  reg       op1_01_inv00;
  reg [3:0] op1_01_in01;
  reg       op1_01_inv01;
  reg [3:0] op1_01_in02;
  reg       op1_01_inv02;
  reg [3:0] op1_01_in03;
  reg       op1_01_inv03;
  reg [3:0] op1_01_in04;
  reg       op1_01_inv04;
  reg [3:0] op1_01_in05;
  reg       op1_01_inv05;
  reg [3:0] op1_01_in06;
  reg       op1_01_inv06;
  reg [3:0] op1_01_in07;
  reg       op1_01_inv07;
  reg [3:0] op1_01_in08;
  reg       op1_01_inv08;
  reg [3:0] op1_01_in09;
  reg       op1_01_inv09;
  reg [3:0] op1_01_in10;
  reg       op1_01_inv10;
  reg [3:0] op1_01_in11;
  reg       op1_01_inv11;
  reg [3:0] op1_01_in12;
  reg       op1_01_inv12;
  reg [3:0] op1_01_in13;
  reg       op1_01_inv13;
  reg [3:0] op1_01_in14;
  reg       op1_01_inv14;
  reg [3:0] op1_01_in15;
  reg       op1_01_inv15;
  reg [3:0] op1_01_in16;
  reg       op1_01_inv16;
  reg [3:0] op1_01_in17;
  reg       op1_01_inv17;
  reg [3:0] op1_01_in18;
  reg       op1_01_inv18;
  reg [3:0] op1_01_in19;
  reg       op1_01_inv19;
  reg [3:0] op1_01_in20;
  reg       op1_01_inv20;
  reg [3:0] op1_01_in21;
  reg       op1_01_inv21;
  reg [3:0] op1_01_in22;
  reg       op1_01_inv22;
  reg [3:0] op1_01_in23;
  reg       op1_01_inv23;
  reg [3:0] op1_01_in24;
  reg       op1_01_inv24;
  reg [3:0] op1_01_in25;
  reg       op1_01_inv25;
  reg [3:0] op1_01_in26;
  reg       op1_01_inv26;
  reg [3:0] op1_01_in27;
  reg       op1_01_inv27;
  reg [3:0] op1_01_in28;
  reg       op1_01_inv28;
  reg [3:0] op1_01_in29;
  reg       op1_01_inv29;
  reg [3:0] op1_01_in30;
  reg       op1_01_inv30;
  reg [3:0] op1_01_in31;
  reg       op1_01_inv31;
  wire [8:0] op1_01_out;
  op1 op1_01(
    .data0_in(op1_01_in00),
    .inv0_in(op1_01_inv00),
    .data1_in(op1_01_in01),
    .inv1_in(op1_01_inv01),
    .data2_in(op1_01_in02),
    .inv2_in(op1_01_inv02),
    .data3_in(op1_01_in03),
    .inv3_in(op1_01_inv03),
    .data4_in(op1_01_in04),
    .inv4_in(op1_01_inv04),
    .data5_in(op1_01_in05),
    .inv5_in(op1_01_inv05),
    .data6_in(op1_01_in06),
    .inv6_in(op1_01_inv06),
    .data7_in(op1_01_in07),
    .inv7_in(op1_01_inv07),
    .data8_in(op1_01_in08),
    .inv8_in(op1_01_inv08),
    .data9_in(op1_01_in09),
    .inv9_in(op1_01_inv09),
    .data10_in(op1_01_in10),
    .inv10_in(op1_01_inv10),
    .data11_in(op1_01_in11),
    .inv11_in(op1_01_inv11),
    .data12_in(op1_01_in12),
    .inv12_in(op1_01_inv12),
    .data13_in(op1_01_in13),
    .inv13_in(op1_01_inv13),
    .data14_in(op1_01_in14),
    .inv14_in(op1_01_inv14),
    .data15_in(op1_01_in15),
    .inv15_in(op1_01_inv15),
    .data16_in(op1_01_in16),
    .inv16_in(op1_01_inv16),
    .data17_in(op1_01_in17),
    .inv17_in(op1_01_inv17),
    .data18_in(op1_01_in18),
    .inv18_in(op1_01_inv18),
    .data19_in(op1_01_in19),
    .inv19_in(op1_01_inv19),
    .data20_in(op1_01_in20),
    .inv20_in(op1_01_inv20),
    .data21_in(op1_01_in21),
    .inv21_in(op1_01_inv21),
    .data22_in(op1_01_in22),
    .inv22_in(op1_01_inv22),
    .data23_in(op1_01_in23),
    .inv23_in(op1_01_inv23),
    .data24_in(op1_01_in24),
    .inv24_in(op1_01_inv24),
    .data25_in(op1_01_in25),
    .inv25_in(op1_01_inv25),
    .data26_in(op1_01_in26),
    .inv26_in(op1_01_inv26),
    .data27_in(op1_01_in27),
    .inv27_in(op1_01_inv27),
    .data28_in(op1_01_in28),
    .inv28_in(op1_01_inv28),
    .data29_in(op1_01_in29),
    .inv29_in(op1_01_inv29),
    .data30_in(op1_01_in30),
    .inv30_in(op1_01_inv30),
    .data31_in(op1_01_in31),
    .inv31_in(op1_01_inv31),
    .data_out(op1_01_out));

  // 2 番目の OP1
  reg [3:0] op1_02_in00;
  reg       op1_02_inv00;
  reg [3:0] op1_02_in01;
  reg       op1_02_inv01;
  reg [3:0] op1_02_in02;
  reg       op1_02_inv02;
  reg [3:0] op1_02_in03;
  reg       op1_02_inv03;
  reg [3:0] op1_02_in04;
  reg       op1_02_inv04;
  reg [3:0] op1_02_in05;
  reg       op1_02_inv05;
  reg [3:0] op1_02_in06;
  reg       op1_02_inv06;
  reg [3:0] op1_02_in07;
  reg       op1_02_inv07;
  reg [3:0] op1_02_in08;
  reg       op1_02_inv08;
  reg [3:0] op1_02_in09;
  reg       op1_02_inv09;
  reg [3:0] op1_02_in10;
  reg       op1_02_inv10;
  reg [3:0] op1_02_in11;
  reg       op1_02_inv11;
  reg [3:0] op1_02_in12;
  reg       op1_02_inv12;
  reg [3:0] op1_02_in13;
  reg       op1_02_inv13;
  reg [3:0] op1_02_in14;
  reg       op1_02_inv14;
  reg [3:0] op1_02_in15;
  reg       op1_02_inv15;
  reg [3:0] op1_02_in16;
  reg       op1_02_inv16;
  reg [3:0] op1_02_in17;
  reg       op1_02_inv17;
  reg [3:0] op1_02_in18;
  reg       op1_02_inv18;
  reg [3:0] op1_02_in19;
  reg       op1_02_inv19;
  reg [3:0] op1_02_in20;
  reg       op1_02_inv20;
  reg [3:0] op1_02_in21;
  reg       op1_02_inv21;
  reg [3:0] op1_02_in22;
  reg       op1_02_inv22;
  reg [3:0] op1_02_in23;
  reg       op1_02_inv23;
  reg [3:0] op1_02_in24;
  reg       op1_02_inv24;
  reg [3:0] op1_02_in25;
  reg       op1_02_inv25;
  reg [3:0] op1_02_in26;
  reg       op1_02_inv26;
  reg [3:0] op1_02_in27;
  reg       op1_02_inv27;
  reg [3:0] op1_02_in28;
  reg       op1_02_inv28;
  reg [3:0] op1_02_in29;
  reg       op1_02_inv29;
  reg [3:0] op1_02_in30;
  reg       op1_02_inv30;
  reg [3:0] op1_02_in31;
  reg       op1_02_inv31;
  wire [8:0] op1_02_out;
  op1 op1_02(
    .data0_in(op1_02_in00),
    .inv0_in(op1_02_inv00),
    .data1_in(op1_02_in01),
    .inv1_in(op1_02_inv01),
    .data2_in(op1_02_in02),
    .inv2_in(op1_02_inv02),
    .data3_in(op1_02_in03),
    .inv3_in(op1_02_inv03),
    .data4_in(op1_02_in04),
    .inv4_in(op1_02_inv04),
    .data5_in(op1_02_in05),
    .inv5_in(op1_02_inv05),
    .data6_in(op1_02_in06),
    .inv6_in(op1_02_inv06),
    .data7_in(op1_02_in07),
    .inv7_in(op1_02_inv07),
    .data8_in(op1_02_in08),
    .inv8_in(op1_02_inv08),
    .data9_in(op1_02_in09),
    .inv9_in(op1_02_inv09),
    .data10_in(op1_02_in10),
    .inv10_in(op1_02_inv10),
    .data11_in(op1_02_in11),
    .inv11_in(op1_02_inv11),
    .data12_in(op1_02_in12),
    .inv12_in(op1_02_inv12),
    .data13_in(op1_02_in13),
    .inv13_in(op1_02_inv13),
    .data14_in(op1_02_in14),
    .inv14_in(op1_02_inv14),
    .data15_in(op1_02_in15),
    .inv15_in(op1_02_inv15),
    .data16_in(op1_02_in16),
    .inv16_in(op1_02_inv16),
    .data17_in(op1_02_in17),
    .inv17_in(op1_02_inv17),
    .data18_in(op1_02_in18),
    .inv18_in(op1_02_inv18),
    .data19_in(op1_02_in19),
    .inv19_in(op1_02_inv19),
    .data20_in(op1_02_in20),
    .inv20_in(op1_02_inv20),
    .data21_in(op1_02_in21),
    .inv21_in(op1_02_inv21),
    .data22_in(op1_02_in22),
    .inv22_in(op1_02_inv22),
    .data23_in(op1_02_in23),
    .inv23_in(op1_02_inv23),
    .data24_in(op1_02_in24),
    .inv24_in(op1_02_inv24),
    .data25_in(op1_02_in25),
    .inv25_in(op1_02_inv25),
    .data26_in(op1_02_in26),
    .inv26_in(op1_02_inv26),
    .data27_in(op1_02_in27),
    .inv27_in(op1_02_inv27),
    .data28_in(op1_02_in28),
    .inv28_in(op1_02_inv28),
    .data29_in(op1_02_in29),
    .inv29_in(op1_02_inv29),
    .data30_in(op1_02_in30),
    .inv30_in(op1_02_inv30),
    .data31_in(op1_02_in31),
    .inv31_in(op1_02_inv31),
    .data_out(op1_02_out));

  // 3 番目の OP1
  reg [3:0] op1_03_in00;
  reg       op1_03_inv00;
  reg [3:0] op1_03_in01;
  reg       op1_03_inv01;
  reg [3:0] op1_03_in02;
  reg       op1_03_inv02;
  reg [3:0] op1_03_in03;
  reg       op1_03_inv03;
  reg [3:0] op1_03_in04;
  reg       op1_03_inv04;
  reg [3:0] op1_03_in05;
  reg       op1_03_inv05;
  reg [3:0] op1_03_in06;
  reg       op1_03_inv06;
  reg [3:0] op1_03_in07;
  reg       op1_03_inv07;
  reg [3:0] op1_03_in08;
  reg       op1_03_inv08;
  reg [3:0] op1_03_in09;
  reg       op1_03_inv09;
  reg [3:0] op1_03_in10;
  reg       op1_03_inv10;
  reg [3:0] op1_03_in11;
  reg       op1_03_inv11;
  reg [3:0] op1_03_in12;
  reg       op1_03_inv12;
  reg [3:0] op1_03_in13;
  reg       op1_03_inv13;
  reg [3:0] op1_03_in14;
  reg       op1_03_inv14;
  reg [3:0] op1_03_in15;
  reg       op1_03_inv15;
  reg [3:0] op1_03_in16;
  reg       op1_03_inv16;
  reg [3:0] op1_03_in17;
  reg       op1_03_inv17;
  reg [3:0] op1_03_in18;
  reg       op1_03_inv18;
  reg [3:0] op1_03_in19;
  reg       op1_03_inv19;
  reg [3:0] op1_03_in20;
  reg       op1_03_inv20;
  reg [3:0] op1_03_in21;
  reg       op1_03_inv21;
  reg [3:0] op1_03_in22;
  reg       op1_03_inv22;
  reg [3:0] op1_03_in23;
  reg       op1_03_inv23;
  reg [3:0] op1_03_in24;
  reg       op1_03_inv24;
  reg [3:0] op1_03_in25;
  reg       op1_03_inv25;
  reg [3:0] op1_03_in26;
  reg       op1_03_inv26;
  reg [3:0] op1_03_in27;
  reg       op1_03_inv27;
  reg [3:0] op1_03_in28;
  reg       op1_03_inv28;
  reg [3:0] op1_03_in29;
  reg       op1_03_inv29;
  reg [3:0] op1_03_in30;
  reg       op1_03_inv30;
  reg [3:0] op1_03_in31;
  reg       op1_03_inv31;
  wire [8:0] op1_03_out;
  op1 op1_03(
    .data0_in(op1_03_in00),
    .inv0_in(op1_03_inv00),
    .data1_in(op1_03_in01),
    .inv1_in(op1_03_inv01),
    .data2_in(op1_03_in02),
    .inv2_in(op1_03_inv02),
    .data3_in(op1_03_in03),
    .inv3_in(op1_03_inv03),
    .data4_in(op1_03_in04),
    .inv4_in(op1_03_inv04),
    .data5_in(op1_03_in05),
    .inv5_in(op1_03_inv05),
    .data6_in(op1_03_in06),
    .inv6_in(op1_03_inv06),
    .data7_in(op1_03_in07),
    .inv7_in(op1_03_inv07),
    .data8_in(op1_03_in08),
    .inv8_in(op1_03_inv08),
    .data9_in(op1_03_in09),
    .inv9_in(op1_03_inv09),
    .data10_in(op1_03_in10),
    .inv10_in(op1_03_inv10),
    .data11_in(op1_03_in11),
    .inv11_in(op1_03_inv11),
    .data12_in(op1_03_in12),
    .inv12_in(op1_03_inv12),
    .data13_in(op1_03_in13),
    .inv13_in(op1_03_inv13),
    .data14_in(op1_03_in14),
    .inv14_in(op1_03_inv14),
    .data15_in(op1_03_in15),
    .inv15_in(op1_03_inv15),
    .data16_in(op1_03_in16),
    .inv16_in(op1_03_inv16),
    .data17_in(op1_03_in17),
    .inv17_in(op1_03_inv17),
    .data18_in(op1_03_in18),
    .inv18_in(op1_03_inv18),
    .data19_in(op1_03_in19),
    .inv19_in(op1_03_inv19),
    .data20_in(op1_03_in20),
    .inv20_in(op1_03_inv20),
    .data21_in(op1_03_in21),
    .inv21_in(op1_03_inv21),
    .data22_in(op1_03_in22),
    .inv22_in(op1_03_inv22),
    .data23_in(op1_03_in23),
    .inv23_in(op1_03_inv23),
    .data24_in(op1_03_in24),
    .inv24_in(op1_03_inv24),
    .data25_in(op1_03_in25),
    .inv25_in(op1_03_inv25),
    .data26_in(op1_03_in26),
    .inv26_in(op1_03_inv26),
    .data27_in(op1_03_in27),
    .inv27_in(op1_03_inv27),
    .data28_in(op1_03_in28),
    .inv28_in(op1_03_inv28),
    .data29_in(op1_03_in29),
    .inv29_in(op1_03_inv29),
    .data30_in(op1_03_in30),
    .inv30_in(op1_03_inv30),
    .data31_in(op1_03_in31),
    .inv31_in(op1_03_inv31),
    .data_out(op1_03_out));

  // 4 番目の OP1
  reg [3:0] op1_04_in00;
  reg       op1_04_inv00;
  reg [3:0] op1_04_in01;
  reg       op1_04_inv01;
  reg [3:0] op1_04_in02;
  reg       op1_04_inv02;
  reg [3:0] op1_04_in03;
  reg       op1_04_inv03;
  reg [3:0] op1_04_in04;
  reg       op1_04_inv04;
  reg [3:0] op1_04_in05;
  reg       op1_04_inv05;
  reg [3:0] op1_04_in06;
  reg       op1_04_inv06;
  reg [3:0] op1_04_in07;
  reg       op1_04_inv07;
  reg [3:0] op1_04_in08;
  reg       op1_04_inv08;
  reg [3:0] op1_04_in09;
  reg       op1_04_inv09;
  reg [3:0] op1_04_in10;
  reg       op1_04_inv10;
  reg [3:0] op1_04_in11;
  reg       op1_04_inv11;
  reg [3:0] op1_04_in12;
  reg       op1_04_inv12;
  reg [3:0] op1_04_in13;
  reg       op1_04_inv13;
  reg [3:0] op1_04_in14;
  reg       op1_04_inv14;
  reg [3:0] op1_04_in15;
  reg       op1_04_inv15;
  reg [3:0] op1_04_in16;
  reg       op1_04_inv16;
  reg [3:0] op1_04_in17;
  reg       op1_04_inv17;
  reg [3:0] op1_04_in18;
  reg       op1_04_inv18;
  reg [3:0] op1_04_in19;
  reg       op1_04_inv19;
  reg [3:0] op1_04_in20;
  reg       op1_04_inv20;
  reg [3:0] op1_04_in21;
  reg       op1_04_inv21;
  reg [3:0] op1_04_in22;
  reg       op1_04_inv22;
  reg [3:0] op1_04_in23;
  reg       op1_04_inv23;
  reg [3:0] op1_04_in24;
  reg       op1_04_inv24;
  reg [3:0] op1_04_in25;
  reg       op1_04_inv25;
  reg [3:0] op1_04_in26;
  reg       op1_04_inv26;
  reg [3:0] op1_04_in27;
  reg       op1_04_inv27;
  reg [3:0] op1_04_in28;
  reg       op1_04_inv28;
  reg [3:0] op1_04_in29;
  reg       op1_04_inv29;
  reg [3:0] op1_04_in30;
  reg       op1_04_inv30;
  reg [3:0] op1_04_in31;
  reg       op1_04_inv31;
  wire [8:0] op1_04_out;
  op1 op1_04(
    .data0_in(op1_04_in00),
    .inv0_in(op1_04_inv00),
    .data1_in(op1_04_in01),
    .inv1_in(op1_04_inv01),
    .data2_in(op1_04_in02),
    .inv2_in(op1_04_inv02),
    .data3_in(op1_04_in03),
    .inv3_in(op1_04_inv03),
    .data4_in(op1_04_in04),
    .inv4_in(op1_04_inv04),
    .data5_in(op1_04_in05),
    .inv5_in(op1_04_inv05),
    .data6_in(op1_04_in06),
    .inv6_in(op1_04_inv06),
    .data7_in(op1_04_in07),
    .inv7_in(op1_04_inv07),
    .data8_in(op1_04_in08),
    .inv8_in(op1_04_inv08),
    .data9_in(op1_04_in09),
    .inv9_in(op1_04_inv09),
    .data10_in(op1_04_in10),
    .inv10_in(op1_04_inv10),
    .data11_in(op1_04_in11),
    .inv11_in(op1_04_inv11),
    .data12_in(op1_04_in12),
    .inv12_in(op1_04_inv12),
    .data13_in(op1_04_in13),
    .inv13_in(op1_04_inv13),
    .data14_in(op1_04_in14),
    .inv14_in(op1_04_inv14),
    .data15_in(op1_04_in15),
    .inv15_in(op1_04_inv15),
    .data16_in(op1_04_in16),
    .inv16_in(op1_04_inv16),
    .data17_in(op1_04_in17),
    .inv17_in(op1_04_inv17),
    .data18_in(op1_04_in18),
    .inv18_in(op1_04_inv18),
    .data19_in(op1_04_in19),
    .inv19_in(op1_04_inv19),
    .data20_in(op1_04_in20),
    .inv20_in(op1_04_inv20),
    .data21_in(op1_04_in21),
    .inv21_in(op1_04_inv21),
    .data22_in(op1_04_in22),
    .inv22_in(op1_04_inv22),
    .data23_in(op1_04_in23),
    .inv23_in(op1_04_inv23),
    .data24_in(op1_04_in24),
    .inv24_in(op1_04_inv24),
    .data25_in(op1_04_in25),
    .inv25_in(op1_04_inv25),
    .data26_in(op1_04_in26),
    .inv26_in(op1_04_inv26),
    .data27_in(op1_04_in27),
    .inv27_in(op1_04_inv27),
    .data28_in(op1_04_in28),
    .inv28_in(op1_04_inv28),
    .data29_in(op1_04_in29),
    .inv29_in(op1_04_inv29),
    .data30_in(op1_04_in30),
    .inv30_in(op1_04_inv30),
    .data31_in(op1_04_in31),
    .inv31_in(op1_04_inv31),
    .data_out(op1_04_out));

  // 5 番目の OP1
  reg [3:0] op1_05_in00;
  reg       op1_05_inv00;
  reg [3:0] op1_05_in01;
  reg       op1_05_inv01;
  reg [3:0] op1_05_in02;
  reg       op1_05_inv02;
  reg [3:0] op1_05_in03;
  reg       op1_05_inv03;
  reg [3:0] op1_05_in04;
  reg       op1_05_inv04;
  reg [3:0] op1_05_in05;
  reg       op1_05_inv05;
  reg [3:0] op1_05_in06;
  reg       op1_05_inv06;
  reg [3:0] op1_05_in07;
  reg       op1_05_inv07;
  reg [3:0] op1_05_in08;
  reg       op1_05_inv08;
  reg [3:0] op1_05_in09;
  reg       op1_05_inv09;
  reg [3:0] op1_05_in10;
  reg       op1_05_inv10;
  reg [3:0] op1_05_in11;
  reg       op1_05_inv11;
  reg [3:0] op1_05_in12;
  reg       op1_05_inv12;
  reg [3:0] op1_05_in13;
  reg       op1_05_inv13;
  reg [3:0] op1_05_in14;
  reg       op1_05_inv14;
  reg [3:0] op1_05_in15;
  reg       op1_05_inv15;
  reg [3:0] op1_05_in16;
  reg       op1_05_inv16;
  reg [3:0] op1_05_in17;
  reg       op1_05_inv17;
  reg [3:0] op1_05_in18;
  reg       op1_05_inv18;
  reg [3:0] op1_05_in19;
  reg       op1_05_inv19;
  reg [3:0] op1_05_in20;
  reg       op1_05_inv20;
  reg [3:0] op1_05_in21;
  reg       op1_05_inv21;
  reg [3:0] op1_05_in22;
  reg       op1_05_inv22;
  reg [3:0] op1_05_in23;
  reg       op1_05_inv23;
  reg [3:0] op1_05_in24;
  reg       op1_05_inv24;
  reg [3:0] op1_05_in25;
  reg       op1_05_inv25;
  reg [3:0] op1_05_in26;
  reg       op1_05_inv26;
  reg [3:0] op1_05_in27;
  reg       op1_05_inv27;
  reg [3:0] op1_05_in28;
  reg       op1_05_inv28;
  reg [3:0] op1_05_in29;
  reg       op1_05_inv29;
  reg [3:0] op1_05_in30;
  reg       op1_05_inv30;
  reg [3:0] op1_05_in31;
  reg       op1_05_inv31;
  wire [8:0] op1_05_out;
  op1 op1_05(
    .data0_in(op1_05_in00),
    .inv0_in(op1_05_inv00),
    .data1_in(op1_05_in01),
    .inv1_in(op1_05_inv01),
    .data2_in(op1_05_in02),
    .inv2_in(op1_05_inv02),
    .data3_in(op1_05_in03),
    .inv3_in(op1_05_inv03),
    .data4_in(op1_05_in04),
    .inv4_in(op1_05_inv04),
    .data5_in(op1_05_in05),
    .inv5_in(op1_05_inv05),
    .data6_in(op1_05_in06),
    .inv6_in(op1_05_inv06),
    .data7_in(op1_05_in07),
    .inv7_in(op1_05_inv07),
    .data8_in(op1_05_in08),
    .inv8_in(op1_05_inv08),
    .data9_in(op1_05_in09),
    .inv9_in(op1_05_inv09),
    .data10_in(op1_05_in10),
    .inv10_in(op1_05_inv10),
    .data11_in(op1_05_in11),
    .inv11_in(op1_05_inv11),
    .data12_in(op1_05_in12),
    .inv12_in(op1_05_inv12),
    .data13_in(op1_05_in13),
    .inv13_in(op1_05_inv13),
    .data14_in(op1_05_in14),
    .inv14_in(op1_05_inv14),
    .data15_in(op1_05_in15),
    .inv15_in(op1_05_inv15),
    .data16_in(op1_05_in16),
    .inv16_in(op1_05_inv16),
    .data17_in(op1_05_in17),
    .inv17_in(op1_05_inv17),
    .data18_in(op1_05_in18),
    .inv18_in(op1_05_inv18),
    .data19_in(op1_05_in19),
    .inv19_in(op1_05_inv19),
    .data20_in(op1_05_in20),
    .inv20_in(op1_05_inv20),
    .data21_in(op1_05_in21),
    .inv21_in(op1_05_inv21),
    .data22_in(op1_05_in22),
    .inv22_in(op1_05_inv22),
    .data23_in(op1_05_in23),
    .inv23_in(op1_05_inv23),
    .data24_in(op1_05_in24),
    .inv24_in(op1_05_inv24),
    .data25_in(op1_05_in25),
    .inv25_in(op1_05_inv25),
    .data26_in(op1_05_in26),
    .inv26_in(op1_05_inv26),
    .data27_in(op1_05_in27),
    .inv27_in(op1_05_inv27),
    .data28_in(op1_05_in28),
    .inv28_in(op1_05_inv28),
    .data29_in(op1_05_in29),
    .inv29_in(op1_05_inv29),
    .data30_in(op1_05_in30),
    .inv30_in(op1_05_inv30),
    .data31_in(op1_05_in31),
    .inv31_in(op1_05_inv31),
    .data_out(op1_05_out));

  // 6 番目の OP1
  reg [3:0] op1_06_in00;
  reg       op1_06_inv00;
  reg [3:0] op1_06_in01;
  reg       op1_06_inv01;
  reg [3:0] op1_06_in02;
  reg       op1_06_inv02;
  reg [3:0] op1_06_in03;
  reg       op1_06_inv03;
  reg [3:0] op1_06_in04;
  reg       op1_06_inv04;
  reg [3:0] op1_06_in05;
  reg       op1_06_inv05;
  reg [3:0] op1_06_in06;
  reg       op1_06_inv06;
  reg [3:0] op1_06_in07;
  reg       op1_06_inv07;
  reg [3:0] op1_06_in08;
  reg       op1_06_inv08;
  reg [3:0] op1_06_in09;
  reg       op1_06_inv09;
  reg [3:0] op1_06_in10;
  reg       op1_06_inv10;
  reg [3:0] op1_06_in11;
  reg       op1_06_inv11;
  reg [3:0] op1_06_in12;
  reg       op1_06_inv12;
  reg [3:0] op1_06_in13;
  reg       op1_06_inv13;
  reg [3:0] op1_06_in14;
  reg       op1_06_inv14;
  reg [3:0] op1_06_in15;
  reg       op1_06_inv15;
  reg [3:0] op1_06_in16;
  reg       op1_06_inv16;
  reg [3:0] op1_06_in17;
  reg       op1_06_inv17;
  reg [3:0] op1_06_in18;
  reg       op1_06_inv18;
  reg [3:0] op1_06_in19;
  reg       op1_06_inv19;
  reg [3:0] op1_06_in20;
  reg       op1_06_inv20;
  reg [3:0] op1_06_in21;
  reg       op1_06_inv21;
  reg [3:0] op1_06_in22;
  reg       op1_06_inv22;
  reg [3:0] op1_06_in23;
  reg       op1_06_inv23;
  reg [3:0] op1_06_in24;
  reg       op1_06_inv24;
  reg [3:0] op1_06_in25;
  reg       op1_06_inv25;
  reg [3:0] op1_06_in26;
  reg       op1_06_inv26;
  reg [3:0] op1_06_in27;
  reg       op1_06_inv27;
  reg [3:0] op1_06_in28;
  reg       op1_06_inv28;
  reg [3:0] op1_06_in29;
  reg       op1_06_inv29;
  reg [3:0] op1_06_in30;
  reg       op1_06_inv30;
  reg [3:0] op1_06_in31;
  reg       op1_06_inv31;
  wire [8:0] op1_06_out;
  op1 op1_06(
    .data0_in(op1_06_in00),
    .inv0_in(op1_06_inv00),
    .data1_in(op1_06_in01),
    .inv1_in(op1_06_inv01),
    .data2_in(op1_06_in02),
    .inv2_in(op1_06_inv02),
    .data3_in(op1_06_in03),
    .inv3_in(op1_06_inv03),
    .data4_in(op1_06_in04),
    .inv4_in(op1_06_inv04),
    .data5_in(op1_06_in05),
    .inv5_in(op1_06_inv05),
    .data6_in(op1_06_in06),
    .inv6_in(op1_06_inv06),
    .data7_in(op1_06_in07),
    .inv7_in(op1_06_inv07),
    .data8_in(op1_06_in08),
    .inv8_in(op1_06_inv08),
    .data9_in(op1_06_in09),
    .inv9_in(op1_06_inv09),
    .data10_in(op1_06_in10),
    .inv10_in(op1_06_inv10),
    .data11_in(op1_06_in11),
    .inv11_in(op1_06_inv11),
    .data12_in(op1_06_in12),
    .inv12_in(op1_06_inv12),
    .data13_in(op1_06_in13),
    .inv13_in(op1_06_inv13),
    .data14_in(op1_06_in14),
    .inv14_in(op1_06_inv14),
    .data15_in(op1_06_in15),
    .inv15_in(op1_06_inv15),
    .data16_in(op1_06_in16),
    .inv16_in(op1_06_inv16),
    .data17_in(op1_06_in17),
    .inv17_in(op1_06_inv17),
    .data18_in(op1_06_in18),
    .inv18_in(op1_06_inv18),
    .data19_in(op1_06_in19),
    .inv19_in(op1_06_inv19),
    .data20_in(op1_06_in20),
    .inv20_in(op1_06_inv20),
    .data21_in(op1_06_in21),
    .inv21_in(op1_06_inv21),
    .data22_in(op1_06_in22),
    .inv22_in(op1_06_inv22),
    .data23_in(op1_06_in23),
    .inv23_in(op1_06_inv23),
    .data24_in(op1_06_in24),
    .inv24_in(op1_06_inv24),
    .data25_in(op1_06_in25),
    .inv25_in(op1_06_inv25),
    .data26_in(op1_06_in26),
    .inv26_in(op1_06_inv26),
    .data27_in(op1_06_in27),
    .inv27_in(op1_06_inv27),
    .data28_in(op1_06_in28),
    .inv28_in(op1_06_inv28),
    .data29_in(op1_06_in29),
    .inv29_in(op1_06_inv29),
    .data30_in(op1_06_in30),
    .inv30_in(op1_06_inv30),
    .data31_in(op1_06_in31),
    .inv31_in(op1_06_inv31),
    .data_out(op1_06_out));

  // 7 番目の OP1
  reg [3:0] op1_07_in00;
  reg       op1_07_inv00;
  reg [3:0] op1_07_in01;
  reg       op1_07_inv01;
  reg [3:0] op1_07_in02;
  reg       op1_07_inv02;
  reg [3:0] op1_07_in03;
  reg       op1_07_inv03;
  reg [3:0] op1_07_in04;
  reg       op1_07_inv04;
  reg [3:0] op1_07_in05;
  reg       op1_07_inv05;
  reg [3:0] op1_07_in06;
  reg       op1_07_inv06;
  reg [3:0] op1_07_in07;
  reg       op1_07_inv07;
  reg [3:0] op1_07_in08;
  reg       op1_07_inv08;
  reg [3:0] op1_07_in09;
  reg       op1_07_inv09;
  reg [3:0] op1_07_in10;
  reg       op1_07_inv10;
  reg [3:0] op1_07_in11;
  reg       op1_07_inv11;
  reg [3:0] op1_07_in12;
  reg       op1_07_inv12;
  reg [3:0] op1_07_in13;
  reg       op1_07_inv13;
  reg [3:0] op1_07_in14;
  reg       op1_07_inv14;
  reg [3:0] op1_07_in15;
  reg       op1_07_inv15;
  reg [3:0] op1_07_in16;
  reg       op1_07_inv16;
  reg [3:0] op1_07_in17;
  reg       op1_07_inv17;
  reg [3:0] op1_07_in18;
  reg       op1_07_inv18;
  reg [3:0] op1_07_in19;
  reg       op1_07_inv19;
  reg [3:0] op1_07_in20;
  reg       op1_07_inv20;
  reg [3:0] op1_07_in21;
  reg       op1_07_inv21;
  reg [3:0] op1_07_in22;
  reg       op1_07_inv22;
  reg [3:0] op1_07_in23;
  reg       op1_07_inv23;
  reg [3:0] op1_07_in24;
  reg       op1_07_inv24;
  reg [3:0] op1_07_in25;
  reg       op1_07_inv25;
  reg [3:0] op1_07_in26;
  reg       op1_07_inv26;
  reg [3:0] op1_07_in27;
  reg       op1_07_inv27;
  reg [3:0] op1_07_in28;
  reg       op1_07_inv28;
  reg [3:0] op1_07_in29;
  reg       op1_07_inv29;
  reg [3:0] op1_07_in30;
  reg       op1_07_inv30;
  reg [3:0] op1_07_in31;
  reg       op1_07_inv31;
  wire [8:0] op1_07_out;
  op1 op1_07(
    .data0_in(op1_07_in00),
    .inv0_in(op1_07_inv00),
    .data1_in(op1_07_in01),
    .inv1_in(op1_07_inv01),
    .data2_in(op1_07_in02),
    .inv2_in(op1_07_inv02),
    .data3_in(op1_07_in03),
    .inv3_in(op1_07_inv03),
    .data4_in(op1_07_in04),
    .inv4_in(op1_07_inv04),
    .data5_in(op1_07_in05),
    .inv5_in(op1_07_inv05),
    .data6_in(op1_07_in06),
    .inv6_in(op1_07_inv06),
    .data7_in(op1_07_in07),
    .inv7_in(op1_07_inv07),
    .data8_in(op1_07_in08),
    .inv8_in(op1_07_inv08),
    .data9_in(op1_07_in09),
    .inv9_in(op1_07_inv09),
    .data10_in(op1_07_in10),
    .inv10_in(op1_07_inv10),
    .data11_in(op1_07_in11),
    .inv11_in(op1_07_inv11),
    .data12_in(op1_07_in12),
    .inv12_in(op1_07_inv12),
    .data13_in(op1_07_in13),
    .inv13_in(op1_07_inv13),
    .data14_in(op1_07_in14),
    .inv14_in(op1_07_inv14),
    .data15_in(op1_07_in15),
    .inv15_in(op1_07_inv15),
    .data16_in(op1_07_in16),
    .inv16_in(op1_07_inv16),
    .data17_in(op1_07_in17),
    .inv17_in(op1_07_inv17),
    .data18_in(op1_07_in18),
    .inv18_in(op1_07_inv18),
    .data19_in(op1_07_in19),
    .inv19_in(op1_07_inv19),
    .data20_in(op1_07_in20),
    .inv20_in(op1_07_inv20),
    .data21_in(op1_07_in21),
    .inv21_in(op1_07_inv21),
    .data22_in(op1_07_in22),
    .inv22_in(op1_07_inv22),
    .data23_in(op1_07_in23),
    .inv23_in(op1_07_inv23),
    .data24_in(op1_07_in24),
    .inv24_in(op1_07_inv24),
    .data25_in(op1_07_in25),
    .inv25_in(op1_07_inv25),
    .data26_in(op1_07_in26),
    .inv26_in(op1_07_inv26),
    .data27_in(op1_07_in27),
    .inv27_in(op1_07_inv27),
    .data28_in(op1_07_in28),
    .inv28_in(op1_07_inv28),
    .data29_in(op1_07_in29),
    .inv29_in(op1_07_inv29),
    .data30_in(op1_07_in30),
    .inv30_in(op1_07_inv30),
    .data31_in(op1_07_in31),
    .inv31_in(op1_07_inv31),
    .data_out(op1_07_out));

  // 8 番目の OP1
  reg [3:0] op1_08_in00;
  reg       op1_08_inv00;
  reg [3:0] op1_08_in01;
  reg       op1_08_inv01;
  reg [3:0] op1_08_in02;
  reg       op1_08_inv02;
  reg [3:0] op1_08_in03;
  reg       op1_08_inv03;
  reg [3:0] op1_08_in04;
  reg       op1_08_inv04;
  reg [3:0] op1_08_in05;
  reg       op1_08_inv05;
  reg [3:0] op1_08_in06;
  reg       op1_08_inv06;
  reg [3:0] op1_08_in07;
  reg       op1_08_inv07;
  reg [3:0] op1_08_in08;
  reg       op1_08_inv08;
  reg [3:0] op1_08_in09;
  reg       op1_08_inv09;
  reg [3:0] op1_08_in10;
  reg       op1_08_inv10;
  reg [3:0] op1_08_in11;
  reg       op1_08_inv11;
  reg [3:0] op1_08_in12;
  reg       op1_08_inv12;
  reg [3:0] op1_08_in13;
  reg       op1_08_inv13;
  reg [3:0] op1_08_in14;
  reg       op1_08_inv14;
  reg [3:0] op1_08_in15;
  reg       op1_08_inv15;
  reg [3:0] op1_08_in16;
  reg       op1_08_inv16;
  reg [3:0] op1_08_in17;
  reg       op1_08_inv17;
  reg [3:0] op1_08_in18;
  reg       op1_08_inv18;
  reg [3:0] op1_08_in19;
  reg       op1_08_inv19;
  reg [3:0] op1_08_in20;
  reg       op1_08_inv20;
  reg [3:0] op1_08_in21;
  reg       op1_08_inv21;
  reg [3:0] op1_08_in22;
  reg       op1_08_inv22;
  reg [3:0] op1_08_in23;
  reg       op1_08_inv23;
  reg [3:0] op1_08_in24;
  reg       op1_08_inv24;
  reg [3:0] op1_08_in25;
  reg       op1_08_inv25;
  reg [3:0] op1_08_in26;
  reg       op1_08_inv26;
  reg [3:0] op1_08_in27;
  reg       op1_08_inv27;
  reg [3:0] op1_08_in28;
  reg       op1_08_inv28;
  reg [3:0] op1_08_in29;
  reg       op1_08_inv29;
  reg [3:0] op1_08_in30;
  reg       op1_08_inv30;
  reg [3:0] op1_08_in31;
  reg       op1_08_inv31;
  wire [8:0] op1_08_out;
  op1 op1_08(
    .data0_in(op1_08_in00),
    .inv0_in(op1_08_inv00),
    .data1_in(op1_08_in01),
    .inv1_in(op1_08_inv01),
    .data2_in(op1_08_in02),
    .inv2_in(op1_08_inv02),
    .data3_in(op1_08_in03),
    .inv3_in(op1_08_inv03),
    .data4_in(op1_08_in04),
    .inv4_in(op1_08_inv04),
    .data5_in(op1_08_in05),
    .inv5_in(op1_08_inv05),
    .data6_in(op1_08_in06),
    .inv6_in(op1_08_inv06),
    .data7_in(op1_08_in07),
    .inv7_in(op1_08_inv07),
    .data8_in(op1_08_in08),
    .inv8_in(op1_08_inv08),
    .data9_in(op1_08_in09),
    .inv9_in(op1_08_inv09),
    .data10_in(op1_08_in10),
    .inv10_in(op1_08_inv10),
    .data11_in(op1_08_in11),
    .inv11_in(op1_08_inv11),
    .data12_in(op1_08_in12),
    .inv12_in(op1_08_inv12),
    .data13_in(op1_08_in13),
    .inv13_in(op1_08_inv13),
    .data14_in(op1_08_in14),
    .inv14_in(op1_08_inv14),
    .data15_in(op1_08_in15),
    .inv15_in(op1_08_inv15),
    .data16_in(op1_08_in16),
    .inv16_in(op1_08_inv16),
    .data17_in(op1_08_in17),
    .inv17_in(op1_08_inv17),
    .data18_in(op1_08_in18),
    .inv18_in(op1_08_inv18),
    .data19_in(op1_08_in19),
    .inv19_in(op1_08_inv19),
    .data20_in(op1_08_in20),
    .inv20_in(op1_08_inv20),
    .data21_in(op1_08_in21),
    .inv21_in(op1_08_inv21),
    .data22_in(op1_08_in22),
    .inv22_in(op1_08_inv22),
    .data23_in(op1_08_in23),
    .inv23_in(op1_08_inv23),
    .data24_in(op1_08_in24),
    .inv24_in(op1_08_inv24),
    .data25_in(op1_08_in25),
    .inv25_in(op1_08_inv25),
    .data26_in(op1_08_in26),
    .inv26_in(op1_08_inv26),
    .data27_in(op1_08_in27),
    .inv27_in(op1_08_inv27),
    .data28_in(op1_08_in28),
    .inv28_in(op1_08_inv28),
    .data29_in(op1_08_in29),
    .inv29_in(op1_08_inv29),
    .data30_in(op1_08_in30),
    .inv30_in(op1_08_inv30),
    .data31_in(op1_08_in31),
    .inv31_in(op1_08_inv31),
    .data_out(op1_08_out));

  // 9 番目の OP1
  reg [3:0] op1_09_in00;
  reg       op1_09_inv00;
  reg [3:0] op1_09_in01;
  reg       op1_09_inv01;
  reg [3:0] op1_09_in02;
  reg       op1_09_inv02;
  reg [3:0] op1_09_in03;
  reg       op1_09_inv03;
  reg [3:0] op1_09_in04;
  reg       op1_09_inv04;
  reg [3:0] op1_09_in05;
  reg       op1_09_inv05;
  reg [3:0] op1_09_in06;
  reg       op1_09_inv06;
  reg [3:0] op1_09_in07;
  reg       op1_09_inv07;
  reg [3:0] op1_09_in08;
  reg       op1_09_inv08;
  reg [3:0] op1_09_in09;
  reg       op1_09_inv09;
  reg [3:0] op1_09_in10;
  reg       op1_09_inv10;
  reg [3:0] op1_09_in11;
  reg       op1_09_inv11;
  reg [3:0] op1_09_in12;
  reg       op1_09_inv12;
  reg [3:0] op1_09_in13;
  reg       op1_09_inv13;
  reg [3:0] op1_09_in14;
  reg       op1_09_inv14;
  reg [3:0] op1_09_in15;
  reg       op1_09_inv15;
  reg [3:0] op1_09_in16;
  reg       op1_09_inv16;
  reg [3:0] op1_09_in17;
  reg       op1_09_inv17;
  reg [3:0] op1_09_in18;
  reg       op1_09_inv18;
  reg [3:0] op1_09_in19;
  reg       op1_09_inv19;
  reg [3:0] op1_09_in20;
  reg       op1_09_inv20;
  reg [3:0] op1_09_in21;
  reg       op1_09_inv21;
  reg [3:0] op1_09_in22;
  reg       op1_09_inv22;
  reg [3:0] op1_09_in23;
  reg       op1_09_inv23;
  reg [3:0] op1_09_in24;
  reg       op1_09_inv24;
  reg [3:0] op1_09_in25;
  reg       op1_09_inv25;
  reg [3:0] op1_09_in26;
  reg       op1_09_inv26;
  reg [3:0] op1_09_in27;
  reg       op1_09_inv27;
  reg [3:0] op1_09_in28;
  reg       op1_09_inv28;
  reg [3:0] op1_09_in29;
  reg       op1_09_inv29;
  reg [3:0] op1_09_in30;
  reg       op1_09_inv30;
  reg [3:0] op1_09_in31;
  reg       op1_09_inv31;
  wire [8:0] op1_09_out;
  op1 op1_09(
    .data0_in(op1_09_in00),
    .inv0_in(op1_09_inv00),
    .data1_in(op1_09_in01),
    .inv1_in(op1_09_inv01),
    .data2_in(op1_09_in02),
    .inv2_in(op1_09_inv02),
    .data3_in(op1_09_in03),
    .inv3_in(op1_09_inv03),
    .data4_in(op1_09_in04),
    .inv4_in(op1_09_inv04),
    .data5_in(op1_09_in05),
    .inv5_in(op1_09_inv05),
    .data6_in(op1_09_in06),
    .inv6_in(op1_09_inv06),
    .data7_in(op1_09_in07),
    .inv7_in(op1_09_inv07),
    .data8_in(op1_09_in08),
    .inv8_in(op1_09_inv08),
    .data9_in(op1_09_in09),
    .inv9_in(op1_09_inv09),
    .data10_in(op1_09_in10),
    .inv10_in(op1_09_inv10),
    .data11_in(op1_09_in11),
    .inv11_in(op1_09_inv11),
    .data12_in(op1_09_in12),
    .inv12_in(op1_09_inv12),
    .data13_in(op1_09_in13),
    .inv13_in(op1_09_inv13),
    .data14_in(op1_09_in14),
    .inv14_in(op1_09_inv14),
    .data15_in(op1_09_in15),
    .inv15_in(op1_09_inv15),
    .data16_in(op1_09_in16),
    .inv16_in(op1_09_inv16),
    .data17_in(op1_09_in17),
    .inv17_in(op1_09_inv17),
    .data18_in(op1_09_in18),
    .inv18_in(op1_09_inv18),
    .data19_in(op1_09_in19),
    .inv19_in(op1_09_inv19),
    .data20_in(op1_09_in20),
    .inv20_in(op1_09_inv20),
    .data21_in(op1_09_in21),
    .inv21_in(op1_09_inv21),
    .data22_in(op1_09_in22),
    .inv22_in(op1_09_inv22),
    .data23_in(op1_09_in23),
    .inv23_in(op1_09_inv23),
    .data24_in(op1_09_in24),
    .inv24_in(op1_09_inv24),
    .data25_in(op1_09_in25),
    .inv25_in(op1_09_inv25),
    .data26_in(op1_09_in26),
    .inv26_in(op1_09_inv26),
    .data27_in(op1_09_in27),
    .inv27_in(op1_09_inv27),
    .data28_in(op1_09_in28),
    .inv28_in(op1_09_inv28),
    .data29_in(op1_09_in29),
    .inv29_in(op1_09_inv29),
    .data30_in(op1_09_in30),
    .inv30_in(op1_09_inv30),
    .data31_in(op1_09_in31),
    .inv31_in(op1_09_inv31),
    .data_out(op1_09_out));

  // 10 番目の OP1
  reg [3:0] op1_10_in00;
  reg       op1_10_inv00;
  reg [3:0] op1_10_in01;
  reg       op1_10_inv01;
  reg [3:0] op1_10_in02;
  reg       op1_10_inv02;
  reg [3:0] op1_10_in03;
  reg       op1_10_inv03;
  reg [3:0] op1_10_in04;
  reg       op1_10_inv04;
  reg [3:0] op1_10_in05;
  reg       op1_10_inv05;
  reg [3:0] op1_10_in06;
  reg       op1_10_inv06;
  reg [3:0] op1_10_in07;
  reg       op1_10_inv07;
  reg [3:0] op1_10_in08;
  reg       op1_10_inv08;
  reg [3:0] op1_10_in09;
  reg       op1_10_inv09;
  reg [3:0] op1_10_in10;
  reg       op1_10_inv10;
  reg [3:0] op1_10_in11;
  reg       op1_10_inv11;
  reg [3:0] op1_10_in12;
  reg       op1_10_inv12;
  reg [3:0] op1_10_in13;
  reg       op1_10_inv13;
  reg [3:0] op1_10_in14;
  reg       op1_10_inv14;
  reg [3:0] op1_10_in15;
  reg       op1_10_inv15;
  reg [3:0] op1_10_in16;
  reg       op1_10_inv16;
  reg [3:0] op1_10_in17;
  reg       op1_10_inv17;
  reg [3:0] op1_10_in18;
  reg       op1_10_inv18;
  reg [3:0] op1_10_in19;
  reg       op1_10_inv19;
  reg [3:0] op1_10_in20;
  reg       op1_10_inv20;
  reg [3:0] op1_10_in21;
  reg       op1_10_inv21;
  reg [3:0] op1_10_in22;
  reg       op1_10_inv22;
  reg [3:0] op1_10_in23;
  reg       op1_10_inv23;
  reg [3:0] op1_10_in24;
  reg       op1_10_inv24;
  reg [3:0] op1_10_in25;
  reg       op1_10_inv25;
  reg [3:0] op1_10_in26;
  reg       op1_10_inv26;
  reg [3:0] op1_10_in27;
  reg       op1_10_inv27;
  reg [3:0] op1_10_in28;
  reg       op1_10_inv28;
  reg [3:0] op1_10_in29;
  reg       op1_10_inv29;
  reg [3:0] op1_10_in30;
  reg       op1_10_inv30;
  reg [3:0] op1_10_in31;
  reg       op1_10_inv31;
  wire [8:0] op1_10_out;
  op1 op1_10(
    .data0_in(op1_10_in00),
    .inv0_in(op1_10_inv00),
    .data1_in(op1_10_in01),
    .inv1_in(op1_10_inv01),
    .data2_in(op1_10_in02),
    .inv2_in(op1_10_inv02),
    .data3_in(op1_10_in03),
    .inv3_in(op1_10_inv03),
    .data4_in(op1_10_in04),
    .inv4_in(op1_10_inv04),
    .data5_in(op1_10_in05),
    .inv5_in(op1_10_inv05),
    .data6_in(op1_10_in06),
    .inv6_in(op1_10_inv06),
    .data7_in(op1_10_in07),
    .inv7_in(op1_10_inv07),
    .data8_in(op1_10_in08),
    .inv8_in(op1_10_inv08),
    .data9_in(op1_10_in09),
    .inv9_in(op1_10_inv09),
    .data10_in(op1_10_in10),
    .inv10_in(op1_10_inv10),
    .data11_in(op1_10_in11),
    .inv11_in(op1_10_inv11),
    .data12_in(op1_10_in12),
    .inv12_in(op1_10_inv12),
    .data13_in(op1_10_in13),
    .inv13_in(op1_10_inv13),
    .data14_in(op1_10_in14),
    .inv14_in(op1_10_inv14),
    .data15_in(op1_10_in15),
    .inv15_in(op1_10_inv15),
    .data16_in(op1_10_in16),
    .inv16_in(op1_10_inv16),
    .data17_in(op1_10_in17),
    .inv17_in(op1_10_inv17),
    .data18_in(op1_10_in18),
    .inv18_in(op1_10_inv18),
    .data19_in(op1_10_in19),
    .inv19_in(op1_10_inv19),
    .data20_in(op1_10_in20),
    .inv20_in(op1_10_inv20),
    .data21_in(op1_10_in21),
    .inv21_in(op1_10_inv21),
    .data22_in(op1_10_in22),
    .inv22_in(op1_10_inv22),
    .data23_in(op1_10_in23),
    .inv23_in(op1_10_inv23),
    .data24_in(op1_10_in24),
    .inv24_in(op1_10_inv24),
    .data25_in(op1_10_in25),
    .inv25_in(op1_10_inv25),
    .data26_in(op1_10_in26),
    .inv26_in(op1_10_inv26),
    .data27_in(op1_10_in27),
    .inv27_in(op1_10_inv27),
    .data28_in(op1_10_in28),
    .inv28_in(op1_10_inv28),
    .data29_in(op1_10_in29),
    .inv29_in(op1_10_inv29),
    .data30_in(op1_10_in30),
    .inv30_in(op1_10_inv30),
    .data31_in(op1_10_in31),
    .inv31_in(op1_10_inv31),
    .data_out(op1_10_out));

  // 11 番目の OP1
  reg [3:0] op1_11_in00;
  reg       op1_11_inv00;
  reg [3:0] op1_11_in01;
  reg       op1_11_inv01;
  reg [3:0] op1_11_in02;
  reg       op1_11_inv02;
  reg [3:0] op1_11_in03;
  reg       op1_11_inv03;
  reg [3:0] op1_11_in04;
  reg       op1_11_inv04;
  reg [3:0] op1_11_in05;
  reg       op1_11_inv05;
  reg [3:0] op1_11_in06;
  reg       op1_11_inv06;
  reg [3:0] op1_11_in07;
  reg       op1_11_inv07;
  reg [3:0] op1_11_in08;
  reg       op1_11_inv08;
  reg [3:0] op1_11_in09;
  reg       op1_11_inv09;
  reg [3:0] op1_11_in10;
  reg       op1_11_inv10;
  reg [3:0] op1_11_in11;
  reg       op1_11_inv11;
  reg [3:0] op1_11_in12;
  reg       op1_11_inv12;
  reg [3:0] op1_11_in13;
  reg       op1_11_inv13;
  reg [3:0] op1_11_in14;
  reg       op1_11_inv14;
  reg [3:0] op1_11_in15;
  reg       op1_11_inv15;
  reg [3:0] op1_11_in16;
  reg       op1_11_inv16;
  reg [3:0] op1_11_in17;
  reg       op1_11_inv17;
  reg [3:0] op1_11_in18;
  reg       op1_11_inv18;
  reg [3:0] op1_11_in19;
  reg       op1_11_inv19;
  reg [3:0] op1_11_in20;
  reg       op1_11_inv20;
  reg [3:0] op1_11_in21;
  reg       op1_11_inv21;
  reg [3:0] op1_11_in22;
  reg       op1_11_inv22;
  reg [3:0] op1_11_in23;
  reg       op1_11_inv23;
  reg [3:0] op1_11_in24;
  reg       op1_11_inv24;
  reg [3:0] op1_11_in25;
  reg       op1_11_inv25;
  reg [3:0] op1_11_in26;
  reg       op1_11_inv26;
  reg [3:0] op1_11_in27;
  reg       op1_11_inv27;
  reg [3:0] op1_11_in28;
  reg       op1_11_inv28;
  reg [3:0] op1_11_in29;
  reg       op1_11_inv29;
  reg [3:0] op1_11_in30;
  reg       op1_11_inv30;
  reg [3:0] op1_11_in31;
  reg       op1_11_inv31;
  wire [8:0] op1_11_out;
  op1 op1_11(
    .data0_in(op1_11_in00),
    .inv0_in(op1_11_inv00),
    .data1_in(op1_11_in01),
    .inv1_in(op1_11_inv01),
    .data2_in(op1_11_in02),
    .inv2_in(op1_11_inv02),
    .data3_in(op1_11_in03),
    .inv3_in(op1_11_inv03),
    .data4_in(op1_11_in04),
    .inv4_in(op1_11_inv04),
    .data5_in(op1_11_in05),
    .inv5_in(op1_11_inv05),
    .data6_in(op1_11_in06),
    .inv6_in(op1_11_inv06),
    .data7_in(op1_11_in07),
    .inv7_in(op1_11_inv07),
    .data8_in(op1_11_in08),
    .inv8_in(op1_11_inv08),
    .data9_in(op1_11_in09),
    .inv9_in(op1_11_inv09),
    .data10_in(op1_11_in10),
    .inv10_in(op1_11_inv10),
    .data11_in(op1_11_in11),
    .inv11_in(op1_11_inv11),
    .data12_in(op1_11_in12),
    .inv12_in(op1_11_inv12),
    .data13_in(op1_11_in13),
    .inv13_in(op1_11_inv13),
    .data14_in(op1_11_in14),
    .inv14_in(op1_11_inv14),
    .data15_in(op1_11_in15),
    .inv15_in(op1_11_inv15),
    .data16_in(op1_11_in16),
    .inv16_in(op1_11_inv16),
    .data17_in(op1_11_in17),
    .inv17_in(op1_11_inv17),
    .data18_in(op1_11_in18),
    .inv18_in(op1_11_inv18),
    .data19_in(op1_11_in19),
    .inv19_in(op1_11_inv19),
    .data20_in(op1_11_in20),
    .inv20_in(op1_11_inv20),
    .data21_in(op1_11_in21),
    .inv21_in(op1_11_inv21),
    .data22_in(op1_11_in22),
    .inv22_in(op1_11_inv22),
    .data23_in(op1_11_in23),
    .inv23_in(op1_11_inv23),
    .data24_in(op1_11_in24),
    .inv24_in(op1_11_inv24),
    .data25_in(op1_11_in25),
    .inv25_in(op1_11_inv25),
    .data26_in(op1_11_in26),
    .inv26_in(op1_11_inv26),
    .data27_in(op1_11_in27),
    .inv27_in(op1_11_inv27),
    .data28_in(op1_11_in28),
    .inv28_in(op1_11_inv28),
    .data29_in(op1_11_in29),
    .inv29_in(op1_11_inv29),
    .data30_in(op1_11_in30),
    .inv30_in(op1_11_inv30),
    .data31_in(op1_11_in31),
    .inv31_in(op1_11_inv31),
    .data_out(op1_11_out));

  // 12 番目の OP1
  reg [3:0] op1_12_in00;
  reg       op1_12_inv00;
  reg [3:0] op1_12_in01;
  reg       op1_12_inv01;
  reg [3:0] op1_12_in02;
  reg       op1_12_inv02;
  reg [3:0] op1_12_in03;
  reg       op1_12_inv03;
  reg [3:0] op1_12_in04;
  reg       op1_12_inv04;
  reg [3:0] op1_12_in05;
  reg       op1_12_inv05;
  reg [3:0] op1_12_in06;
  reg       op1_12_inv06;
  reg [3:0] op1_12_in07;
  reg       op1_12_inv07;
  reg [3:0] op1_12_in08;
  reg       op1_12_inv08;
  reg [3:0] op1_12_in09;
  reg       op1_12_inv09;
  reg [3:0] op1_12_in10;
  reg       op1_12_inv10;
  reg [3:0] op1_12_in11;
  reg       op1_12_inv11;
  reg [3:0] op1_12_in12;
  reg       op1_12_inv12;
  reg [3:0] op1_12_in13;
  reg       op1_12_inv13;
  reg [3:0] op1_12_in14;
  reg       op1_12_inv14;
  reg [3:0] op1_12_in15;
  reg       op1_12_inv15;
  reg [3:0] op1_12_in16;
  reg       op1_12_inv16;
  reg [3:0] op1_12_in17;
  reg       op1_12_inv17;
  reg [3:0] op1_12_in18;
  reg       op1_12_inv18;
  reg [3:0] op1_12_in19;
  reg       op1_12_inv19;
  reg [3:0] op1_12_in20;
  reg       op1_12_inv20;
  reg [3:0] op1_12_in21;
  reg       op1_12_inv21;
  reg [3:0] op1_12_in22;
  reg       op1_12_inv22;
  reg [3:0] op1_12_in23;
  reg       op1_12_inv23;
  reg [3:0] op1_12_in24;
  reg       op1_12_inv24;
  reg [3:0] op1_12_in25;
  reg       op1_12_inv25;
  reg [3:0] op1_12_in26;
  reg       op1_12_inv26;
  reg [3:0] op1_12_in27;
  reg       op1_12_inv27;
  reg [3:0] op1_12_in28;
  reg       op1_12_inv28;
  reg [3:0] op1_12_in29;
  reg       op1_12_inv29;
  reg [3:0] op1_12_in30;
  reg       op1_12_inv30;
  reg [3:0] op1_12_in31;
  reg       op1_12_inv31;
  wire [8:0] op1_12_out;
  op1 op1_12(
    .data0_in(op1_12_in00),
    .inv0_in(op1_12_inv00),
    .data1_in(op1_12_in01),
    .inv1_in(op1_12_inv01),
    .data2_in(op1_12_in02),
    .inv2_in(op1_12_inv02),
    .data3_in(op1_12_in03),
    .inv3_in(op1_12_inv03),
    .data4_in(op1_12_in04),
    .inv4_in(op1_12_inv04),
    .data5_in(op1_12_in05),
    .inv5_in(op1_12_inv05),
    .data6_in(op1_12_in06),
    .inv6_in(op1_12_inv06),
    .data7_in(op1_12_in07),
    .inv7_in(op1_12_inv07),
    .data8_in(op1_12_in08),
    .inv8_in(op1_12_inv08),
    .data9_in(op1_12_in09),
    .inv9_in(op1_12_inv09),
    .data10_in(op1_12_in10),
    .inv10_in(op1_12_inv10),
    .data11_in(op1_12_in11),
    .inv11_in(op1_12_inv11),
    .data12_in(op1_12_in12),
    .inv12_in(op1_12_inv12),
    .data13_in(op1_12_in13),
    .inv13_in(op1_12_inv13),
    .data14_in(op1_12_in14),
    .inv14_in(op1_12_inv14),
    .data15_in(op1_12_in15),
    .inv15_in(op1_12_inv15),
    .data16_in(op1_12_in16),
    .inv16_in(op1_12_inv16),
    .data17_in(op1_12_in17),
    .inv17_in(op1_12_inv17),
    .data18_in(op1_12_in18),
    .inv18_in(op1_12_inv18),
    .data19_in(op1_12_in19),
    .inv19_in(op1_12_inv19),
    .data20_in(op1_12_in20),
    .inv20_in(op1_12_inv20),
    .data21_in(op1_12_in21),
    .inv21_in(op1_12_inv21),
    .data22_in(op1_12_in22),
    .inv22_in(op1_12_inv22),
    .data23_in(op1_12_in23),
    .inv23_in(op1_12_inv23),
    .data24_in(op1_12_in24),
    .inv24_in(op1_12_inv24),
    .data25_in(op1_12_in25),
    .inv25_in(op1_12_inv25),
    .data26_in(op1_12_in26),
    .inv26_in(op1_12_inv26),
    .data27_in(op1_12_in27),
    .inv27_in(op1_12_inv27),
    .data28_in(op1_12_in28),
    .inv28_in(op1_12_inv28),
    .data29_in(op1_12_in29),
    .inv29_in(op1_12_inv29),
    .data30_in(op1_12_in30),
    .inv30_in(op1_12_inv30),
    .data31_in(op1_12_in31),
    .inv31_in(op1_12_inv31),
    .data_out(op1_12_out));

  // 13 番目の OP1
  reg [3:0] op1_13_in00;
  reg       op1_13_inv00;
  reg [3:0] op1_13_in01;
  reg       op1_13_inv01;
  reg [3:0] op1_13_in02;
  reg       op1_13_inv02;
  reg [3:0] op1_13_in03;
  reg       op1_13_inv03;
  reg [3:0] op1_13_in04;
  reg       op1_13_inv04;
  reg [3:0] op1_13_in05;
  reg       op1_13_inv05;
  reg [3:0] op1_13_in06;
  reg       op1_13_inv06;
  reg [3:0] op1_13_in07;
  reg       op1_13_inv07;
  reg [3:0] op1_13_in08;
  reg       op1_13_inv08;
  reg [3:0] op1_13_in09;
  reg       op1_13_inv09;
  reg [3:0] op1_13_in10;
  reg       op1_13_inv10;
  reg [3:0] op1_13_in11;
  reg       op1_13_inv11;
  reg [3:0] op1_13_in12;
  reg       op1_13_inv12;
  reg [3:0] op1_13_in13;
  reg       op1_13_inv13;
  reg [3:0] op1_13_in14;
  reg       op1_13_inv14;
  reg [3:0] op1_13_in15;
  reg       op1_13_inv15;
  reg [3:0] op1_13_in16;
  reg       op1_13_inv16;
  reg [3:0] op1_13_in17;
  reg       op1_13_inv17;
  reg [3:0] op1_13_in18;
  reg       op1_13_inv18;
  reg [3:0] op1_13_in19;
  reg       op1_13_inv19;
  reg [3:0] op1_13_in20;
  reg       op1_13_inv20;
  reg [3:0] op1_13_in21;
  reg       op1_13_inv21;
  reg [3:0] op1_13_in22;
  reg       op1_13_inv22;
  reg [3:0] op1_13_in23;
  reg       op1_13_inv23;
  reg [3:0] op1_13_in24;
  reg       op1_13_inv24;
  reg [3:0] op1_13_in25;
  reg       op1_13_inv25;
  reg [3:0] op1_13_in26;
  reg       op1_13_inv26;
  reg [3:0] op1_13_in27;
  reg       op1_13_inv27;
  reg [3:0] op1_13_in28;
  reg       op1_13_inv28;
  reg [3:0] op1_13_in29;
  reg       op1_13_inv29;
  reg [3:0] op1_13_in30;
  reg       op1_13_inv30;
  reg [3:0] op1_13_in31;
  reg       op1_13_inv31;
  wire [8:0] op1_13_out;
  op1 op1_13(
    .data0_in(op1_13_in00),
    .inv0_in(op1_13_inv00),
    .data1_in(op1_13_in01),
    .inv1_in(op1_13_inv01),
    .data2_in(op1_13_in02),
    .inv2_in(op1_13_inv02),
    .data3_in(op1_13_in03),
    .inv3_in(op1_13_inv03),
    .data4_in(op1_13_in04),
    .inv4_in(op1_13_inv04),
    .data5_in(op1_13_in05),
    .inv5_in(op1_13_inv05),
    .data6_in(op1_13_in06),
    .inv6_in(op1_13_inv06),
    .data7_in(op1_13_in07),
    .inv7_in(op1_13_inv07),
    .data8_in(op1_13_in08),
    .inv8_in(op1_13_inv08),
    .data9_in(op1_13_in09),
    .inv9_in(op1_13_inv09),
    .data10_in(op1_13_in10),
    .inv10_in(op1_13_inv10),
    .data11_in(op1_13_in11),
    .inv11_in(op1_13_inv11),
    .data12_in(op1_13_in12),
    .inv12_in(op1_13_inv12),
    .data13_in(op1_13_in13),
    .inv13_in(op1_13_inv13),
    .data14_in(op1_13_in14),
    .inv14_in(op1_13_inv14),
    .data15_in(op1_13_in15),
    .inv15_in(op1_13_inv15),
    .data16_in(op1_13_in16),
    .inv16_in(op1_13_inv16),
    .data17_in(op1_13_in17),
    .inv17_in(op1_13_inv17),
    .data18_in(op1_13_in18),
    .inv18_in(op1_13_inv18),
    .data19_in(op1_13_in19),
    .inv19_in(op1_13_inv19),
    .data20_in(op1_13_in20),
    .inv20_in(op1_13_inv20),
    .data21_in(op1_13_in21),
    .inv21_in(op1_13_inv21),
    .data22_in(op1_13_in22),
    .inv22_in(op1_13_inv22),
    .data23_in(op1_13_in23),
    .inv23_in(op1_13_inv23),
    .data24_in(op1_13_in24),
    .inv24_in(op1_13_inv24),
    .data25_in(op1_13_in25),
    .inv25_in(op1_13_inv25),
    .data26_in(op1_13_in26),
    .inv26_in(op1_13_inv26),
    .data27_in(op1_13_in27),
    .inv27_in(op1_13_inv27),
    .data28_in(op1_13_in28),
    .inv28_in(op1_13_inv28),
    .data29_in(op1_13_in29),
    .inv29_in(op1_13_inv29),
    .data30_in(op1_13_in30),
    .inv30_in(op1_13_inv30),
    .data31_in(op1_13_in31),
    .inv31_in(op1_13_inv31),
    .data_out(op1_13_out));

  // 14 番目の OP1
  reg [3:0] op1_14_in00;
  reg       op1_14_inv00;
  reg [3:0] op1_14_in01;
  reg       op1_14_inv01;
  reg [3:0] op1_14_in02;
  reg       op1_14_inv02;
  reg [3:0] op1_14_in03;
  reg       op1_14_inv03;
  reg [3:0] op1_14_in04;
  reg       op1_14_inv04;
  reg [3:0] op1_14_in05;
  reg       op1_14_inv05;
  reg [3:0] op1_14_in06;
  reg       op1_14_inv06;
  reg [3:0] op1_14_in07;
  reg       op1_14_inv07;
  reg [3:0] op1_14_in08;
  reg       op1_14_inv08;
  reg [3:0] op1_14_in09;
  reg       op1_14_inv09;
  reg [3:0] op1_14_in10;
  reg       op1_14_inv10;
  reg [3:0] op1_14_in11;
  reg       op1_14_inv11;
  reg [3:0] op1_14_in12;
  reg       op1_14_inv12;
  reg [3:0] op1_14_in13;
  reg       op1_14_inv13;
  reg [3:0] op1_14_in14;
  reg       op1_14_inv14;
  reg [3:0] op1_14_in15;
  reg       op1_14_inv15;
  reg [3:0] op1_14_in16;
  reg       op1_14_inv16;
  reg [3:0] op1_14_in17;
  reg       op1_14_inv17;
  reg [3:0] op1_14_in18;
  reg       op1_14_inv18;
  reg [3:0] op1_14_in19;
  reg       op1_14_inv19;
  reg [3:0] op1_14_in20;
  reg       op1_14_inv20;
  reg [3:0] op1_14_in21;
  reg       op1_14_inv21;
  reg [3:0] op1_14_in22;
  reg       op1_14_inv22;
  reg [3:0] op1_14_in23;
  reg       op1_14_inv23;
  reg [3:0] op1_14_in24;
  reg       op1_14_inv24;
  reg [3:0] op1_14_in25;
  reg       op1_14_inv25;
  reg [3:0] op1_14_in26;
  reg       op1_14_inv26;
  reg [3:0] op1_14_in27;
  reg       op1_14_inv27;
  reg [3:0] op1_14_in28;
  reg       op1_14_inv28;
  reg [3:0] op1_14_in29;
  reg       op1_14_inv29;
  reg [3:0] op1_14_in30;
  reg       op1_14_inv30;
  reg [3:0] op1_14_in31;
  reg       op1_14_inv31;
  wire [8:0] op1_14_out;
  op1 op1_14(
    .data0_in(op1_14_in00),
    .inv0_in(op1_14_inv00),
    .data1_in(op1_14_in01),
    .inv1_in(op1_14_inv01),
    .data2_in(op1_14_in02),
    .inv2_in(op1_14_inv02),
    .data3_in(op1_14_in03),
    .inv3_in(op1_14_inv03),
    .data4_in(op1_14_in04),
    .inv4_in(op1_14_inv04),
    .data5_in(op1_14_in05),
    .inv5_in(op1_14_inv05),
    .data6_in(op1_14_in06),
    .inv6_in(op1_14_inv06),
    .data7_in(op1_14_in07),
    .inv7_in(op1_14_inv07),
    .data8_in(op1_14_in08),
    .inv8_in(op1_14_inv08),
    .data9_in(op1_14_in09),
    .inv9_in(op1_14_inv09),
    .data10_in(op1_14_in10),
    .inv10_in(op1_14_inv10),
    .data11_in(op1_14_in11),
    .inv11_in(op1_14_inv11),
    .data12_in(op1_14_in12),
    .inv12_in(op1_14_inv12),
    .data13_in(op1_14_in13),
    .inv13_in(op1_14_inv13),
    .data14_in(op1_14_in14),
    .inv14_in(op1_14_inv14),
    .data15_in(op1_14_in15),
    .inv15_in(op1_14_inv15),
    .data16_in(op1_14_in16),
    .inv16_in(op1_14_inv16),
    .data17_in(op1_14_in17),
    .inv17_in(op1_14_inv17),
    .data18_in(op1_14_in18),
    .inv18_in(op1_14_inv18),
    .data19_in(op1_14_in19),
    .inv19_in(op1_14_inv19),
    .data20_in(op1_14_in20),
    .inv20_in(op1_14_inv20),
    .data21_in(op1_14_in21),
    .inv21_in(op1_14_inv21),
    .data22_in(op1_14_in22),
    .inv22_in(op1_14_inv22),
    .data23_in(op1_14_in23),
    .inv23_in(op1_14_inv23),
    .data24_in(op1_14_in24),
    .inv24_in(op1_14_inv24),
    .data25_in(op1_14_in25),
    .inv25_in(op1_14_inv25),
    .data26_in(op1_14_in26),
    .inv26_in(op1_14_inv26),
    .data27_in(op1_14_in27),
    .inv27_in(op1_14_inv27),
    .data28_in(op1_14_in28),
    .inv28_in(op1_14_inv28),
    .data29_in(op1_14_in29),
    .inv29_in(op1_14_inv29),
    .data30_in(op1_14_in30),
    .inv30_in(op1_14_inv30),
    .data31_in(op1_14_in31),
    .inv31_in(op1_14_inv31),
    .data_out(op1_14_out));

  // 15 番目の OP1
  reg [3:0] op1_15_in00;
  reg       op1_15_inv00;
  reg [3:0] op1_15_in01;
  reg       op1_15_inv01;
  reg [3:0] op1_15_in02;
  reg       op1_15_inv02;
  reg [3:0] op1_15_in03;
  reg       op1_15_inv03;
  reg [3:0] op1_15_in04;
  reg       op1_15_inv04;
  reg [3:0] op1_15_in05;
  reg       op1_15_inv05;
  reg [3:0] op1_15_in06;
  reg       op1_15_inv06;
  reg [3:0] op1_15_in07;
  reg       op1_15_inv07;
  reg [3:0] op1_15_in08;
  reg       op1_15_inv08;
  reg [3:0] op1_15_in09;
  reg       op1_15_inv09;
  reg [3:0] op1_15_in10;
  reg       op1_15_inv10;
  reg [3:0] op1_15_in11;
  reg       op1_15_inv11;
  reg [3:0] op1_15_in12;
  reg       op1_15_inv12;
  reg [3:0] op1_15_in13;
  reg       op1_15_inv13;
  reg [3:0] op1_15_in14;
  reg       op1_15_inv14;
  reg [3:0] op1_15_in15;
  reg       op1_15_inv15;
  reg [3:0] op1_15_in16;
  reg       op1_15_inv16;
  reg [3:0] op1_15_in17;
  reg       op1_15_inv17;
  reg [3:0] op1_15_in18;
  reg       op1_15_inv18;
  reg [3:0] op1_15_in19;
  reg       op1_15_inv19;
  reg [3:0] op1_15_in20;
  reg       op1_15_inv20;
  reg [3:0] op1_15_in21;
  reg       op1_15_inv21;
  reg [3:0] op1_15_in22;
  reg       op1_15_inv22;
  reg [3:0] op1_15_in23;
  reg       op1_15_inv23;
  reg [3:0] op1_15_in24;
  reg       op1_15_inv24;
  reg [3:0] op1_15_in25;
  reg       op1_15_inv25;
  reg [3:0] op1_15_in26;
  reg       op1_15_inv26;
  reg [3:0] op1_15_in27;
  reg       op1_15_inv27;
  reg [3:0] op1_15_in28;
  reg       op1_15_inv28;
  reg [3:0] op1_15_in29;
  reg       op1_15_inv29;
  reg [3:0] op1_15_in30;
  reg       op1_15_inv30;
  reg [3:0] op1_15_in31;
  reg       op1_15_inv31;
  wire [8:0] op1_15_out;
  op1 op1_15(
    .data0_in(op1_15_in00),
    .inv0_in(op1_15_inv00),
    .data1_in(op1_15_in01),
    .inv1_in(op1_15_inv01),
    .data2_in(op1_15_in02),
    .inv2_in(op1_15_inv02),
    .data3_in(op1_15_in03),
    .inv3_in(op1_15_inv03),
    .data4_in(op1_15_in04),
    .inv4_in(op1_15_inv04),
    .data5_in(op1_15_in05),
    .inv5_in(op1_15_inv05),
    .data6_in(op1_15_in06),
    .inv6_in(op1_15_inv06),
    .data7_in(op1_15_in07),
    .inv7_in(op1_15_inv07),
    .data8_in(op1_15_in08),
    .inv8_in(op1_15_inv08),
    .data9_in(op1_15_in09),
    .inv9_in(op1_15_inv09),
    .data10_in(op1_15_in10),
    .inv10_in(op1_15_inv10),
    .data11_in(op1_15_in11),
    .inv11_in(op1_15_inv11),
    .data12_in(op1_15_in12),
    .inv12_in(op1_15_inv12),
    .data13_in(op1_15_in13),
    .inv13_in(op1_15_inv13),
    .data14_in(op1_15_in14),
    .inv14_in(op1_15_inv14),
    .data15_in(op1_15_in15),
    .inv15_in(op1_15_inv15),
    .data16_in(op1_15_in16),
    .inv16_in(op1_15_inv16),
    .data17_in(op1_15_in17),
    .inv17_in(op1_15_inv17),
    .data18_in(op1_15_in18),
    .inv18_in(op1_15_inv18),
    .data19_in(op1_15_in19),
    .inv19_in(op1_15_inv19),
    .data20_in(op1_15_in20),
    .inv20_in(op1_15_inv20),
    .data21_in(op1_15_in21),
    .inv21_in(op1_15_inv21),
    .data22_in(op1_15_in22),
    .inv22_in(op1_15_inv22),
    .data23_in(op1_15_in23),
    .inv23_in(op1_15_inv23),
    .data24_in(op1_15_in24),
    .inv24_in(op1_15_inv24),
    .data25_in(op1_15_in25),
    .inv25_in(op1_15_inv25),
    .data26_in(op1_15_in26),
    .inv26_in(op1_15_inv26),
    .data27_in(op1_15_in27),
    .inv27_in(op1_15_inv27),
    .data28_in(op1_15_in28),
    .inv28_in(op1_15_inv28),
    .data29_in(op1_15_in29),
    .inv29_in(op1_15_inv29),
    .data30_in(op1_15_in30),
    .inv30_in(op1_15_inv30),
    .data31_in(op1_15_in31),
    .inv31_in(op1_15_inv31),
    .data_out(op1_15_out));

  // 0 番目の OP2
  reg [8:0] op2_00_in00;
  reg [8:0] op2_00_in01;
  reg [8:0] op2_00_in02;
  reg [8:0] op2_00_in03;
  reg [8:0] op2_00_in04;
  reg [8:0] op2_00_in05;
  reg [8:0] op2_00_in06;
  reg [8:0] op2_00_in07;
  reg [8:0] op2_00_in08;
  reg [8:0] op2_00_in09;
  reg [8:0] op2_00_in10;
  reg [8:0] op2_00_in11;
  reg [8:0] op2_00_in12;
  reg [8:0] op2_00_in13;
  reg [8:0] op2_00_in14;
  reg [8:0] op2_00_in15;
  reg [8:0] op2_00_in16;
  reg [8:0] op2_00_in17;
  reg [8:0] op2_00_in18;
  reg [8:0] op2_00_in19;
  reg [8:0] op2_00_in20;
  reg [8:0] op2_00_in21;
  reg [8:0] op2_00_in22;
  reg [8:0] op2_00_in23;
  reg [8:0] op2_00_in24;
  reg [8:0] op2_00_in25;
  reg [8:0] op2_00_in26;
  reg [8:0] op2_00_in27;
  reg [8:0] op2_00_in28;
  reg [8:0] op2_00_in29;
  reg [8:0] op2_00_in30;
  reg [8:0] op2_00_bias;
  wire [8:0] op2_00_out;
  op2 op2_00(
    .data0_in(op2_00_in00),
    .data1_in(op2_00_in01),
    .data2_in(op2_00_in02),
    .data3_in(op2_00_in03),
    .data4_in(op2_00_in04),
    .data5_in(op2_00_in05),
    .data6_in(op2_00_in06),
    .data7_in(op2_00_in07),
    .data8_in(op2_00_in08),
    .data9_in(op2_00_in09),
    .data10_in(op2_00_in10),
    .data11_in(op2_00_in11),
    .data12_in(op2_00_in12),
    .data13_in(op2_00_in13),
    .data14_in(op2_00_in14),
    .data15_in(op2_00_in15),
    .data16_in(op2_00_in16),
    .data17_in(op2_00_in17),
    .data18_in(op2_00_in18),
    .data19_in(op2_00_in19),
    .data20_in(op2_00_in20),
    .data21_in(op2_00_in21),
    .data22_in(op2_00_in22),
    .data23_in(op2_00_in23),
    .data24_in(op2_00_in24),
    .data25_in(op2_00_in25),
    .data26_in(op2_00_in26),
    .data27_in(op2_00_in27),
    .data28_in(op2_00_in28),
    .data29_in(op2_00_in29),
    .data30_in(op2_00_in30),
    .data31_in(op2_00_bias),
    .data_out(op2_00_out));

  // 1 番目の OP2
  reg [8:0] op2_01_in00;
  reg [8:0] op2_01_in01;
  reg [8:0] op2_01_in02;
  reg [8:0] op2_01_in03;
  reg [8:0] op2_01_in04;
  reg [8:0] op2_01_in05;
  reg [8:0] op2_01_in06;
  reg [8:0] op2_01_in07;
  reg [8:0] op2_01_in08;
  reg [8:0] op2_01_in09;
  reg [8:0] op2_01_in10;
  reg [8:0] op2_01_in11;
  reg [8:0] op2_01_in12;
  reg [8:0] op2_01_in13;
  reg [8:0] op2_01_in14;
  reg [8:0] op2_01_in15;
  reg [8:0] op2_01_in16;
  reg [8:0] op2_01_in17;
  reg [8:0] op2_01_in18;
  reg [8:0] op2_01_in19;
  reg [8:0] op2_01_in20;
  reg [8:0] op2_01_in21;
  reg [8:0] op2_01_in22;
  reg [8:0] op2_01_in23;
  reg [8:0] op2_01_in24;
  reg [8:0] op2_01_in25;
  reg [8:0] op2_01_in26;
  reg [8:0] op2_01_in27;
  reg [8:0] op2_01_in28;
  reg [8:0] op2_01_in29;
  reg [8:0] op2_01_in30;
  reg [8:0] op2_01_bias;
  wire [8:0] op2_01_out;
  op2 op2_01(
    .data0_in(op2_01_in00),
    .data1_in(op2_01_in01),
    .data2_in(op2_01_in02),
    .data3_in(op2_01_in03),
    .data4_in(op2_01_in04),
    .data5_in(op2_01_in05),
    .data6_in(op2_01_in06),
    .data7_in(op2_01_in07),
    .data8_in(op2_01_in08),
    .data9_in(op2_01_in09),
    .data10_in(op2_01_in10),
    .data11_in(op2_01_in11),
    .data12_in(op2_01_in12),
    .data13_in(op2_01_in13),
    .data14_in(op2_01_in14),
    .data15_in(op2_01_in15),
    .data16_in(op2_01_in16),
    .data17_in(op2_01_in17),
    .data18_in(op2_01_in18),
    .data19_in(op2_01_in19),
    .data20_in(op2_01_in20),
    .data21_in(op2_01_in21),
    .data22_in(op2_01_in22),
    .data23_in(op2_01_in23),
    .data24_in(op2_01_in24),
    .data25_in(op2_01_in25),
    .data26_in(op2_01_in26),
    .data27_in(op2_01_in27),
    .data28_in(op2_01_in28),
    .data29_in(op2_01_in29),
    .data30_in(op2_01_in30),
    .data31_in(op2_01_bias),
    .data_out(op2_01_out));

  // 2 番目の OP2
  reg [8:0] op2_02_in00;
  reg [8:0] op2_02_in01;
  reg [8:0] op2_02_in02;
  reg [8:0] op2_02_in03;
  reg [8:0] op2_02_in04;
  reg [8:0] op2_02_in05;
  reg [8:0] op2_02_in06;
  reg [8:0] op2_02_in07;
  reg [8:0] op2_02_in08;
  reg [8:0] op2_02_in09;
  reg [8:0] op2_02_in10;
  reg [8:0] op2_02_in11;
  reg [8:0] op2_02_in12;
  reg [8:0] op2_02_in13;
  reg [8:0] op2_02_in14;
  reg [8:0] op2_02_in15;
  reg [8:0] op2_02_in16;
  reg [8:0] op2_02_in17;
  reg [8:0] op2_02_in18;
  reg [8:0] op2_02_in19;
  reg [8:0] op2_02_in20;
  reg [8:0] op2_02_in21;
  reg [8:0] op2_02_in22;
  reg [8:0] op2_02_in23;
  reg [8:0] op2_02_in24;
  reg [8:0] op2_02_in25;
  reg [8:0] op2_02_in26;
  reg [8:0] op2_02_in27;
  reg [8:0] op2_02_in28;
  reg [8:0] op2_02_in29;
  reg [8:0] op2_02_in30;
  reg [8:0] op2_02_bias;
  wire [8:0] op2_02_out;
  op2 op2_02(
    .data0_in(op2_02_in00),
    .data1_in(op2_02_in01),
    .data2_in(op2_02_in02),
    .data3_in(op2_02_in03),
    .data4_in(op2_02_in04),
    .data5_in(op2_02_in05),
    .data6_in(op2_02_in06),
    .data7_in(op2_02_in07),
    .data8_in(op2_02_in08),
    .data9_in(op2_02_in09),
    .data10_in(op2_02_in10),
    .data11_in(op2_02_in11),
    .data12_in(op2_02_in12),
    .data13_in(op2_02_in13),
    .data14_in(op2_02_in14),
    .data15_in(op2_02_in15),
    .data16_in(op2_02_in16),
    .data17_in(op2_02_in17),
    .data18_in(op2_02_in18),
    .data19_in(op2_02_in19),
    .data20_in(op2_02_in20),
    .data21_in(op2_02_in21),
    .data22_in(op2_02_in22),
    .data23_in(op2_02_in23),
    .data24_in(op2_02_in24),
    .data25_in(op2_02_in25),
    .data26_in(op2_02_in26),
    .data27_in(op2_02_in27),
    .data28_in(op2_02_in28),
    .data29_in(op2_02_in29),
    .data30_in(op2_02_in30),
    .data31_in(op2_02_bias),
    .data_out(op2_02_out));

  // 3 番目の OP2
  reg [8:0] op2_03_in00;
  reg [8:0] op2_03_in01;
  reg [8:0] op2_03_in02;
  reg [8:0] op2_03_in03;
  reg [8:0] op2_03_in04;
  reg [8:0] op2_03_in05;
  reg [8:0] op2_03_in06;
  reg [8:0] op2_03_in07;
  reg [8:0] op2_03_in08;
  reg [8:0] op2_03_in09;
  reg [8:0] op2_03_in10;
  reg [8:0] op2_03_in11;
  reg [8:0] op2_03_in12;
  reg [8:0] op2_03_in13;
  reg [8:0] op2_03_in14;
  reg [8:0] op2_03_in15;
  reg [8:0] op2_03_in16;
  reg [8:0] op2_03_in17;
  reg [8:0] op2_03_in18;
  reg [8:0] op2_03_in19;
  reg [8:0] op2_03_in20;
  reg [8:0] op2_03_in21;
  reg [8:0] op2_03_in22;
  reg [8:0] op2_03_in23;
  reg [8:0] op2_03_in24;
  reg [8:0] op2_03_in25;
  reg [8:0] op2_03_in26;
  reg [8:0] op2_03_in27;
  reg [8:0] op2_03_in28;
  reg [8:0] op2_03_in29;
  reg [8:0] op2_03_in30;
  reg [8:0] op2_03_bias;
  wire [8:0] op2_03_out;
  op2 op2_03(
    .data0_in(op2_03_in00),
    .data1_in(op2_03_in01),
    .data2_in(op2_03_in02),
    .data3_in(op2_03_in03),
    .data4_in(op2_03_in04),
    .data5_in(op2_03_in05),
    .data6_in(op2_03_in06),
    .data7_in(op2_03_in07),
    .data8_in(op2_03_in08),
    .data9_in(op2_03_in09),
    .data10_in(op2_03_in10),
    .data11_in(op2_03_in11),
    .data12_in(op2_03_in12),
    .data13_in(op2_03_in13),
    .data14_in(op2_03_in14),
    .data15_in(op2_03_in15),
    .data16_in(op2_03_in16),
    .data17_in(op2_03_in17),
    .data18_in(op2_03_in18),
    .data19_in(op2_03_in19),
    .data20_in(op2_03_in20),
    .data21_in(op2_03_in21),
    .data22_in(op2_03_in22),
    .data23_in(op2_03_in23),
    .data24_in(op2_03_in24),
    .data25_in(op2_03_in25),
    .data26_in(op2_03_in26),
    .data27_in(op2_03_in27),
    .data28_in(op2_03_in28),
    .data29_in(op2_03_in29),
    .data30_in(op2_03_in30),
    .data31_in(op2_03_bias),
    .data_out(op2_03_out));

  // 中間レジスタ
  reg [8:0] reg_0000;
  reg [8:0] reg_0001;
  reg [8:0] reg_0002;
  reg [8:0] reg_0003;
  reg [8:0] reg_0004;
  reg [8:0] reg_0005;
  reg [8:0] reg_0006;
  reg [8:0] reg_0007;
  reg [8:0] reg_0008;
  reg [8:0] reg_0009;
  reg [8:0] reg_0010;
  reg [8:0] reg_0011;
  reg [8:0] reg_0012;
  reg [8:0] reg_0013;
  reg [8:0] reg_0014;
  reg [8:0] reg_0015;
  reg [8:0] reg_0016;
  reg [8:0] reg_0017;
  reg [8:0] reg_0018;
  reg [8:0] reg_0019;
  reg [8:0] reg_0020;
  reg [8:0] reg_0021;
  reg [8:0] reg_0022;
  reg [8:0] reg_0023;
  reg [8:0] reg_0024;
  reg [8:0] reg_0025;
  reg [8:0] reg_0026;
  reg [8:0] reg_0027;
  reg [8:0] reg_0028;
  reg [8:0] reg_0029;
  reg [8:0] reg_0030;
  reg [8:0] reg_0031;
  reg [8:0] reg_0032;
  reg [8:0] reg_0033;
  reg [8:0] reg_0034;
  reg [8:0] reg_0035;
  reg [8:0] reg_0036;
  reg [8:0] reg_0037;
  reg [8:0] reg_0038;
  reg [8:0] reg_0039;
  reg [8:0] reg_0040;
  reg [8:0] reg_0041;
  reg [8:0] reg_0042;
  reg [8:0] reg_0043;
  reg [8:0] reg_0044;
  reg [8:0] reg_0045;
  reg [8:0] reg_0046;
  reg [8:0] reg_0047;
  reg [8:0] reg_0048;
  reg [8:0] reg_0049;
  reg [8:0] reg_0050;
  reg [8:0] reg_0051;
  reg [8:0] reg_0052;
  reg [8:0] reg_0053;
  reg [8:0] reg_0054;
  reg [8:0] reg_0055;
  reg [8:0] reg_0056;
  reg [8:0] reg_0057;
  reg [8:0] reg_0058;
  reg [8:0] reg_0059;
  reg [8:0] reg_0060;
  reg [8:0] reg_0061;
  reg [8:0] reg_0062;
  reg [8:0] reg_0063;
  reg [8:0] reg_0064;
  reg [8:0] reg_0065;
  reg [8:0] reg_0066;
  reg [8:0] reg_0067;
  reg [8:0] reg_0068;
  reg [8:0] reg_0069;
  reg [8:0] reg_0070;
  reg [8:0] reg_0071;
  reg [8:0] reg_0072;
  reg [8:0] reg_0073;
  reg [8:0] reg_0074;
  reg [8:0] reg_0075;
  reg [8:0] reg_0076;
  reg [8:0] reg_0077;
  reg [8:0] reg_0078;
  reg [8:0] reg_0079;
  reg [8:0] reg_0080;
  reg [8:0] reg_0081;
  reg [8:0] reg_0082;
  reg [8:0] reg_0083;
  reg [8:0] reg_0084;
  reg [8:0] reg_0085;
  reg [8:0] reg_0086;
  reg [8:0] reg_0087;
  reg [8:0] reg_0088;
  reg [8:0] reg_0089;
  reg [8:0] reg_0090;
  reg [8:0] reg_0091;
  reg [8:0] reg_0092;
  reg [8:0] reg_0093;
  reg [8:0] reg_0094;
  reg [8:0] reg_0095;
  reg [8:0] reg_0096;
  reg [8:0] reg_0097;
  reg [8:0] reg_0098;
  reg [8:0] reg_0099;
  reg [8:0] reg_0100;
  reg [8:0] reg_0101;
  reg [8:0] reg_0102;
  reg [8:0] reg_0103;
  reg [8:0] reg_0104;
  reg [8:0] reg_0105;
  reg [8:0] reg_0106;
  reg [8:0] reg_0107;
  reg [8:0] reg_0108;
  reg [8:0] reg_0109;
  reg [8:0] reg_0110;
  reg [8:0] reg_0111;
  reg [8:0] reg_0112;
  reg [8:0] reg_0113;
  reg [8:0] reg_0114;
  reg [8:0] reg_0115;
  reg [8:0] reg_0116;
  reg [8:0] reg_0117;
  reg [8:0] reg_0118;
  reg [8:0] reg_0119;
  reg [8:0] reg_0120;
  reg [8:0] reg_0121;
  reg [8:0] reg_0122;
  reg [8:0] reg_0123;
  reg [8:0] reg_0124;
  reg [8:0] reg_0125;
  reg [8:0] reg_0126;
  reg [8:0] reg_0127;
  reg [8:0] reg_0128;
  reg [8:0] reg_0129;
  reg [8:0] reg_0130;
  reg [8:0] reg_0131;
  reg [8:0] reg_0132;
  reg [8:0] reg_0133;
  reg [8:0] reg_0134;
  reg [8:0] reg_0135;
  reg [8:0] reg_0136;
  reg [8:0] reg_0137;
  reg [8:0] reg_0138;
  reg [8:0] reg_0139;
  reg [8:0] reg_0140;
  reg [8:0] reg_0141;
  reg [8:0] reg_0142;
  reg [8:0] reg_0143;
  reg [8:0] reg_0144;
  reg [8:0] reg_0145;
  reg [8:0] reg_0146;
  reg [8:0] reg_0147;
  reg [8:0] reg_0148;
  reg [8:0] reg_0149;
  reg [8:0] reg_0150;
  reg [8:0] reg_0151;
  reg [8:0] reg_0152;
  reg [8:0] reg_0153;
  reg [8:0] reg_0154;
  reg [8:0] reg_0155;
  reg [8:0] reg_0156;
  reg [8:0] reg_0157;
  reg [8:0] reg_0158;
  reg [8:0] reg_0159;
  reg [8:0] reg_0160;
  reg [8:0] reg_0161;
  reg [8:0] reg_0162;
  reg [8:0] reg_0163;
  reg [8:0] reg_0164;
  reg [8:0] reg_0165;
  reg [8:0] reg_0166;
  reg [8:0] reg_0167;
  reg [8:0] reg_0168;
  reg [8:0] reg_0169;
  reg [8:0] reg_0170;
  reg [8:0] reg_0171;
  reg [8:0] reg_0172;
  reg [8:0] reg_0173;
  reg [8:0] reg_0174;
  reg [8:0] reg_0175;
  reg [8:0] reg_0176;
  reg [8:0] reg_0177;
  reg [8:0] reg_0178;
  reg [8:0] reg_0179;
  reg [8:0] reg_0180;
  reg [8:0] reg_0181;
  reg [8:0] reg_0182;
  reg [8:0] reg_0183;
  reg [8:0] reg_0184;
  reg [8:0] reg_0185;
  reg [8:0] reg_0186;
  reg [8:0] reg_0187;
  reg [8:0] reg_0188;
  reg [8:0] reg_0189;
  reg [8:0] reg_0190;
  reg [8:0] reg_0191;
  reg [8:0] reg_0192;
  reg [8:0] reg_0193;
  reg [8:0] reg_0194;
  reg [8:0] reg_0195;
  reg [8:0] reg_0196;
  reg [8:0] reg_0197;
  reg [8:0] reg_0198;
  reg [8:0] reg_0199;
  reg [8:0] reg_0200;
  reg [8:0] reg_0201;
  reg [8:0] reg_0202;
  reg [8:0] reg_0203;
  reg [8:0] reg_0204;
  reg [8:0] reg_0205;
  reg [8:0] reg_0206;
  reg [8:0] reg_0207;
  reg [8:0] reg_0208;
  reg [8:0] reg_0209;
  reg [8:0] reg_0210;
  reg [8:0] reg_0211;
  reg [8:0] reg_0212;
  reg [8:0] reg_0213;
  reg [8:0] reg_0214;
  reg [8:0] reg_0215;
  reg [8:0] reg_0216;
  reg [8:0] reg_0217;
  reg [8:0] reg_0218;
  reg [8:0] reg_0219;
  reg [8:0] reg_0220;
  reg [8:0] reg_0221;
  reg [8:0] reg_0222;
  reg [8:0] reg_0223;
  reg [8:0] reg_0224;
  reg [8:0] reg_0225;
  reg [8:0] reg_0226;
  reg [8:0] reg_0227;
  reg [8:0] reg_0228;
  reg [8:0] reg_0229;
  reg [8:0] reg_0230;
  reg [8:0] reg_0231;
  reg [8:0] reg_0232;
  reg [8:0] reg_0233;
  reg [8:0] reg_0234;
  reg [8:0] reg_0235;
  reg [8:0] reg_0236;
  reg [8:0] reg_0237;
  reg [8:0] reg_0238;
  reg [8:0] reg_0239;
  reg [8:0] reg_0240;
  reg [8:0] reg_0241;
  reg [8:0] reg_0242;
  reg [8:0] reg_0243;
  reg [8:0] reg_0244;
  reg [8:0] reg_0245;
  reg [8:0] reg_0246;
  reg [8:0] reg_0247;
  reg [8:0] reg_0248;
  reg [8:0] reg_0249;
  reg [8:0] reg_0250;
  reg [8:0] reg_0251;
  reg [8:0] reg_0252;
  reg [8:0] reg_0253;
  reg [8:0] reg_0254;
  reg [8:0] reg_0255;
  reg [8:0] reg_0256;
  reg [8:0] reg_0257;
  reg [8:0] reg_0258;
  reg [8:0] reg_0259;
  reg [8:0] reg_0260;
  reg [8:0] reg_0261;
  reg [8:0] reg_0262;
  reg [8:0] reg_0263;
  reg [8:0] reg_0264;
  reg [8:0] reg_0265;
  reg [8:0] reg_0266;
  reg [8:0] reg_0267;
  reg [8:0] reg_0268;
  reg [8:0] reg_0269;
  reg [8:0] reg_0270;
  reg [8:0] reg_0271;
  reg [8:0] reg_0272;
  reg [8:0] reg_0273;
  reg [8:0] reg_0274;
  reg [8:0] reg_0275;
  reg [8:0] reg_0276;
  reg [8:0] reg_0277;
  reg [8:0] reg_0278;
  reg [8:0] reg_0279;
  reg [8:0] reg_0280;
  reg [8:0] reg_0281;
  reg [8:0] reg_0282;
  reg [8:0] reg_0283;
  reg [8:0] reg_0284;
  reg [8:0] reg_0285;
  reg [8:0] reg_0286;
  reg [8:0] reg_0287;
  reg [8:0] reg_0288;
  reg [8:0] reg_0289;
  reg [8:0] reg_0290;
  reg [8:0] reg_0291;
  reg [8:0] reg_0292;
  reg [8:0] reg_0293;
  reg [8:0] reg_0294;
  reg [8:0] reg_0295;
  reg [8:0] reg_0296;
  reg [8:0] reg_0297;
  reg [8:0] reg_0298;
  reg [8:0] reg_0299;
  reg [8:0] reg_0300;
  reg [8:0] reg_0301;
  reg [8:0] reg_0302;
  reg [8:0] reg_0303;
  reg [8:0] reg_0304;
  reg [8:0] reg_0305;
  reg [8:0] reg_0306;
  reg [8:0] reg_0307;
  reg [8:0] reg_0308;
  reg [8:0] reg_0309;
  reg [8:0] reg_0310;
  reg [8:0] reg_0311;
  reg [8:0] reg_0312;
  reg [8:0] reg_0313;
  reg [8:0] reg_0314;
  reg [8:0] reg_0315;
  reg [8:0] reg_0316;
  reg [8:0] reg_0317;
  reg [8:0] reg_0318;
  reg [8:0] reg_0319;
  reg [8:0] reg_0320;
  reg [8:0] reg_0321;
  reg [8:0] reg_0322;
  reg [8:0] reg_0323;
  reg [8:0] reg_0324;
  reg [8:0] reg_0325;
  reg [8:0] reg_0326;
  reg [8:0] reg_0327;
  reg [8:0] reg_0328;
  reg [8:0] reg_0329;
  reg [8:0] reg_0330;
  reg [8:0] reg_0331;
  reg [8:0] reg_0332;
  reg [8:0] reg_0333;
  reg [8:0] reg_0334;
  reg [8:0] reg_0335;
  reg [8:0] reg_0336;
  reg [8:0] reg_0337;
  reg [8:0] reg_0338;
  reg [8:0] reg_0339;
  reg [8:0] reg_0340;
  reg [8:0] reg_0341;
  reg [8:0] reg_0342;
  reg [8:0] reg_0343;
  reg [8:0] reg_0344;
  reg [8:0] reg_0345;
  reg [8:0] reg_0346;
  reg [8:0] reg_0347;
  reg [8:0] reg_0348;
  reg [8:0] reg_0349;
  reg [8:0] reg_0350;
  reg [8:0] reg_0351;
  reg [8:0] reg_0352;
  reg [8:0] reg_0353;
  reg [8:0] reg_0354;
  reg [8:0] reg_0355;
  reg [8:0] reg_0356;
  reg [8:0] reg_0357;
  reg [8:0] reg_0358;
  reg [8:0] reg_0359;
  reg [8:0] reg_0360;
  reg [8:0] reg_0361;
  reg [8:0] reg_0362;
  reg [8:0] reg_0363;
  reg [8:0] reg_0364;
  reg [8:0] reg_0365;
  reg [8:0] reg_0366;
  reg [8:0] reg_0367;
  reg [8:0] reg_0368;
  reg [8:0] reg_0369;
  reg [8:0] reg_0370;
  reg [8:0] reg_0371;
  reg [8:0] reg_0372;
  reg [8:0] reg_0373;
  reg [8:0] reg_0374;
  reg [8:0] reg_0375;
  reg [8:0] reg_0376;
  reg [8:0] reg_0377;
  reg [8:0] reg_0378;
  reg [8:0] reg_0379;
  reg [8:0] reg_0380;
  reg [8:0] reg_0381;
  reg [8:0] reg_0382;
  reg [8:0] reg_0383;
  reg [8:0] reg_0384;
  reg [8:0] reg_0385;
  reg [8:0] reg_0386;
  reg [8:0] reg_0387;
  reg [8:0] reg_0388;
  reg [8:0] reg_0389;
  reg [8:0] reg_0390;
  reg [8:0] reg_0391;
  reg [8:0] reg_0392;
  reg [8:0] reg_0393;
  reg [8:0] reg_0394;
  reg [8:0] reg_0395;
  reg [8:0] reg_0396;
  reg [8:0] reg_0397;
  reg [8:0] reg_0398;
  reg [8:0] reg_0399;
  reg [8:0] reg_0400;
  reg [8:0] reg_0401;
  reg [8:0] reg_0402;
  reg [8:0] reg_0403;
  reg [8:0] reg_0404;
  reg [8:0] reg_0405;
  reg [8:0] reg_0406;
  reg [8:0] reg_0407;
  reg [8:0] reg_0408;
  reg [8:0] reg_0409;
  reg [8:0] reg_0410;
  reg [8:0] reg_0411;
  reg [8:0] reg_0412;
  reg [8:0] reg_0413;
  reg [8:0] reg_0414;
  reg [8:0] reg_0415;
  reg [8:0] reg_0416;
  reg [8:0] reg_0417;
  reg [8:0] reg_0418;
  reg [8:0] reg_0419;
  reg [8:0] reg_0420;
  reg [8:0] reg_0421;
  reg [8:0] reg_0422;
  reg [8:0] reg_0423;
  reg [8:0] reg_0424;
  reg [8:0] reg_0425;
  reg [8:0] reg_0426;
  reg [8:0] reg_0427;
  reg [8:0] reg_0428;
  reg [8:0] reg_0429;
  reg [8:0] reg_0430;
  reg [8:0] reg_0431;
  reg [8:0] reg_0432;
  reg [8:0] reg_0433;
  reg [8:0] reg_0434;
  reg [8:0] reg_0435;
  reg [8:0] reg_0436;
  reg [8:0] reg_0437;
  reg [8:0] reg_0438;
  reg [8:0] reg_0439;
  reg [8:0] reg_0440;
  reg [8:0] reg_0441;
  reg [8:0] reg_0442;
  reg [8:0] reg_0443;
  reg [8:0] reg_0444;
  reg [8:0] reg_0445;
  reg [8:0] reg_0446;
  reg [8:0] reg_0447;
  reg [8:0] reg_0448;
  reg [8:0] reg_0449;
  reg [8:0] reg_0450;
  reg [8:0] reg_0451;
  reg [8:0] reg_0452;
  reg [8:0] reg_0453;
  reg [8:0] reg_0454;
  reg [8:0] reg_0455;
  reg [8:0] reg_0456;
  reg [8:0] reg_0457;
  reg [8:0] reg_0458;
  reg [8:0] reg_0459;
  reg [8:0] reg_0460;
  reg [8:0] reg_0461;
  reg [8:0] reg_0462;
  reg [8:0] reg_0463;
  reg [8:0] reg_0464;
  reg [8:0] reg_0465;
  reg [8:0] reg_0466;
  reg [8:0] reg_0467;
  reg [8:0] reg_0468;
  reg [8:0] reg_0469;
  reg [8:0] reg_0470;
  reg [8:0] reg_0471;
  reg [8:0] reg_0472;
  reg [8:0] reg_0473;
  reg [8:0] reg_0474;
  reg [8:0] reg_0475;
  reg [8:0] reg_0476;
  reg [8:0] reg_0477;
  reg [8:0] reg_0478;
  reg [8:0] reg_0479;
  reg [8:0] reg_0480;
  reg [8:0] reg_0481;
  reg [8:0] reg_0482;
  reg [8:0] reg_0483;
  reg [8:0] reg_0484;
  reg [8:0] reg_0485;
  reg [8:0] reg_0486;
  reg [8:0] reg_0487;
  reg [8:0] reg_0488;
  reg [8:0] reg_0489;
  reg [8:0] reg_0490;
  reg [8:0] reg_0491;
  reg [8:0] reg_0492;
  reg [8:0] reg_0493;
  reg [8:0] reg_0494;
  reg [8:0] reg_0495;
  reg [8:0] reg_0496;
  reg [8:0] reg_0497;
  reg [8:0] reg_0498;
  reg [8:0] reg_0499;
  reg [8:0] reg_0500;
  reg [8:0] reg_0501;
  reg [8:0] reg_0502;
  reg [8:0] reg_0503;
  reg [8:0] reg_0504;
  reg [8:0] reg_0505;
  reg [8:0] reg_0506;
  reg [8:0] reg_0507;
  reg [8:0] reg_0508;
  reg [8:0] reg_0509;
  reg [8:0] reg_0510;
  reg [8:0] reg_0511;
  reg [8:0] reg_0512;
  reg [8:0] reg_0513;
  reg [8:0] reg_0514;
  reg [8:0] reg_0515;
  reg [8:0] reg_0516;
  reg [8:0] reg_0517;
  reg [8:0] reg_0518;
  reg [8:0] reg_0519;
  reg [8:0] reg_0520;
  reg [8:0] reg_0521;
  reg [8:0] reg_0522;
  reg [8:0] reg_0523;
  reg [8:0] reg_0524;
  reg [8:0] reg_0525;
  reg [8:0] reg_0526;
  reg [8:0] reg_0527;
  reg [8:0] reg_0528;
  reg [8:0] reg_0529;
  reg [8:0] reg_0530;
  reg [8:0] reg_0531;
  reg [8:0] reg_0532;
  reg [8:0] reg_0533;
  reg [8:0] reg_0534;
  reg [8:0] reg_0535;
  reg [8:0] reg_0536;
  reg [8:0] reg_0537;
  reg [8:0] reg_0538;
  reg [8:0] reg_0539;
  reg [8:0] reg_0540;
  reg [8:0] reg_0541;
  reg [8:0] reg_0542;
  reg [8:0] reg_0543;
  reg [8:0] reg_0544;
  reg [8:0] reg_0545;
  reg [8:0] reg_0546;
  reg [8:0] reg_0547;
  reg [8:0] reg_0548;
  reg [8:0] reg_0549;
  reg [8:0] reg_0550;
  reg [8:0] reg_0551;
  reg [8:0] reg_0552;
  reg [8:0] reg_0553;
  reg [8:0] reg_0554;
  reg [8:0] reg_0555;
  reg [8:0] reg_0556;
  reg [8:0] reg_0557;
  reg [8:0] reg_0558;
  reg [8:0] reg_0559;
  reg [8:0] reg_0560;
  reg [8:0] reg_0561;
  reg [8:0] reg_0562;
  reg [8:0] reg_0563;
  reg [8:0] reg_0564;
  reg [8:0] reg_0565;
  reg [8:0] reg_0566;
  reg [8:0] reg_0567;
  reg [8:0] reg_0568;
  reg [8:0] reg_0569;
  reg [8:0] reg_0570;
  reg [8:0] reg_0571;
  reg [8:0] reg_0572;
  reg [8:0] reg_0573;
  reg [8:0] reg_0574;
  reg [8:0] reg_0575;
  reg [8:0] reg_0576;
  reg [8:0] reg_0577;
  reg [8:0] reg_0578;
  reg [8:0] reg_0579;
  reg [8:0] reg_0580;
  reg [8:0] reg_0581;
  reg [8:0] reg_0582;
  reg [8:0] reg_0583;
  reg [8:0] reg_0584;
  reg [8:0] reg_0585;
  reg [8:0] reg_0586;
  reg [8:0] reg_0587;
  reg [8:0] reg_0588;
  reg [8:0] reg_0589;
  reg [8:0] reg_0590;
  reg [8:0] reg_0591;
  reg [8:0] reg_0592;
  reg [8:0] reg_0593;
  reg [8:0] reg_0594;
  reg [8:0] reg_0595;
  reg [8:0] reg_0596;
  reg [8:0] reg_0597;
  reg [8:0] reg_0598;
  reg [8:0] reg_0599;
  reg [8:0] reg_0600;
  reg [8:0] reg_0601;
  reg [8:0] reg_0602;
  reg [8:0] reg_0603;
  reg [8:0] reg_0604;
  reg [8:0] reg_0605;
  reg [8:0] reg_0606;
  reg [8:0] reg_0607;
  reg [8:0] reg_0608;
  reg [8:0] reg_0609;
  reg [8:0] reg_0610;
  reg [8:0] reg_0611;
  reg [8:0] reg_0612;
  reg [8:0] reg_0613;
  reg [8:0] reg_0614;
  reg [8:0] reg_0615;
  reg [8:0] reg_0616;
  reg [8:0] reg_0617;
  reg [8:0] reg_0618;
  reg [8:0] reg_0619;
  reg [8:0] reg_0620;
  reg [8:0] reg_0621;
  reg [8:0] reg_0622;
  reg [8:0] reg_0623;
  reg [8:0] reg_0624;
  reg [8:0] reg_0625;
  reg [8:0] reg_0626;
  reg [8:0] reg_0627;
  reg [8:0] reg_0628;
  reg [8:0] reg_0629;
  reg [8:0] reg_0630;
  reg [8:0] reg_0631;
  reg [8:0] reg_0632;
  reg [8:0] reg_0633;
  reg [8:0] reg_0634;
  reg [8:0] reg_0635;
  reg [8:0] reg_0636;
  reg [8:0] reg_0637;
  reg [8:0] reg_0638;
  reg [8:0] reg_0639;
  reg [8:0] reg_0640;
  reg [8:0] reg_0641;
  reg [8:0] reg_0642;
  reg [8:0] reg_0643;
  reg [8:0] reg_0644;
  reg [8:0] reg_0645;
  reg [8:0] reg_0646;
  reg [8:0] reg_0647;
  reg [8:0] reg_0648;
  reg [8:0] reg_0649;
  reg [8:0] reg_0650;
  reg [8:0] reg_0651;
  reg [8:0] reg_0652;
  reg [8:0] reg_0653;
  reg [8:0] reg_0654;
  reg [8:0] reg_0655;
  reg [8:0] reg_0656;
  reg [8:0] reg_0657;
  reg [8:0] reg_0658;
  reg [8:0] reg_0659;
  reg [8:0] reg_0660;
  reg [8:0] reg_0661;
  reg [8:0] reg_0662;
  reg [8:0] reg_0663;
  reg [8:0] reg_0664;
  reg [8:0] reg_0665;
  reg [8:0] reg_0666;
  reg [8:0] reg_0667;
  reg [8:0] reg_0668;
  reg [8:0] reg_0669;
  reg [8:0] reg_0670;
  reg [8:0] reg_0671;
  reg [8:0] reg_0672;
  reg [8:0] reg_0673;
  reg [8:0] reg_0674;
  reg [8:0] reg_0675;
  reg [8:0] reg_0676;
  reg [8:0] reg_0677;
  reg [8:0] reg_0678;
  reg [8:0] reg_0679;
  reg [8:0] reg_0680;
  reg [8:0] reg_0681;
  reg [8:0] reg_0682;
  reg [8:0] reg_0683;
  reg [8:0] reg_0684;
  reg [8:0] reg_0685;
  reg [8:0] reg_0686;
  reg [8:0] reg_0687;
  reg [8:0] reg_0688;
  reg [8:0] reg_0689;
  reg [8:0] reg_0690;
  reg [8:0] reg_0691;
  reg [8:0] reg_0692;
  reg [8:0] reg_0693;
  reg [8:0] reg_0694;
  reg [8:0] reg_0695;
  reg [8:0] reg_0696;
  reg [8:0] reg_0697;
  reg [8:0] reg_0698;
  reg [8:0] reg_0699;
  reg [8:0] reg_0700;
  reg [8:0] reg_0701;
  reg [8:0] reg_0702;
  reg [8:0] reg_0703;
  reg [8:0] reg_0704;
  reg [8:0] reg_0705;
  reg [8:0] reg_0706;
  reg [8:0] reg_0707;
  reg [8:0] reg_0708;
  reg [8:0] reg_0709;
  reg [8:0] reg_0710;
  reg [8:0] reg_0711;
  reg [8:0] reg_0712;
  reg [8:0] reg_0713;
  reg [8:0] reg_0714;
  reg [8:0] reg_0715;
  reg [8:0] reg_0716;
  reg [8:0] reg_0717;
  reg [8:0] reg_0718;
  reg [8:0] reg_0719;
  reg [8:0] reg_0720;
  reg [8:0] reg_0721;
  reg [8:0] reg_0722;
  reg [8:0] reg_0723;
  reg [8:0] reg_0724;
  reg [8:0] reg_0725;
  reg [8:0] reg_0726;
  reg [8:0] reg_0727;
  reg [8:0] reg_0728;
  reg [8:0] reg_0729;
  reg [8:0] reg_0730;
  reg [8:0] reg_0731;
  reg [8:0] reg_0732;
  reg [8:0] reg_0733;
  reg [8:0] reg_0734;
  reg [8:0] reg_0735;
  reg [8:0] reg_0736;
  reg [8:0] reg_0737;
  reg [8:0] reg_0738;
  reg [8:0] reg_0739;
  reg [8:0] reg_0740;
  reg [8:0] reg_0741;
  reg [8:0] reg_0742;
  reg [8:0] reg_0743;
  reg [8:0] reg_0744;
  reg [8:0] reg_0745;
  reg [8:0] reg_0746;
  reg [8:0] reg_0747;
  reg [8:0] reg_0748;
  reg [8:0] reg_0749;
  reg [8:0] reg_0750;
  reg [8:0] reg_0751;
  reg [8:0] reg_0752;
  reg [8:0] reg_0753;
  reg [8:0] reg_0754;
  reg [8:0] reg_0755;
  reg [8:0] reg_0756;
  reg [8:0] reg_0757;
  reg [8:0] reg_0758;
  reg [8:0] reg_0759;
  reg [8:0] reg_0760;
  reg [8:0] reg_0761;
  reg [8:0] reg_0762;
  reg [8:0] reg_0763;
  reg [8:0] reg_0764;
  reg [8:0] reg_0765;
  reg [8:0] reg_0766;
  reg [8:0] reg_0767;
  reg [8:0] reg_0768;
  reg [8:0] reg_0769;
  reg [8:0] reg_0770;
  reg [8:0] reg_0771;
  reg [8:0] reg_0772;
  reg [8:0] reg_0773;
  reg [8:0] reg_0774;
  reg [8:0] reg_0775;
  reg [8:0] reg_0776;
  reg [8:0] reg_0777;
  reg [8:0] reg_0778;
  reg [8:0] reg_0779;
  reg [8:0] reg_0780;
  reg [8:0] reg_0781;
  reg [8:0] reg_0782;
  reg [8:0] reg_0783;
  reg [8:0] reg_0784;
  reg [8:0] reg_0785;
  reg [8:0] reg_0786;
  reg [8:0] reg_0787;
  reg [8:0] reg_0788;
  reg [8:0] reg_0789;
  reg [8:0] reg_0790;
  reg [8:0] reg_0791;
  reg [8:0] reg_0792;
  reg [8:0] reg_0793;
  reg [8:0] reg_0794;
  reg [8:0] reg_0795;
  reg [8:0] reg_0796;
  reg [8:0] reg_0797;
  reg [8:0] reg_0798;
  reg [8:0] reg_0799;
  reg [8:0] reg_0800;
  reg [8:0] reg_0801;
  reg [8:0] reg_0802;
  reg [8:0] reg_0803;
  reg [8:0] reg_0804;
  reg [8:0] reg_0805;
  reg [8:0] reg_0806;
  reg [8:0] reg_0807;
  reg [8:0] reg_0808;
  reg [8:0] reg_0809;
  reg [8:0] reg_0810;
  reg [8:0] reg_0811;
  reg [8:0] reg_0812;
  reg [8:0] reg_0813;
  reg [8:0] reg_0814;
  reg [8:0] reg_0815;
  reg [8:0] reg_0816;
  reg [8:0] reg_0817;
  reg [8:0] reg_0818;
  reg [8:0] reg_0819;
  reg [8:0] reg_0820;
  reg [8:0] reg_0821;
  reg [8:0] reg_0822;
  reg [8:0] reg_0823;
  reg [8:0] reg_0824;
  reg [8:0] reg_0825;
  reg [8:0] reg_0826;
  reg [8:0] reg_0827;
  reg [8:0] reg_0828;
  reg [8:0] reg_0829;
  reg [8:0] reg_0830;
  reg [8:0] reg_0831;

  // 制御マシンの状態
  reg [7:0] state;
  reg _busy;
  assign busy = _busy;
  // 制御マシンの動作
  always @ ( posedge clock or negedge reset ) begin
    if ( !reset ) begin
      _busy <= 0;
      state <= 0;
    end
    else if ( _busy ) begin
      if ( state < 137 ) begin
        state <= state + 1;
      end
      else begin
        _busy <= 0;
        state <= 0;
      end
    end
    else if ( start ) begin
      _busy <= 1;
    end
  end

  // 0番目の入力用メモリブロックの制御
  reg [1:0] _imem00_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem00_bank = 0;
    2: _imem00_bank = 1;
    1: _imem00_bank = 2;
    0: _imem00_bank = 3;
    4: _imem00_bank = 0;
    5: _imem00_bank = 0;
    6: _imem00_bank = 0;
    7: _imem00_bank = 0;
    8: _imem00_bank = 0;
    9: _imem00_bank = 0;
    10: _imem00_bank = 0;
    11: _imem00_bank = 0;
    12: _imem00_bank = 0;
    13: _imem00_bank = 0;
    14: _imem00_bank = 0;
    15: _imem00_bank = 0;
    16: _imem00_bank = 0;
    17: _imem00_bank = 0;
    18: _imem00_bank = 0;
    19: _imem00_bank = 0;
    20: _imem00_bank = 0;
    21: _imem00_bank = 0;
    22: _imem00_bank = 0;
    23: _imem00_bank = 0;
    24: _imem00_bank = 0;
    25: _imem00_bank = 0;
    26: _imem00_bank = 0;
    27: _imem00_bank = 0;
    28: _imem00_bank = 0;
    29: _imem00_bank = 0;
    30: _imem00_bank = 0;
    31: _imem00_bank = 0;
    32: _imem00_bank = 0;
    33: _imem00_bank = 0;
    34: _imem00_bank = 0;
    35: _imem00_bank = 0;
    36: _imem00_bank = 0;
    37: _imem00_bank = 0;
    38: _imem00_bank = 0;
    39: _imem00_bank = 0;
    40: _imem00_bank = 0;
    41: _imem00_bank = 0;
    42: _imem00_bank = 0;
    43: _imem00_bank = 0;
    44: _imem00_bank = 0;
    45: _imem00_bank = 0;
    46: _imem00_bank = 0;
    47: _imem00_bank = 0;
    48: _imem00_bank = 0;
    49: _imem00_bank = 0;
    50: _imem00_bank = 0;
    51: _imem00_bank = 0;
    52: _imem00_bank = 0;
    53: _imem00_bank = 1;
    54: _imem00_bank = 0;
    55: _imem00_bank = 0;
    56: _imem00_bank = 0;
    57: _imem00_bank = 0;
    58: _imem00_bank = 0;
    59: _imem00_bank = 0;
    60: _imem00_bank = 0;
    61: _imem00_bank = 0;
    62: _imem00_bank = 0;
    63: _imem00_bank = 0;
    64: _imem00_bank = 0;
    65: _imem00_bank = 0;
    66: _imem00_bank = 0;
    67: _imem00_bank = 0;
    68: _imem00_bank = 0;
    69: _imem00_bank = 0;
    70: _imem00_bank = 0;
    71: _imem00_bank = 0;
    72: _imem00_bank = 0;
    73: _imem00_bank = 0;
    74: _imem00_bank = 0;
    75: _imem00_bank = 0;
    76: _imem00_bank = 0;
    77: _imem00_bank = 0;
    78: _imem00_bank = 0;
    79: _imem00_bank = 0;
    80: _imem00_bank = 0;
    81: _imem00_bank = 0;
    82: _imem00_bank = 0;
    83: _imem00_bank = 0;
    84: _imem00_bank = 0;
    85: _imem00_bank = 0;
    86: _imem00_bank = 0;
    87: _imem00_bank = 0;
    88: _imem00_bank = 0;
    89: _imem00_bank = 1;
    90: _imem00_bank = 0;
    91: _imem00_bank = 0;
    92: _imem00_bank = 0;
    93: _imem00_bank = 0;
    94: _imem00_bank = 0;
    95: _imem00_bank = 0;
    default: _imem00_bank = 0;
    endcase
  end // always @ ( * )
  assign imem00_bank = _imem00_bank;
  reg _imem00_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem00_rd = 1;
    2: _imem00_rd = 1;
    1: _imem00_rd = 1;
    0: _imem00_rd = 1;
    4: _imem00_rd = 1;
    5: _imem00_rd = 1;
    6: _imem00_rd = 1;
    7: _imem00_rd = 1;
    8: _imem00_rd = 1;
    9: _imem00_rd = 1;
    10: _imem00_rd = 1;
    11: _imem00_rd = 1;
    12: _imem00_rd = 1;
    13: _imem00_rd = 1;
    14: _imem00_rd = 1;
    15: _imem00_rd = 1;
    16: _imem00_rd = 1;
    17: _imem00_rd = 1;
    18: _imem00_rd = 1;
    19: _imem00_rd = 1;
    20: _imem00_rd = 1;
    21: _imem00_rd = 1;
    22: _imem00_rd = 1;
    23: _imem00_rd = 1;
    24: _imem00_rd = 1;
    25: _imem00_rd = 1;
    26: _imem00_rd = 1;
    27: _imem00_rd = 1;
    28: _imem00_rd = 1;
    29: _imem00_rd = 1;
    30: _imem00_rd = 1;
    31: _imem00_rd = 1;
    32: _imem00_rd = 1;
    33: _imem00_rd = 1;
    34: _imem00_rd = 1;
    35: _imem00_rd = 1;
    36: _imem00_rd = 1;
    37: _imem00_rd = 1;
    38: _imem00_rd = 1;
    39: _imem00_rd = 1;
    40: _imem00_rd = 1;
    41: _imem00_rd = 1;
    42: _imem00_rd = 1;
    43: _imem00_rd = 1;
    44: _imem00_rd = 1;
    45: _imem00_rd = 1;
    46: _imem00_rd = 1;
    47: _imem00_rd = 1;
    48: _imem00_rd = 1;
    49: _imem00_rd = 1;
    50: _imem00_rd = 1;
    51: _imem00_rd = 1;
    52: _imem00_rd = 1;
    53: _imem00_rd = 1;
    54: _imem00_rd = 1;
    55: _imem00_rd = 1;
    56: _imem00_rd = 1;
    57: _imem00_rd = 1;
    58: _imem00_rd = 1;
    59: _imem00_rd = 1;
    60: _imem00_rd = 1;
    61: _imem00_rd = 1;
    62: _imem00_rd = 1;
    63: _imem00_rd = 1;
    64: _imem00_rd = 1;
    65: _imem00_rd = 1;
    66: _imem00_rd = 1;
    67: _imem00_rd = 1;
    68: _imem00_rd = 1;
    69: _imem00_rd = 1;
    70: _imem00_rd = 1;
    71: _imem00_rd = 1;
    72: _imem00_rd = 1;
    73: _imem00_rd = 1;
    74: _imem00_rd = 1;
    75: _imem00_rd = 1;
    76: _imem00_rd = 1;
    77: _imem00_rd = 1;
    78: _imem00_rd = 1;
    79: _imem00_rd = 1;
    80: _imem00_rd = 1;
    81: _imem00_rd = 1;
    82: _imem00_rd = 1;
    83: _imem00_rd = 1;
    84: _imem00_rd = 1;
    85: _imem00_rd = 1;
    86: _imem00_rd = 1;
    87: _imem00_rd = 1;
    88: _imem00_rd = 1;
    89: _imem00_rd = 1;
    90: _imem00_rd = 1;
    91: _imem00_rd = 1;
    92: _imem00_rd = 1;
    93: _imem00_rd = 1;
    94: _imem00_rd = 1;
    95: _imem00_rd = 1;
    default: _imem00_rd = 0;
    endcase
  end // always @ ( * )
  assign imem00_rd = _imem00_rd;

  // 1番目の入力用メモリブロックの制御
  reg [1:0] _imem01_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem01_bank = 0;
    2: _imem01_bank = 1;
    1: _imem01_bank = 2;
    0: _imem01_bank = 3;
    4: _imem01_bank = 0;
    5: _imem01_bank = 0;
    6: _imem01_bank = 0;
    7: _imem01_bank = 0;
    8: _imem01_bank = 2;
    9: _imem01_bank = 1;
    10: _imem01_bank = 0;
    11: _imem01_bank = 0;
    12: _imem01_bank = 0;
    13: _imem01_bank = 0;
    14: _imem01_bank = 0;
    15: _imem01_bank = 0;
    16: _imem01_bank = 0;
    17: _imem01_bank = 0;
    18: _imem01_bank = 0;
    19: _imem01_bank = 0;
    20: _imem01_bank = 0;
    21: _imem01_bank = 0;
    22: _imem01_bank = 0;
    23: _imem01_bank = 1;
    24: _imem01_bank = 0;
    25: _imem01_bank = 0;
    26: _imem01_bank = 0;
    27: _imem01_bank = 0;
    28: _imem01_bank = 0;
    29: _imem01_bank = 0;
    30: _imem01_bank = 0;
    31: _imem01_bank = 0;
    32: _imem01_bank = 0;
    33: _imem01_bank = 0;
    34: _imem01_bank = 0;
    35: _imem01_bank = 0;
    36: _imem01_bank = 0;
    37: _imem01_bank = 0;
    38: _imem01_bank = 2;
    39: _imem01_bank = 2;
    40: _imem01_bank = 0;
    41: _imem01_bank = 0;
    42: _imem01_bank = 0;
    43: _imem01_bank = 0;
    44: _imem01_bank = 0;
    45: _imem01_bank = 0;
    46: _imem01_bank = 1;
    47: _imem01_bank = 1;
    48: _imem01_bank = 0;
    49: _imem01_bank = 0;
    50: _imem01_bank = 0;
    51: _imem01_bank = 3;
    52: _imem01_bank = 0;
    53: _imem01_bank = 0;
    54: _imem01_bank = 0;
    55: _imem01_bank = 0;
    56: _imem01_bank = 0;
    57: _imem01_bank = 0;
    58: _imem01_bank = 0;
    59: _imem01_bank = 0;
    60: _imem01_bank = 0;
    61: _imem01_bank = 0;
    62: _imem01_bank = 0;
    63: _imem01_bank = 0;
    64: _imem01_bank = 0;
    65: _imem01_bank = 0;
    66: _imem01_bank = 0;
    67: _imem01_bank = 1;
    68: _imem01_bank = 0;
    69: _imem01_bank = 0;
    70: _imem01_bank = 0;
    71: _imem01_bank = 0;
    72: _imem01_bank = 0;
    73: _imem01_bank = 0;
    74: _imem01_bank = 0;
    75: _imem01_bank = 0;
    76: _imem01_bank = 0;
    77: _imem01_bank = 0;
    78: _imem01_bank = 0;
    79: _imem01_bank = 0;
    80: _imem01_bank = 0;
    81: _imem01_bank = 0;
    82: _imem01_bank = 0;
    83: _imem01_bank = 0;
    84: _imem01_bank = 0;
    85: _imem01_bank = 0;
    86: _imem01_bank = 0;
    87: _imem01_bank = 0;
    88: _imem01_bank = 0;
    89: _imem01_bank = 0;
    90: _imem01_bank = 0;
    91: _imem01_bank = 2;
    92: _imem01_bank = 1;
    93: _imem01_bank = 2;
    94: _imem01_bank = 1;
    95: _imem01_bank = 0;
    default: _imem01_bank = 0;
    endcase
  end // always @ ( * )
  assign imem01_bank = _imem01_bank;
  reg _imem01_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem01_rd = 1;
    2: _imem01_rd = 1;
    1: _imem01_rd = 1;
    0: _imem01_rd = 1;
    4: _imem01_rd = 1;
    5: _imem01_rd = 1;
    6: _imem01_rd = 1;
    7: _imem01_rd = 1;
    8: _imem01_rd = 1;
    9: _imem01_rd = 1;
    10: _imem01_rd = 1;
    11: _imem01_rd = 1;
    12: _imem01_rd = 1;
    13: _imem01_rd = 1;
    14: _imem01_rd = 1;
    15: _imem01_rd = 1;
    16: _imem01_rd = 1;
    17: _imem01_rd = 1;
    18: _imem01_rd = 1;
    19: _imem01_rd = 1;
    20: _imem01_rd = 1;
    21: _imem01_rd = 1;
    22: _imem01_rd = 1;
    23: _imem01_rd = 1;
    24: _imem01_rd = 1;
    25: _imem01_rd = 1;
    26: _imem01_rd = 1;
    27: _imem01_rd = 1;
    28: _imem01_rd = 1;
    29: _imem01_rd = 1;
    30: _imem01_rd = 1;
    31: _imem01_rd = 1;
    32: _imem01_rd = 1;
    33: _imem01_rd = 1;
    34: _imem01_rd = 1;
    35: _imem01_rd = 1;
    36: _imem01_rd = 1;
    37: _imem01_rd = 1;
    38: _imem01_rd = 1;
    39: _imem01_rd = 1;
    40: _imem01_rd = 1;
    41: _imem01_rd = 1;
    42: _imem01_rd = 1;
    43: _imem01_rd = 1;
    44: _imem01_rd = 1;
    45: _imem01_rd = 1;
    46: _imem01_rd = 1;
    47: _imem01_rd = 1;
    48: _imem01_rd = 1;
    49: _imem01_rd = 1;
    50: _imem01_rd = 1;
    51: _imem01_rd = 1;
    52: _imem01_rd = 1;
    53: _imem01_rd = 1;
    54: _imem01_rd = 1;
    55: _imem01_rd = 1;
    56: _imem01_rd = 1;
    57: _imem01_rd = 1;
    58: _imem01_rd = 1;
    59: _imem01_rd = 1;
    60: _imem01_rd = 1;
    61: _imem01_rd = 1;
    62: _imem01_rd = 1;
    63: _imem01_rd = 1;
    64: _imem01_rd = 1;
    65: _imem01_rd = 1;
    66: _imem01_rd = 1;
    67: _imem01_rd = 1;
    68: _imem01_rd = 1;
    69: _imem01_rd = 1;
    70: _imem01_rd = 1;
    71: _imem01_rd = 1;
    72: _imem01_rd = 1;
    73: _imem01_rd = 1;
    74: _imem01_rd = 1;
    75: _imem01_rd = 1;
    76: _imem01_rd = 1;
    77: _imem01_rd = 1;
    78: _imem01_rd = 1;
    79: _imem01_rd = 1;
    80: _imem01_rd = 1;
    81: _imem01_rd = 1;
    82: _imem01_rd = 1;
    83: _imem01_rd = 1;
    84: _imem01_rd = 1;
    85: _imem01_rd = 1;
    86: _imem01_rd = 1;
    87: _imem01_rd = 1;
    88: _imem01_rd = 1;
    89: _imem01_rd = 1;
    90: _imem01_rd = 1;
    91: _imem01_rd = 1;
    92: _imem01_rd = 1;
    93: _imem01_rd = 1;
    94: _imem01_rd = 1;
    95: _imem01_rd = 1;
    default: _imem01_rd = 0;
    endcase
  end // always @ ( * )
  assign imem01_rd = _imem01_rd;

  // 2番目の入力用メモリブロックの制御
  reg [1:0] _imem02_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem02_bank = 0;
    2: _imem02_bank = 1;
    1: _imem02_bank = 2;
    0: _imem02_bank = 3;
    4: _imem02_bank = 0;
    5: _imem02_bank = 0;
    6: _imem02_bank = 0;
    7: _imem02_bank = 0;
    8: _imem02_bank = 0;
    9: _imem02_bank = 0;
    10: _imem02_bank = 0;
    11: _imem02_bank = 0;
    12: _imem02_bank = 0;
    13: _imem02_bank = 0;
    14: _imem02_bank = 0;
    15: _imem02_bank = 0;
    16: _imem02_bank = 0;
    17: _imem02_bank = 0;
    18: _imem02_bank = 0;
    19: _imem02_bank = 3;
    20: _imem02_bank = 0;
    21: _imem02_bank = 0;
    22: _imem02_bank = 0;
    23: _imem02_bank = 0;
    24: _imem02_bank = 2;
    25: _imem02_bank = 0;
    26: _imem02_bank = 0;
    27: _imem02_bank = 0;
    28: _imem02_bank = 0;
    29: _imem02_bank = 0;
    30: _imem02_bank = 0;
    31: _imem02_bank = 0;
    32: _imem02_bank = 0;
    33: _imem02_bank = 0;
    34: _imem02_bank = 0;
    35: _imem02_bank = 0;
    36: _imem02_bank = 0;
    37: _imem02_bank = 0;
    38: _imem02_bank = 0;
    39: _imem02_bank = 0;
    40: _imem02_bank = 0;
    41: _imem02_bank = 0;
    42: _imem02_bank = 0;
    43: _imem02_bank = 1;
    44: _imem02_bank = 0;
    45: _imem02_bank = 0;
    46: _imem02_bank = 0;
    47: _imem02_bank = 0;
    48: _imem02_bank = 0;
    49: _imem02_bank = 0;
    50: _imem02_bank = 2;
    51: _imem02_bank = 0;
    52: _imem02_bank = 0;
    53: _imem02_bank = 0;
    54: _imem02_bank = 0;
    55: _imem02_bank = 0;
    56: _imem02_bank = 0;
    57: _imem02_bank = 0;
    58: _imem02_bank = 0;
    59: _imem02_bank = 0;
    60: _imem02_bank = 0;
    61: _imem02_bank = 1;
    62: _imem02_bank = 0;
    63: _imem02_bank = 0;
    64: _imem02_bank = 0;
    65: _imem02_bank = 0;
    66: _imem02_bank = 0;
    67: _imem02_bank = 0;
    68: _imem02_bank = 0;
    69: _imem02_bank = 0;
    70: _imem02_bank = 1;
    71: _imem02_bank = 0;
    72: _imem02_bank = 0;
    73: _imem02_bank = 0;
    74: _imem02_bank = 0;
    75: _imem02_bank = 0;
    76: _imem02_bank = 0;
    77: _imem02_bank = 0;
    78: _imem02_bank = 0;
    79: _imem02_bank = 0;
    80: _imem02_bank = 0;
    81: _imem02_bank = 0;
    82: _imem02_bank = 1;
    83: _imem02_bank = 3;
    84: _imem02_bank = 0;
    85: _imem02_bank = 0;
    86: _imem02_bank = 0;
    87: _imem02_bank = 0;
    88: _imem02_bank = 0;
    89: _imem02_bank = 0;
    90: _imem02_bank = 0;
    91: _imem02_bank = 0;
    92: _imem02_bank = 0;
    93: _imem02_bank = 0;
    94: _imem02_bank = 0;
    95: _imem02_bank = 0;
    default: _imem02_bank = 0;
    endcase
  end // always @ ( * )
  assign imem02_bank = _imem02_bank;
  reg _imem02_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem02_rd = 1;
    2: _imem02_rd = 1;
    1: _imem02_rd = 1;
    0: _imem02_rd = 1;
    4: _imem02_rd = 1;
    5: _imem02_rd = 1;
    6: _imem02_rd = 1;
    7: _imem02_rd = 1;
    8: _imem02_rd = 1;
    9: _imem02_rd = 1;
    10: _imem02_rd = 1;
    11: _imem02_rd = 1;
    12: _imem02_rd = 1;
    13: _imem02_rd = 1;
    14: _imem02_rd = 1;
    15: _imem02_rd = 1;
    16: _imem02_rd = 1;
    17: _imem02_rd = 1;
    18: _imem02_rd = 1;
    19: _imem02_rd = 1;
    20: _imem02_rd = 1;
    21: _imem02_rd = 1;
    22: _imem02_rd = 1;
    23: _imem02_rd = 1;
    24: _imem02_rd = 1;
    25: _imem02_rd = 1;
    26: _imem02_rd = 1;
    27: _imem02_rd = 1;
    28: _imem02_rd = 1;
    29: _imem02_rd = 1;
    30: _imem02_rd = 1;
    31: _imem02_rd = 1;
    32: _imem02_rd = 1;
    33: _imem02_rd = 1;
    34: _imem02_rd = 1;
    35: _imem02_rd = 1;
    36: _imem02_rd = 1;
    37: _imem02_rd = 1;
    38: _imem02_rd = 1;
    39: _imem02_rd = 1;
    40: _imem02_rd = 1;
    41: _imem02_rd = 1;
    42: _imem02_rd = 1;
    43: _imem02_rd = 1;
    44: _imem02_rd = 1;
    45: _imem02_rd = 1;
    46: _imem02_rd = 1;
    47: _imem02_rd = 1;
    48: _imem02_rd = 1;
    49: _imem02_rd = 1;
    50: _imem02_rd = 1;
    51: _imem02_rd = 1;
    52: _imem02_rd = 1;
    53: _imem02_rd = 1;
    54: _imem02_rd = 1;
    55: _imem02_rd = 1;
    56: _imem02_rd = 1;
    57: _imem02_rd = 1;
    58: _imem02_rd = 1;
    59: _imem02_rd = 1;
    60: _imem02_rd = 1;
    61: _imem02_rd = 1;
    62: _imem02_rd = 1;
    63: _imem02_rd = 1;
    64: _imem02_rd = 1;
    65: _imem02_rd = 1;
    66: _imem02_rd = 1;
    67: _imem02_rd = 1;
    68: _imem02_rd = 1;
    69: _imem02_rd = 1;
    70: _imem02_rd = 1;
    71: _imem02_rd = 1;
    72: _imem02_rd = 1;
    73: _imem02_rd = 1;
    74: _imem02_rd = 1;
    75: _imem02_rd = 1;
    76: _imem02_rd = 1;
    77: _imem02_rd = 1;
    78: _imem02_rd = 1;
    79: _imem02_rd = 1;
    80: _imem02_rd = 1;
    81: _imem02_rd = 1;
    82: _imem02_rd = 1;
    83: _imem02_rd = 1;
    84: _imem02_rd = 1;
    85: _imem02_rd = 1;
    86: _imem02_rd = 1;
    87: _imem02_rd = 1;
    88: _imem02_rd = 1;
    89: _imem02_rd = 1;
    90: _imem02_rd = 1;
    91: _imem02_rd = 1;
    92: _imem02_rd = 1;
    93: _imem02_rd = 1;
    94: _imem02_rd = 1;
    95: _imem02_rd = 1;
    default: _imem02_rd = 0;
    endcase
  end // always @ ( * )
  assign imem02_rd = _imem02_rd;

  // 3番目の入力用メモリブロックの制御
  reg [1:0] _imem03_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem03_bank = 0;
    2: _imem03_bank = 1;
    1: _imem03_bank = 2;
    0: _imem03_bank = 3;
    4: _imem03_bank = 3;
    5: _imem03_bank = 0;
    6: _imem03_bank = 0;
    7: _imem03_bank = 0;
    8: _imem03_bank = 0;
    9: _imem03_bank = 0;
    10: _imem03_bank = 0;
    11: _imem03_bank = 0;
    12: _imem03_bank = 0;
    13: _imem03_bank = 0;
    14: _imem03_bank = 0;
    15: _imem03_bank = 0;
    16: _imem03_bank = 0;
    17: _imem03_bank = 0;
    18: _imem03_bank = 0;
    19: _imem03_bank = 0;
    20: _imem03_bank = 0;
    21: _imem03_bank = 0;
    22: _imem03_bank = 0;
    23: _imem03_bank = 0;
    24: _imem03_bank = 0;
    25: _imem03_bank = 0;
    26: _imem03_bank = 2;
    27: _imem03_bank = 0;
    28: _imem03_bank = 0;
    29: _imem03_bank = 1;
    30: _imem03_bank = 0;
    31: _imem03_bank = 0;
    32: _imem03_bank = 0;
    33: _imem03_bank = 0;
    34: _imem03_bank = 0;
    35: _imem03_bank = 0;
    36: _imem03_bank = 0;
    37: _imem03_bank = 0;
    38: _imem03_bank = 0;
    39: _imem03_bank = 0;
    40: _imem03_bank = 0;
    41: _imem03_bank = 0;
    42: _imem03_bank = 0;
    43: _imem03_bank = 0;
    44: _imem03_bank = 0;
    45: _imem03_bank = 0;
    46: _imem03_bank = 0;
    47: _imem03_bank = 0;
    48: _imem03_bank = 0;
    49: _imem03_bank = 0;
    50: _imem03_bank = 0;
    51: _imem03_bank = 0;
    52: _imem03_bank = 1;
    53: _imem03_bank = 1;
    54: _imem03_bank = 0;
    55: _imem03_bank = 0;
    56: _imem03_bank = 0;
    57: _imem03_bank = 0;
    58: _imem03_bank = 0;
    59: _imem03_bank = 0;
    60: _imem03_bank = 0;
    61: _imem03_bank = 0;
    62: _imem03_bank = 0;
    63: _imem03_bank = 0;
    64: _imem03_bank = 0;
    65: _imem03_bank = 0;
    66: _imem03_bank = 0;
    67: _imem03_bank = 0;
    68: _imem03_bank = 2;
    69: _imem03_bank = 0;
    70: _imem03_bank = 0;
    71: _imem03_bank = 0;
    72: _imem03_bank = 0;
    73: _imem03_bank = 0;
    74: _imem03_bank = 0;
    75: _imem03_bank = 0;
    76: _imem03_bank = 0;
    77: _imem03_bank = 0;
    78: _imem03_bank = 0;
    79: _imem03_bank = 0;
    80: _imem03_bank = 0;
    81: _imem03_bank = 0;
    82: _imem03_bank = 0;
    83: _imem03_bank = 0;
    84: _imem03_bank = 0;
    85: _imem03_bank = 0;
    86: _imem03_bank = 1;
    87: _imem03_bank = 0;
    88: _imem03_bank = 3;
    89: _imem03_bank = 0;
    90: _imem03_bank = 0;
    91: _imem03_bank = 0;
    92: _imem03_bank = 0;
    93: _imem03_bank = 0;
    94: _imem03_bank = 0;
    95: _imem03_bank = 0;
    default: _imem03_bank = 0;
    endcase
  end // always @ ( * )
  assign imem03_bank = _imem03_bank;
  reg _imem03_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem03_rd = 1;
    2: _imem03_rd = 1;
    1: _imem03_rd = 1;
    0: _imem03_rd = 1;
    4: _imem03_rd = 1;
    5: _imem03_rd = 1;
    6: _imem03_rd = 1;
    7: _imem03_rd = 1;
    8: _imem03_rd = 1;
    9: _imem03_rd = 1;
    10: _imem03_rd = 1;
    11: _imem03_rd = 1;
    12: _imem03_rd = 1;
    13: _imem03_rd = 1;
    14: _imem03_rd = 1;
    15: _imem03_rd = 1;
    16: _imem03_rd = 1;
    17: _imem03_rd = 1;
    18: _imem03_rd = 1;
    19: _imem03_rd = 1;
    20: _imem03_rd = 1;
    21: _imem03_rd = 1;
    22: _imem03_rd = 1;
    23: _imem03_rd = 1;
    24: _imem03_rd = 1;
    25: _imem03_rd = 1;
    26: _imem03_rd = 1;
    27: _imem03_rd = 1;
    28: _imem03_rd = 1;
    29: _imem03_rd = 1;
    30: _imem03_rd = 1;
    31: _imem03_rd = 1;
    32: _imem03_rd = 1;
    33: _imem03_rd = 1;
    34: _imem03_rd = 1;
    35: _imem03_rd = 1;
    36: _imem03_rd = 1;
    37: _imem03_rd = 1;
    38: _imem03_rd = 1;
    39: _imem03_rd = 1;
    40: _imem03_rd = 1;
    41: _imem03_rd = 1;
    42: _imem03_rd = 1;
    43: _imem03_rd = 1;
    44: _imem03_rd = 1;
    45: _imem03_rd = 1;
    46: _imem03_rd = 1;
    47: _imem03_rd = 1;
    48: _imem03_rd = 1;
    49: _imem03_rd = 1;
    50: _imem03_rd = 1;
    51: _imem03_rd = 1;
    52: _imem03_rd = 1;
    53: _imem03_rd = 1;
    54: _imem03_rd = 1;
    55: _imem03_rd = 1;
    56: _imem03_rd = 1;
    57: _imem03_rd = 1;
    58: _imem03_rd = 1;
    59: _imem03_rd = 1;
    60: _imem03_rd = 1;
    61: _imem03_rd = 1;
    62: _imem03_rd = 1;
    63: _imem03_rd = 1;
    64: _imem03_rd = 1;
    65: _imem03_rd = 1;
    66: _imem03_rd = 1;
    67: _imem03_rd = 1;
    68: _imem03_rd = 1;
    69: _imem03_rd = 1;
    70: _imem03_rd = 1;
    71: _imem03_rd = 1;
    72: _imem03_rd = 1;
    73: _imem03_rd = 1;
    74: _imem03_rd = 1;
    75: _imem03_rd = 1;
    76: _imem03_rd = 1;
    77: _imem03_rd = 1;
    78: _imem03_rd = 1;
    79: _imem03_rd = 1;
    80: _imem03_rd = 1;
    81: _imem03_rd = 1;
    82: _imem03_rd = 1;
    83: _imem03_rd = 1;
    84: _imem03_rd = 1;
    85: _imem03_rd = 1;
    86: _imem03_rd = 1;
    87: _imem03_rd = 1;
    88: _imem03_rd = 1;
    89: _imem03_rd = 1;
    90: _imem03_rd = 1;
    91: _imem03_rd = 1;
    92: _imem03_rd = 1;
    93: _imem03_rd = 1;
    94: _imem03_rd = 1;
    95: _imem03_rd = 1;
    default: _imem03_rd = 0;
    endcase
  end // always @ ( * )
  assign imem03_rd = _imem03_rd;

  // 4番目の入力用メモリブロックの制御
  reg [1:0] _imem04_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem04_bank = 0;
    2: _imem04_bank = 1;
    1: _imem04_bank = 2;
    0: _imem04_bank = 3;
    4: _imem04_bank = 0;
    5: _imem04_bank = 0;
    6: _imem04_bank = 0;
    7: _imem04_bank = 0;
    8: _imem04_bank = 0;
    9: _imem04_bank = 0;
    10: _imem04_bank = 0;
    11: _imem04_bank = 0;
    12: _imem04_bank = 0;
    13: _imem04_bank = 0;
    14: _imem04_bank = 0;
    15: _imem04_bank = 0;
    16: _imem04_bank = 3;
    17: _imem04_bank = 2;
    18: _imem04_bank = 0;
    19: _imem04_bank = 0;
    20: _imem04_bank = 1;
    21: _imem04_bank = 0;
    22: _imem04_bank = 1;
    23: _imem04_bank = 0;
    24: _imem04_bank = 0;
    25: _imem04_bank = 0;
    26: _imem04_bank = 0;
    27: _imem04_bank = 0;
    28: _imem04_bank = 0;
    29: _imem04_bank = 0;
    30: _imem04_bank = 0;
    31: _imem04_bank = 0;
    32: _imem04_bank = 0;
    33: _imem04_bank = 0;
    34: _imem04_bank = 0;
    35: _imem04_bank = 0;
    36: _imem04_bank = 0;
    37: _imem04_bank = 0;
    38: _imem04_bank = 0;
    39: _imem04_bank = 0;
    40: _imem04_bank = 2;
    41: _imem04_bank = 0;
    42: _imem04_bank = 0;
    43: _imem04_bank = 0;
    44: _imem04_bank = 3;
    45: _imem04_bank = 0;
    46: _imem04_bank = 0;
    47: _imem04_bank = 3;
    48: _imem04_bank = 0;
    49: _imem04_bank = 0;
    50: _imem04_bank = 0;
    51: _imem04_bank = 0;
    52: _imem04_bank = 0;
    53: _imem04_bank = 0;
    54: _imem04_bank = 0;
    55: _imem04_bank = 0;
    56: _imem04_bank = 0;
    57: _imem04_bank = 3;
    58: _imem04_bank = 0;
    59: _imem04_bank = 0;
    60: _imem04_bank = 0;
    61: _imem04_bank = 0;
    62: _imem04_bank = 0;
    63: _imem04_bank = 0;
    64: _imem04_bank = 0;
    65: _imem04_bank = 0;
    66: _imem04_bank = 0;
    67: _imem04_bank = 0;
    68: _imem04_bank = 0;
    69: _imem04_bank = 0;
    70: _imem04_bank = 0;
    71: _imem04_bank = 0;
    72: _imem04_bank = 0;
    73: _imem04_bank = 0;
    74: _imem04_bank = 0;
    75: _imem04_bank = 0;
    76: _imem04_bank = 0;
    77: _imem04_bank = 0;
    78: _imem04_bank = 0;
    79: _imem04_bank = 0;
    80: _imem04_bank = 0;
    81: _imem04_bank = 1;
    82: _imem04_bank = 0;
    83: _imem04_bank = 0;
    84: _imem04_bank = 0;
    85: _imem04_bank = 0;
    86: _imem04_bank = 0;
    87: _imem04_bank = 0;
    88: _imem04_bank = 0;
    89: _imem04_bank = 0;
    90: _imem04_bank = 0;
    91: _imem04_bank = 0;
    92: _imem04_bank = 0;
    93: _imem04_bank = 0;
    94: _imem04_bank = 0;
    95: _imem04_bank = 0;
    default: _imem04_bank = 0;
    endcase
  end // always @ ( * )
  assign imem04_bank = _imem04_bank;
  reg _imem04_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem04_rd = 1;
    2: _imem04_rd = 1;
    1: _imem04_rd = 1;
    0: _imem04_rd = 1;
    4: _imem04_rd = 1;
    5: _imem04_rd = 1;
    6: _imem04_rd = 1;
    7: _imem04_rd = 1;
    8: _imem04_rd = 1;
    9: _imem04_rd = 1;
    10: _imem04_rd = 1;
    11: _imem04_rd = 1;
    12: _imem04_rd = 1;
    13: _imem04_rd = 1;
    14: _imem04_rd = 1;
    15: _imem04_rd = 1;
    16: _imem04_rd = 1;
    17: _imem04_rd = 1;
    18: _imem04_rd = 1;
    19: _imem04_rd = 1;
    20: _imem04_rd = 1;
    21: _imem04_rd = 1;
    22: _imem04_rd = 1;
    23: _imem04_rd = 1;
    24: _imem04_rd = 1;
    25: _imem04_rd = 1;
    26: _imem04_rd = 1;
    27: _imem04_rd = 1;
    28: _imem04_rd = 1;
    29: _imem04_rd = 1;
    30: _imem04_rd = 1;
    31: _imem04_rd = 1;
    32: _imem04_rd = 1;
    33: _imem04_rd = 1;
    34: _imem04_rd = 1;
    35: _imem04_rd = 1;
    36: _imem04_rd = 1;
    37: _imem04_rd = 1;
    38: _imem04_rd = 1;
    39: _imem04_rd = 1;
    40: _imem04_rd = 1;
    41: _imem04_rd = 1;
    42: _imem04_rd = 1;
    43: _imem04_rd = 1;
    44: _imem04_rd = 1;
    45: _imem04_rd = 1;
    46: _imem04_rd = 1;
    47: _imem04_rd = 1;
    48: _imem04_rd = 1;
    49: _imem04_rd = 1;
    50: _imem04_rd = 1;
    51: _imem04_rd = 1;
    52: _imem04_rd = 1;
    53: _imem04_rd = 1;
    54: _imem04_rd = 1;
    55: _imem04_rd = 1;
    56: _imem04_rd = 1;
    57: _imem04_rd = 1;
    58: _imem04_rd = 1;
    59: _imem04_rd = 1;
    60: _imem04_rd = 1;
    61: _imem04_rd = 1;
    62: _imem04_rd = 1;
    63: _imem04_rd = 1;
    64: _imem04_rd = 1;
    65: _imem04_rd = 1;
    66: _imem04_rd = 1;
    67: _imem04_rd = 1;
    68: _imem04_rd = 1;
    69: _imem04_rd = 1;
    70: _imem04_rd = 1;
    71: _imem04_rd = 1;
    72: _imem04_rd = 1;
    73: _imem04_rd = 1;
    74: _imem04_rd = 1;
    75: _imem04_rd = 1;
    76: _imem04_rd = 1;
    77: _imem04_rd = 1;
    78: _imem04_rd = 1;
    79: _imem04_rd = 1;
    80: _imem04_rd = 1;
    81: _imem04_rd = 1;
    82: _imem04_rd = 1;
    83: _imem04_rd = 1;
    84: _imem04_rd = 1;
    85: _imem04_rd = 1;
    86: _imem04_rd = 1;
    87: _imem04_rd = 1;
    88: _imem04_rd = 1;
    89: _imem04_rd = 1;
    90: _imem04_rd = 1;
    91: _imem04_rd = 1;
    92: _imem04_rd = 1;
    93: _imem04_rd = 1;
    94: _imem04_rd = 1;
    95: _imem04_rd = 1;
    default: _imem04_rd = 0;
    endcase
  end // always @ ( * )
  assign imem04_rd = _imem04_rd;

  // 5番目の入力用メモリブロックの制御
  reg [1:0] _imem05_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem05_bank = 0;
    2: _imem05_bank = 1;
    1: _imem05_bank = 2;
    0: _imem05_bank = 3;
    4: _imem05_bank = 1;
    5: _imem05_bank = 0;
    6: _imem05_bank = 0;
    7: _imem05_bank = 0;
    8: _imem05_bank = 0;
    9: _imem05_bank = 0;
    10: _imem05_bank = 2;
    11: _imem05_bank = 0;
    12: _imem05_bank = 0;
    13: _imem05_bank = 0;
    14: _imem05_bank = 0;
    15: _imem05_bank = 0;
    16: _imem05_bank = 0;
    17: _imem05_bank = 0;
    18: _imem05_bank = 2;
    19: _imem05_bank = 0;
    20: _imem05_bank = 0;
    21: _imem05_bank = 0;
    22: _imem05_bank = 0;
    23: _imem05_bank = 0;
    24: _imem05_bank = 0;
    25: _imem05_bank = 0;
    26: _imem05_bank = 0;
    27: _imem05_bank = 0;
    28: _imem05_bank = 0;
    29: _imem05_bank = 0;
    30: _imem05_bank = 0;
    31: _imem05_bank = 0;
    32: _imem05_bank = 0;
    33: _imem05_bank = 0;
    34: _imem05_bank = 0;
    35: _imem05_bank = 0;
    36: _imem05_bank = 0;
    37: _imem05_bank = 0;
    38: _imem05_bank = 0;
    39: _imem05_bank = 0;
    40: _imem05_bank = 0;
    41: _imem05_bank = 0;
    42: _imem05_bank = 0;
    43: _imem05_bank = 0;
    44: _imem05_bank = 0;
    45: _imem05_bank = 0;
    46: _imem05_bank = 0;
    47: _imem05_bank = 0;
    48: _imem05_bank = 2;
    49: _imem05_bank = 0;
    50: _imem05_bank = 0;
    51: _imem05_bank = 0;
    52: _imem05_bank = 0;
    53: _imem05_bank = 0;
    54: _imem05_bank = 1;
    55: _imem05_bank = 0;
    56: _imem05_bank = 0;
    57: _imem05_bank = 0;
    58: _imem05_bank = 0;
    59: _imem05_bank = 1;
    60: _imem05_bank = 0;
    61: _imem05_bank = 0;
    62: _imem05_bank = 0;
    63: _imem05_bank = 1;
    64: _imem05_bank = 2;
    65: _imem05_bank = 0;
    66: _imem05_bank = 1;
    67: _imem05_bank = 0;
    68: _imem05_bank = 0;
    69: _imem05_bank = 0;
    70: _imem05_bank = 0;
    71: _imem05_bank = 1;
    72: _imem05_bank = 3;
    73: _imem05_bank = 0;
    74: _imem05_bank = 0;
    75: _imem05_bank = 0;
    76: _imem05_bank = 0;
    77: _imem05_bank = 2;
    78: _imem05_bank = 0;
    79: _imem05_bank = 0;
    80: _imem05_bank = 0;
    81: _imem05_bank = 0;
    82: _imem05_bank = 0;
    83: _imem05_bank = 0;
    84: _imem05_bank = 0;
    85: _imem05_bank = 2;
    86: _imem05_bank = 0;
    87: _imem05_bank = 0;
    88: _imem05_bank = 0;
    89: _imem05_bank = 0;
    90: _imem05_bank = 0;
    91: _imem05_bank = 0;
    92: _imem05_bank = 0;
    93: _imem05_bank = 0;
    94: _imem05_bank = 0;
    95: _imem05_bank = 0;
    default: _imem05_bank = 0;
    endcase
  end // always @ ( * )
  assign imem05_bank = _imem05_bank;
  reg _imem05_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem05_rd = 1;
    2: _imem05_rd = 1;
    1: _imem05_rd = 1;
    0: _imem05_rd = 1;
    4: _imem05_rd = 1;
    5: _imem05_rd = 1;
    6: _imem05_rd = 1;
    7: _imem05_rd = 1;
    8: _imem05_rd = 1;
    9: _imem05_rd = 1;
    10: _imem05_rd = 1;
    11: _imem05_rd = 1;
    12: _imem05_rd = 1;
    13: _imem05_rd = 1;
    14: _imem05_rd = 1;
    15: _imem05_rd = 1;
    16: _imem05_rd = 1;
    17: _imem05_rd = 1;
    18: _imem05_rd = 1;
    19: _imem05_rd = 1;
    20: _imem05_rd = 1;
    21: _imem05_rd = 1;
    22: _imem05_rd = 1;
    23: _imem05_rd = 1;
    24: _imem05_rd = 1;
    25: _imem05_rd = 1;
    26: _imem05_rd = 1;
    27: _imem05_rd = 1;
    28: _imem05_rd = 1;
    29: _imem05_rd = 1;
    30: _imem05_rd = 1;
    31: _imem05_rd = 1;
    32: _imem05_rd = 1;
    33: _imem05_rd = 1;
    34: _imem05_rd = 1;
    35: _imem05_rd = 1;
    36: _imem05_rd = 1;
    37: _imem05_rd = 1;
    38: _imem05_rd = 1;
    39: _imem05_rd = 1;
    40: _imem05_rd = 1;
    41: _imem05_rd = 1;
    42: _imem05_rd = 1;
    43: _imem05_rd = 1;
    44: _imem05_rd = 1;
    45: _imem05_rd = 1;
    46: _imem05_rd = 1;
    47: _imem05_rd = 1;
    48: _imem05_rd = 1;
    49: _imem05_rd = 1;
    50: _imem05_rd = 1;
    51: _imem05_rd = 1;
    52: _imem05_rd = 1;
    53: _imem05_rd = 1;
    54: _imem05_rd = 1;
    55: _imem05_rd = 1;
    56: _imem05_rd = 1;
    57: _imem05_rd = 1;
    58: _imem05_rd = 1;
    59: _imem05_rd = 1;
    60: _imem05_rd = 1;
    61: _imem05_rd = 1;
    62: _imem05_rd = 1;
    63: _imem05_rd = 1;
    64: _imem05_rd = 1;
    65: _imem05_rd = 1;
    66: _imem05_rd = 1;
    67: _imem05_rd = 1;
    68: _imem05_rd = 1;
    69: _imem05_rd = 1;
    70: _imem05_rd = 1;
    71: _imem05_rd = 1;
    72: _imem05_rd = 1;
    73: _imem05_rd = 1;
    74: _imem05_rd = 1;
    75: _imem05_rd = 1;
    76: _imem05_rd = 1;
    77: _imem05_rd = 1;
    78: _imem05_rd = 1;
    79: _imem05_rd = 1;
    80: _imem05_rd = 1;
    81: _imem05_rd = 1;
    82: _imem05_rd = 1;
    83: _imem05_rd = 1;
    84: _imem05_rd = 1;
    85: _imem05_rd = 1;
    86: _imem05_rd = 1;
    87: _imem05_rd = 1;
    88: _imem05_rd = 1;
    89: _imem05_rd = 1;
    90: _imem05_rd = 1;
    91: _imem05_rd = 1;
    92: _imem05_rd = 1;
    93: _imem05_rd = 1;
    94: _imem05_rd = 1;
    95: _imem05_rd = 1;
    default: _imem05_rd = 0;
    endcase
  end // always @ ( * )
  assign imem05_rd = _imem05_rd;

  // 6番目の入力用メモリブロックの制御
  reg [1:0] _imem06_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem06_bank = 0;
    2: _imem06_bank = 1;
    1: _imem06_bank = 2;
    0: _imem06_bank = 3;
    4: _imem06_bank = 0;
    5: _imem06_bank = 0;
    6: _imem06_bank = 0;
    7: _imem06_bank = 3;
    8: _imem06_bank = 0;
    9: _imem06_bank = 0;
    10: _imem06_bank = 0;
    11: _imem06_bank = 0;
    12: _imem06_bank = 0;
    13: _imem06_bank = 0;
    14: _imem06_bank = 0;
    15: _imem06_bank = 0;
    16: _imem06_bank = 0;
    17: _imem06_bank = 0;
    18: _imem06_bank = 0;
    19: _imem06_bank = 0;
    20: _imem06_bank = 0;
    21: _imem06_bank = 0;
    22: _imem06_bank = 0;
    23: _imem06_bank = 0;
    24: _imem06_bank = 0;
    25: _imem06_bank = 0;
    26: _imem06_bank = 0;
    27: _imem06_bank = 2;
    28: _imem06_bank = 0;
    29: _imem06_bank = 0;
    30: _imem06_bank = 3;
    31: _imem06_bank = 0;
    32: _imem06_bank = 0;
    33: _imem06_bank = 0;
    34: _imem06_bank = 1;
    35: _imem06_bank = 3;
    36: _imem06_bank = 0;
    37: _imem06_bank = 1;
    38: _imem06_bank = 0;
    39: _imem06_bank = 0;
    40: _imem06_bank = 0;
    41: _imem06_bank = 0;
    42: _imem06_bank = 0;
    43: _imem06_bank = 0;
    44: _imem06_bank = 0;
    45: _imem06_bank = 0;
    46: _imem06_bank = 0;
    47: _imem06_bank = 0;
    48: _imem06_bank = 0;
    49: _imem06_bank = 0;
    50: _imem06_bank = 0;
    51: _imem06_bank = 0;
    52: _imem06_bank = 0;
    53: _imem06_bank = 0;
    54: _imem06_bank = 0;
    55: _imem06_bank = 1;
    56: _imem06_bank = 2;
    57: _imem06_bank = 0;
    58: _imem06_bank = 0;
    59: _imem06_bank = 3;
    60: _imem06_bank = 0;
    61: _imem06_bank = 0;
    62: _imem06_bank = 0;
    63: _imem06_bank = 0;
    64: _imem06_bank = 0;
    65: _imem06_bank = 0;
    66: _imem06_bank = 0;
    67: _imem06_bank = 0;
    68: _imem06_bank = 0;
    69: _imem06_bank = 3;
    70: _imem06_bank = 0;
    71: _imem06_bank = 0;
    72: _imem06_bank = 0;
    73: _imem06_bank = 0;
    74: _imem06_bank = 0;
    75: _imem06_bank = 0;
    76: _imem06_bank = 0;
    77: _imem06_bank = 0;
    78: _imem06_bank = 0;
    79: _imem06_bank = 0;
    80: _imem06_bank = 0;
    81: _imem06_bank = 0;
    82: _imem06_bank = 0;
    83: _imem06_bank = 0;
    84: _imem06_bank = 2;
    85: _imem06_bank = 0;
    86: _imem06_bank = 0;
    87: _imem06_bank = 3;
    88: _imem06_bank = 0;
    89: _imem06_bank = 0;
    90: _imem06_bank = 0;
    91: _imem06_bank = 0;
    92: _imem06_bank = 0;
    93: _imem06_bank = 0;
    94: _imem06_bank = 0;
    95: _imem06_bank = 0;
    default: _imem06_bank = 0;
    endcase
  end // always @ ( * )
  assign imem06_bank = _imem06_bank;
  reg _imem06_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem06_rd = 1;
    2: _imem06_rd = 1;
    1: _imem06_rd = 1;
    0: _imem06_rd = 1;
    4: _imem06_rd = 1;
    5: _imem06_rd = 1;
    6: _imem06_rd = 1;
    7: _imem06_rd = 1;
    8: _imem06_rd = 1;
    9: _imem06_rd = 1;
    10: _imem06_rd = 1;
    11: _imem06_rd = 1;
    12: _imem06_rd = 1;
    13: _imem06_rd = 1;
    14: _imem06_rd = 1;
    15: _imem06_rd = 1;
    16: _imem06_rd = 1;
    17: _imem06_rd = 1;
    18: _imem06_rd = 1;
    19: _imem06_rd = 1;
    20: _imem06_rd = 1;
    21: _imem06_rd = 1;
    22: _imem06_rd = 1;
    23: _imem06_rd = 1;
    24: _imem06_rd = 1;
    25: _imem06_rd = 1;
    26: _imem06_rd = 1;
    27: _imem06_rd = 1;
    28: _imem06_rd = 1;
    29: _imem06_rd = 1;
    30: _imem06_rd = 1;
    31: _imem06_rd = 1;
    32: _imem06_rd = 1;
    33: _imem06_rd = 1;
    34: _imem06_rd = 1;
    35: _imem06_rd = 1;
    36: _imem06_rd = 1;
    37: _imem06_rd = 1;
    38: _imem06_rd = 1;
    39: _imem06_rd = 1;
    40: _imem06_rd = 1;
    41: _imem06_rd = 1;
    42: _imem06_rd = 1;
    43: _imem06_rd = 1;
    44: _imem06_rd = 1;
    45: _imem06_rd = 1;
    46: _imem06_rd = 1;
    47: _imem06_rd = 1;
    48: _imem06_rd = 1;
    49: _imem06_rd = 1;
    50: _imem06_rd = 1;
    51: _imem06_rd = 1;
    52: _imem06_rd = 1;
    53: _imem06_rd = 1;
    54: _imem06_rd = 1;
    55: _imem06_rd = 1;
    56: _imem06_rd = 1;
    57: _imem06_rd = 1;
    58: _imem06_rd = 1;
    59: _imem06_rd = 1;
    60: _imem06_rd = 1;
    61: _imem06_rd = 1;
    62: _imem06_rd = 1;
    63: _imem06_rd = 1;
    64: _imem06_rd = 1;
    65: _imem06_rd = 1;
    66: _imem06_rd = 1;
    67: _imem06_rd = 1;
    68: _imem06_rd = 1;
    69: _imem06_rd = 1;
    70: _imem06_rd = 1;
    71: _imem06_rd = 1;
    72: _imem06_rd = 1;
    73: _imem06_rd = 1;
    74: _imem06_rd = 1;
    75: _imem06_rd = 1;
    76: _imem06_rd = 1;
    77: _imem06_rd = 1;
    78: _imem06_rd = 1;
    79: _imem06_rd = 1;
    80: _imem06_rd = 1;
    81: _imem06_rd = 1;
    82: _imem06_rd = 1;
    83: _imem06_rd = 1;
    84: _imem06_rd = 1;
    85: _imem06_rd = 1;
    86: _imem06_rd = 1;
    87: _imem06_rd = 1;
    88: _imem06_rd = 1;
    89: _imem06_rd = 1;
    90: _imem06_rd = 1;
    91: _imem06_rd = 1;
    92: _imem06_rd = 1;
    93: _imem06_rd = 1;
    94: _imem06_rd = 1;
    95: _imem06_rd = 1;
    default: _imem06_rd = 0;
    endcase
  end // always @ ( * )
  assign imem06_rd = _imem06_rd;

  // 7番目の入力用メモリブロックの制御
  reg [1:0] _imem07_bank;
  always @ ( * ) begin
    case ( state )
    3: _imem07_bank = 0;
    2: _imem07_bank = 1;
    1: _imem07_bank = 2;
    0: _imem07_bank = 3;
    4: _imem07_bank = 0;
    5: _imem07_bank = 0;
    6: _imem07_bank = 0;
    7: _imem07_bank = 0;
    8: _imem07_bank = 0;
    9: _imem07_bank = 0;
    10: _imem07_bank = 0;
    11: _imem07_bank = 0;
    12: _imem07_bank = 0;
    13: _imem07_bank = 0;
    14: _imem07_bank = 0;
    15: _imem07_bank = 0;
    16: _imem07_bank = 0;
    17: _imem07_bank = 0;
    18: _imem07_bank = 0;
    19: _imem07_bank = 0;
    20: _imem07_bank = 0;
    21: _imem07_bank = 0;
    22: _imem07_bank = 0;
    23: _imem07_bank = 0;
    24: _imem07_bank = 0;
    25: _imem07_bank = 0;
    26: _imem07_bank = 0;
    27: _imem07_bank = 0;
    28: _imem07_bank = 0;
    29: _imem07_bank = 0;
    30: _imem07_bank = 0;
    31: _imem07_bank = 0;
    32: _imem07_bank = 0;
    33: _imem07_bank = 0;
    34: _imem07_bank = 0;
    35: _imem07_bank = 0;
    36: _imem07_bank = 0;
    37: _imem07_bank = 0;
    38: _imem07_bank = 0;
    39: _imem07_bank = 0;
    40: _imem07_bank = 0;
    41: _imem07_bank = 2;
    42: _imem07_bank = 0;
    43: _imem07_bank = 0;
    44: _imem07_bank = 0;
    45: _imem07_bank = 0;
    46: _imem07_bank = 0;
    47: _imem07_bank = 0;
    48: _imem07_bank = 0;
    49: _imem07_bank = 0;
    50: _imem07_bank = 0;
    51: _imem07_bank = 0;
    52: _imem07_bank = 0;
    53: _imem07_bank = 0;
    54: _imem07_bank = 0;
    55: _imem07_bank = 0;
    56: _imem07_bank = 0;
    57: _imem07_bank = 0;
    58: _imem07_bank = 0;
    59: _imem07_bank = 0;
    60: _imem07_bank = 0;
    61: _imem07_bank = 0;
    62: _imem07_bank = 0;
    63: _imem07_bank = 0;
    64: _imem07_bank = 0;
    65: _imem07_bank = 0;
    66: _imem07_bank = 0;
    67: _imem07_bank = 0;
    68: _imem07_bank = 0;
    69: _imem07_bank = 0;
    70: _imem07_bank = 0;
    71: _imem07_bank = 0;
    72: _imem07_bank = 0;
    73: _imem07_bank = 1;
    74: _imem07_bank = 0;
    75: _imem07_bank = 0;
    76: _imem07_bank = 0;
    77: _imem07_bank = 1;
    78: _imem07_bank = 0;
    79: _imem07_bank = 3;
    80: _imem07_bank = 3;
    81: _imem07_bank = 0;
    82: _imem07_bank = 0;
    83: _imem07_bank = 0;
    84: _imem07_bank = 0;
    85: _imem07_bank = 0;
    86: _imem07_bank = 0;
    87: _imem07_bank = 0;
    88: _imem07_bank = 0;
    89: _imem07_bank = 0;
    90: _imem07_bank = 0;
    91: _imem07_bank = 0;
    92: _imem07_bank = 0;
    93: _imem07_bank = 0;
    94: _imem07_bank = 0;
    95: _imem07_bank = 0;
    default: _imem07_bank = 0;
    endcase
  end // always @ ( * )
  assign imem07_bank = _imem07_bank;
  reg _imem07_rd;
  always @ ( * ) begin
    case ( state )
    3: _imem07_rd = 1;
    2: _imem07_rd = 1;
    1: _imem07_rd = 1;
    0: _imem07_rd = 1;
    4: _imem07_rd = 1;
    5: _imem07_rd = 1;
    6: _imem07_rd = 1;
    7: _imem07_rd = 1;
    8: _imem07_rd = 1;
    9: _imem07_rd = 1;
    10: _imem07_rd = 1;
    11: _imem07_rd = 1;
    12: _imem07_rd = 1;
    13: _imem07_rd = 1;
    14: _imem07_rd = 1;
    15: _imem07_rd = 1;
    16: _imem07_rd = 1;
    17: _imem07_rd = 1;
    18: _imem07_rd = 1;
    19: _imem07_rd = 1;
    20: _imem07_rd = 1;
    21: _imem07_rd = 1;
    22: _imem07_rd = 1;
    23: _imem07_rd = 1;
    24: _imem07_rd = 1;
    25: _imem07_rd = 1;
    26: _imem07_rd = 1;
    27: _imem07_rd = 1;
    28: _imem07_rd = 1;
    29: _imem07_rd = 1;
    30: _imem07_rd = 1;
    31: _imem07_rd = 1;
    32: _imem07_rd = 1;
    33: _imem07_rd = 1;
    34: _imem07_rd = 1;
    35: _imem07_rd = 1;
    36: _imem07_rd = 1;
    37: _imem07_rd = 1;
    38: _imem07_rd = 1;
    39: _imem07_rd = 1;
    40: _imem07_rd = 1;
    41: _imem07_rd = 1;
    42: _imem07_rd = 1;
    43: _imem07_rd = 1;
    44: _imem07_rd = 1;
    45: _imem07_rd = 1;
    46: _imem07_rd = 1;
    47: _imem07_rd = 1;
    48: _imem07_rd = 1;
    49: _imem07_rd = 1;
    50: _imem07_rd = 1;
    51: _imem07_rd = 1;
    52: _imem07_rd = 1;
    53: _imem07_rd = 1;
    54: _imem07_rd = 1;
    55: _imem07_rd = 1;
    56: _imem07_rd = 1;
    57: _imem07_rd = 1;
    58: _imem07_rd = 1;
    59: _imem07_rd = 1;
    60: _imem07_rd = 1;
    61: _imem07_rd = 1;
    62: _imem07_rd = 1;
    63: _imem07_rd = 1;
    64: _imem07_rd = 1;
    65: _imem07_rd = 1;
    66: _imem07_rd = 1;
    67: _imem07_rd = 1;
    68: _imem07_rd = 1;
    69: _imem07_rd = 1;
    70: _imem07_rd = 1;
    71: _imem07_rd = 1;
    72: _imem07_rd = 1;
    73: _imem07_rd = 1;
    74: _imem07_rd = 1;
    75: _imem07_rd = 1;
    76: _imem07_rd = 1;
    77: _imem07_rd = 1;
    78: _imem07_rd = 1;
    79: _imem07_rd = 1;
    80: _imem07_rd = 1;
    81: _imem07_rd = 1;
    82: _imem07_rd = 1;
    83: _imem07_rd = 1;
    84: _imem07_rd = 1;
    85: _imem07_rd = 1;
    86: _imem07_rd = 1;
    87: _imem07_rd = 1;
    88: _imem07_rd = 1;
    89: _imem07_rd = 1;
    90: _imem07_rd = 1;
    91: _imem07_rd = 1;
    92: _imem07_rd = 1;
    93: _imem07_rd = 1;
    94: _imem07_rd = 1;
    95: _imem07_rd = 1;
    default: _imem07_rd = 0;
    endcase
  end // always @ ( * )
  assign imem07_rd = _imem07_rd;

  // 0番目の出力用メモリブロックの制御
  reg [5:0] _omem00_bank;
  always @ ( * ) begin
    case ( state )
    6: _omem00_bank = 0;
    7: _omem00_bank = 1;
    8: _omem00_bank = 2;
    9: _omem00_bank = 3;
    10: _omem00_bank = 4;
    11: _omem00_bank = 5;
    12: _omem00_bank = 6;
    13: _omem00_bank = 7;
    14: _omem00_bank = 8;
    15: _omem00_bank = 9;
    16: _omem00_bank = 10;
    17: _omem00_bank = 11;
    18: _omem00_bank = 12;
    19: _omem00_bank = 13;
    20: _omem00_bank = 14;
    21: _omem00_bank = 15;
    22: _omem00_bank = 16;
    23: _omem00_bank = 17;
    24: _omem00_bank = 18;
    25: _omem00_bank = 19;
    26: _omem00_bank = 20;
    27: _omem00_bank = 21;
    28: _omem00_bank = 22;
    29: _omem00_bank = 23;
    30: _omem00_bank = 24;
    31: _omem00_bank = 25;
    32: _omem00_bank = 26;
    33: _omem00_bank = 27;
    34: _omem00_bank = 28;
    35: _omem00_bank = 29;
    36: _omem00_bank = 30;
    37: _omem00_bank = 31;
    38: _omem00_bank = 32;
    39: _omem00_bank = 33;
    40: _omem00_bank = 34;
    41: _omem00_bank = 35;
    42: _omem00_bank = 36;
    43: _omem00_bank = 37;
    44: _omem00_bank = 38;
    45: _omem00_bank = 39;
    46: _omem00_bank = 40;
    47: _omem00_bank = 41;
    48: _omem00_bank = 42;
    49: _omem00_bank = 43;
    50: _omem00_bank = 44;
    51: _omem00_bank = 45;
    52: _omem00_bank = 46;
    53: _omem00_bank = 47;
    54: _omem00_bank = 48;
    55: _omem00_bank = 49;
    56: _omem00_bank = 50;
    57: _omem00_bank = 51;
    58: _omem00_bank = 52;
    59: _omem00_bank = 53;
    60: _omem00_bank = 54;
    61: _omem00_bank = 55;
    62: _omem00_bank = 56;
    63: _omem00_bank = 57;
    64: _omem00_bank = 58;
    65: _omem00_bank = 59;
    default: _omem00_bank = 0;
    endcase
  end // always @ ( * )
  assign omem00_bank = _omem00_bank;
  reg _omem00_wr;
  always @ ( * ) begin
    case ( state )
    6: _omem00_wr = 1;
    7: _omem00_wr = 1;
    8: _omem00_wr = 1;
    9: _omem00_wr = 1;
    10: _omem00_wr = 1;
    11: _omem00_wr = 1;
    12: _omem00_wr = 1;
    13: _omem00_wr = 1;
    14: _omem00_wr = 1;
    15: _omem00_wr = 1;
    16: _omem00_wr = 1;
    17: _omem00_wr = 1;
    18: _omem00_wr = 1;
    19: _omem00_wr = 1;
    20: _omem00_wr = 1;
    21: _omem00_wr = 1;
    22: _omem00_wr = 1;
    23: _omem00_wr = 1;
    24: _omem00_wr = 1;
    25: _omem00_wr = 1;
    26: _omem00_wr = 1;
    27: _omem00_wr = 1;
    28: _omem00_wr = 1;
    29: _omem00_wr = 1;
    30: _omem00_wr = 1;
    31: _omem00_wr = 1;
    32: _omem00_wr = 1;
    33: _omem00_wr = 1;
    34: _omem00_wr = 1;
    35: _omem00_wr = 1;
    36: _omem00_wr = 1;
    37: _omem00_wr = 1;
    38: _omem00_wr = 1;
    39: _omem00_wr = 1;
    40: _omem00_wr = 1;
    41: _omem00_wr = 1;
    42: _omem00_wr = 1;
    43: _omem00_wr = 1;
    44: _omem00_wr = 1;
    45: _omem00_wr = 1;
    46: _omem00_wr = 1;
    47: _omem00_wr = 1;
    48: _omem00_wr = 1;
    49: _omem00_wr = 1;
    50: _omem00_wr = 1;
    51: _omem00_wr = 1;
    52: _omem00_wr = 1;
    53: _omem00_wr = 1;
    54: _omem00_wr = 1;
    55: _omem00_wr = 1;
    56: _omem00_wr = 1;
    57: _omem00_wr = 1;
    58: _omem00_wr = 1;
    59: _omem00_wr = 1;
    60: _omem00_wr = 1;
    61: _omem00_wr = 1;
    62: _omem00_wr = 1;
    63: _omem00_wr = 1;
    64: _omem00_wr = 1;
    65: _omem00_wr = 1;
    default: _omem00_wr = 0;
    endcase
  end // always @ ( * )
  assign omem00_wr = _omem00_wr;

  // 1番目の出力用メモリブロックの制御
  reg [5:0] _omem01_bank;
  always @ ( * ) begin
    case ( state )
    23: _omem01_bank = 0;
    24: _omem01_bank = 1;
    25: _omem01_bank = 2;
    26: _omem01_bank = 3;
    27: _omem01_bank = 4;
    28: _omem01_bank = 5;
    29: _omem01_bank = 6;
    30: _omem01_bank = 7;
    31: _omem01_bank = 8;
    32: _omem01_bank = 9;
    33: _omem01_bank = 10;
    34: _omem01_bank = 11;
    35: _omem01_bank = 12;
    36: _omem01_bank = 13;
    37: _omem01_bank = 14;
    38: _omem01_bank = 15;
    39: _omem01_bank = 16;
    40: _omem01_bank = 17;
    41: _omem01_bank = 18;
    42: _omem01_bank = 19;
    43: _omem01_bank = 20;
    44: _omem01_bank = 21;
    45: _omem01_bank = 22;
    46: _omem01_bank = 23;
    47: _omem01_bank = 24;
    48: _omem01_bank = 25;
    49: _omem01_bank = 26;
    50: _omem01_bank = 27;
    51: _omem01_bank = 28;
    52: _omem01_bank = 29;
    53: _omem01_bank = 30;
    54: _omem01_bank = 31;
    55: _omem01_bank = 32;
    56: _omem01_bank = 33;
    57: _omem01_bank = 34;
    58: _omem01_bank = 35;
    59: _omem01_bank = 36;
    60: _omem01_bank = 37;
    61: _omem01_bank = 38;
    62: _omem01_bank = 39;
    63: _omem01_bank = 40;
    64: _omem01_bank = 41;
    65: _omem01_bank = 42;
    66: _omem01_bank = 43;
    67: _omem01_bank = 44;
    68: _omem01_bank = 45;
    69: _omem01_bank = 46;
    70: _omem01_bank = 47;
    71: _omem01_bank = 48;
    72: _omem01_bank = 49;
    73: _omem01_bank = 50;
    74: _omem01_bank = 51;
    75: _omem01_bank = 52;
    76: _omem01_bank = 53;
    77: _omem01_bank = 54;
    78: _omem01_bank = 55;
    79: _omem01_bank = 56;
    80: _omem01_bank = 57;
    81: _omem01_bank = 58;
    82: _omem01_bank = 59;
    default: _omem01_bank = 0;
    endcase
  end // always @ ( * )
  assign omem01_bank = _omem01_bank;
  reg _omem01_wr;
  always @ ( * ) begin
    case ( state )
    23: _omem01_wr = 1;
    24: _omem01_wr = 1;
    25: _omem01_wr = 1;
    26: _omem01_wr = 1;
    27: _omem01_wr = 1;
    28: _omem01_wr = 1;
    29: _omem01_wr = 1;
    30: _omem01_wr = 1;
    31: _omem01_wr = 1;
    32: _omem01_wr = 1;
    33: _omem01_wr = 1;
    34: _omem01_wr = 1;
    35: _omem01_wr = 1;
    36: _omem01_wr = 1;
    37: _omem01_wr = 1;
    38: _omem01_wr = 1;
    39: _omem01_wr = 1;
    40: _omem01_wr = 1;
    41: _omem01_wr = 1;
    42: _omem01_wr = 1;
    43: _omem01_wr = 1;
    44: _omem01_wr = 1;
    45: _omem01_wr = 1;
    46: _omem01_wr = 1;
    47: _omem01_wr = 1;
    48: _omem01_wr = 1;
    49: _omem01_wr = 1;
    50: _omem01_wr = 1;
    51: _omem01_wr = 1;
    52: _omem01_wr = 1;
    53: _omem01_wr = 1;
    54: _omem01_wr = 1;
    55: _omem01_wr = 1;
    56: _omem01_wr = 1;
    57: _omem01_wr = 1;
    58: _omem01_wr = 1;
    59: _omem01_wr = 1;
    60: _omem01_wr = 1;
    61: _omem01_wr = 1;
    62: _omem01_wr = 1;
    63: _omem01_wr = 1;
    64: _omem01_wr = 1;
    65: _omem01_wr = 1;
    66: _omem01_wr = 1;
    67: _omem01_wr = 1;
    68: _omem01_wr = 1;
    69: _omem01_wr = 1;
    70: _omem01_wr = 1;
    71: _omem01_wr = 1;
    72: _omem01_wr = 1;
    73: _omem01_wr = 1;
    74: _omem01_wr = 1;
    75: _omem01_wr = 1;
    76: _omem01_wr = 1;
    77: _omem01_wr = 1;
    78: _omem01_wr = 1;
    79: _omem01_wr = 1;
    80: _omem01_wr = 1;
    81: _omem01_wr = 1;
    82: _omem01_wr = 1;
    default: _omem01_wr = 0;
    endcase
  end // always @ ( * )
  assign omem01_wr = _omem01_wr;

  // 2番目の出力用メモリブロックの制御
  reg [5:0] _omem02_bank;
  always @ ( * ) begin
    case ( state )
    42: _omem02_bank = 0;
    43: _omem02_bank = 1;
    44: _omem02_bank = 2;
    45: _omem02_bank = 3;
    46: _omem02_bank = 4;
    47: _omem02_bank = 5;
    48: _omem02_bank = 6;
    49: _omem02_bank = 7;
    50: _omem02_bank = 8;
    51: _omem02_bank = 9;
    52: _omem02_bank = 10;
    53: _omem02_bank = 11;
    54: _omem02_bank = 12;
    55: _omem02_bank = 13;
    56: _omem02_bank = 14;
    57: _omem02_bank = 15;
    58: _omem02_bank = 16;
    59: _omem02_bank = 17;
    60: _omem02_bank = 18;
    61: _omem02_bank = 19;
    62: _omem02_bank = 20;
    63: _omem02_bank = 21;
    64: _omem02_bank = 22;
    65: _omem02_bank = 23;
    66: _omem02_bank = 24;
    67: _omem02_bank = 25;
    68: _omem02_bank = 26;
    69: _omem02_bank = 27;
    70: _omem02_bank = 28;
    71: _omem02_bank = 29;
    72: _omem02_bank = 30;
    73: _omem02_bank = 31;
    74: _omem02_bank = 32;
    75: _omem02_bank = 33;
    76: _omem02_bank = 34;
    77: _omem02_bank = 35;
    78: _omem02_bank = 36;
    79: _omem02_bank = 37;
    80: _omem02_bank = 38;
    81: _omem02_bank = 39;
    82: _omem02_bank = 40;
    83: _omem02_bank = 41;
    84: _omem02_bank = 42;
    85: _omem02_bank = 43;
    86: _omem02_bank = 44;
    87: _omem02_bank = 45;
    88: _omem02_bank = 46;
    89: _omem02_bank = 47;
    90: _omem02_bank = 48;
    91: _omem02_bank = 49;
    92: _omem02_bank = 50;
    93: _omem02_bank = 51;
    94: _omem02_bank = 52;
    95: _omem02_bank = 53;
    96: _omem02_bank = 54;
    97: _omem02_bank = 55;
    98: _omem02_bank = 56;
    99: _omem02_bank = 57;
    100: _omem02_bank = 58;
    101: _omem02_bank = 59;
    default: _omem02_bank = 0;
    endcase
  end // always @ ( * )
  assign omem02_bank = _omem02_bank;
  reg _omem02_wr;
  always @ ( * ) begin
    case ( state )
    42: _omem02_wr = 1;
    43: _omem02_wr = 1;
    44: _omem02_wr = 1;
    45: _omem02_wr = 1;
    46: _omem02_wr = 1;
    47: _omem02_wr = 1;
    48: _omem02_wr = 1;
    49: _omem02_wr = 1;
    50: _omem02_wr = 1;
    51: _omem02_wr = 1;
    52: _omem02_wr = 1;
    53: _omem02_wr = 1;
    54: _omem02_wr = 1;
    55: _omem02_wr = 1;
    56: _omem02_wr = 1;
    57: _omem02_wr = 1;
    58: _omem02_wr = 1;
    59: _omem02_wr = 1;
    60: _omem02_wr = 1;
    61: _omem02_wr = 1;
    62: _omem02_wr = 1;
    63: _omem02_wr = 1;
    64: _omem02_wr = 1;
    65: _omem02_wr = 1;
    66: _omem02_wr = 1;
    67: _omem02_wr = 1;
    68: _omem02_wr = 1;
    69: _omem02_wr = 1;
    70: _omem02_wr = 1;
    71: _omem02_wr = 1;
    72: _omem02_wr = 1;
    73: _omem02_wr = 1;
    74: _omem02_wr = 1;
    75: _omem02_wr = 1;
    76: _omem02_wr = 1;
    77: _omem02_wr = 1;
    78: _omem02_wr = 1;
    79: _omem02_wr = 1;
    80: _omem02_wr = 1;
    81: _omem02_wr = 1;
    82: _omem02_wr = 1;
    83: _omem02_wr = 1;
    84: _omem02_wr = 1;
    85: _omem02_wr = 1;
    86: _omem02_wr = 1;
    87: _omem02_wr = 1;
    88: _omem02_wr = 1;
    89: _omem02_wr = 1;
    90: _omem02_wr = 1;
    91: _omem02_wr = 1;
    92: _omem02_wr = 1;
    93: _omem02_wr = 1;
    94: _omem02_wr = 1;
    95: _omem02_wr = 1;
    96: _omem02_wr = 1;
    97: _omem02_wr = 1;
    98: _omem02_wr = 1;
    99: _omem02_wr = 1;
    100: _omem02_wr = 1;
    101: _omem02_wr = 1;
    default: _omem02_wr = 0;
    endcase
  end // always @ ( * )
  assign omem02_wr = _omem02_wr;

  // 3番目の出力用メモリブロックの制御
  reg [5:0] _omem03_bank;
  always @ ( * ) begin
    case ( state )
    61: _omem03_bank = 0;
    62: _omem03_bank = 1;
    63: _omem03_bank = 2;
    64: _omem03_bank = 3;
    65: _omem03_bank = 4;
    66: _omem03_bank = 5;
    67: _omem03_bank = 6;
    68: _omem03_bank = 7;
    69: _omem03_bank = 8;
    70: _omem03_bank = 9;
    71: _omem03_bank = 10;
    72: _omem03_bank = 11;
    73: _omem03_bank = 12;
    74: _omem03_bank = 13;
    75: _omem03_bank = 14;
    76: _omem03_bank = 15;
    77: _omem03_bank = 16;
    78: _omem03_bank = 17;
    79: _omem03_bank = 18;
    80: _omem03_bank = 19;
    81: _omem03_bank = 20;
    82: _omem03_bank = 21;
    83: _omem03_bank = 22;
    84: _omem03_bank = 23;
    85: _omem03_bank = 24;
    86: _omem03_bank = 25;
    87: _omem03_bank = 26;
    88: _omem03_bank = 27;
    89: _omem03_bank = 28;
    90: _omem03_bank = 29;
    91: _omem03_bank = 30;
    92: _omem03_bank = 31;
    93: _omem03_bank = 32;
    94: _omem03_bank = 33;
    95: _omem03_bank = 34;
    96: _omem03_bank = 35;
    97: _omem03_bank = 36;
    98: _omem03_bank = 37;
    99: _omem03_bank = 38;
    100: _omem03_bank = 39;
    101: _omem03_bank = 40;
    102: _omem03_bank = 41;
    103: _omem03_bank = 42;
    104: _omem03_bank = 43;
    105: _omem03_bank = 44;
    106: _omem03_bank = 45;
    107: _omem03_bank = 46;
    108: _omem03_bank = 47;
    109: _omem03_bank = 48;
    110: _omem03_bank = 49;
    111: _omem03_bank = 50;
    112: _omem03_bank = 51;
    113: _omem03_bank = 52;
    114: _omem03_bank = 53;
    115: _omem03_bank = 54;
    116: _omem03_bank = 55;
    117: _omem03_bank = 56;
    118: _omem03_bank = 57;
    119: _omem03_bank = 58;
    120: _omem03_bank = 59;
    default: _omem03_bank = 0;
    endcase
  end // always @ ( * )
  assign omem03_bank = _omem03_bank;
  reg _omem03_wr;
  always @ ( * ) begin
    case ( state )
    61: _omem03_wr = 1;
    62: _omem03_wr = 1;
    63: _omem03_wr = 1;
    64: _omem03_wr = 1;
    65: _omem03_wr = 1;
    66: _omem03_wr = 1;
    67: _omem03_wr = 1;
    68: _omem03_wr = 1;
    69: _omem03_wr = 1;
    70: _omem03_wr = 1;
    71: _omem03_wr = 1;
    72: _omem03_wr = 1;
    73: _omem03_wr = 1;
    74: _omem03_wr = 1;
    75: _omem03_wr = 1;
    76: _omem03_wr = 1;
    77: _omem03_wr = 1;
    78: _omem03_wr = 1;
    79: _omem03_wr = 1;
    80: _omem03_wr = 1;
    81: _omem03_wr = 1;
    82: _omem03_wr = 1;
    83: _omem03_wr = 1;
    84: _omem03_wr = 1;
    85: _omem03_wr = 1;
    86: _omem03_wr = 1;
    87: _omem03_wr = 1;
    88: _omem03_wr = 1;
    89: _omem03_wr = 1;
    90: _omem03_wr = 1;
    91: _omem03_wr = 1;
    92: _omem03_wr = 1;
    93: _omem03_wr = 1;
    94: _omem03_wr = 1;
    95: _omem03_wr = 1;
    96: _omem03_wr = 1;
    97: _omem03_wr = 1;
    98: _omem03_wr = 1;
    99: _omem03_wr = 1;
    100: _omem03_wr = 1;
    101: _omem03_wr = 1;
    102: _omem03_wr = 1;
    103: _omem03_wr = 1;
    104: _omem03_wr = 1;
    105: _omem03_wr = 1;
    106: _omem03_wr = 1;
    107: _omem03_wr = 1;
    108: _omem03_wr = 1;
    109: _omem03_wr = 1;
    110: _omem03_wr = 1;
    111: _omem03_wr = 1;
    112: _omem03_wr = 1;
    113: _omem03_wr = 1;
    114: _omem03_wr = 1;
    115: _omem03_wr = 1;
    116: _omem03_wr = 1;
    117: _omem03_wr = 1;
    118: _omem03_wr = 1;
    119: _omem03_wr = 1;
    120: _omem03_wr = 1;
    default: _omem03_wr = 0;
    endcase
  end // always @ ( * )
  assign omem03_wr = _omem03_wr;

  // 4番目の出力用メモリブロックの制御
  reg [5:0] _omem04_bank;
  always @ ( * ) begin
    case ( state )
    80: _omem04_bank = 0;
    81: _omem04_bank = 1;
    82: _omem04_bank = 2;
    83: _omem04_bank = 3;
    84: _omem04_bank = 4;
    85: _omem04_bank = 5;
    86: _omem04_bank = 6;
    87: _omem04_bank = 7;
    88: _omem04_bank = 8;
    89: _omem04_bank = 9;
    90: _omem04_bank = 10;
    91: _omem04_bank = 11;
    92: _omem04_bank = 12;
    93: _omem04_bank = 13;
    94: _omem04_bank = 14;
    95: _omem04_bank = 15;
    96: _omem04_bank = 16;
    97: _omem04_bank = 17;
    98: _omem04_bank = 18;
    99: _omem04_bank = 19;
    100: _omem04_bank = 20;
    101: _omem04_bank = 21;
    102: _omem04_bank = 22;
    103: _omem04_bank = 23;
    104: _omem04_bank = 24;
    105: _omem04_bank = 25;
    106: _omem04_bank = 26;
    107: _omem04_bank = 27;
    108: _omem04_bank = 28;
    109: _omem04_bank = 29;
    110: _omem04_bank = 30;
    111: _omem04_bank = 31;
    112: _omem04_bank = 32;
    113: _omem04_bank = 33;
    114: _omem04_bank = 34;
    115: _omem04_bank = 35;
    116: _omem04_bank = 36;
    117: _omem04_bank = 37;
    118: _omem04_bank = 38;
    119: _omem04_bank = 39;
    120: _omem04_bank = 40;
    121: _omem04_bank = 41;
    122: _omem04_bank = 42;
    123: _omem04_bank = 43;
    124: _omem04_bank = 44;
    125: _omem04_bank = 45;
    126: _omem04_bank = 46;
    127: _omem04_bank = 47;
    128: _omem04_bank = 48;
    129: _omem04_bank = 49;
    130: _omem04_bank = 50;
    131: _omem04_bank = 51;
    132: _omem04_bank = 52;
    133: _omem04_bank = 53;
    134: _omem04_bank = 54;
    135: _omem04_bank = 55;
    136: _omem04_bank = 56;
    137: _omem04_bank = 57;
    default: _omem04_bank = 0;
    endcase
  end // always @ ( * )
  assign omem04_bank = _omem04_bank;
  reg _omem04_wr;
  always @ ( * ) begin
    case ( state )
    80: _omem04_wr = 1;
    81: _omem04_wr = 1;
    82: _omem04_wr = 1;
    83: _omem04_wr = 1;
    84: _omem04_wr = 1;
    85: _omem04_wr = 1;
    86: _omem04_wr = 1;
    87: _omem04_wr = 1;
    88: _omem04_wr = 1;
    89: _omem04_wr = 1;
    90: _omem04_wr = 1;
    91: _omem04_wr = 1;
    92: _omem04_wr = 1;
    93: _omem04_wr = 1;
    94: _omem04_wr = 1;
    95: _omem04_wr = 1;
    96: _omem04_wr = 1;
    97: _omem04_wr = 1;
    98: _omem04_wr = 1;
    99: _omem04_wr = 1;
    100: _omem04_wr = 1;
    101: _omem04_wr = 1;
    102: _omem04_wr = 1;
    103: _omem04_wr = 1;
    104: _omem04_wr = 1;
    105: _omem04_wr = 1;
    106: _omem04_wr = 1;
    107: _omem04_wr = 1;
    108: _omem04_wr = 1;
    109: _omem04_wr = 1;
    110: _omem04_wr = 1;
    111: _omem04_wr = 1;
    112: _omem04_wr = 1;
    113: _omem04_wr = 1;
    114: _omem04_wr = 1;
    115: _omem04_wr = 1;
    116: _omem04_wr = 1;
    117: _omem04_wr = 1;
    118: _omem04_wr = 1;
    119: _omem04_wr = 1;
    120: _omem04_wr = 1;
    121: _omem04_wr = 1;
    122: _omem04_wr = 1;
    123: _omem04_wr = 1;
    124: _omem04_wr = 1;
    125: _omem04_wr = 1;
    126: _omem04_wr = 1;
    127: _omem04_wr = 1;
    128: _omem04_wr = 1;
    129: _omem04_wr = 1;
    130: _omem04_wr = 1;
    131: _omem04_wr = 1;
    132: _omem04_wr = 1;
    133: _omem04_wr = 1;
    134: _omem04_wr = 1;
    135: _omem04_wr = 1;
    136: _omem04_wr = 1;
    137: _omem04_wr = 1;
    default: _omem04_wr = 0;
    endcase
  end // always @ ( * )
  assign omem04_wr = _omem04_wr;
  reg [8:0] _omem00_out;
  always @ ( * ) begin
    case ( state )
    6: _omem00_out = reg_0022;
    7: _omem00_out = reg_0023;
    8: _omem00_out = reg_0024;
    9: _omem00_out = reg_0022;
    10: _omem00_out = reg_0221;
    11: _omem00_out = reg_0222;
    12: _omem00_out = reg_0223;
    13: _omem00_out = reg_0745;
    14: _omem00_out = reg_0023;
    15: _omem00_out = reg_0746;
    16: _omem00_out = reg_0026;
    17: _omem00_out = reg_0027;
    18: _omem00_out = reg_0024;
    19: _omem00_out = reg_0022;
    20: _omem00_out = reg_0524;
    21: _omem00_out = reg_0754;
    22: _omem00_out = reg_0823;
    23: _omem00_out = reg_0738;
    24: _omem00_out = reg_0221;
    25: _omem00_out = reg_0739;
    26: _omem00_out = reg_0045;
    27: _omem00_out = reg_0250;
    28: _omem00_out = reg_0222;
    29: _omem00_out = reg_0044;
    30: _omem00_out = reg_0046;
    31: _omem00_out = reg_0251;
    32: _omem00_out = reg_0223;
    33: _omem00_out = reg_0745;
    34: _omem00_out = reg_0047;
    35: _omem00_out = reg_0252;
    36: _omem00_out = reg_0042;
    37: _omem00_out = reg_0023;
    38: _omem00_out = reg_0048;
    39: _omem00_out = reg_0049;
    40: _omem00_out = reg_0228;
    41: _omem00_out = reg_0230;
    42: _omem00_out = reg_0746;
    43: _omem00_out = reg_0026;
    44: _omem00_out = reg_0261;
    45: _omem00_out = reg_0263;
    46: _omem00_out = reg_0287;
    47: _omem00_out = reg_0027;
    48: _omem00_out = reg_0300;
    49: _omem00_out = reg_0310;
    50: _omem00_out = reg_0509;
    51: _omem00_out = reg_0024;
    52: _omem00_out = reg_0528;
    53: _omem00_out = reg_0022;
    54: _omem00_out = reg_0312;
    55: _omem00_out = reg_0313;
    56: _omem00_out = reg_0522;
    57: _omem00_out = reg_0524;
    58: _omem00_out = reg_0543;
    59: _omem00_out = reg_0546;
    60: _omem00_out = reg_0521;
    61: _omem00_out = reg_0525;
    62: _omem00_out = reg_0754;
    63: _omem00_out = reg_0325;
    64: _omem00_out = reg_0326;
    65: _omem00_out = reg_0327;
    default: _omem00_out = 0;
    endcase
  end // always @ ( * )
  assign omem00_out = _omem00_out[8:0];
  reg [8:0] _omem01_out;
  always @ ( * ) begin
    case ( state )
    23: _omem01_out = reg_0823;
    24: _omem01_out = reg_0738;
    25: _omem01_out = reg_0331;
    26: _omem01_out = reg_0332;
    27: _omem01_out = reg_0738;
    28: _omem01_out = reg_0221;
    29: _omem01_out = reg_0034;
    30: _omem01_out = reg_0823;
    31: _omem01_out = reg_0330;
    32: _omem01_out = reg_0335;
    33: _omem01_out = reg_0739;
    34: _omem01_out = reg_0045;
    35: _omem01_out = reg_0379;
    36: _omem01_out = reg_0332;
    37: _omem01_out = reg_0382;
    38: _omem01_out = reg_0738;
    39: _omem01_out = reg_0250;
    40: _omem01_out = reg_0264;
    41: _omem01_out = reg_0390;
    42: _omem01_out = reg_0221;
    43: _omem01_out = reg_0222;
    44: _omem01_out = reg_0044;
    45: _omem01_out = reg_0036;
    46: _omem01_out = reg_0034;
    47: _omem01_out = reg_0399;
    48: _omem01_out = reg_0823;
    49: _omem01_out = reg_0046;
    50: _omem01_out = reg_0826;
    51: _omem01_out = reg_0330;
    52: _omem01_out = reg_0033;
    53: _omem01_out = reg_0251;
    54: _omem01_out = reg_0030;
    55: _omem01_out = reg_0335;
    56: _omem01_out = reg_0035;
    57: _omem01_out = reg_0223;
    58: _omem01_out = reg_0745;
    59: _omem01_out = reg_0534;
    60: _omem01_out = reg_0739;
    61: _omem01_out = reg_0045;
    62: _omem01_out = reg_0047;
    63: _omem01_out = reg_0381;
    64: _omem01_out = reg_0284;
    65: _omem01_out = reg_0379;
    66: _omem01_out = reg_0252;
    67: _omem01_out = reg_0042;
    68: _omem01_out = reg_0072;
    69: _omem01_out = reg_0332;
    70: _omem01_out = reg_0380;
    71: _omem01_out = reg_0023;
    72: _omem01_out = reg_0415;
    73: _omem01_out = reg_0382;
    74: _omem01_out = reg_0738;
    75: _omem01_out = reg_0041;
    76: _omem01_out = reg_0048;
    77: _omem01_out = reg_0273;
    78: _omem01_out = reg_0250;
    79: _omem01_out = reg_0274;
    80: _omem01_out = reg_0228;
    81: _omem01_out = reg_0428;
    82: _omem01_out = reg_0264;
    default: _omem01_out = 0;
    endcase
  end // always @ ( * )
  assign omem01_out = _omem01_out[8:0];
  reg [8:0] _omem02_out;
  always @ ( * ) begin
    case ( state )
    42: _omem02_out = reg_0390;
    43: _omem02_out = reg_0230;
    44: _omem02_out = reg_0049;
    45: _omem02_out = reg_0390;
    46: _omem02_out = reg_0221;
    47: _omem02_out = reg_0746;
    48: _omem02_out = reg_0026;
    49: _omem02_out = reg_0230;
    50: _omem02_out = reg_0222;
    51: _omem02_out = reg_0281;
    52: _omem02_out = reg_0044;
    53: _omem02_out = reg_0261;
    54: _omem02_out = reg_0049;
    55: _omem02_out = reg_0390;
    56: _omem02_out = reg_0036;
    57: _omem02_out = reg_0263;
    58: _omem02_out = reg_0287;
    59: _omem02_out = reg_0221;
    60: _omem02_out = reg_0034;
    61: _omem02_out = reg_0271;
    62: _omem02_out = reg_0648;
    63: _omem02_out = reg_0027;
    64: _omem02_out = reg_0746;
    65: _omem02_out = reg_0026;
    66: _omem02_out = reg_0282;
    67: _omem02_out = reg_0300;
    68: _omem02_out = reg_0310;
    69: _omem02_out = reg_0046;
    70: _omem02_out = reg_0254;
    71: _omem02_out = reg_0823;
    72: _omem02_out = reg_0272;
    73: _omem02_out = reg_0222;
    74: _omem02_out = reg_0330;
    75: _omem02_out = reg_0230;
    76: _omem02_out = reg_0024;
    77: _omem02_out = reg_0044;
    78: _omem02_out = reg_0033;
    79: _omem02_out = reg_0826;
    80: _omem02_out = reg_0022;
    81: _omem02_out = reg_0261;
    82: _omem02_out = reg_0251;
    83: _omem02_out = reg_0030;
    84: _omem02_out = reg_0312;
    85: _omem02_out = reg_0049;
    86: _omem02_out = reg_0390;
    87: _omem02_out = reg_0335;
    88: _omem02_out = reg_0313;
    89: _omem02_out = reg_0522;
    90: _omem02_out = reg_0036;
    91: _omem02_out = reg_0662;
    92: _omem02_out = reg_0286;
    93: _omem02_out = reg_0524;
    94: _omem02_out = reg_0263;
    95: _omem02_out = reg_0287;
    96: _omem02_out = reg_0482;
    97: _omem02_out = reg_0543;
    98: _omem02_out = reg_0745;
    99: _omem02_out = reg_0221;
    100: _omem02_out = reg_0798;
    101: _omem02_out = reg_0546;
    default: _omem02_out = 0;
    endcase
  end // always @ ( * )
  assign omem02_out = _omem02_out[8:0];
  reg [8:0] _omem03_out;
  always @ ( * ) begin
    case ( state )
    61: _omem03_out = reg_0521;
    62: _omem03_out = reg_0269;
    63: _omem03_out = reg_0521;
    64: _omem03_out = reg_0525;
    65: _omem03_out = reg_0034;
    66: _omem03_out = reg_0271;
    67: _omem03_out = reg_0648;
    68: _omem03_out = reg_0047;
    69: _omem03_out = reg_0754;
    70: _omem03_out = reg_0325;
    71: _omem03_out = reg_0027;
    72: _omem03_out = reg_0381;
    73: _omem03_out = reg_0284;
    74: _omem03_out = reg_0269;
    75: _omem03_out = reg_0746;
    76: _omem03_out = reg_0026;
    77: _omem03_out = reg_0379;
    78: _omem03_out = reg_0327;
    79: _omem03_out = reg_0521;
    80: _omem03_out = reg_0525;
    81: _omem03_out = reg_0561;
    82: _omem03_out = reg_0042;
    83: _omem03_out = reg_0129;
    84: _omem03_out = reg_0300;
    85: _omem03_out = reg_0310;
    86: _omem03_out = reg_0047;
    87: _omem03_out = reg_0373;
    88: _omem03_out = reg_0271;
    89: _omem03_out = reg_0701;
    90: _omem03_out = reg_0046;
    91: _omem03_out = reg_0332;
    92: _omem03_out = reg_0380;
    93: _omem03_out = reg_0072;
    94: _omem03_out = reg_0034;
    95: _omem03_out = reg_0823;
    96: _omem03_out = reg_0023;
    97: _omem03_out = reg_0706;
    98: _omem03_out = reg_0707;
    99: _omem03_out = reg_0831;
    100: _omem03_out = reg_0272;
    101: _omem03_out = reg_0381;
    102: _omem03_out = reg_0284;
    103: _omem03_out = reg_0282;
    104: _omem03_out = reg_0222;
    105: _omem03_out = reg_0330;
    106: _omem03_out = reg_0269;
    107: _omem03_out = reg_0082;
    108: _omem03_out = reg_0738;
    109: _omem03_out = reg_0041;
    110: _omem03_out = reg_0415;
    111: _omem03_out = reg_0040;
    112: _omem03_out = reg_0026;
    113: _omem03_out = reg_0230;
    114: _omem03_out = reg_0024;
    115: _omem03_out = reg_0273;
    116: _omem03_out = reg_0379;
    117: _omem03_out = reg_0746;
    118: _omem03_out = reg_0172;
    119: _omem03_out = reg_0033;
    120: _omem03_out = reg_0048;
    default: _omem03_out = 0;
    endcase
  end // always @ ( * )
  assign omem03_out = _omem03_out[8:0];
  reg [8:0] _omem04_out;
  always @ ( * ) begin
    case ( state )
    80: _omem04_out = reg_0521;
    81: _omem04_out = reg_0250;
    82: _omem04_out = reg_0274;
    83: _omem04_out = reg_0022;
    84: _omem04_out = reg_0525;
    85: _omem04_out = reg_0254;
    86: _omem04_out = reg_0045;
    87: _omem04_out = reg_0250;
    88: _omem04_out = reg_0561;
    89: _omem04_out = reg_0521;
    90: _omem04_out = reg_0428;
    91: _omem04_out = reg_0035;
    92: _omem04_out = reg_0022;
    93: _omem04_out = reg_0129;
    94: _omem04_out = reg_0739;
    95: _omem04_out = reg_0044;
    96: _omem04_out = reg_0312;
    97: _omem04_out = reg_0300;
    98: _omem04_out = reg_0310;
    99: _omem04_out = reg_0525;
    100: _omem04_out = reg_0049;
    101: _omem04_out = reg_0045;
    102: _omem04_out = reg_0047;
    103: _omem04_out = reg_0826;
    104: _omem04_out = reg_0682;
    105: _omem04_out = reg_0250;
    106: _omem04_out = reg_0373;
    107: _omem04_out = reg_0390;
    108: _omem04_out = reg_0652;
    109: _omem04_out = reg_0313;
    110: _omem04_out = reg_0521;
    111: _omem04_out = reg_0187;
    112: _omem04_out = reg_0754;
    113: _omem04_out = reg_0223;
    114: _omem04_out = reg_0701;
    115: _omem04_out = reg_0036;
    116: _omem04_out = reg_0270;
    117: _omem04_out = reg_0103;
    118: _omem04_out = reg_0428;
    119: _omem04_out = reg_0035;
    120: _omem04_out = reg_0022;
    121: _omem04_out = reg_0027;
    122: _omem04_out = reg_0252;
    123: _omem04_out = reg_0399;
    124: _omem04_out = reg_0042;
    125: _omem04_out = reg_0046;
    126: _omem04_out = reg_0254;
    127: _omem04_out = reg_0030;
    128: _omem04_out = reg_0072;
    129: _omem04_out = reg_0034;
    130: _omem04_out = reg_0044;
    131: _omem04_out = reg_0129;
    132: _omem04_out = reg_0263;
    133: _omem04_out = reg_0228;
    134: _omem04_out = reg_0023;
    135: _omem04_out = reg_0251;
    136: _omem04_out = reg_0286;
    137: _omem04_out = reg_0261;
    default: _omem04_out = 0;
    endcase
  end // always @ ( * )
  assign omem04_out = _omem04_out[8:0];

  // OP1#0の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in00 = imem00_in[59:56];
    2: op1_00_in00 = imem07_in[123:120];
    5: op1_00_in00 = imem03_in[95:92];
    3: op1_00_in00 = imem07_in[91:88];
    6: op1_00_in00 = imem00_in[23:20];
    1: op1_00_in00 = imem07_in[115:112];
    7: op1_00_in00 = imem04_in[103:100];
    8: op1_00_in00 = imem06_in[107:104];
    9: op1_00_in00 = imem01_in[107:104];
    10: op1_00_in00 = imem01_in[83:80];
    24: op1_00_in00 = imem01_in[83:80];
    11: op1_00_in00 = imem05_in[99:96];
    12: op1_00_in00 = imem00_in[7:4];
    13: op1_00_in00 = imem05_in[103:100];
    14: op1_00_in00 = imem00_in[27:24];
    29: op1_00_in00 = imem00_in[27:24];
    59: op1_00_in00 = imem00_in[27:24];
    76: op1_00_in00 = imem00_in[27:24];
    15: op1_00_in00 = imem00_in[11:8];
    38: op1_00_in00 = imem00_in[11:8];
    16: op1_00_in00 = imem03_in[91:88];
    17: op1_00_in00 = imem04_in[115:112];
    18: op1_00_in00 = imem04_in[31:28];
    19: op1_00_in00 = imem05_in[35:32];
    20: op1_00_in00 = imem02_in[15:12];
    21: op1_00_in00 = imem06_in[95:92];
    57: op1_00_in00 = imem06_in[95:92];
    22: op1_00_in00 = imem00_in[107:104];
    23: op1_00_in00 = imem04_in[111:108];
    25: op1_00_in00 = imem02_in[119:116];
    26: op1_00_in00 = imem00_in[3:0];
    37: op1_00_in00 = imem00_in[3:0];
    27: op1_00_in00 = imem03_in[127:124];
    28: op1_00_in00 = imem06_in[11:8];
    30: op1_00_in00 = imem03_in[99:96];
    54: op1_00_in00 = imem03_in[99:96];
    31: op1_00_in00 = imem06_in[15:12];
    66: op1_00_in00 = imem06_in[15:12];
    32: op1_00_in00 = imem00_in[35:32];
    46: op1_00_in00 = imem00_in[35:32];
    33: op1_00_in00 = imem00_in[43:40];
    34: op1_00_in00 = imem06_in[111:108];
    35: op1_00_in00 = imem06_in[63:60];
    70: op1_00_in00 = imem06_in[63:60];
    36: op1_00_in00 = imem06_in[103:100];
    39: op1_00_in00 = imem01_in[119:116];
    40: op1_00_in00 = imem01_in[79:76];
    41: op1_00_in00 = imem04_in[59:56];
    42: op1_00_in00 = imem07_in[107:104];
    43: op1_00_in00 = imem00_in[19:16];
    44: op1_00_in00 = imem02_in[63:60];
    71: op1_00_in00 = imem02_in[63:60];
    45: op1_00_in00 = imem04_in[23:20];
    47: op1_00_in00 = imem01_in[71:68];
    48: op1_00_in00 = imem04_in[79:76];
    49: op1_00_in00 = imem05_in[95:92];
    50: op1_00_in00 = imem04_in[95:92];
    51: op1_00_in00 = imem02_in[39:36];
    52: op1_00_in00 = imem01_in[99:96];
    53: op1_00_in00 = imem03_in[55:52];
    55: op1_00_in00 = imem05_in[19:16];
    65: op1_00_in00 = imem05_in[19:16];
    56: op1_00_in00 = imem07_in[111:108];
    58: op1_00_in00 = imem04_in[47:44];
    82: op1_00_in00 = imem04_in[47:44];
    60: op1_00_in00 = imem06_in[35:32];
    88: op1_00_in00 = imem06_in[35:32];
    61: op1_00_in00 = imem00_in[91:88];
    62: op1_00_in00 = imem02_in[7:4];
    63: op1_00_in00 = imem04_in[127:124];
    64: op1_00_in00 = imem05_in[83:80];
    67: op1_00_in00 = imem05_in[47:44];
    68: op1_00_in00 = imem01_in[31:28];
    69: op1_00_in00 = imem03_in[103:100];
    72: op1_00_in00 = imem05_in[59:56];
    73: op1_00_in00 = imem05_in[111:108];
    79: op1_00_in00 = imem05_in[111:108];
    74: op1_00_in00 = imem07_in[43:40];
    75: op1_00_in00 = imem00_in[75:72];
    77: op1_00_in00 = imem03_in[11:8];
    89: op1_00_in00 = imem03_in[11:8];
    78: op1_00_in00 = imem05_in[71:68];
    80: op1_00_in00 = imem07_in[47:44];
    81: op1_00_in00 = imem07_in[35:32];
    83: op1_00_in00 = imem02_in[75:72];
    84: op1_00_in00 = imem02_in[55:52];
    85: op1_00_in00 = imem06_in[75:72];
    86: op1_00_in00 = imem05_in[115:112];
    87: op1_00_in00 = imem03_in[47:44];
    90: op1_00_in00 = imem05_in[123:120];
    91: op1_00_in00 = imem06_in[3:0];
    92: op1_00_in00 = imem01_in[95:92];
    93: op1_00_in00 = imem01_in[27:24];
    94: op1_00_in00 = imem01_in[67:64];
    95: op1_00_in00 = imem00_in[79:76];
    96: op1_00_in00 = imem00_in[15:12];
    default: op1_00_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv00 = 1;
    9: op1_00_inv00 = 1;
    10: op1_00_inv00 = 1;
    13: op1_00_inv00 = 1;
    14: op1_00_inv00 = 1;
    15: op1_00_inv00 = 1;
    16: op1_00_inv00 = 1;
    17: op1_00_inv00 = 1;
    18: op1_00_inv00 = 1;
    19: op1_00_inv00 = 1;
    20: op1_00_inv00 = 1;
    21: op1_00_inv00 = 1;
    24: op1_00_inv00 = 1;
    26: op1_00_inv00 = 1;
    27: op1_00_inv00 = 1;
    28: op1_00_inv00 = 1;
    32: op1_00_inv00 = 1;
    34: op1_00_inv00 = 1;
    39: op1_00_inv00 = 1;
    41: op1_00_inv00 = 1;
    42: op1_00_inv00 = 1;
    43: op1_00_inv00 = 1;
    46: op1_00_inv00 = 1;
    48: op1_00_inv00 = 1;
    49: op1_00_inv00 = 1;
    53: op1_00_inv00 = 1;
    55: op1_00_inv00 = 1;
    56: op1_00_inv00 = 1;
    58: op1_00_inv00 = 1;
    59: op1_00_inv00 = 1;
    60: op1_00_inv00 = 1;
    61: op1_00_inv00 = 1;
    62: op1_00_inv00 = 1;
    63: op1_00_inv00 = 1;
    64: op1_00_inv00 = 1;
    66: op1_00_inv00 = 1;
    68: op1_00_inv00 = 1;
    69: op1_00_inv00 = 1;
    72: op1_00_inv00 = 1;
    73: op1_00_inv00 = 1;
    74: op1_00_inv00 = 1;
    76: op1_00_inv00 = 1;
    77: op1_00_inv00 = 1;
    82: op1_00_inv00 = 1;
    86: op1_00_inv00 = 1;
    87: op1_00_inv00 = 1;
    89: op1_00_inv00 = 1;
    91: op1_00_inv00 = 1;
    93: op1_00_inv00 = 1;
    94: op1_00_inv00 = 1;
    default: op1_00_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in01 = imem00_in[111:108];
    22: op1_00_in01 = imem00_in[111:108];
    32: op1_00_in01 = imem00_in[111:108];
    75: op1_00_in01 = imem00_in[111:108];
    2: op1_00_in01 = reg_0181;
    5: op1_00_in01 = imem04_in[67:64];
    3: op1_00_in01 = reg_0441;
    6: op1_00_in01 = imem00_in[27:24];
    37: op1_00_in01 = imem00_in[27:24];
    7: op1_00_in01 = imem04_in[115:112];
    8: op1_00_in01 = imem07_in[27:24];
    9: op1_00_in01 = imem01_in[111:108];
    52: op1_00_in01 = imem01_in[111:108];
    10: op1_00_in01 = imem01_in[95:92];
    24: op1_00_in01 = imem01_in[95:92];
    94: op1_00_in01 = imem01_in[95:92];
    11: op1_00_in01 = imem05_in[119:116];
    12: op1_00_in01 = imem00_in[39:36];
    14: op1_00_in01 = imem00_in[39:36];
    29: op1_00_in01 = imem00_in[39:36];
    96: op1_00_in01 = imem00_in[39:36];
    13: op1_00_in01 = imem05_in[111:108];
    15: op1_00_in01 = imem00_in[107:104];
    61: op1_00_in01 = imem00_in[107:104];
    16: op1_00_in01 = imem03_in[103:100];
    17: op1_00_in01 = imem05_in[47:44];
    18: op1_00_in01 = imem04_in[51:48];
    58: op1_00_in01 = imem04_in[51:48];
    19: op1_00_in01 = imem05_in[87:84];
    78: op1_00_in01 = imem05_in[87:84];
    20: op1_00_in01 = imem02_in[19:16];
    21: op1_00_in01 = imem06_in[99:96];
    23: op1_00_in01 = reg_0301;
    25: op1_00_in01 = reg_0314;
    26: op1_00_in01 = imem00_in[31:28];
    27: op1_00_in01 = reg_0012;
    28: op1_00_in01 = imem06_in[19:16];
    30: op1_00_in01 = imem03_in[115:112];
    54: op1_00_in01 = imem03_in[115:112];
    31: op1_00_in01 = imem06_in[83:80];
    33: op1_00_in01 = imem00_in[75:72];
    34: op1_00_in01 = reg_0629;
    35: op1_00_in01 = imem06_in[107:104];
    36: op1_00_in01 = imem06_in[111:108];
    38: op1_00_in01 = imem00_in[23:20];
    39: op1_00_in01 = reg_0102;
    40: op1_00_in01 = imem01_in[87:84];
    41: op1_00_in01 = reg_0078;
    42: op1_00_in01 = imem07_in[119:116];
    43: op1_00_in01 = imem00_in[63:60];
    44: op1_00_in01 = imem02_in[79:76];
    45: op1_00_in01 = imem04_in[39:36];
    46: op1_00_in01 = imem00_in[43:40];
    47: op1_00_in01 = imem01_in[75:72];
    48: op1_00_in01 = imem04_in[83:80];
    49: op1_00_in01 = imem05_in[107:104];
    50: op1_00_in01 = reg_0315;
    51: op1_00_in01 = imem02_in[43:40];
    53: op1_00_in01 = imem03_in[59:56];
    89: op1_00_in01 = imem03_in[59:56];
    55: op1_00_in01 = imem05_in[31:28];
    56: op1_00_in01 = imem07_in[115:112];
    57: op1_00_in01 = imem06_in[103:100];
    60: op1_00_in01 = imem06_in[103:100];
    59: op1_00_in01 = imem00_in[51:48];
    76: op1_00_in01 = imem00_in[51:48];
    62: op1_00_in01 = imem02_in[47:44];
    63: op1_00_in01 = reg_0043;
    64: op1_00_in01 = imem05_in[99:96];
    65: op1_00_in01 = imem05_in[43:40];
    66: op1_00_in01 = imem06_in[51:48];
    67: op1_00_in01 = imem05_in[55:52];
    68: op1_00_in01 = imem01_in[43:40];
    69: op1_00_in01 = reg_0006;
    70: op1_00_in01 = imem06_in[95:92];
    71: op1_00_in01 = imem02_in[71:68];
    72: op1_00_in01 = imem05_in[91:88];
    73: op1_00_in01 = imem06_in[43:40];
    74: op1_00_in01 = imem07_in[55:52];
    77: op1_00_in01 = imem03_in[19:16];
    79: op1_00_in01 = reg_0135;
    80: op1_00_in01 = imem07_in[51:48];
    81: op1_00_in01 = imem07_in[59:56];
    82: op1_00_in01 = imem04_in[55:52];
    83: op1_00_in01 = imem02_in[99:96];
    84: op1_00_in01 = imem02_in[91:88];
    85: op1_00_in01 = imem06_in[79:76];
    86: op1_00_in01 = reg_0812;
    87: op1_00_in01 = imem03_in[123:120];
    88: op1_00_in01 = imem06_in[55:52];
    90: op1_00_in01 = reg_0550;
    91: op1_00_in01 = imem06_in[7:4];
    92: op1_00_in01 = imem01_in[115:112];
    93: op1_00_in01 = imem01_in[31:28];
    95: op1_00_in01 = reg_0683;
    default: op1_00_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    3: op1_00_inv01 = 1;
    6: op1_00_inv01 = 1;
    8: op1_00_inv01 = 1;
    9: op1_00_inv01 = 1;
    12: op1_00_inv01 = 1;
    14: op1_00_inv01 = 1;
    17: op1_00_inv01 = 1;
    23: op1_00_inv01 = 1;
    25: op1_00_inv01 = 1;
    26: op1_00_inv01 = 1;
    29: op1_00_inv01 = 1;
    30: op1_00_inv01 = 1;
    31: op1_00_inv01 = 1;
    33: op1_00_inv01 = 1;
    36: op1_00_inv01 = 1;
    37: op1_00_inv01 = 1;
    38: op1_00_inv01 = 1;
    39: op1_00_inv01 = 1;
    40: op1_00_inv01 = 1;
    43: op1_00_inv01 = 1;
    44: op1_00_inv01 = 1;
    45: op1_00_inv01 = 1;
    46: op1_00_inv01 = 1;
    48: op1_00_inv01 = 1;
    49: op1_00_inv01 = 1;
    51: op1_00_inv01 = 1;
    57: op1_00_inv01 = 1;
    58: op1_00_inv01 = 1;
    60: op1_00_inv01 = 1;
    64: op1_00_inv01 = 1;
    66: op1_00_inv01 = 1;
    70: op1_00_inv01 = 1;
    71: op1_00_inv01 = 1;
    72: op1_00_inv01 = 1;
    73: op1_00_inv01 = 1;
    74: op1_00_inv01 = 1;
    75: op1_00_inv01 = 1;
    76: op1_00_inv01 = 1;
    78: op1_00_inv01 = 1;
    79: op1_00_inv01 = 1;
    80: op1_00_inv01 = 1;
    81: op1_00_inv01 = 1;
    82: op1_00_inv01 = 1;
    84: op1_00_inv01 = 1;
    86: op1_00_inv01 = 1;
    87: op1_00_inv01 = 1;
    89: op1_00_inv01 = 1;
    91: op1_00_inv01 = 1;
    92: op1_00_inv01 = 1;
    93: op1_00_inv01 = 1;
    94: op1_00_inv01 = 1;
    95: op1_00_inv01 = 1;
    default: op1_00_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in02 = imem00_in[115:112];
    15: op1_00_in02 = imem00_in[115:112];
    2: op1_00_in02 = reg_0169;
    5: op1_00_in02 = imem04_in[103:100];
    18: op1_00_in02 = imem04_in[103:100];
    3: op1_00_in02 = reg_0428;
    6: op1_00_in02 = imem00_in[63:60];
    7: op1_00_in02 = reg_0545;
    8: op1_00_in02 = imem07_in[95:92];
    9: op1_00_in02 = imem01_in[115:112];
    24: op1_00_in02 = imem01_in[115:112];
    40: op1_00_in02 = imem01_in[115:112];
    10: op1_00_in02 = reg_0232;
    11: op1_00_in02 = reg_0132;
    12: op1_00_in02 = imem00_in[59:56];
    29: op1_00_in02 = imem00_in[59:56];
    13: op1_00_in02 = reg_0798;
    14: op1_00_in02 = imem00_in[47:44];
    96: op1_00_in02 = imem00_in[47:44];
    16: op1_00_in02 = imem03_in[119:116];
    54: op1_00_in02 = imem03_in[119:116];
    17: op1_00_in02 = imem05_in[59:56];
    19: op1_00_in02 = reg_0147;
    20: op1_00_in02 = imem02_in[75:72];
    71: op1_00_in02 = imem02_in[75:72];
    21: op1_00_in02 = imem06_in[103:100];
    22: op1_00_in02 = reg_0684;
    23: op1_00_in02 = reg_0266;
    25: op1_00_in02 = reg_0770;
    26: op1_00_in02 = imem00_in[55:52];
    46: op1_00_in02 = imem00_in[55:52];
    27: op1_00_in02 = reg_0803;
    28: op1_00_in02 = imem06_in[23:20];
    91: op1_00_in02 = imem06_in[23:20];
    30: op1_00_in02 = reg_0569;
    31: op1_00_in02 = imem07_in[3:0];
    32: op1_00_in02 = reg_0689;
    33: op1_00_in02 = imem00_in[79:76];
    34: op1_00_in02 = reg_0630;
    35: op1_00_in02 = reg_0025;
    36: op1_00_in02 = imem06_in[115:112];
    37: op1_00_in02 = imem00_in[31:28];
    38: op1_00_in02 = imem00_in[91:88];
    39: op1_00_in02 = reg_0114;
    41: op1_00_in02 = reg_0062;
    42: op1_00_in02 = reg_0179;
    43: op1_00_in02 = imem00_in[67:64];
    76: op1_00_in02 = imem00_in[67:64];
    44: op1_00_in02 = imem02_in[87:84];
    45: op1_00_in02 = imem04_in[67:64];
    47: op1_00_in02 = imem01_in[95:92];
    48: op1_00_in02 = imem04_in[87:84];
    49: op1_00_in02 = imem05_in[115:112];
    50: op1_00_in02 = reg_0553;
    51: op1_00_in02 = imem02_in[59:56];
    52: op1_00_in02 = imem02_in[35:32];
    53: op1_00_in02 = imem03_in[71:68];
    55: op1_00_in02 = imem05_in[71:68];
    56: op1_00_in02 = reg_0721;
    57: op1_00_in02 = imem06_in[127:124];
    58: op1_00_in02 = imem04_in[55:52];
    59: op1_00_in02 = imem00_in[95:92];
    60: op1_00_in02 = imem07_in[19:16];
    61: op1_00_in02 = imem00_in[119:116];
    62: op1_00_in02 = imem02_in[83:80];
    63: op1_00_in02 = reg_0555;
    64: op1_00_in02 = imem05_in[111:108];
    65: op1_00_in02 = imem05_in[83:80];
    66: op1_00_in02 = imem06_in[55:52];
    67: op1_00_in02 = imem05_in[87:84];
    68: op1_00_in02 = imem01_in[91:88];
    69: op1_00_in02 = reg_0811;
    70: op1_00_in02 = imem06_in[99:96];
    72: op1_00_in02 = imem05_in[107:104];
    73: op1_00_in02 = imem06_in[59:56];
    74: op1_00_in02 = reg_0295;
    75: op1_00_in02 = reg_0683;
    77: op1_00_in02 = imem03_in[23:20];
    78: op1_00_in02 = imem05_in[119:116];
    79: op1_00_in02 = reg_0227;
    80: op1_00_in02 = imem07_in[59:56];
    81: op1_00_in02 = imem07_in[63:60];
    82: op1_00_in02 = imem04_in[123:120];
    83: op1_00_in02 = imem02_in[111:108];
    84: op1_00_in02 = imem03_in[43:40];
    85: op1_00_in02 = reg_0573;
    86: op1_00_in02 = reg_0148;
    87: op1_00_in02 = reg_0549;
    88: op1_00_in02 = imem06_in[79:76];
    89: op1_00_in02 = imem03_in[63:60];
    90: op1_00_in02 = reg_0231;
    92: op1_00_in02 = reg_0105;
    93: op1_00_in02 = imem01_in[55:52];
    94: op1_00_in02 = imem01_in[111:108];
    95: op1_00_in02 = reg_0112;
    default: op1_00_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv02 = 1;
    5: op1_00_inv02 = 1;
    6: op1_00_inv02 = 1;
    8: op1_00_inv02 = 1;
    10: op1_00_inv02 = 1;
    11: op1_00_inv02 = 1;
    12: op1_00_inv02 = 1;
    16: op1_00_inv02 = 1;
    18: op1_00_inv02 = 1;
    19: op1_00_inv02 = 1;
    21: op1_00_inv02 = 1;
    23: op1_00_inv02 = 1;
    24: op1_00_inv02 = 1;
    26: op1_00_inv02 = 1;
    27: op1_00_inv02 = 1;
    28: op1_00_inv02 = 1;
    31: op1_00_inv02 = 1;
    32: op1_00_inv02 = 1;
    34: op1_00_inv02 = 1;
    35: op1_00_inv02 = 1;
    36: op1_00_inv02 = 1;
    38: op1_00_inv02 = 1;
    41: op1_00_inv02 = 1;
    44: op1_00_inv02 = 1;
    45: op1_00_inv02 = 1;
    50: op1_00_inv02 = 1;
    52: op1_00_inv02 = 1;
    53: op1_00_inv02 = 1;
    55: op1_00_inv02 = 1;
    56: op1_00_inv02 = 1;
    57: op1_00_inv02 = 1;
    58: op1_00_inv02 = 1;
    59: op1_00_inv02 = 1;
    62: op1_00_inv02 = 1;
    63: op1_00_inv02 = 1;
    66: op1_00_inv02 = 1;
    67: op1_00_inv02 = 1;
    68: op1_00_inv02 = 1;
    69: op1_00_inv02 = 1;
    70: op1_00_inv02 = 1;
    71: op1_00_inv02 = 1;
    73: op1_00_inv02 = 1;
    74: op1_00_inv02 = 1;
    77: op1_00_inv02 = 1;
    79: op1_00_inv02 = 1;
    82: op1_00_inv02 = 1;
    89: op1_00_inv02 = 1;
    91: op1_00_inv02 = 1;
    95: op1_00_inv02 = 1;
    96: op1_00_inv02 = 1;
    default: op1_00_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in03 = reg_0683;
    2: op1_00_in03 = reg_0160;
    5: op1_00_in03 = imem04_in[107:104];
    18: op1_00_in03 = imem04_in[107:104];
    3: op1_00_in03 = reg_0442;
    6: op1_00_in03 = imem00_in[95:92];
    38: op1_00_in03 = imem00_in[95:92];
    7: op1_00_in03 = reg_0557;
    8: op1_00_in03 = imem07_in[107:104];
    9: op1_00_in03 = imem01_in[119:116];
    10: op1_00_in03 = reg_0220;
    11: op1_00_in03 = reg_0146;
    12: op1_00_in03 = imem00_in[67:64];
    13: op1_00_in03 = reg_0788;
    14: op1_00_in03 = imem00_in[51:48];
    37: op1_00_in03 = imem00_in[51:48];
    15: op1_00_in03 = reg_0694;
    75: op1_00_in03 = reg_0694;
    16: op1_00_in03 = reg_0573;
    17: op1_00_in03 = imem05_in[99:96];
    19: op1_00_in03 = reg_0148;
    20: op1_00_in03 = imem02_in[87:84];
    21: op1_00_in03 = imem06_in[111:108];
    22: op1_00_in03 = reg_0670;
    23: op1_00_in03 = reg_0284;
    24: op1_00_in03 = reg_0217;
    25: op1_00_in03 = reg_0526;
    26: op1_00_in03 = imem00_in[91:88];
    27: op1_00_in03 = reg_0807;
    28: op1_00_in03 = imem06_in[55:52];
    29: op1_00_in03 = imem00_in[71:68];
    30: op1_00_in03 = reg_0572;
    31: op1_00_in03 = imem07_in[23:20];
    32: op1_00_in03 = reg_0679;
    33: op1_00_in03 = imem00_in[83:80];
    34: op1_00_in03 = reg_0633;
    35: op1_00_in03 = reg_0331;
    36: op1_00_in03 = imem07_in[3:0];
    70: op1_00_in03 = imem07_in[3:0];
    39: op1_00_in03 = reg_0107;
    40: op1_00_in03 = reg_0123;
    41: op1_00_in03 = reg_0255;
    42: op1_00_in03 = reg_0169;
    43: op1_00_in03 = imem00_in[119:116];
    44: op1_00_in03 = imem02_in[119:116];
    45: op1_00_in03 = imem05_in[3:0];
    46: op1_00_in03 = imem00_in[59:56];
    47: op1_00_in03 = imem01_in[99:96];
    48: op1_00_in03 = imem04_in[111:108];
    49: op1_00_in03 = reg_0145;
    50: op1_00_in03 = reg_0328;
    51: op1_00_in03 = imem02_in[95:92];
    62: op1_00_in03 = imem02_in[95:92];
    52: op1_00_in03 = imem02_in[43:40];
    53: op1_00_in03 = imem03_in[87:84];
    89: op1_00_in03 = imem03_in[87:84];
    54: op1_00_in03 = reg_0395;
    55: op1_00_in03 = imem05_in[91:88];
    56: op1_00_in03 = reg_0713;
    57: op1_00_in03 = reg_0614;
    58: op1_00_in03 = imem04_in[59:56];
    59: op1_00_in03 = imem00_in[123:120];
    60: op1_00_in03 = imem07_in[27:24];
    61: op1_00_in03 = imem00_in[127:124];
    63: op1_00_in03 = reg_0052;
    64: op1_00_in03 = reg_0736;
    65: op1_00_in03 = imem05_in[119:116];
    66: op1_00_in03 = imem06_in[67:64];
    67: op1_00_in03 = imem05_in[95:92];
    68: op1_00_in03 = reg_0232;
    69: op1_00_in03 = reg_0002;
    71: op1_00_in03 = reg_0414;
    72: op1_00_in03 = reg_0279;
    73: op1_00_in03 = imem06_in[63:60];
    74: op1_00_in03 = reg_0067;
    76: op1_00_in03 = imem00_in[75:72];
    77: op1_00_in03 = imem03_in[67:64];
    78: op1_00_in03 = imem05_in[123:120];
    79: op1_00_in03 = reg_0666;
    80: op1_00_in03 = imem07_in[79:76];
    81: op1_00_in03 = imem07_in[115:112];
    82: op1_00_in03 = reg_0079;
    83: op1_00_in03 = reg_0587;
    84: op1_00_in03 = reg_0528;
    85: op1_00_in03 = reg_0563;
    86: op1_00_in03 = reg_0154;
    87: op1_00_in03 = reg_0747;
    88: op1_00_in03 = imem06_in[83:80];
    90: op1_00_in03 = reg_0134;
    91: op1_00_in03 = reg_0817;
    92: op1_00_in03 = reg_0124;
    93: op1_00_in03 = imem01_in[63:60];
    94: op1_00_in03 = reg_0673;
    95: op1_00_in03 = reg_0685;
    96: op1_00_in03 = imem00_in[99:96];
    default: op1_00_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    2: op1_00_inv03 = 1;
    5: op1_00_inv03 = 1;
    3: op1_00_inv03 = 1;
    6: op1_00_inv03 = 1;
    7: op1_00_inv03 = 1;
    9: op1_00_inv03 = 1;
    10: op1_00_inv03 = 1;
    11: op1_00_inv03 = 1;
    14: op1_00_inv03 = 1;
    17: op1_00_inv03 = 1;
    20: op1_00_inv03 = 1;
    22: op1_00_inv03 = 1;
    24: op1_00_inv03 = 1;
    25: op1_00_inv03 = 1;
    27: op1_00_inv03 = 1;
    33: op1_00_inv03 = 1;
    35: op1_00_inv03 = 1;
    37: op1_00_inv03 = 1;
    39: op1_00_inv03 = 1;
    41: op1_00_inv03 = 1;
    42: op1_00_inv03 = 1;
    45: op1_00_inv03 = 1;
    48: op1_00_inv03 = 1;
    50: op1_00_inv03 = 1;
    52: op1_00_inv03 = 1;
    54: op1_00_inv03 = 1;
    61: op1_00_inv03 = 1;
    63: op1_00_inv03 = 1;
    64: op1_00_inv03 = 1;
    68: op1_00_inv03 = 1;
    69: op1_00_inv03 = 1;
    74: op1_00_inv03 = 1;
    75: op1_00_inv03 = 1;
    76: op1_00_inv03 = 1;
    79: op1_00_inv03 = 1;
    83: op1_00_inv03 = 1;
    88: op1_00_inv03 = 1;
    90: op1_00_inv03 = 1;
    93: op1_00_inv03 = 1;
    94: op1_00_inv03 = 1;
    96: op1_00_inv03 = 1;
    default: op1_00_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in04 = reg_0684;
    5: op1_00_in04 = reg_0545;
    3: op1_00_in04 = reg_0443;
    6: op1_00_in04 = imem00_in[107:104];
    29: op1_00_in04 = imem00_in[107:104];
    7: op1_00_in04 = reg_0530;
    8: op1_00_in04 = imem07_in[115:112];
    9: op1_00_in04 = reg_0123;
    10: op1_00_in04 = reg_0247;
    24: op1_00_in04 = reg_0247;
    11: op1_00_in04 = reg_0155;
    12: op1_00_in04 = imem00_in[87:84];
    46: op1_00_in04 = imem00_in[87:84];
    13: op1_00_in04 = reg_0793;
    14: op1_00_in04 = imem00_in[59:56];
    15: op1_00_in04 = reg_0677;
    16: op1_00_in04 = reg_0596;
    17: op1_00_in04 = imem05_in[123:120];
    18: op1_00_in04 = reg_0299;
    19: op1_00_in04 = reg_0153;
    20: op1_00_in04 = imem03_in[27:24];
    21: op1_00_in04 = imem06_in[123:120];
    22: op1_00_in04 = reg_0680;
    23: op1_00_in04 = reg_0278;
    25: op1_00_in04 = reg_0740;
    26: op1_00_in04 = imem00_in[103:100];
    37: op1_00_in04 = imem00_in[103:100];
    27: op1_00_in04 = reg_0801;
    28: op1_00_in04 = reg_0039;
    30: op1_00_in04 = reg_0499;
    31: op1_00_in04 = imem07_in[39:36];
    32: op1_00_in04 = reg_0678;
    33: op1_00_in04 = imem00_in[127:124];
    34: op1_00_in04 = reg_0632;
    35: op1_00_in04 = reg_0409;
    36: op1_00_in04 = imem07_in[15:12];
    38: op1_00_in04 = reg_0683;
    39: op1_00_in04 = imem02_in[47:44];
    40: op1_00_in04 = reg_0103;
    41: op1_00_in04 = reg_0068;
    42: op1_00_in04 = reg_0185;
    43: op1_00_in04 = reg_0681;
    44: op1_00_in04 = reg_0320;
    83: op1_00_in04 = reg_0320;
    45: op1_00_in04 = imem05_in[11:8];
    47: op1_00_in04 = reg_0423;
    48: op1_00_in04 = imem05_in[15:12];
    49: op1_00_in04 = reg_0129;
    50: op1_00_in04 = reg_0552;
    51: op1_00_in04 = imem02_in[107:104];
    52: op1_00_in04 = imem02_in[51:48];
    53: op1_00_in04 = imem03_in[91:88];
    54: op1_00_in04 = reg_0572;
    55: op1_00_in04 = reg_0090;
    56: op1_00_in04 = reg_0707;
    57: op1_00_in04 = reg_0620;
    58: op1_00_in04 = imem05_in[3:0];
    59: op1_00_in04 = reg_0696;
    61: op1_00_in04 = reg_0696;
    60: op1_00_in04 = imem07_in[59:56];
    62: op1_00_in04 = imem02_in[119:116];
    63: op1_00_in04 = reg_0615;
    64: op1_00_in04 = reg_0246;
    65: op1_00_in04 = imem05_in[127:124];
    66: op1_00_in04 = imem06_in[83:80];
    73: op1_00_in04 = imem06_in[83:80];
    67: op1_00_in04 = imem05_in[107:104];
    68: op1_00_in04 = reg_0240;
    69: op1_00_in04 = reg_0007;
    70: op1_00_in04 = imem07_in[11:8];
    71: op1_00_in04 = reg_0533;
    72: op1_00_in04 = reg_0276;
    74: op1_00_in04 = reg_0061;
    75: op1_00_in04 = reg_0690;
    76: op1_00_in04 = imem00_in[115:112];
    77: op1_00_in04 = imem03_in[99:96];
    89: op1_00_in04 = imem03_in[99:96];
    78: op1_00_in04 = reg_0785;
    79: op1_00_in04 = reg_0146;
    80: op1_00_in04 = imem07_in[83:80];
    82: op1_00_in04 = reg_0052;
    84: op1_00_in04 = reg_0399;
    85: op1_00_in04 = reg_0819;
    86: op1_00_in04 = reg_0829;
    87: op1_00_in04 = reg_0396;
    88: op1_00_in04 = imem07_in[7:4];
    90: op1_00_in04 = reg_0386;
    91: op1_00_in04 = reg_0618;
    92: op1_00_in04 = reg_0119;
    94: op1_00_in04 = reg_0119;
    93: op1_00_in04 = reg_0574;
    95: op1_00_in04 = reg_0077;
    96: op1_00_in04 = imem00_in[123:120];
    default: op1_00_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv04 = 1;
    5: op1_00_inv04 = 1;
    7: op1_00_inv04 = 1;
    8: op1_00_inv04 = 1;
    9: op1_00_inv04 = 1;
    10: op1_00_inv04 = 1;
    12: op1_00_inv04 = 1;
    14: op1_00_inv04 = 1;
    15: op1_00_inv04 = 1;
    16: op1_00_inv04 = 1;
    17: op1_00_inv04 = 1;
    19: op1_00_inv04 = 1;
    21: op1_00_inv04 = 1;
    24: op1_00_inv04 = 1;
    25: op1_00_inv04 = 1;
    29: op1_00_inv04 = 1;
    30: op1_00_inv04 = 1;
    31: op1_00_inv04 = 1;
    33: op1_00_inv04 = 1;
    37: op1_00_inv04 = 1;
    38: op1_00_inv04 = 1;
    39: op1_00_inv04 = 1;
    40: op1_00_inv04 = 1;
    42: op1_00_inv04 = 1;
    43: op1_00_inv04 = 1;
    45: op1_00_inv04 = 1;
    46: op1_00_inv04 = 1;
    48: op1_00_inv04 = 1;
    49: op1_00_inv04 = 1;
    50: op1_00_inv04 = 1;
    51: op1_00_inv04 = 1;
    53: op1_00_inv04 = 1;
    54: op1_00_inv04 = 1;
    57: op1_00_inv04 = 1;
    58: op1_00_inv04 = 1;
    59: op1_00_inv04 = 1;
    60: op1_00_inv04 = 1;
    61: op1_00_inv04 = 1;
    63: op1_00_inv04 = 1;
    67: op1_00_inv04 = 1;
    69: op1_00_inv04 = 1;
    70: op1_00_inv04 = 1;
    71: op1_00_inv04 = 1;
    73: op1_00_inv04 = 1;
    75: op1_00_inv04 = 1;
    76: op1_00_inv04 = 1;
    85: op1_00_inv04 = 1;
    86: op1_00_inv04 = 1;
    87: op1_00_inv04 = 1;
    95: op1_00_inv04 = 1;
    default: op1_00_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in05 = reg_0679;
    5: op1_00_in05 = reg_0551;
    3: op1_00_in05 = reg_0172;
    6: op1_00_in05 = imem00_in[123:120];
    7: op1_00_in05 = reg_0550;
    8: op1_00_in05 = reg_0722;
    9: op1_00_in05 = reg_0124;
    10: op1_00_in05 = reg_0236;
    24: op1_00_in05 = reg_0236;
    11: op1_00_in05 = imem06_in[3:0];
    12: op1_00_in05 = reg_0697;
    13: op1_00_in05 = reg_0780;
    14: op1_00_in05 = imem00_in[63:60];
    15: op1_00_in05 = reg_0678;
    16: op1_00_in05 = reg_0583;
    17: op1_00_in05 = reg_0791;
    18: op1_00_in05 = reg_0256;
    19: op1_00_in05 = reg_0134;
    20: op1_00_in05 = imem03_in[43:40];
    21: op1_00_in05 = reg_0604;
    22: op1_00_in05 = reg_0477;
    23: op1_00_in05 = reg_0079;
    25: op1_00_in05 = imem03_in[35:32];
    26: op1_00_in05 = reg_0684;
    27: op1_00_in05 = reg_0015;
    28: op1_00_in05 = reg_0814;
    29: op1_00_in05 = reg_0685;
    33: op1_00_in05 = reg_0685;
    43: op1_00_in05 = reg_0685;
    59: op1_00_in05 = reg_0685;
    30: op1_00_in05 = reg_0397;
    31: op1_00_in05 = imem07_in[43:40];
    32: op1_00_in05 = reg_0688;
    34: op1_00_in05 = reg_0623;
    35: op1_00_in05 = reg_0773;
    36: op1_00_in05 = imem07_in[59:56];
    37: op1_00_in05 = reg_0682;
    38: op1_00_in05 = reg_0681;
    39: op1_00_in05 = imem02_in[51:48];
    40: op1_00_in05 = reg_0118;
    41: op1_00_in05 = imem05_in[15:12];
    42: op1_00_in05 = reg_0173;
    44: op1_00_in05 = reg_0341;
    45: op1_00_in05 = imem05_in[27:24];
    46: op1_00_in05 = imem00_in[119:116];
    47: op1_00_in05 = reg_0054;
    48: op1_00_in05 = imem05_in[19:16];
    49: op1_00_in05 = imem06_in[59:56];
    50: op1_00_in05 = reg_0537;
    51: op1_00_in05 = imem02_in[115:112];
    52: op1_00_in05 = imem02_in[83:80];
    53: op1_00_in05 = imem03_in[103:100];
    77: op1_00_in05 = imem03_in[103:100];
    54: op1_00_in05 = reg_0376;
    55: op1_00_in05 = reg_0103;
    56: op1_00_in05 = reg_0434;
    57: op1_00_in05 = reg_0040;
    58: op1_00_in05 = imem05_in[91:88];
    60: op1_00_in05 = imem07_in[67:64];
    88: op1_00_in05 = imem07_in[67:64];
    61: op1_00_in05 = reg_0686;
    62: op1_00_in05 = imem02_in[127:124];
    63: op1_00_in05 = reg_0076;
    64: op1_00_in05 = reg_0309;
    65: op1_00_in05 = reg_0147;
    66: op1_00_in05 = imem06_in[87:84];
    67: op1_00_in05 = imem05_in[115:112];
    68: op1_00_in05 = reg_0248;
    69: op1_00_in05 = reg_0807;
    70: op1_00_in05 = imem07_in[91:88];
    71: op1_00_in05 = reg_0757;
    72: op1_00_in05 = reg_0257;
    73: op1_00_in05 = imem06_in[95:92];
    74: op1_00_in05 = reg_0446;
    75: op1_00_in05 = reg_0634;
    76: op1_00_in05 = reg_0696;
    78: op1_00_in05 = reg_0152;
    79: op1_00_in05 = reg_0641;
    82: op1_00_in05 = reg_0433;
    83: op1_00_in05 = reg_0359;
    84: op1_00_in05 = reg_0588;
    85: op1_00_in05 = reg_0657;
    86: op1_00_in05 = reg_0783;
    87: op1_00_in05 = reg_0649;
    89: op1_00_in05 = imem03_in[115:112];
    90: op1_00_in05 = reg_0399;
    91: op1_00_in05 = reg_0276;
    92: op1_00_in05 = reg_0120;
    93: op1_00_in05 = reg_0240;
    94: op1_00_in05 = reg_0660;
    95: op1_00_in05 = reg_0689;
    96: op1_00_in05 = reg_0695;
    default: op1_00_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv05 = 1;
    6: op1_00_inv05 = 1;
    8: op1_00_inv05 = 1;
    10: op1_00_inv05 = 1;
    11: op1_00_inv05 = 1;
    13: op1_00_inv05 = 1;
    14: op1_00_inv05 = 1;
    15: op1_00_inv05 = 1;
    16: op1_00_inv05 = 1;
    17: op1_00_inv05 = 1;
    24: op1_00_inv05 = 1;
    31: op1_00_inv05 = 1;
    32: op1_00_inv05 = 1;
    35: op1_00_inv05 = 1;
    42: op1_00_inv05 = 1;
    46: op1_00_inv05 = 1;
    47: op1_00_inv05 = 1;
    48: op1_00_inv05 = 1;
    51: op1_00_inv05 = 1;
    54: op1_00_inv05 = 1;
    55: op1_00_inv05 = 1;
    56: op1_00_inv05 = 1;
    59: op1_00_inv05 = 1;
    64: op1_00_inv05 = 1;
    66: op1_00_inv05 = 1;
    67: op1_00_inv05 = 1;
    68: op1_00_inv05 = 1;
    69: op1_00_inv05 = 1;
    70: op1_00_inv05 = 1;
    73: op1_00_inv05 = 1;
    74: op1_00_inv05 = 1;
    75: op1_00_inv05 = 1;
    76: op1_00_inv05 = 1;
    79: op1_00_inv05 = 1;
    83: op1_00_inv05 = 1;
    87: op1_00_inv05 = 1;
    88: op1_00_inv05 = 1;
    91: op1_00_inv05 = 1;
    default: op1_00_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in06 = reg_0668;
    5: op1_00_in06 = reg_0281;
    3: op1_00_in06 = reg_0157;
    6: op1_00_in06 = reg_0689;
    7: op1_00_in06 = reg_0548;
    8: op1_00_in06 = reg_0709;
    9: op1_00_in06 = reg_0103;
    10: op1_00_in06 = reg_0245;
    24: op1_00_in06 = reg_0245;
    11: op1_00_in06 = imem06_in[115:112];
    12: op1_00_in06 = reg_0451;
    13: op1_00_in06 = reg_0786;
    14: op1_00_in06 = imem00_in[83:80];
    15: op1_00_in06 = reg_0673;
    16: op1_00_in06 = reg_0572;
    17: op1_00_in06 = reg_0792;
    18: op1_00_in06 = imem05_in[87:84];
    45: op1_00_in06 = imem05_in[87:84];
    19: op1_00_in06 = imem06_in[7:4];
    20: op1_00_in06 = imem03_in[55:52];
    21: op1_00_in06 = reg_0609;
    22: op1_00_in06 = reg_0481;
    23: op1_00_in06 = reg_0066;
    25: op1_00_in06 = imem03_in[47:44];
    26: op1_00_in06 = reg_0677;
    27: op1_00_in06 = reg_0010;
    28: op1_00_in06 = reg_0037;
    29: op1_00_in06 = reg_0694;
    30: op1_00_in06 = reg_0013;
    31: op1_00_in06 = imem07_in[51:48];
    32: op1_00_in06 = reg_0463;
    33: op1_00_in06 = reg_0674;
    34: op1_00_in06 = reg_0317;
    35: op1_00_in06 = reg_0270;
    36: op1_00_in06 = imem07_in[91:88];
    37: op1_00_in06 = reg_0697;
    38: op1_00_in06 = reg_0685;
    39: op1_00_in06 = imem02_in[95:92];
    40: op1_00_in06 = reg_0116;
    41: op1_00_in06 = imem05_in[39:36];
    43: op1_00_in06 = reg_0684;
    59: op1_00_in06 = reg_0684;
    44: op1_00_in06 = reg_0353;
    46: op1_00_in06 = reg_0672;
    47: op1_00_in06 = reg_0567;
    48: op1_00_in06 = imem05_in[31:28];
    49: op1_00_in06 = reg_0625;
    50: op1_00_in06 = reg_0055;
    51: op1_00_in06 = reg_0518;
    52: op1_00_in06 = imem02_in[115:112];
    53: op1_00_in06 = reg_0387;
    54: op1_00_in06 = reg_0393;
    55: op1_00_in06 = reg_0249;
    56: op1_00_in06 = reg_0084;
    57: op1_00_in06 = imem07_in[11:8];
    58: op1_00_in06 = imem05_in[95:92];
    60: op1_00_in06 = imem07_in[71:68];
    61: op1_00_in06 = reg_0688;
    62: op1_00_in06 = reg_0362;
    63: op1_00_in06 = reg_0529;
    64: op1_00_in06 = reg_0229;
    65: op1_00_in06 = reg_0136;
    66: op1_00_in06 = imem06_in[95:92];
    67: op1_00_in06 = reg_0386;
    68: op1_00_in06 = reg_0234;
    69: op1_00_in06 = reg_0799;
    70: op1_00_in06 = imem07_in[99:96];
    88: op1_00_in06 = imem07_in[99:96];
    71: op1_00_in06 = imem03_in[43:40];
    72: op1_00_in06 = reg_0307;
    73: op1_00_in06 = reg_0299;
    74: op1_00_in06 = reg_0165;
    75: op1_00_in06 = reg_0465;
    76: op1_00_in06 = reg_0492;
    77: op1_00_in06 = imem03_in[111:108];
    78: op1_00_in06 = reg_0830;
    79: op1_00_in06 = reg_0782;
    82: op1_00_in06 = reg_0076;
    83: op1_00_in06 = reg_0324;
    84: op1_00_in06 = reg_0648;
    85: op1_00_in06 = reg_0752;
    86: op1_00_in06 = reg_0765;
    87: op1_00_in06 = reg_0570;
    89: op1_00_in06 = imem04_in[71:68];
    90: op1_00_in06 = reg_0531;
    91: op1_00_in06 = reg_0484;
    92: op1_00_in06 = reg_0675;
    93: op1_00_in06 = reg_0051;
    94: op1_00_in06 = reg_0669;
    95: op1_00_in06 = reg_0749;
    96: op1_00_in06 = reg_0693;
    default: op1_00_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv06 = 1;
    7: op1_00_inv06 = 1;
    10: op1_00_inv06 = 1;
    12: op1_00_inv06 = 1;
    14: op1_00_inv06 = 1;
    17: op1_00_inv06 = 1;
    18: op1_00_inv06 = 1;
    19: op1_00_inv06 = 1;
    20: op1_00_inv06 = 1;
    24: op1_00_inv06 = 1;
    25: op1_00_inv06 = 1;
    27: op1_00_inv06 = 1;
    30: op1_00_inv06 = 1;
    32: op1_00_inv06 = 1;
    33: op1_00_inv06 = 1;
    37: op1_00_inv06 = 1;
    41: op1_00_inv06 = 1;
    46: op1_00_inv06 = 1;
    47: op1_00_inv06 = 1;
    48: op1_00_inv06 = 1;
    49: op1_00_inv06 = 1;
    51: op1_00_inv06 = 1;
    53: op1_00_inv06 = 1;
    55: op1_00_inv06 = 1;
    56: op1_00_inv06 = 1;
    59: op1_00_inv06 = 1;
    60: op1_00_inv06 = 1;
    62: op1_00_inv06 = 1;
    63: op1_00_inv06 = 1;
    65: op1_00_inv06 = 1;
    68: op1_00_inv06 = 1;
    70: op1_00_inv06 = 1;
    71: op1_00_inv06 = 1;
    73: op1_00_inv06 = 1;
    74: op1_00_inv06 = 1;
    75: op1_00_inv06 = 1;
    76: op1_00_inv06 = 1;
    79: op1_00_inv06 = 1;
    84: op1_00_inv06 = 1;
    85: op1_00_inv06 = 1;
    88: op1_00_inv06 = 1;
    92: op1_00_inv06 = 1;
    93: op1_00_inv06 = 1;
    95: op1_00_inv06 = 1;
    default: op1_00_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in07 = reg_0680;
    26: op1_00_in07 = reg_0680;
    5: op1_00_in07 = reg_0305;
    3: op1_00_in07 = reg_0173;
    6: op1_00_in07 = reg_0677;
    7: op1_00_in07 = reg_0549;
    8: op1_00_in07 = reg_0421;
    9: op1_00_in07 = reg_0116;
    10: op1_00_in07 = reg_0238;
    11: op1_00_in07 = imem06_in[119:116];
    12: op1_00_in07 = reg_0462;
    13: op1_00_in07 = reg_0268;
    14: op1_00_in07 = imem00_in[115:112];
    15: op1_00_in07 = reg_0457;
    16: op1_00_in07 = reg_0593;
    17: op1_00_in07 = reg_0488;
    18: op1_00_in07 = imem05_in[107:104];
    19: op1_00_in07 = imem06_in[23:20];
    20: op1_00_in07 = imem03_in[87:84];
    21: op1_00_in07 = reg_0611;
    22: op1_00_in07 = reg_0480;
    23: op1_00_in07 = reg_0071;
    24: op1_00_in07 = reg_0041;
    25: op1_00_in07 = imem03_in[51:48];
    27: op1_00_in07 = imem04_in[7:4];
    28: op1_00_in07 = reg_0750;
    29: op1_00_in07 = reg_0668;
    30: op1_00_in07 = reg_0800;
    31: op1_00_in07 = imem07_in[71:68];
    32: op1_00_in07 = reg_0454;
    33: op1_00_in07 = reg_0463;
    34: op1_00_in07 = reg_0763;
    35: op1_00_in07 = reg_0404;
    36: op1_00_in07 = imem07_in[111:108];
    37: op1_00_in07 = reg_0690;
    38: op1_00_in07 = reg_0684;
    39: op1_00_in07 = imem02_in[127:124];
    40: op1_00_in07 = reg_0120;
    41: op1_00_in07 = imem05_in[47:44];
    43: op1_00_in07 = reg_0674;
    44: op1_00_in07 = reg_0323;
    45: op1_00_in07 = imem05_in[123:120];
    46: op1_00_in07 = reg_0686;
    59: op1_00_in07 = reg_0686;
    76: op1_00_in07 = reg_0686;
    47: op1_00_in07 = reg_0234;
    48: op1_00_in07 = imem05_in[43:40];
    49: op1_00_in07 = reg_0604;
    50: op1_00_in07 = reg_0060;
    51: op1_00_in07 = reg_0092;
    52: op1_00_in07 = reg_0637;
    53: op1_00_in07 = reg_0575;
    54: op1_00_in07 = reg_0570;
    55: op1_00_in07 = reg_0285;
    56: op1_00_in07 = reg_0438;
    57: op1_00_in07 = imem07_in[35:32];
    58: op1_00_in07 = imem05_in[99:96];
    60: op1_00_in07 = imem07_in[91:88];
    61: op1_00_in07 = reg_0455;
    62: op1_00_in07 = reg_0359;
    63: op1_00_in07 = reg_0077;
    64: op1_00_in07 = reg_0145;
    65: op1_00_in07 = reg_0152;
    66: op1_00_in07 = reg_0289;
    67: op1_00_in07 = reg_0075;
    68: op1_00_in07 = reg_0506;
    69: op1_00_in07 = reg_0016;
    70: op1_00_in07 = reg_0716;
    71: op1_00_in07 = imem03_in[47:44];
    72: op1_00_in07 = reg_0783;
    73: op1_00_in07 = reg_0577;
    74: op1_00_in07 = reg_0159;
    75: op1_00_in07 = reg_0464;
    77: op1_00_in07 = reg_0599;
    78: op1_00_in07 = reg_0143;
    79: op1_00_in07 = reg_0665;
    82: op1_00_in07 = reg_0529;
    83: op1_00_in07 = reg_0406;
    84: op1_00_in07 = reg_0395;
    85: op1_00_in07 = reg_0367;
    86: op1_00_in07 = imem06_in[3:0];
    87: op1_00_in07 = reg_0000;
    88: op1_00_in07 = imem07_in[103:100];
    89: op1_00_in07 = imem04_in[119:116];
    90: op1_00_in07 = reg_0547;
    91: op1_00_in07 = reg_0608;
    92: op1_00_in07 = reg_0106;
    93: op1_00_in07 = reg_0054;
    94: op1_00_in07 = reg_0601;
    95: op1_00_in07 = reg_0130;
    96: op1_00_in07 = reg_0189;
    default: op1_00_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv07 = 1;
    3: op1_00_inv07 = 1;
    6: op1_00_inv07 = 1;
    11: op1_00_inv07 = 1;
    12: op1_00_inv07 = 1;
    14: op1_00_inv07 = 1;
    16: op1_00_inv07 = 1;
    18: op1_00_inv07 = 1;
    24: op1_00_inv07 = 1;
    27: op1_00_inv07 = 1;
    28: op1_00_inv07 = 1;
    29: op1_00_inv07 = 1;
    30: op1_00_inv07 = 1;
    31: op1_00_inv07 = 1;
    32: op1_00_inv07 = 1;
    37: op1_00_inv07 = 1;
    40: op1_00_inv07 = 1;
    41: op1_00_inv07 = 1;
    43: op1_00_inv07 = 1;
    44: op1_00_inv07 = 1;
    45: op1_00_inv07 = 1;
    46: op1_00_inv07 = 1;
    47: op1_00_inv07 = 1;
    50: op1_00_inv07 = 1;
    52: op1_00_inv07 = 1;
    54: op1_00_inv07 = 1;
    57: op1_00_inv07 = 1;
    58: op1_00_inv07 = 1;
    59: op1_00_inv07 = 1;
    61: op1_00_inv07 = 1;
    62: op1_00_inv07 = 1;
    64: op1_00_inv07 = 1;
    67: op1_00_inv07 = 1;
    68: op1_00_inv07 = 1;
    70: op1_00_inv07 = 1;
    71: op1_00_inv07 = 1;
    72: op1_00_inv07 = 1;
    73: op1_00_inv07 = 1;
    74: op1_00_inv07 = 1;
    75: op1_00_inv07 = 1;
    78: op1_00_inv07 = 1;
    79: op1_00_inv07 = 1;
    83: op1_00_inv07 = 1;
    86: op1_00_inv07 = 1;
    87: op1_00_inv07 = 1;
    88: op1_00_inv07 = 1;
    89: op1_00_inv07 = 1;
    90: op1_00_inv07 = 1;
    91: op1_00_inv07 = 1;
    93: op1_00_inv07 = 1;
    94: op1_00_inv07 = 1;
    95: op1_00_inv07 = 1;
    96: op1_00_inv07 = 1;
    default: op1_00_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in08 = reg_0688;
    5: op1_00_in08 = reg_0277;
    6: op1_00_in08 = reg_0453;
    7: op1_00_in08 = reg_0554;
    8: op1_00_in08 = reg_0426;
    9: op1_00_in08 = reg_0099;
    10: op1_00_in08 = reg_0243;
    24: op1_00_in08 = reg_0243;
    11: op1_00_in08 = reg_0625;
    12: op1_00_in08 = reg_0467;
    13: op1_00_in08 = reg_0259;
    14: op1_00_in08 = reg_0679;
    15: op1_00_in08 = reg_0479;
    16: op1_00_in08 = reg_0321;
    17: op1_00_in08 = reg_0526;
    18: op1_00_in08 = reg_0796;
    19: op1_00_in08 = imem06_in[27:24];
    86: op1_00_in08 = imem06_in[27:24];
    20: op1_00_in08 = imem03_in[99:96];
    21: op1_00_in08 = reg_0632;
    22: op1_00_in08 = reg_0452;
    23: op1_00_in08 = imem05_in[11:8];
    25: op1_00_in08 = imem03_in[79:76];
    26: op1_00_in08 = reg_0692;
    38: op1_00_in08 = reg_0692;
    27: op1_00_in08 = imem04_in[15:12];
    28: op1_00_in08 = reg_0005;
    29: op1_00_in08 = reg_0673;
    30: op1_00_in08 = reg_0014;
    31: op1_00_in08 = imem07_in[79:76];
    32: op1_00_in08 = reg_0466;
    75: op1_00_in08 = reg_0466;
    33: op1_00_in08 = reg_0450;
    34: op1_00_in08 = reg_0403;
    35: op1_00_in08 = reg_0319;
    36: op1_00_in08 = reg_0704;
    37: op1_00_in08 = reg_0475;
    39: op1_00_in08 = reg_0650;
    40: op1_00_in08 = reg_0112;
    41: op1_00_in08 = imem05_in[87:84];
    48: op1_00_in08 = imem05_in[87:84];
    43: op1_00_in08 = reg_0675;
    44: op1_00_in08 = reg_0095;
    51: op1_00_in08 = reg_0095;
    45: op1_00_in08 = reg_0791;
    46: op1_00_in08 = reg_0677;
    47: op1_00_in08 = reg_0506;
    49: op1_00_in08 = reg_0291;
    50: op1_00_in08 = reg_0523;
    52: op1_00_in08 = reg_0355;
    53: op1_00_in08 = reg_0572;
    54: op1_00_in08 = reg_0002;
    55: op1_00_in08 = reg_0143;
    56: op1_00_in08 = reg_0448;
    57: op1_00_in08 = imem07_in[51:48];
    58: op1_00_in08 = imem05_in[119:116];
    59: op1_00_in08 = reg_0690;
    60: op1_00_in08 = reg_0728;
    61: op1_00_in08 = reg_0474;
    62: op1_00_in08 = reg_0342;
    63: op1_00_in08 = reg_0629;
    64: op1_00_in08 = reg_0135;
    65: op1_00_in08 = reg_0142;
    66: op1_00_in08 = reg_0348;
    67: op1_00_in08 = reg_0491;
    68: op1_00_in08 = reg_0424;
    69: op1_00_in08 = reg_0806;
    70: op1_00_in08 = reg_0720;
    71: op1_00_in08 = imem03_in[59:56];
    72: op1_00_in08 = reg_0147;
    73: op1_00_in08 = reg_0605;
    74: op1_00_in08 = reg_0177;
    76: op1_00_in08 = reg_0758;
    77: op1_00_in08 = reg_0595;
    78: op1_00_in08 = reg_0153;
    79: op1_00_in08 = reg_0517;
    82: op1_00_in08 = reg_0302;
    83: op1_00_in08 = reg_0514;
    84: op1_00_in08 = reg_0028;
    85: op1_00_in08 = imem07_in[11:8];
    87: op1_00_in08 = reg_0807;
    88: op1_00_in08 = reg_0716;
    89: op1_00_in08 = reg_0262;
    90: op1_00_in08 = reg_0149;
    91: op1_00_in08 = reg_0638;
    92: op1_00_in08 = reg_0669;
    93: op1_00_in08 = reg_0124;
    94: op1_00_in08 = reg_0671;
    95: op1_00_in08 = reg_0171;
    96: op1_00_in08 = reg_0163;
    default: op1_00_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv08 = 1;
    5: op1_00_inv08 = 1;
    6: op1_00_inv08 = 1;
    8: op1_00_inv08 = 1;
    10: op1_00_inv08 = 1;
    13: op1_00_inv08 = 1;
    14: op1_00_inv08 = 1;
    15: op1_00_inv08 = 1;
    17: op1_00_inv08 = 1;
    20: op1_00_inv08 = 1;
    21: op1_00_inv08 = 1;
    23: op1_00_inv08 = 1;
    24: op1_00_inv08 = 1;
    25: op1_00_inv08 = 1;
    26: op1_00_inv08 = 1;
    29: op1_00_inv08 = 1;
    30: op1_00_inv08 = 1;
    34: op1_00_inv08 = 1;
    35: op1_00_inv08 = 1;
    36: op1_00_inv08 = 1;
    37: op1_00_inv08 = 1;
    38: op1_00_inv08 = 1;
    41: op1_00_inv08 = 1;
    44: op1_00_inv08 = 1;
    45: op1_00_inv08 = 1;
    46: op1_00_inv08 = 1;
    47: op1_00_inv08 = 1;
    50: op1_00_inv08 = 1;
    53: op1_00_inv08 = 1;
    54: op1_00_inv08 = 1;
    55: op1_00_inv08 = 1;
    56: op1_00_inv08 = 1;
    57: op1_00_inv08 = 1;
    59: op1_00_inv08 = 1;
    60: op1_00_inv08 = 1;
    62: op1_00_inv08 = 1;
    64: op1_00_inv08 = 1;
    65: op1_00_inv08 = 1;
    66: op1_00_inv08 = 1;
    67: op1_00_inv08 = 1;
    69: op1_00_inv08 = 1;
    70: op1_00_inv08 = 1;
    72: op1_00_inv08 = 1;
    74: op1_00_inv08 = 1;
    76: op1_00_inv08 = 1;
    78: op1_00_inv08 = 1;
    79: op1_00_inv08 = 1;
    83: op1_00_inv08 = 1;
    84: op1_00_inv08 = 1;
    85: op1_00_inv08 = 1;
    92: op1_00_inv08 = 1;
    93: op1_00_inv08 = 1;
    95: op1_00_inv08 = 1;
    default: op1_00_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in09 = reg_0673;
    93: op1_00_in09 = reg_0673;
    5: op1_00_in09 = reg_0306;
    6: op1_00_in09 = reg_0200;
    7: op1_00_in09 = reg_0546;
    8: op1_00_in09 = reg_0418;
    9: op1_00_in09 = reg_0112;
    10: op1_00_in09 = reg_0122;
    68: op1_00_in09 = reg_0122;
    11: op1_00_in09 = reg_0612;
    12: op1_00_in09 = reg_0479;
    13: op1_00_in09 = reg_0273;
    14: op1_00_in09 = reg_0691;
    46: op1_00_in09 = reg_0691;
    15: op1_00_in09 = reg_0478;
    16: op1_00_in09 = reg_0311;
    17: op1_00_in09 = reg_0147;
    18: op1_00_in09 = reg_0789;
    19: op1_00_in09 = imem06_in[91:88];
    20: op1_00_in09 = imem03_in[107:104];
    21: op1_00_in09 = reg_0622;
    22: op1_00_in09 = reg_0214;
    23: op1_00_in09 = imem05_in[19:16];
    24: op1_00_in09 = reg_0249;
    25: op1_00_in09 = imem03_in[103:100];
    26: op1_00_in09 = reg_0457;
    38: op1_00_in09 = reg_0457;
    27: op1_00_in09 = imem04_in[51:48];
    28: op1_00_in09 = imem07_in[23:20];
    29: op1_00_in09 = reg_0477;
    30: op1_00_in09 = reg_0799;
    31: op1_00_in09 = imem07_in[115:112];
    32: op1_00_in09 = reg_0462;
    33: op1_00_in09 = reg_0476;
    34: op1_00_in09 = reg_0776;
    35: op1_00_in09 = reg_0406;
    36: op1_00_in09 = reg_0719;
    60: op1_00_in09 = reg_0719;
    37: op1_00_in09 = reg_0480;
    39: op1_00_in09 = reg_0645;
    40: op1_00_in09 = reg_0108;
    41: op1_00_in09 = imem05_in[107:104];
    43: op1_00_in09 = reg_0687;
    44: op1_00_in09 = reg_0082;
    45: op1_00_in09 = reg_0488;
    47: op1_00_in09 = reg_0243;
    48: op1_00_in09 = imem05_in[95:92];
    49: op1_00_in09 = reg_0605;
    50: op1_00_in09 = reg_0516;
    51: op1_00_in09 = reg_0540;
    52: op1_00_in09 = reg_0365;
    53: op1_00_in09 = reg_0570;
    54: op1_00_in09 = reg_0807;
    55: op1_00_in09 = imem06_in[27:24];
    56: op1_00_in09 = reg_0175;
    57: op1_00_in09 = imem07_in[59:56];
    58: op1_00_in09 = reg_0798;
    59: op1_00_in09 = reg_0658;
    61: op1_00_in09 = reg_0459;
    62: op1_00_in09 = reg_0590;
    63: op1_00_in09 = reg_0643;
    64: op1_00_in09 = reg_0128;
    65: op1_00_in09 = reg_0156;
    66: op1_00_in09 = reg_0346;
    67: op1_00_in09 = reg_0257;
    69: op1_00_in09 = reg_0009;
    70: op1_00_in09 = reg_0726;
    88: op1_00_in09 = reg_0726;
    71: op1_00_in09 = imem03_in[75:72];
    72: op1_00_in09 = reg_0148;
    73: op1_00_in09 = reg_0370;
    74: op1_00_in09 = reg_0164;
    75: op1_00_in09 = reg_0475;
    76: op1_00_in09 = reg_0247;
    77: op1_00_in09 = reg_0588;
    78: op1_00_in09 = reg_0761;
    90: op1_00_in09 = reg_0761;
    79: op1_00_in09 = reg_0075;
    82: op1_00_in09 = reg_0074;
    83: op1_00_in09 = reg_0092;
    84: op1_00_in09 = reg_0368;
    85: op1_00_in09 = imem07_in[43:40];
    86: op1_00_in09 = imem06_in[83:80];
    87: op1_00_in09 = reg_0804;
    89: op1_00_in09 = reg_0058;
    91: op1_00_in09 = reg_0777;
    92: op1_00_in09 = reg_0678;
    94: op1_00_in09 = reg_0121;
    95: op1_00_in09 = reg_0070;
    96: op1_00_in09 = reg_0686;
    default: op1_00_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv09 = 1;
    7: op1_00_inv09 = 1;
    10: op1_00_inv09 = 1;
    12: op1_00_inv09 = 1;
    14: op1_00_inv09 = 1;
    16: op1_00_inv09 = 1;
    17: op1_00_inv09 = 1;
    20: op1_00_inv09 = 1;
    23: op1_00_inv09 = 1;
    26: op1_00_inv09 = 1;
    32: op1_00_inv09 = 1;
    34: op1_00_inv09 = 1;
    36: op1_00_inv09 = 1;
    39: op1_00_inv09 = 1;
    40: op1_00_inv09 = 1;
    44: op1_00_inv09 = 1;
    46: op1_00_inv09 = 1;
    47: op1_00_inv09 = 1;
    49: op1_00_inv09 = 1;
    53: op1_00_inv09 = 1;
    54: op1_00_inv09 = 1;
    56: op1_00_inv09 = 1;
    65: op1_00_inv09 = 1;
    66: op1_00_inv09 = 1;
    72: op1_00_inv09 = 1;
    74: op1_00_inv09 = 1;
    75: op1_00_inv09 = 1;
    79: op1_00_inv09 = 1;
    82: op1_00_inv09 = 1;
    85: op1_00_inv09 = 1;
    87: op1_00_inv09 = 1;
    89: op1_00_inv09 = 1;
    92: op1_00_inv09 = 1;
    default: op1_00_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in10 = reg_0669;
    5: op1_00_in10 = reg_0292;
    6: op1_00_in10 = reg_0189;
    7: op1_00_in10 = reg_0558;
    8: op1_00_in10 = reg_0445;
    9: op1_00_in10 = reg_0108;
    10: op1_00_in10 = reg_0119;
    24: op1_00_in10 = reg_0119;
    47: op1_00_in10 = reg_0119;
    11: op1_00_in10 = reg_0402;
    12: op1_00_in10 = reg_0459;
    33: op1_00_in10 = reg_0459;
    75: op1_00_in10 = reg_0459;
    13: op1_00_in10 = reg_0042;
    14: op1_00_in10 = reg_0678;
    15: op1_00_in10 = reg_0208;
    16: op1_00_in10 = reg_0385;
    17: op1_00_in10 = reg_0136;
    18: op1_00_in10 = reg_0491;
    19: op1_00_in10 = reg_0620;
    20: op1_00_in10 = reg_0569;
    21: op1_00_in10 = reg_0405;
    22: op1_00_in10 = reg_0193;
    23: op1_00_in10 = imem05_in[31:28];
    25: op1_00_in10 = imem03_in[115:112];
    26: op1_00_in10 = reg_0466;
    27: op1_00_in10 = imem04_in[91:88];
    28: op1_00_in10 = imem07_in[27:24];
    29: op1_00_in10 = reg_0456;
    30: op1_00_in10 = reg_0016;
    31: op1_00_in10 = imem07_in[127:124];
    32: op1_00_in10 = reg_0480;
    34: op1_00_in10 = reg_0604;
    35: op1_00_in10 = reg_0814;
    36: op1_00_in10 = reg_0700;
    37: op1_00_in10 = reg_0473;
    38: op1_00_in10 = reg_0461;
    39: op1_00_in10 = reg_0646;
    40: op1_00_in10 = reg_0110;
    41: op1_00_in10 = reg_0791;
    43: op1_00_in10 = reg_0454;
    44: op1_00_in10 = reg_0539;
    45: op1_00_in10 = reg_0793;
    46: op1_00_in10 = reg_0674;
    48: op1_00_in10 = imem05_in[103:100];
    49: op1_00_in10 = reg_0608;
    50: op1_00_in10 = reg_0357;
    51: op1_00_in10 = reg_0770;
    52: op1_00_in10 = reg_0541;
    53: op1_00_in10 = reg_0803;
    54: op1_00_in10 = reg_0804;
    55: op1_00_in10 = imem06_in[35:32];
    56: op1_00_in10 = reg_0164;
    57: op1_00_in10 = imem07_in[71:68];
    58: op1_00_in10 = reg_0111;
    59: op1_00_in10 = reg_0407;
    60: op1_00_in10 = reg_0720;
    61: op1_00_in10 = reg_0191;
    62: op1_00_in10 = reg_0514;
    63: op1_00_in10 = reg_0771;
    64: op1_00_in10 = reg_0152;
    65: op1_00_in10 = reg_0144;
    66: op1_00_in10 = reg_0291;
    67: op1_00_in10 = reg_0307;
    68: op1_00_in10 = reg_0671;
    69: op1_00_in10 = imem04_in[11:8];
    70: op1_00_in10 = reg_0705;
    71: op1_00_in10 = imem03_in[103:100];
    72: op1_00_in10 = reg_0150;
    73: op1_00_in10 = reg_0354;
    76: op1_00_in10 = reg_0453;
    77: op1_00_in10 = reg_0331;
    78: op1_00_in10 = imem06_in[23:20];
    79: op1_00_in10 = reg_0486;
    82: op1_00_in10 = reg_0065;
    83: op1_00_in10 = reg_0096;
    84: op1_00_in10 = reg_0562;
    85: op1_00_in10 = imem07_in[47:44];
    86: op1_00_in10 = imem06_in[95:92];
    87: op1_00_in10 = imem04_in[15:12];
    88: op1_00_in10 = reg_0784;
    89: op1_00_in10 = reg_0179;
    90: op1_00_in10 = imem06_in[71:68];
    91: op1_00_in10 = reg_0609;
    92: op1_00_in10 = imem02_in[23:20];
    93: op1_00_in10 = reg_0670;
    94: op1_00_in10 = imem02_in[31:28];
    95: op1_00_in10 = reg_0692;
    96: op1_00_in10 = reg_0131;
    default: op1_00_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_00_inv10 = 1;
    9: op1_00_inv10 = 1;
    11: op1_00_inv10 = 1;
    12: op1_00_inv10 = 1;
    14: op1_00_inv10 = 1;
    16: op1_00_inv10 = 1;
    17: op1_00_inv10 = 1;
    19: op1_00_inv10 = 1;
    20: op1_00_inv10 = 1;
    21: op1_00_inv10 = 1;
    22: op1_00_inv10 = 1;
    23: op1_00_inv10 = 1;
    25: op1_00_inv10 = 1;
    26: op1_00_inv10 = 1;
    27: op1_00_inv10 = 1;
    28: op1_00_inv10 = 1;
    33: op1_00_inv10 = 1;
    36: op1_00_inv10 = 1;
    40: op1_00_inv10 = 1;
    45: op1_00_inv10 = 1;
    46: op1_00_inv10 = 1;
    50: op1_00_inv10 = 1;
    52: op1_00_inv10 = 1;
    54: op1_00_inv10 = 1;
    58: op1_00_inv10 = 1;
    59: op1_00_inv10 = 1;
    61: op1_00_inv10 = 1;
    66: op1_00_inv10 = 1;
    67: op1_00_inv10 = 1;
    68: op1_00_inv10 = 1;
    69: op1_00_inv10 = 1;
    71: op1_00_inv10 = 1;
    73: op1_00_inv10 = 1;
    75: op1_00_inv10 = 1;
    78: op1_00_inv10 = 1;
    82: op1_00_inv10 = 1;
    84: op1_00_inv10 = 1;
    91: op1_00_inv10 = 1;
    93: op1_00_inv10 = 1;
    94: op1_00_inv10 = 1;
    95: op1_00_inv10 = 1;
    96: op1_00_inv10 = 1;
    default: op1_00_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in11 = reg_0465;
    95: op1_00_in11 = reg_0465;
    5: op1_00_in11 = reg_0275;
    6: op1_00_in11 = reg_0204;
    7: op1_00_in11 = reg_0304;
    8: op1_00_in11 = reg_0446;
    9: op1_00_in11 = reg_0114;
    10: op1_00_in11 = reg_0112;
    11: op1_00_in11 = reg_0405;
    12: op1_00_in11 = reg_0214;
    13: op1_00_in11 = reg_0735;
    14: op1_00_in11 = reg_0668;
    15: op1_00_in11 = reg_0188;
    16: op1_00_in11 = reg_0376;
    17: op1_00_in11 = reg_0142;
    64: op1_00_in11 = reg_0142;
    18: op1_00_in11 = reg_0785;
    19: op1_00_in11 = reg_0621;
    20: op1_00_in11 = reg_0563;
    21: op1_00_in11 = reg_0404;
    22: op1_00_in11 = reg_0201;
    33: op1_00_in11 = reg_0201;
    23: op1_00_in11 = imem05_in[59:56];
    24: op1_00_in11 = reg_0110;
    25: op1_00_in11 = reg_0583;
    26: op1_00_in11 = reg_0467;
    27: op1_00_in11 = imem04_in[103:100];
    28: op1_00_in11 = imem07_in[31:28];
    29: op1_00_in11 = reg_0458;
    30: op1_00_in11 = reg_0004;
    31: op1_00_in11 = reg_0729;
    32: op1_00_in11 = reg_0473;
    34: op1_00_in11 = reg_0777;
    35: op1_00_in11 = reg_0372;
    36: op1_00_in11 = reg_0419;
    37: op1_00_in11 = reg_0468;
    38: op1_00_in11 = reg_0460;
    39: op1_00_in11 = reg_0638;
    40: op1_00_in11 = imem02_in[19:16];
    41: op1_00_in11 = reg_0796;
    43: op1_00_in11 = reg_0466;
    44: op1_00_in11 = reg_0098;
    45: op1_00_in11 = reg_0790;
    46: op1_00_in11 = reg_0671;
    47: op1_00_in11 = reg_0108;
    48: op1_00_in11 = imem05_in[115:112];
    49: op1_00_in11 = reg_0622;
    50: op1_00_in11 = reg_0078;
    51: op1_00_in11 = reg_0082;
    52: op1_00_in11 = reg_0097;
    53: op1_00_in11 = reg_0800;
    54: op1_00_in11 = reg_0008;
    55: op1_00_in11 = imem06_in[59:56];
    56: op1_00_in11 = reg_0157;
    57: op1_00_in11 = imem07_in[83:80];
    58: op1_00_in11 = reg_0752;
    59: op1_00_in11 = reg_0494;
    60: op1_00_in11 = reg_0730;
    61: op1_00_in11 = reg_0210;
    62: op1_00_in11 = reg_0532;
    63: op1_00_in11 = reg_0776;
    65: op1_00_in11 = imem06_in[3:0];
    66: op1_00_in11 = reg_0624;
    67: op1_00_in11 = reg_0135;
    68: op1_00_in11 = imem02_in[31:28];
    69: op1_00_in11 = imem04_in[59:56];
    70: op1_00_in11 = reg_0441;
    71: op1_00_in11 = reg_0602;
    72: op1_00_in11 = imem06_in[7:4];
    73: op1_00_in11 = reg_0377;
    75: op1_00_in11 = reg_0209;
    76: op1_00_in11 = reg_0457;
    77: op1_00_in11 = reg_0417;
    78: op1_00_in11 = imem06_in[63:60];
    79: op1_00_in11 = reg_0500;
    82: op1_00_in11 = reg_0513;
    83: op1_00_in11 = reg_0770;
    84: op1_00_in11 = reg_0637;
    85: op1_00_in11 = imem07_in[51:48];
    86: op1_00_in11 = imem06_in[103:100];
    87: op1_00_in11 = imem04_in[19:16];
    88: op1_00_in11 = reg_0382;
    89: op1_00_in11 = reg_0060;
    90: op1_00_in11 = imem06_in[83:80];
    91: op1_00_in11 = reg_0501;
    92: op1_00_in11 = imem02_in[107:104];
    93: op1_00_in11 = reg_0675;
    94: op1_00_in11 = imem02_in[39:36];
    96: op1_00_in11 = reg_0688;
    default: op1_00_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv11 = 1;
    5: op1_00_inv11 = 1;
    6: op1_00_inv11 = 1;
    7: op1_00_inv11 = 1;
    8: op1_00_inv11 = 1;
    9: op1_00_inv11 = 1;
    10: op1_00_inv11 = 1;
    11: op1_00_inv11 = 1;
    14: op1_00_inv11 = 1;
    15: op1_00_inv11 = 1;
    16: op1_00_inv11 = 1;
    17: op1_00_inv11 = 1;
    18: op1_00_inv11 = 1;
    20: op1_00_inv11 = 1;
    22: op1_00_inv11 = 1;
    23: op1_00_inv11 = 1;
    26: op1_00_inv11 = 1;
    27: op1_00_inv11 = 1;
    28: op1_00_inv11 = 1;
    29: op1_00_inv11 = 1;
    33: op1_00_inv11 = 1;
    34: op1_00_inv11 = 1;
    37: op1_00_inv11 = 1;
    40: op1_00_inv11 = 1;
    43: op1_00_inv11 = 1;
    44: op1_00_inv11 = 1;
    45: op1_00_inv11 = 1;
    50: op1_00_inv11 = 1;
    52: op1_00_inv11 = 1;
    53: op1_00_inv11 = 1;
    54: op1_00_inv11 = 1;
    56: op1_00_inv11 = 1;
    57: op1_00_inv11 = 1;
    58: op1_00_inv11 = 1;
    62: op1_00_inv11 = 1;
    64: op1_00_inv11 = 1;
    65: op1_00_inv11 = 1;
    66: op1_00_inv11 = 1;
    68: op1_00_inv11 = 1;
    71: op1_00_inv11 = 1;
    73: op1_00_inv11 = 1;
    75: op1_00_inv11 = 1;
    77: op1_00_inv11 = 1;
    78: op1_00_inv11 = 1;
    83: op1_00_inv11 = 1;
    84: op1_00_inv11 = 1;
    85: op1_00_inv11 = 1;
    90: op1_00_inv11 = 1;
    92: op1_00_inv11 = 1;
    default: op1_00_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in12 = reg_0451;
    14: op1_00_in12 = reg_0451;
    59: op1_00_in12 = reg_0451;
    5: op1_00_in12 = reg_0041;
    6: op1_00_in12 = reg_0193;
    75: op1_00_in12 = reg_0193;
    7: op1_00_in12 = reg_0292;
    8: op1_00_in12 = reg_0442;
    9: op1_00_in12 = reg_0101;
    10: op1_00_in12 = reg_0115;
    11: op1_00_in12 = reg_0409;
    12: op1_00_in12 = reg_0200;
    13: op1_00_in12 = reg_0274;
    15: op1_00_in12 = reg_0213;
    16: op1_00_in12 = reg_0007;
    17: op1_00_in12 = reg_0146;
    18: op1_00_in12 = reg_0783;
    19: op1_00_in12 = reg_0622;
    20: op1_00_in12 = reg_0391;
    21: op1_00_in12 = reg_0035;
    22: op1_00_in12 = reg_0202;
    23: op1_00_in12 = imem05_in[95:92];
    24: op1_00_in12 = imem02_in[7:4];
    25: op1_00_in12 = reg_0572;
    26: op1_00_in12 = reg_0468;
    27: op1_00_in12 = imem04_in[107:104];
    28: op1_00_in12 = imem07_in[35:32];
    29: op1_00_in12 = reg_0204;
    30: op1_00_in12 = imem04_in[3:0];
    31: op1_00_in12 = reg_0432;
    32: op1_00_in12 = reg_0474;
    33: op1_00_in12 = imem01_in[39:36];
    34: op1_00_in12 = reg_0817;
    35: op1_00_in12 = reg_0778;
    36: op1_00_in12 = reg_0434;
    37: op1_00_in12 = reg_0214;
    38: op1_00_in12 = reg_0473;
    39: op1_00_in12 = reg_0665;
    40: op1_00_in12 = imem02_in[47:44];
    41: op1_00_in12 = reg_0781;
    43: op1_00_in12 = reg_0475;
    44: op1_00_in12 = reg_0498;
    45: op1_00_in12 = reg_0787;
    46: op1_00_in12 = reg_0680;
    47: op1_00_in12 = reg_0114;
    48: op1_00_in12 = reg_0482;
    49: op1_00_in12 = reg_0278;
    50: op1_00_in12 = reg_0515;
    51: op1_00_in12 = reg_0531;
    52: op1_00_in12 = imem03_in[7:4];
    53: op1_00_in12 = reg_0014;
    54: op1_00_in12 = reg_0015;
    55: op1_00_in12 = imem06_in[63:60];
    56: op1_00_in12 = reg_0176;
    57: op1_00_in12 = imem07_in[103:100];
    58: op1_00_in12 = reg_0256;
    60: op1_00_in12 = reg_0726;
    61: op1_00_in12 = reg_0188;
    62: op1_00_in12 = imem03_in[87:84];
    63: op1_00_in12 = reg_0416;
    64: op1_00_in12 = reg_0156;
    65: op1_00_in12 = imem06_in[31:28];
    66: op1_00_in12 = reg_0370;
    67: op1_00_in12 = reg_0136;
    68: op1_00_in12 = imem02_in[59:56];
    69: op1_00_in12 = imem04_in[63:60];
    70: op1_00_in12 = reg_0051;
    71: op1_00_in12 = reg_0347;
    72: op1_00_in12 = imem06_in[11:8];
    73: op1_00_in12 = reg_0608;
    76: op1_00_in12 = reg_0461;
    77: op1_00_in12 = reg_0755;
    78: op1_00_in12 = imem06_in[119:116];
    79: op1_00_in12 = reg_0139;
    82: op1_00_in12 = reg_0644;
    83: op1_00_in12 = imem03_in[39:36];
    84: op1_00_in12 = reg_0799;
    85: op1_00_in12 = imem07_in[67:64];
    86: op1_00_in12 = imem06_in[107:104];
    87: op1_00_in12 = imem04_in[51:48];
    88: op1_00_in12 = reg_0166;
    89: op1_00_in12 = reg_0331;
    90: op1_00_in12 = imem06_in[99:96];
    91: op1_00_in12 = reg_0633;
    92: op1_00_in12 = reg_0042;
    93: op1_00_in12 = reg_0106;
    94: op1_00_in12 = imem02_in[71:68];
    95: op1_00_in12 = reg_0472;
    96: op1_00_in12 = reg_0477;
    default: op1_00_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv12 = 1;
    7: op1_00_inv12 = 1;
    8: op1_00_inv12 = 1;
    9: op1_00_inv12 = 1;
    10: op1_00_inv12 = 1;
    11: op1_00_inv12 = 1;
    12: op1_00_inv12 = 1;
    14: op1_00_inv12 = 1;
    15: op1_00_inv12 = 1;
    16: op1_00_inv12 = 1;
    17: op1_00_inv12 = 1;
    18: op1_00_inv12 = 1;
    19: op1_00_inv12 = 1;
    21: op1_00_inv12 = 1;
    22: op1_00_inv12 = 1;
    23: op1_00_inv12 = 1;
    24: op1_00_inv12 = 1;
    26: op1_00_inv12 = 1;
    27: op1_00_inv12 = 1;
    30: op1_00_inv12 = 1;
    31: op1_00_inv12 = 1;
    33: op1_00_inv12 = 1;
    36: op1_00_inv12 = 1;
    37: op1_00_inv12 = 1;
    39: op1_00_inv12 = 1;
    43: op1_00_inv12 = 1;
    45: op1_00_inv12 = 1;
    48: op1_00_inv12 = 1;
    50: op1_00_inv12 = 1;
    52: op1_00_inv12 = 1;
    54: op1_00_inv12 = 1;
    55: op1_00_inv12 = 1;
    59: op1_00_inv12 = 1;
    60: op1_00_inv12 = 1;
    61: op1_00_inv12 = 1;
    63: op1_00_inv12 = 1;
    66: op1_00_inv12 = 1;
    67: op1_00_inv12 = 1;
    69: op1_00_inv12 = 1;
    70: op1_00_inv12 = 1;
    72: op1_00_inv12 = 1;
    75: op1_00_inv12 = 1;
    77: op1_00_inv12 = 1;
    78: op1_00_inv12 = 1;
    85: op1_00_inv12 = 1;
    86: op1_00_inv12 = 1;
    87: op1_00_inv12 = 1;
    88: op1_00_inv12 = 1;
    89: op1_00_inv12 = 1;
    90: op1_00_inv12 = 1;
    92: op1_00_inv12 = 1;
    93: op1_00_inv12 = 1;
    94: op1_00_inv12 = 1;
    95: op1_00_inv12 = 1;
    96: op1_00_inv12 = 1;
    default: op1_00_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in13 = reg_0455;
    5: op1_00_in13 = reg_0065;
    6: op1_00_in13 = reg_0195;
    7: op1_00_in13 = reg_0295;
    8: op1_00_in13 = reg_0443;
    9: op1_00_in13 = reg_0109;
    10: op1_00_in13 = reg_0110;
    11: op1_00_in13 = reg_0337;
    12: op1_00_in13 = reg_0203;
    13: op1_00_in13 = reg_0260;
    14: op1_00_in13 = reg_0466;
    15: op1_00_in13 = reg_0205;
    16: op1_00_in13 = reg_0008;
    17: op1_00_in13 = reg_0143;
    64: op1_00_in13 = reg_0143;
    18: op1_00_in13 = reg_0271;
    19: op1_00_in13 = reg_0348;
    20: op1_00_in13 = reg_0321;
    21: op1_00_in13 = reg_0036;
    22: op1_00_in13 = reg_0199;
    23: op1_00_in13 = imem05_in[103:100];
    24: op1_00_in13 = imem02_in[23:20];
    25: op1_00_in13 = reg_0576;
    26: op1_00_in13 = reg_0459;
    27: op1_00_in13 = reg_0315;
    28: op1_00_in13 = imem07_in[39:36];
    29: op1_00_in13 = reg_0207;
    30: op1_00_in13 = imem04_in[63:60];
    31: op1_00_in13 = reg_0422;
    32: op1_00_in13 = reg_0456;
    33: op1_00_in13 = imem01_in[87:84];
    34: op1_00_in13 = reg_0606;
    35: op1_00_in13 = reg_0817;
    78: op1_00_in13 = reg_0817;
    36: op1_00_in13 = reg_0446;
    37: op1_00_in13 = reg_0210;
    38: op1_00_in13 = reg_0470;
    39: op1_00_in13 = reg_0229;
    40: op1_00_in13 = imem02_in[71:68];
    41: op1_00_in13 = reg_0491;
    48: op1_00_in13 = reg_0491;
    43: op1_00_in13 = reg_0481;
    44: op1_00_in13 = reg_0094;
    45: op1_00_in13 = reg_0091;
    46: op1_00_in13 = reg_0673;
    47: op1_00_in13 = reg_0113;
    49: op1_00_in13 = reg_0774;
    50: op1_00_in13 = reg_0288;
    51: op1_00_in13 = reg_0526;
    52: op1_00_in13 = imem03_in[15:12];
    53: op1_00_in13 = imem04_in[7:4];
    54: op1_00_in13 = imem04_in[27:24];
    55: op1_00_in13 = imem06_in[71:68];
    56: op1_00_in13 = reg_0171;
    57: op1_00_in13 = reg_0728;
    58: op1_00_in13 = reg_0148;
    59: op1_00_in13 = reg_0457;
    60: op1_00_in13 = reg_0717;
    61: op1_00_in13 = reg_0201;
    62: op1_00_in13 = imem03_in[123:120];
    63: op1_00_in13 = imem05_in[19:16];
    65: op1_00_in13 = imem06_in[67:64];
    66: op1_00_in13 = reg_0609;
    67: op1_00_in13 = reg_0141;
    68: op1_00_in13 = imem02_in[75:72];
    69: op1_00_in13 = imem04_in[75:72];
    70: op1_00_in13 = reg_0333;
    71: op1_00_in13 = reg_0750;
    72: op1_00_in13 = imem06_in[19:16];
    73: op1_00_in13 = reg_0638;
    75: op1_00_in13 = reg_0186;
    76: op1_00_in13 = reg_0475;
    77: op1_00_in13 = reg_0568;
    79: op1_00_in13 = reg_0307;
    82: op1_00_in13 = imem05_in[11:8];
    83: op1_00_in13 = imem03_in[51:48];
    84: op1_00_in13 = reg_0016;
    85: op1_00_in13 = imem07_in[87:84];
    86: op1_00_in13 = imem06_in[127:124];
    87: op1_00_in13 = reg_0247;
    88: op1_00_in13 = reg_0712;
    89: op1_00_in13 = reg_0615;
    90: op1_00_in13 = imem06_in[103:100];
    91: op1_00_in13 = imem07_in[3:0];
    92: op1_00_in13 = reg_0392;
    93: op1_00_in13 = reg_0126;
    94: op1_00_in13 = imem02_in[91:88];
    95: op1_00_in13 = reg_0480;
    96: op1_00_in13 = reg_0476;
    default: op1_00_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv13 = 1;
    5: op1_00_inv13 = 1;
    7: op1_00_inv13 = 1;
    8: op1_00_inv13 = 1;
    14: op1_00_inv13 = 1;
    15: op1_00_inv13 = 1;
    16: op1_00_inv13 = 1;
    17: op1_00_inv13 = 1;
    18: op1_00_inv13 = 1;
    19: op1_00_inv13 = 1;
    22: op1_00_inv13 = 1;
    24: op1_00_inv13 = 1;
    25: op1_00_inv13 = 1;
    27: op1_00_inv13 = 1;
    31: op1_00_inv13 = 1;
    32: op1_00_inv13 = 1;
    34: op1_00_inv13 = 1;
    37: op1_00_inv13 = 1;
    38: op1_00_inv13 = 1;
    43: op1_00_inv13 = 1;
    47: op1_00_inv13 = 1;
    48: op1_00_inv13 = 1;
    49: op1_00_inv13 = 1;
    51: op1_00_inv13 = 1;
    52: op1_00_inv13 = 1;
    54: op1_00_inv13 = 1;
    57: op1_00_inv13 = 1;
    58: op1_00_inv13 = 1;
    59: op1_00_inv13 = 1;
    66: op1_00_inv13 = 1;
    68: op1_00_inv13 = 1;
    70: op1_00_inv13 = 1;
    71: op1_00_inv13 = 1;
    73: op1_00_inv13 = 1;
    79: op1_00_inv13 = 1;
    82: op1_00_inv13 = 1;
    84: op1_00_inv13 = 1;
    85: op1_00_inv13 = 1;
    87: op1_00_inv13 = 1;
    90: op1_00_inv13 = 1;
    94: op1_00_inv13 = 1;
    95: op1_00_inv13 = 1;
    default: op1_00_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in14 = reg_0466;
    5: op1_00_in14 = imem05_in[19:16];
    6: op1_00_in14 = imem01_in[3:0];
    7: op1_00_in14 = reg_0065;
    8: op1_00_in14 = reg_0165;
    9: op1_00_in14 = reg_0117;
    10: op1_00_in14 = imem02_in[47:44];
    93: op1_00_in14 = imem02_in[47:44];
    11: op1_00_in14 = reg_0813;
    12: op1_00_in14 = reg_0194;
    13: op1_00_in14 = reg_0145;
    14: op1_00_in14 = reg_0460;
    15: op1_00_in14 = imem01_in[27:24];
    16: op1_00_in14 = imem04_in[47:44];
    54: op1_00_in14 = imem04_in[47:44];
    17: op1_00_in14 = reg_0138;
    18: op1_00_in14 = reg_0737;
    19: op1_00_in14 = reg_0356;
    20: op1_00_in14 = reg_0369;
    21: op1_00_in14 = reg_0029;
    22: op1_00_in14 = imem01_in[19:16];
    23: op1_00_in14 = imem05_in[119:116];
    24: op1_00_in14 = imem02_in[59:56];
    25: op1_00_in14 = reg_0385;
    26: op1_00_in14 = reg_0452;
    27: op1_00_in14 = reg_0056;
    28: op1_00_in14 = imem07_in[59:56];
    29: op1_00_in14 = reg_0196;
    30: op1_00_in14 = imem04_in[67:64];
    31: op1_00_in14 = reg_0419;
    32: op1_00_in14 = reg_0200;
    33: op1_00_in14 = imem01_in[91:88];
    34: op1_00_in14 = imem07_in[7:4];
    91: op1_00_in14 = imem07_in[7:4];
    35: op1_00_in14 = reg_0375;
    36: op1_00_in14 = reg_0444;
    37: op1_00_in14 = reg_0209;
    38: op1_00_in14 = reg_0468;
    76: op1_00_in14 = reg_0468;
    39: op1_00_in14 = reg_0363;
    40: op1_00_in14 = imem02_in[79:76];
    41: op1_00_in14 = reg_0780;
    43: op1_00_in14 = reg_0480;
    44: op1_00_in14 = imem03_in[27:24];
    45: op1_00_in14 = reg_0304;
    46: op1_00_in14 = reg_0450;
    47: op1_00_in14 = imem02_in[3:0];
    48: op1_00_in14 = reg_0492;
    49: op1_00_in14 = reg_0317;
    50: op1_00_in14 = imem05_in[47:44];
    51: op1_00_in14 = reg_0094;
    52: op1_00_in14 = imem03_in[51:48];
    53: op1_00_in14 = imem04_in[31:28];
    55: op1_00_in14 = imem06_in[83:80];
    65: op1_00_in14 = imem06_in[83:80];
    56: op1_00_in14 = reg_0184;
    57: op1_00_in14 = reg_0064;
    58: op1_00_in14 = reg_0154;
    59: op1_00_in14 = reg_0469;
    60: op1_00_in14 = reg_0705;
    61: op1_00_in14 = reg_0212;
    62: op1_00_in14 = reg_0281;
    63: op1_00_in14 = imem05_in[71:68];
    64: op1_00_in14 = imem06_in[35:32];
    66: op1_00_in14 = reg_0298;
    67: op1_00_in14 = reg_0144;
    68: op1_00_in14 = imem02_in[111:108];
    69: op1_00_in14 = imem04_in[123:120];
    70: op1_00_in14 = reg_0084;
    71: op1_00_in14 = reg_0350;
    72: op1_00_in14 = imem06_in[47:44];
    73: op1_00_in14 = reg_0764;
    75: op1_00_in14 = reg_0198;
    77: op1_00_in14 = reg_0572;
    78: op1_00_in14 = reg_0260;
    79: op1_00_in14 = reg_0149;
    82: op1_00_in14 = imem05_in[43:40];
    83: op1_00_in14 = imem03_in[55:52];
    84: op1_00_in14 = reg_0810;
    85: op1_00_in14 = imem07_in[99:96];
    86: op1_00_in14 = reg_0289;
    87: op1_00_in14 = reg_0553;
    88: op1_00_in14 = reg_0158;
    89: op1_00_in14 = reg_0077;
    90: op1_00_in14 = reg_0348;
    92: op1_00_in14 = reg_0358;
    94: op1_00_in14 = imem02_in[119:116];
    95: op1_00_in14 = imem01_in[39:36];
    96: op1_00_in14 = reg_0475;
    default: op1_00_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv14 = 1;
    7: op1_00_inv14 = 1;
    8: op1_00_inv14 = 1;
    9: op1_00_inv14 = 1;
    10: op1_00_inv14 = 1;
    12: op1_00_inv14 = 1;
    14: op1_00_inv14 = 1;
    17: op1_00_inv14 = 1;
    18: op1_00_inv14 = 1;
    19: op1_00_inv14 = 1;
    21: op1_00_inv14 = 1;
    22: op1_00_inv14 = 1;
    23: op1_00_inv14 = 1;
    26: op1_00_inv14 = 1;
    27: op1_00_inv14 = 1;
    32: op1_00_inv14 = 1;
    33: op1_00_inv14 = 1;
    36: op1_00_inv14 = 1;
    37: op1_00_inv14 = 1;
    38: op1_00_inv14 = 1;
    39: op1_00_inv14 = 1;
    43: op1_00_inv14 = 1;
    44: op1_00_inv14 = 1;
    48: op1_00_inv14 = 1;
    49: op1_00_inv14 = 1;
    53: op1_00_inv14 = 1;
    54: op1_00_inv14 = 1;
    55: op1_00_inv14 = 1;
    57: op1_00_inv14 = 1;
    61: op1_00_inv14 = 1;
    67: op1_00_inv14 = 1;
    69: op1_00_inv14 = 1;
    72: op1_00_inv14 = 1;
    73: op1_00_inv14 = 1;
    77: op1_00_inv14 = 1;
    83: op1_00_inv14 = 1;
    85: op1_00_inv14 = 1;
    87: op1_00_inv14 = 1;
    88: op1_00_inv14 = 1;
    89: op1_00_inv14 = 1;
    92: op1_00_inv14 = 1;
    93: op1_00_inv14 = 1;
    94: op1_00_inv14 = 1;
    95: op1_00_inv14 = 1;
    default: op1_00_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in15 = reg_0473;
    5: op1_00_in15 = imem05_in[35:32];
    6: op1_00_in15 = imem01_in[51:48];
    7: op1_00_in15 = reg_0053;
    57: op1_00_in15 = reg_0053;
    9: op1_00_in15 = imem02_in[3:0];
    10: op1_00_in15 = imem02_in[51:48];
    11: op1_00_in15 = reg_0815;
    12: op1_00_in15 = reg_0206;
    13: op1_00_in15 = reg_0133;
    14: op1_00_in15 = reg_0209;
    15: op1_00_in15 = imem01_in[127:124];
    16: op1_00_in15 = imem04_in[99:96];
    17: op1_00_in15 = imem06_in[19:16];
    67: op1_00_in15 = imem06_in[19:16];
    18: op1_00_in15 = reg_0735;
    19: op1_00_in15 = reg_0383;
    20: op1_00_in15 = reg_0808;
    21: op1_00_in15 = imem07_in[15:12];
    22: op1_00_in15 = imem01_in[23:20];
    23: op1_00_in15 = reg_0789;
    24: op1_00_in15 = imem02_in[67:64];
    93: op1_00_in15 = imem02_in[67:64];
    25: op1_00_in15 = reg_0374;
    26: op1_00_in15 = reg_0456;
    27: op1_00_in15 = reg_0060;
    28: op1_00_in15 = imem07_in[63:60];
    29: op1_00_in15 = reg_0202;
    30: op1_00_in15 = reg_0059;
    69: op1_00_in15 = reg_0059;
    31: op1_00_in15 = reg_0431;
    32: op1_00_in15 = reg_0211;
    33: op1_00_in15 = imem01_in[103:100];
    34: op1_00_in15 = imem07_in[59:56];
    35: op1_00_in15 = reg_0779;
    36: op1_00_in15 = reg_0437;
    37: op1_00_in15 = reg_0188;
    38: op1_00_in15 = reg_0459;
    43: op1_00_in15 = reg_0459;
    39: op1_00_in15 = reg_0322;
    40: op1_00_in15 = reg_0666;
    41: op1_00_in15 = reg_0495;
    44: op1_00_in15 = imem03_in[39:36];
    45: op1_00_in15 = reg_0275;
    46: op1_00_in15 = reg_0469;
    47: op1_00_in15 = imem02_in[15:12];
    48: op1_00_in15 = reg_0494;
    49: op1_00_in15 = reg_0577;
    50: op1_00_in15 = imem05_in[103:100];
    51: op1_00_in15 = imem03_in[7:4];
    52: op1_00_in15 = imem03_in[95:92];
    53: op1_00_in15 = imem04_in[47:44];
    54: op1_00_in15 = imem04_in[59:56];
    55: op1_00_in15 = imem06_in[115:112];
    58: op1_00_in15 = reg_0139;
    59: op1_00_in15 = reg_0467;
    60: op1_00_in15 = reg_0713;
    61: op1_00_in15 = imem01_in[71:68];
    62: op1_00_in15 = reg_0572;
    63: op1_00_in15 = imem05_in[91:88];
    64: op1_00_in15 = imem06_in[47:44];
    65: op1_00_in15 = imem06_in[91:88];
    66: op1_00_in15 = reg_0606;
    68: op1_00_in15 = reg_0089;
    70: op1_00_in15 = reg_0438;
    71: op1_00_in15 = reg_0329;
    72: op1_00_in15 = reg_0605;
    73: op1_00_in15 = reg_0573;
    75: op1_00_in15 = reg_0196;
    76: op1_00_in15 = reg_0191;
    77: op1_00_in15 = reg_0637;
    78: op1_00_in15 = reg_0402;
    79: op1_00_in15 = reg_0765;
    82: op1_00_in15 = imem05_in[55:52];
    83: op1_00_in15 = imem03_in[63:60];
    84: op1_00_in15 = reg_0010;
    85: op1_00_in15 = imem07_in[115:112];
    86: op1_00_in15 = reg_0348;
    87: op1_00_in15 = reg_0551;
    88: op1_00_in15 = reg_0253;
    89: op1_00_in15 = reg_0616;
    90: op1_00_in15 = reg_0346;
    91: op1_00_in15 = imem07_in[55:52];
    92: op1_00_in15 = reg_0345;
    94: op1_00_in15 = reg_0642;
    95: op1_00_in15 = imem01_in[67:64];
    96: op1_00_in15 = reg_0480;
    default: op1_00_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv15 = 1;
    5: op1_00_inv15 = 1;
    11: op1_00_inv15 = 1;
    15: op1_00_inv15 = 1;
    17: op1_00_inv15 = 1;
    18: op1_00_inv15 = 1;
    20: op1_00_inv15 = 1;
    23: op1_00_inv15 = 1;
    26: op1_00_inv15 = 1;
    28: op1_00_inv15 = 1;
    29: op1_00_inv15 = 1;
    30: op1_00_inv15 = 1;
    33: op1_00_inv15 = 1;
    34: op1_00_inv15 = 1;
    40: op1_00_inv15 = 1;
    41: op1_00_inv15 = 1;
    44: op1_00_inv15 = 1;
    45: op1_00_inv15 = 1;
    47: op1_00_inv15 = 1;
    51: op1_00_inv15 = 1;
    53: op1_00_inv15 = 1;
    54: op1_00_inv15 = 1;
    55: op1_00_inv15 = 1;
    57: op1_00_inv15 = 1;
    58: op1_00_inv15 = 1;
    59: op1_00_inv15 = 1;
    60: op1_00_inv15 = 1;
    62: op1_00_inv15 = 1;
    64: op1_00_inv15 = 1;
    65: op1_00_inv15 = 1;
    66: op1_00_inv15 = 1;
    67: op1_00_inv15 = 1;
    68: op1_00_inv15 = 1;
    72: op1_00_inv15 = 1;
    73: op1_00_inv15 = 1;
    76: op1_00_inv15 = 1;
    83: op1_00_inv15 = 1;
    84: op1_00_inv15 = 1;
    85: op1_00_inv15 = 1;
    87: op1_00_inv15 = 1;
    89: op1_00_inv15 = 1;
    91: op1_00_inv15 = 1;
    92: op1_00_inv15 = 1;
    93: op1_00_inv15 = 1;
    94: op1_00_inv15 = 1;
    96: op1_00_inv15 = 1;
    default: op1_00_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in16 = reg_0467;
    5: op1_00_in16 = imem05_in[79:76];
    6: op1_00_in16 = imem01_in[123:120];
    7: op1_00_in16 = reg_0068;
    9: op1_00_in16 = imem02_in[19:16];
    10: op1_00_in16 = imem02_in[91:88];
    11: op1_00_in16 = reg_0040;
    12: op1_00_in16 = imem01_in[39:36];
    13: op1_00_in16 = reg_0139;
    14: op1_00_in16 = reg_0203;
    15: op1_00_in16 = reg_0497;
    16: op1_00_in16 = reg_0544;
    17: op1_00_in16 = imem06_in[27:24];
    18: op1_00_in16 = reg_0260;
    19: op1_00_in16 = reg_0032;
    20: op1_00_in16 = reg_0810;
    21: op1_00_in16 = imem07_in[19:16];
    22: op1_00_in16 = imem01_in[47:44];
    23: op1_00_in16 = reg_0494;
    24: op1_00_in16 = imem02_in[75:72];
    93: op1_00_in16 = imem02_in[75:72];
    25: op1_00_in16 = reg_0389;
    26: op1_00_in16 = reg_0214;
    27: op1_00_in16 = reg_0554;
    28: op1_00_in16 = imem07_in[127:124];
    29: op1_00_in16 = imem01_in[19:16];
    30: op1_00_in16 = reg_0087;
    31: op1_00_in16 = reg_0159;
    32: op1_00_in16 = reg_0198;
    33: op1_00_in16 = reg_0501;
    34: op1_00_in16 = imem07_in[67:64];
    35: op1_00_in16 = imem07_in[11:8];
    36: op1_00_in16 = reg_0420;
    37: op1_00_in16 = imem01_in[59:56];
    38: op1_00_in16 = reg_0478;
    39: op1_00_in16 = reg_0518;
    40: op1_00_in16 = reg_0655;
    41: op1_00_in16 = reg_0794;
    43: op1_00_in16 = reg_0191;
    44: op1_00_in16 = imem03_in[51:48];
    45: op1_00_in16 = reg_0224;
    46: op1_00_in16 = reg_0481;
    47: op1_00_in16 = imem02_in[43:40];
    48: op1_00_in16 = reg_0495;
    49: op1_00_in16 = reg_0405;
    50: op1_00_in16 = reg_0791;
    51: op1_00_in16 = imem03_in[27:24];
    52: op1_00_in16 = imem03_in[99:96];
    53: op1_00_in16 = imem04_in[91:88];
    84: op1_00_in16 = imem04_in[91:88];
    54: op1_00_in16 = imem04_in[63:60];
    55: op1_00_in16 = imem06_in[119:116];
    57: op1_00_in16 = reg_0447;
    58: op1_00_in16 = imem06_in[19:16];
    59: op1_00_in16 = reg_0468;
    60: op1_00_in16 = reg_0715;
    61: op1_00_in16 = reg_0646;
    62: op1_00_in16 = reg_0393;
    63: op1_00_in16 = imem05_in[99:96];
    64: op1_00_in16 = imem06_in[87:84];
    65: op1_00_in16 = imem06_in[107:104];
    66: op1_00_in16 = reg_0238;
    67: op1_00_in16 = imem06_in[31:28];
    68: op1_00_in16 = reg_0739;
    69: op1_00_in16 = reg_0262;
    70: op1_00_in16 = reg_0268;
    71: op1_00_in16 = reg_0357;
    72: op1_00_in16 = reg_0038;
    73: op1_00_in16 = reg_0777;
    75: op1_00_in16 = reg_0202;
    76: op1_00_in16 = reg_0209;
    77: op1_00_in16 = reg_0557;
    78: op1_00_in16 = reg_0628;
    79: op1_00_in16 = reg_0137;
    82: op1_00_in16 = imem05_in[59:56];
    83: op1_00_in16 = imem03_in[75:72];
    85: op1_00_in16 = reg_0391;
    86: op1_00_in16 = reg_0625;
    87: op1_00_in16 = reg_0303;
    88: op1_00_in16 = reg_0333;
    89: op1_00_in16 = reg_0679;
    90: op1_00_in16 = reg_0762;
    91: op1_00_in16 = imem07_in[91:88];
    92: op1_00_in16 = reg_0414;
    94: op1_00_in16 = reg_0088;
    95: op1_00_in16 = imem01_in[71:68];
    96: op1_00_in16 = reg_0479;
    default: op1_00_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv16 = 1;
    7: op1_00_inv16 = 1;
    10: op1_00_inv16 = 1;
    11: op1_00_inv16 = 1;
    14: op1_00_inv16 = 1;
    16: op1_00_inv16 = 1;
    18: op1_00_inv16 = 1;
    20: op1_00_inv16 = 1;
    23: op1_00_inv16 = 1;
    26: op1_00_inv16 = 1;
    28: op1_00_inv16 = 1;
    29: op1_00_inv16 = 1;
    30: op1_00_inv16 = 1;
    31: op1_00_inv16 = 1;
    32: op1_00_inv16 = 1;
    34: op1_00_inv16 = 1;
    38: op1_00_inv16 = 1;
    40: op1_00_inv16 = 1;
    44: op1_00_inv16 = 1;
    49: op1_00_inv16 = 1;
    52: op1_00_inv16 = 1;
    54: op1_00_inv16 = 1;
    55: op1_00_inv16 = 1;
    57: op1_00_inv16 = 1;
    59: op1_00_inv16 = 1;
    62: op1_00_inv16 = 1;
    63: op1_00_inv16 = 1;
    64: op1_00_inv16 = 1;
    65: op1_00_inv16 = 1;
    66: op1_00_inv16 = 1;
    69: op1_00_inv16 = 1;
    70: op1_00_inv16 = 1;
    71: op1_00_inv16 = 1;
    72: op1_00_inv16 = 1;
    73: op1_00_inv16 = 1;
    75: op1_00_inv16 = 1;
    77: op1_00_inv16 = 1;
    83: op1_00_inv16 = 1;
    84: op1_00_inv16 = 1;
    85: op1_00_inv16 = 1;
    86: op1_00_inv16 = 1;
    88: op1_00_inv16 = 1;
    89: op1_00_inv16 = 1;
    90: op1_00_inv16 = 1;
    91: op1_00_inv16 = 1;
    93: op1_00_inv16 = 1;
    96: op1_00_inv16 = 1;
    default: op1_00_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in17 = reg_0474;
    5: op1_00_in17 = imem05_in[115:112];
    6: op1_00_in17 = reg_0501;
    7: op1_00_in17 = reg_0074;
    9: op1_00_in17 = imem02_in[27:24];
    10: op1_00_in17 = reg_0658;
    11: op1_00_in17 = reg_0819;
    12: op1_00_in17 = imem01_in[59:56];
    13: op1_00_in17 = reg_0140;
    14: op1_00_in17 = reg_0193;
    15: op1_00_in17 = reg_0509;
    16: op1_00_in17 = reg_0553;
    17: op1_00_in17 = imem06_in[35:32];
    18: op1_00_in17 = reg_0269;
    19: op1_00_in17 = reg_0035;
    20: op1_00_in17 = reg_0004;
    21: op1_00_in17 = imem07_in[27:24];
    22: op1_00_in17 = imem01_in[63:60];
    23: op1_00_in17 = reg_0785;
    24: op1_00_in17 = reg_0666;
    25: op1_00_in17 = reg_0003;
    26: op1_00_in17 = reg_0194;
    27: op1_00_in17 = reg_0558;
    28: op1_00_in17 = reg_0728;
    91: op1_00_in17 = reg_0728;
    29: op1_00_in17 = imem01_in[31:28];
    30: op1_00_in17 = reg_0542;
    31: op1_00_in17 = reg_0173;
    32: op1_00_in17 = reg_0190;
    33: op1_00_in17 = reg_0824;
    34: op1_00_in17 = imem07_in[87:84];
    35: op1_00_in17 = imem07_in[15:12];
    36: op1_00_in17 = reg_0162;
    37: op1_00_in17 = reg_0520;
    38: op1_00_in17 = reg_0189;
    39: op1_00_in17 = reg_0541;
    40: op1_00_in17 = reg_0653;
    41: op1_00_in17 = reg_0784;
    43: op1_00_in17 = reg_0206;
    44: op1_00_in17 = imem03_in[63:60];
    45: op1_00_in17 = reg_0138;
    46: op1_00_in17 = reg_0468;
    47: op1_00_in17 = imem02_in[51:48];
    48: op1_00_in17 = reg_0742;
    49: op1_00_in17 = reg_0748;
    50: op1_00_in17 = reg_0798;
    51: op1_00_in17 = imem03_in[59:56];
    52: op1_00_in17 = reg_0599;
    53: op1_00_in17 = reg_0544;
    84: op1_00_in17 = reg_0544;
    54: op1_00_in17 = reg_0088;
    55: op1_00_in17 = reg_0628;
    57: op1_00_in17 = reg_0160;
    58: op1_00_in17 = imem06_in[27:24];
    59: op1_00_in17 = reg_0458;
    60: op1_00_in17 = reg_0718;
    61: op1_00_in17 = reg_0741;
    62: op1_00_in17 = reg_0001;
    63: op1_00_in17 = reg_0796;
    64: op1_00_in17 = imem06_in[103:100];
    65: op1_00_in17 = imem06_in[119:116];
    66: op1_00_in17 = reg_0618;
    67: op1_00_in17 = imem06_in[43:40];
    68: op1_00_in17 = reg_0637;
    69: op1_00_in17 = reg_0560;
    70: op1_00_in17 = reg_0164;
    71: op1_00_in17 = reg_0331;
    72: op1_00_in17 = reg_0401;
    73: op1_00_in17 = reg_0661;
    75: op1_00_in17 = reg_0199;
    76: op1_00_in17 = reg_0201;
    77: op1_00_in17 = reg_0006;
    78: op1_00_in17 = reg_0659;
    79: op1_00_in17 = imem06_in[19:16];
    82: op1_00_in17 = imem05_in[71:68];
    83: op1_00_in17 = imem03_in[91:88];
    85: op1_00_in17 = reg_0161;
    86: op1_00_in17 = reg_0115;
    87: op1_00_in17 = reg_0429;
    88: op1_00_in17 = reg_0434;
    89: op1_00_in17 = reg_0776;
    90: op1_00_in17 = reg_0298;
    92: op1_00_in17 = reg_0132;
    93: op1_00_in17 = imem02_in[79:76];
    94: op1_00_in17 = reg_0533;
    95: op1_00_in17 = imem01_in[103:100];
    96: op1_00_in17 = reg_0214;
    default: op1_00_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv17 = 1;
    9: op1_00_inv17 = 1;
    13: op1_00_inv17 = 1;
    16: op1_00_inv17 = 1;
    19: op1_00_inv17 = 1;
    20: op1_00_inv17 = 1;
    27: op1_00_inv17 = 1;
    29: op1_00_inv17 = 1;
    30: op1_00_inv17 = 1;
    31: op1_00_inv17 = 1;
    35: op1_00_inv17 = 1;
    36: op1_00_inv17 = 1;
    38: op1_00_inv17 = 1;
    39: op1_00_inv17 = 1;
    43: op1_00_inv17 = 1;
    48: op1_00_inv17 = 1;
    49: op1_00_inv17 = 1;
    58: op1_00_inv17 = 1;
    59: op1_00_inv17 = 1;
    66: op1_00_inv17 = 1;
    68: op1_00_inv17 = 1;
    69: op1_00_inv17 = 1;
    71: op1_00_inv17 = 1;
    75: op1_00_inv17 = 1;
    76: op1_00_inv17 = 1;
    79: op1_00_inv17 = 1;
    83: op1_00_inv17 = 1;
    84: op1_00_inv17 = 1;
    86: op1_00_inv17 = 1;
    88: op1_00_inv17 = 1;
    89: op1_00_inv17 = 1;
    90: op1_00_inv17 = 1;
    95: op1_00_inv17 = 1;
    96: op1_00_inv17 = 1;
    default: op1_00_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in18 = reg_0452;
    5: op1_00_in18 = imem05_in[127:124];
    6: op1_00_in18 = reg_0522;
    7: op1_00_in18 = reg_0064;
    9: op1_00_in18 = imem02_in[39:36];
    10: op1_00_in18 = reg_0653;
    11: op1_00_in18 = imem07_in[7:4];
    12: op1_00_in18 = imem01_in[75:72];
    13: op1_00_in18 = imem06_in[11:8];
    14: op1_00_in18 = reg_0205;
    15: op1_00_in18 = reg_0514;
    16: op1_00_in18 = reg_0552;
    17: op1_00_in18 = imem06_in[39:36];
    18: op1_00_in18 = reg_0145;
    19: op1_00_in18 = reg_0748;
    20: op1_00_in18 = imem04_in[59:56];
    21: op1_00_in18 = imem07_in[39:36];
    22: op1_00_in18 = imem01_in[79:76];
    23: op1_00_in18 = reg_0495;
    24: op1_00_in18 = reg_0667;
    25: op1_00_in18 = reg_0016;
    62: op1_00_in18 = reg_0016;
    26: op1_00_in18 = reg_0201;
    27: op1_00_in18 = reg_0516;
    28: op1_00_in18 = reg_0731;
    29: op1_00_in18 = imem01_in[35:32];
    30: op1_00_in18 = reg_0060;
    32: op1_00_in18 = imem01_in[51:48];
    33: op1_00_in18 = reg_0227;
    34: op1_00_in18 = reg_0710;
    35: op1_00_in18 = imem07_in[19:16];
    36: op1_00_in18 = reg_0167;
    37: op1_00_in18 = reg_0515;
    38: op1_00_in18 = reg_0193;
    39: op1_00_in18 = reg_0081;
    40: op1_00_in18 = reg_0656;
    41: op1_00_in18 = reg_0489;
    43: op1_00_in18 = reg_0197;
    44: op1_00_in18 = imem03_in[99:96];
    45: op1_00_in18 = reg_0153;
    46: op1_00_in18 = reg_0459;
    47: op1_00_in18 = imem02_in[67:64];
    48: op1_00_in18 = reg_0136;
    49: op1_00_in18 = reg_0404;
    50: op1_00_in18 = reg_0490;
    51: op1_00_in18 = imem03_in[107:104];
    52: op1_00_in18 = reg_0591;
    53: op1_00_in18 = reg_0055;
    54: op1_00_in18 = reg_0555;
    55: op1_00_in18 = reg_0625;
    57: op1_00_in18 = reg_0163;
    58: op1_00_in18 = imem06_in[75:72];
    59: op1_00_in18 = reg_0189;
    60: op1_00_in18 = reg_0701;
    61: op1_00_in18 = reg_0563;
    63: op1_00_in18 = reg_0278;
    64: op1_00_in18 = imem06_in[127:124];
    65: op1_00_in18 = imem06_in[127:124];
    66: op1_00_in18 = reg_0401;
    67: op1_00_in18 = imem06_in[47:44];
    68: op1_00_in18 = reg_0417;
    69: op1_00_in18 = reg_0536;
    70: op1_00_in18 = reg_0170;
    71: op1_00_in18 = reg_0648;
    72: op1_00_in18 = reg_0402;
    73: op1_00_in18 = reg_0367;
    75: op1_00_in18 = imem01_in[23:20];
    76: op1_00_in18 = reg_0190;
    77: op1_00_in18 = reg_0012;
    78: op1_00_in18 = reg_0775;
    79: op1_00_in18 = imem06_in[31:28];
    82: op1_00_in18 = imem05_in[99:96];
    83: op1_00_in18 = imem03_in[103:100];
    84: op1_00_in18 = reg_0548;
    85: op1_00_in18 = reg_0295;
    86: op1_00_in18 = reg_0349;
    87: op1_00_in18 = reg_0076;
    88: op1_00_in18 = reg_0110;
    89: op1_00_in18 = reg_0233;
    90: op1_00_in18 = reg_0618;
    91: op1_00_in18 = reg_0391;
    92: op1_00_in18 = reg_0756;
    93: op1_00_in18 = imem02_in[111:108];
    94: op1_00_in18 = reg_0080;
    95: op1_00_in18 = reg_0098;
    96: op1_00_in18 = reg_0208;
    default: op1_00_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv18 = 1;
    5: op1_00_inv18 = 1;
    7: op1_00_inv18 = 1;
    9: op1_00_inv18 = 1;
    10: op1_00_inv18 = 1;
    11: op1_00_inv18 = 1;
    13: op1_00_inv18 = 1;
    15: op1_00_inv18 = 1;
    21: op1_00_inv18 = 1;
    23: op1_00_inv18 = 1;
    24: op1_00_inv18 = 1;
    27: op1_00_inv18 = 1;
    28: op1_00_inv18 = 1;
    29: op1_00_inv18 = 1;
    30: op1_00_inv18 = 1;
    37: op1_00_inv18 = 1;
    39: op1_00_inv18 = 1;
    40: op1_00_inv18 = 1;
    41: op1_00_inv18 = 1;
    45: op1_00_inv18 = 1;
    46: op1_00_inv18 = 1;
    48: op1_00_inv18 = 1;
    54: op1_00_inv18 = 1;
    55: op1_00_inv18 = 1;
    57: op1_00_inv18 = 1;
    58: op1_00_inv18 = 1;
    60: op1_00_inv18 = 1;
    67: op1_00_inv18 = 1;
    69: op1_00_inv18 = 1;
    71: op1_00_inv18 = 1;
    72: op1_00_inv18 = 1;
    73: op1_00_inv18 = 1;
    75: op1_00_inv18 = 1;
    76: op1_00_inv18 = 1;
    78: op1_00_inv18 = 1;
    82: op1_00_inv18 = 1;
    84: op1_00_inv18 = 1;
    86: op1_00_inv18 = 1;
    87: op1_00_inv18 = 1;
    89: op1_00_inv18 = 1;
    94: op1_00_inv18 = 1;
    default: op1_00_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in19 = reg_0189;
    5: op1_00_in19 = reg_0241;
    6: op1_00_in19 = reg_0520;
    7: op1_00_in19 = imem05_in[15:12];
    9: op1_00_in19 = imem02_in[59:56];
    10: op1_00_in19 = reg_0654;
    11: op1_00_in19 = imem07_in[15:12];
    12: op1_00_in19 = reg_0500;
    27: op1_00_in19 = reg_0500;
    13: op1_00_in19 = imem06_in[15:12];
    14: op1_00_in19 = imem01_in[31:28];
    15: op1_00_in19 = reg_0776;
    16: op1_00_in19 = reg_0540;
    17: op1_00_in19 = imem06_in[119:116];
    18: op1_00_in19 = imem06_in[127:124];
    19: op1_00_in19 = reg_0751;
    20: op1_00_in19 = imem04_in[71:68];
    21: op1_00_in19 = imem07_in[43:40];
    22: op1_00_in19 = imem01_in[107:104];
    23: op1_00_in19 = reg_0226;
    24: op1_00_in19 = reg_0352;
    25: op1_00_in19 = imem04_in[23:20];
    26: op1_00_in19 = reg_0206;
    28: op1_00_in19 = reg_0721;
    34: op1_00_in19 = reg_0721;
    29: op1_00_in19 = imem01_in[83:80];
    30: op1_00_in19 = reg_0554;
    32: op1_00_in19 = imem01_in[63:60];
    33: op1_00_in19 = reg_0771;
    35: op1_00_in19 = imem07_in[67:64];
    36: op1_00_in19 = reg_0163;
    37: op1_00_in19 = reg_0235;
    38: op1_00_in19 = reg_0212;
    39: op1_00_in19 = reg_0539;
    40: op1_00_in19 = reg_0649;
    41: op1_00_in19 = reg_0736;
    43: op1_00_in19 = imem01_in[59:56];
    44: op1_00_in19 = imem03_in[103:100];
    45: op1_00_in19 = imem06_in[39:36];
    79: op1_00_in19 = imem06_in[39:36];
    46: op1_00_in19 = reg_0458;
    47: op1_00_in19 = imem02_in[83:80];
    48: op1_00_in19 = reg_0133;
    49: op1_00_in19 = reg_0406;
    50: op1_00_in19 = reg_0783;
    51: op1_00_in19 = reg_0602;
    52: op1_00_in19 = reg_0589;
    53: op1_00_in19 = reg_0060;
    54: op1_00_in19 = reg_0523;
    55: op1_00_in19 = reg_0630;
    57: op1_00_in19 = reg_0166;
    58: op1_00_in19 = imem06_in[103:100];
    59: op1_00_in19 = reg_0194;
    60: op1_00_in19 = reg_0706;
    61: op1_00_in19 = reg_0550;
    62: op1_00_in19 = reg_0010;
    63: op1_00_in19 = reg_0784;
    64: op1_00_in19 = reg_0289;
    65: op1_00_in19 = reg_0346;
    66: op1_00_in19 = reg_0031;
    67: op1_00_in19 = imem06_in[91:88];
    68: op1_00_in19 = reg_0641;
    69: op1_00_in19 = reg_0058;
    71: op1_00_in19 = reg_0403;
    72: op1_00_in19 = reg_0369;
    73: op1_00_in19 = reg_0256;
    75: op1_00_in19 = imem01_in[35:32];
    76: op1_00_in19 = reg_0199;
    77: op1_00_in19 = reg_0003;
    78: op1_00_in19 = reg_0638;
    82: op1_00_in19 = imem05_in[103:100];
    83: op1_00_in19 = reg_0063;
    84: op1_00_in19 = reg_0331;
    85: op1_00_in19 = reg_0333;
    86: op1_00_in19 = reg_0815;
    87: op1_00_in19 = reg_0292;
    88: op1_00_in19 = reg_0142;
    89: op1_00_in19 = imem05_in[47:44];
    90: op1_00_in19 = reg_0265;
    91: op1_00_in19 = reg_0723;
    92: op1_00_in19 = reg_0526;
    93: op1_00_in19 = imem02_in[119:116];
    94: op1_00_in19 = reg_0392;
    95: op1_00_in19 = reg_0240;
    96: op1_00_in19 = reg_0210;
    default: op1_00_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_00_inv19 = 1;
    10: op1_00_inv19 = 1;
    14: op1_00_inv19 = 1;
    17: op1_00_inv19 = 1;
    18: op1_00_inv19 = 1;
    21: op1_00_inv19 = 1;
    22: op1_00_inv19 = 1;
    25: op1_00_inv19 = 1;
    29: op1_00_inv19 = 1;
    35: op1_00_inv19 = 1;
    40: op1_00_inv19 = 1;
    43: op1_00_inv19 = 1;
    44: op1_00_inv19 = 1;
    45: op1_00_inv19 = 1;
    46: op1_00_inv19 = 1;
    53: op1_00_inv19 = 1;
    55: op1_00_inv19 = 1;
    57: op1_00_inv19 = 1;
    66: op1_00_inv19 = 1;
    71: op1_00_inv19 = 1;
    76: op1_00_inv19 = 1;
    79: op1_00_inv19 = 1;
    84: op1_00_inv19 = 1;
    86: op1_00_inv19 = 1;
    87: op1_00_inv19 = 1;
    88: op1_00_inv19 = 1;
    89: op1_00_inv19 = 1;
    93: op1_00_inv19 = 1;
    94: op1_00_inv19 = 1;
    95: op1_00_inv19 = 1;
    default: op1_00_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in20 = reg_0207;
    5: op1_00_in20 = reg_0264;
    6: op1_00_in20 = reg_0499;
    7: op1_00_in20 = imem05_in[23:20];
    9: op1_00_in20 = imem02_in[103:100];
    47: op1_00_in20 = imem02_in[103:100];
    10: op1_00_in20 = reg_0664;
    11: op1_00_in20 = imem07_in[75:72];
    12: op1_00_in20 = reg_0824;
    13: op1_00_in20 = imem06_in[71:68];
    14: op1_00_in20 = imem01_in[75:72];
    15: op1_00_in20 = reg_0525;
    16: op1_00_in20 = reg_0532;
    17: op1_00_in20 = reg_0368;
    18: op1_00_in20 = reg_0617;
    19: op1_00_in20 = reg_0749;
    20: op1_00_in20 = imem04_in[83:80];
    21: op1_00_in20 = imem07_in[59:56];
    22: op1_00_in20 = reg_0497;
    23: op1_00_in20 = reg_0744;
    24: op1_00_in20 = reg_0357;
    25: op1_00_in20 = imem04_in[59:56];
    26: op1_00_in20 = reg_0192;
    27: op1_00_in20 = reg_0547;
    28: op1_00_in20 = reg_0725;
    29: op1_00_in20 = imem01_in[87:84];
    30: op1_00_in20 = reg_0510;
    32: op1_00_in20 = imem01_in[95:92];
    33: op1_00_in20 = reg_0515;
    34: op1_00_in20 = reg_0715;
    35: op1_00_in20 = imem07_in[79:76];
    36: op1_00_in20 = reg_0164;
    37: op1_00_in20 = reg_0241;
    38: op1_00_in20 = reg_0205;
    39: op1_00_in20 = reg_0757;
    40: op1_00_in20 = reg_0665;
    41: op1_00_in20 = reg_0276;
    43: op1_00_in20 = imem01_in[115:112];
    44: op1_00_in20 = reg_0587;
    45: op1_00_in20 = imem06_in[43:40];
    46: op1_00_in20 = reg_0198;
    48: op1_00_in20 = reg_0154;
    49: op1_00_in20 = reg_0038;
    50: op1_00_in20 = reg_0787;
    51: op1_00_in20 = reg_0583;
    52: op1_00_in20 = reg_0600;
    53: op1_00_in20 = reg_0554;
    54: op1_00_in20 = reg_0058;
    55: op1_00_in20 = reg_0613;
    57: op1_00_in20 = reg_0157;
    58: op1_00_in20 = imem06_in[111:108];
    59: op1_00_in20 = imem01_in[3:0];
    60: op1_00_in20 = reg_0441;
    61: op1_00_in20 = reg_0760;
    95: op1_00_in20 = reg_0760;
    62: op1_00_in20 = imem04_in[3:0];
    63: op1_00_in20 = reg_0309;
    64: op1_00_in20 = reg_0291;
    65: op1_00_in20 = reg_0298;
    66: op1_00_in20 = reg_0519;
    67: op1_00_in20 = imem06_in[127:124];
    68: op1_00_in20 = reg_0275;
    69: op1_00_in20 = reg_0076;
    71: op1_00_in20 = reg_0747;
    72: op1_00_in20 = reg_0816;
    73: op1_00_in20 = imem07_in[15:12];
    75: op1_00_in20 = imem01_in[63:60];
    76: op1_00_in20 = imem01_in[43:40];
    77: op1_00_in20 = reg_0807;
    78: op1_00_in20 = reg_0025;
    79: op1_00_in20 = imem06_in[83:80];
    82: op1_00_in20 = imem05_in[123:120];
    83: op1_00_in20 = reg_0317;
    84: op1_00_in20 = reg_0249;
    85: op1_00_in20 = reg_0445;
    86: op1_00_in20 = reg_0817;
    87: op1_00_in20 = reg_0598;
    88: op1_00_in20 = reg_0183;
    89: op1_00_in20 = imem05_in[55:52];
    90: op1_00_in20 = reg_0260;
    91: op1_00_in20 = reg_0161;
    92: op1_00_in20 = imem03_in[3:0];
    93: op1_00_in20 = reg_0042;
    94: op1_00_in20 = reg_0083;
    96: op1_00_in20 = reg_0209;
    default: op1_00_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv20 = 1;
    5: op1_00_inv20 = 1;
    9: op1_00_inv20 = 1;
    11: op1_00_inv20 = 1;
    15: op1_00_inv20 = 1;
    19: op1_00_inv20 = 1;
    20: op1_00_inv20 = 1;
    23: op1_00_inv20 = 1;
    24: op1_00_inv20 = 1;
    27: op1_00_inv20 = 1;
    29: op1_00_inv20 = 1;
    33: op1_00_inv20 = 1;
    34: op1_00_inv20 = 1;
    35: op1_00_inv20 = 1;
    36: op1_00_inv20 = 1;
    38: op1_00_inv20 = 1;
    41: op1_00_inv20 = 1;
    43: op1_00_inv20 = 1;
    44: op1_00_inv20 = 1;
    45: op1_00_inv20 = 1;
    47: op1_00_inv20 = 1;
    53: op1_00_inv20 = 1;
    57: op1_00_inv20 = 1;
    58: op1_00_inv20 = 1;
    59: op1_00_inv20 = 1;
    64: op1_00_inv20 = 1;
    67: op1_00_inv20 = 1;
    68: op1_00_inv20 = 1;
    69: op1_00_inv20 = 1;
    73: op1_00_inv20 = 1;
    77: op1_00_inv20 = 1;
    82: op1_00_inv20 = 1;
    83: op1_00_inv20 = 1;
    84: op1_00_inv20 = 1;
    86: op1_00_inv20 = 1;
    87: op1_00_inv20 = 1;
    89: op1_00_inv20 = 1;
    90: op1_00_inv20 = 1;
    94: op1_00_inv20 = 1;
    96: op1_00_inv20 = 1;
    default: op1_00_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in21 = reg_0194;
    5: op1_00_in21 = reg_0265;
    6: op1_00_in21 = reg_0498;
    7: op1_00_in21 = imem05_in[27:24];
    9: op1_00_in21 = imem02_in[119:116];
    10: op1_00_in21 = reg_0660;
    11: op1_00_in21 = imem07_in[99:96];
    12: op1_00_in21 = reg_0499;
    13: op1_00_in21 = imem06_in[99:96];
    14: op1_00_in21 = imem01_in[83:80];
    15: op1_00_in21 = reg_0215;
    50: op1_00_in21 = reg_0215;
    16: op1_00_in21 = reg_0559;
    17: op1_00_in21 = reg_0039;
    18: op1_00_in21 = reg_0618;
    19: op1_00_in21 = imem07_in[31:28];
    20: op1_00_in21 = imem04_in[87:84];
    21: op1_00_in21 = imem07_in[107:104];
    22: op1_00_in21 = reg_0500;
    23: op1_00_in21 = reg_0734;
    24: op1_00_in21 = reg_0358;
    25: op1_00_in21 = imem04_in[71:68];
    26: op1_00_in21 = imem01_in[63:60];
    27: op1_00_in21 = reg_0301;
    28: op1_00_in21 = reg_0709;
    29: op1_00_in21 = imem01_in[99:96];
    75: op1_00_in21 = imem01_in[99:96];
    30: op1_00_in21 = reg_0283;
    32: op1_00_in21 = reg_0512;
    33: op1_00_in21 = reg_0487;
    34: op1_00_in21 = reg_0700;
    78: op1_00_in21 = reg_0700;
    35: op1_00_in21 = reg_0712;
    36: op1_00_in21 = reg_0170;
    37: op1_00_in21 = reg_0505;
    38: op1_00_in21 = reg_0202;
    39: op1_00_in21 = imem03_in[7:4];
    40: op1_00_in21 = reg_0348;
    41: op1_00_in21 = reg_0224;
    43: op1_00_in21 = reg_0501;
    44: op1_00_in21 = reg_0589;
    45: op1_00_in21 = imem06_in[63:60];
    46: op1_00_in21 = reg_0201;
    47: op1_00_in21 = imem02_in[107:104];
    48: op1_00_in21 = reg_0143;
    49: op1_00_in21 = reg_0764;
    51: op1_00_in21 = reg_0592;
    52: op1_00_in21 = reg_0595;
    53: op1_00_in21 = reg_0536;
    54: op1_00_in21 = reg_0305;
    55: op1_00_in21 = reg_0577;
    57: op1_00_in21 = reg_0176;
    58: op1_00_in21 = reg_0115;
    59: op1_00_in21 = imem01_in[27:24];
    60: op1_00_in21 = reg_0449;
    61: op1_00_in21 = reg_0306;
    62: op1_00_in21 = imem04_in[15:12];
    63: op1_00_in21 = reg_0102;
    64: op1_00_in21 = reg_0624;
    65: op1_00_in21 = reg_0606;
    66: op1_00_in21 = reg_0578;
    67: op1_00_in21 = reg_0299;
    68: op1_00_in21 = reg_0352;
    69: op1_00_in21 = reg_0071;
    71: op1_00_in21 = reg_0007;
    72: op1_00_in21 = reg_0270;
    73: op1_00_in21 = imem07_in[43:40];
    76: op1_00_in21 = imem01_in[75:72];
    77: op1_00_in21 = reg_0801;
    79: op1_00_in21 = imem06_in[87:84];
    82: op1_00_in21 = imem05_in[127:124];
    83: op1_00_in21 = reg_0493;
    84: op1_00_in21 = reg_0432;
    85: op1_00_in21 = reg_0448;
    86: op1_00_in21 = reg_0238;
    87: op1_00_in21 = imem05_in[3:0];
    88: op1_00_in21 = reg_0279;
    89: op1_00_in21 = imem05_in[63:60];
    90: op1_00_in21 = reg_0408;
    91: op1_00_in21 = reg_0167;
    92: op1_00_in21 = imem03_in[31:28];
    93: op1_00_in21 = reg_0530;
    94: op1_00_in21 = reg_0702;
    95: op1_00_in21 = reg_0673;
    96: op1_00_in21 = reg_0207;
    default: op1_00_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv21 = 1;
    12: op1_00_inv21 = 1;
    15: op1_00_inv21 = 1;
    16: op1_00_inv21 = 1;
    17: op1_00_inv21 = 1;
    21: op1_00_inv21 = 1;
    22: op1_00_inv21 = 1;
    23: op1_00_inv21 = 1;
    25: op1_00_inv21 = 1;
    28: op1_00_inv21 = 1;
    33: op1_00_inv21 = 1;
    34: op1_00_inv21 = 1;
    35: op1_00_inv21 = 1;
    36: op1_00_inv21 = 1;
    37: op1_00_inv21 = 1;
    38: op1_00_inv21 = 1;
    39: op1_00_inv21 = 1;
    40: op1_00_inv21 = 1;
    41: op1_00_inv21 = 1;
    43: op1_00_inv21 = 1;
    44: op1_00_inv21 = 1;
    45: op1_00_inv21 = 1;
    46: op1_00_inv21 = 1;
    47: op1_00_inv21 = 1;
    50: op1_00_inv21 = 1;
    54: op1_00_inv21 = 1;
    55: op1_00_inv21 = 1;
    57: op1_00_inv21 = 1;
    58: op1_00_inv21 = 1;
    59: op1_00_inv21 = 1;
    61: op1_00_inv21 = 1;
    62: op1_00_inv21 = 1;
    64: op1_00_inv21 = 1;
    65: op1_00_inv21 = 1;
    67: op1_00_inv21 = 1;
    68: op1_00_inv21 = 1;
    69: op1_00_inv21 = 1;
    75: op1_00_inv21 = 1;
    77: op1_00_inv21 = 1;
    78: op1_00_inv21 = 1;
    79: op1_00_inv21 = 1;
    83: op1_00_inv21 = 1;
    84: op1_00_inv21 = 1;
    85: op1_00_inv21 = 1;
    86: op1_00_inv21 = 1;
    88: op1_00_inv21 = 1;
    89: op1_00_inv21 = 1;
    92: op1_00_inv21 = 1;
    93: op1_00_inv21 = 1;
    94: op1_00_inv21 = 1;
    default: op1_00_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in22 = reg_0201;
    5: op1_00_in22 = reg_0266;
    6: op1_00_in22 = reg_0218;
    7: op1_00_in22 = imem05_in[63:60];
    9: op1_00_in22 = reg_0666;
    10: op1_00_in22 = reg_0639;
    11: op1_00_in22 = reg_0704;
    21: op1_00_in22 = reg_0704;
    12: op1_00_in22 = reg_0825;
    13: op1_00_in22 = imem06_in[115:112];
    14: op1_00_in22 = imem01_in[103:100];
    15: op1_00_in22 = reg_0216;
    16: op1_00_in22 = reg_0556;
    17: op1_00_in22 = reg_0813;
    18: op1_00_in22 = reg_0627;
    19: op1_00_in22 = imem07_in[39:36];
    20: op1_00_in22 = imem04_in[99:96];
    22: op1_00_in22 = reg_0499;
    23: op1_00_in22 = reg_0128;
    24: op1_00_in22 = reg_0354;
    25: op1_00_in22 = imem04_in[79:76];
    26: op1_00_in22 = imem01_in[71:68];
    27: op1_00_in22 = reg_0280;
    28: op1_00_in22 = reg_0718;
    29: op1_00_in22 = imem01_in[127:124];
    30: op1_00_in22 = reg_0534;
    32: op1_00_in22 = reg_0772;
    33: op1_00_in22 = reg_0548;
    34: op1_00_in22 = reg_0436;
    35: op1_00_in22 = reg_0729;
    37: op1_00_in22 = reg_0233;
    38: op1_00_in22 = imem01_in[7:4];
    39: op1_00_in22 = imem03_in[15:12];
    40: op1_00_in22 = reg_0356;
    41: op1_00_in22 = reg_0132;
    43: op1_00_in22 = reg_0497;
    44: op1_00_in22 = reg_0600;
    45: op1_00_in22 = imem06_in[67:64];
    46: op1_00_in22 = reg_0196;
    47: op1_00_in22 = reg_0337;
    48: op1_00_in22 = imem06_in[51:48];
    49: op1_00_in22 = reg_0242;
    50: op1_00_in22 = reg_0742;
    51: op1_00_in22 = reg_0750;
    90: op1_00_in22 = reg_0750;
    52: op1_00_in22 = reg_0568;
    53: op1_00_in22 = reg_0516;
    54: op1_00_in22 = reg_0501;
    55: op1_00_in22 = reg_0773;
    57: op1_00_in22 = reg_0158;
    58: op1_00_in22 = reg_0349;
    59: op1_00_in22 = imem01_in[59:56];
    60: op1_00_in22 = reg_0160;
    61: op1_00_in22 = reg_0217;
    62: op1_00_in22 = imem04_in[71:68];
    63: op1_00_in22 = reg_0257;
    64: op1_00_in22 = reg_0370;
    65: op1_00_in22 = reg_0619;
    66: op1_00_in22 = reg_0405;
    67: op1_00_in22 = reg_0369;
    68: op1_00_in22 = reg_0365;
    69: op1_00_in22 = reg_0617;
    71: op1_00_in22 = reg_0800;
    72: op1_00_in22 = reg_0375;
    73: op1_00_in22 = imem07_in[75:72];
    75: op1_00_in22 = imem01_in[115:112];
    76: op1_00_in22 = imem01_in[115:112];
    77: op1_00_in22 = imem04_in[3:0];
    78: op1_00_in22 = reg_0777;
    79: op1_00_in22 = reg_0291;
    82: op1_00_in22 = reg_0791;
    83: op1_00_in22 = reg_0319;
    84: op1_00_in22 = reg_0305;
    85: op1_00_in22 = reg_0181;
    86: op1_00_in22 = reg_0038;
    87: op1_00_in22 = imem05_in[23:20];
    89: op1_00_in22 = imem05_in[75:72];
    91: op1_00_in22 = reg_0784;
    92: op1_00_in22 = imem03_in[43:40];
    93: op1_00_in22 = reg_0647;
    94: op1_00_in22 = reg_0362;
    95: op1_00_in22 = reg_0672;
    96: op1_00_in22 = reg_0211;
    default: op1_00_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv22 = 1;
    7: op1_00_inv22 = 1;
    9: op1_00_inv22 = 1;
    11: op1_00_inv22 = 1;
    12: op1_00_inv22 = 1;
    14: op1_00_inv22 = 1;
    15: op1_00_inv22 = 1;
    16: op1_00_inv22 = 1;
    17: op1_00_inv22 = 1;
    19: op1_00_inv22 = 1;
    21: op1_00_inv22 = 1;
    22: op1_00_inv22 = 1;
    24: op1_00_inv22 = 1;
    27: op1_00_inv22 = 1;
    28: op1_00_inv22 = 1;
    29: op1_00_inv22 = 1;
    32: op1_00_inv22 = 1;
    33: op1_00_inv22 = 1;
    35: op1_00_inv22 = 1;
    37: op1_00_inv22 = 1;
    39: op1_00_inv22 = 1;
    40: op1_00_inv22 = 1;
    48: op1_00_inv22 = 1;
    50: op1_00_inv22 = 1;
    54: op1_00_inv22 = 1;
    55: op1_00_inv22 = 1;
    57: op1_00_inv22 = 1;
    58: op1_00_inv22 = 1;
    59: op1_00_inv22 = 1;
    60: op1_00_inv22 = 1;
    62: op1_00_inv22 = 1;
    63: op1_00_inv22 = 1;
    64: op1_00_inv22 = 1;
    71: op1_00_inv22 = 1;
    72: op1_00_inv22 = 1;
    75: op1_00_inv22 = 1;
    78: op1_00_inv22 = 1;
    79: op1_00_inv22 = 1;
    82: op1_00_inv22 = 1;
    84: op1_00_inv22 = 1;
    85: op1_00_inv22 = 1;
    86: op1_00_inv22 = 1;
    87: op1_00_inv22 = 1;
    89: op1_00_inv22 = 1;
    90: op1_00_inv22 = 1;
    91: op1_00_inv22 = 1;
    92: op1_00_inv22 = 1;
    93: op1_00_inv22 = 1;
    95: op1_00_inv22 = 1;
    96: op1_00_inv22 = 1;
    default: op1_00_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in23 = reg_0190;
    5: op1_00_in23 = reg_0139;
    6: op1_00_in23 = reg_0219;
    7: op1_00_in23 = imem05_in[75:72];
    9: op1_00_in23 = reg_0653;
    75: op1_00_in23 = reg_0653;
    10: op1_00_in23 = reg_0640;
    11: op1_00_in23 = reg_0723;
    12: op1_00_in23 = reg_0778;
    13: op1_00_in23 = reg_0628;
    14: op1_00_in23 = imem01_in[107:104];
    15: op1_00_in23 = reg_0248;
    37: op1_00_in23 = reg_0248;
    16: op1_00_in23 = reg_0294;
    17: op1_00_in23 = reg_0815;
    18: op1_00_in23 = reg_0622;
    19: op1_00_in23 = imem07_in[83:80];
    73: op1_00_in23 = imem07_in[83:80];
    20: op1_00_in23 = imem04_in[107:104];
    21: op1_00_in23 = reg_0703;
    22: op1_00_in23 = reg_0825;
    23: op1_00_in23 = reg_0130;
    24: op1_00_in23 = reg_0346;
    47: op1_00_in23 = reg_0346;
    25: op1_00_in23 = reg_0315;
    26: op1_00_in23 = imem01_in[87:84];
    27: op1_00_in23 = reg_0050;
    28: op1_00_in23 = reg_0421;
    29: op1_00_in23 = reg_0758;
    30: op1_00_in23 = reg_0529;
    32: op1_00_in23 = reg_0514;
    33: op1_00_in23 = reg_0233;
    34: op1_00_in23 = reg_0418;
    35: op1_00_in23 = reg_0715;
    38: op1_00_in23 = imem01_in[23:20];
    39: op1_00_in23 = imem03_in[47:44];
    40: op1_00_in23 = reg_0092;
    41: op1_00_in23 = reg_0145;
    43: op1_00_in23 = reg_0771;
    44: op1_00_in23 = reg_0597;
    45: op1_00_in23 = reg_0286;
    46: op1_00_in23 = reg_0195;
    48: op1_00_in23 = imem06_in[63:60];
    49: op1_00_in23 = reg_0812;
    50: op1_00_in23 = reg_0229;
    51: op1_00_in23 = reg_0578;
    67: op1_00_in23 = reg_0578;
    52: op1_00_in23 = reg_0385;
    53: op1_00_in23 = reg_0547;
    54: op1_00_in23 = reg_0075;
    55: op1_00_in23 = reg_0763;
    57: op1_00_in23 = reg_0173;
    58: op1_00_in23 = reg_0766;
    65: op1_00_in23 = reg_0766;
    59: op1_00_in23 = imem01_in[75:72];
    60: op1_00_in23 = reg_0166;
    61: op1_00_in23 = reg_0567;
    62: op1_00_in23 = imem04_in[79:76];
    63: op1_00_in23 = reg_0732;
    64: op1_00_in23 = reg_0609;
    66: op1_00_in23 = reg_0583;
    68: op1_00_in23 = reg_0081;
    69: op1_00_in23 = reg_0626;
    71: op1_00_in23 = reg_0008;
    72: op1_00_in23 = reg_0576;
    76: op1_00_in23 = imem01_in[119:116];
    77: op1_00_in23 = imem04_in[35:32];
    78: op1_00_in23 = reg_0657;
    79: op1_00_in23 = reg_0619;
    82: op1_00_in23 = reg_0337;
    83: op1_00_in23 = reg_0350;
    84: op1_00_in23 = reg_0629;
    85: op1_00_in23 = reg_0099;
    86: op1_00_in23 = reg_0293;
    87: op1_00_in23 = imem05_in[31:28];
    89: op1_00_in23 = imem05_in[91:88];
    90: op1_00_in23 = reg_0608;
    91: op1_00_in23 = reg_0712;
    92: op1_00_in23 = imem03_in[67:64];
    93: op1_00_in23 = reg_0753;
    94: op1_00_in23 = reg_0341;
    95: op1_00_in23 = reg_0677;
    96: op1_00_in23 = reg_0213;
    default: op1_00_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    12: op1_00_inv23 = 1;
    15: op1_00_inv23 = 1;
    16: op1_00_inv23 = 1;
    19: op1_00_inv23 = 1;
    22: op1_00_inv23 = 1;
    23: op1_00_inv23 = 1;
    24: op1_00_inv23 = 1;
    28: op1_00_inv23 = 1;
    34: op1_00_inv23 = 1;
    35: op1_00_inv23 = 1;
    40: op1_00_inv23 = 1;
    43: op1_00_inv23 = 1;
    48: op1_00_inv23 = 1;
    50: op1_00_inv23 = 1;
    51: op1_00_inv23 = 1;
    52: op1_00_inv23 = 1;
    53: op1_00_inv23 = 1;
    55: op1_00_inv23 = 1;
    57: op1_00_inv23 = 1;
    58: op1_00_inv23 = 1;
    61: op1_00_inv23 = 1;
    62: op1_00_inv23 = 1;
    64: op1_00_inv23 = 1;
    66: op1_00_inv23 = 1;
    67: op1_00_inv23 = 1;
    69: op1_00_inv23 = 1;
    73: op1_00_inv23 = 1;
    75: op1_00_inv23 = 1;
    76: op1_00_inv23 = 1;
    79: op1_00_inv23 = 1;
    82: op1_00_inv23 = 1;
    83: op1_00_inv23 = 1;
    85: op1_00_inv23 = 1;
    90: op1_00_inv23 = 1;
    91: op1_00_inv23 = 1;
    94: op1_00_inv23 = 1;
    95: op1_00_inv23 = 1;
    96: op1_00_inv23 = 1;
    default: op1_00_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in24 = reg_0202;
    5: op1_00_in24 = imem06_in[3:0];
    6: op1_00_in24 = reg_0123;
    7: op1_00_in24 = imem05_in[99:96];
    9: op1_00_in24 = reg_0664;
    78: op1_00_in24 = reg_0664;
    10: op1_00_in24 = reg_0662;
    11: op1_00_in24 = reg_0425;
    12: op1_00_in24 = reg_0232;
    13: op1_00_in24 = reg_0625;
    14: op1_00_in24 = reg_0501;
    15: op1_00_in24 = reg_0237;
    16: op1_00_in24 = reg_0297;
    17: op1_00_in24 = reg_0005;
    18: op1_00_in24 = reg_0392;
    52: op1_00_in24 = reg_0392;
    19: op1_00_in24 = imem07_in[103:100];
    20: op1_00_in24 = imem04_in[115:112];
    21: op1_00_in24 = reg_0712;
    22: op1_00_in24 = reg_0778;
    23: op1_00_in24 = reg_0131;
    24: op1_00_in24 = reg_0347;
    25: op1_00_in24 = reg_0328;
    26: op1_00_in24 = reg_0336;
    27: op1_00_in24 = reg_0065;
    28: op1_00_in24 = reg_0440;
    29: op1_00_in24 = reg_0496;
    30: op1_00_in24 = reg_0265;
    32: op1_00_in24 = reg_0519;
    33: op1_00_in24 = reg_0217;
    34: op1_00_in24 = reg_0419;
    35: op1_00_in24 = reg_0441;
    37: op1_00_in24 = reg_0243;
    38: op1_00_in24 = imem01_in[43:40];
    96: op1_00_in24 = imem01_in[43:40];
    39: op1_00_in24 = imem03_in[127:124];
    40: op1_00_in24 = reg_0770;
    41: op1_00_in24 = reg_0154;
    43: op1_00_in24 = reg_0515;
    44: op1_00_in24 = reg_0755;
    45: op1_00_in24 = reg_0633;
    46: op1_00_in24 = imem01_in[7:4];
    47: op1_00_in24 = reg_0638;
    66: op1_00_in24 = reg_0638;
    48: op1_00_in24 = imem06_in[71:68];
    49: op1_00_in24 = reg_0372;
    50: op1_00_in24 = reg_0224;
    51: op1_00_in24 = reg_0384;
    53: op1_00_in24 = reg_0303;
    54: op1_00_in24 = reg_0549;
    55: op1_00_in24 = reg_0764;
    58: op1_00_in24 = reg_0369;
    65: op1_00_in24 = reg_0369;
    59: op1_00_in24 = imem01_in[107:104];
    60: op1_00_in24 = reg_0157;
    61: op1_00_in24 = reg_0502;
    62: op1_00_in24 = imem04_in[87:84];
    63: op1_00_in24 = reg_0086;
    64: op1_00_in24 = reg_0339;
    67: op1_00_in24 = reg_0608;
    68: op1_00_in24 = reg_0095;
    69: op1_00_in24 = reg_0614;
    71: op1_00_in24 = reg_0009;
    72: op1_00_in24 = reg_0573;
    73: op1_00_in24 = reg_0728;
    75: op1_00_in24 = reg_0741;
    76: op1_00_in24 = reg_0376;
    77: op1_00_in24 = imem04_in[103:100];
    79: op1_00_in24 = reg_0238;
    82: op1_00_in24 = reg_0736;
    83: op1_00_in24 = reg_0329;
    84: op1_00_in24 = reg_0050;
    85: op1_00_in24 = reg_0185;
    86: op1_00_in24 = reg_0260;
    87: op1_00_in24 = imem05_in[55:52];
    89: op1_00_in24 = imem05_in[111:108];
    90: op1_00_in24 = reg_0512;
    91: op1_00_in24 = reg_0103;
    92: op1_00_in24 = imem03_in[75:72];
    93: op1_00_in24 = reg_0322;
    94: op1_00_in24 = reg_0345;
    95: op1_00_in24 = reg_0121;
    default: op1_00_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv24 = 1;
    9: op1_00_inv24 = 1;
    10: op1_00_inv24 = 1;
    13: op1_00_inv24 = 1;
    14: op1_00_inv24 = 1;
    19: op1_00_inv24 = 1;
    20: op1_00_inv24 = 1;
    21: op1_00_inv24 = 1;
    22: op1_00_inv24 = 1;
    23: op1_00_inv24 = 1;
    24: op1_00_inv24 = 1;
    25: op1_00_inv24 = 1;
    27: op1_00_inv24 = 1;
    29: op1_00_inv24 = 1;
    30: op1_00_inv24 = 1;
    33: op1_00_inv24 = 1;
    34: op1_00_inv24 = 1;
    38: op1_00_inv24 = 1;
    39: op1_00_inv24 = 1;
    40: op1_00_inv24 = 1;
    43: op1_00_inv24 = 1;
    47: op1_00_inv24 = 1;
    48: op1_00_inv24 = 1;
    50: op1_00_inv24 = 1;
    52: op1_00_inv24 = 1;
    53: op1_00_inv24 = 1;
    54: op1_00_inv24 = 1;
    60: op1_00_inv24 = 1;
    61: op1_00_inv24 = 1;
    63: op1_00_inv24 = 1;
    65: op1_00_inv24 = 1;
    66: op1_00_inv24 = 1;
    67: op1_00_inv24 = 1;
    68: op1_00_inv24 = 1;
    71: op1_00_inv24 = 1;
    72: op1_00_inv24 = 1;
    77: op1_00_inv24 = 1;
    79: op1_00_inv24 = 1;
    84: op1_00_inv24 = 1;
    86: op1_00_inv24 = 1;
    87: op1_00_inv24 = 1;
    90: op1_00_inv24 = 1;
    91: op1_00_inv24 = 1;
    96: op1_00_inv24 = 1;
    default: op1_00_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in25 = reg_0195;
    5: op1_00_in25 = imem06_in[7:4];
    6: op1_00_in25 = imem02_in[39:36];
    7: op1_00_in25 = imem05_in[107:104];
    9: op1_00_in25 = reg_0657;
    10: op1_00_in25 = reg_0665;
    11: op1_00_in25 = reg_0441;
    12: op1_00_in25 = reg_0233;
    13: op1_00_in25 = reg_0616;
    14: op1_00_in25 = reg_0514;
    15: op1_00_in25 = reg_0245;
    16: op1_00_in25 = reg_0295;
    17: op1_00_in25 = imem07_in[63:60];
    18: op1_00_in25 = reg_0383;
    19: op1_00_in25 = imem07_in[107:104];
    20: op1_00_in25 = reg_0544;
    21: op1_00_in25 = reg_0706;
    22: op1_00_in25 = reg_0516;
    23: op1_00_in25 = imem06_in[15:12];
    24: op1_00_in25 = reg_0092;
    25: op1_00_in25 = reg_0542;
    26: op1_00_in25 = reg_0496;
    27: op1_00_in25 = reg_0077;
    28: op1_00_in25 = reg_0435;
    29: op1_00_in25 = reg_0822;
    30: op1_00_in25 = reg_0286;
    32: op1_00_in25 = reg_0825;
    33: op1_00_in25 = reg_0502;
    34: op1_00_in25 = reg_0439;
    35: op1_00_in25 = reg_0445;
    37: op1_00_in25 = reg_0249;
    38: op1_00_in25 = imem01_in[47:44];
    39: op1_00_in25 = reg_0582;
    40: op1_00_in25 = reg_0082;
    41: op1_00_in25 = reg_0139;
    43: op1_00_in25 = reg_0548;
    44: op1_00_in25 = reg_0569;
    45: op1_00_in25 = reg_0278;
    46: op1_00_in25 = imem01_in[31:28];
    47: op1_00_in25 = reg_0662;
    48: op1_00_in25 = imem06_in[111:108];
    49: op1_00_in25 = reg_0620;
    50: op1_00_in25 = reg_0277;
    51: op1_00_in25 = reg_0564;
    52: op1_00_in25 = reg_0397;
    53: op1_00_in25 = reg_0050;
    54: op1_00_in25 = reg_0296;
    55: op1_00_in25 = reg_0777;
    58: op1_00_in25 = reg_0578;
    59: op1_00_in25 = imem01_in[115:112];
    61: op1_00_in25 = reg_0290;
    62: op1_00_in25 = imem04_in[95:92];
    63: op1_00_in25 = reg_0151;
    64: op1_00_in25 = reg_0613;
    86: op1_00_in25 = reg_0613;
    65: op1_00_in25 = reg_0408;
    66: op1_00_in25 = reg_0593;
    67: op1_00_in25 = imem07_in[67:64];
    68: op1_00_in25 = reg_0769;
    69: op1_00_in25 = reg_0078;
    71: op1_00_in25 = imem04_in[15:12];
    72: op1_00_in25 = reg_0652;
    73: op1_00_in25 = reg_0720;
    75: op1_00_in25 = reg_0131;
    76: op1_00_in25 = reg_0111;
    77: op1_00_in25 = imem04_in[107:104];
    78: op1_00_in25 = reg_0752;
    79: op1_00_in25 = reg_0404;
    82: op1_00_in25 = reg_0788;
    83: op1_00_in25 = reg_0648;
    84: op1_00_in25 = reg_0065;
    87: op1_00_in25 = imem05_in[103:100];
    89: op1_00_in25 = imem05_in[115:112];
    90: op1_00_in25 = reg_0663;
    91: op1_00_in25 = reg_0051;
    92: op1_00_in25 = imem03_in[87:84];
    93: op1_00_in25 = reg_0344;
    94: op1_00_in25 = reg_0342;
    95: op1_00_in25 = imem02_in[11:8];
    96: op1_00_in25 = imem01_in[55:52];
    default: op1_00_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv25 = 1;
    5: op1_00_inv25 = 1;
    7: op1_00_inv25 = 1;
    15: op1_00_inv25 = 1;
    16: op1_00_inv25 = 1;
    18: op1_00_inv25 = 1;
    20: op1_00_inv25 = 1;
    21: op1_00_inv25 = 1;
    22: op1_00_inv25 = 1;
    23: op1_00_inv25 = 1;
    26: op1_00_inv25 = 1;
    28: op1_00_inv25 = 1;
    29: op1_00_inv25 = 1;
    34: op1_00_inv25 = 1;
    37: op1_00_inv25 = 1;
    38: op1_00_inv25 = 1;
    40: op1_00_inv25 = 1;
    45: op1_00_inv25 = 1;
    46: op1_00_inv25 = 1;
    47: op1_00_inv25 = 1;
    49: op1_00_inv25 = 1;
    50: op1_00_inv25 = 1;
    53: op1_00_inv25 = 1;
    54: op1_00_inv25 = 1;
    55: op1_00_inv25 = 1;
    58: op1_00_inv25 = 1;
    59: op1_00_inv25 = 1;
    61: op1_00_inv25 = 1;
    64: op1_00_inv25 = 1;
    65: op1_00_inv25 = 1;
    66: op1_00_inv25 = 1;
    67: op1_00_inv25 = 1;
    69: op1_00_inv25 = 1;
    73: op1_00_inv25 = 1;
    75: op1_00_inv25 = 1;
    77: op1_00_inv25 = 1;
    78: op1_00_inv25 = 1;
    79: op1_00_inv25 = 1;
    82: op1_00_inv25 = 1;
    84: op1_00_inv25 = 1;
    86: op1_00_inv25 = 1;
    87: op1_00_inv25 = 1;
    89: op1_00_inv25 = 1;
    90: op1_00_inv25 = 1;
    91: op1_00_inv25 = 1;
    94: op1_00_inv25 = 1;
    95: op1_00_inv25 = 1;
    96: op1_00_inv25 = 1;
    default: op1_00_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in26 = imem01_in[47:44];
    5: op1_00_in26 = imem06_in[15:12];
    6: op1_00_in26 = imem02_in[75:72];
    7: op1_00_in26 = reg_0488;
    9: op1_00_in26 = reg_0639;
    10: op1_00_in26 = reg_0659;
    86: op1_00_in26 = reg_0659;
    11: op1_00_in26 = reg_0421;
    12: op1_00_in26 = reg_0511;
    13: op1_00_in26 = reg_0626;
    14: op1_00_in26 = reg_0820;
    15: op1_00_in26 = reg_0249;
    16: op1_00_in26 = reg_0298;
    17: op1_00_in26 = imem07_in[71:68];
    18: op1_00_in26 = reg_0406;
    19: op1_00_in26 = imem07_in[111:108];
    67: op1_00_in26 = imem07_in[111:108];
    20: op1_00_in26 = reg_0560;
    21: op1_00_in26 = reg_0424;
    22: op1_00_in26 = reg_0502;
    23: op1_00_in26 = imem06_in[95:92];
    24: op1_00_in26 = reg_0533;
    25: op1_00_in26 = reg_0500;
    26: op1_00_in26 = reg_0563;
    27: op1_00_in26 = reg_0063;
    28: op1_00_in26 = reg_0175;
    29: op1_00_in26 = reg_0514;
    30: op1_00_in26 = reg_0258;
    32: op1_00_in26 = reg_0333;
    33: op1_00_in26 = reg_0220;
    34: op1_00_in26 = reg_0446;
    35: op1_00_in26 = reg_0428;
    37: op1_00_in26 = reg_0124;
    38: op1_00_in26 = imem01_in[51:48];
    39: op1_00_in26 = reg_0579;
    40: op1_00_in26 = reg_0740;
    41: op1_00_in26 = imem06_in[3:0];
    43: op1_00_in26 = reg_0559;
    44: op1_00_in26 = reg_0562;
    45: op1_00_in26 = reg_0402;
    46: op1_00_in26 = imem01_in[87:84];
    47: op1_00_in26 = reg_0349;
    48: op1_00_in26 = reg_0289;
    49: op1_00_in26 = reg_0368;
    50: op1_00_in26 = reg_0285;
    51: op1_00_in26 = reg_0517;
    52: op1_00_in26 = reg_0393;
    53: op1_00_in26 = reg_0357;
    54: op1_00_in26 = reg_0288;
    55: op1_00_in26 = reg_0620;
    58: op1_00_in26 = reg_0773;
    59: op1_00_in26 = reg_0085;
    61: op1_00_in26 = reg_0506;
    62: op1_00_in26 = reg_0316;
    63: op1_00_in26 = reg_0156;
    64: op1_00_in26 = reg_0377;
    65: op1_00_in26 = reg_0813;
    90: op1_00_in26 = reg_0813;
    66: op1_00_in26 = reg_0580;
    68: op1_00_in26 = reg_0539;
    69: op1_00_in26 = reg_0065;
    71: op1_00_in26 = imem04_in[55:52];
    72: op1_00_in26 = imem07_in[3:0];
    73: op1_00_in26 = reg_0723;
    75: op1_00_in26 = reg_0241;
    76: op1_00_in26 = reg_0131;
    77: op1_00_in26 = reg_0059;
    78: op1_00_in26 = reg_0367;
    79: op1_00_in26 = reg_0038;
    82: op1_00_in26 = reg_0795;
    83: op1_00_in26 = reg_0575;
    84: op1_00_in26 = reg_0780;
    87: op1_00_in26 = imem05_in[127:124];
    89: op1_00_in26 = reg_0736;
    91: op1_00_in26 = reg_0445;
    92: op1_00_in26 = reg_0509;
    93: op1_00_in26 = reg_0359;
    94: op1_00_in26 = reg_0590;
    95: op1_00_in26 = imem02_in[27:24];
    96: op1_00_in26 = imem01_in[71:68];
    default: op1_00_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_00_inv26 = 1;
    9: op1_00_inv26 = 1;
    11: op1_00_inv26 = 1;
    12: op1_00_inv26 = 1;
    13: op1_00_inv26 = 1;
    14: op1_00_inv26 = 1;
    16: op1_00_inv26 = 1;
    17: op1_00_inv26 = 1;
    18: op1_00_inv26 = 1;
    20: op1_00_inv26 = 1;
    25: op1_00_inv26 = 1;
    27: op1_00_inv26 = 1;
    28: op1_00_inv26 = 1;
    30: op1_00_inv26 = 1;
    32: op1_00_inv26 = 1;
    33: op1_00_inv26 = 1;
    35: op1_00_inv26 = 1;
    39: op1_00_inv26 = 1;
    48: op1_00_inv26 = 1;
    52: op1_00_inv26 = 1;
    53: op1_00_inv26 = 1;
    55: op1_00_inv26 = 1;
    59: op1_00_inv26 = 1;
    61: op1_00_inv26 = 1;
    62: op1_00_inv26 = 1;
    65: op1_00_inv26 = 1;
    66: op1_00_inv26 = 1;
    67: op1_00_inv26 = 1;
    71: op1_00_inv26 = 1;
    72: op1_00_inv26 = 1;
    75: op1_00_inv26 = 1;
    78: op1_00_inv26 = 1;
    79: op1_00_inv26 = 1;
    82: op1_00_inv26 = 1;
    86: op1_00_inv26 = 1;
    87: op1_00_inv26 = 1;
    90: op1_00_inv26 = 1;
    93: op1_00_inv26 = 1;
    95: op1_00_inv26 = 1;
    default: op1_00_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in27 = imem01_in[59:56];
    5: op1_00_in27 = imem06_in[71:68];
    6: op1_00_in27 = reg_0658;
    7: op1_00_in27 = reg_0484;
    9: op1_00_in27 = reg_0640;
    10: op1_00_in27 = reg_0667;
    11: op1_00_in27 = reg_0434;
    35: op1_00_in27 = reg_0434;
    12: op1_00_in27 = reg_0240;
    13: op1_00_in27 = reg_0618;
    14: op1_00_in27 = reg_0825;
    15: op1_00_in27 = reg_0103;
    37: op1_00_in27 = reg_0103;
    16: op1_00_in27 = reg_0288;
    17: op1_00_in27 = reg_0724;
    18: op1_00_in27 = reg_0401;
    19: op1_00_in27 = imem07_in[119:116];
    20: op1_00_in27 = reg_0546;
    21: op1_00_in27 = reg_0430;
    22: op1_00_in27 = reg_0220;
    23: op1_00_in27 = imem06_in[103:100];
    24: op1_00_in27 = reg_0081;
    25: op1_00_in27 = reg_0305;
    26: op1_00_in27 = reg_0761;
    27: op1_00_in27 = reg_0256;
    78: op1_00_in27 = reg_0256;
    28: op1_00_in27 = reg_0162;
    29: op1_00_in27 = reg_0515;
    32: op1_00_in27 = reg_0515;
    30: op1_00_in27 = reg_0281;
    33: op1_00_in27 = reg_0105;
    34: op1_00_in27 = reg_0440;
    38: op1_00_in27 = imem01_in[95:92];
    39: op1_00_in27 = reg_0565;
    40: op1_00_in27 = imem03_in[3:0];
    41: op1_00_in27 = imem06_in[23:20];
    43: op1_00_in27 = reg_0306;
    44: op1_00_in27 = reg_0376;
    51: op1_00_in27 = reg_0376;
    45: op1_00_in27 = reg_0577;
    46: op1_00_in27 = reg_0501;
    47: op1_00_in27 = reg_0358;
    48: op1_00_in27 = reg_0624;
    49: op1_00_in27 = reg_0375;
    50: op1_00_in27 = reg_0146;
    52: op1_00_in27 = reg_0747;
    53: op1_00_in27 = reg_0520;
    54: op1_00_in27 = imem05_in[83:80];
    55: op1_00_in27 = reg_0815;
    58: op1_00_in27 = reg_0821;
    59: op1_00_in27 = reg_0733;
    61: op1_00_in27 = reg_0505;
    62: op1_00_in27 = reg_0537;
    63: op1_00_in27 = reg_0154;
    64: op1_00_in27 = reg_0405;
    86: op1_00_in27 = reg_0405;
    65: op1_00_in27 = reg_0032;
    66: op1_00_in27 = reg_0512;
    67: op1_00_in27 = reg_0728;
    68: op1_00_in27 = reg_0098;
    69: op1_00_in27 = reg_0598;
    71: op1_00_in27 = imem04_in[67:64];
    72: op1_00_in27 = imem07_in[11:8];
    73: op1_00_in27 = reg_0717;
    75: op1_00_in27 = reg_0418;
    76: op1_00_in27 = reg_0388;
    77: op1_00_in27 = reg_0262;
    79: op1_00_in27 = reg_0408;
    82: op1_00_in27 = reg_0550;
    83: op1_00_in27 = reg_0417;
    84: op1_00_in27 = imem05_in[47:44];
    87: op1_00_in27 = reg_0133;
    89: op1_00_in27 = reg_0135;
    90: op1_00_in27 = reg_0612;
    91: op1_00_in27 = reg_0267;
    92: op1_00_in27 = reg_0003;
    93: op1_00_in27 = reg_0360;
    94: op1_00_in27 = reg_0343;
    95: op1_00_in27 = imem02_in[63:60];
    96: op1_00_in27 = imem01_in[87:84];
    default: op1_00_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv27 = 1;
    9: op1_00_inv27 = 1;
    10: op1_00_inv27 = 1;
    12: op1_00_inv27 = 1;
    13: op1_00_inv27 = 1;
    16: op1_00_inv27 = 1;
    18: op1_00_inv27 = 1;
    19: op1_00_inv27 = 1;
    20: op1_00_inv27 = 1;
    21: op1_00_inv27 = 1;
    22: op1_00_inv27 = 1;
    23: op1_00_inv27 = 1;
    25: op1_00_inv27 = 1;
    26: op1_00_inv27 = 1;
    28: op1_00_inv27 = 1;
    30: op1_00_inv27 = 1;
    32: op1_00_inv27 = 1;
    41: op1_00_inv27 = 1;
    44: op1_00_inv27 = 1;
    45: op1_00_inv27 = 1;
    47: op1_00_inv27 = 1;
    48: op1_00_inv27 = 1;
    49: op1_00_inv27 = 1;
    51: op1_00_inv27 = 1;
    55: op1_00_inv27 = 1;
    58: op1_00_inv27 = 1;
    59: op1_00_inv27 = 1;
    61: op1_00_inv27 = 1;
    62: op1_00_inv27 = 1;
    65: op1_00_inv27 = 1;
    67: op1_00_inv27 = 1;
    68: op1_00_inv27 = 1;
    73: op1_00_inv27 = 1;
    75: op1_00_inv27 = 1;
    76: op1_00_inv27 = 1;
    77: op1_00_inv27 = 1;
    79: op1_00_inv27 = 1;
    82: op1_00_inv27 = 1;
    83: op1_00_inv27 = 1;
    84: op1_00_inv27 = 1;
    87: op1_00_inv27 = 1;
    89: op1_00_inv27 = 1;
    90: op1_00_inv27 = 1;
    92: op1_00_inv27 = 1;
    94: op1_00_inv27 = 1;
    96: op1_00_inv27 = 1;
    default: op1_00_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in28 = imem01_in[83:80];
    5: op1_00_in28 = imem06_in[75:72];
    6: op1_00_in28 = reg_0654;
    7: op1_00_in28 = reg_0793;
    82: op1_00_in28 = reg_0793;
    9: op1_00_in28 = reg_0648;
    10: op1_00_in28 = reg_0341;
    11: op1_00_in28 = reg_0166;
    12: op1_00_in28 = reg_0236;
    13: op1_00_in28 = reg_0348;
    14: op1_00_in28 = reg_0517;
    15: op1_00_in28 = reg_0111;
    16: op1_00_in28 = reg_0061;
    17: op1_00_in28 = reg_0729;
    18: op1_00_in28 = reg_0033;
    19: op1_00_in28 = reg_0716;
    20: op1_00_in28 = reg_0052;
    21: op1_00_in28 = reg_0436;
    22: op1_00_in28 = reg_0122;
    23: op1_00_in28 = imem06_in[119:116];
    24: op1_00_in28 = reg_0097;
    25: op1_00_in28 = reg_0265;
    26: op1_00_in28 = reg_0511;
    27: op1_00_in28 = imem05_in[87:84];
    28: op1_00_in28 = reg_0163;
    29: op1_00_in28 = reg_0507;
    32: op1_00_in28 = reg_0507;
    30: op1_00_in28 = reg_0076;
    33: op1_00_in28 = reg_0118;
    37: op1_00_in28 = reg_0118;
    34: op1_00_in28 = reg_0443;
    35: op1_00_in28 = reg_0444;
    38: op1_00_in28 = reg_0336;
    39: op1_00_in28 = reg_0039;
    40: op1_00_in28 = imem03_in[11:8];
    68: op1_00_in28 = imem03_in[11:8];
    41: op1_00_in28 = imem06_in[71:68];
    43: op1_00_in28 = reg_0054;
    44: op1_00_in28 = reg_0393;
    45: op1_00_in28 = reg_0405;
    46: op1_00_in28 = reg_0772;
    47: op1_00_in28 = reg_0350;
    48: op1_00_in28 = reg_0286;
    49: op1_00_in28 = reg_0231;
    50: op1_00_in28 = reg_0139;
    51: op1_00_in28 = reg_0389;
    52: op1_00_in28 = reg_0807;
    53: op1_00_in28 = reg_0065;
    54: op1_00_in28 = imem05_in[107:104];
    55: op1_00_in28 = reg_0040;
    58: op1_00_in28 = reg_0638;
    59: op1_00_in28 = reg_0761;
    61: op1_00_in28 = reg_0420;
    62: op1_00_in28 = reg_0554;
    63: op1_00_in28 = reg_0153;
    64: op1_00_in28 = reg_0375;
    65: op1_00_in28 = reg_0656;
    66: op1_00_in28 = reg_0028;
    67: op1_00_in28 = reg_0719;
    69: op1_00_in28 = reg_0780;
    71: op1_00_in28 = imem04_in[123:120];
    72: op1_00_in28 = imem07_in[31:28];
    73: op1_00_in28 = reg_0725;
    75: op1_00_in28 = reg_0574;
    76: op1_00_in28 = reg_0397;
    77: op1_00_in28 = reg_0553;
    78: op1_00_in28 = imem07_in[11:8];
    79: op1_00_in28 = reg_0816;
    83: op1_00_in28 = reg_0403;
    84: op1_00_in28 = reg_0791;
    86: op1_00_in28 = reg_0307;
    87: op1_00_in28 = reg_0128;
    89: op1_00_in28 = reg_0070;
    90: op1_00_in28 = reg_0657;
    91: op1_00_in28 = reg_0181;
    92: op1_00_in28 = reg_0559;
    93: op1_00_in28 = reg_0406;
    94: op1_00_in28 = reg_0132;
    95: op1_00_in28 = imem02_in[87:84];
    96: op1_00_in28 = imem01_in[115:112];
    default: op1_00_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv28 = 1;
    6: op1_00_inv28 = 1;
    7: op1_00_inv28 = 1;
    10: op1_00_inv28 = 1;
    12: op1_00_inv28 = 1;
    16: op1_00_inv28 = 1;
    17: op1_00_inv28 = 1;
    20: op1_00_inv28 = 1;
    22: op1_00_inv28 = 1;
    23: op1_00_inv28 = 1;
    26: op1_00_inv28 = 1;
    28: op1_00_inv28 = 1;
    34: op1_00_inv28 = 1;
    39: op1_00_inv28 = 1;
    43: op1_00_inv28 = 1;
    44: op1_00_inv28 = 1;
    46: op1_00_inv28 = 1;
    47: op1_00_inv28 = 1;
    49: op1_00_inv28 = 1;
    54: op1_00_inv28 = 1;
    55: op1_00_inv28 = 1;
    58: op1_00_inv28 = 1;
    61: op1_00_inv28 = 1;
    63: op1_00_inv28 = 1;
    64: op1_00_inv28 = 1;
    65: op1_00_inv28 = 1;
    67: op1_00_inv28 = 1;
    68: op1_00_inv28 = 1;
    69: op1_00_inv28 = 1;
    71: op1_00_inv28 = 1;
    75: op1_00_inv28 = 1;
    76: op1_00_inv28 = 1;
    77: op1_00_inv28 = 1;
    82: op1_00_inv28 = 1;
    84: op1_00_inv28 = 1;
    87: op1_00_inv28 = 1;
    89: op1_00_inv28 = 1;
    91: op1_00_inv28 = 1;
    93: op1_00_inv28 = 1;
    94: op1_00_inv28 = 1;
    95: op1_00_inv28 = 1;
    default: op1_00_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in29 = imem01_in[91:88];
    5: op1_00_in29 = imem06_in[79:76];
    6: op1_00_in29 = reg_0660;
    7: op1_00_in29 = reg_0495;
    9: op1_00_in29 = reg_0364;
    10: op1_00_in29 = reg_0318;
    11: op1_00_in29 = reg_0168;
    12: op1_00_in29 = reg_0508;
    13: op1_00_in29 = reg_0381;
    14: op1_00_in29 = reg_0776;
    15: op1_00_in29 = reg_0116;
    33: op1_00_in29 = reg_0116;
    16: op1_00_in29 = reg_0078;
    17: op1_00_in29 = reg_0705;
    18: op1_00_in29 = reg_0032;
    19: op1_00_in29 = reg_0731;
    20: op1_00_in29 = reg_0274;
    21: op1_00_in29 = reg_0422;
    22: op1_00_in29 = reg_0124;
    46: op1_00_in29 = reg_0124;
    23: op1_00_in29 = reg_0628;
    24: op1_00_in29 = reg_0540;
    25: op1_00_in29 = reg_0051;
    26: op1_00_in29 = reg_0248;
    27: op1_00_in29 = imem05_in[91:88];
    28: op1_00_in29 = reg_0166;
    29: op1_00_in29 = reg_0505;
    32: op1_00_in29 = reg_0505;
    30: op1_00_in29 = reg_0256;
    34: op1_00_in29 = reg_0183;
    35: op1_00_in29 = reg_0448;
    37: op1_00_in29 = reg_0100;
    38: op1_00_in29 = reg_0496;
    39: op1_00_in29 = reg_0750;
    40: op1_00_in29 = imem03_in[39:36];
    41: op1_00_in29 = imem06_in[99:96];
    43: op1_00_in29 = reg_0419;
    44: op1_00_in29 = reg_0006;
    83: op1_00_in29 = reg_0006;
    45: op1_00_in29 = reg_0775;
    47: op1_00_in29 = reg_0081;
    48: op1_00_in29 = reg_0609;
    49: op1_00_in29 = imem07_in[23:20];
    78: op1_00_in29 = imem07_in[23:20];
    50: op1_00_in29 = imem06_in[15:12];
    51: op1_00_in29 = reg_0810;
    52: op1_00_in29 = reg_0801;
    53: op1_00_in29 = reg_0075;
    54: op1_00_in29 = reg_0791;
    55: op1_00_in29 = reg_0029;
    58: op1_00_in29 = reg_0040;
    59: op1_00_in29 = reg_0649;
    61: op1_00_in29 = reg_0123;
    62: op1_00_in29 = reg_0057;
    63: op1_00_in29 = reg_0137;
    64: op1_00_in29 = reg_0638;
    65: op1_00_in29 = reg_0819;
    66: op1_00_in29 = reg_0607;
    67: op1_00_in29 = reg_0711;
    68: op1_00_in29 = imem03_in[27:24];
    69: op1_00_in29 = reg_0259;
    71: op1_00_in29 = reg_0544;
    72: op1_00_in29 = imem07_in[51:48];
    73: op1_00_in29 = reg_0729;
    75: op1_00_in29 = reg_0243;
    76: op1_00_in29 = reg_0737;
    77: op1_00_in29 = reg_0056;
    79: op1_00_in29 = reg_0512;
    82: op1_00_in29 = reg_0732;
    84: op1_00_in29 = reg_0736;
    86: op1_00_in29 = reg_0484;
    87: op1_00_in29 = reg_0090;
    89: op1_00_in29 = reg_0386;
    90: op1_00_in29 = reg_0037;
    91: op1_00_in29 = reg_0327;
    92: op1_00_in29 = reg_0591;
    93: op1_00_in29 = reg_0743;
    94: op1_00_in29 = reg_0770;
    95: op1_00_in29 = imem02_in[115:112];
    96: op1_00_in29 = imem01_in[119:116];
    default: op1_00_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_00_inv29 = 1;
    6: op1_00_inv29 = 1;
    9: op1_00_inv29 = 1;
    11: op1_00_inv29 = 1;
    12: op1_00_inv29 = 1;
    13: op1_00_inv29 = 1;
    16: op1_00_inv29 = 1;
    17: op1_00_inv29 = 1;
    19: op1_00_inv29 = 1;
    22: op1_00_inv29 = 1;
    26: op1_00_inv29 = 1;
    27: op1_00_inv29 = 1;
    28: op1_00_inv29 = 1;
    33: op1_00_inv29 = 1;
    35: op1_00_inv29 = 1;
    37: op1_00_inv29 = 1;
    38: op1_00_inv29 = 1;
    39: op1_00_inv29 = 1;
    40: op1_00_inv29 = 1;
    41: op1_00_inv29 = 1;
    43: op1_00_inv29 = 1;
    44: op1_00_inv29 = 1;
    45: op1_00_inv29 = 1;
    46: op1_00_inv29 = 1;
    47: op1_00_inv29 = 1;
    48: op1_00_inv29 = 1;
    50: op1_00_inv29 = 1;
    52: op1_00_inv29 = 1;
    53: op1_00_inv29 = 1;
    54: op1_00_inv29 = 1;
    55: op1_00_inv29 = 1;
    59: op1_00_inv29 = 1;
    62: op1_00_inv29 = 1;
    64: op1_00_inv29 = 1;
    65: op1_00_inv29 = 1;
    68: op1_00_inv29 = 1;
    71: op1_00_inv29 = 1;
    73: op1_00_inv29 = 1;
    78: op1_00_inv29 = 1;
    82: op1_00_inv29 = 1;
    86: op1_00_inv29 = 1;
    87: op1_00_inv29 = 1;
    89: op1_00_inv29 = 1;
    90: op1_00_inv29 = 1;
    91: op1_00_inv29 = 1;
    92: op1_00_inv29 = 1;
    95: op1_00_inv29 = 1;
    default: op1_00_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_00_in30 = reg_0513;
    5: op1_00_in30 = imem06_in[87:84];
    6: op1_00_in30 = reg_0661;
    7: op1_00_in30 = reg_0787;
    9: op1_00_in30 = reg_0359;
    10: op1_00_in30 = reg_0338;
    12: op1_00_in30 = reg_0111;
    13: op1_00_in30 = reg_0367;
    14: op1_00_in30 = reg_0507;
    15: op1_00_in30 = reg_0117;
    16: op1_00_in30 = reg_0066;
    17: op1_00_in30 = reg_0727;
    18: op1_00_in30 = reg_0040;
    19: op1_00_in30 = reg_0708;
    20: op1_00_in30 = reg_0302;
    21: op1_00_in30 = reg_0433;
    22: op1_00_in30 = reg_0103;
    23: op1_00_in30 = reg_0607;
    24: op1_00_in30 = reg_0531;
    25: op1_00_in30 = reg_0069;
    26: op1_00_in30 = reg_0105;
    61: op1_00_in30 = reg_0105;
    27: op1_00_in30 = imem05_in[95:92];
    28: op1_00_in30 = reg_0164;
    34: op1_00_in30 = reg_0164;
    29: op1_00_in30 = reg_0245;
    30: op1_00_in30 = imem05_in[99:96];
    32: op1_00_in30 = reg_0511;
    33: op1_00_in30 = reg_0120;
    35: op1_00_in30 = reg_0162;
    37: op1_00_in30 = imem02_in[7:4];
    38: op1_00_in30 = reg_0512;
    64: op1_00_in30 = reg_0512;
    39: op1_00_in30 = reg_0581;
    40: op1_00_in30 = imem03_in[43:40];
    41: op1_00_in30 = reg_0289;
    43: op1_00_in30 = reg_0124;
    44: op1_00_in30 = reg_0019;
    45: op1_00_in30 = reg_0329;
    46: op1_00_in30 = reg_0116;
    47: op1_00_in30 = reg_0540;
    48: op1_00_in30 = reg_0633;
    49: op1_00_in30 = imem07_in[39:36];
    50: op1_00_in30 = imem06_in[103:100];
    51: op1_00_in30 = reg_0809;
    52: op1_00_in30 = reg_0800;
    53: op1_00_in30 = reg_0399;
    54: op1_00_in30 = reg_0792;
    55: op1_00_in30 = reg_0632;
    58: op1_00_in30 = reg_0621;
    59: op1_00_in30 = reg_0825;
    62: op1_00_in30 = reg_0305;
    63: op1_00_in30 = imem06_in[7:4];
    65: op1_00_in30 = reg_0368;
    66: op1_00_in30 = reg_0813;
    67: op1_00_in30 = reg_0253;
    68: op1_00_in30 = imem03_in[63:60];
    69: op1_00_in30 = reg_0644;
    71: op1_00_in30 = reg_0087;
    72: op1_00_in30 = imem07_in[63:60];
    73: op1_00_in30 = reg_0061;
    75: op1_00_in30 = reg_0505;
    76: op1_00_in30 = reg_0110;
    77: op1_00_in30 = reg_0523;
    78: op1_00_in30 = imem07_in[47:44];
    79: op1_00_in30 = reg_0573;
    82: op1_00_in30 = reg_0386;
    83: op1_00_in30 = reg_0803;
    84: op1_00_in30 = reg_0788;
    86: op1_00_in30 = reg_0215;
    87: op1_00_in30 = reg_0489;
    89: op1_00_in30 = reg_0518;
    90: op1_00_in30 = reg_0680;
    91: op1_00_in30 = reg_0183;
    92: op1_00_in30 = reg_0318;
    93: op1_00_in30 = reg_0109;
    94: op1_00_in30 = reg_0255;
    95: op1_00_in30 = imem02_in[119:116];
    96: op1_00_in30 = imem01_in[123:120];
    default: op1_00_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_00_inv30 = 1;
    5: op1_00_inv30 = 1;
    7: op1_00_inv30 = 1;
    10: op1_00_inv30 = 1;
    18: op1_00_inv30 = 1;
    19: op1_00_inv30 = 1;
    27: op1_00_inv30 = 1;
    33: op1_00_inv30 = 1;
    35: op1_00_inv30 = 1;
    39: op1_00_inv30 = 1;
    40: op1_00_inv30 = 1;
    41: op1_00_inv30 = 1;
    43: op1_00_inv30 = 1;
    44: op1_00_inv30 = 1;
    46: op1_00_inv30 = 1;
    48: op1_00_inv30 = 1;
    49: op1_00_inv30 = 1;
    50: op1_00_inv30 = 1;
    52: op1_00_inv30 = 1;
    54: op1_00_inv30 = 1;
    61: op1_00_inv30 = 1;
    62: op1_00_inv30 = 1;
    66: op1_00_inv30 = 1;
    67: op1_00_inv30 = 1;
    69: op1_00_inv30 = 1;
    73: op1_00_inv30 = 1;
    75: op1_00_inv30 = 1;
    76: op1_00_inv30 = 1;
    78: op1_00_inv30 = 1;
    86: op1_00_inv30 = 1;
    89: op1_00_inv30 = 1;
    93: op1_00_inv30 = 1;
    default: op1_00_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_00_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_00_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in00 = reg_0514;
    5: op1_01_in00 = imem06_in[127:124];
    6: op1_01_in00 = reg_0640;
    7: op1_01_in00 = reg_0486;
    3: op1_01_in00 = imem07_in[47:44];
    8: op1_01_in00 = imem00_in[19:16];
    74: op1_01_in00 = imem00_in[19:16];
    2: op1_01_in00 = imem07_in[103:100];
    72: op1_01_in00 = imem07_in[103:100];
    9: op1_01_in00 = reg_0324;
    10: op1_01_in00 = reg_0335;
    11: op1_01_in00 = imem00_in[43:40];
    12: op1_01_in00 = reg_0099;
    1: op1_01_in00 = imem07_in[15:12];
    13: op1_01_in00 = reg_0380;
    14: op1_01_in00 = reg_0225;
    76: op1_01_in00 = reg_0225;
    15: op1_01_in00 = imem02_in[31:28];
    16: op1_01_in00 = reg_0070;
    17: op1_01_in00 = imem00_in[3:0];
    19: op1_01_in00 = imem00_in[3:0];
    57: op1_01_in00 = imem00_in[3:0];
    70: op1_01_in00 = imem00_in[3:0];
    18: op1_01_in00 = reg_0751;
    20: op1_01_in00 = reg_0290;
    21: op1_01_in00 = imem00_in[51:48];
    28: op1_01_in00 = imem00_in[51:48];
    85: op1_01_in00 = imem00_in[51:48];
    22: op1_01_in00 = reg_0104;
    23: op1_01_in00 = reg_0616;
    24: op1_01_in00 = imem03_in[3:0];
    25: op1_01_in00 = reg_0064;
    26: op1_01_in00 = reg_0122;
    27: op1_01_in00 = imem05_in[123:120];
    30: op1_01_in00 = imem05_in[123:120];
    29: op1_01_in00 = reg_0041;
    31: op1_01_in00 = imem00_in[27:24];
    32: op1_01_in00 = reg_0218;
    33: op1_01_in00 = reg_0108;
    34: op1_01_in00 = imem00_in[55:52];
    88: op1_01_in00 = imem00_in[55:52];
    35: op1_01_in00 = reg_0182;
    36: op1_01_in00 = imem00_in[39:36];
    37: op1_01_in00 = imem02_in[19:16];
    38: op1_01_in00 = reg_0771;
    39: op1_01_in00 = reg_0561;
    40: op1_01_in00 = reg_0599;
    41: op1_01_in00 = reg_0608;
    48: op1_01_in00 = reg_0608;
    42: op1_01_in00 = imem00_in[59:56];
    43: op1_01_in00 = reg_0118;
    75: op1_01_in00 = reg_0118;
    44: op1_01_in00 = reg_0012;
    45: op1_01_in00 = reg_0038;
    46: op1_01_in00 = reg_0114;
    47: op1_01_in00 = reg_0770;
    49: op1_01_in00 = imem07_in[63:60];
    50: op1_01_in00 = reg_0625;
    51: op1_01_in00 = reg_0004;
    52: op1_01_in00 = reg_0016;
    53: op1_01_in00 = reg_0068;
    54: op1_01_in00 = reg_0482;
    55: op1_01_in00 = imem07_in[11:8];
    56: op1_01_in00 = imem00_in[15:12];
    81: op1_01_in00 = imem00_in[15:12];
    58: op1_01_in00 = reg_0037;
    59: op1_01_in00 = reg_0760;
    60: op1_01_in00 = imem00_in[7:4];
    61: op1_01_in00 = reg_0073;
    62: op1_01_in00 = reg_0280;
    63: op1_01_in00 = imem06_in[43:40];
    64: op1_01_in00 = reg_0520;
    65: op1_01_in00 = imem07_in[83:80];
    66: op1_01_in00 = reg_0620;
    67: op1_01_in00 = reg_0635;
    68: op1_01_in00 = imem03_in[87:84];
    69: op1_01_in00 = imem05_in[51:48];
    71: op1_01_in00 = reg_0551;
    73: op1_01_in00 = reg_0333;
    77: op1_01_in00 = reg_0058;
    78: op1_01_in00 = imem07_in[55:52];
    79: op1_01_in00 = reg_0813;
    80: op1_01_in00 = imem00_in[31:28];
    82: op1_01_in00 = reg_0309;
    83: op1_01_in00 = reg_0007;
    84: op1_01_in00 = reg_0641;
    86: op1_01_in00 = reg_0638;
    87: op1_01_in00 = reg_0517;
    89: op1_01_in00 = reg_0399;
    90: op1_01_in00 = reg_0661;
    91: op1_01_in00 = reg_0170;
    92: op1_01_in00 = reg_0528;
    93: op1_01_in00 = reg_0095;
    94: op1_01_in00 = reg_0055;
    95: op1_01_in00 = reg_0031;
    96: op1_01_in00 = reg_0013;
    default: op1_01_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv00 = 1;
    5: op1_01_inv00 = 1;
    6: op1_01_inv00 = 1;
    17: op1_01_inv00 = 1;
    20: op1_01_inv00 = 1;
    21: op1_01_inv00 = 1;
    22: op1_01_inv00 = 1;
    24: op1_01_inv00 = 1;
    25: op1_01_inv00 = 1;
    27: op1_01_inv00 = 1;
    29: op1_01_inv00 = 1;
    30: op1_01_inv00 = 1;
    32: op1_01_inv00 = 1;
    33: op1_01_inv00 = 1;
    34: op1_01_inv00 = 1;
    35: op1_01_inv00 = 1;
    37: op1_01_inv00 = 1;
    40: op1_01_inv00 = 1;
    42: op1_01_inv00 = 1;
    43: op1_01_inv00 = 1;
    45: op1_01_inv00 = 1;
    48: op1_01_inv00 = 1;
    50: op1_01_inv00 = 1;
    51: op1_01_inv00 = 1;
    53: op1_01_inv00 = 1;
    55: op1_01_inv00 = 1;
    57: op1_01_inv00 = 1;
    58: op1_01_inv00 = 1;
    59: op1_01_inv00 = 1;
    61: op1_01_inv00 = 1;
    63: op1_01_inv00 = 1;
    67: op1_01_inv00 = 1;
    68: op1_01_inv00 = 1;
    69: op1_01_inv00 = 1;
    70: op1_01_inv00 = 1;
    71: op1_01_inv00 = 1;
    73: op1_01_inv00 = 1;
    74: op1_01_inv00 = 1;
    79: op1_01_inv00 = 1;
    82: op1_01_inv00 = 1;
    86: op1_01_inv00 = 1;
    87: op1_01_inv00 = 1;
    88: op1_01_inv00 = 1;
    89: op1_01_inv00 = 1;
    default: op1_01_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in01 = reg_0502;
    5: op1_01_in01 = reg_0625;
    6: op1_01_in01 = reg_0649;
    7: op1_01_in01 = reg_0260;
    3: op1_01_in01 = imem07_in[51:48];
    8: op1_01_in01 = imem00_in[59:56];
    36: op1_01_in01 = imem00_in[59:56];
    88: op1_01_in01 = imem00_in[59:56];
    2: op1_01_in01 = imem07_in[115:112];
    9: op1_01_in01 = reg_0353;
    10: op1_01_in01 = reg_0328;
    11: op1_01_in01 = imem00_in[99:96];
    12: op1_01_in01 = reg_0108;
    1: op1_01_in01 = imem07_in[27:24];
    13: op1_01_in01 = reg_0028;
    14: op1_01_in01 = reg_0215;
    48: op1_01_in01 = reg_0215;
    15: op1_01_in01 = imem02_in[79:76];
    16: op1_01_in01 = imem05_in[27:24];
    17: op1_01_in01 = imem00_in[27:24];
    74: op1_01_in01 = imem00_in[27:24];
    18: op1_01_in01 = imem07_in[87:84];
    65: op1_01_in01 = imem07_in[87:84];
    19: op1_01_in01 = imem00_in[55:52];
    20: op1_01_in01 = reg_0051;
    21: op1_01_in01 = imem00_in[127:124];
    22: op1_01_in01 = imem02_in[23:20];
    23: op1_01_in01 = reg_0609;
    24: op1_01_in01 = imem03_in[55:52];
    25: op1_01_in01 = imem05_in[19:16];
    26: op1_01_in01 = reg_0124;
    27: op1_01_in01 = imem05_in[127:124];
    28: op1_01_in01 = imem00_in[83:80];
    42: op1_01_in01 = imem00_in[83:80];
    29: op1_01_in01 = reg_0219;
    30: op1_01_in01 = reg_0791;
    31: op1_01_in01 = imem00_in[39:36];
    57: op1_01_in01 = imem00_in[39:36];
    32: op1_01_in01 = reg_0506;
    33: op1_01_in01 = imem02_in[7:4];
    34: op1_01_in01 = imem00_in[79:76];
    85: op1_01_in01 = imem00_in[79:76];
    35: op1_01_in01 = reg_0160;
    37: op1_01_in01 = imem02_in[51:48];
    38: op1_01_in01 = reg_0761;
    39: op1_01_in01 = reg_0568;
    40: op1_01_in01 = reg_0583;
    41: op1_01_in01 = reg_0618;
    43: op1_01_in01 = reg_0114;
    44: op1_01_in01 = reg_0002;
    45: op1_01_in01 = reg_0031;
    46: op1_01_in01 = reg_0106;
    47: op1_01_in01 = reg_0531;
    49: op1_01_in01 = imem07_in[71:68];
    50: op1_01_in01 = reg_0291;
    51: op1_01_in01 = imem04_in[59:56];
    52: op1_01_in01 = reg_0806;
    53: op1_01_in01 = reg_0275;
    54: op1_01_in01 = reg_0797;
    55: op1_01_in01 = imem07_in[83:80];
    56: op1_01_in01 = imem00_in[51:48];
    58: op1_01_in01 = reg_0236;
    59: op1_01_in01 = reg_0423;
    76: op1_01_in01 = reg_0423;
    60: op1_01_in01 = imem00_in[11:8];
    61: op1_01_in01 = reg_0104;
    75: op1_01_in01 = reg_0104;
    62: op1_01_in01 = reg_0508;
    63: op1_01_in01 = imem06_in[91:88];
    64: op1_01_in01 = reg_0700;
    66: op1_01_in01 = reg_0656;
    67: op1_01_in01 = reg_0445;
    68: op1_01_in01 = reg_0317;
    69: op1_01_in01 = imem05_in[59:56];
    70: op1_01_in01 = imem00_in[15:12];
    71: op1_01_in01 = reg_0052;
    72: op1_01_in01 = imem07_in[123:120];
    73: op1_01_in01 = reg_0439;
    77: op1_01_in01 = reg_0283;
    78: op1_01_in01 = imem07_in[67:64];
    79: op1_01_in01 = reg_0620;
    80: op1_01_in01 = imem00_in[47:44];
    81: op1_01_in01 = imem00_in[23:20];
    82: op1_01_in01 = reg_0491;
    83: op1_01_in01 = reg_0800;
    84: op1_01_in01 = reg_0793;
    86: op1_01_in01 = reg_0169;
    87: op1_01_in01 = reg_0538;
    89: op1_01_in01 = reg_0827;
    90: op1_01_in01 = reg_0632;
    91: op1_01_in01 = reg_0091;
    92: op1_01_in01 = reg_0493;
    93: op1_01_in01 = reg_0757;
    94: op1_01_in01 = reg_0526;
    95: op1_01_in01 = reg_0264;
    96: op1_01_in01 = reg_0499;
    default: op1_01_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv01 = 1;
    6: op1_01_inv01 = 1;
    7: op1_01_inv01 = 1;
    9: op1_01_inv01 = 1;
    10: op1_01_inv01 = 1;
    11: op1_01_inv01 = 1;
    12: op1_01_inv01 = 1;
    1: op1_01_inv01 = 1;
    13: op1_01_inv01 = 1;
    14: op1_01_inv01 = 1;
    18: op1_01_inv01 = 1;
    23: op1_01_inv01 = 1;
    29: op1_01_inv01 = 1;
    31: op1_01_inv01 = 1;
    35: op1_01_inv01 = 1;
    36: op1_01_inv01 = 1;
    37: op1_01_inv01 = 1;
    38: op1_01_inv01 = 1;
    40: op1_01_inv01 = 1;
    41: op1_01_inv01 = 1;
    44: op1_01_inv01 = 1;
    45: op1_01_inv01 = 1;
    47: op1_01_inv01 = 1;
    49: op1_01_inv01 = 1;
    56: op1_01_inv01 = 1;
    57: op1_01_inv01 = 1;
    58: op1_01_inv01 = 1;
    59: op1_01_inv01 = 1;
    63: op1_01_inv01 = 1;
    68: op1_01_inv01 = 1;
    70: op1_01_inv01 = 1;
    73: op1_01_inv01 = 1;
    74: op1_01_inv01 = 1;
    75: op1_01_inv01 = 1;
    77: op1_01_inv01 = 1;
    78: op1_01_inv01 = 1;
    80: op1_01_inv01 = 1;
    81: op1_01_inv01 = 1;
    82: op1_01_inv01 = 1;
    83: op1_01_inv01 = 1;
    86: op1_01_inv01 = 1;
    88: op1_01_inv01 = 1;
    90: op1_01_inv01 = 1;
    92: op1_01_inv01 = 1;
    93: op1_01_inv01 = 1;
    94: op1_01_inv01 = 1;
    96: op1_01_inv01 = 1;
    default: op1_01_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in02 = reg_0503;
    5: op1_01_in02 = reg_0604;
    6: op1_01_in02 = reg_0652;
    7: op1_01_in02 = reg_0253;
    3: op1_01_in02 = imem07_in[75:72];
    49: op1_01_in02 = imem07_in[75:72];
    8: op1_01_in02 = imem00_in[75:72];
    2: op1_01_in02 = reg_0179;
    9: op1_01_in02 = reg_0310;
    10: op1_01_in02 = reg_0347;
    11: op1_01_in02 = reg_0682;
    21: op1_01_in02 = reg_0682;
    42: op1_01_in02 = reg_0682;
    12: op1_01_in02 = reg_0100;
    43: op1_01_in02 = reg_0100;
    1: op1_01_in02 = imem07_in[31:28];
    13: op1_01_in02 = reg_0031;
    14: op1_01_in02 = reg_0239;
    67: op1_01_in02 = reg_0239;
    15: op1_01_in02 = imem02_in[87:84];
    16: op1_01_in02 = imem05_in[39:36];
    17: op1_01_in02 = imem00_in[31:28];
    74: op1_01_in02 = imem00_in[31:28];
    18: op1_01_in02 = reg_0716;
    19: op1_01_in02 = imem00_in[87:84];
    28: op1_01_in02 = imem00_in[87:84];
    20: op1_01_in02 = reg_0278;
    41: op1_01_in02 = reg_0278;
    22: op1_01_in02 = imem02_in[35:32];
    23: op1_01_in02 = reg_0615;
    24: op1_01_in02 = imem03_in[63:60];
    25: op1_01_in02 = imem05_in[31:28];
    26: op1_01_in02 = reg_0102;
    27: op1_01_in02 = reg_0797;
    87: op1_01_in02 = reg_0797;
    29: op1_01_in02 = reg_0116;
    30: op1_01_in02 = reg_0490;
    54: op1_01_in02 = reg_0490;
    31: op1_01_in02 = imem00_in[103:100];
    85: op1_01_in02 = imem00_in[103:100];
    32: op1_01_in02 = reg_0242;
    33: op1_01_in02 = imem02_in[59:56];
    34: op1_01_in02 = imem00_in[83:80];
    36: op1_01_in02 = imem00_in[67:64];
    37: op1_01_in02 = imem02_in[111:108];
    38: op1_01_in02 = reg_0507;
    39: op1_01_in02 = reg_0517;
    40: op1_01_in02 = reg_0585;
    62: op1_01_in02 = reg_0585;
    44: op1_01_in02 = reg_0803;
    45: op1_01_in02 = reg_0231;
    46: op1_01_in02 = reg_0107;
    47: op1_01_in02 = reg_0740;
    48: op1_01_in02 = reg_0766;
    50: op1_01_in02 = reg_0218;
    79: op1_01_in02 = reg_0218;
    51: op1_01_in02 = imem04_in[71:68];
    52: op1_01_in02 = reg_0010;
    53: op1_01_in02 = imem05_in[11:8];
    55: op1_01_in02 = imem07_in[123:120];
    56: op1_01_in02 = imem00_in[79:76];
    88: op1_01_in02 = imem00_in[79:76];
    57: op1_01_in02 = imem00_in[55:52];
    81: op1_01_in02 = imem00_in[55:52];
    58: op1_01_in02 = imem07_in[15:12];
    59: op1_01_in02 = reg_0420;
    60: op1_01_in02 = imem00_in[71:68];
    61: op1_01_in02 = reg_0106;
    63: op1_01_in02 = imem06_in[127:124];
    64: op1_01_in02 = reg_0368;
    65: op1_01_in02 = imem07_in[91:88];
    66: op1_01_in02 = reg_0029;
    68: op1_01_in02 = reg_0493;
    69: op1_01_in02 = imem05_in[79:76];
    70: op1_01_in02 = imem00_in[27:24];
    71: op1_01_in02 = reg_0050;
    72: op1_01_in02 = reg_0720;
    82: op1_01_in02 = reg_0720;
    73: op1_01_in02 = reg_0438;
    75: op1_01_in02 = reg_0672;
    76: op1_01_in02 = reg_0306;
    77: op1_01_in02 = reg_0280;
    78: op1_01_in02 = imem07_in[83:80];
    80: op1_01_in02 = imem00_in[63:60];
    83: op1_01_in02 = reg_0806;
    84: op1_01_in02 = reg_0499;
    86: op1_01_in02 = reg_0512;
    89: op1_01_in02 = reg_0150;
    90: op1_01_in02 = imem07_in[3:0];
    91: op1_01_in02 = reg_0184;
    92: op1_01_in02 = reg_0009;
    93: op1_01_in02 = reg_0094;
    94: op1_01_in02 = reg_0094;
    95: op1_01_in02 = reg_0374;
    96: op1_01_in02 = reg_0019;
    default: op1_01_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv02 = 1;
    6: op1_01_inv02 = 1;
    7: op1_01_inv02 = 1;
    8: op1_01_inv02 = 1;
    10: op1_01_inv02 = 1;
    12: op1_01_inv02 = 1;
    1: op1_01_inv02 = 1;
    13: op1_01_inv02 = 1;
    14: op1_01_inv02 = 1;
    15: op1_01_inv02 = 1;
    16: op1_01_inv02 = 1;
    20: op1_01_inv02 = 1;
    21: op1_01_inv02 = 1;
    23: op1_01_inv02 = 1;
    24: op1_01_inv02 = 1;
    26: op1_01_inv02 = 1;
    27: op1_01_inv02 = 1;
    29: op1_01_inv02 = 1;
    31: op1_01_inv02 = 1;
    33: op1_01_inv02 = 1;
    36: op1_01_inv02 = 1;
    38: op1_01_inv02 = 1;
    39: op1_01_inv02 = 1;
    40: op1_01_inv02 = 1;
    49: op1_01_inv02 = 1;
    51: op1_01_inv02 = 1;
    52: op1_01_inv02 = 1;
    55: op1_01_inv02 = 1;
    56: op1_01_inv02 = 1;
    57: op1_01_inv02 = 1;
    59: op1_01_inv02 = 1;
    60: op1_01_inv02 = 1;
    61: op1_01_inv02 = 1;
    62: op1_01_inv02 = 1;
    64: op1_01_inv02 = 1;
    67: op1_01_inv02 = 1;
    70: op1_01_inv02 = 1;
    71: op1_01_inv02 = 1;
    74: op1_01_inv02 = 1;
    76: op1_01_inv02 = 1;
    78: op1_01_inv02 = 1;
    80: op1_01_inv02 = 1;
    81: op1_01_inv02 = 1;
    83: op1_01_inv02 = 1;
    84: op1_01_inv02 = 1;
    85: op1_01_inv02 = 1;
    87: op1_01_inv02 = 1;
    89: op1_01_inv02 = 1;
    91: op1_01_inv02 = 1;
    92: op1_01_inv02 = 1;
    96: op1_01_inv02 = 1;
    default: op1_01_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in03 = reg_0515;
    5: op1_01_in03 = reg_0617;
    6: op1_01_in03 = reg_0334;
    7: op1_01_in03 = reg_0132;
    3: op1_01_in03 = imem07_in[79:76];
    8: op1_01_in03 = imem00_in[79:76];
    2: op1_01_in03 = reg_0161;
    9: op1_01_in03 = reg_0342;
    10: op1_01_in03 = reg_0092;
    11: op1_01_in03 = reg_0689;
    12: op1_01_in03 = reg_0115;
    1: op1_01_in03 = imem07_in[39:36];
    13: op1_01_in03 = reg_0753;
    14: op1_01_in03 = reg_0217;
    15: op1_01_in03 = imem02_in[123:120];
    16: op1_01_in03 = imem05_in[55:52];
    25: op1_01_in03 = imem05_in[55:52];
    17: op1_01_in03 = imem00_in[51:48];
    18: op1_01_in03 = reg_0704;
    19: op1_01_in03 = imem00_in[127:124];
    20: op1_01_in03 = reg_0066;
    21: op1_01_in03 = reg_0693;
    22: op1_01_in03 = imem02_in[127:124];
    23: op1_01_in03 = reg_0344;
    24: op1_01_in03 = imem03_in[91:88];
    26: op1_01_in03 = reg_0117;
    27: op1_01_in03 = reg_0788;
    30: op1_01_in03 = reg_0788;
    28: op1_01_in03 = reg_0671;
    29: op1_01_in03 = reg_0104;
    96: op1_01_in03 = reg_0104;
    31: op1_01_in03 = imem00_in[111:108];
    32: op1_01_in03 = reg_0216;
    33: op1_01_in03 = imem02_in[115:112];
    37: op1_01_in03 = imem02_in[115:112];
    34: op1_01_in03 = imem00_in[99:96];
    36: op1_01_in03 = imem00_in[123:120];
    81: op1_01_in03 = imem00_in[123:120];
    38: op1_01_in03 = reg_0760;
    39: op1_01_in03 = reg_0811;
    40: op1_01_in03 = reg_0593;
    41: op1_01_in03 = reg_0318;
    42: op1_01_in03 = reg_0672;
    43: op1_01_in03 = reg_0101;
    44: op1_01_in03 = reg_0807;
    45: op1_01_in03 = reg_0029;
    46: op1_01_in03 = reg_0127;
    47: op1_01_in03 = imem03_in[59:56];
    48: op1_01_in03 = reg_0612;
    49: op1_01_in03 = imem07_in[87:84];
    58: op1_01_in03 = imem07_in[87:84];
    50: op1_01_in03 = reg_0605;
    51: op1_01_in03 = imem04_in[87:84];
    52: op1_01_in03 = imem04_in[3:0];
    53: op1_01_in03 = imem05_in[71:68];
    54: op1_01_in03 = reg_0484;
    55: op1_01_in03 = reg_0710;
    56: op1_01_in03 = imem00_in[83:80];
    88: op1_01_in03 = imem00_in[83:80];
    57: op1_01_in03 = imem00_in[63:60];
    59: op1_01_in03 = reg_0105;
    60: op1_01_in03 = imem00_in[87:84];
    61: op1_01_in03 = reg_0121;
    62: op1_01_in03 = reg_0622;
    63: op1_01_in03 = reg_0348;
    64: op1_01_in03 = imem07_in[23:20];
    65: op1_01_in03 = imem07_in[95:92];
    66: op1_01_in03 = imem07_in[51:48];
    67: op1_01_in03 = reg_0443;
    68: op1_01_in03 = reg_0596;
    69: op1_01_in03 = imem05_in[119:116];
    70: op1_01_in03 = imem00_in[67:64];
    71: op1_01_in03 = reg_0614;
    72: op1_01_in03 = reg_0721;
    73: op1_01_in03 = reg_0180;
    74: op1_01_in03 = imem00_in[35:32];
    75: op1_01_in03 = imem02_in[3:0];
    76: op1_01_in03 = reg_0511;
    77: op1_01_in03 = reg_0631;
    78: op1_01_in03 = imem07_in[99:96];
    79: op1_01_in03 = reg_0657;
    80: op1_01_in03 = reg_0492;
    82: op1_01_in03 = reg_0276;
    83: op1_01_in03 = reg_0009;
    84: op1_01_in03 = reg_0246;
    85: op1_01_in03 = reg_0758;
    86: op1_01_in03 = reg_0573;
    87: op1_01_in03 = reg_0245;
    89: op1_01_in03 = reg_0152;
    90: op1_01_in03 = imem07_in[15:12];
    92: op1_01_in03 = reg_0486;
    93: op1_01_in03 = imem03_in[39:36];
    94: op1_01_in03 = reg_0740;
    95: op1_01_in03 = reg_0587;
    default: op1_01_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_01_inv03 = 1;
    9: op1_01_inv03 = 1;
    12: op1_01_inv03 = 1;
    13: op1_01_inv03 = 1;
    15: op1_01_inv03 = 1;
    19: op1_01_inv03 = 1;
    21: op1_01_inv03 = 1;
    22: op1_01_inv03 = 1;
    23: op1_01_inv03 = 1;
    24: op1_01_inv03 = 1;
    26: op1_01_inv03 = 1;
    27: op1_01_inv03 = 1;
    28: op1_01_inv03 = 1;
    33: op1_01_inv03 = 1;
    37: op1_01_inv03 = 1;
    39: op1_01_inv03 = 1;
    40: op1_01_inv03 = 1;
    41: op1_01_inv03 = 1;
    44: op1_01_inv03 = 1;
    46: op1_01_inv03 = 1;
    50: op1_01_inv03 = 1;
    53: op1_01_inv03 = 1;
    56: op1_01_inv03 = 1;
    60: op1_01_inv03 = 1;
    61: op1_01_inv03 = 1;
    62: op1_01_inv03 = 1;
    63: op1_01_inv03 = 1;
    64: op1_01_inv03 = 1;
    67: op1_01_inv03 = 1;
    70: op1_01_inv03 = 1;
    71: op1_01_inv03 = 1;
    72: op1_01_inv03 = 1;
    73: op1_01_inv03 = 1;
    74: op1_01_inv03 = 1;
    75: op1_01_inv03 = 1;
    76: op1_01_inv03 = 1;
    77: op1_01_inv03 = 1;
    78: op1_01_inv03 = 1;
    81: op1_01_inv03 = 1;
    84: op1_01_inv03 = 1;
    85: op1_01_inv03 = 1;
    87: op1_01_inv03 = 1;
    95: op1_01_inv03 = 1;
    96: op1_01_inv03 = 1;
    default: op1_01_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in04 = reg_0498;
    5: op1_01_in04 = reg_0605;
    6: op1_01_in04 = reg_0357;
    7: op1_01_in04 = reg_0147;
    3: op1_01_in04 = imem07_in[83:80];
    8: op1_01_in04 = imem00_in[111:108];
    2: op1_01_in04 = reg_0169;
    9: op1_01_in04 = reg_0350;
    10: op1_01_in04 = reg_0045;
    11: op1_01_in04 = reg_0684;
    12: op1_01_in04 = reg_0113;
    46: op1_01_in04 = reg_0113;
    1: op1_01_in04 = imem07_in[63:60];
    13: op1_01_in04 = reg_0035;
    14: op1_01_in04 = reg_0242;
    15: op1_01_in04 = imem02_in[127:124];
    16: op1_01_in04 = imem05_in[63:60];
    17: op1_01_in04 = imem00_in[59:56];
    18: op1_01_in04 = reg_0702;
    19: op1_01_in04 = reg_0681;
    60: op1_01_in04 = reg_0681;
    20: op1_01_in04 = reg_0064;
    21: op1_01_in04 = reg_0683;
    22: op1_01_in04 = reg_0654;
    23: op1_01_in04 = reg_0372;
    24: op1_01_in04 = reg_0586;
    25: op1_01_in04 = imem05_in[119:116];
    26: op1_01_in04 = reg_0110;
    27: op1_01_in04 = reg_0795;
    54: op1_01_in04 = reg_0795;
    28: op1_01_in04 = reg_0678;
    59: op1_01_in04 = reg_0678;
    29: op1_01_in04 = reg_0115;
    63: op1_01_in04 = reg_0115;
    30: op1_01_in04 = reg_0785;
    31: op1_01_in04 = imem00_in[115:112];
    32: op1_01_in04 = reg_0247;
    33: op1_01_in04 = imem02_in[119:116];
    37: op1_01_in04 = imem02_in[119:116];
    34: op1_01_in04 = reg_0697;
    36: op1_01_in04 = reg_0695;
    38: op1_01_in04 = reg_0506;
    39: op1_01_in04 = imem04_in[43:40];
    40: op1_01_in04 = reg_0580;
    87: op1_01_in04 = reg_0580;
    41: op1_01_in04 = reg_0331;
    50: op1_01_in04 = reg_0331;
    42: op1_01_in04 = reg_0679;
    43: op1_01_in04 = reg_0117;
    44: op1_01_in04 = reg_0010;
    45: op1_01_in04 = reg_0367;
    47: op1_01_in04 = imem03_in[67:64];
    48: op1_01_in04 = reg_0402;
    49: op1_01_in04 = reg_0717;
    51: op1_01_in04 = imem04_in[91:88];
    52: op1_01_in04 = imem04_in[11:8];
    53: op1_01_in04 = imem05_in[87:84];
    55: op1_01_in04 = reg_0729;
    56: op1_01_in04 = imem00_in[91:88];
    88: op1_01_in04 = imem00_in[91:88];
    57: op1_01_in04 = imem00_in[71:68];
    70: op1_01_in04 = imem00_in[71:68];
    58: op1_01_in04 = reg_0728;
    61: op1_01_in04 = reg_0126;
    62: op1_01_in04 = reg_0068;
    64: op1_01_in04 = imem07_in[119:116];
    78: op1_01_in04 = imem07_in[119:116];
    65: op1_01_in04 = imem07_in[107:104];
    66: op1_01_in04 = imem07_in[59:56];
    67: op1_01_in04 = reg_0174;
    68: op1_01_in04 = reg_0319;
    69: op1_01_in04 = reg_0392;
    71: op1_01_in04 = reg_0078;
    72: op1_01_in04 = reg_0723;
    73: op1_01_in04 = reg_0162;
    74: op1_01_in04 = imem00_in[39:36];
    75: op1_01_in04 = imem02_in[23:20];
    76: op1_01_in04 = reg_0675;
    77: op1_01_in04 = reg_0629;
    79: op1_01_in04 = reg_0664;
    80: op1_01_in04 = reg_0689;
    81: op1_01_in04 = reg_0693;
    82: op1_01_in04 = reg_0277;
    83: op1_01_in04 = imem04_in[3:0];
    84: op1_01_in04 = reg_0278;
    85: op1_01_in04 = reg_0407;
    86: op1_01_in04 = reg_0029;
    89: op1_01_in04 = imem06_in[7:4];
    90: op1_01_in04 = imem07_in[19:16];
    92: op1_01_in04 = reg_0389;
    93: op1_01_in04 = imem03_in[43:40];
    94: op1_01_in04 = imem03_in[11:8];
    95: op1_01_in04 = reg_0581;
    96: op1_01_in04 = reg_0119;
    default: op1_01_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv04 = 1;
    2: op1_01_inv04 = 1;
    11: op1_01_inv04 = 1;
    12: op1_01_inv04 = 1;
    1: op1_01_inv04 = 1;
    13: op1_01_inv04 = 1;
    15: op1_01_inv04 = 1;
    17: op1_01_inv04 = 1;
    18: op1_01_inv04 = 1;
    19: op1_01_inv04 = 1;
    22: op1_01_inv04 = 1;
    25: op1_01_inv04 = 1;
    27: op1_01_inv04 = 1;
    30: op1_01_inv04 = 1;
    34: op1_01_inv04 = 1;
    39: op1_01_inv04 = 1;
    40: op1_01_inv04 = 1;
    42: op1_01_inv04 = 1;
    43: op1_01_inv04 = 1;
    44: op1_01_inv04 = 1;
    47: op1_01_inv04 = 1;
    48: op1_01_inv04 = 1;
    49: op1_01_inv04 = 1;
    50: op1_01_inv04 = 1;
    53: op1_01_inv04 = 1;
    54: op1_01_inv04 = 1;
    57: op1_01_inv04 = 1;
    58: op1_01_inv04 = 1;
    59: op1_01_inv04 = 1;
    63: op1_01_inv04 = 1;
    64: op1_01_inv04 = 1;
    65: op1_01_inv04 = 1;
    66: op1_01_inv04 = 1;
    69: op1_01_inv04 = 1;
    72: op1_01_inv04 = 1;
    74: op1_01_inv04 = 1;
    75: op1_01_inv04 = 1;
    77: op1_01_inv04 = 1;
    78: op1_01_inv04 = 1;
    79: op1_01_inv04 = 1;
    85: op1_01_inv04 = 1;
    89: op1_01_inv04 = 1;
    90: op1_01_inv04 = 1;
    92: op1_01_inv04 = 1;
    94: op1_01_inv04 = 1;
    95: op1_01_inv04 = 1;
    96: op1_01_inv04 = 1;
    default: op1_01_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in05 = reg_0232;
    5: op1_01_in05 = reg_0626;
    6: op1_01_in05 = reg_0346;
    7: op1_01_in05 = reg_0149;
    3: op1_01_in05 = imem07_in[119:116];
    8: op1_01_in05 = imem00_in[115:112];
    2: op1_01_in05 = reg_0183;
    9: op1_01_in05 = reg_0081;
    10: op1_01_in05 = reg_0087;
    11: op1_01_in05 = reg_0686;
    12: op1_01_in05 = reg_0121;
    43: op1_01_in05 = reg_0121;
    13: op1_01_in05 = reg_0750;
    14: op1_01_in05 = reg_0503;
    15: op1_01_in05 = reg_0658;
    16: op1_01_in05 = imem05_in[83:80];
    17: op1_01_in05 = imem00_in[95:92];
    88: op1_01_in05 = imem00_in[95:92];
    18: op1_01_in05 = reg_0708;
    19: op1_01_in05 = reg_0696;
    20: op1_01_in05 = reg_0256;
    21: op1_01_in05 = reg_0685;
    36: op1_01_in05 = reg_0685;
    22: op1_01_in05 = reg_0640;
    23: op1_01_in05 = reg_0337;
    24: op1_01_in05 = reg_0587;
    25: op1_01_in05 = reg_0798;
    26: op1_01_in05 = imem02_in[15:12];
    27: op1_01_in05 = reg_0793;
    28: op1_01_in05 = reg_0675;
    29: op1_01_in05 = reg_0107;
    30: op1_01_in05 = reg_0794;
    31: op1_01_in05 = reg_0693;
    32: op1_01_in05 = reg_0236;
    33: op1_01_in05 = imem02_in[123:120];
    34: op1_01_in05 = reg_0676;
    37: op1_01_in05 = reg_0645;
    38: op1_01_in05 = reg_0244;
    39: op1_01_in05 = imem04_in[47:44];
    40: op1_01_in05 = reg_0597;
    41: op1_01_in05 = reg_0370;
    42: op1_01_in05 = reg_0691;
    44: op1_01_in05 = reg_0809;
    45: op1_01_in05 = imem07_in[23:20];
    46: op1_01_in05 = imem02_in[7:4];
    47: op1_01_in05 = imem03_in[91:88];
    48: op1_01_in05 = reg_0774;
    71: op1_01_in05 = reg_0774;
    49: op1_01_in05 = reg_0718;
    50: op1_01_in05 = reg_0577;
    51: op1_01_in05 = imem04_in[123:120];
    52: op1_01_in05 = imem04_in[31:28];
    53: op1_01_in05 = imem05_in[103:100];
    54: op1_01_in05 = reg_0489;
    55: op1_01_in05 = reg_0705;
    56: op1_01_in05 = imem00_in[107:104];
    57: op1_01_in05 = imem00_in[107:104];
    58: op1_01_in05 = reg_0720;
    59: op1_01_in05 = imem02_in[27:24];
    60: op1_01_in05 = reg_0749;
    61: op1_01_in05 = imem02_in[19:16];
    62: op1_01_in05 = reg_0233;
    63: op1_01_in05 = reg_0238;
    64: op1_01_in05 = imem07_in[123:120];
    65: op1_01_in05 = imem07_in[127:124];
    78: op1_01_in05 = imem07_in[127:124];
    66: op1_01_in05 = imem07_in[99:96];
    67: op1_01_in05 = reg_0175;
    68: op1_01_in05 = reg_0318;
    69: op1_01_in05 = reg_0326;
    70: op1_01_in05 = imem00_in[99:96];
    72: op1_01_in05 = reg_0714;
    73: op1_01_in05 = reg_0167;
    74: op1_01_in05 = imem00_in[71:68];
    75: op1_01_in05 = imem02_in[103:100];
    76: op1_01_in05 = reg_0106;
    77: op1_01_in05 = reg_0679;
    79: op1_01_in05 = reg_0632;
    80: op1_01_in05 = reg_0478;
    81: op1_01_in05 = reg_0690;
    82: op1_01_in05 = reg_0389;
    83: op1_01_in05 = imem04_in[19:16];
    84: op1_01_in05 = reg_0307;
    85: op1_01_in05 = reg_0634;
    86: op1_01_in05 = reg_0663;
    87: op1_01_in05 = reg_0399;
    89: op1_01_in05 = imem06_in[23:20];
    90: op1_01_in05 = imem07_in[27:24];
    92: op1_01_in05 = reg_0575;
    93: op1_01_in05 = imem03_in[47:44];
    94: op1_01_in05 = imem03_in[39:36];
    95: op1_01_in05 = reg_0594;
    96: op1_01_in05 = reg_0115;
    default: op1_01_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_01_inv05 = 1;
    13: op1_01_inv05 = 1;
    15: op1_01_inv05 = 1;
    17: op1_01_inv05 = 1;
    18: op1_01_inv05 = 1;
    20: op1_01_inv05 = 1;
    24: op1_01_inv05 = 1;
    26: op1_01_inv05 = 1;
    27: op1_01_inv05 = 1;
    28: op1_01_inv05 = 1;
    29: op1_01_inv05 = 1;
    30: op1_01_inv05 = 1;
    33: op1_01_inv05 = 1;
    34: op1_01_inv05 = 1;
    36: op1_01_inv05 = 1;
    37: op1_01_inv05 = 1;
    38: op1_01_inv05 = 1;
    39: op1_01_inv05 = 1;
    40: op1_01_inv05 = 1;
    42: op1_01_inv05 = 1;
    44: op1_01_inv05 = 1;
    45: op1_01_inv05 = 1;
    46: op1_01_inv05 = 1;
    47: op1_01_inv05 = 1;
    48: op1_01_inv05 = 1;
    49: op1_01_inv05 = 1;
    55: op1_01_inv05 = 1;
    57: op1_01_inv05 = 1;
    60: op1_01_inv05 = 1;
    66: op1_01_inv05 = 1;
    67: op1_01_inv05 = 1;
    68: op1_01_inv05 = 1;
    69: op1_01_inv05 = 1;
    71: op1_01_inv05 = 1;
    72: op1_01_inv05 = 1;
    74: op1_01_inv05 = 1;
    75: op1_01_inv05 = 1;
    79: op1_01_inv05 = 1;
    81: op1_01_inv05 = 1;
    82: op1_01_inv05 = 1;
    84: op1_01_inv05 = 1;
    86: op1_01_inv05 = 1;
    88: op1_01_inv05 = 1;
    89: op1_01_inv05 = 1;
    90: op1_01_inv05 = 1;
    92: op1_01_inv05 = 1;
    95: op1_01_inv05 = 1;
    96: op1_01_inv05 = 1;
    default: op1_01_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in06 = reg_0226;
    5: op1_01_in06 = reg_0627;
    6: op1_01_in06 = reg_0324;
    7: op1_01_in06 = reg_0153;
    3: op1_01_in06 = imem07_in[123:120];
    8: op1_01_in06 = reg_0682;
    2: op1_01_in06 = reg_0178;
    9: op1_01_in06 = reg_0095;
    10: op1_01_in06 = reg_0093;
    11: op1_01_in06 = reg_0679;
    12: op1_01_in06 = imem02_in[23:20];
    13: op1_01_in06 = imem07_in[3:0];
    14: op1_01_in06 = reg_0236;
    15: op1_01_in06 = reg_0358;
    16: op1_01_in06 = imem05_in[95:92];
    17: op1_01_in06 = imem00_in[127:124];
    70: op1_01_in06 = imem00_in[127:124];
    18: op1_01_in06 = reg_0715;
    19: op1_01_in06 = reg_0688;
    42: op1_01_in06 = reg_0688;
    81: op1_01_in06 = reg_0688;
    20: op1_01_in06 = imem05_in[7:4];
    21: op1_01_in06 = reg_0684;
    22: op1_01_in06 = reg_0641;
    23: op1_01_in06 = reg_0033;
    24: op1_01_in06 = reg_0592;
    25: op1_01_in06 = reg_0488;
    26: op1_01_in06 = imem02_in[43:40];
    27: op1_01_in06 = reg_0785;
    28: op1_01_in06 = reg_0692;
    29: op1_01_in06 = reg_0126;
    30: op1_01_in06 = reg_0790;
    31: op1_01_in06 = reg_0697;
    32: op1_01_in06 = reg_0248;
    33: op1_01_in06 = reg_0637;
    34: op1_01_in06 = reg_0698;
    36: op1_01_in06 = reg_0677;
    37: op1_01_in06 = reg_0658;
    38: op1_01_in06 = reg_0216;
    39: op1_01_in06 = imem04_in[55:52];
    40: op1_01_in06 = reg_0394;
    41: op1_01_in06 = reg_0762;
    43: op1_01_in06 = imem02_in[7:4];
    44: op1_01_in06 = imem04_in[35:32];
    45: op1_01_in06 = imem07_in[43:40];
    46: op1_01_in06 = imem02_in[55:52];
    47: op1_01_in06 = imem03_in[127:124];
    48: op1_01_in06 = reg_0317;
    49: op1_01_in06 = reg_0711;
    50: op1_01_in06 = reg_0775;
    51: op1_01_in06 = reg_0316;
    52: op1_01_in06 = imem04_in[47:44];
    53: op1_01_in06 = imem05_in[127:124];
    54: op1_01_in06 = reg_0309;
    55: op1_01_in06 = reg_0713;
    56: op1_01_in06 = imem00_in[115:112];
    57: op1_01_in06 = reg_0689;
    58: op1_01_in06 = reg_0731;
    59: op1_01_in06 = imem02_in[87:84];
    60: op1_01_in06 = reg_0463;
    61: op1_01_in06 = imem02_in[47:44];
    62: op1_01_in06 = imem05_in[27:24];
    63: op1_01_in06 = reg_0405;
    64: op1_01_in06 = reg_0704;
    65: op1_01_in06 = reg_0730;
    66: op1_01_in06 = imem07_in[103:100];
    67: op1_01_in06 = reg_0163;
    68: op1_01_in06 = reg_0751;
    69: op1_01_in06 = reg_0257;
    71: op1_01_in06 = imem05_in[63:60];
    72: op1_01_in06 = reg_0718;
    73: op1_01_in06 = reg_0169;
    74: op1_01_in06 = reg_0693;
    75: op1_01_in06 = imem02_in[107:104];
    76: op1_01_in06 = imem02_in[3:0];
    77: op1_01_in06 = reg_0223;
    78: op1_01_in06 = reg_0051;
    79: op1_01_in06 = imem07_in[39:36];
    80: op1_01_in06 = reg_0214;
    82: op1_01_in06 = reg_0812;
    83: op1_01_in06 = imem04_in[43:40];
    84: op1_01_in06 = reg_0719;
    85: op1_01_in06 = reg_0455;
    86: op1_01_in06 = reg_0620;
    87: op1_01_in06 = reg_0277;
    88: op1_01_in06 = imem00_in[119:116];
    89: op1_01_in06 = imem06_in[43:40];
    90: op1_01_in06 = imem07_in[59:56];
    92: op1_01_in06 = reg_0568;
    93: op1_01_in06 = imem03_in[67:64];
    94: op1_01_in06 = imem03_in[91:88];
    95: op1_01_in06 = reg_0566;
    96: op1_01_in06 = reg_0574;
    default: op1_01_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv06 = 1;
    6: op1_01_inv06 = 1;
    7: op1_01_inv06 = 1;
    3: op1_01_inv06 = 1;
    8: op1_01_inv06 = 1;
    2: op1_01_inv06 = 1;
    12: op1_01_inv06 = 1;
    13: op1_01_inv06 = 1;
    18: op1_01_inv06 = 1;
    22: op1_01_inv06 = 1;
    25: op1_01_inv06 = 1;
    27: op1_01_inv06 = 1;
    30: op1_01_inv06 = 1;
    31: op1_01_inv06 = 1;
    37: op1_01_inv06 = 1;
    38: op1_01_inv06 = 1;
    40: op1_01_inv06 = 1;
    44: op1_01_inv06 = 1;
    49: op1_01_inv06 = 1;
    50: op1_01_inv06 = 1;
    51: op1_01_inv06 = 1;
    52: op1_01_inv06 = 1;
    53: op1_01_inv06 = 1;
    54: op1_01_inv06 = 1;
    56: op1_01_inv06 = 1;
    60: op1_01_inv06 = 1;
    61: op1_01_inv06 = 1;
    62: op1_01_inv06 = 1;
    63: op1_01_inv06 = 1;
    64: op1_01_inv06 = 1;
    65: op1_01_inv06 = 1;
    67: op1_01_inv06 = 1;
    71: op1_01_inv06 = 1;
    72: op1_01_inv06 = 1;
    74: op1_01_inv06 = 1;
    76: op1_01_inv06 = 1;
    78: op1_01_inv06 = 1;
    80: op1_01_inv06 = 1;
    82: op1_01_inv06 = 1;
    83: op1_01_inv06 = 1;
    85: op1_01_inv06 = 1;
    87: op1_01_inv06 = 1;
    88: op1_01_inv06 = 1;
    92: op1_01_inv06 = 1;
    93: op1_01_inv06 = 1;
    94: op1_01_inv06 = 1;
    default: op1_01_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in07 = reg_0233;
    5: op1_01_in07 = reg_0348;
    6: op1_01_in07 = reg_0342;
    7: op1_01_in07 = reg_0140;
    3: op1_01_in07 = reg_0425;
    8: op1_01_in07 = reg_0693;
    2: op1_01_in07 = reg_0157;
    9: op1_01_in07 = reg_0060;
    10: op1_01_in07 = reg_0073;
    11: op1_01_in07 = reg_0677;
    12: op1_01_in07 = imem02_in[39:36];
    13: op1_01_in07 = imem07_in[15:12];
    14: op1_01_in07 = reg_0245;
    15: op1_01_in07 = reg_0364;
    16: op1_01_in07 = reg_0798;
    17: op1_01_in07 = reg_0698;
    18: op1_01_in07 = reg_0701;
    19: op1_01_in07 = reg_0692;
    20: op1_01_in07 = imem05_in[19:16];
    21: op1_01_in07 = reg_0690;
    22: op1_01_in07 = reg_0320;
    23: op1_01_in07 = reg_0032;
    24: op1_01_in07 = reg_0585;
    25: op1_01_in07 = reg_0793;
    26: op1_01_in07 = imem02_in[107:104];
    27: op1_01_in07 = reg_0091;
    28: op1_01_in07 = reg_0465;
    57: op1_01_in07 = reg_0465;
    29: op1_01_in07 = imem02_in[11:8];
    30: op1_01_in07 = reg_0787;
    31: op1_01_in07 = reg_0674;
    32: op1_01_in07 = reg_0243;
    33: op1_01_in07 = reg_0660;
    34: op1_01_in07 = reg_0679;
    36: op1_01_in07 = reg_0450;
    37: op1_01_in07 = reg_0656;
    38: op1_01_in07 = reg_0234;
    39: op1_01_in07 = imem04_in[71:68];
    40: op1_01_in07 = reg_0561;
    41: op1_01_in07 = reg_0405;
    42: op1_01_in07 = reg_0453;
    60: op1_01_in07 = reg_0453;
    43: op1_01_in07 = imem02_in[23:20];
    44: op1_01_in07 = imem04_in[87:84];
    45: op1_01_in07 = imem07_in[47:44];
    46: op1_01_in07 = imem02_in[99:96];
    47: op1_01_in07 = reg_0602;
    48: op1_01_in07 = reg_0577;
    49: op1_01_in07 = reg_0706;
    50: op1_01_in07 = reg_0773;
    51: op1_01_in07 = reg_0552;
    52: op1_01_in07 = imem04_in[107:104];
    53: op1_01_in07 = reg_0483;
    54: op1_01_in07 = reg_0249;
    69: op1_01_in07 = reg_0249;
    55: op1_01_in07 = reg_0266;
    56: op1_01_in07 = reg_0695;
    88: op1_01_in07 = reg_0695;
    58: op1_01_in07 = reg_0721;
    59: op1_01_in07 = imem02_in[119:116];
    61: op1_01_in07 = imem02_in[91:88];
    62: op1_01_in07 = imem05_in[47:44];
    63: op1_01_in07 = reg_0515;
    64: op1_01_in07 = reg_0719;
    65: op1_01_in07 = reg_0723;
    66: op1_01_in07 = imem07_in[115:112];
    67: op1_01_in07 = reg_0176;
    68: op1_01_in07 = reg_0387;
    70: op1_01_in07 = reg_0683;
    71: op1_01_in07 = imem05_in[67:64];
    72: op1_01_in07 = reg_0727;
    73: op1_01_in07 = reg_0166;
    74: op1_01_in07 = reg_0612;
    75: op1_01_in07 = reg_0534;
    76: op1_01_in07 = imem02_in[15:12];
    77: op1_01_in07 = reg_0301;
    78: op1_01_in07 = reg_0434;
    79: op1_01_in07 = imem07_in[79:76];
    80: op1_01_in07 = reg_0191;
    81: op1_01_in07 = reg_0247;
    82: op1_01_in07 = reg_0829;
    83: op1_01_in07 = imem04_in[51:48];
    84: op1_01_in07 = reg_0389;
    85: op1_01_in07 = reg_0481;
    86: op1_01_in07 = reg_0794;
    87: op1_01_in07 = reg_0812;
    89: op1_01_in07 = imem06_in[71:68];
    90: op1_01_in07 = imem07_in[67:64];
    92: op1_01_in07 = reg_0569;
    93: op1_01_in07 = imem03_in[75:72];
    94: op1_01_in07 = imem03_in[99:96];
    95: op1_01_in07 = reg_0584;
    96: op1_01_in07 = reg_0054;
    default: op1_01_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv07 = 1;
    5: op1_01_inv07 = 1;
    3: op1_01_inv07 = 1;
    9: op1_01_inv07 = 1;
    12: op1_01_inv07 = 1;
    15: op1_01_inv07 = 1;
    16: op1_01_inv07 = 1;
    17: op1_01_inv07 = 1;
    18: op1_01_inv07 = 1;
    23: op1_01_inv07 = 1;
    24: op1_01_inv07 = 1;
    28: op1_01_inv07 = 1;
    31: op1_01_inv07 = 1;
    34: op1_01_inv07 = 1;
    36: op1_01_inv07 = 1;
    37: op1_01_inv07 = 1;
    41: op1_01_inv07 = 1;
    42: op1_01_inv07 = 1;
    43: op1_01_inv07 = 1;
    44: op1_01_inv07 = 1;
    49: op1_01_inv07 = 1;
    50: op1_01_inv07 = 1;
    51: op1_01_inv07 = 1;
    52: op1_01_inv07 = 1;
    53: op1_01_inv07 = 1;
    54: op1_01_inv07 = 1;
    56: op1_01_inv07 = 1;
    58: op1_01_inv07 = 1;
    65: op1_01_inv07 = 1;
    66: op1_01_inv07 = 1;
    68: op1_01_inv07 = 1;
    70: op1_01_inv07 = 1;
    71: op1_01_inv07 = 1;
    72: op1_01_inv07 = 1;
    73: op1_01_inv07 = 1;
    75: op1_01_inv07 = 1;
    77: op1_01_inv07 = 1;
    78: op1_01_inv07 = 1;
    79: op1_01_inv07 = 1;
    80: op1_01_inv07 = 1;
    81: op1_01_inv07 = 1;
    82: op1_01_inv07 = 1;
    84: op1_01_inv07 = 1;
    90: op1_01_inv07 = 1;
    93: op1_01_inv07 = 1;
    96: op1_01_inv07 = 1;
    default: op1_01_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in08 = reg_0218;
    5: op1_01_in08 = reg_0386;
    6: op1_01_in08 = reg_0338;
    7: op1_01_in08 = imem06_in[7:4];
    3: op1_01_in08 = reg_0418;
    8: op1_01_in08 = reg_0697;
    2: op1_01_in08 = reg_0171;
    9: op1_01_in08 = reg_0094;
    10: op1_01_in08 = imem03_in[31:28];
    11: op1_01_in08 = reg_0688;
    12: op1_01_in08 = imem02_in[51:48];
    13: op1_01_in08 = imem07_in[23:20];
    14: op1_01_in08 = reg_0219;
    15: op1_01_in08 = reg_0324;
    16: op1_01_in08 = reg_0483;
    17: op1_01_in08 = reg_0670;
    18: op1_01_in08 = reg_0441;
    19: op1_01_in08 = reg_0669;
    20: op1_01_in08 = imem05_in[31:28];
    21: op1_01_in08 = reg_0677;
    22: op1_01_in08 = reg_0326;
    23: op1_01_in08 = reg_0034;
    24: op1_01_in08 = reg_0570;
    25: op1_01_in08 = reg_0784;
    26: op1_01_in08 = imem02_in[119:116];
    27: op1_01_in08 = reg_0304;
    28: op1_01_in08 = reg_0451;
    29: op1_01_in08 = imem02_in[43:40];
    43: op1_01_in08 = imem02_in[43:40];
    30: op1_01_in08 = reg_0091;
    31: op1_01_in08 = reg_0678;
    32: op1_01_in08 = reg_0108;
    33: op1_01_in08 = reg_0647;
    37: op1_01_in08 = reg_0647;
    34: op1_01_in08 = reg_0680;
    36: op1_01_in08 = reg_0462;
    38: op1_01_in08 = reg_0122;
    39: op1_01_in08 = reg_0315;
    40: op1_01_in08 = reg_0564;
    41: op1_01_in08 = reg_0401;
    42: op1_01_in08 = reg_0454;
    44: op1_01_in08 = imem04_in[95:92];
    45: op1_01_in08 = imem07_in[75:72];
    46: op1_01_in08 = imem02_in[107:104];
    47: op1_01_in08 = reg_0565;
    48: op1_01_in08 = reg_0777;
    49: op1_01_in08 = reg_0636;
    50: op1_01_in08 = reg_0406;
    51: op1_01_in08 = reg_0087;
    52: op1_01_in08 = imem04_in[123:120];
    53: op1_01_in08 = reg_0488;
    54: op1_01_in08 = reg_0307;
    55: op1_01_in08 = reg_0295;
    56: op1_01_in08 = reg_0492;
    57: op1_01_in08 = reg_0476;
    58: op1_01_in08 = reg_0714;
    59: op1_01_in08 = imem02_in[123:120];
    60: op1_01_in08 = reg_0457;
    61: op1_01_in08 = imem02_in[115:112];
    62: op1_01_in08 = imem05_in[79:76];
    63: op1_01_in08 = reg_0028;
    64: op1_01_in08 = reg_0730;
    65: op1_01_in08 = reg_0712;
    66: op1_01_in08 = reg_0722;
    67: op1_01_in08 = reg_0158;
    68: op1_01_in08 = reg_0571;
    69: op1_01_in08 = reg_0383;
    70: op1_01_in08 = reg_0407;
    71: op1_01_in08 = reg_0231;
    72: op1_01_in08 = reg_0447;
    73: op1_01_in08 = reg_0164;
    74: op1_01_in08 = reg_0749;
    75: op1_01_in08 = reg_0427;
    76: op1_01_in08 = imem02_in[75:72];
    77: op1_01_in08 = reg_0416;
    78: op1_01_in08 = reg_0444;
    79: op1_01_in08 = imem07_in[115:112];
    80: op1_01_in08 = reg_0212;
    81: op1_01_in08 = reg_0699;
    82: op1_01_in08 = reg_0783;
    83: op1_01_in08 = imem04_in[67:64];
    84: op1_01_in08 = reg_0285;
    85: op1_01_in08 = reg_0471;
    86: op1_01_in08 = reg_0651;
    87: op1_01_in08 = reg_0147;
    88: op1_01_in08 = reg_0463;
    89: op1_01_in08 = imem06_in[95:92];
    90: op1_01_in08 = imem07_in[83:80];
    92: op1_01_in08 = reg_0398;
    93: op1_01_in08 = imem03_in[83:80];
    94: op1_01_in08 = imem03_in[107:104];
    95: op1_01_in08 = reg_0096;
    96: op1_01_in08 = reg_0567;
    default: op1_01_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv08 = 1;
    9: op1_01_inv08 = 1;
    14: op1_01_inv08 = 1;
    21: op1_01_inv08 = 1;
    24: op1_01_inv08 = 1;
    25: op1_01_inv08 = 1;
    28: op1_01_inv08 = 1;
    31: op1_01_inv08 = 1;
    32: op1_01_inv08 = 1;
    39: op1_01_inv08 = 1;
    40: op1_01_inv08 = 1;
    43: op1_01_inv08 = 1;
    47: op1_01_inv08 = 1;
    48: op1_01_inv08 = 1;
    51: op1_01_inv08 = 1;
    53: op1_01_inv08 = 1;
    55: op1_01_inv08 = 1;
    58: op1_01_inv08 = 1;
    65: op1_01_inv08 = 1;
    67: op1_01_inv08 = 1;
    68: op1_01_inv08 = 1;
    70: op1_01_inv08 = 1;
    74: op1_01_inv08 = 1;
    77: op1_01_inv08 = 1;
    78: op1_01_inv08 = 1;
    79: op1_01_inv08 = 1;
    81: op1_01_inv08 = 1;
    84: op1_01_inv08 = 1;
    88: op1_01_inv08 = 1;
    90: op1_01_inv08 = 1;
    93: op1_01_inv08 = 1;
    96: op1_01_inv08 = 1;
    default: op1_01_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in09 = reg_0234;
    5: op1_01_in09 = reg_0033;
    6: op1_01_in09 = reg_0355;
    7: op1_01_in09 = imem06_in[15:12];
    3: op1_01_in09 = reg_0428;
    8: op1_01_in09 = reg_0698;
    9: op1_01_in09 = imem03_in[15:12];
    10: op1_01_in09 = imem03_in[59:56];
    11: op1_01_in09 = reg_0463;
    12: op1_01_in09 = imem02_in[107:104];
    13: op1_01_in09 = imem07_in[43:40];
    14: op1_01_in09 = reg_0249;
    15: op1_01_in09 = reg_0338;
    16: op1_01_in09 = reg_0795;
    17: op1_01_in09 = reg_0679;
    18: op1_01_in09 = reg_0446;
    19: op1_01_in09 = reg_0454;
    20: op1_01_in09 = imem05_in[63:60];
    21: op1_01_in09 = reg_0674;
    22: op1_01_in09 = reg_0359;
    23: op1_01_in09 = reg_0749;
    56: op1_01_in09 = reg_0749;
    24: op1_01_in09 = reg_0360;
    25: op1_01_in09 = reg_0309;
    27: op1_01_in09 = reg_0309;
    26: op1_01_in09 = reg_0661;
    28: op1_01_in09 = reg_0472;
    29: op1_01_in09 = imem02_in[59:56];
    30: op1_01_in09 = reg_0741;
    31: op1_01_in09 = reg_0688;
    32: op1_01_in09 = imem02_in[23:20];
    33: op1_01_in09 = reg_0659;
    34: op1_01_in09 = reg_0450;
    36: op1_01_in09 = reg_0481;
    37: op1_01_in09 = reg_0640;
    38: op1_01_in09 = reg_0116;
    39: op1_01_in09 = reg_0087;
    40: op1_01_in09 = reg_0388;
    41: op1_01_in09 = reg_0375;
    42: op1_01_in09 = reg_0451;
    43: op1_01_in09 = imem02_in[47:44];
    44: op1_01_in09 = imem04_in[115:112];
    45: op1_01_in09 = imem07_in[115:112];
    46: op1_01_in09 = reg_0337;
    59: op1_01_in09 = reg_0337;
    47: op1_01_in09 = reg_0600;
    48: op1_01_in09 = reg_0040;
    49: op1_01_in09 = reg_0174;
    50: op1_01_in09 = reg_0401;
    51: op1_01_in09 = reg_0060;
    52: op1_01_in09 = reg_0315;
    95: op1_01_in09 = reg_0315;
    53: op1_01_in09 = reg_0788;
    54: op1_01_in09 = reg_0277;
    55: op1_01_in09 = reg_0635;
    57: op1_01_in09 = reg_0462;
    58: op1_01_in09 = reg_0729;
    60: op1_01_in09 = reg_0458;
    61: op1_01_in09 = reg_0655;
    62: op1_01_in09 = imem05_in[107:104];
    63: op1_01_in09 = reg_0813;
    64: op1_01_in09 = reg_0710;
    65: op1_01_in09 = reg_0707;
    66: op1_01_in09 = reg_0719;
    68: op1_01_in09 = reg_0811;
    69: op1_01_in09 = reg_0145;
    70: op1_01_in09 = reg_0680;
    71: op1_01_in09 = reg_0742;
    72: op1_01_in09 = reg_0239;
    73: op1_01_in09 = reg_0157;
    74: op1_01_in09 = reg_0658;
    75: op1_01_in09 = reg_0352;
    76: op1_01_in09 = imem02_in[127:124];
    77: op1_01_in09 = imem05_in[7:4];
    78: op1_01_in09 = reg_0437;
    79: op1_01_in09 = reg_0722;
    80: op1_01_in09 = reg_0199;
    81: op1_01_in09 = reg_0453;
    82: op1_01_in09 = imem06_in[3:0];
    83: op1_01_in09 = imem04_in[79:76];
    84: op1_01_in09 = reg_0827;
    85: op1_01_in09 = reg_0468;
    86: op1_01_in09 = reg_0652;
    87: op1_01_in09 = reg_0781;
    88: op1_01_in09 = reg_0475;
    89: op1_01_in09 = reg_0409;
    90: op1_01_in09 = imem07_in[87:84];
    92: op1_01_in09 = reg_0733;
    93: op1_01_in09 = reg_0602;
    94: op1_01_in09 = imem03_in[123:120];
    96: op1_01_in09 = reg_0240;
    default: op1_01_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv09 = 1;
    5: op1_01_inv09 = 1;
    6: op1_01_inv09 = 1;
    7: op1_01_inv09 = 1;
    3: op1_01_inv09 = 1;
    11: op1_01_inv09 = 1;
    12: op1_01_inv09 = 1;
    14: op1_01_inv09 = 1;
    15: op1_01_inv09 = 1;
    17: op1_01_inv09 = 1;
    18: op1_01_inv09 = 1;
    22: op1_01_inv09 = 1;
    23: op1_01_inv09 = 1;
    27: op1_01_inv09 = 1;
    29: op1_01_inv09 = 1;
    30: op1_01_inv09 = 1;
    36: op1_01_inv09 = 1;
    37: op1_01_inv09 = 1;
    38: op1_01_inv09 = 1;
    39: op1_01_inv09 = 1;
    42: op1_01_inv09 = 1;
    43: op1_01_inv09 = 1;
    44: op1_01_inv09 = 1;
    46: op1_01_inv09 = 1;
    49: op1_01_inv09 = 1;
    51: op1_01_inv09 = 1;
    52: op1_01_inv09 = 1;
    55: op1_01_inv09 = 1;
    56: op1_01_inv09 = 1;
    57: op1_01_inv09 = 1;
    58: op1_01_inv09 = 1;
    59: op1_01_inv09 = 1;
    60: op1_01_inv09 = 1;
    65: op1_01_inv09 = 1;
    69: op1_01_inv09 = 1;
    71: op1_01_inv09 = 1;
    74: op1_01_inv09 = 1;
    75: op1_01_inv09 = 1;
    76: op1_01_inv09 = 1;
    82: op1_01_inv09 = 1;
    83: op1_01_inv09 = 1;
    88: op1_01_inv09 = 1;
    89: op1_01_inv09 = 1;
    default: op1_01_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in10 = reg_0219;
    5: op1_01_in10 = reg_0028;
    50: op1_01_in10 = reg_0028;
    6: op1_01_in10 = reg_0335;
    7: op1_01_in10 = imem06_in[19:16];
    3: op1_01_in10 = reg_0444;
    8: op1_01_in10 = reg_0684;
    9: op1_01_in10 = imem03_in[23:20];
    10: op1_01_in10 = imem03_in[111:108];
    11: op1_01_in10 = reg_0453;
    12: op1_01_in10 = reg_0645;
    13: op1_01_in10 = imem07_in[75:72];
    14: op1_01_in10 = reg_0118;
    15: op1_01_in10 = reg_0355;
    16: op1_01_in10 = reg_0785;
    17: op1_01_in10 = reg_0678;
    18: op1_01_in10 = reg_0440;
    19: op1_01_in10 = reg_0455;
    20: op1_01_in10 = imem05_in[67:64];
    21: op1_01_in10 = reg_0450;
    81: op1_01_in10 = reg_0450;
    22: op1_01_in10 = reg_0329;
    23: op1_01_in10 = imem07_in[11:8];
    24: op1_01_in10 = reg_0343;
    25: op1_01_in10 = reg_0735;
    26: op1_01_in10 = reg_0357;
    27: op1_01_in10 = reg_0086;
    28: op1_01_in10 = reg_0480;
    29: op1_01_in10 = imem02_in[95:92];
    30: op1_01_in10 = reg_0085;
    31: op1_01_in10 = reg_0464;
    34: op1_01_in10 = reg_0464;
    42: op1_01_in10 = reg_0464;
    32: op1_01_in10 = imem02_in[27:24];
    33: op1_01_in10 = reg_0361;
    36: op1_01_in10 = reg_0470;
    37: op1_01_in10 = reg_0641;
    38: op1_01_in10 = reg_0114;
    39: op1_01_in10 = reg_0554;
    40: op1_01_in10 = reg_0571;
    41: op1_01_in10 = reg_0037;
    43: op1_01_in10 = imem02_in[55:52];
    44: op1_01_in10 = reg_0544;
    45: op1_01_in10 = reg_0720;
    46: op1_01_in10 = reg_0655;
    47: op1_01_in10 = reg_0597;
    48: op1_01_in10 = reg_0368;
    49: op1_01_in10 = reg_0175;
    51: op1_01_in10 = reg_0516;
    52: op1_01_in10 = reg_0328;
    53: op1_01_in10 = reg_0795;
    54: op1_01_in10 = reg_0101;
    55: op1_01_in10 = reg_0239;
    56: op1_01_in10 = reg_0688;
    57: op1_01_in10 = reg_0473;
    58: op1_01_in10 = reg_0718;
    59: op1_01_in10 = reg_0656;
    60: op1_01_in10 = reg_0194;
    61: op1_01_in10 = reg_0657;
    62: op1_01_in10 = imem05_in[123:120];
    63: op1_01_in10 = reg_0623;
    64: op1_01_in10 = reg_0703;
    65: op1_01_in10 = reg_0706;
    66: op1_01_in10 = reg_0717;
    68: op1_01_in10 = reg_0012;
    93: op1_01_in10 = reg_0012;
    69: op1_01_in10 = reg_0135;
    70: op1_01_in10 = reg_0451;
    71: op1_01_in10 = reg_0226;
    72: op1_01_in10 = reg_0434;
    74: op1_01_in10 = reg_0691;
    75: op1_01_in10 = reg_0320;
    76: op1_01_in10 = reg_0139;
    77: op1_01_in10 = imem05_in[31:28];
    78: op1_01_in10 = reg_0174;
    79: op1_01_in10 = reg_0710;
    80: op1_01_in10 = reg_0192;
    82: op1_01_in10 = imem06_in[39:36];
    83: op1_01_in10 = imem04_in[111:108];
    84: op1_01_in10 = imem06_in[87:84];
    85: op1_01_in10 = reg_0210;
    86: op1_01_in10 = reg_0787;
    87: op1_01_in10 = reg_0155;
    88: op1_01_in10 = reg_0460;
    89: op1_01_in10 = reg_0298;
    90: op1_01_in10 = reg_0726;
    92: op1_01_in10 = reg_0747;
    94: op1_01_in10 = reg_0582;
    95: op1_01_in10 = reg_0532;
    96: op1_01_in10 = reg_0260;
    default: op1_01_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv10 = 1;
    6: op1_01_inv10 = 1;
    7: op1_01_inv10 = 1;
    9: op1_01_inv10 = 1;
    10: op1_01_inv10 = 1;
    11: op1_01_inv10 = 1;
    13: op1_01_inv10 = 1;
    14: op1_01_inv10 = 1;
    18: op1_01_inv10 = 1;
    23: op1_01_inv10 = 1;
    24: op1_01_inv10 = 1;
    27: op1_01_inv10 = 1;
    28: op1_01_inv10 = 1;
    29: op1_01_inv10 = 1;
    31: op1_01_inv10 = 1;
    32: op1_01_inv10 = 1;
    33: op1_01_inv10 = 1;
    36: op1_01_inv10 = 1;
    38: op1_01_inv10 = 1;
    40: op1_01_inv10 = 1;
    41: op1_01_inv10 = 1;
    42: op1_01_inv10 = 1;
    43: op1_01_inv10 = 1;
    44: op1_01_inv10 = 1;
    45: op1_01_inv10 = 1;
    48: op1_01_inv10 = 1;
    50: op1_01_inv10 = 1;
    55: op1_01_inv10 = 1;
    56: op1_01_inv10 = 1;
    60: op1_01_inv10 = 1;
    61: op1_01_inv10 = 1;
    62: op1_01_inv10 = 1;
    63: op1_01_inv10 = 1;
    64: op1_01_inv10 = 1;
    65: op1_01_inv10 = 1;
    68: op1_01_inv10 = 1;
    70: op1_01_inv10 = 1;
    74: op1_01_inv10 = 1;
    76: op1_01_inv10 = 1;
    78: op1_01_inv10 = 1;
    80: op1_01_inv10 = 1;
    81: op1_01_inv10 = 1;
    82: op1_01_inv10 = 1;
    83: op1_01_inv10 = 1;
    84: op1_01_inv10 = 1;
    85: op1_01_inv10 = 1;
    88: op1_01_inv10 = 1;
    89: op1_01_inv10 = 1;
    90: op1_01_inv10 = 1;
    92: op1_01_inv10 = 1;
    93: op1_01_inv10 = 1;
    95: op1_01_inv10 = 1;
    96: op1_01_inv10 = 1;
    default: op1_01_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in11 = reg_0118;
    5: op1_01_in11 = reg_0025;
    6: op1_01_in11 = reg_0336;
    7: op1_01_in11 = imem06_in[27:24];
    87: op1_01_in11 = imem06_in[27:24];
    3: op1_01_in11 = reg_0175;
    78: op1_01_in11 = reg_0175;
    8: op1_01_in11 = reg_0671;
    9: op1_01_in11 = imem03_in[39:36];
    10: op1_01_in11 = reg_0602;
    11: op1_01_in11 = reg_0454;
    12: op1_01_in11 = reg_0653;
    13: op1_01_in11 = imem07_in[123:120];
    14: op1_01_in11 = reg_0116;
    15: op1_01_in11 = reg_0052;
    16: op1_01_in11 = reg_0264;
    17: op1_01_in11 = reg_0669;
    18: op1_01_in11 = reg_0427;
    19: op1_01_in11 = reg_0457;
    20: op1_01_in11 = imem05_in[83:80];
    21: op1_01_in11 = reg_0464;
    22: op1_01_in11 = reg_0363;
    23: op1_01_in11 = imem07_in[35:32];
    24: op1_01_in11 = reg_0388;
    25: op1_01_in11 = reg_0226;
    26: op1_01_in11 = reg_0769;
    27: op1_01_in11 = reg_0089;
    28: op1_01_in11 = reg_0467;
    42: op1_01_in11 = reg_0467;
    29: op1_01_in11 = imem02_in[99:96];
    30: op1_01_in11 = reg_0285;
    31: op1_01_in11 = reg_0461;
    32: op1_01_in11 = imem02_in[75:72];
    43: op1_01_in11 = imem02_in[75:72];
    33: op1_01_in11 = reg_0360;
    34: op1_01_in11 = reg_0472;
    36: op1_01_in11 = reg_0468;
    37: op1_01_in11 = reg_0643;
    38: op1_01_in11 = imem02_in[3:0];
    39: op1_01_in11 = reg_0523;
    40: op1_01_in11 = reg_0002;
    41: op1_01_in11 = imem07_in[59:56];
    44: op1_01_in11 = reg_0043;
    45: op1_01_in11 = reg_0724;
    64: op1_01_in11 = reg_0724;
    46: op1_01_in11 = reg_0637;
    47: op1_01_in11 = reg_0395;
    48: op1_01_in11 = reg_0231;
    49: op1_01_in11 = reg_0180;
    50: op1_01_in11 = reg_0242;
    51: op1_01_in11 = reg_0308;
    52: op1_01_in11 = reg_0555;
    53: op1_01_in11 = reg_0793;
    54: op1_01_in11 = reg_0132;
    55: op1_01_in11 = reg_0434;
    56: op1_01_in11 = reg_0465;
    57: op1_01_in11 = reg_0191;
    58: op1_01_in11 = reg_0707;
    59: op1_01_in11 = reg_0651;
    60: op1_01_in11 = reg_0201;
    61: op1_01_in11 = reg_0641;
    62: op1_01_in11 = reg_0781;
    63: op1_01_in11 = imem07_in[11:8];
    65: op1_01_in11 = reg_0445;
    66: op1_01_in11 = reg_0702;
    68: op1_01_in11 = reg_0803;
    69: op1_01_in11 = reg_0133;
    70: op1_01_in11 = reg_0455;
    71: op1_01_in11 = reg_0489;
    72: op1_01_in11 = reg_0166;
    90: op1_01_in11 = reg_0166;
    74: op1_01_in11 = reg_0688;
    75: op1_01_in11 = reg_0581;
    76: op1_01_in11 = reg_0548;
    77: op1_01_in11 = imem05_in[35:32];
    79: op1_01_in11 = reg_0159;
    80: op1_01_in11 = imem01_in[11:8];
    81: op1_01_in11 = reg_0462;
    82: op1_01_in11 = imem06_in[67:64];
    83: op1_01_in11 = reg_0171;
    84: op1_01_in11 = imem06_in[107:104];
    85: op1_01_in11 = reg_0195;
    86: op1_01_in11 = reg_0767;
    88: op1_01_in11 = reg_0479;
    89: op1_01_in11 = reg_0038;
    92: op1_01_in11 = reg_0557;
    93: op1_01_in11 = reg_0801;
    94: op1_01_in11 = reg_0367;
    95: op1_01_in11 = imem03_in[31:28];
    96: op1_01_in11 = reg_0304;
    default: op1_01_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv11 = 1;
    3: op1_01_inv11 = 1;
    9: op1_01_inv11 = 1;
    12: op1_01_inv11 = 1;
    13: op1_01_inv11 = 1;
    15: op1_01_inv11 = 1;
    16: op1_01_inv11 = 1;
    17: op1_01_inv11 = 1;
    18: op1_01_inv11 = 1;
    21: op1_01_inv11 = 1;
    22: op1_01_inv11 = 1;
    25: op1_01_inv11 = 1;
    26: op1_01_inv11 = 1;
    27: op1_01_inv11 = 1;
    28: op1_01_inv11 = 1;
    29: op1_01_inv11 = 1;
    30: op1_01_inv11 = 1;
    31: op1_01_inv11 = 1;
    33: op1_01_inv11 = 1;
    36: op1_01_inv11 = 1;
    38: op1_01_inv11 = 1;
    39: op1_01_inv11 = 1;
    40: op1_01_inv11 = 1;
    43: op1_01_inv11 = 1;
    48: op1_01_inv11 = 1;
    54: op1_01_inv11 = 1;
    57: op1_01_inv11 = 1;
    58: op1_01_inv11 = 1;
    59: op1_01_inv11 = 1;
    60: op1_01_inv11 = 1;
    64: op1_01_inv11 = 1;
    66: op1_01_inv11 = 1;
    68: op1_01_inv11 = 1;
    69: op1_01_inv11 = 1;
    71: op1_01_inv11 = 1;
    74: op1_01_inv11 = 1;
    76: op1_01_inv11 = 1;
    77: op1_01_inv11 = 1;
    78: op1_01_inv11 = 1;
    81: op1_01_inv11 = 1;
    86: op1_01_inv11 = 1;
    90: op1_01_inv11 = 1;
    default: op1_01_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in12 = reg_0104;
    14: op1_01_in12 = reg_0104;
    5: op1_01_in12 = imem07_in[47:44];
    23: op1_01_in12 = imem07_in[47:44];
    6: op1_01_in12 = reg_0089;
    7: op1_01_in12 = imem06_in[91:88];
    3: op1_01_in12 = reg_0180;
    8: op1_01_in12 = reg_0688;
    9: op1_01_in12 = imem03_in[47:44];
    10: op1_01_in12 = reg_0582;
    11: op1_01_in12 = reg_0469;
    21: op1_01_in12 = reg_0469;
    12: op1_01_in12 = reg_0637;
    13: op1_01_in12 = imem07_in[127:124];
    15: op1_01_in12 = reg_0086;
    16: op1_01_in12 = reg_0732;
    17: op1_01_in12 = reg_0481;
    81: op1_01_in12 = reg_0481;
    18: op1_01_in12 = reg_0181;
    49: op1_01_in12 = reg_0181;
    19: op1_01_in12 = reg_0464;
    20: op1_01_in12 = reg_0792;
    22: op1_01_in12 = reg_0338;
    24: op1_01_in12 = reg_0362;
    25: op1_01_in12 = reg_0733;
    26: op1_01_in12 = reg_0539;
    27: op1_01_in12 = reg_0134;
    28: op1_01_in12 = reg_0200;
    29: op1_01_in12 = imem02_in[103:100];
    30: op1_01_in12 = reg_0156;
    31: op1_01_in12 = reg_0466;
    32: op1_01_in12 = reg_0645;
    33: op1_01_in12 = reg_0346;
    34: op1_01_in12 = reg_0479;
    36: op1_01_in12 = reg_0459;
    37: op1_01_in12 = reg_0659;
    38: op1_01_in12 = imem02_in[31:28];
    39: op1_01_in12 = reg_0558;
    40: op1_01_in12 = reg_0803;
    41: op1_01_in12 = imem07_in[83:80];
    42: op1_01_in12 = reg_0214;
    43: op1_01_in12 = imem02_in[91:88];
    44: op1_01_in12 = reg_0088;
    45: op1_01_in12 = reg_0715;
    46: op1_01_in12 = reg_0664;
    47: op1_01_in12 = reg_0384;
    48: op1_01_in12 = imem07_in[11:8];
    50: op1_01_in12 = reg_0031;
    51: op1_01_in12 = reg_0076;
    52: op1_01_in12 = reg_0057;
    53: op1_01_in12 = reg_0786;
    54: op1_01_in12 = reg_0149;
    55: op1_01_in12 = reg_0435;
    56: op1_01_in12 = reg_0476;
    57: op1_01_in12 = reg_0204;
    58: op1_01_in12 = reg_0700;
    59: op1_01_in12 = reg_0345;
    60: op1_01_in12 = reg_0205;
    61: op1_01_in12 = reg_0427;
    62: op1_01_in12 = reg_0789;
    63: op1_01_in12 = imem07_in[31:28];
    64: op1_01_in12 = reg_0729;
    65: op1_01_in12 = reg_0440;
    66: op1_01_in12 = reg_0712;
    68: op1_01_in12 = reg_0008;
    69: op1_01_in12 = reg_0152;
    70: op1_01_in12 = reg_0461;
    71: op1_01_in12 = reg_0246;
    74: op1_01_in12 = reg_0247;
    75: op1_01_in12 = reg_0514;
    76: op1_01_in12 = reg_0702;
    77: op1_01_in12 = imem05_in[47:44];
    78: op1_01_in12 = reg_0172;
    79: op1_01_in12 = reg_0784;
    80: op1_01_in12 = imem01_in[23:20];
    82: op1_01_in12 = imem06_in[75:72];
    83: op1_01_in12 = reg_0173;
    84: op1_01_in12 = imem06_in[119:116];
    85: op1_01_in12 = reg_0206;
    86: op1_01_in12 = reg_0661;
    87: op1_01_in12 = imem06_in[59:56];
    88: op1_01_in12 = reg_0452;
    89: op1_01_in12 = reg_0402;
    90: op1_01_in12 = reg_0711;
    92: op1_01_in12 = reg_0570;
    93: op1_01_in12 = reg_0799;
    94: op1_01_in12 = reg_0003;
    95: op1_01_in12 = imem03_in[91:88];
    96: op1_01_in12 = reg_0000;
    default: op1_01_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv12 = 1;
    6: op1_01_inv12 = 1;
    7: op1_01_inv12 = 1;
    3: op1_01_inv12 = 1;
    9: op1_01_inv12 = 1;
    11: op1_01_inv12 = 1;
    14: op1_01_inv12 = 1;
    16: op1_01_inv12 = 1;
    17: op1_01_inv12 = 1;
    18: op1_01_inv12 = 1;
    20: op1_01_inv12 = 1;
    22: op1_01_inv12 = 1;
    25: op1_01_inv12 = 1;
    26: op1_01_inv12 = 1;
    27: op1_01_inv12 = 1;
    28: op1_01_inv12 = 1;
    29: op1_01_inv12 = 1;
    30: op1_01_inv12 = 1;
    34: op1_01_inv12 = 1;
    39: op1_01_inv12 = 1;
    40: op1_01_inv12 = 1;
    42: op1_01_inv12 = 1;
    45: op1_01_inv12 = 1;
    46: op1_01_inv12 = 1;
    47: op1_01_inv12 = 1;
    49: op1_01_inv12 = 1;
    50: op1_01_inv12 = 1;
    54: op1_01_inv12 = 1;
    55: op1_01_inv12 = 1;
    57: op1_01_inv12 = 1;
    59: op1_01_inv12 = 1;
    60: op1_01_inv12 = 1;
    61: op1_01_inv12 = 1;
    64: op1_01_inv12 = 1;
    65: op1_01_inv12 = 1;
    69: op1_01_inv12 = 1;
    71: op1_01_inv12 = 1;
    74: op1_01_inv12 = 1;
    76: op1_01_inv12 = 1;
    77: op1_01_inv12 = 1;
    82: op1_01_inv12 = 1;
    84: op1_01_inv12 = 1;
    87: op1_01_inv12 = 1;
    92: op1_01_inv12 = 1;
    94: op1_01_inv12 = 1;
    95: op1_01_inv12 = 1;
    96: op1_01_inv12 = 1;
    default: op1_01_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in13 = reg_0100;
    5: op1_01_in13 = imem07_in[123:120];
    6: op1_01_in13 = reg_0096;
    7: op1_01_in13 = imem06_in[95:92];
    3: op1_01_in13 = reg_0162;
    49: op1_01_in13 = reg_0162;
    8: op1_01_in13 = reg_0462;
    9: op1_01_in13 = imem03_in[51:48];
    10: op1_01_in13 = reg_0572;
    11: op1_01_in13 = reg_0472;
    12: op1_01_in13 = reg_0651;
    13: op1_01_in13 = reg_0729;
    14: op1_01_in13 = reg_0119;
    15: op1_01_in13 = reg_0055;
    16: op1_01_in13 = reg_0132;
    17: op1_01_in13 = reg_0473;
    18: op1_01_in13 = reg_0179;
    19: op1_01_in13 = reg_0469;
    20: op1_01_in13 = reg_0490;
    21: op1_01_in13 = reg_0467;
    22: op1_01_in13 = reg_0355;
    23: op1_01_in13 = imem07_in[55:52];
    24: op1_01_in13 = reg_0369;
    25: op1_01_in13 = reg_0282;
    26: op1_01_in13 = reg_0740;
    27: op1_01_in13 = imem06_in[63:60];
    28: op1_01_in13 = reg_0203;
    29: op1_01_in13 = imem02_in[111:108];
    30: op1_01_in13 = reg_0139;
    31: op1_01_in13 = reg_0480;
    81: op1_01_in13 = reg_0480;
    32: op1_01_in13 = reg_0658;
    33: op1_01_in13 = reg_0342;
    34: op1_01_in13 = reg_0452;
    36: op1_01_in13 = reg_0200;
    37: op1_01_in13 = reg_0352;
    61: op1_01_in13 = reg_0352;
    38: op1_01_in13 = imem02_in[39:36];
    39: op1_01_in13 = reg_0516;
    40: op1_01_in13 = reg_0805;
    41: op1_01_in13 = reg_0713;
    64: op1_01_in13 = reg_0713;
    42: op1_01_in13 = reg_0208;
    43: op1_01_in13 = imem02_in[95:92];
    44: op1_01_in13 = reg_0280;
    45: op1_01_in13 = reg_0707;
    46: op1_01_in13 = reg_0657;
    47: op1_01_in13 = reg_0575;
    48: op1_01_in13 = imem07_in[51:48];
    50: op1_01_in13 = reg_0753;
    51: op1_01_in13 = reg_0077;
    52: op1_01_in13 = reg_0536;
    53: op1_01_in13 = reg_0091;
    54: op1_01_in13 = reg_0142;
    55: op1_01_in13 = reg_0180;
    56: op1_01_in13 = reg_0466;
    57: op1_01_in13 = reg_0211;
    58: op1_01_in13 = reg_0441;
    59: op1_01_in13 = reg_0361;
    60: op1_01_in13 = reg_0202;
    62: op1_01_in13 = reg_0491;
    63: op1_01_in13 = imem07_in[47:44];
    65: op1_01_in13 = reg_0437;
    66: op1_01_in13 = reg_0709;
    68: op1_01_in13 = reg_0004;
    69: op1_01_in13 = reg_0153;
    70: op1_01_in13 = reg_0477;
    71: op1_01_in13 = reg_0276;
    74: op1_01_in13 = reg_0692;
    75: op1_01_in13 = reg_0743;
    76: op1_01_in13 = reg_0358;
    77: op1_01_in13 = imem05_in[63:60];
    78: op1_01_in13 = reg_0171;
    79: op1_01_in13 = reg_0382;
    80: op1_01_in13 = imem01_in[51:48];
    82: op1_01_in13 = imem06_in[83:80];
    83: op1_01_in13 = reg_0275;
    84: op1_01_in13 = imem06_in[127:124];
    85: op1_01_in13 = imem01_in[3:0];
    86: op1_01_in13 = reg_0367;
    87: op1_01_in13 = imem06_in[99:96];
    88: op1_01_in13 = reg_0189;
    89: op1_01_in13 = reg_0405;
    90: op1_01_in13 = reg_0103;
    92: op1_01_in13 = reg_0811;
    93: op1_01_in13 = reg_0589;
    94: op1_01_in13 = reg_0595;
    95: op1_01_in13 = reg_0509;
    96: op1_01_in13 = reg_0498;
    default: op1_01_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_01_inv13 = 1;
    10: op1_01_inv13 = 1;
    12: op1_01_inv13 = 1;
    14: op1_01_inv13 = 1;
    15: op1_01_inv13 = 1;
    16: op1_01_inv13 = 1;
    17: op1_01_inv13 = 1;
    19: op1_01_inv13 = 1;
    20: op1_01_inv13 = 1;
    22: op1_01_inv13 = 1;
    23: op1_01_inv13 = 1;
    25: op1_01_inv13 = 1;
    26: op1_01_inv13 = 1;
    27: op1_01_inv13 = 1;
    28: op1_01_inv13 = 1;
    31: op1_01_inv13 = 1;
    32: op1_01_inv13 = 1;
    33: op1_01_inv13 = 1;
    34: op1_01_inv13 = 1;
    36: op1_01_inv13 = 1;
    37: op1_01_inv13 = 1;
    38: op1_01_inv13 = 1;
    39: op1_01_inv13 = 1;
    41: op1_01_inv13 = 1;
    42: op1_01_inv13 = 1;
    43: op1_01_inv13 = 1;
    49: op1_01_inv13 = 1;
    50: op1_01_inv13 = 1;
    52: op1_01_inv13 = 1;
    53: op1_01_inv13 = 1;
    58: op1_01_inv13 = 1;
    59: op1_01_inv13 = 1;
    62: op1_01_inv13 = 1;
    63: op1_01_inv13 = 1;
    64: op1_01_inv13 = 1;
    65: op1_01_inv13 = 1;
    66: op1_01_inv13 = 1;
    71: op1_01_inv13 = 1;
    75: op1_01_inv13 = 1;
    81: op1_01_inv13 = 1;
    83: op1_01_inv13 = 1;
    84: op1_01_inv13 = 1;
    90: op1_01_inv13 = 1;
    92: op1_01_inv13 = 1;
    93: op1_01_inv13 = 1;
    94: op1_01_inv13 = 1;
    95: op1_01_inv13 = 1;
    96: op1_01_inv13 = 1;
    default: op1_01_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in14 = reg_0109;
    5: op1_01_in14 = reg_0717;
    6: op1_01_in14 = reg_0082;
    7: op1_01_in14 = reg_0614;
    3: op1_01_in14 = reg_0169;
    8: op1_01_in14 = reg_0206;
    60: op1_01_in14 = reg_0206;
    9: op1_01_in14 = imem03_in[71:68];
    10: op1_01_in14 = reg_0587;
    11: op1_01_in14 = reg_0473;
    12: op1_01_in14 = reg_0662;
    13: op1_01_in14 = reg_0706;
    45: op1_01_in14 = reg_0706;
    14: op1_01_in14 = reg_0115;
    15: op1_01_in14 = reg_0060;
    16: op1_01_in14 = reg_0148;
    17: op1_01_in14 = reg_0456;
    81: op1_01_in14 = reg_0456;
    18: op1_01_in14 = reg_0167;
    49: op1_01_in14 = reg_0167;
    19: op1_01_in14 = reg_0466;
    20: op1_01_in14 = reg_0491;
    21: op1_01_in14 = reg_0468;
    22: op1_01_in14 = reg_0336;
    23: op1_01_in14 = imem07_in[63:60];
    24: op1_01_in14 = reg_0393;
    25: op1_01_in14 = reg_0744;
    26: op1_01_in14 = imem03_in[43:40];
    27: op1_01_in14 = imem06_in[95:92];
    28: op1_01_in14 = reg_0193;
    42: op1_01_in14 = reg_0193;
    29: op1_01_in14 = imem02_in[123:120];
    30: op1_01_in14 = reg_0138;
    31: op1_01_in14 = reg_0470;
    74: op1_01_in14 = reg_0470;
    32: op1_01_in14 = reg_0653;
    33: op1_01_in14 = reg_0321;
    34: op1_01_in14 = reg_0478;
    36: op1_01_in14 = reg_0187;
    37: op1_01_in14 = reg_0349;
    38: op1_01_in14 = imem02_in[47:44];
    39: op1_01_in14 = reg_0303;
    40: op1_01_in14 = reg_0008;
    41: op1_01_in14 = reg_0436;
    43: op1_01_in14 = reg_0664;
    44: op1_01_in14 = reg_0430;
    46: op1_01_in14 = reg_0301;
    47: op1_01_in14 = reg_0564;
    48: op1_01_in14 = imem07_in[95:92];
    50: op1_01_in14 = reg_0777;
    51: op1_01_in14 = reg_0626;
    52: op1_01_in14 = reg_0556;
    53: op1_01_in14 = reg_0246;
    54: op1_01_in14 = imem06_in[7:4];
    55: op1_01_in14 = reg_0159;
    56: op1_01_in14 = reg_0480;
    57: op1_01_in14 = reg_0205;
    58: op1_01_in14 = reg_0434;
    59: op1_01_in14 = reg_0365;
    61: op1_01_in14 = reg_0358;
    62: op1_01_in14 = reg_0782;
    63: op1_01_in14 = imem07_in[51:48];
    64: op1_01_in14 = reg_0701;
    65: op1_01_in14 = reg_0175;
    66: op1_01_in14 = reg_0705;
    68: op1_01_in14 = imem04_in[7:4];
    69: op1_01_in14 = reg_0137;
    70: op1_01_in14 = reg_0474;
    71: op1_01_in14 = reg_0249;
    75: op1_01_in14 = reg_0095;
    76: op1_01_in14 = reg_0363;
    77: op1_01_in14 = imem05_in[87:84];
    78: op1_01_in14 = reg_0184;
    79: op1_01_in14 = reg_0709;
    80: op1_01_in14 = imem01_in[83:80];
    82: op1_01_in14 = reg_0289;
    83: op1_01_in14 = reg_0058;
    84: op1_01_in14 = reg_0293;
    85: op1_01_in14 = imem01_in[23:20];
    86: op1_01_in14 = imem07_in[3:0];
    87: op1_01_in14 = reg_0577;
    88: op1_01_in14 = reg_0188;
    89: op1_01_in14 = reg_0763;
    90: op1_01_in14 = reg_0727;
    92: op1_01_in14 = reg_0561;
    93: op1_01_in14 = reg_0389;
    94: op1_01_in14 = reg_0575;
    95: op1_01_in14 = reg_0003;
    96: op1_01_in14 = reg_0219;
    default: op1_01_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_01_inv14 = 1;
    3: op1_01_inv14 = 1;
    10: op1_01_inv14 = 1;
    11: op1_01_inv14 = 1;
    15: op1_01_inv14 = 1;
    17: op1_01_inv14 = 1;
    19: op1_01_inv14 = 1;
    20: op1_01_inv14 = 1;
    21: op1_01_inv14 = 1;
    22: op1_01_inv14 = 1;
    26: op1_01_inv14 = 1;
    28: op1_01_inv14 = 1;
    29: op1_01_inv14 = 1;
    31: op1_01_inv14 = 1;
    34: op1_01_inv14 = 1;
    36: op1_01_inv14 = 1;
    44: op1_01_inv14 = 1;
    47: op1_01_inv14 = 1;
    52: op1_01_inv14 = 1;
    53: op1_01_inv14 = 1;
    55: op1_01_inv14 = 1;
    57: op1_01_inv14 = 1;
    62: op1_01_inv14 = 1;
    64: op1_01_inv14 = 1;
    66: op1_01_inv14 = 1;
    70: op1_01_inv14 = 1;
    71: op1_01_inv14 = 1;
    80: op1_01_inv14 = 1;
    83: op1_01_inv14 = 1;
    87: op1_01_inv14 = 1;
    88: op1_01_inv14 = 1;
    93: op1_01_inv14 = 1;
    default: op1_01_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in15 = imem02_in[23:20];
    5: op1_01_in15 = reg_0725;
    6: op1_01_in15 = reg_0091;
    7: op1_01_in15 = reg_0607;
    3: op1_01_in15 = reg_0177;
    83: op1_01_in15 = reg_0177;
    8: op1_01_in15 = reg_0199;
    57: op1_01_in15 = reg_0199;
    9: op1_01_in15 = imem03_in[83:80];
    10: op1_01_in15 = reg_0600;
    11: op1_01_in15 = reg_0452;
    12: op1_01_in15 = reg_0644;
    13: op1_01_in15 = reg_0432;
    52: op1_01_in15 = reg_0432;
    14: op1_01_in15 = reg_0110;
    15: op1_01_in15 = reg_0094;
    16: op1_01_in15 = reg_0135;
    17: op1_01_in15 = reg_0188;
    81: op1_01_in15 = reg_0188;
    19: op1_01_in15 = reg_0467;
    20: op1_01_in15 = reg_0795;
    21: op1_01_in15 = reg_0459;
    22: op1_01_in15 = reg_0518;
    23: op1_01_in15 = imem07_in[75:72];
    24: op1_01_in15 = reg_0396;
    25: op1_01_in15 = reg_0734;
    26: op1_01_in15 = imem03_in[47:44];
    27: op1_01_in15 = imem06_in[107:104];
    28: op1_01_in15 = reg_0194;
    34: op1_01_in15 = reg_0194;
    29: op1_01_in15 = reg_0666;
    30: op1_01_in15 = reg_0140;
    31: op1_01_in15 = reg_0456;
    32: op1_01_in15 = reg_0639;
    33: op1_01_in15 = reg_0323;
    36: op1_01_in15 = reg_0211;
    37: op1_01_in15 = reg_0357;
    38: op1_01_in15 = imem02_in[59:56];
    39: op1_01_in15 = reg_0280;
    40: op1_01_in15 = reg_0806;
    41: op1_01_in15 = reg_0445;
    42: op1_01_in15 = reg_0207;
    88: op1_01_in15 = reg_0207;
    43: op1_01_in15 = reg_0659;
    44: op1_01_in15 = reg_0617;
    45: op1_01_in15 = reg_0700;
    46: op1_01_in15 = reg_0638;
    47: op1_01_in15 = reg_0569;
    48: op1_01_in15 = reg_0722;
    49: op1_01_in15 = reg_0163;
    50: op1_01_in15 = reg_0368;
    51: op1_01_in15 = reg_0610;
    53: op1_01_in15 = reg_0304;
    54: op1_01_in15 = imem06_in[15:12];
    55: op1_01_in15 = reg_0183;
    56: op1_01_in15 = reg_0471;
    58: op1_01_in15 = reg_0444;
    59: op1_01_in15 = reg_0527;
    60: op1_01_in15 = imem01_in[7:4];
    61: op1_01_in15 = reg_0341;
    62: op1_01_in15 = reg_0786;
    63: op1_01_in15 = imem07_in[63:60];
    64: op1_01_in15 = reg_0253;
    65: op1_01_in15 = reg_0181;
    66: op1_01_in15 = reg_0436;
    68: op1_01_in15 = imem04_in[15:12];
    69: op1_01_in15 = imem06_in[19:16];
    70: op1_01_in15 = reg_0214;
    71: op1_01_in15 = reg_0383;
    74: op1_01_in15 = reg_0209;
    75: op1_01_in15 = reg_0535;
    76: op1_01_in15 = reg_0324;
    77: op1_01_in15 = imem05_in[111:108];
    79: op1_01_in15 = reg_0731;
    80: op1_01_in15 = imem01_in[107:104];
    82: op1_01_in15 = reg_0346;
    84: op1_01_in15 = reg_0270;
    85: op1_01_in15 = imem01_in[87:84];
    86: op1_01_in15 = imem07_in[35:32];
    87: op1_01_in15 = reg_0370;
    89: op1_01_in15 = reg_0242;
    90: op1_01_in15 = reg_0061;
    92: op1_01_in15 = reg_0248;
    93: op1_01_in15 = reg_0575;
    94: op1_01_in15 = reg_0417;
    95: op1_01_in15 = reg_0595;
    96: op1_01_in15 = reg_0106;
    default: op1_01_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_01_inv15 = 1;
    3: op1_01_inv15 = 1;
    8: op1_01_inv15 = 1;
    10: op1_01_inv15 = 1;
    12: op1_01_inv15 = 1;
    14: op1_01_inv15 = 1;
    15: op1_01_inv15 = 1;
    16: op1_01_inv15 = 1;
    22: op1_01_inv15 = 1;
    23: op1_01_inv15 = 1;
    24: op1_01_inv15 = 1;
    26: op1_01_inv15 = 1;
    27: op1_01_inv15 = 1;
    29: op1_01_inv15 = 1;
    32: op1_01_inv15 = 1;
    33: op1_01_inv15 = 1;
    34: op1_01_inv15 = 1;
    36: op1_01_inv15 = 1;
    37: op1_01_inv15 = 1;
    38: op1_01_inv15 = 1;
    39: op1_01_inv15 = 1;
    40: op1_01_inv15 = 1;
    42: op1_01_inv15 = 1;
    43: op1_01_inv15 = 1;
    45: op1_01_inv15 = 1;
    52: op1_01_inv15 = 1;
    53: op1_01_inv15 = 1;
    54: op1_01_inv15 = 1;
    56: op1_01_inv15 = 1;
    58: op1_01_inv15 = 1;
    60: op1_01_inv15 = 1;
    61: op1_01_inv15 = 1;
    66: op1_01_inv15 = 1;
    71: op1_01_inv15 = 1;
    75: op1_01_inv15 = 1;
    80: op1_01_inv15 = 1;
    81: op1_01_inv15 = 1;
    82: op1_01_inv15 = 1;
    83: op1_01_inv15 = 1;
    84: op1_01_inv15 = 1;
    85: op1_01_inv15 = 1;
    89: op1_01_inv15 = 1;
    90: op1_01_inv15 = 1;
    92: op1_01_inv15 = 1;
    94: op1_01_inv15 = 1;
    96: op1_01_inv15 = 1;
    default: op1_01_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in16 = imem02_in[43:40];
    5: op1_01_in16 = reg_0701;
    6: op1_01_in16 = reg_0094;
    7: op1_01_in16 = reg_0608;
    3: op1_01_in16 = reg_0170;
    8: op1_01_in16 = imem01_in[23:20];
    60: op1_01_in16 = imem01_in[23:20];
    9: op1_01_in16 = imem03_in[87:84];
    10: op1_01_in16 = reg_0578;
    11: op1_01_in16 = reg_0478;
    21: op1_01_in16 = reg_0478;
    12: op1_01_in16 = reg_0643;
    13: op1_01_in16 = reg_0426;
    14: op1_01_in16 = imem02_in[31:28];
    15: op1_01_in16 = imem03_in[7:4];
    16: op1_01_in16 = reg_0143;
    17: op1_01_in16 = reg_0198;
    19: op1_01_in16 = reg_0471;
    20: op1_01_in16 = reg_0485;
    22: op1_01_in16 = reg_0314;
    33: op1_01_in16 = reg_0314;
    23: op1_01_in16 = imem07_in[91:88];
    24: op1_01_in16 = reg_0374;
    25: op1_01_in16 = reg_0149;
    26: op1_01_in16 = imem03_in[67:64];
    27: op1_01_in16 = imem06_in[123:120];
    28: op1_01_in16 = imem01_in[15:12];
    29: op1_01_in16 = reg_0646;
    94: op1_01_in16 = reg_0646;
    30: op1_01_in16 = reg_0155;
    31: op1_01_in16 = reg_0187;
    70: op1_01_in16 = reg_0187;
    32: op1_01_in16 = reg_0662;
    34: op1_01_in16 = reg_0199;
    36: op1_01_in16 = reg_0194;
    37: op1_01_in16 = reg_0356;
    38: op1_01_in16 = imem02_in[83:80];
    39: op1_01_in16 = reg_0294;
    40: op1_01_in16 = reg_0010;
    41: op1_01_in16 = reg_0439;
    42: op1_01_in16 = reg_0211;
    43: op1_01_in16 = reg_0667;
    44: op1_01_in16 = reg_0258;
    45: op1_01_in16 = reg_0334;
    46: op1_01_in16 = reg_0357;
    51: op1_01_in16 = reg_0357;
    47: op1_01_in16 = reg_0562;
    48: op1_01_in16 = reg_0728;
    49: op1_01_in16 = reg_0168;
    50: op1_01_in16 = reg_0375;
    52: op1_01_in16 = reg_0302;
    53: op1_01_in16 = reg_0742;
    54: op1_01_in16 = imem06_in[35:32];
    55: op1_01_in16 = reg_0166;
    56: op1_01_in16 = reg_0479;
    57: op1_01_in16 = imem01_in[3:0];
    58: op1_01_in16 = reg_0442;
    59: op1_01_in16 = reg_0518;
    61: op1_01_in16 = reg_0345;
    62: op1_01_in16 = reg_0489;
    63: op1_01_in16 = imem07_in[67:64];
    64: op1_01_in16 = reg_0635;
    65: op1_01_in16 = reg_0164;
    66: op1_01_in16 = reg_0636;
    68: op1_01_in16 = imem04_in[47:44];
    69: op1_01_in16 = imem06_in[23:20];
    71: op1_01_in16 = reg_0145;
    74: op1_01_in16 = reg_0193;
    75: op1_01_in16 = imem03_in[31:28];
    76: op1_01_in16 = reg_0351;
    77: op1_01_in16 = imem05_in[119:116];
    79: op1_01_in16 = reg_0064;
    80: op1_01_in16 = reg_0653;
    81: op1_01_in16 = reg_0207;
    82: op1_01_in16 = reg_0624;
    83: op1_01_in16 = reg_0542;
    84: op1_01_in16 = reg_0029;
    85: op1_01_in16 = imem01_in[91:88];
    86: op1_01_in16 = imem07_in[39:36];
    87: op1_01_in16 = reg_0609;
    88: op1_01_in16 = imem01_in[39:36];
    89: op1_01_in16 = reg_0515;
    90: op1_01_in16 = reg_0239;
    92: op1_01_in16 = reg_0013;
    93: op1_01_in16 = reg_0372;
    95: op1_01_in16 = reg_0747;
    96: op1_01_in16 = reg_0676;
    default: op1_01_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv16 = 1;
    5: op1_01_inv16 = 1;
    7: op1_01_inv16 = 1;
    8: op1_01_inv16 = 1;
    10: op1_01_inv16 = 1;
    12: op1_01_inv16 = 1;
    13: op1_01_inv16 = 1;
    15: op1_01_inv16 = 1;
    22: op1_01_inv16 = 1;
    23: op1_01_inv16 = 1;
    25: op1_01_inv16 = 1;
    29: op1_01_inv16 = 1;
    30: op1_01_inv16 = 1;
    32: op1_01_inv16 = 1;
    33: op1_01_inv16 = 1;
    37: op1_01_inv16 = 1;
    38: op1_01_inv16 = 1;
    40: op1_01_inv16 = 1;
    41: op1_01_inv16 = 1;
    42: op1_01_inv16 = 1;
    44: op1_01_inv16 = 1;
    45: op1_01_inv16 = 1;
    46: op1_01_inv16 = 1;
    48: op1_01_inv16 = 1;
    50: op1_01_inv16 = 1;
    51: op1_01_inv16 = 1;
    53: op1_01_inv16 = 1;
    55: op1_01_inv16 = 1;
    56: op1_01_inv16 = 1;
    57: op1_01_inv16 = 1;
    65: op1_01_inv16 = 1;
    66: op1_01_inv16 = 1;
    76: op1_01_inv16 = 1;
    80: op1_01_inv16 = 1;
    82: op1_01_inv16 = 1;
    84: op1_01_inv16 = 1;
    85: op1_01_inv16 = 1;
    87: op1_01_inv16 = 1;
    88: op1_01_inv16 = 1;
    89: op1_01_inv16 = 1;
    90: op1_01_inv16 = 1;
    92: op1_01_inv16 = 1;
    95: op1_01_inv16 = 1;
    default: op1_01_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in17 = imem02_in[71:68];
    5: op1_01_in17 = reg_0436;
    6: op1_01_in17 = reg_0073;
    7: op1_01_in17 = reg_0618;
    8: op1_01_in17 = imem01_in[43:40];
    9: op1_01_in17 = imem03_in[123:120];
    10: op1_01_in17 = reg_0597;
    11: op1_01_in17 = reg_0210;
    12: op1_01_in17 = reg_0665;
    13: op1_01_in17 = reg_0175;
    14: op1_01_in17 = imem02_in[39:36];
    15: op1_01_in17 = imem03_in[79:76];
    16: op1_01_in17 = reg_0130;
    17: op1_01_in17 = reg_0196;
    19: op1_01_in17 = reg_0459;
    20: op1_01_in17 = reg_0741;
    21: op1_01_in17 = imem01_in[31:28];
    22: op1_01_in17 = reg_0080;
    23: op1_01_in17 = imem07_in[99:96];
    24: op1_01_in17 = reg_0012;
    25: op1_01_in17 = reg_0150;
    26: op1_01_in17 = imem03_in[119:116];
    27: op1_01_in17 = imem06_in[127:124];
    28: op1_01_in17 = imem01_in[99:96];
    29: op1_01_in17 = reg_0647;
    30: op1_01_in17 = imem06_in[7:4];
    71: op1_01_in17 = imem06_in[7:4];
    31: op1_01_in17 = reg_0209;
    32: op1_01_in17 = reg_0362;
    33: op1_01_in17 = reg_0770;
    34: op1_01_in17 = imem01_in[15:12];
    57: op1_01_in17 = imem01_in[15:12];
    36: op1_01_in17 = reg_0198;
    37: op1_01_in17 = reg_0342;
    38: op1_01_in17 = reg_0660;
    39: op1_01_in17 = reg_0050;
    40: op1_01_in17 = imem04_in[35:32];
    41: op1_01_in17 = reg_0446;
    42: op1_01_in17 = reg_0213;
    43: op1_01_in17 = reg_0358;
    44: op1_01_in17 = reg_0256;
    45: op1_01_in17 = reg_0636;
    46: op1_01_in17 = reg_0341;
    47: op1_01_in17 = reg_0747;
    48: op1_01_in17 = reg_0704;
    49: op1_01_in17 = reg_0170;
    50: op1_01_in17 = reg_0029;
    51: op1_01_in17 = reg_0520;
    52: op1_01_in17 = reg_0503;
    53: op1_01_in17 = reg_0103;
    54: op1_01_in17 = imem06_in[59:56];
    55: op1_01_in17 = reg_0158;
    56: op1_01_in17 = reg_0214;
    58: op1_01_in17 = reg_0162;
    59: op1_01_in17 = imem03_in[11:8];
    60: op1_01_in17 = imem01_in[87:84];
    61: op1_01_in17 = reg_0594;
    62: op1_01_in17 = reg_0090;
    63: op1_01_in17 = imem07_in[91:88];
    64: op1_01_in17 = reg_0434;
    65: op1_01_in17 = reg_0168;
    66: op1_01_in17 = reg_0437;
    68: op1_01_in17 = imem04_in[51:48];
    69: op1_01_in17 = imem06_in[39:36];
    70: op1_01_in17 = reg_0203;
    74: op1_01_in17 = reg_0190;
    75: op1_01_in17 = imem03_in[103:100];
    76: op1_01_in17 = reg_0518;
    77: op1_01_in17 = imem05_in[123:120];
    79: op1_01_in17 = reg_0266;
    80: op1_01_in17 = reg_0668;
    81: op1_01_in17 = reg_0201;
    82: op1_01_in17 = reg_0609;
    83: op1_01_in17 = reg_0534;
    84: op1_01_in17 = reg_0657;
    85: op1_01_in17 = imem01_in[119:116];
    86: op1_01_in17 = imem07_in[59:56];
    87: op1_01_in17 = reg_0619;
    88: op1_01_in17 = imem01_in[123:120];
    89: op1_01_in17 = reg_0512;
    90: op1_01_in17 = reg_0084;
    92: op1_01_in17 = reg_0216;
    93: op1_01_in17 = reg_0403;
    94: op1_01_in17 = reg_0398;
    95: op1_01_in17 = reg_0623;
    96: op1_01_in17 = reg_0678;
    default: op1_01_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv17 = 1;
    6: op1_01_inv17 = 1;
    14: op1_01_inv17 = 1;
    15: op1_01_inv17 = 1;
    16: op1_01_inv17 = 1;
    17: op1_01_inv17 = 1;
    20: op1_01_inv17 = 1;
    21: op1_01_inv17 = 1;
    22: op1_01_inv17 = 1;
    23: op1_01_inv17 = 1;
    24: op1_01_inv17 = 1;
    26: op1_01_inv17 = 1;
    27: op1_01_inv17 = 1;
    28: op1_01_inv17 = 1;
    31: op1_01_inv17 = 1;
    32: op1_01_inv17 = 1;
    34: op1_01_inv17 = 1;
    38: op1_01_inv17 = 1;
    40: op1_01_inv17 = 1;
    41: op1_01_inv17 = 1;
    45: op1_01_inv17 = 1;
    47: op1_01_inv17 = 1;
    49: op1_01_inv17 = 1;
    50: op1_01_inv17 = 1;
    55: op1_01_inv17 = 1;
    56: op1_01_inv17 = 1;
    57: op1_01_inv17 = 1;
    58: op1_01_inv17 = 1;
    60: op1_01_inv17 = 1;
    65: op1_01_inv17 = 1;
    66: op1_01_inv17 = 1;
    68: op1_01_inv17 = 1;
    75: op1_01_inv17 = 1;
    82: op1_01_inv17 = 1;
    84: op1_01_inv17 = 1;
    85: op1_01_inv17 = 1;
    86: op1_01_inv17 = 1;
    87: op1_01_inv17 = 1;
    89: op1_01_inv17 = 1;
    92: op1_01_inv17 = 1;
    95: op1_01_inv17 = 1;
    default: op1_01_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in18 = imem02_in[75:72];
    5: op1_01_in18 = reg_0434;
    6: op1_01_in18 = imem03_in[3:0];
    7: op1_01_in18 = reg_0405;
    8: op1_01_in18 = imem01_in[63:60];
    9: op1_01_in18 = reg_0598;
    10: op1_01_in18 = reg_0319;
    11: op1_01_in18 = reg_0188;
    12: op1_01_in18 = reg_0329;
    13: op1_01_in18 = reg_0172;
    14: op1_01_in18 = imem02_in[51:48];
    15: op1_01_in18 = reg_0602;
    16: op1_01_in18 = reg_0155;
    17: op1_01_in18 = imem01_in[3:0];
    19: op1_01_in18 = reg_0208;
    20: op1_01_in18 = reg_0279;
    21: op1_01_in18 = imem01_in[39:36];
    22: op1_01_in18 = reg_0540;
    23: op1_01_in18 = reg_0722;
    24: op1_01_in18 = reg_0003;
    25: op1_01_in18 = reg_0154;
    26: op1_01_in18 = reg_0586;
    27: op1_01_in18 = reg_0614;
    28: op1_01_in18 = reg_0496;
    29: op1_01_in18 = reg_0662;
    30: op1_01_in18 = imem06_in[35:32];
    31: op1_01_in18 = reg_0193;
    32: op1_01_in18 = reg_0354;
    33: op1_01_in18 = imem03_in[51:48];
    34: op1_01_in18 = imem01_in[55:52];
    36: op1_01_in18 = reg_0205;
    37: op1_01_in18 = reg_0092;
    76: op1_01_in18 = reg_0092;
    38: op1_01_in18 = reg_0643;
    39: op1_01_in18 = reg_0257;
    40: op1_01_in18 = imem04_in[43:40];
    41: op1_01_in18 = reg_0440;
    42: op1_01_in18 = reg_0199;
    81: op1_01_in18 = reg_0199;
    43: op1_01_in18 = reg_0361;
    44: op1_01_in18 = imem05_in[3:0];
    45: op1_01_in18 = reg_0051;
    46: op1_01_in18 = reg_0324;
    61: op1_01_in18 = reg_0324;
    47: op1_01_in18 = reg_0803;
    48: op1_01_in18 = reg_0726;
    49: op1_01_in18 = reg_0157;
    65: op1_01_in18 = reg_0157;
    50: op1_01_in18 = imem07_in[19:16];
    84: op1_01_in18 = imem07_in[19:16];
    51: op1_01_in18 = reg_0513;
    52: op1_01_in18 = reg_0629;
    53: op1_01_in18 = reg_0276;
    54: op1_01_in18 = imem06_in[67:64];
    56: op1_01_in18 = reg_0194;
    57: op1_01_in18 = imem01_in[35:32];
    58: op1_01_in18 = reg_0166;
    59: op1_01_in18 = imem03_in[15:12];
    60: op1_01_in18 = imem01_in[107:104];
    62: op1_01_in18 = reg_0099;
    63: op1_01_in18 = imem07_in[95:92];
    64: op1_01_in18 = reg_0442;
    66: op1_01_in18 = reg_0448;
    68: op1_01_in18 = imem04_in[67:64];
    69: op1_01_in18 = imem06_in[95:92];
    70: op1_01_in18 = reg_0211;
    71: op1_01_in18 = imem06_in[51:48];
    74: op1_01_in18 = imem01_in[15:12];
    75: op1_01_in18 = imem03_in[111:108];
    77: op1_01_in18 = reg_0792;
    79: op1_01_in18 = reg_0436;
    80: op1_01_in18 = reg_0102;
    82: op1_01_in18 = reg_0238;
    83: op1_01_in18 = reg_0179;
    85: op1_01_in18 = reg_0336;
    86: op1_01_in18 = imem07_in[123:120];
    87: op1_01_in18 = reg_0404;
    88: op1_01_in18 = reg_0760;
    89: op1_01_in18 = reg_0657;
    90: op1_01_in18 = reg_0267;
    92: op1_01_in18 = imem04_in[3:0];
    93: op1_01_in18 = reg_0490;
    94: op1_01_in18 = reg_0607;
    95: op1_01_in18 = reg_0418;
    96: op1_01_in18 = imem02_in[11:8];
    default: op1_01_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv18 = 1;
    5: op1_01_inv18 = 1;
    6: op1_01_inv18 = 1;
    8: op1_01_inv18 = 1;
    9: op1_01_inv18 = 1;
    11: op1_01_inv18 = 1;
    13: op1_01_inv18 = 1;
    14: op1_01_inv18 = 1;
    17: op1_01_inv18 = 1;
    19: op1_01_inv18 = 1;
    22: op1_01_inv18 = 1;
    25: op1_01_inv18 = 1;
    29: op1_01_inv18 = 1;
    30: op1_01_inv18 = 1;
    31: op1_01_inv18 = 1;
    37: op1_01_inv18 = 1;
    39: op1_01_inv18 = 1;
    42: op1_01_inv18 = 1;
    43: op1_01_inv18 = 1;
    48: op1_01_inv18 = 1;
    49: op1_01_inv18 = 1;
    51: op1_01_inv18 = 1;
    52: op1_01_inv18 = 1;
    53: op1_01_inv18 = 1;
    57: op1_01_inv18 = 1;
    59: op1_01_inv18 = 1;
    60: op1_01_inv18 = 1;
    61: op1_01_inv18 = 1;
    63: op1_01_inv18 = 1;
    66: op1_01_inv18 = 1;
    69: op1_01_inv18 = 1;
    70: op1_01_inv18 = 1;
    75: op1_01_inv18 = 1;
    79: op1_01_inv18 = 1;
    82: op1_01_inv18 = 1;
    87: op1_01_inv18 = 1;
    88: op1_01_inv18 = 1;
    89: op1_01_inv18 = 1;
    92: op1_01_inv18 = 1;
    94: op1_01_inv18 = 1;
    96: op1_01_inv18 = 1;
    default: op1_01_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in19 = reg_0658;
    5: op1_01_in19 = reg_0437;
    41: op1_01_in19 = reg_0437;
    6: op1_01_in19 = imem03_in[75:72];
    7: op1_01_in19 = reg_0404;
    8: op1_01_in19 = imem01_in[71:68];
    9: op1_01_in19 = reg_0586;
    10: op1_01_in19 = reg_0398;
    11: op1_01_in19 = reg_0207;
    12: op1_01_in19 = reg_0353;
    13: op1_01_in19 = reg_0181;
    14: op1_01_in19 = imem02_in[111:108];
    15: op1_01_in19 = reg_0579;
    16: op1_01_in19 = imem06_in[31:28];
    17: op1_01_in19 = imem01_in[75:72];
    19: op1_01_in19 = reg_0210;
    20: op1_01_in19 = reg_0733;
    21: op1_01_in19 = imem01_in[63:60];
    22: op1_01_in19 = reg_0531;
    23: op1_01_in19 = reg_0716;
    24: op1_01_in19 = reg_0014;
    25: op1_01_in19 = reg_0139;
    26: op1_01_in19 = reg_0572;
    27: op1_01_in19 = reg_0624;
    28: op1_01_in19 = reg_0759;
    29: op1_01_in19 = reg_0636;
    30: op1_01_in19 = imem06_in[67:64];
    31: op1_01_in19 = reg_0198;
    70: op1_01_in19 = reg_0198;
    32: op1_01_in19 = reg_0341;
    33: op1_01_in19 = reg_0587;
    34: op1_01_in19 = imem01_in[83:80];
    36: op1_01_in19 = imem01_in[11:8];
    37: op1_01_in19 = reg_0314;
    38: op1_01_in19 = reg_0652;
    39: op1_01_in19 = reg_0253;
    40: op1_01_in19 = imem04_in[63:60];
    42: op1_01_in19 = reg_0197;
    43: op1_01_in19 = reg_0342;
    44: op1_01_in19 = imem05_in[51:48];
    45: op1_01_in19 = reg_0239;
    79: op1_01_in19 = reg_0239;
    46: op1_01_in19 = reg_0347;
    47: op1_01_in19 = reg_0007;
    48: op1_01_in19 = reg_0709;
    49: op1_01_in19 = reg_0158;
    50: op1_01_in19 = imem07_in[23:20];
    51: op1_01_in19 = reg_0065;
    52: op1_01_in19 = imem05_in[63:60];
    53: op1_01_in19 = reg_0224;
    54: op1_01_in19 = imem06_in[83:80];
    56: op1_01_in19 = reg_0213;
    57: op1_01_in19 = imem01_in[99:96];
    59: op1_01_in19 = imem03_in[19:16];
    60: op1_01_in19 = reg_0741;
    85: op1_01_in19 = reg_0741;
    61: op1_01_in19 = reg_0770;
    62: op1_01_in19 = reg_0304;
    63: op1_01_in19 = reg_0710;
    64: op1_01_in19 = reg_0448;
    65: op1_01_in19 = reg_0173;
    66: op1_01_in19 = reg_0435;
    68: op1_01_in19 = imem04_in[83:80];
    69: op1_01_in19 = reg_0814;
    71: op1_01_in19 = imem06_in[63:60];
    74: op1_01_in19 = imem01_in[31:28];
    75: op1_01_in19 = imem03_in[119:116];
    76: op1_01_in19 = imem03_in[7:4];
    77: op1_01_in19 = reg_0144;
    80: op1_01_in19 = reg_0241;
    81: op1_01_in19 = imem01_in[51:48];
    82: op1_01_in19 = reg_0260;
    83: op1_01_in19 = reg_0536;
    84: op1_01_in19 = imem07_in[79:76];
    86: op1_01_in19 = imem07_in[127:124];
    87: op1_01_in19 = reg_0168;
    88: op1_01_in19 = reg_0225;
    89: op1_01_in19 = reg_0680;
    90: op1_01_in19 = reg_0268;
    92: op1_01_in19 = imem04_in[15:12];
    93: op1_01_in19 = reg_0562;
    94: op1_01_in19 = reg_0001;
    95: op1_01_in19 = reg_0278;
    96: op1_01_in19 = imem02_in[31:28];
    default: op1_01_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_01_inv19 = 1;
    8: op1_01_inv19 = 1;
    9: op1_01_inv19 = 1;
    10: op1_01_inv19 = 1;
    12: op1_01_inv19 = 1;
    13: op1_01_inv19 = 1;
    14: op1_01_inv19 = 1;
    15: op1_01_inv19 = 1;
    17: op1_01_inv19 = 1;
    19: op1_01_inv19 = 1;
    21: op1_01_inv19 = 1;
    26: op1_01_inv19 = 1;
    27: op1_01_inv19 = 1;
    28: op1_01_inv19 = 1;
    33: op1_01_inv19 = 1;
    36: op1_01_inv19 = 1;
    38: op1_01_inv19 = 1;
    39: op1_01_inv19 = 1;
    40: op1_01_inv19 = 1;
    47: op1_01_inv19 = 1;
    52: op1_01_inv19 = 1;
    53: op1_01_inv19 = 1;
    56: op1_01_inv19 = 1;
    61: op1_01_inv19 = 1;
    63: op1_01_inv19 = 1;
    64: op1_01_inv19 = 1;
    66: op1_01_inv19 = 1;
    69: op1_01_inv19 = 1;
    70: op1_01_inv19 = 1;
    71: op1_01_inv19 = 1;
    79: op1_01_inv19 = 1;
    81: op1_01_inv19 = 1;
    83: op1_01_inv19 = 1;
    84: op1_01_inv19 = 1;
    85: op1_01_inv19 = 1;
    86: op1_01_inv19 = 1;
    87: op1_01_inv19 = 1;
    90: op1_01_inv19 = 1;
    92: op1_01_inv19 = 1;
    96: op1_01_inv19 = 1;
    default: op1_01_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in20 = reg_0646;
    5: op1_01_in20 = reg_0438;
    41: op1_01_in20 = reg_0438;
    6: op1_01_in20 = imem03_in[107:104];
    7: op1_01_in20 = reg_0406;
    8: op1_01_in20 = imem01_in[75:72];
    81: op1_01_in20 = imem01_in[75:72];
    9: op1_01_in20 = reg_0582;
    75: op1_01_in20 = reg_0582;
    10: op1_01_in20 = reg_0374;
    11: op1_01_in20 = reg_0201;
    12: op1_01_in20 = reg_0342;
    13: op1_01_in20 = reg_0169;
    14: op1_01_in20 = reg_0650;
    15: op1_01_in20 = reg_0563;
    16: op1_01_in20 = imem06_in[79:76];
    17: op1_01_in20 = imem01_in[115:112];
    19: op1_01_in20 = reg_0189;
    20: op1_01_in20 = reg_0282;
    21: op1_01_in20 = imem01_in[103:100];
    22: op1_01_in20 = reg_0538;
    23: op1_01_in20 = reg_0704;
    24: op1_01_in20 = reg_0809;
    25: op1_01_in20 = reg_0138;
    26: op1_01_in20 = reg_0569;
    27: op1_01_in20 = reg_0617;
    28: op1_01_in20 = reg_0760;
    29: op1_01_in20 = reg_0324;
    30: op1_01_in20 = reg_0605;
    31: op1_01_in20 = imem01_in[3:0];
    32: op1_01_in20 = reg_0321;
    33: op1_01_in20 = reg_0589;
    34: op1_01_in20 = imem01_in[107:104];
    36: op1_01_in20 = imem01_in[39:36];
    74: op1_01_in20 = imem01_in[39:36];
    37: op1_01_in20 = reg_0080;
    46: op1_01_in20 = reg_0080;
    38: op1_01_in20 = reg_0352;
    39: op1_01_in20 = reg_0066;
    40: op1_01_in20 = imem04_in[71:68];
    42: op1_01_in20 = imem01_in[23:20];
    43: op1_01_in20 = reg_0350;
    44: op1_01_in20 = imem05_in[63:60];
    45: op1_01_in20 = reg_0434;
    47: op1_01_in20 = reg_0804;
    48: op1_01_in20 = reg_0067;
    50: op1_01_in20 = imem07_in[39:36];
    51: op1_01_in20 = reg_0507;
    52: op1_01_in20 = imem05_in[103:100];
    53: op1_01_in20 = reg_0249;
    54: op1_01_in20 = imem06_in[103:100];
    56: op1_01_in20 = reg_0199;
    57: op1_01_in20 = imem01_in[119:116];
    59: op1_01_in20 = imem03_in[47:44];
    60: op1_01_in20 = reg_0550;
    61: op1_01_in20 = reg_0098;
    62: op1_01_in20 = reg_0256;
    63: op1_01_in20 = reg_0731;
    64: op1_01_in20 = reg_0435;
    66: op1_01_in20 = reg_0268;
    68: op1_01_in20 = imem04_in[95:92];
    69: op1_01_in20 = reg_0618;
    70: op1_01_in20 = reg_0202;
    71: op1_01_in20 = imem06_in[67:64];
    76: op1_01_in20 = imem03_in[67:64];
    77: op1_01_in20 = reg_0386;
    79: op1_01_in20 = reg_0440;
    80: op1_01_in20 = reg_0574;
    82: op1_01_in20 = reg_0031;
    83: op1_01_in20 = reg_0510;
    84: op1_01_in20 = imem07_in[107:104];
    85: op1_01_in20 = reg_0394;
    86: op1_01_in20 = reg_0726;
    87: op1_01_in20 = reg_0578;
    88: op1_01_in20 = reg_0232;
    89: op1_01_in20 = imem07_in[19:16];
    90: op1_01_in20 = reg_0182;
    92: op1_01_in20 = imem04_in[35:32];
    93: op1_01_in20 = reg_0557;
    94: op1_01_in20 = reg_0002;
    95: op1_01_in20 = reg_0806;
    96: op1_01_in20 = imem02_in[79:76];
    default: op1_01_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv20 = 1;
    6: op1_01_inv20 = 1;
    7: op1_01_inv20 = 1;
    8: op1_01_inv20 = 1;
    9: op1_01_inv20 = 1;
    14: op1_01_inv20 = 1;
    19: op1_01_inv20 = 1;
    20: op1_01_inv20 = 1;
    21: op1_01_inv20 = 1;
    22: op1_01_inv20 = 1;
    28: op1_01_inv20 = 1;
    31: op1_01_inv20 = 1;
    32: op1_01_inv20 = 1;
    33: op1_01_inv20 = 1;
    34: op1_01_inv20 = 1;
    36: op1_01_inv20 = 1;
    37: op1_01_inv20 = 1;
    39: op1_01_inv20 = 1;
    42: op1_01_inv20 = 1;
    43: op1_01_inv20 = 1;
    44: op1_01_inv20 = 1;
    45: op1_01_inv20 = 1;
    46: op1_01_inv20 = 1;
    47: op1_01_inv20 = 1;
    48: op1_01_inv20 = 1;
    50: op1_01_inv20 = 1;
    52: op1_01_inv20 = 1;
    54: op1_01_inv20 = 1;
    57: op1_01_inv20 = 1;
    60: op1_01_inv20 = 1;
    61: op1_01_inv20 = 1;
    68: op1_01_inv20 = 1;
    69: op1_01_inv20 = 1;
    70: op1_01_inv20 = 1;
    74: op1_01_inv20 = 1;
    75: op1_01_inv20 = 1;
    76: op1_01_inv20 = 1;
    77: op1_01_inv20 = 1;
    81: op1_01_inv20 = 1;
    82: op1_01_inv20 = 1;
    83: op1_01_inv20 = 1;
    85: op1_01_inv20 = 1;
    87: op1_01_inv20 = 1;
    88: op1_01_inv20 = 1;
    89: op1_01_inv20 = 1;
    90: op1_01_inv20 = 1;
    92: op1_01_inv20 = 1;
    93: op1_01_inv20 = 1;
    95: op1_01_inv20 = 1;
    default: op1_01_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in21 = reg_0647;
    5: op1_01_in21 = reg_0162;
    41: op1_01_in21 = reg_0162;
    6: op1_01_in21 = reg_0591;
    7: op1_01_in21 = reg_0028;
    8: op1_01_in21 = imem01_in[95:92];
    9: op1_01_in21 = reg_0596;
    10: op1_01_in21 = reg_0001;
    11: op1_01_in21 = imem01_in[31:28];
    42: op1_01_in21 = imem01_in[31:28];
    12: op1_01_in21 = reg_0082;
    13: op1_01_in21 = reg_0183;
    14: op1_01_in21 = reg_0658;
    15: op1_01_in21 = reg_0576;
    16: op1_01_in21 = imem06_in[83:80];
    17: op1_01_in21 = reg_0523;
    19: op1_01_in21 = reg_0201;
    20: op1_01_in21 = reg_0272;
    21: op1_01_in21 = imem01_in[107:104];
    22: op1_01_in21 = reg_0532;
    23: op1_01_in21 = reg_0721;
    24: op1_01_in21 = imem04_in[15:12];
    25: op1_01_in21 = imem06_in[23:20];
    26: op1_01_in21 = reg_0594;
    27: op1_01_in21 = reg_0621;
    28: op1_01_in21 = reg_0235;
    29: op1_01_in21 = reg_0353;
    30: op1_01_in21 = reg_0606;
    31: op1_01_in21 = imem01_in[27:24];
    32: op1_01_in21 = reg_0092;
    33: op1_01_in21 = reg_0517;
    34: op1_01_in21 = reg_0758;
    36: op1_01_in21 = imem01_in[67:64];
    37: op1_01_in21 = reg_0530;
    38: op1_01_in21 = reg_0356;
    39: op1_01_in21 = reg_0071;
    40: op1_01_in21 = imem04_in[91:88];
    43: op1_01_in21 = reg_0321;
    44: op1_01_in21 = imem05_in[71:68];
    45: op1_01_in21 = reg_0449;
    46: op1_01_in21 = reg_0539;
    47: op1_01_in21 = reg_0806;
    48: op1_01_in21 = reg_0447;
    50: op1_01_in21 = imem07_in[127:124];
    51: op1_01_in21 = reg_0296;
    52: op1_01_in21 = reg_0792;
    53: op1_01_in21 = reg_0101;
    54: op1_01_in21 = imem06_in[107:104];
    56: op1_01_in21 = imem01_in[47:44];
    57: op1_01_in21 = reg_0646;
    59: op1_01_in21 = imem03_in[87:84];
    60: op1_01_in21 = reg_0760;
    61: op1_01_in21 = reg_0757;
    62: op1_01_in21 = reg_0742;
    63: op1_01_in21 = reg_0725;
    64: op1_01_in21 = reg_0268;
    66: op1_01_in21 = reg_0180;
    68: op1_01_in21 = imem04_in[107:104];
    69: op1_01_in21 = reg_0659;
    70: op1_01_in21 = imem01_in[15:12];
    71: op1_01_in21 = imem06_in[95:92];
    74: op1_01_in21 = imem01_in[63:60];
    75: op1_01_in21 = reg_0750;
    76: op1_01_in21 = imem03_in[119:116];
    77: op1_01_in21 = reg_0246;
    79: op1_01_in21 = reg_0181;
    80: op1_01_in21 = reg_0054;
    81: op1_01_in21 = imem01_in[79:76];
    82: op1_01_in21 = reg_0405;
    83: op1_01_in21 = reg_0516;
    84: op1_01_in21 = reg_0159;
    85: op1_01_in21 = reg_0507;
    86: op1_01_in21 = reg_0382;
    87: op1_01_in21 = reg_0408;
    88: op1_01_in21 = reg_0216;
    89: op1_01_in21 = imem07_in[31:28];
    92: op1_01_in21 = imem04_in[51:48];
    93: op1_01_in21 = reg_0248;
    94: op1_01_in21 = reg_0418;
    95: op1_01_in21 = reg_0809;
    96: op1_01_in21 = imem02_in[95:92];
    default: op1_01_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    12: op1_01_inv21 = 1;
    13: op1_01_inv21 = 1;
    14: op1_01_inv21 = 1;
    20: op1_01_inv21 = 1;
    22: op1_01_inv21 = 1;
    24: op1_01_inv21 = 1;
    28: op1_01_inv21 = 1;
    29: op1_01_inv21 = 1;
    32: op1_01_inv21 = 1;
    33: op1_01_inv21 = 1;
    34: op1_01_inv21 = 1;
    36: op1_01_inv21 = 1;
    37: op1_01_inv21 = 1;
    39: op1_01_inv21 = 1;
    40: op1_01_inv21 = 1;
    46: op1_01_inv21 = 1;
    54: op1_01_inv21 = 1;
    56: op1_01_inv21 = 1;
    57: op1_01_inv21 = 1;
    59: op1_01_inv21 = 1;
    62: op1_01_inv21 = 1;
    63: op1_01_inv21 = 1;
    64: op1_01_inv21 = 1;
    66: op1_01_inv21 = 1;
    68: op1_01_inv21 = 1;
    70: op1_01_inv21 = 1;
    76: op1_01_inv21 = 1;
    80: op1_01_inv21 = 1;
    81: op1_01_inv21 = 1;
    84: op1_01_inv21 = 1;
    85: op1_01_inv21 = 1;
    89: op1_01_inv21 = 1;
    95: op1_01_inv21 = 1;
    default: op1_01_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in22 = reg_0648;
    5: op1_01_in22 = reg_0163;
    6: op1_01_in22 = reg_0589;
    7: op1_01_in22 = reg_0037;
    8: op1_01_in22 = reg_0506;
    9: op1_01_in22 = reg_0583;
    10: op1_01_in22 = reg_0808;
    11: op1_01_in22 = imem01_in[39:36];
    12: op1_01_in22 = imem03_in[71:68];
    13: op1_01_in22 = reg_0166;
    14: op1_01_in22 = reg_0653;
    15: op1_01_in22 = reg_0394;
    16: op1_01_in22 = imem06_in[91:88];
    17: op1_01_in22 = reg_0822;
    19: op1_01_in22 = reg_0213;
    20: op1_01_in22 = reg_0277;
    21: op1_01_in22 = reg_0523;
    22: op1_01_in22 = imem03_in[23:20];
    61: op1_01_in22 = imem03_in[23:20];
    23: op1_01_in22 = reg_0713;
    24: op1_01_in22 = imem04_in[19:16];
    25: op1_01_in22 = imem06_in[59:56];
    26: op1_01_in22 = reg_0597;
    27: op1_01_in22 = reg_0611;
    28: op1_01_in22 = reg_0215;
    29: op1_01_in22 = reg_0073;
    30: op1_01_in22 = reg_0609;
    31: op1_01_in22 = imem01_in[107:104];
    32: op1_01_in22 = reg_0743;
    33: op1_01_in22 = reg_0001;
    34: op1_01_in22 = reg_0336;
    36: op1_01_in22 = imem01_in[111:108];
    37: op1_01_in22 = reg_0526;
    38: op1_01_in22 = reg_0353;
    39: op1_01_in22 = reg_0075;
    40: op1_01_in22 = imem04_in[107:104];
    41: op1_01_in22 = reg_0168;
    42: op1_01_in22 = imem01_in[51:48];
    43: op1_01_in22 = reg_0095;
    44: op1_01_in22 = imem05_in[75:72];
    45: op1_01_in22 = reg_0268;
    46: op1_01_in22 = reg_0756;
    47: op1_01_in22 = imem04_in[11:8];
    48: op1_01_in22 = reg_0434;
    50: op1_01_in22 = reg_0728;
    51: op1_01_in22 = reg_0519;
    52: op1_01_in22 = reg_0099;
    53: op1_01_in22 = reg_0130;
    54: op1_01_in22 = imem06_in[123:120];
    56: op1_01_in22 = imem01_in[55:52];
    57: op1_01_in22 = reg_0735;
    59: op1_01_in22 = imem03_in[95:92];
    60: op1_01_in22 = reg_0248;
    62: op1_01_in22 = reg_0066;
    63: op1_01_in22 = reg_0712;
    64: op1_01_in22 = reg_0180;
    66: op1_01_in22 = reg_0164;
    68: op1_01_in22 = imem04_in[115:112];
    69: op1_01_in22 = reg_0816;
    70: op1_01_in22 = imem01_in[31:28];
    71: op1_01_in22 = imem06_in[103:100];
    74: op1_01_in22 = imem01_in[71:68];
    75: op1_01_in22 = reg_0600;
    76: op1_01_in22 = imem03_in[123:120];
    77: op1_01_in22 = reg_0150;
    79: op1_01_in22 = reg_0184;
    80: op1_01_in22 = reg_0240;
    81: op1_01_in22 = imem01_in[99:96];
    82: op1_01_in22 = reg_0375;
    83: op1_01_in22 = reg_0556;
    84: op1_01_in22 = reg_0382;
    85: op1_01_in22 = reg_0225;
    86: op1_01_in22 = reg_0789;
    87: op1_01_in22 = reg_0775;
    88: op1_01_in22 = reg_0294;
    89: op1_01_in22 = imem07_in[43:40];
    92: op1_01_in22 = imem04_in[55:52];
    93: op1_01_in22 = reg_0319;
    94: op1_01_in22 = reg_0368;
    95: op1_01_in22 = imem04_in[7:4];
    96: op1_01_in22 = imem02_in[119:116];
    default: op1_01_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_01_inv22 = 1;
    8: op1_01_inv22 = 1;
    9: op1_01_inv22 = 1;
    10: op1_01_inv22 = 1;
    12: op1_01_inv22 = 1;
    15: op1_01_inv22 = 1;
    16: op1_01_inv22 = 1;
    19: op1_01_inv22 = 1;
    20: op1_01_inv22 = 1;
    21: op1_01_inv22 = 1;
    22: op1_01_inv22 = 1;
    23: op1_01_inv22 = 1;
    24: op1_01_inv22 = 1;
    26: op1_01_inv22 = 1;
    27: op1_01_inv22 = 1;
    31: op1_01_inv22 = 1;
    36: op1_01_inv22 = 1;
    38: op1_01_inv22 = 1;
    40: op1_01_inv22 = 1;
    41: op1_01_inv22 = 1;
    43: op1_01_inv22 = 1;
    47: op1_01_inv22 = 1;
    50: op1_01_inv22 = 1;
    51: op1_01_inv22 = 1;
    59: op1_01_inv22 = 1;
    60: op1_01_inv22 = 1;
    62: op1_01_inv22 = 1;
    64: op1_01_inv22 = 1;
    66: op1_01_inv22 = 1;
    70: op1_01_inv22 = 1;
    74: op1_01_inv22 = 1;
    76: op1_01_inv22 = 1;
    77: op1_01_inv22 = 1;
    80: op1_01_inv22 = 1;
    82: op1_01_inv22 = 1;
    84: op1_01_inv22 = 1;
    85: op1_01_inv22 = 1;
    86: op1_01_inv22 = 1;
    87: op1_01_inv22 = 1;
    88: op1_01_inv22 = 1;
    89: op1_01_inv22 = 1;
    92: op1_01_inv22 = 1;
    93: op1_01_inv22 = 1;
    94: op1_01_inv22 = 1;
    95: op1_01_inv22 = 1;
    default: op1_01_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in23 = reg_0649;
    5: op1_01_in23 = reg_0168;
    6: op1_01_in23 = reg_0593;
    7: op1_01_in23 = reg_0029;
    8: op1_01_in23 = reg_0510;
    9: op1_01_in23 = reg_0585;
    10: op1_01_in23 = reg_0803;
    11: op1_01_in23 = imem01_in[71:68];
    42: op1_01_in23 = imem01_in[71:68];
    12: op1_01_in23 = reg_0598;
    13: op1_01_in23 = reg_0157;
    41: op1_01_in23 = reg_0157;
    14: op1_01_in23 = reg_0654;
    15: op1_01_in23 = reg_0362;
    16: op1_01_in23 = reg_0613;
    17: op1_01_in23 = reg_0755;
    19: op1_01_in23 = reg_0190;
    20: op1_01_in23 = reg_0285;
    21: op1_01_in23 = reg_0520;
    22: op1_01_in23 = imem03_in[43:40];
    23: op1_01_in23 = reg_0430;
    24: op1_01_in23 = imem04_in[51:48];
    25: op1_01_in23 = imem06_in[119:116];
    26: op1_01_in23 = reg_0570;
    27: op1_01_in23 = reg_0633;
    28: op1_01_in23 = reg_0244;
    29: op1_01_in23 = reg_0096;
    30: op1_01_in23 = reg_0618;
    31: op1_01_in23 = imem01_in[119:116];
    32: op1_01_in23 = reg_0540;
    33: op1_01_in23 = reg_0008;
    34: op1_01_in23 = reg_0497;
    36: op1_01_in23 = imem01_in[115:112];
    37: op1_01_in23 = reg_0538;
    38: op1_01_in23 = reg_0322;
    39: op1_01_in23 = imem05_in[83:80];
    40: op1_01_in23 = imem04_in[111:108];
    43: op1_01_in23 = reg_0530;
    44: op1_01_in23 = reg_0798;
    45: op1_01_in23 = reg_0181;
    46: op1_01_in23 = reg_0531;
    47: op1_01_in23 = imem04_in[55:52];
    48: op1_01_in23 = reg_0158;
    84: op1_01_in23 = reg_0158;
    50: op1_01_in23 = reg_0716;
    51: op1_01_in23 = reg_0233;
    52: op1_01_in23 = reg_0070;
    53: op1_01_in23 = imem06_in[3:0];
    54: op1_01_in23 = reg_0218;
    56: op1_01_in23 = imem01_in[75:72];
    57: op1_01_in23 = reg_0653;
    59: op1_01_in23 = reg_0602;
    60: op1_01_in23 = reg_0506;
    61: op1_01_in23 = imem03_in[39:36];
    62: op1_01_in23 = reg_0153;
    63: op1_01_in23 = reg_0705;
    64: op1_01_in23 = reg_0160;
    66: op1_01_in23 = reg_0185;
    68: op1_01_in23 = reg_0544;
    69: op1_01_in23 = reg_0638;
    70: op1_01_in23 = imem01_in[63:60];
    71: op1_01_in23 = reg_0815;
    74: op1_01_in23 = imem01_in[87:84];
    75: op1_01_in23 = reg_0595;
    76: op1_01_in23 = reg_0063;
    77: op1_01_in23 = reg_0143;
    80: op1_01_in23 = reg_0420;
    81: op1_01_in23 = imem01_in[107:104];
    82: op1_01_in23 = reg_0583;
    83: op1_01_in23 = reg_0432;
    85: op1_01_in23 = reg_0232;
    86: op1_01_in23 = reg_0724;
    87: op1_01_in23 = reg_0484;
    88: op1_01_in23 = reg_0219;
    89: op1_01_in23 = imem07_in[67:64];
    92: op1_01_in23 = imem04_in[59:56];
    93: op1_01_in23 = imem04_in[7:4];
    94: op1_01_in23 = reg_0319;
    95: op1_01_in23 = imem04_in[15:12];
    96: op1_01_in23 = reg_0057;
    default: op1_01_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv23 = 1;
    13: op1_01_inv23 = 1;
    15: op1_01_inv23 = 1;
    16: op1_01_inv23 = 1;
    21: op1_01_inv23 = 1;
    22: op1_01_inv23 = 1;
    23: op1_01_inv23 = 1;
    24: op1_01_inv23 = 1;
    27: op1_01_inv23 = 1;
    28: op1_01_inv23 = 1;
    32: op1_01_inv23 = 1;
    34: op1_01_inv23 = 1;
    36: op1_01_inv23 = 1;
    37: op1_01_inv23 = 1;
    38: op1_01_inv23 = 1;
    39: op1_01_inv23 = 1;
    41: op1_01_inv23 = 1;
    47: op1_01_inv23 = 1;
    52: op1_01_inv23 = 1;
    54: op1_01_inv23 = 1;
    56: op1_01_inv23 = 1;
    57: op1_01_inv23 = 1;
    59: op1_01_inv23 = 1;
    63: op1_01_inv23 = 1;
    64: op1_01_inv23 = 1;
    69: op1_01_inv23 = 1;
    70: op1_01_inv23 = 1;
    80: op1_01_inv23 = 1;
    82: op1_01_inv23 = 1;
    83: op1_01_inv23 = 1;
    84: op1_01_inv23 = 1;
    86: op1_01_inv23 = 1;
    87: op1_01_inv23 = 1;
    88: op1_01_inv23 = 1;
    89: op1_01_inv23 = 1;
    92: op1_01_inv23 = 1;
    94: op1_01_inv23 = 1;
    95: op1_01_inv23 = 1;
    96: op1_01_inv23 = 1;
    default: op1_01_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in24 = reg_0659;
    5: op1_01_in24 = reg_0170;
    6: op1_01_in24 = reg_0580;
    9: op1_01_in24 = reg_0580;
    7: op1_01_in24 = reg_0038;
    8: op1_01_in24 = reg_0232;
    10: op1_01_in24 = reg_0014;
    11: op1_01_in24 = imem01_in[95:92];
    12: op1_01_in24 = reg_0602;
    13: op1_01_in24 = reg_0173;
    48: op1_01_in24 = reg_0173;
    14: op1_01_in24 = reg_0656;
    15: op1_01_in24 = reg_0373;
    16: op1_01_in24 = reg_0605;
    54: op1_01_in24 = reg_0605;
    17: op1_01_in24 = reg_0235;
    19: op1_01_in24 = imem01_in[51:48];
    20: op1_01_in24 = reg_0089;
    21: op1_01_in24 = reg_0514;
    22: op1_01_in24 = imem03_in[83:80];
    61: op1_01_in24 = imem03_in[83:80];
    23: op1_01_in24 = reg_0419;
    24: op1_01_in24 = imem04_in[67:64];
    92: op1_01_in24 = imem04_in[67:64];
    25: op1_01_in24 = imem06_in[127:124];
    26: op1_01_in24 = reg_0394;
    27: op1_01_in24 = reg_0618;
    28: op1_01_in24 = reg_0220;
    29: op1_01_in24 = reg_0770;
    30: op1_01_in24 = reg_0627;
    31: op1_01_in24 = reg_0337;
    32: op1_01_in24 = reg_0094;
    37: op1_01_in24 = reg_0094;
    33: op1_01_in24 = reg_0015;
    34: op1_01_in24 = reg_0520;
    36: op1_01_in24 = imem01_in[119:116];
    74: op1_01_in24 = imem01_in[119:116];
    38: op1_01_in24 = reg_0343;
    39: op1_01_in24 = reg_0792;
    40: op1_01_in24 = reg_0553;
    42: op1_01_in24 = imem01_in[87:84];
    43: op1_01_in24 = reg_0498;
    44: op1_01_in24 = reg_0483;
    45: op1_01_in24 = reg_0161;
    46: op1_01_in24 = reg_0532;
    47: op1_01_in24 = imem04_in[59:56];
    50: op1_01_in24 = reg_0710;
    51: op1_01_in24 = imem05_in[7:4];
    52: op1_01_in24 = reg_0269;
    53: op1_01_in24 = imem06_in[11:8];
    56: op1_01_in24 = imem01_in[99:96];
    57: op1_01_in24 = reg_0778;
    59: op1_01_in24 = reg_0582;
    60: op1_01_in24 = reg_0124;
    80: op1_01_in24 = reg_0124;
    62: op1_01_in24 = imem06_in[3:0];
    63: op1_01_in24 = reg_0706;
    64: op1_01_in24 = reg_0185;
    66: op1_01_in24 = reg_0176;
    68: op1_01_in24 = reg_0560;
    69: op1_01_in24 = reg_0764;
    70: op1_01_in24 = imem01_in[79:76];
    71: op1_01_in24 = reg_0354;
    75: op1_01_in24 = reg_0509;
    76: op1_01_in24 = reg_0597;
    77: op1_01_in24 = reg_0783;
    81: op1_01_in24 = reg_0085;
    82: op1_01_in24 = reg_0035;
    83: op1_01_in24 = reg_0079;
    84: op1_01_in24 = reg_0727;
    85: op1_01_in24 = reg_0241;
    86: op1_01_in24 = reg_0103;
    87: op1_01_in24 = reg_0661;
    88: op1_01_in24 = reg_0073;
    89: op1_01_in24 = reg_0726;
    93: op1_01_in24 = imem04_in[19:16];
    94: op1_01_in24 = reg_0278;
    95: op1_01_in24 = imem04_in[27:24];
    96: op1_01_in24 = reg_0081;
    default: op1_01_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv24 = 1;
    5: op1_01_inv24 = 1;
    8: op1_01_inv24 = 1;
    11: op1_01_inv24 = 1;
    14: op1_01_inv24 = 1;
    16: op1_01_inv24 = 1;
    20: op1_01_inv24 = 1;
    21: op1_01_inv24 = 1;
    23: op1_01_inv24 = 1;
    24: op1_01_inv24 = 1;
    25: op1_01_inv24 = 1;
    32: op1_01_inv24 = 1;
    33: op1_01_inv24 = 1;
    36: op1_01_inv24 = 1;
    38: op1_01_inv24 = 1;
    44: op1_01_inv24 = 1;
    48: op1_01_inv24 = 1;
    50: op1_01_inv24 = 1;
    53: op1_01_inv24 = 1;
    54: op1_01_inv24 = 1;
    56: op1_01_inv24 = 1;
    59: op1_01_inv24 = 1;
    61: op1_01_inv24 = 1;
    66: op1_01_inv24 = 1;
    68: op1_01_inv24 = 1;
    77: op1_01_inv24 = 1;
    80: op1_01_inv24 = 1;
    81: op1_01_inv24 = 1;
    82: op1_01_inv24 = 1;
    83: op1_01_inv24 = 1;
    84: op1_01_inv24 = 1;
    86: op1_01_inv24 = 1;
    87: op1_01_inv24 = 1;
    88: op1_01_inv24 = 1;
    92: op1_01_inv24 = 1;
    94: op1_01_inv24 = 1;
    96: op1_01_inv24 = 1;
    default: op1_01_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in25 = reg_0320;
    5: op1_01_in25 = reg_0171;
    6: op1_01_in25 = reg_0576;
    7: op1_01_in25 = imem07_in[39:36];
    8: op1_01_in25 = reg_0249;
    9: op1_01_in25 = reg_0578;
    10: op1_01_in25 = reg_0810;
    11: op1_01_in25 = imem01_in[127:124];
    12: op1_01_in25 = reg_0579;
    14: op1_01_in25 = reg_0665;
    15: op1_01_in25 = reg_0327;
    16: op1_01_in25 = reg_0611;
    17: op1_01_in25 = reg_0503;
    19: op1_01_in25 = imem01_in[71:68];
    20: op1_01_in25 = reg_0147;
    21: op1_01_in25 = reg_0820;
    34: op1_01_in25 = reg_0820;
    22: op1_01_in25 = imem03_in[99:96];
    23: op1_01_in25 = reg_0434;
    24: op1_01_in25 = imem04_in[71:68];
    47: op1_01_in25 = imem04_in[71:68];
    25: op1_01_in25 = reg_0610;
    26: op1_01_in25 = reg_0391;
    27: op1_01_in25 = reg_0632;
    28: op1_01_in25 = reg_0041;
    29: op1_01_in25 = reg_0539;
    30: op1_01_in25 = reg_0623;
    31: op1_01_in25 = reg_0514;
    32: op1_01_in25 = reg_0093;
    33: op1_01_in25 = reg_0016;
    36: op1_01_in25 = reg_0501;
    37: op1_01_in25 = imem03_in[43:40];
    38: op1_01_in25 = reg_0314;
    39: op1_01_in25 = reg_0483;
    40: op1_01_in25 = reg_0552;
    42: op1_01_in25 = imem01_in[103:100];
    43: op1_01_in25 = imem03_in[7:4];
    44: op1_01_in25 = reg_0488;
    45: op1_01_in25 = reg_0169;
    46: op1_01_in25 = imem03_in[3:0];
    50: op1_01_in25 = reg_0714;
    51: op1_01_in25 = imem05_in[11:8];
    52: op1_01_in25 = reg_0744;
    53: op1_01_in25 = imem06_in[23:20];
    54: op1_01_in25 = reg_0286;
    56: op1_01_in25 = imem01_in[111:108];
    57: op1_01_in25 = reg_0557;
    59: op1_01_in25 = reg_0599;
    60: op1_01_in25 = reg_0118;
    61: op1_01_in25 = imem03_in[91:88];
    62: op1_01_in25 = imem06_in[63:60];
    63: op1_01_in25 = reg_0266;
    66: op1_01_in25 = reg_0184;
    68: op1_01_in25 = reg_0087;
    69: op1_01_in25 = reg_0667;
    70: op1_01_in25 = imem01_in[83:80];
    71: op1_01_in25 = reg_0766;
    74: op1_01_in25 = reg_0497;
    75: op1_01_in25 = reg_0028;
    76: op1_01_in25 = reg_0559;
    77: op1_01_in25 = reg_0765;
    80: op1_01_in25 = reg_0673;
    81: op1_01_in25 = reg_0645;
    82: op1_01_in25 = reg_0512;
    83: op1_01_in25 = reg_0305;
    84: op1_01_in25 = reg_0439;
    85: op1_01_in25 = reg_0423;
    86: op1_01_in25 = reg_0436;
    87: op1_01_in25 = imem07_in[3:0];
    88: op1_01_in25 = reg_0677;
    89: op1_01_in25 = reg_0784;
    92: op1_01_in25 = imem04_in[75:72];
    93: op1_01_in25 = imem04_in[43:40];
    94: op1_01_in25 = reg_0290;
    95: op1_01_in25 = imem04_in[35:32];
    96: op1_01_in25 = reg_0753;
    default: op1_01_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_01_inv25 = 1;
    11: op1_01_inv25 = 1;
    12: op1_01_inv25 = 1;
    14: op1_01_inv25 = 1;
    20: op1_01_inv25 = 1;
    21: op1_01_inv25 = 1;
    23: op1_01_inv25 = 1;
    24: op1_01_inv25 = 1;
    25: op1_01_inv25 = 1;
    29: op1_01_inv25 = 1;
    31: op1_01_inv25 = 1;
    32: op1_01_inv25 = 1;
    37: op1_01_inv25 = 1;
    39: op1_01_inv25 = 1;
    43: op1_01_inv25 = 1;
    44: op1_01_inv25 = 1;
    45: op1_01_inv25 = 1;
    46: op1_01_inv25 = 1;
    47: op1_01_inv25 = 1;
    50: op1_01_inv25 = 1;
    51: op1_01_inv25 = 1;
    53: op1_01_inv25 = 1;
    56: op1_01_inv25 = 1;
    57: op1_01_inv25 = 1;
    59: op1_01_inv25 = 1;
    60: op1_01_inv25 = 1;
    68: op1_01_inv25 = 1;
    69: op1_01_inv25 = 1;
    70: op1_01_inv25 = 1;
    74: op1_01_inv25 = 1;
    75: op1_01_inv25 = 1;
    76: op1_01_inv25 = 1;
    77: op1_01_inv25 = 1;
    81: op1_01_inv25 = 1;
    83: op1_01_inv25 = 1;
    84: op1_01_inv25 = 1;
    86: op1_01_inv25 = 1;
    87: op1_01_inv25 = 1;
    92: op1_01_inv25 = 1;
    93: op1_01_inv25 = 1;
    94: op1_01_inv25 = 1;
    default: op1_01_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in26 = reg_0341;
    14: op1_01_in26 = reg_0341;
    6: op1_01_in26 = reg_0321;
    7: op1_01_in26 = imem07_in[43:40];
    8: op1_01_in26 = imem02_in[15:12];
    9: op1_01_in26 = reg_0394;
    10: op1_01_in26 = imem04_in[7:4];
    11: op1_01_in26 = reg_0520;
    12: op1_01_in26 = reg_0568;
    15: op1_01_in26 = reg_0000;
    16: op1_01_in26 = reg_0615;
    83: op1_01_in26 = reg_0615;
    17: op1_01_in26 = reg_0504;
    19: op1_01_in26 = imem01_in[75:72];
    20: op1_01_in26 = reg_0133;
    21: op1_01_in26 = reg_0755;
    22: op1_01_in26 = imem03_in[123:120];
    23: op1_01_in26 = reg_0446;
    24: op1_01_in26 = imem04_in[83:80];
    25: op1_01_in26 = reg_0607;
    26: op1_01_in26 = reg_0388;
    27: op1_01_in26 = reg_0408;
    28: op1_01_in26 = reg_0243;
    29: op1_01_in26 = reg_0098;
    30: op1_01_in26 = reg_0612;
    31: op1_01_in26 = reg_0825;
    32: op1_01_in26 = imem03_in[3:0];
    33: op1_01_in26 = reg_0009;
    34: op1_01_in26 = reg_0505;
    36: op1_01_in26 = reg_0550;
    37: op1_01_in26 = imem03_in[71:68];
    38: op1_01_in26 = reg_0081;
    39: op1_01_in26 = reg_0780;
    40: op1_01_in26 = reg_0087;
    42: op1_01_in26 = reg_0515;
    43: op1_01_in26 = imem03_in[27:24];
    44: op1_01_in26 = reg_0491;
    45: op1_01_in26 = reg_0178;
    46: op1_01_in26 = imem03_in[11:8];
    47: op1_01_in26 = imem04_in[99:96];
    50: op1_01_in26 = reg_0729;
    51: op1_01_in26 = imem05_in[71:68];
    52: op1_01_in26 = reg_0147;
    53: op1_01_in26 = imem06_in[67:64];
    54: op1_01_in26 = reg_0622;
    56: op1_01_in26 = reg_0653;
    57: op1_01_in26 = reg_0652;
    59: op1_01_in26 = reg_0604;
    60: op1_01_in26 = reg_0677;
    61: op1_01_in26 = imem03_in[115:112];
    62: op1_01_in26 = imem06_in[75:72];
    63: op1_01_in26 = reg_0295;
    68: op1_01_in26 = reg_0056;
    69: op1_01_in26 = reg_0777;
    70: op1_01_in26 = imem01_in[95:92];
    71: op1_01_in26 = reg_0260;
    74: op1_01_in26 = reg_0111;
    75: op1_01_in26 = reg_0387;
    76: op1_01_in26 = reg_0318;
    77: op1_01_in26 = imem06_in[39:36];
    80: op1_01_in26 = reg_0073;
    81: op1_01_in26 = reg_0759;
    82: op1_01_in26 = reg_0813;
    84: op1_01_in26 = reg_0449;
    85: op1_01_in26 = reg_0248;
    86: op1_01_in26 = reg_0239;
    87: op1_01_in26 = imem07_in[19:16];
    88: op1_01_in26 = reg_0601;
    89: op1_01_in26 = reg_0158;
    92: op1_01_in26 = imem04_in[91:88];
    93: op1_01_in26 = imem04_in[47:44];
    95: op1_01_in26 = imem04_in[47:44];
    94: op1_01_in26 = imem04_in[3:0];
    96: op1_01_in26 = reg_0256;
    default: op1_01_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv26 = 1;
    6: op1_01_inv26 = 1;
    9: op1_01_inv26 = 1;
    11: op1_01_inv26 = 1;
    12: op1_01_inv26 = 1;
    16: op1_01_inv26 = 1;
    17: op1_01_inv26 = 1;
    21: op1_01_inv26 = 1;
    23: op1_01_inv26 = 1;
    24: op1_01_inv26 = 1;
    28: op1_01_inv26 = 1;
    30: op1_01_inv26 = 1;
    31: op1_01_inv26 = 1;
    33: op1_01_inv26 = 1;
    34: op1_01_inv26 = 1;
    37: op1_01_inv26 = 1;
    39: op1_01_inv26 = 1;
    40: op1_01_inv26 = 1;
    42: op1_01_inv26 = 1;
    46: op1_01_inv26 = 1;
    51: op1_01_inv26 = 1;
    53: op1_01_inv26 = 1;
    54: op1_01_inv26 = 1;
    56: op1_01_inv26 = 1;
    57: op1_01_inv26 = 1;
    59: op1_01_inv26 = 1;
    60: op1_01_inv26 = 1;
    62: op1_01_inv26 = 1;
    63: op1_01_inv26 = 1;
    68: op1_01_inv26 = 1;
    71: op1_01_inv26 = 1;
    76: op1_01_inv26 = 1;
    80: op1_01_inv26 = 1;
    82: op1_01_inv26 = 1;
    84: op1_01_inv26 = 1;
    85: op1_01_inv26 = 1;
    86: op1_01_inv26 = 1;
    87: op1_01_inv26 = 1;
    88: op1_01_inv26 = 1;
    89: op1_01_inv26 = 1;
    92: op1_01_inv26 = 1;
    93: op1_01_inv26 = 1;
    default: op1_01_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in27 = reg_0329;
    6: op1_01_in27 = reg_0369;
    7: op1_01_in27 = imem07_in[59:56];
    8: op1_01_in27 = imem02_in[39:36];
    9: op1_01_in27 = reg_0387;
    10: op1_01_in27 = imem04_in[43:40];
    11: op1_01_in27 = reg_0514;
    12: op1_01_in27 = reg_0592;
    14: op1_01_in27 = reg_0359;
    15: op1_01_in27 = reg_0808;
    16: op1_01_in27 = reg_0356;
    17: op1_01_in27 = reg_0119;
    19: op1_01_in27 = imem01_in[95:92];
    20: op1_01_in27 = reg_0155;
    21: op1_01_in27 = reg_0511;
    22: op1_01_in27 = reg_0598;
    23: op1_01_in27 = reg_0443;
    24: op1_01_in27 = imem04_in[91:88];
    25: op1_01_in27 = reg_0630;
    26: op1_01_in27 = reg_0397;
    27: op1_01_in27 = reg_0407;
    28: op1_01_in27 = reg_0108;
    29: op1_01_in27 = reg_0093;
    30: op1_01_in27 = reg_0025;
    31: op1_01_in27 = reg_0515;
    32: op1_01_in27 = imem03_in[31:28];
    33: op1_01_in27 = reg_0809;
    34: op1_01_in27 = reg_0217;
    36: op1_01_in27 = reg_0215;
    37: op1_01_in27 = reg_0599;
    38: op1_01_in27 = reg_0532;
    39: op1_01_in27 = reg_0790;
    40: op1_01_in27 = reg_0542;
    42: op1_01_in27 = reg_0548;
    43: op1_01_in27 = imem03_in[51:48];
    44: op1_01_in27 = reg_0737;
    45: op1_01_in27 = reg_0157;
    46: op1_01_in27 = imem03_in[23:20];
    47: op1_01_in27 = imem04_in[115:112];
    50: op1_01_in27 = reg_0715;
    51: op1_01_in27 = imem05_in[87:84];
    52: op1_01_in27 = reg_0128;
    53: op1_01_in27 = imem06_in[111:108];
    54: op1_01_in27 = reg_0293;
    56: op1_01_in27 = reg_0733;
    57: op1_01_in27 = reg_0423;
    59: op1_01_in27 = reg_0399;
    60: op1_01_in27 = reg_0675;
    61: op1_01_in27 = reg_0063;
    62: op1_01_in27 = imem06_in[119:116];
    63: op1_01_in27 = reg_0447;
    68: op1_01_in27 = reg_0043;
    69: op1_01_in27 = reg_0620;
    70: op1_01_in27 = imem01_in[115:112];
    71: op1_01_in27 = reg_0242;
    74: op1_01_in27 = reg_0668;
    75: op1_01_in27 = reg_0557;
    76: op1_01_in27 = reg_0350;
    77: op1_01_in27 = imem06_in[79:76];
    80: op1_01_in27 = reg_0118;
    81: op1_01_in27 = reg_0241;
    82: op1_01_in27 = reg_0563;
    83: op1_01_in27 = reg_0292;
    84: op1_01_in27 = reg_0444;
    85: op1_01_in27 = reg_0506;
    86: op1_01_in27 = reg_0442;
    87: op1_01_in27 = imem07_in[31:28];
    88: op1_01_in27 = reg_0671;
    89: op1_01_in27 = reg_0064;
    92: op1_01_in27 = imem04_in[107:104];
    93: op1_01_in27 = imem04_in[123:120];
    94: op1_01_in27 = imem04_in[71:68];
    95: op1_01_in27 = imem04_in[55:52];
    96: op1_01_in27 = reg_0587;
    default: op1_01_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv27 = 1;
    6: op1_01_inv27 = 1;
    7: op1_01_inv27 = 1;
    10: op1_01_inv27 = 1;
    11: op1_01_inv27 = 1;
    12: op1_01_inv27 = 1;
    16: op1_01_inv27 = 1;
    17: op1_01_inv27 = 1;
    19: op1_01_inv27 = 1;
    21: op1_01_inv27 = 1;
    23: op1_01_inv27 = 1;
    27: op1_01_inv27 = 1;
    33: op1_01_inv27 = 1;
    39: op1_01_inv27 = 1;
    44: op1_01_inv27 = 1;
    47: op1_01_inv27 = 1;
    52: op1_01_inv27 = 1;
    53: op1_01_inv27 = 1;
    54: op1_01_inv27 = 1;
    56: op1_01_inv27 = 1;
    59: op1_01_inv27 = 1;
    60: op1_01_inv27 = 1;
    61: op1_01_inv27 = 1;
    68: op1_01_inv27 = 1;
    69: op1_01_inv27 = 1;
    70: op1_01_inv27 = 1;
    71: op1_01_inv27 = 1;
    77: op1_01_inv27 = 1;
    80: op1_01_inv27 = 1;
    83: op1_01_inv27 = 1;
    84: op1_01_inv27 = 1;
    85: op1_01_inv27 = 1;
    87: op1_01_inv27 = 1;
    88: op1_01_inv27 = 1;
    89: op1_01_inv27 = 1;
    94: op1_01_inv27 = 1;
    95: op1_01_inv27 = 1;
    default: op1_01_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in28 = reg_0330;
    6: op1_01_in28 = reg_0361;
    7: op1_01_in28 = imem07_in[75:72];
    8: op1_01_in28 = imem02_in[83:80];
    9: op1_01_in28 = reg_0370;
    10: op1_01_in28 = imem04_in[59:56];
    11: op1_01_in28 = reg_0227;
    12: op1_01_in28 = reg_0589;
    14: op1_01_in28 = reg_0318;
    15: op1_01_in28 = reg_0801;
    16: op1_01_in28 = reg_0406;
    17: op1_01_in28 = reg_0120;
    19: op1_01_in28 = imem01_in[99:96];
    20: op1_01_in28 = reg_0134;
    21: op1_01_in28 = reg_0237;
    22: op1_01_in28 = reg_0573;
    23: op1_01_in28 = reg_0437;
    24: op1_01_in28 = imem04_in[107:104];
    25: op1_01_in28 = reg_0633;
    26: op1_01_in28 = reg_0393;
    27: op1_01_in28 = reg_0405;
    30: op1_01_in28 = reg_0405;
    28: op1_01_in28 = reg_0100;
    29: op1_01_in28 = imem03_in[15:12];
    31: op1_01_in28 = reg_0761;
    32: op1_01_in28 = imem03_in[39:36];
    33: op1_01_in28 = imem04_in[39:36];
    34: op1_01_in28 = reg_0216;
    36: op1_01_in28 = reg_0506;
    37: op1_01_in28 = reg_0596;
    38: op1_01_in28 = imem03_in[31:28];
    39: op1_01_in28 = reg_0735;
    40: op1_01_in28 = reg_0056;
    42: op1_01_in28 = reg_0760;
    43: op1_01_in28 = imem03_in[55:52];
    46: op1_01_in28 = imem03_in[55:52];
    44: op1_01_in28 = reg_0148;
    45: op1_01_in28 = reg_0176;
    47: op1_01_in28 = reg_0315;
    50: op1_01_in28 = reg_0706;
    51: op1_01_in28 = imem05_in[91:88];
    52: op1_01_in28 = reg_0152;
    53: op1_01_in28 = imem06_in[127:124];
    54: op1_01_in28 = reg_0278;
    56: op1_01_in28 = reg_0668;
    57: op1_01_in28 = reg_0504;
    59: op1_01_in28 = reg_0751;
    60: op1_01_in28 = imem02_in[23:20];
    61: op1_01_in28 = reg_0582;
    62: op1_01_in28 = reg_0625;
    63: op1_01_in28 = reg_0061;
    68: op1_01_in28 = reg_0055;
    69: op1_01_in28 = reg_0218;
    70: op1_01_in28 = reg_0336;
    71: op1_01_in28 = reg_0369;
    74: op1_01_in28 = reg_0520;
    75: op1_01_in28 = reg_0570;
    76: op1_01_in28 = reg_0384;
    77: op1_01_in28 = imem06_in[91:88];
    80: op1_01_in28 = reg_0119;
    81: op1_01_in28 = reg_0244;
    82: op1_01_in28 = reg_0664;
    83: op1_01_in28 = reg_0431;
    84: op1_01_in28 = reg_0435;
    85: op1_01_in28 = reg_0123;
    86: op1_01_in28 = reg_0084;
    87: op1_01_in28 = reg_0725;
    88: op1_01_in28 = imem02_in[35:32];
    89: op1_01_in28 = reg_0253;
    92: op1_01_in28 = reg_0262;
    93: op1_01_in28 = reg_0247;
    94: op1_01_in28 = imem04_in[99:96];
    95: op1_01_in28 = imem04_in[63:60];
    96: op1_01_in28 = reg_0362;
    default: op1_01_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_01_inv28 = 1;
    6: op1_01_inv28 = 1;
    11: op1_01_inv28 = 1;
    12: op1_01_inv28 = 1;
    14: op1_01_inv28 = 1;
    16: op1_01_inv28 = 1;
    20: op1_01_inv28 = 1;
    21: op1_01_inv28 = 1;
    26: op1_01_inv28 = 1;
    28: op1_01_inv28 = 1;
    31: op1_01_inv28 = 1;
    32: op1_01_inv28 = 1;
    33: op1_01_inv28 = 1;
    34: op1_01_inv28 = 1;
    36: op1_01_inv28 = 1;
    38: op1_01_inv28 = 1;
    39: op1_01_inv28 = 1;
    40: op1_01_inv28 = 1;
    42: op1_01_inv28 = 1;
    46: op1_01_inv28 = 1;
    50: op1_01_inv28 = 1;
    54: op1_01_inv28 = 1;
    59: op1_01_inv28 = 1;
    62: op1_01_inv28 = 1;
    68: op1_01_inv28 = 1;
    69: op1_01_inv28 = 1;
    70: op1_01_inv28 = 1;
    71: op1_01_inv28 = 1;
    75: op1_01_inv28 = 1;
    77: op1_01_inv28 = 1;
    81: op1_01_inv28 = 1;
    82: op1_01_inv28 = 1;
    83: op1_01_inv28 = 1;
    84: op1_01_inv28 = 1;
    85: op1_01_inv28 = 1;
    86: op1_01_inv28 = 1;
    88: op1_01_inv28 = 1;
    89: op1_01_inv28 = 1;
    92: op1_01_inv28 = 1;
    93: op1_01_inv28 = 1;
    95: op1_01_inv28 = 1;
    default: op1_01_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in29 = reg_0342;
    6: op1_01_in29 = reg_0389;
    7: op1_01_in29 = reg_0728;
    8: op1_01_in29 = imem02_in[95:92];
    9: op1_01_in29 = reg_0343;
    10: op1_01_in29 = imem04_in[83:80];
    11: op1_01_in29 = reg_0518;
    12: op1_01_in29 = reg_0594;
    14: op1_01_in29 = reg_0310;
    15: op1_01_in29 = reg_0800;
    16: op1_01_in29 = reg_0367;
    17: op1_01_in29 = reg_0109;
    19: op1_01_in29 = reg_0233;
    20: op1_01_in29 = reg_0144;
    21: op1_01_in29 = reg_0504;
    22: op1_01_in29 = reg_0591;
    23: op1_01_in29 = reg_0162;
    24: op1_01_in29 = reg_0315;
    25: op1_01_in29 = reg_0618;
    26: op1_01_in29 = reg_0807;
    27: op1_01_in29 = reg_0403;
    30: op1_01_in29 = reg_0403;
    28: op1_01_in29 = imem02_in[3:0];
    29: op1_01_in29 = imem03_in[27:24];
    31: op1_01_in29 = reg_0241;
    32: op1_01_in29 = imem03_in[47:44];
    38: op1_01_in29 = imem03_in[47:44];
    33: op1_01_in29 = imem04_in[47:44];
    34: op1_01_in29 = reg_0247;
    36: op1_01_in29 = reg_0240;
    37: op1_01_in29 = reg_0592;
    39: op1_01_in29 = reg_0152;
    40: op1_01_in29 = reg_0057;
    42: op1_01_in29 = reg_0423;
    43: op1_01_in29 = imem03_in[107:104];
    44: op1_01_in29 = reg_0145;
    46: op1_01_in29 = imem03_in[83:80];
    47: op1_01_in29 = reg_0055;
    50: op1_01_in29 = reg_0727;
    51: op1_01_in29 = imem05_in[99:96];
    52: op1_01_in29 = reg_0143;
    53: op1_01_in29 = reg_0289;
    54: op1_01_in29 = reg_0370;
    56: op1_01_in29 = reg_0734;
    57: op1_01_in29 = reg_0419;
    59: op1_01_in29 = reg_0387;
    60: op1_01_in29 = imem02_in[71:68];
    61: op1_01_in29 = reg_0559;
    62: op1_01_in29 = reg_0291;
    63: op1_01_in29 = reg_0446;
    68: op1_01_in29 = reg_0058;
    69: op1_01_in29 = reg_0794;
    70: op1_01_in29 = reg_0085;
    71: op1_01_in29 = reg_0578;
    74: op1_01_in29 = reg_0102;
    75: op1_01_in29 = reg_0003;
    76: op1_01_in29 = reg_0564;
    77: op1_01_in29 = imem06_in[111:108];
    80: op1_01_in29 = reg_0601;
    81: op1_01_in29 = reg_0234;
    82: op1_01_in29 = reg_0652;
    83: op1_01_in29 = reg_0050;
    84: op1_01_in29 = reg_0110;
    85: op1_01_in29 = reg_0122;
    86: op1_01_in29 = reg_0267;
    87: op1_01_in29 = reg_0708;
    88: op1_01_in29 = imem02_in[115:112];
    89: op1_01_in29 = reg_0439;
    92: op1_01_in29 = reg_0177;
    93: op1_01_in29 = reg_0179;
    94: op1_01_in29 = imem04_in[119:116];
    95: op1_01_in29 = imem04_in[71:68];
    96: op1_01_in29 = reg_0320;
    default: op1_01_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_01_inv29 = 1;
    9: op1_01_inv29 = 1;
    12: op1_01_inv29 = 1;
    16: op1_01_inv29 = 1;
    17: op1_01_inv29 = 1;
    22: op1_01_inv29 = 1;
    25: op1_01_inv29 = 1;
    27: op1_01_inv29 = 1;
    30: op1_01_inv29 = 1;
    33: op1_01_inv29 = 1;
    34: op1_01_inv29 = 1;
    36: op1_01_inv29 = 1;
    37: op1_01_inv29 = 1;
    38: op1_01_inv29 = 1;
    40: op1_01_inv29 = 1;
    43: op1_01_inv29 = 1;
    50: op1_01_inv29 = 1;
    51: op1_01_inv29 = 1;
    52: op1_01_inv29 = 1;
    53: op1_01_inv29 = 1;
    54: op1_01_inv29 = 1;
    56: op1_01_inv29 = 1;
    57: op1_01_inv29 = 1;
    59: op1_01_inv29 = 1;
    60: op1_01_inv29 = 1;
    71: op1_01_inv29 = 1;
    74: op1_01_inv29 = 1;
    77: op1_01_inv29 = 1;
    83: op1_01_inv29 = 1;
    85: op1_01_inv29 = 1;
    86: op1_01_inv29 = 1;
    87: op1_01_inv29 = 1;
    89: op1_01_inv29 = 1;
    94: op1_01_inv29 = 1;
    96: op1_01_inv29 = 1;
    default: op1_01_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_01_in30 = reg_0083;
    6: op1_01_in30 = reg_0002;
    7: op1_01_in30 = reg_0719;
    8: op1_01_in30 = imem02_in[111:108];
    9: op1_01_in30 = reg_0385;
    10: op1_01_in30 = imem04_in[91:88];
    33: op1_01_in30 = imem04_in[91:88];
    95: op1_01_in30 = imem04_in[91:88];
    11: op1_01_in30 = reg_0515;
    12: op1_01_in30 = reg_0581;
    96: op1_01_in30 = reg_0581;
    14: op1_01_in30 = reg_0092;
    15: op1_01_in30 = reg_0805;
    75: op1_01_in30 = reg_0805;
    16: op1_01_in30 = reg_0747;
    17: op1_01_in30 = reg_0107;
    19: op1_01_in30 = reg_0119;
    85: op1_01_in30 = reg_0119;
    20: op1_01_in30 = imem06_in[123:120];
    21: op1_01_in30 = reg_0124;
    22: op1_01_in30 = reg_0563;
    23: op1_01_in30 = reg_0158;
    24: op1_01_in30 = reg_0553;
    25: op1_01_in30 = reg_0623;
    26: op1_01_in30 = reg_0804;
    27: op1_01_in30 = reg_0406;
    28: op1_01_in30 = imem02_in[43:40];
    29: op1_01_in30 = imem03_in[47:44];
    30: op1_01_in30 = reg_0038;
    31: op1_01_in30 = reg_0215;
    32: op1_01_in30 = imem03_in[51:48];
    34: op1_01_in30 = reg_0249;
    36: op1_01_in30 = reg_0219;
    57: op1_01_in30 = reg_0219;
    37: op1_01_in30 = reg_0591;
    38: op1_01_in30 = imem03_in[59:56];
    39: op1_01_in30 = reg_0129;
    40: op1_01_in30 = reg_0052;
    42: op1_01_in30 = reg_0424;
    81: op1_01_in30 = reg_0424;
    43: op1_01_in30 = reg_0589;
    44: op1_01_in30 = reg_0142;
    46: op1_01_in30 = imem03_in[99:96];
    47: op1_01_in30 = reg_0057;
    50: op1_01_in30 = reg_0051;
    51: op1_01_in30 = imem05_in[107:104];
    52: op1_01_in30 = reg_0153;
    53: op1_01_in30 = reg_0020;
    54: op1_01_in30 = reg_0409;
    56: op1_01_in30 = reg_0557;
    59: op1_01_in30 = reg_0569;
    60: op1_01_in30 = imem02_in[95:92];
    61: op1_01_in30 = reg_0493;
    62: op1_01_in30 = reg_0349;
    63: op1_01_in30 = reg_0440;
    68: op1_01_in30 = reg_0500;
    69: op1_01_in30 = reg_0787;
    82: op1_01_in30 = reg_0787;
    70: op1_01_in30 = reg_0388;
    71: op1_01_in30 = reg_0775;
    74: op1_01_in30 = reg_0394;
    76: op1_01_in30 = reg_0372;
    77: op1_01_in30 = reg_0625;
    80: op1_01_in30 = imem02_in[51:48];
    83: op1_01_in30 = reg_0585;
    84: op1_01_in30 = reg_0170;
    86: op1_01_in30 = reg_0438;
    87: op1_01_in30 = reg_0157;
    88: op1_01_in30 = reg_0031;
    89: op1_01_in30 = reg_0449;
    92: op1_01_in30 = reg_0537;
    93: op1_01_in30 = reg_0535;
    94: op1_01_in30 = imem04_in[123:120];
    default: op1_01_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_01_inv30 = 1;
    8: op1_01_inv30 = 1;
    9: op1_01_inv30 = 1;
    12: op1_01_inv30 = 1;
    14: op1_01_inv30 = 1;
    15: op1_01_inv30 = 1;
    19: op1_01_inv30 = 1;
    23: op1_01_inv30 = 1;
    25: op1_01_inv30 = 1;
    27: op1_01_inv30 = 1;
    28: op1_01_inv30 = 1;
    29: op1_01_inv30 = 1;
    32: op1_01_inv30 = 1;
    37: op1_01_inv30 = 1;
    42: op1_01_inv30 = 1;
    44: op1_01_inv30 = 1;
    50: op1_01_inv30 = 1;
    52: op1_01_inv30 = 1;
    56: op1_01_inv30 = 1;
    57: op1_01_inv30 = 1;
    60: op1_01_inv30 = 1;
    61: op1_01_inv30 = 1;
    63: op1_01_inv30 = 1;
    68: op1_01_inv30 = 1;
    69: op1_01_inv30 = 1;
    76: op1_01_inv30 = 1;
    80: op1_01_inv30 = 1;
    85: op1_01_inv30 = 1;
    89: op1_01_inv30 = 1;
    96: op1_01_inv30 = 1;
    default: op1_01_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_01_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in00 = reg_0042;
    5: op1_02_in00 = imem00_in[43:40];
    6: op1_02_in00 = reg_0807;
    7: op1_02_in00 = imem00_in[27:24];
    67: op1_02_in00 = imem00_in[27:24];
    8: op1_02_in00 = imem02_in[115:112];
    3: op1_02_in00 = imem07_in[75:72];
    9: op1_02_in00 = reg_0322;
    2: op1_02_in00 = imem07_in[43:40];
    10: op1_02_in00 = imem04_in[107:104];
    11: op1_02_in00 = reg_0776;
    12: op1_02_in00 = reg_0387;
    13: op1_02_in00 = imem00_in[15:12];
    72: op1_02_in00 = imem00_in[15:12];
    90: op1_02_in00 = imem00_in[15:12];
    14: op1_02_in00 = reg_0089;
    1: op1_02_in00 = imem07_in[23:20];
    15: op1_02_in00 = reg_0802;
    16: op1_02_in00 = reg_0035;
    17: op1_02_in00 = imem02_in[27:24];
    18: op1_02_in00 = imem00_in[3:0];
    55: op1_02_in00 = imem00_in[3:0];
    73: op1_02_in00 = imem00_in[3:0];
    89: op1_02_in00 = imem00_in[3:0];
    91: op1_02_in00 = imem00_in[3:0];
    19: op1_02_in00 = reg_0115;
    20: op1_02_in00 = reg_0628;
    21: op1_02_in00 = reg_0108;
    22: op1_02_in00 = reg_0585;
    23: op1_02_in00 = imem00_in[111:108];
    24: op1_02_in00 = reg_0060;
    25: op1_02_in00 = reg_0615;
    26: op1_02_in00 = imem04_in[15:12];
    27: op1_02_in00 = reg_0039;
    28: op1_02_in00 = reg_0661;
    82: op1_02_in00 = reg_0661;
    29: op1_02_in00 = imem03_in[119:116];
    30: op1_02_in00 = reg_0031;
    31: op1_02_in00 = reg_0502;
    32: op1_02_in00 = imem03_in[55:52];
    33: op1_02_in00 = imem04_in[115:112];
    34: op1_02_in00 = reg_0124;
    35: op1_02_in00 = imem00_in[87:84];
    36: op1_02_in00 = reg_0118;
    37: op1_02_in00 = reg_0581;
    38: op1_02_in00 = imem03_in[115:112];
    46: op1_02_in00 = imem03_in[115:112];
    39: op1_02_in00 = reg_0130;
    40: op1_02_in00 = reg_0297;
    41: op1_02_in00 = imem00_in[59:56];
    42: op1_02_in00 = reg_0219;
    43: op1_02_in00 = reg_0580;
    44: op1_02_in00 = reg_0146;
    45: op1_02_in00 = imem00_in[39:36];
    48: op1_02_in00 = imem00_in[39:36];
    47: op1_02_in00 = reg_0516;
    49: op1_02_in00 = imem00_in[7:4];
    65: op1_02_in00 = imem00_in[7:4];
    79: op1_02_in00 = imem00_in[7:4];
    50: op1_02_in00 = reg_0434;
    51: op1_02_in00 = reg_0791;
    52: op1_02_in00 = imem06_in[11:8];
    53: op1_02_in00 = reg_0371;
    54: op1_02_in00 = reg_0576;
    71: op1_02_in00 = reg_0576;
    56: op1_02_in00 = reg_0574;
    57: op1_02_in00 = reg_0105;
    58: op1_02_in00 = imem00_in[35:32];
    78: op1_02_in00 = imem00_in[35:32];
    59: op1_02_in00 = reg_0562;
    60: op1_02_in00 = imem02_in[99:96];
    61: op1_02_in00 = reg_0591;
    62: op1_02_in00 = reg_0619;
    63: op1_02_in00 = reg_0084;
    64: op1_02_in00 = imem00_in[19:16];
    66: op1_02_in00 = imem00_in[75:72];
    68: op1_02_in00 = reg_0283;
    69: op1_02_in00 = reg_0029;
    70: op1_02_in00 = reg_0737;
    74: op1_02_in00 = reg_0294;
    75: op1_02_in00 = reg_0806;
    76: op1_02_in00 = reg_0549;
    77: op1_02_in00 = reg_0346;
    80: op1_02_in00 = imem02_in[59:56];
    81: op1_02_in00 = reg_0420;
    83: op1_02_in00 = reg_0311;
    84: op1_02_in00 = imem00_in[31:28];
    85: op1_02_in00 = reg_0672;
    86: op1_02_in00 = reg_0116;
    87: op1_02_in00 = reg_0731;
    88: op1_02_in00 = reg_0639;
    92: op1_02_in00 = reg_0554;
    93: op1_02_in00 = reg_0554;
    94: op1_02_in00 = reg_0173;
    95: op1_02_in00 = imem04_in[123:120];
    96: op1_02_in00 = reg_0594;
    default: op1_02_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv00 = 1;
    5: op1_02_inv00 = 1;
    6: op1_02_inv00 = 1;
    8: op1_02_inv00 = 1;
    11: op1_02_inv00 = 1;
    13: op1_02_inv00 = 1;
    14: op1_02_inv00 = 1;
    15: op1_02_inv00 = 1;
    19: op1_02_inv00 = 1;
    20: op1_02_inv00 = 1;
    21: op1_02_inv00 = 1;
    22: op1_02_inv00 = 1;
    23: op1_02_inv00 = 1;
    24: op1_02_inv00 = 1;
    25: op1_02_inv00 = 1;
    27: op1_02_inv00 = 1;
    29: op1_02_inv00 = 1;
    32: op1_02_inv00 = 1;
    33: op1_02_inv00 = 1;
    36: op1_02_inv00 = 1;
    37: op1_02_inv00 = 1;
    39: op1_02_inv00 = 1;
    40: op1_02_inv00 = 1;
    43: op1_02_inv00 = 1;
    45: op1_02_inv00 = 1;
    49: op1_02_inv00 = 1;
    52: op1_02_inv00 = 1;
    53: op1_02_inv00 = 1;
    54: op1_02_inv00 = 1;
    56: op1_02_inv00 = 1;
    58: op1_02_inv00 = 1;
    59: op1_02_inv00 = 1;
    62: op1_02_inv00 = 1;
    63: op1_02_inv00 = 1;
    66: op1_02_inv00 = 1;
    68: op1_02_inv00 = 1;
    69: op1_02_inv00 = 1;
    70: op1_02_inv00 = 1;
    73: op1_02_inv00 = 1;
    76: op1_02_inv00 = 1;
    77: op1_02_inv00 = 1;
    78: op1_02_inv00 = 1;
    80: op1_02_inv00 = 1;
    81: op1_02_inv00 = 1;
    85: op1_02_inv00 = 1;
    86: op1_02_inv00 = 1;
    87: op1_02_inv00 = 1;
    89: op1_02_inv00 = 1;
    91: op1_02_inv00 = 1;
    93: op1_02_inv00 = 1;
    95: op1_02_inv00 = 1;
    96: op1_02_inv00 = 1;
    default: op1_02_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in01 = reg_0080;
    14: op1_02_in01 = reg_0080;
    5: op1_02_in01 = imem00_in[127:124];
    6: op1_02_in01 = reg_0801;
    7: op1_02_in01 = imem00_in[51:48];
    13: op1_02_in01 = imem00_in[51:48];
    48: op1_02_in01 = imem00_in[51:48];
    8: op1_02_in01 = imem02_in[119:116];
    3: op1_02_in01 = reg_0425;
    9: op1_02_in01 = reg_0398;
    2: op1_02_in01 = imem07_in[71:68];
    10: op1_02_in01 = imem04_in[119:116];
    11: op1_02_in01 = reg_0755;
    12: op1_02_in01 = reg_0391;
    1: op1_02_in01 = imem07_in[27:24];
    15: op1_02_in01 = imem04_in[7:4];
    16: op1_02_in01 = reg_0750;
    17: op1_02_in01 = imem02_in[87:84];
    80: op1_02_in01 = imem02_in[87:84];
    18: op1_02_in01 = imem00_in[23:20];
    49: op1_02_in01 = imem00_in[23:20];
    19: op1_02_in01 = reg_0127;
    20: op1_02_in01 = reg_0610;
    21: op1_02_in01 = reg_0126;
    85: op1_02_in01 = reg_0126;
    22: op1_02_in01 = reg_0597;
    23: op1_02_in01 = imem00_in[119:116];
    24: op1_02_in01 = reg_0554;
    25: op1_02_in01 = reg_0381;
    26: op1_02_in01 = imem04_in[19:16];
    27: op1_02_in01 = reg_0753;
    28: op1_02_in01 = reg_0639;
    29: op1_02_in01 = imem03_in[123:120];
    38: op1_02_in01 = imem03_in[123:120];
    30: op1_02_in01 = reg_0818;
    31: op1_02_in01 = reg_0216;
    32: op1_02_in01 = imem03_in[59:56];
    33: op1_02_in01 = reg_0553;
    34: op1_02_in01 = reg_0107;
    35: op1_02_in01 = imem00_in[99:96];
    36: op1_02_in01 = reg_0112;
    37: op1_02_in01 = reg_0588;
    43: op1_02_in01 = reg_0588;
    39: op1_02_in01 = reg_0140;
    40: op1_02_in01 = reg_0079;
    41: op1_02_in01 = imem00_in[79:76];
    42: op1_02_in01 = reg_0099;
    44: op1_02_in01 = reg_0154;
    45: op1_02_in01 = imem00_in[63:60];
    58: op1_02_in01 = imem00_in[63:60];
    46: op1_02_in01 = reg_0598;
    47: op1_02_in01 = reg_0303;
    50: op1_02_in01 = reg_0443;
    51: op1_02_in01 = reg_0796;
    52: op1_02_in01 = imem06_in[47:44];
    53: op1_02_in01 = reg_0606;
    54: op1_02_in01 = reg_0620;
    55: op1_02_in01 = imem00_in[47:44];
    78: op1_02_in01 = imem00_in[47:44];
    89: op1_02_in01 = imem00_in[47:44];
    90: op1_02_in01 = imem00_in[47:44];
    56: op1_02_in01 = reg_0054;
    57: op1_02_in01 = reg_0124;
    74: op1_02_in01 = reg_0124;
    59: op1_02_in01 = reg_0572;
    60: op1_02_in01 = reg_0664;
    61: op1_02_in01 = reg_0329;
    62: op1_02_in01 = reg_0618;
    63: op1_02_in01 = reg_0438;
    64: op1_02_in01 = imem00_in[31:28];
    73: op1_02_in01 = imem00_in[31:28];
    65: op1_02_in01 = imem00_in[27:24];
    79: op1_02_in01 = imem00_in[27:24];
    66: op1_02_in01 = imem00_in[87:84];
    72: op1_02_in01 = imem00_in[87:84];
    67: op1_02_in01 = imem00_in[67:64];
    68: op1_02_in01 = reg_0611;
    69: op1_02_in01 = reg_0752;
    82: op1_02_in01 = reg_0752;
    70: op1_02_in01 = reg_0511;
    71: op1_02_in01 = reg_0512;
    75: op1_02_in01 = reg_0810;
    76: op1_02_in01 = reg_0012;
    77: op1_02_in01 = reg_0291;
    81: op1_02_in01 = reg_0104;
    83: op1_02_in01 = reg_0233;
    84: op1_02_in01 = imem00_in[59:56];
    86: op1_02_in01 = reg_0181;
    87: op1_02_in01 = reg_0727;
    88: op1_02_in01 = reg_0647;
    91: op1_02_in01 = imem00_in[35:32];
    92: op1_02_in01 = reg_0523;
    93: op1_02_in01 = reg_0261;
    94: op1_02_in01 = reg_0275;
    95: op1_02_in01 = reg_0060;
    96: op1_02_in01 = reg_0281;
    default: op1_02_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_02_inv01 = 1;
    8: op1_02_inv01 = 1;
    3: op1_02_inv01 = 1;
    2: op1_02_inv01 = 1;
    10: op1_02_inv01 = 1;
    12: op1_02_inv01 = 1;
    18: op1_02_inv01 = 1;
    19: op1_02_inv01 = 1;
    26: op1_02_inv01 = 1;
    30: op1_02_inv01 = 1;
    31: op1_02_inv01 = 1;
    32: op1_02_inv01 = 1;
    34: op1_02_inv01 = 1;
    35: op1_02_inv01 = 1;
    37: op1_02_inv01 = 1;
    38: op1_02_inv01 = 1;
    41: op1_02_inv01 = 1;
    42: op1_02_inv01 = 1;
    43: op1_02_inv01 = 1;
    44: op1_02_inv01 = 1;
    45: op1_02_inv01 = 1;
    48: op1_02_inv01 = 1;
    49: op1_02_inv01 = 1;
    53: op1_02_inv01 = 1;
    55: op1_02_inv01 = 1;
    56: op1_02_inv01 = 1;
    58: op1_02_inv01 = 1;
    60: op1_02_inv01 = 1;
    62: op1_02_inv01 = 1;
    63: op1_02_inv01 = 1;
    65: op1_02_inv01 = 1;
    67: op1_02_inv01 = 1;
    68: op1_02_inv01 = 1;
    70: op1_02_inv01 = 1;
    71: op1_02_inv01 = 1;
    72: op1_02_inv01 = 1;
    73: op1_02_inv01 = 1;
    75: op1_02_inv01 = 1;
    79: op1_02_inv01 = 1;
    80: op1_02_inv01 = 1;
    81: op1_02_inv01 = 1;
    83: op1_02_inv01 = 1;
    88: op1_02_inv01 = 1;
    89: op1_02_inv01 = 1;
    92: op1_02_inv01 = 1;
    94: op1_02_inv01 = 1;
    default: op1_02_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in02 = imem03_in[7:4];
    5: op1_02_in02 = reg_0675;
    6: op1_02_in02 = reg_0800;
    7: op1_02_in02 = imem00_in[71:68];
    45: op1_02_in02 = imem00_in[71:68];
    64: op1_02_in02 = imem00_in[71:68];
    8: op1_02_in02 = reg_0649;
    3: op1_02_in02 = reg_0430;
    9: op1_02_in02 = reg_0312;
    2: op1_02_in02 = imem07_in[115:112];
    10: op1_02_in02 = imem04_in[127:124];
    11: op1_02_in02 = reg_0218;
    12: op1_02_in02 = reg_0370;
    13: op1_02_in02 = imem00_in[91:88];
    67: op1_02_in02 = imem00_in[91:88];
    14: op1_02_in02 = reg_0095;
    1: op1_02_in02 = imem07_in[87:84];
    15: op1_02_in02 = imem04_in[11:8];
    16: op1_02_in02 = reg_0030;
    30: op1_02_in02 = reg_0030;
    17: op1_02_in02 = imem02_in[99:96];
    18: op1_02_in02 = imem00_in[35:32];
    19: op1_02_in02 = imem02_in[43:40];
    34: op1_02_in02 = imem02_in[43:40];
    20: op1_02_in02 = reg_0629;
    21: op1_02_in02 = imem02_in[7:4];
    22: op1_02_in02 = reg_0581;
    23: op1_02_in02 = reg_0698;
    24: op1_02_in02 = reg_0558;
    25: op1_02_in02 = reg_0372;
    26: op1_02_in02 = imem04_in[51:48];
    27: op1_02_in02 = reg_0812;
    28: op1_02_in02 = reg_0647;
    29: op1_02_in02 = reg_0602;
    32: op1_02_in02 = reg_0602;
    38: op1_02_in02 = reg_0602;
    31: op1_02_in02 = reg_0236;
    86: op1_02_in02 = reg_0236;
    33: op1_02_in02 = reg_0542;
    35: op1_02_in02 = imem00_in[103:100];
    41: op1_02_in02 = imem00_in[103:100];
    36: op1_02_in02 = reg_0106;
    37: op1_02_in02 = reg_0751;
    43: op1_02_in02 = reg_0751;
    39: op1_02_in02 = reg_0144;
    40: op1_02_in02 = reg_0076;
    42: op1_02_in02 = reg_0120;
    81: op1_02_in02 = reg_0120;
    44: op1_02_in02 = reg_0140;
    46: op1_02_in02 = reg_0583;
    47: op1_02_in02 = reg_0280;
    48: op1_02_in02 = imem00_in[75:72];
    90: op1_02_in02 = imem00_in[75:72];
    49: op1_02_in02 = imem00_in[31:28];
    50: op1_02_in02 = reg_0437;
    51: op1_02_in02 = reg_0488;
    52: op1_02_in02 = imem06_in[67:64];
    53: op1_02_in02 = reg_0619;
    54: op1_02_in02 = reg_0040;
    55: op1_02_in02 = imem00_in[55:52];
    91: op1_02_in02 = imem00_in[55:52];
    56: op1_02_in02 = reg_0567;
    57: op1_02_in02 = reg_0073;
    58: op1_02_in02 = imem00_in[95:92];
    72: op1_02_in02 = imem00_in[95:92];
    59: op1_02_in02 = reg_0397;
    60: op1_02_in02 = reg_0417;
    61: op1_02_in02 = reg_0399;
    62: op1_02_in02 = reg_0401;
    63: op1_02_in02 = reg_0169;
    65: op1_02_in02 = imem00_in[39:36];
    66: op1_02_in02 = imem00_in[107:104];
    68: op1_02_in02 = reg_0077;
    69: op1_02_in02 = reg_0367;
    70: op1_02_in02 = reg_0422;
    71: op1_02_in02 = reg_0777;
    73: op1_02_in02 = imem00_in[59:56];
    78: op1_02_in02 = imem00_in[59:56];
    74: op1_02_in02 = reg_0670;
    75: op1_02_in02 = imem04_in[31:28];
    76: op1_02_in02 = reg_0007;
    77: op1_02_in02 = reg_0815;
    79: op1_02_in02 = imem00_in[63:60];
    80: op1_02_in02 = imem02_in[103:100];
    82: op1_02_in02 = reg_0011;
    83: op1_02_in02 = imem05_in[7:4];
    84: op1_02_in02 = imem00_in[83:80];
    85: op1_02_in02 = imem02_in[31:28];
    87: op1_02_in02 = reg_0295;
    88: op1_02_in02 = reg_0498;
    89: op1_02_in02 = imem00_in[115:112];
    92: op1_02_in02 = reg_0432;
    93: op1_02_in02 = reg_0536;
    94: op1_02_in02 = reg_0058;
    95: op1_02_in02 = reg_0174;
    96: op1_02_in02 = reg_0097;
    default: op1_02_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv02 = 1;
    5: op1_02_inv02 = 1;
    6: op1_02_inv02 = 1;
    7: op1_02_inv02 = 1;
    9: op1_02_inv02 = 1;
    2: op1_02_inv02 = 1;
    10: op1_02_inv02 = 1;
    13: op1_02_inv02 = 1;
    14: op1_02_inv02 = 1;
    1: op1_02_inv02 = 1;
    15: op1_02_inv02 = 1;
    17: op1_02_inv02 = 1;
    20: op1_02_inv02 = 1;
    26: op1_02_inv02 = 1;
    27: op1_02_inv02 = 1;
    28: op1_02_inv02 = 1;
    30: op1_02_inv02 = 1;
    31: op1_02_inv02 = 1;
    32: op1_02_inv02 = 1;
    33: op1_02_inv02 = 1;
    35: op1_02_inv02 = 1;
    36: op1_02_inv02 = 1;
    37: op1_02_inv02 = 1;
    39: op1_02_inv02 = 1;
    41: op1_02_inv02 = 1;
    42: op1_02_inv02 = 1;
    46: op1_02_inv02 = 1;
    49: op1_02_inv02 = 1;
    51: op1_02_inv02 = 1;
    52: op1_02_inv02 = 1;
    54: op1_02_inv02 = 1;
    55: op1_02_inv02 = 1;
    57: op1_02_inv02 = 1;
    58: op1_02_inv02 = 1;
    61: op1_02_inv02 = 1;
    62: op1_02_inv02 = 1;
    67: op1_02_inv02 = 1;
    71: op1_02_inv02 = 1;
    72: op1_02_inv02 = 1;
    73: op1_02_inv02 = 1;
    75: op1_02_inv02 = 1;
    76: op1_02_inv02 = 1;
    77: op1_02_inv02 = 1;
    78: op1_02_inv02 = 1;
    79: op1_02_inv02 = 1;
    80: op1_02_inv02 = 1;
    82: op1_02_inv02 = 1;
    88: op1_02_inv02 = 1;
    89: op1_02_inv02 = 1;
    90: op1_02_inv02 = 1;
    91: op1_02_inv02 = 1;
    93: op1_02_inv02 = 1;
    94: op1_02_inv02 = 1;
    96: op1_02_inv02 = 1;
    default: op1_02_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in03 = imem03_in[39:36];
    5: op1_02_in03 = reg_0680;
    6: op1_02_in03 = reg_0004;
    7: op1_02_in03 = imem00_in[79:76];
    79: op1_02_in03 = imem00_in[79:76];
    8: op1_02_in03 = reg_0320;
    3: op1_02_in03 = reg_0431;
    9: op1_02_in03 = reg_0361;
    2: op1_02_in03 = imem07_in[119:116];
    10: op1_02_in03 = reg_0545;
    11: op1_02_in03 = reg_0242;
    12: op1_02_in03 = reg_0388;
    13: op1_02_in03 = imem00_in[111:108];
    41: op1_02_in03 = imem00_in[111:108];
    84: op1_02_in03 = imem00_in[111:108];
    14: op1_02_in03 = reg_0090;
    1: op1_02_in03 = imem07_in[91:88];
    15: op1_02_in03 = imem04_in[51:48];
    16: op1_02_in03 = imem07_in[71:68];
    17: op1_02_in03 = imem02_in[103:100];
    18: op1_02_in03 = imem00_in[39:36];
    19: op1_02_in03 = imem02_in[47:44];
    20: op1_02_in03 = reg_0607;
    21: op1_02_in03 = imem02_in[67:64];
    22: op1_02_in03 = reg_0391;
    23: op1_02_in03 = reg_0688;
    24: op1_02_in03 = reg_0516;
    93: op1_02_in03 = reg_0516;
    25: op1_02_in03 = reg_0408;
    26: op1_02_in03 = imem04_in[127:124];
    27: op1_02_in03 = reg_0813;
    28: op1_02_in03 = reg_0636;
    29: op1_02_in03 = reg_0586;
    30: op1_02_in03 = imem07_in[47:44];
    31: op1_02_in03 = reg_0248;
    32: op1_02_in03 = reg_0601;
    33: op1_02_in03 = reg_0500;
    34: op1_02_in03 = imem02_in[55:52];
    35: op1_02_in03 = reg_0681;
    36: op1_02_in03 = reg_0110;
    37: op1_02_in03 = reg_0394;
    38: op1_02_in03 = reg_0039;
    39: op1_02_in03 = imem06_in[63:60];
    40: op1_02_in03 = reg_0071;
    47: op1_02_in03 = reg_0071;
    42: op1_02_in03 = imem02_in[7:4];
    43: op1_02_in03 = reg_0387;
    44: op1_02_in03 = imem06_in[43:40];
    45: op1_02_in03 = imem00_in[83:80];
    64: op1_02_in03 = imem00_in[83:80];
    46: op1_02_in03 = reg_0589;
    48: op1_02_in03 = imem00_in[87:84];
    49: op1_02_in03 = imem00_in[35:32];
    50: op1_02_in03 = reg_0174;
    51: op1_02_in03 = reg_0795;
    52: op1_02_in03 = imem06_in[95:92];
    53: op1_02_in03 = reg_0622;
    54: op1_02_in03 = reg_0814;
    55: op1_02_in03 = imem00_in[91:88];
    56: op1_02_in03 = reg_0216;
    57: op1_02_in03 = reg_0121;
    58: op1_02_in03 = imem00_in[107:104];
    59: op1_02_in03 = reg_0374;
    60: op1_02_in03 = reg_0665;
    61: op1_02_in03 = reg_0281;
    62: op1_02_in03 = reg_0519;
    63: op1_02_in03 = reg_0182;
    65: op1_02_in03 = imem00_in[47:44];
    66: op1_02_in03 = imem00_in[127:124];
    67: op1_02_in03 = imem00_in[103:100];
    68: op1_02_in03 = reg_0627;
    69: op1_02_in03 = imem07_in[7:4];
    70: op1_02_in03 = reg_0054;
    71: op1_02_in03 = reg_0484;
    72: op1_02_in03 = imem00_in[99:96];
    73: op1_02_in03 = imem00_in[75:72];
    74: op1_02_in03 = reg_0669;
    75: op1_02_in03 = reg_0553;
    76: op1_02_in03 = reg_0807;
    77: op1_02_in03 = reg_0605;
    78: op1_02_in03 = imem00_in[63:60];
    80: op1_02_in03 = reg_0254;
    81: op1_02_in03 = reg_0126;
    82: op1_02_in03 = reg_0367;
    83: op1_02_in03 = imem05_in[71:68];
    85: op1_02_in03 = imem02_in[63:60];
    86: op1_02_in03 = reg_0142;
    87: op1_02_in03 = reg_0053;
    88: op1_02_in03 = reg_0087;
    89: op1_02_in03 = reg_0693;
    90: op1_02_in03 = imem00_in[95:92];
    91: op1_02_in03 = imem00_in[59:56];
    92: op1_02_in03 = reg_0433;
    94: op1_02_in03 = reg_0523;
    95: op1_02_in03 = reg_0611;
    96: op1_02_in03 = reg_0487;
    default: op1_02_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_02_inv03 = 1;
    8: op1_02_inv03 = 1;
    9: op1_02_inv03 = 1;
    10: op1_02_inv03 = 1;
    11: op1_02_inv03 = 1;
    12: op1_02_inv03 = 1;
    14: op1_02_inv03 = 1;
    16: op1_02_inv03 = 1;
    18: op1_02_inv03 = 1;
    19: op1_02_inv03 = 1;
    20: op1_02_inv03 = 1;
    21: op1_02_inv03 = 1;
    25: op1_02_inv03 = 1;
    26: op1_02_inv03 = 1;
    27: op1_02_inv03 = 1;
    29: op1_02_inv03 = 1;
    31: op1_02_inv03 = 1;
    35: op1_02_inv03 = 1;
    36: op1_02_inv03 = 1;
    37: op1_02_inv03 = 1;
    39: op1_02_inv03 = 1;
    42: op1_02_inv03 = 1;
    43: op1_02_inv03 = 1;
    47: op1_02_inv03 = 1;
    50: op1_02_inv03 = 1;
    54: op1_02_inv03 = 1;
    58: op1_02_inv03 = 1;
    59: op1_02_inv03 = 1;
    60: op1_02_inv03 = 1;
    62: op1_02_inv03 = 1;
    63: op1_02_inv03 = 1;
    64: op1_02_inv03 = 1;
    65: op1_02_inv03 = 1;
    67: op1_02_inv03 = 1;
    74: op1_02_inv03 = 1;
    75: op1_02_inv03 = 1;
    78: op1_02_inv03 = 1;
    81: op1_02_inv03 = 1;
    83: op1_02_inv03 = 1;
    86: op1_02_inv03 = 1;
    87: op1_02_inv03 = 1;
    90: op1_02_inv03 = 1;
    91: op1_02_inv03 = 1;
    92: op1_02_inv03 = 1;
    95: op1_02_inv03 = 1;
    default: op1_02_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in04 = imem03_in[43:40];
    5: op1_02_in04 = reg_0692;
    6: op1_02_in04 = imem04_in[123:120];
    7: op1_02_in04 = imem00_in[83:80];
    91: op1_02_in04 = imem00_in[83:80];
    8: op1_02_in04 = reg_0318;
    3: op1_02_in04 = reg_0184;
    9: op1_02_in04 = reg_0396;
    2: op1_02_in04 = reg_0175;
    50: op1_02_in04 = reg_0175;
    10: op1_02_in04 = reg_0550;
    11: op1_02_in04 = reg_0216;
    12: op1_02_in04 = reg_0362;
    13: op1_02_in04 = reg_0695;
    66: op1_02_in04 = reg_0695;
    14: op1_02_in04 = reg_0087;
    1: op1_02_in04 = imem07_in[103:100];
    15: op1_02_in04 = imem04_in[67:64];
    16: op1_02_in04 = imem07_in[115:112];
    17: op1_02_in04 = imem02_in[119:116];
    18: op1_02_in04 = imem00_in[43:40];
    19: op1_02_in04 = reg_0658;
    20: op1_02_in04 = reg_0605;
    21: op1_02_in04 = imem02_in[83:80];
    22: op1_02_in04 = reg_0321;
    23: op1_02_in04 = reg_0463;
    24: op1_02_in04 = reg_0308;
    25: op1_02_in04 = reg_0405;
    26: op1_02_in04 = reg_0328;
    27: op1_02_in04 = reg_0748;
    28: op1_02_in04 = reg_0663;
    29: op1_02_in04 = reg_0599;
    30: op1_02_in04 = imem07_in[67:64];
    31: op1_02_in04 = reg_0041;
    32: op1_02_in04 = reg_0592;
    33: op1_02_in04 = reg_0556;
    34: op1_02_in04 = imem02_in[59:56];
    35: op1_02_in04 = reg_0676;
    36: op1_02_in04 = imem02_in[11:8];
    37: op1_02_in04 = reg_0564;
    38: op1_02_in04 = reg_0387;
    39: op1_02_in04 = imem06_in[71:68];
    40: op1_02_in04 = reg_0070;
    41: op1_02_in04 = reg_0682;
    42: op1_02_in04 = imem02_in[23:20];
    43: op1_02_in04 = reg_0562;
    44: op1_02_in04 = imem06_in[47:44];
    45: op1_02_in04 = imem00_in[99:96];
    46: op1_02_in04 = reg_0580;
    47: op1_02_in04 = reg_0616;
    95: op1_02_in04 = reg_0616;
    48: op1_02_in04 = imem00_in[95:92];
    73: op1_02_in04 = imem00_in[95:92];
    49: op1_02_in04 = imem00_in[51:48];
    51: op1_02_in04 = reg_0784;
    52: op1_02_in04 = imem06_in[123:120];
    53: op1_02_in04 = reg_0612;
    54: op1_02_in04 = reg_0375;
    55: op1_02_in04 = reg_0697;
    56: op1_02_in04 = reg_0290;
    57: op1_02_in04 = imem02_in[43:40];
    58: op1_02_in04 = imem00_in[119:116];
    59: op1_02_in04 = reg_0001;
    60: op1_02_in04 = reg_0426;
    61: op1_02_in04 = reg_0588;
    62: op1_02_in04 = reg_0654;
    63: op1_02_in04 = reg_0164;
    64: op1_02_in04 = imem00_in[91:88];
    65: op1_02_in04 = imem00_in[71:68];
    67: op1_02_in04 = imem00_in[107:104];
    68: op1_02_in04 = reg_0780;
    69: op1_02_in04 = imem07_in[19:16];
    70: op1_02_in04 = reg_0502;
    71: op1_02_in04 = imem07_in[11:8];
    72: op1_02_in04 = reg_0744;
    74: op1_02_in04 = reg_0121;
    75: op1_02_in04 = reg_0554;
    76: op1_02_in04 = reg_0801;
    77: op1_02_in04 = reg_0370;
    78: op1_02_in04 = imem00_in[75:72];
    79: op1_02_in04 = reg_0696;
    80: op1_02_in04 = reg_0392;
    81: op1_02_in04 = imem02_in[63:60];
    82: op1_02_in04 = imem07_in[7:4];
    83: op1_02_in04 = imem05_in[75:72];
    84: op1_02_in04 = imem00_in[115:112];
    85: op1_02_in04 = imem02_in[87:84];
    86: op1_02_in04 = reg_0327;
    87: op1_02_in04 = reg_0635;
    88: op1_02_in04 = reg_0322;
    89: op1_02_in04 = reg_0685;
    90: op1_02_in04 = imem00_in[103:100];
    92: op1_02_in04 = reg_0302;
    93: op1_02_in04 = reg_0432;
    94: op1_02_in04 = reg_0558;
    96: op1_02_in04 = reg_0540;
    default: op1_02_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv04 = 1;
    3: op1_02_inv04 = 1;
    10: op1_02_inv04 = 1;
    11: op1_02_inv04 = 1;
    12: op1_02_inv04 = 1;
    1: op1_02_inv04 = 1;
    15: op1_02_inv04 = 1;
    16: op1_02_inv04 = 1;
    20: op1_02_inv04 = 1;
    21: op1_02_inv04 = 1;
    25: op1_02_inv04 = 1;
    27: op1_02_inv04 = 1;
    30: op1_02_inv04 = 1;
    31: op1_02_inv04 = 1;
    32: op1_02_inv04 = 1;
    36: op1_02_inv04 = 1;
    37: op1_02_inv04 = 1;
    39: op1_02_inv04 = 1;
    41: op1_02_inv04 = 1;
    42: op1_02_inv04 = 1;
    44: op1_02_inv04 = 1;
    45: op1_02_inv04 = 1;
    46: op1_02_inv04 = 1;
    47: op1_02_inv04 = 1;
    48: op1_02_inv04 = 1;
    51: op1_02_inv04 = 1;
    52: op1_02_inv04 = 1;
    54: op1_02_inv04 = 1;
    55: op1_02_inv04 = 1;
    59: op1_02_inv04 = 1;
    61: op1_02_inv04 = 1;
    63: op1_02_inv04 = 1;
    64: op1_02_inv04 = 1;
    67: op1_02_inv04 = 1;
    68: op1_02_inv04 = 1;
    71: op1_02_inv04 = 1;
    72: op1_02_inv04 = 1;
    73: op1_02_inv04 = 1;
    74: op1_02_inv04 = 1;
    82: op1_02_inv04 = 1;
    84: op1_02_inv04 = 1;
    85: op1_02_inv04 = 1;
    86: op1_02_inv04 = 1;
    88: op1_02_inv04 = 1;
    91: op1_02_inv04 = 1;
    93: op1_02_inv04 = 1;
    94: op1_02_inv04 = 1;
    95: op1_02_inv04 = 1;
    default: op1_02_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in05 = imem03_in[79:76];
    5: op1_02_in05 = reg_0453;
    23: op1_02_in05 = reg_0453;
    6: op1_02_in05 = reg_0529;
    7: op1_02_in05 = imem00_in[107:104];
    8: op1_02_in05 = reg_0338;
    9: op1_02_in05 = reg_0309;
    2: op1_02_in05 = reg_0183;
    86: op1_02_in05 = reg_0183;
    10: op1_02_in05 = reg_0546;
    11: op1_02_in05 = reg_0504;
    12: op1_02_in05 = reg_0369;
    13: op1_02_in05 = reg_0688;
    14: op1_02_in05 = reg_0093;
    15: op1_02_in05 = reg_0560;
    16: op1_02_in05 = reg_0731;
    17: op1_02_in05 = reg_0661;
    19: op1_02_in05 = reg_0661;
    18: op1_02_in05 = imem00_in[71:68];
    20: op1_02_in05 = reg_0609;
    77: op1_02_in05 = reg_0609;
    21: op1_02_in05 = imem02_in[95:92];
    22: op1_02_in05 = reg_0396;
    24: op1_02_in05 = reg_0054;
    25: op1_02_in05 = reg_0371;
    26: op1_02_in05 = reg_0087;
    27: op1_02_in05 = reg_0037;
    28: op1_02_in05 = reg_0349;
    29: op1_02_in05 = reg_0587;
    30: op1_02_in05 = imem07_in[71:68];
    31: op1_02_in05 = reg_0243;
    32: op1_02_in05 = reg_0591;
    33: op1_02_in05 = reg_0547;
    34: op1_02_in05 = imem02_in[99:96];
    35: op1_02_in05 = reg_0698;
    36: op1_02_in05 = imem02_in[23:20];
    37: op1_02_in05 = reg_0392;
    38: op1_02_in05 = reg_0568;
    39: op1_02_in05 = imem06_in[79:76];
    40: op1_02_in05 = reg_0256;
    41: op1_02_in05 = reg_0693;
    45: op1_02_in05 = reg_0693;
    42: op1_02_in05 = imem02_in[31:28];
    43: op1_02_in05 = reg_0398;
    44: op1_02_in05 = imem06_in[67:64];
    46: op1_02_in05 = reg_0578;
    47: op1_02_in05 = reg_0520;
    48: op1_02_in05 = reg_0683;
    49: op1_02_in05 = imem00_in[63:60];
    50: op1_02_in05 = reg_0165;
    51: op1_02_in05 = reg_0736;
    52: op1_02_in05 = reg_0247;
    53: op1_02_in05 = reg_0748;
    54: op1_02_in05 = reg_0623;
    55: op1_02_in05 = reg_0612;
    56: op1_02_in05 = reg_0073;
    57: op1_02_in05 = imem02_in[51:48];
    58: op1_02_in05 = reg_0696;
    59: op1_02_in05 = reg_0013;
    60: op1_02_in05 = reg_0586;
    61: op1_02_in05 = reg_0751;
    62: op1_02_in05 = reg_0775;
    63: op1_02_in05 = reg_0168;
    64: op1_02_in05 = imem00_in[103:100];
    65: op1_02_in05 = imem00_in[119:116];
    66: op1_02_in05 = reg_0681;
    67: op1_02_in05 = imem00_in[115:112];
    68: op1_02_in05 = imem05_in[15:12];
    69: op1_02_in05 = imem07_in[31:28];
    70: op1_02_in05 = reg_0220;
    71: op1_02_in05 = imem07_in[35:32];
    72: op1_02_in05 = reg_0690;
    73: op1_02_in05 = reg_0695;
    74: op1_02_in05 = reg_0678;
    75: op1_02_in05 = reg_0556;
    76: op1_02_in05 = reg_0004;
    78: op1_02_in05 = reg_0694;
    89: op1_02_in05 = reg_0694;
    79: op1_02_in05 = reg_0492;
    80: op1_02_in05 = reg_0584;
    81: op1_02_in05 = reg_0650;
    82: op1_02_in05 = imem07_in[15:12];
    83: op1_02_in05 = imem05_in[83:80];
    84: op1_02_in05 = reg_0455;
    85: op1_02_in05 = imem02_in[107:104];
    87: op1_02_in05 = reg_0333;
    88: op1_02_in05 = reg_0414;
    90: op1_02_in05 = reg_0463;
    91: op1_02_in05 = imem00_in[99:96];
    92: op1_02_in05 = reg_0259;
    93: op1_02_in05 = reg_0631;
    94: op1_02_in05 = reg_0516;
    95: op1_02_in05 = reg_0292;
    96: op1_02_in05 = reg_0770;
    default: op1_02_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv05 = 1;
    7: op1_02_inv05 = 1;
    8: op1_02_inv05 = 1;
    2: op1_02_inv05 = 1;
    13: op1_02_inv05 = 1;
    15: op1_02_inv05 = 1;
    20: op1_02_inv05 = 1;
    22: op1_02_inv05 = 1;
    24: op1_02_inv05 = 1;
    26: op1_02_inv05 = 1;
    28: op1_02_inv05 = 1;
    31: op1_02_inv05 = 1;
    36: op1_02_inv05 = 1;
    39: op1_02_inv05 = 1;
    41: op1_02_inv05 = 1;
    43: op1_02_inv05 = 1;
    44: op1_02_inv05 = 1;
    50: op1_02_inv05 = 1;
    53: op1_02_inv05 = 1;
    54: op1_02_inv05 = 1;
    55: op1_02_inv05 = 1;
    57: op1_02_inv05 = 1;
    60: op1_02_inv05 = 1;
    61: op1_02_inv05 = 1;
    62: op1_02_inv05 = 1;
    63: op1_02_inv05 = 1;
    64: op1_02_inv05 = 1;
    67: op1_02_inv05 = 1;
    69: op1_02_inv05 = 1;
    70: op1_02_inv05 = 1;
    71: op1_02_inv05 = 1;
    73: op1_02_inv05 = 1;
    74: op1_02_inv05 = 1;
    75: op1_02_inv05 = 1;
    76: op1_02_inv05 = 1;
    78: op1_02_inv05 = 1;
    82: op1_02_inv05 = 1;
    83: op1_02_inv05 = 1;
    84: op1_02_inv05 = 1;
    85: op1_02_inv05 = 1;
    87: op1_02_inv05 = 1;
    91: op1_02_inv05 = 1;
    95: op1_02_inv05 = 1;
    default: op1_02_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in06 = imem03_in[99:96];
    5: op1_02_in06 = reg_0461;
    6: op1_02_in06 = reg_0539;
    7: op1_02_in06 = reg_0672;
    8: op1_02_in06 = reg_0335;
    9: op1_02_in06 = reg_0000;
    2: op1_02_in06 = reg_0177;
    10: op1_02_in06 = reg_0531;
    11: op1_02_in06 = reg_0243;
    12: op1_02_in06 = reg_0322;
    13: op1_02_in06 = reg_0687;
    14: op1_02_in06 = reg_0073;
    15: op1_02_in06 = reg_0535;
    16: op1_02_in06 = reg_0721;
    17: op1_02_in06 = reg_0638;
    18: op1_02_in06 = imem00_in[83:80];
    19: op1_02_in06 = reg_0663;
    20: op1_02_in06 = reg_0619;
    21: op1_02_in06 = imem02_in[107:104];
    22: op1_02_in06 = reg_0811;
    23: op1_02_in06 = reg_0457;
    24: op1_02_in06 = reg_0265;
    25: op1_02_in06 = reg_0367;
    26: op1_02_in06 = reg_0294;
    70: op1_02_in06 = reg_0294;
    27: op1_02_in06 = reg_0750;
    28: op1_02_in06 = reg_0344;
    29: op1_02_in06 = reg_0592;
    30: op1_02_in06 = imem07_in[91:88];
    31: op1_02_in06 = reg_0104;
    56: op1_02_in06 = reg_0104;
    32: op1_02_in06 = reg_0581;
    33: op1_02_in06 = reg_0303;
    34: op1_02_in06 = imem02_in[111:108];
    35: op1_02_in06 = reg_0690;
    36: op1_02_in06 = imem02_in[35:32];
    37: op1_02_in06 = reg_0569;
    38: op1_02_in06 = reg_0383;
    39: op1_02_in06 = imem06_in[91:88];
    40: op1_02_in06 = reg_0288;
    41: op1_02_in06 = reg_0683;
    42: op1_02_in06 = imem02_in[43:40];
    43: op1_02_in06 = reg_0396;
    44: op1_02_in06 = imem06_in[71:68];
    45: op1_02_in06 = reg_0676;
    46: op1_02_in06 = reg_0387;
    47: op1_02_in06 = reg_0519;
    48: op1_02_in06 = reg_0681;
    49: op1_02_in06 = imem00_in[71:68];
    50: op1_02_in06 = reg_0162;
    51: op1_02_in06 = reg_0304;
    52: op1_02_in06 = reg_0630;
    53: op1_02_in06 = reg_0576;
    54: op1_02_in06 = imem07_in[11:8];
    55: op1_02_in06 = reg_0744;
    57: op1_02_in06 = imem02_in[71:68];
    58: op1_02_in06 = reg_0686;
    59: op1_02_in06 = reg_0014;
    60: op1_02_in06 = reg_0345;
    61: op1_02_in06 = reg_0573;
    62: op1_02_in06 = reg_0764;
    64: op1_02_in06 = imem00_in[111:108];
    65: op1_02_in06 = reg_0693;
    73: op1_02_in06 = reg_0693;
    66: op1_02_in06 = reg_0694;
    67: op1_02_in06 = reg_0695;
    68: op1_02_in06 = imem05_in[27:24];
    69: op1_02_in06 = imem07_in[35:32];
    71: op1_02_in06 = imem07_in[39:36];
    72: op1_02_in06 = reg_0407;
    74: op1_02_in06 = imem02_in[59:56];
    75: op1_02_in06 = reg_0280;
    76: op1_02_in06 = imem04_in[3:0];
    77: op1_02_in06 = reg_0298;
    78: op1_02_in06 = reg_0612;
    79: op1_02_in06 = reg_0612;
    80: op1_02_in06 = reg_0639;
    81: op1_02_in06 = reg_0534;
    82: op1_02_in06 = imem07_in[59:56];
    83: op1_02_in06 = imem05_in[107:104];
    84: op1_02_in06 = reg_0466;
    85: op1_02_in06 = reg_0086;
    86: op1_02_in06 = reg_0091;
    87: op1_02_in06 = reg_0175;
    88: op1_02_in06 = reg_0590;
    89: op1_02_in06 = reg_0749;
    90: op1_02_in06 = reg_0465;
    91: op1_02_in06 = imem00_in[103:100];
    92: op1_02_in06 = reg_0296;
    93: op1_02_in06 = reg_0302;
    94: op1_02_in06 = reg_0249;
    95: op1_02_in06 = reg_0074;
    96: op1_02_in06 = reg_0757;
    default: op1_02_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv06 = 1;
    7: op1_02_inv06 = 1;
    8: op1_02_inv06 = 1;
    11: op1_02_inv06 = 1;
    16: op1_02_inv06 = 1;
    17: op1_02_inv06 = 1;
    21: op1_02_inv06 = 1;
    22: op1_02_inv06 = 1;
    24: op1_02_inv06 = 1;
    33: op1_02_inv06 = 1;
    34: op1_02_inv06 = 1;
    35: op1_02_inv06 = 1;
    36: op1_02_inv06 = 1;
    37: op1_02_inv06 = 1;
    38: op1_02_inv06 = 1;
    41: op1_02_inv06 = 1;
    42: op1_02_inv06 = 1;
    43: op1_02_inv06 = 1;
    44: op1_02_inv06 = 1;
    45: op1_02_inv06 = 1;
    48: op1_02_inv06 = 1;
    50: op1_02_inv06 = 1;
    51: op1_02_inv06 = 1;
    52: op1_02_inv06 = 1;
    58: op1_02_inv06 = 1;
    60: op1_02_inv06 = 1;
    61: op1_02_inv06 = 1;
    65: op1_02_inv06 = 1;
    67: op1_02_inv06 = 1;
    68: op1_02_inv06 = 1;
    72: op1_02_inv06 = 1;
    73: op1_02_inv06 = 1;
    74: op1_02_inv06 = 1;
    76: op1_02_inv06 = 1;
    79: op1_02_inv06 = 1;
    80: op1_02_inv06 = 1;
    82: op1_02_inv06 = 1;
    83: op1_02_inv06 = 1;
    85: op1_02_inv06 = 1;
    87: op1_02_inv06 = 1;
    88: op1_02_inv06 = 1;
    90: op1_02_inv06 = 1;
    91: op1_02_inv06 = 1;
    95: op1_02_inv06 = 1;
    default: op1_02_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in07 = reg_0582;
    5: op1_02_in07 = reg_0469;
    6: op1_02_in07 = reg_0537;
    7: op1_02_in07 = reg_0679;
    8: op1_02_in07 = reg_0314;
    9: op1_02_in07 = reg_0019;
    2: op1_02_in07 = reg_0164;
    10: op1_02_in07 = reg_0556;
    94: op1_02_in07 = reg_0556;
    11: op1_02_in07 = reg_0118;
    12: op1_02_in07 = reg_0397;
    13: op1_02_in07 = reg_0669;
    14: op1_02_in07 = imem03_in[11:8];
    15: op1_02_in07 = reg_0532;
    16: op1_02_in07 = reg_0714;
    17: op1_02_in07 = reg_0665;
    18: op1_02_in07 = imem00_in[87:84];
    49: op1_02_in07 = imem00_in[87:84];
    19: op1_02_in07 = reg_0352;
    20: op1_02_in07 = reg_0612;
    21: op1_02_in07 = reg_0334;
    22: op1_02_in07 = reg_0007;
    23: op1_02_in07 = reg_0189;
    24: op1_02_in07 = reg_0267;
    25: op1_02_in07 = reg_0033;
    26: op1_02_in07 = reg_0298;
    27: op1_02_in07 = reg_0005;
    28: op1_02_in07 = reg_0358;
    29: op1_02_in07 = reg_0594;
    30: op1_02_in07 = imem07_in[95:92];
    31: op1_02_in07 = reg_0119;
    32: op1_02_in07 = reg_0590;
    33: op1_02_in07 = reg_0053;
    34: op1_02_in07 = reg_0642;
    35: op1_02_in07 = reg_0699;
    36: op1_02_in07 = reg_0653;
    37: op1_02_in07 = reg_0562;
    38: op1_02_in07 = reg_0374;
    39: op1_02_in07 = imem06_in[107:104];
    40: op1_02_in07 = imem05_in[123:120];
    41: op1_02_in07 = reg_0696;
    64: op1_02_in07 = reg_0696;
    42: op1_02_in07 = imem02_in[55:52];
    43: op1_02_in07 = reg_0570;
    44: op1_02_in07 = imem06_in[79:76];
    45: op1_02_in07 = reg_0698;
    78: op1_02_in07 = reg_0698;
    46: op1_02_in07 = reg_0391;
    47: op1_02_in07 = reg_0487;
    48: op1_02_in07 = reg_0672;
    50: op1_02_in07 = reg_0167;
    51: op1_02_in07 = reg_0245;
    52: op1_02_in07 = reg_0624;
    53: op1_02_in07 = reg_0372;
    54: op1_02_in07 = imem07_in[31:28];
    55: op1_02_in07 = reg_0455;
    56: op1_02_in07 = reg_0678;
    57: op1_02_in07 = imem02_in[79:76];
    58: op1_02_in07 = reg_0407;
    59: op1_02_in07 = reg_0015;
    60: op1_02_in07 = reg_0361;
    61: op1_02_in07 = reg_0373;
    62: op1_02_in07 = reg_0520;
    65: op1_02_in07 = reg_0749;
    66: op1_02_in07 = reg_0686;
    67: op1_02_in07 = reg_0494;
    79: op1_02_in07 = reg_0494;
    68: op1_02_in07 = imem05_in[31:28];
    69: op1_02_in07 = imem07_in[83:80];
    70: op1_02_in07 = reg_0504;
    71: op1_02_in07 = imem07_in[47:44];
    72: op1_02_in07 = reg_0463;
    73: op1_02_in07 = reg_0681;
    74: op1_02_in07 = imem02_in[67:64];
    75: op1_02_in07 = reg_0611;
    76: op1_02_in07 = imem04_in[31:28];
    77: op1_02_in07 = reg_0766;
    80: op1_02_in07 = reg_0647;
    81: op1_02_in07 = reg_0621;
    82: op1_02_in07 = imem07_in[87:84];
    83: op1_02_in07 = imem05_in[127:124];
    84: op1_02_in07 = reg_0475;
    85: op1_02_in07 = reg_0702;
    86: op1_02_in07 = reg_0427;
    87: op1_02_in07 = reg_0730;
    88: op1_02_in07 = reg_0096;
    89: op1_02_in07 = reg_0758;
    90: op1_02_in07 = reg_0454;
    91: op1_02_in07 = imem00_in[127:124];
    92: op1_02_in07 = reg_0644;
    93: op1_02_in07 = reg_0627;
    95: op1_02_in07 = reg_0617;
    96: op1_02_in07 = reg_0315;
    default: op1_02_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv07 = 1;
    12: op1_02_inv07 = 1;
    13: op1_02_inv07 = 1;
    14: op1_02_inv07 = 1;
    16: op1_02_inv07 = 1;
    21: op1_02_inv07 = 1;
    23: op1_02_inv07 = 1;
    24: op1_02_inv07 = 1;
    25: op1_02_inv07 = 1;
    27: op1_02_inv07 = 1;
    29: op1_02_inv07 = 1;
    30: op1_02_inv07 = 1;
    32: op1_02_inv07 = 1;
    33: op1_02_inv07 = 1;
    36: op1_02_inv07 = 1;
    38: op1_02_inv07 = 1;
    40: op1_02_inv07 = 1;
    42: op1_02_inv07 = 1;
    45: op1_02_inv07 = 1;
    46: op1_02_inv07 = 1;
    47: op1_02_inv07 = 1;
    48: op1_02_inv07 = 1;
    51: op1_02_inv07 = 1;
    52: op1_02_inv07 = 1;
    55: op1_02_inv07 = 1;
    56: op1_02_inv07 = 1;
    57: op1_02_inv07 = 1;
    59: op1_02_inv07 = 1;
    61: op1_02_inv07 = 1;
    62: op1_02_inv07 = 1;
    64: op1_02_inv07 = 1;
    74: op1_02_inv07 = 1;
    80: op1_02_inv07 = 1;
    82: op1_02_inv07 = 1;
    83: op1_02_inv07 = 1;
    84: op1_02_inv07 = 1;
    85: op1_02_inv07 = 1;
    86: op1_02_inv07 = 1;
    90: op1_02_inv07 = 1;
    91: op1_02_inv07 = 1;
    93: op1_02_inv07 = 1;
    96: op1_02_inv07 = 1;
    default: op1_02_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in08 = reg_0583;
    5: op1_02_in08 = reg_0462;
    6: op1_02_in08 = reg_0301;
    15: op1_02_in08 = reg_0301;
    7: op1_02_in08 = reg_0673;
    8: op1_02_in08 = reg_0083;
    9: op1_02_in08 = reg_0012;
    2: op1_02_in08 = reg_0157;
    10: op1_02_in08 = reg_0304;
    11: op1_02_in08 = reg_0101;
    12: op1_02_in08 = reg_0393;
    13: op1_02_in08 = reg_0453;
    14: op1_02_in08 = imem03_in[19:16];
    16: op1_02_in08 = reg_0729;
    17: op1_02_in08 = reg_0659;
    18: op1_02_in08 = reg_0693;
    19: op1_02_in08 = reg_0358;
    20: op1_02_in08 = reg_0402;
    21: op1_02_in08 = reg_0339;
    22: op1_02_in08 = reg_0810;
    23: op1_02_in08 = reg_0188;
    24: op1_02_in08 = reg_0257;
    25: op1_02_in08 = reg_0039;
    26: op1_02_in08 = reg_0078;
    27: op1_02_in08 = reg_0751;
    28: op1_02_in08 = reg_0359;
    29: op1_02_in08 = reg_0575;
    46: op1_02_in08 = reg_0575;
    30: op1_02_in08 = reg_0717;
    31: op1_02_in08 = reg_0120;
    32: op1_02_in08 = reg_0568;
    33: op1_02_in08 = reg_0054;
    34: op1_02_in08 = reg_0666;
    35: op1_02_in08 = reg_0463;
    36: op1_02_in08 = reg_0661;
    37: op1_02_in08 = reg_0803;
    38: op1_02_in08 = reg_0019;
    39: op1_02_in08 = reg_0289;
    40: op1_02_in08 = reg_0798;
    41: op1_02_in08 = reg_0698;
    73: op1_02_in08 = reg_0698;
    42: op1_02_in08 = imem02_in[59:56];
    43: op1_02_in08 = reg_0808;
    44: op1_02_in08 = imem06_in[87:84];
    45: op1_02_in08 = reg_0684;
    78: op1_02_in08 = reg_0684;
    47: op1_02_in08 = imem05_in[3:0];
    48: op1_02_in08 = reg_0676;
    49: op1_02_in08 = imem00_in[99:96];
    50: op1_02_in08 = reg_0160;
    51: op1_02_in08 = reg_0276;
    52: op1_02_in08 = reg_0298;
    53: op1_02_in08 = reg_0620;
    62: op1_02_in08 = reg_0620;
    54: op1_02_in08 = imem07_in[71:68];
    55: op1_02_in08 = reg_0466;
    56: op1_02_in08 = imem02_in[3:0];
    57: op1_02_in08 = imem02_in[111:108];
    58: op1_02_in08 = reg_0680;
    59: op1_02_in08 = imem04_in[11:8];
    60: op1_02_in08 = reg_0360;
    61: op1_02_in08 = reg_0562;
    64: op1_02_in08 = reg_0694;
    65: op1_02_in08 = reg_0407;
    66: op1_02_in08 = reg_0658;
    67: op1_02_in08 = reg_0460;
    68: op1_02_in08 = imem05_in[75:72];
    69: op1_02_in08 = imem07_in[107:104];
    70: op1_02_in08 = reg_0505;
    71: op1_02_in08 = imem07_in[63:60];
    72: op1_02_in08 = reg_0465;
    74: op1_02_in08 = imem02_in[87:84];
    75: op1_02_in08 = reg_0302;
    76: op1_02_in08 = imem04_in[47:44];
    77: op1_02_in08 = reg_0628;
    79: op1_02_in08 = reg_0247;
    80: op1_02_in08 = reg_0753;
    81: op1_02_in08 = reg_0487;
    82: op1_02_in08 = imem07_in[95:92];
    83: op1_02_in08 = reg_0337;
    84: op1_02_in08 = reg_0470;
    85: op1_02_in08 = reg_0374;
    87: op1_02_in08 = reg_0142;
    88: op1_02_in08 = reg_0540;
    89: op1_02_in08 = reg_0477;
    90: op1_02_in08 = reg_0450;
    91: op1_02_in08 = reg_0697;
    92: op1_02_in08 = imem05_in[7:4];
    93: op1_02_in08 = reg_0050;
    94: op1_02_in08 = reg_0305;
    95: op1_02_in08 = reg_0626;
    96: op1_02_in08 = imem03_in[27:24];
    default: op1_02_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv08 = 1;
    7: op1_02_inv08 = 1;
    8: op1_02_inv08 = 1;
    2: op1_02_inv08 = 1;
    10: op1_02_inv08 = 1;
    14: op1_02_inv08 = 1;
    15: op1_02_inv08 = 1;
    16: op1_02_inv08 = 1;
    17: op1_02_inv08 = 1;
    20: op1_02_inv08 = 1;
    21: op1_02_inv08 = 1;
    24: op1_02_inv08 = 1;
    28: op1_02_inv08 = 1;
    29: op1_02_inv08 = 1;
    30: op1_02_inv08 = 1;
    32: op1_02_inv08 = 1;
    35: op1_02_inv08 = 1;
    37: op1_02_inv08 = 1;
    39: op1_02_inv08 = 1;
    40: op1_02_inv08 = 1;
    43: op1_02_inv08 = 1;
    46: op1_02_inv08 = 1;
    47: op1_02_inv08 = 1;
    48: op1_02_inv08 = 1;
    49: op1_02_inv08 = 1;
    51: op1_02_inv08 = 1;
    52: op1_02_inv08 = 1;
    53: op1_02_inv08 = 1;
    54: op1_02_inv08 = 1;
    55: op1_02_inv08 = 1;
    56: op1_02_inv08 = 1;
    57: op1_02_inv08 = 1;
    58: op1_02_inv08 = 1;
    59: op1_02_inv08 = 1;
    61: op1_02_inv08 = 1;
    64: op1_02_inv08 = 1;
    68: op1_02_inv08 = 1;
    69: op1_02_inv08 = 1;
    71: op1_02_inv08 = 1;
    72: op1_02_inv08 = 1;
    73: op1_02_inv08 = 1;
    77: op1_02_inv08 = 1;
    81: op1_02_inv08 = 1;
    87: op1_02_inv08 = 1;
    89: op1_02_inv08 = 1;
    91: op1_02_inv08 = 1;
    92: op1_02_inv08 = 1;
    93: op1_02_inv08 = 1;
    94: op1_02_inv08 = 1;
    95: op1_02_inv08 = 1;
    96: op1_02_inv08 = 1;
    default: op1_02_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in09 = reg_0568;
    5: op1_02_in09 = reg_0467;
    6: op1_02_in09 = reg_0292;
    7: op1_02_in09 = reg_0687;
    8: op1_02_in09 = reg_0090;
    9: op1_02_in09 = reg_0808;
    2: op1_02_in09 = reg_0173;
    10: op1_02_in09 = reg_0281;
    11: op1_02_in09 = imem02_in[3:0];
    12: op1_02_in09 = reg_0389;
    13: op1_02_in09 = reg_0451;
    72: op1_02_in09 = reg_0451;
    14: op1_02_in09 = imem03_in[47:44];
    15: op1_02_in09 = reg_0283;
    16: op1_02_in09 = reg_0425;
    17: op1_02_in09 = reg_0636;
    18: op1_02_in09 = reg_0676;
    19: op1_02_in09 = reg_0330;
    20: op1_02_in09 = reg_0349;
    21: op1_02_in09 = reg_0342;
    22: op1_02_in09 = imem04_in[15:12];
    23: op1_02_in09 = reg_0207;
    24: op1_02_in09 = reg_0077;
    75: op1_02_in09 = reg_0077;
    25: op1_02_in09 = reg_0753;
    26: op1_02_in09 = reg_0253;
    27: op1_02_in09 = imem07_in[23:20];
    28: op1_02_in09 = reg_0345;
    29: op1_02_in09 = reg_0564;
    30: op1_02_in09 = reg_0709;
    31: op1_02_in09 = reg_0108;
    32: op1_02_in09 = reg_0572;
    33: op1_02_in09 = reg_0274;
    34: op1_02_in09 = reg_0660;
    35: op1_02_in09 = reg_0457;
    36: op1_02_in09 = reg_0639;
    37: op1_02_in09 = reg_0801;
    38: op1_02_in09 = reg_0012;
    39: op1_02_in09 = reg_0817;
    40: op1_02_in09 = reg_0781;
    41: op1_02_in09 = reg_0686;
    42: op1_02_in09 = imem02_in[79:76];
    43: op1_02_in09 = reg_0007;
    44: op1_02_in09 = imem06_in[127:124];
    45: op1_02_in09 = reg_0668;
    46: op1_02_in09 = reg_0385;
    47: op1_02_in09 = imem05_in[7:4];
    48: op1_02_in09 = reg_0684;
    49: op1_02_in09 = imem00_in[123:120];
    50: op1_02_in09 = reg_0163;
    51: op1_02_in09 = reg_0269;
    52: op1_02_in09 = reg_0766;
    53: op1_02_in09 = reg_0368;
    54: op1_02_in09 = imem07_in[79:76];
    55: op1_02_in09 = reg_0479;
    56: op1_02_in09 = imem02_in[35:32];
    57: op1_02_in09 = reg_0637;
    58: op1_02_in09 = reg_0453;
    59: op1_02_in09 = imem04_in[35:32];
    60: op1_02_in09 = reg_0351;
    61: op1_02_in09 = reg_0376;
    62: op1_02_in09 = reg_0642;
    74: op1_02_in09 = reg_0642;
    64: op1_02_in09 = reg_0255;
    65: op1_02_in09 = reg_0680;
    66: op1_02_in09 = reg_0117;
    67: op1_02_in09 = reg_0480;
    68: op1_02_in09 = imem05_in[87:84];
    69: op1_02_in09 = reg_0436;
    70: op1_02_in09 = reg_0105;
    71: op1_02_in09 = imem07_in[99:96];
    73: op1_02_in09 = reg_0689;
    76: op1_02_in09 = imem04_in[55:52];
    77: op1_02_in09 = reg_0519;
    78: op1_02_in09 = reg_0691;
    79: op1_02_in09 = reg_0692;
    80: op1_02_in09 = reg_0304;
    81: op1_02_in09 = reg_0655;
    82: op1_02_in09 = imem07_in[103:100];
    83: op1_02_in09 = reg_0667;
    84: op1_02_in09 = reg_0474;
    85: op1_02_in09 = reg_0341;
    87: op1_02_in09 = reg_0099;
    88: op1_02_in09 = reg_0136;
    89: op1_02_in09 = reg_0472;
    90: op1_02_in09 = reg_0455;
    91: op1_02_in09 = reg_0189;
    92: op1_02_in09 = imem05_in[83:80];
    93: op1_02_in09 = reg_0679;
    95: op1_02_in09 = reg_0679;
    94: op1_02_in09 = reg_0503;
    96: op1_02_in09 = imem03_in[39:36];
    default: op1_02_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv09 = 1;
    6: op1_02_inv09 = 1;
    7: op1_02_inv09 = 1;
    10: op1_02_inv09 = 1;
    14: op1_02_inv09 = 1;
    15: op1_02_inv09 = 1;
    16: op1_02_inv09 = 1;
    17: op1_02_inv09 = 1;
    18: op1_02_inv09 = 1;
    20: op1_02_inv09 = 1;
    21: op1_02_inv09 = 1;
    22: op1_02_inv09 = 1;
    23: op1_02_inv09 = 1;
    24: op1_02_inv09 = 1;
    25: op1_02_inv09 = 1;
    26: op1_02_inv09 = 1;
    27: op1_02_inv09 = 1;
    29: op1_02_inv09 = 1;
    34: op1_02_inv09 = 1;
    35: op1_02_inv09 = 1;
    40: op1_02_inv09 = 1;
    42: op1_02_inv09 = 1;
    44: op1_02_inv09 = 1;
    45: op1_02_inv09 = 1;
    46: op1_02_inv09 = 1;
    48: op1_02_inv09 = 1;
    51: op1_02_inv09 = 1;
    60: op1_02_inv09 = 1;
    67: op1_02_inv09 = 1;
    68: op1_02_inv09 = 1;
    69: op1_02_inv09 = 1;
    71: op1_02_inv09 = 1;
    74: op1_02_inv09 = 1;
    75: op1_02_inv09 = 1;
    77: op1_02_inv09 = 1;
    78: op1_02_inv09 = 1;
    80: op1_02_inv09 = 1;
    82: op1_02_inv09 = 1;
    85: op1_02_inv09 = 1;
    91: op1_02_inv09 = 1;
    93: op1_02_inv09 = 1;
    default: op1_02_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in10 = reg_0569;
    5: op1_02_in10 = reg_0470;
    6: op1_02_in10 = reg_0062;
    7: op1_02_in10 = reg_0451;
    8: op1_02_in10 = imem03_in[31:28];
    9: op1_02_in10 = reg_0803;
    2: op1_02_in10 = reg_0171;
    10: op1_02_in10 = reg_0305;
    11: op1_02_in10 = imem02_in[39:36];
    12: op1_02_in10 = reg_0012;
    13: op1_02_in10 = reg_0455;
    72: op1_02_in10 = reg_0455;
    14: op1_02_in10 = imem03_in[51:48];
    15: op1_02_in10 = reg_0289;
    16: op1_02_in10 = reg_0433;
    17: op1_02_in10 = reg_0663;
    18: op1_02_in10 = reg_0689;
    19: op1_02_in10 = reg_0363;
    20: op1_02_in10 = reg_0403;
    21: op1_02_in10 = reg_0338;
    22: op1_02_in10 = imem04_in[43:40];
    23: op1_02_in10 = reg_0201;
    24: op1_02_in10 = reg_0296;
    25: op1_02_in10 = reg_0812;
    26: op1_02_in10 = reg_0076;
    27: op1_02_in10 = imem07_in[95:92];
    28: op1_02_in10 = reg_0342;
    29: op1_02_in10 = reg_0373;
    30: op1_02_in10 = reg_0727;
    31: op1_02_in10 = reg_0110;
    32: op1_02_in10 = reg_0006;
    33: op1_02_in10 = reg_0534;
    34: op1_02_in10 = reg_0651;
    35: op1_02_in10 = reg_0481;
    36: op1_02_in10 = reg_0638;
    37: op1_02_in10 = reg_0015;
    38: op1_02_in10 = reg_0003;
    39: op1_02_in10 = reg_0371;
    40: op1_02_in10 = reg_0795;
    41: op1_02_in10 = reg_0670;
    48: op1_02_in10 = reg_0670;
    42: op1_02_in10 = imem02_in[119:116];
    43: op1_02_in10 = reg_0806;
    44: op1_02_in10 = reg_0817;
    45: op1_02_in10 = reg_0477;
    46: op1_02_in10 = reg_0562;
    47: op1_02_in10 = imem05_in[39:36];
    49: op1_02_in10 = reg_0693;
    50: op1_02_in10 = reg_0183;
    51: op1_02_in10 = reg_0257;
    52: op1_02_in10 = reg_0612;
    53: op1_02_in10 = reg_0375;
    54: op1_02_in10 = reg_0716;
    71: op1_02_in10 = reg_0716;
    55: op1_02_in10 = reg_0478;
    56: op1_02_in10 = imem02_in[55:52];
    57: op1_02_in10 = reg_0657;
    58: op1_02_in10 = reg_0457;
    90: op1_02_in10 = reg_0457;
    59: op1_02_in10 = imem04_in[59:56];
    60: op1_02_in10 = reg_0323;
    61: op1_02_in10 = reg_0001;
    62: op1_02_in10 = imem07_in[3:0];
    64: op1_02_in10 = reg_0117;
    65: op1_02_in10 = reg_0465;
    66: op1_02_in10 = reg_0463;
    67: op1_02_in10 = reg_0459;
    84: op1_02_in10 = reg_0459;
    68: op1_02_in10 = imem05_in[107:104];
    69: op1_02_in10 = reg_0635;
    70: op1_02_in10 = reg_0125;
    73: op1_02_in10 = reg_0475;
    74: op1_02_in10 = reg_0045;
    75: op1_02_in10 = reg_0629;
    76: op1_02_in10 = imem04_in[79:76];
    77: op1_02_in10 = reg_0578;
    78: op1_02_in10 = reg_0466;
    79: op1_02_in10 = reg_0450;
    80: op1_02_in10 = reg_0702;
    81: op1_02_in10 = reg_0702;
    82: op1_02_in10 = reg_0710;
    83: op1_02_in10 = reg_0666;
    85: op1_02_in10 = reg_0361;
    87: op1_02_in10 = reg_0185;
    88: op1_02_in10 = reg_0098;
    89: op1_02_in10 = reg_0480;
    91: op1_02_in10 = reg_0112;
    92: op1_02_in10 = reg_0227;
    93: op1_02_in10 = reg_0065;
    94: op1_02_in10 = reg_0617;
    95: op1_02_in10 = reg_0622;
    96: op1_02_in10 = imem03_in[83:80];
    default: op1_02_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv10 = 1;
    7: op1_02_inv10 = 1;
    8: op1_02_inv10 = 1;
    9: op1_02_inv10 = 1;
    2: op1_02_inv10 = 1;
    10: op1_02_inv10 = 1;
    13: op1_02_inv10 = 1;
    14: op1_02_inv10 = 1;
    15: op1_02_inv10 = 1;
    16: op1_02_inv10 = 1;
    17: op1_02_inv10 = 1;
    22: op1_02_inv10 = 1;
    23: op1_02_inv10 = 1;
    24: op1_02_inv10 = 1;
    32: op1_02_inv10 = 1;
    33: op1_02_inv10 = 1;
    34: op1_02_inv10 = 1;
    35: op1_02_inv10 = 1;
    36: op1_02_inv10 = 1;
    37: op1_02_inv10 = 1;
    38: op1_02_inv10 = 1;
    40: op1_02_inv10 = 1;
    42: op1_02_inv10 = 1;
    44: op1_02_inv10 = 1;
    46: op1_02_inv10 = 1;
    47: op1_02_inv10 = 1;
    50: op1_02_inv10 = 1;
    51: op1_02_inv10 = 1;
    52: op1_02_inv10 = 1;
    54: op1_02_inv10 = 1;
    55: op1_02_inv10 = 1;
    57: op1_02_inv10 = 1;
    58: op1_02_inv10 = 1;
    60: op1_02_inv10 = 1;
    64: op1_02_inv10 = 1;
    66: op1_02_inv10 = 1;
    67: op1_02_inv10 = 1;
    68: op1_02_inv10 = 1;
    69: op1_02_inv10 = 1;
    70: op1_02_inv10 = 1;
    73: op1_02_inv10 = 1;
    75: op1_02_inv10 = 1;
    76: op1_02_inv10 = 1;
    77: op1_02_inv10 = 1;
    80: op1_02_inv10 = 1;
    81: op1_02_inv10 = 1;
    83: op1_02_inv10 = 1;
    85: op1_02_inv10 = 1;
    87: op1_02_inv10 = 1;
    88: op1_02_inv10 = 1;
    91: op1_02_inv10 = 1;
    95: op1_02_inv10 = 1;
    96: op1_02_inv10 = 1;
    default: op1_02_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in11 = reg_0584;
    5: op1_02_in11 = reg_0474;
    6: op1_02_in11 = reg_0058;
    7: op1_02_in11 = reg_0469;
    45: op1_02_in11 = reg_0469;
    8: op1_02_in11 = imem03_in[47:44];
    9: op1_02_in11 = reg_0801;
    2: op1_02_in11 = reg_0184;
    10: op1_02_in11 = reg_0299;
    11: op1_02_in11 = imem02_in[71:68];
    12: op1_02_in11 = reg_0805;
    13: op1_02_in11 = reg_0461;
    14: op1_02_in11 = imem03_in[67:64];
    15: op1_02_in11 = reg_0290;
    16: op1_02_in11 = reg_0419;
    17: op1_02_in11 = reg_0358;
    18: op1_02_in11 = reg_0684;
    19: op1_02_in11 = reg_0365;
    20: op1_02_in11 = reg_0337;
    21: op1_02_in11 = reg_0518;
    22: op1_02_in11 = imem04_in[99:96];
    23: op1_02_in11 = imem01_in[35:32];
    24: op1_02_in11 = reg_0256;
    25: op1_02_in11 = reg_0035;
    26: op1_02_in11 = reg_0296;
    27: op1_02_in11 = reg_0716;
    28: op1_02_in11 = reg_0092;
    29: op1_02_in11 = reg_0385;
    30: op1_02_in11 = reg_0429;
    31: op1_02_in11 = imem02_in[7:4];
    32: op1_02_in11 = reg_0804;
    33: op1_02_in11 = reg_0529;
    34: op1_02_in11 = reg_0641;
    35: op1_02_in11 = reg_0203;
    36: op1_02_in11 = reg_0636;
    37: op1_02_in11 = reg_0799;
    38: op1_02_in11 = reg_0803;
    39: op1_02_in11 = reg_0618;
    40: op1_02_in11 = reg_0494;
    41: op1_02_in11 = reg_0679;
    42: op1_02_in11 = imem02_in[127:124];
    43: op1_02_in11 = imem04_in[7:4];
    44: op1_02_in11 = reg_0286;
    46: op1_02_in11 = reg_0747;
    47: op1_02_in11 = imem05_in[79:76];
    48: op1_02_in11 = reg_0673;
    49: op1_02_in11 = reg_0672;
    50: op1_02_in11 = reg_0164;
    51: op1_02_in11 = reg_0732;
    52: op1_02_in11 = reg_0318;
    53: op1_02_in11 = reg_0818;
    54: op1_02_in11 = reg_0720;
    55: op1_02_in11 = reg_0189;
    56: op1_02_in11 = imem02_in[59:56];
    57: op1_02_in11 = reg_0651;
    58: op1_02_in11 = reg_0478;
    59: op1_02_in11 = imem04_in[79:76];
    60: op1_02_in11 = reg_0535;
    61: op1_02_in11 = reg_0010;
    62: op1_02_in11 = imem07_in[11:8];
    64: op1_02_in11 = reg_0247;
    65: op1_02_in11 = reg_0475;
    66: op1_02_in11 = reg_0477;
    67: op1_02_in11 = reg_0456;
    68: op1_02_in11 = imem05_in[111:108];
    69: op1_02_in11 = reg_0439;
    70: op1_02_in11 = reg_0120;
    71: op1_02_in11 = reg_0719;
    72: op1_02_in11 = reg_0457;
    73: op1_02_in11 = reg_0460;
    74: op1_02_in11 = reg_0534;
    75: op1_02_in11 = reg_0050;
    76: op1_02_in11 = reg_0544;
    77: op1_02_in11 = reg_0375;
    78: op1_02_in11 = reg_0470;
    79: op1_02_in11 = reg_0451;
    80: op1_02_in11 = reg_0485;
    81: op1_02_in11 = reg_0705;
    82: op1_02_in11 = reg_0162;
    83: op1_02_in11 = reg_0128;
    84: op1_02_in11 = reg_0208;
    85: op1_02_in11 = reg_0343;
    87: op1_02_in11 = reg_0176;
    88: op1_02_in11 = imem03_in[75:72];
    89: op1_02_in11 = reg_0204;
    90: op1_02_in11 = reg_0464;
    91: op1_02_in11 = reg_0688;
    92: op1_02_in11 = reg_0666;
    93: op1_02_in11 = reg_0643;
    94: op1_02_in11 = reg_0610;
    95: op1_02_in11 = reg_0776;
    96: op1_02_in11 = reg_0582;
    default: op1_02_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv11 = 1;
    5: op1_02_inv11 = 1;
    7: op1_02_inv11 = 1;
    8: op1_02_inv11 = 1;
    2: op1_02_inv11 = 1;
    10: op1_02_inv11 = 1;
    11: op1_02_inv11 = 1;
    12: op1_02_inv11 = 1;
    13: op1_02_inv11 = 1;
    20: op1_02_inv11 = 1;
    21: op1_02_inv11 = 1;
    23: op1_02_inv11 = 1;
    25: op1_02_inv11 = 1;
    26: op1_02_inv11 = 1;
    30: op1_02_inv11 = 1;
    31: op1_02_inv11 = 1;
    33: op1_02_inv11 = 1;
    34: op1_02_inv11 = 1;
    36: op1_02_inv11 = 1;
    37: op1_02_inv11 = 1;
    38: op1_02_inv11 = 1;
    40: op1_02_inv11 = 1;
    44: op1_02_inv11 = 1;
    45: op1_02_inv11 = 1;
    46: op1_02_inv11 = 1;
    47: op1_02_inv11 = 1;
    50: op1_02_inv11 = 1;
    51: op1_02_inv11 = 1;
    52: op1_02_inv11 = 1;
    54: op1_02_inv11 = 1;
    56: op1_02_inv11 = 1;
    57: op1_02_inv11 = 1;
    58: op1_02_inv11 = 1;
    59: op1_02_inv11 = 1;
    65: op1_02_inv11 = 1;
    66: op1_02_inv11 = 1;
    68: op1_02_inv11 = 1;
    73: op1_02_inv11 = 1;
    74: op1_02_inv11 = 1;
    80: op1_02_inv11 = 1;
    83: op1_02_inv11 = 1;
    84: op1_02_inv11 = 1;
    85: op1_02_inv11 = 1;
    87: op1_02_inv11 = 1;
    88: op1_02_inv11 = 1;
    91: op1_02_inv11 = 1;
    92: op1_02_inv11 = 1;
    93: op1_02_inv11 = 1;
    default: op1_02_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in12 = reg_0585;
    5: op1_02_in12 = reg_0468;
    65: op1_02_in12 = reg_0468;
    6: op1_02_in12 = reg_0064;
    26: op1_02_in12 = reg_0064;
    7: op1_02_in12 = reg_0480;
    8: op1_02_in12 = imem03_in[87:84];
    9: op1_02_in12 = reg_0014;
    10: op1_02_in12 = reg_0285;
    11: op1_02_in12 = reg_0653;
    12: op1_02_in12 = reg_0008;
    13: op1_02_in12 = reg_0460;
    14: op1_02_in12 = imem03_in[83:80];
    15: op1_02_in12 = reg_0292;
    16: op1_02_in12 = reg_0446;
    17: op1_02_in12 = reg_0320;
    18: op1_02_in12 = reg_0686;
    19: op1_02_in12 = reg_0097;
    20: op1_02_in12 = reg_0401;
    21: op1_02_in12 = reg_0081;
    22: op1_02_in12 = imem04_in[107:104];
    23: op1_02_in12 = imem01_in[47:44];
    24: op1_02_in12 = reg_0288;
    25: op1_02_in12 = reg_0040;
    27: op1_02_in12 = reg_0725;
    28: op1_02_in12 = reg_0541;
    29: op1_02_in12 = reg_0572;
    30: op1_02_in12 = reg_0432;
    31: op1_02_in12 = imem02_in[15:12];
    32: op1_02_in12 = reg_0802;
    33: op1_02_in12 = reg_0290;
    34: op1_02_in12 = reg_0361;
    35: op1_02_in12 = imem01_in[31:28];
    36: op1_02_in12 = reg_0092;
    37: op1_02_in12 = reg_0810;
    38: op1_02_in12 = reg_0801;
    39: op1_02_in12 = reg_0612;
    40: op1_02_in12 = reg_0787;
    41: op1_02_in12 = reg_0675;
    42: op1_02_in12 = reg_0646;
    43: op1_02_in12 = reg_0542;
    44: op1_02_in12 = reg_0339;
    45: op1_02_in12 = reg_0459;
    46: op1_02_in12 = reg_0570;
    47: op1_02_in12 = reg_0792;
    48: op1_02_in12 = reg_0465;
    49: op1_02_in12 = reg_0676;
    50: op1_02_in12 = reg_0168;
    51: op1_02_in12 = reg_0744;
    52: op1_02_in12 = reg_0369;
    53: op1_02_in12 = reg_0029;
    54: op1_02_in12 = reg_0723;
    55: op1_02_in12 = reg_0194;
    56: op1_02_in12 = imem02_in[67:64];
    57: op1_02_in12 = reg_0426;
    58: op1_02_in12 = reg_0458;
    59: op1_02_in12 = imem04_in[119:116];
    60: op1_02_in12 = reg_0539;
    61: op1_02_in12 = imem04_in[7:4];
    62: op1_02_in12 = imem07_in[71:68];
    64: op1_02_in12 = reg_0451;
    66: op1_02_in12 = reg_0476;
    67: op1_02_in12 = reg_0186;
    68: op1_02_in12 = reg_0392;
    69: op1_02_in12 = reg_0180;
    70: op1_02_in12 = reg_0669;
    71: op1_02_in12 = reg_0731;
    72: op1_02_in12 = reg_0477;
    73: op1_02_in12 = reg_0191;
    74: op1_02_in12 = reg_0142;
    75: op1_02_in12 = reg_0626;
    76: op1_02_in12 = reg_0556;
    77: op1_02_in12 = reg_0583;
    78: op1_02_in12 = reg_0452;
    79: op1_02_in12 = reg_0457;
    80: op1_02_in12 = reg_0594;
    81: op1_02_in12 = reg_0275;
    82: op1_02_in12 = reg_0726;
    83: op1_02_in12 = reg_0070;
    84: op1_02_in12 = reg_0193;
    85: op1_02_in12 = reg_0314;
    88: op1_02_in12 = imem03_in[79:76];
    89: op1_02_in12 = reg_0203;
    90: op1_02_in12 = reg_0461;
    91: op1_02_in12 = reg_0455;
    92: op1_02_in12 = reg_0788;
    93: op1_02_in12 = reg_0311;
    94: op1_02_in12 = reg_0301;
    95: op1_02_in12 = imem05_in[7:4];
    96: op1_02_in12 = reg_0003;
    default: op1_02_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv12 = 1;
    7: op1_02_inv12 = 1;
    9: op1_02_inv12 = 1;
    12: op1_02_inv12 = 1;
    13: op1_02_inv12 = 1;
    15: op1_02_inv12 = 1;
    16: op1_02_inv12 = 1;
    19: op1_02_inv12 = 1;
    22: op1_02_inv12 = 1;
    24: op1_02_inv12 = 1;
    25: op1_02_inv12 = 1;
    26: op1_02_inv12 = 1;
    27: op1_02_inv12 = 1;
    29: op1_02_inv12 = 1;
    33: op1_02_inv12 = 1;
    37: op1_02_inv12 = 1;
    38: op1_02_inv12 = 1;
    39: op1_02_inv12 = 1;
    40: op1_02_inv12 = 1;
    41: op1_02_inv12 = 1;
    42: op1_02_inv12 = 1;
    45: op1_02_inv12 = 1;
    46: op1_02_inv12 = 1;
    47: op1_02_inv12 = 1;
    51: op1_02_inv12 = 1;
    52: op1_02_inv12 = 1;
    53: op1_02_inv12 = 1;
    54: op1_02_inv12 = 1;
    56: op1_02_inv12 = 1;
    59: op1_02_inv12 = 1;
    64: op1_02_inv12 = 1;
    68: op1_02_inv12 = 1;
    70: op1_02_inv12 = 1;
    74: op1_02_inv12 = 1;
    76: op1_02_inv12 = 1;
    78: op1_02_inv12 = 1;
    83: op1_02_inv12 = 1;
    84: op1_02_inv12 = 1;
    85: op1_02_inv12 = 1;
    89: op1_02_inv12 = 1;
    91: op1_02_inv12 = 1;
    92: op1_02_inv12 = 1;
    94: op1_02_inv12 = 1;
    95: op1_02_inv12 = 1;
    96: op1_02_inv12 = 1;
    default: op1_02_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in13 = reg_0578;
    5: op1_02_in13 = reg_0459;
    65: op1_02_in13 = reg_0459;
    6: op1_02_in13 = reg_0044;
    7: op1_02_in13 = reg_0468;
    8: op1_02_in13 = imem03_in[103:100];
    9: op1_02_in13 = reg_0805;
    10: op1_02_in13 = reg_0295;
    11: op1_02_in13 = reg_0657;
    12: op1_02_in13 = reg_0009;
    13: op1_02_in13 = reg_0462;
    14: op1_02_in13 = imem03_in[99:96];
    15: op1_02_in13 = reg_0286;
    16: op1_02_in13 = reg_0168;
    17: op1_02_in13 = reg_0363;
    18: op1_02_in13 = reg_0691;
    19: op1_02_in13 = imem03_in[3:0];
    20: op1_02_in13 = reg_0028;
    21: op1_02_in13 = reg_0080;
    28: op1_02_in13 = reg_0080;
    22: op1_02_in13 = imem04_in[123:120];
    23: op1_02_in13 = imem01_in[123:120];
    24: op1_02_in13 = imem05_in[11:8];
    93: op1_02_in13 = imem05_in[11:8];
    25: op1_02_in13 = reg_0814;
    26: op1_02_in13 = reg_0072;
    27: op1_02_in13 = reg_0724;
    29: op1_02_in13 = reg_0804;
    30: op1_02_in13 = reg_0422;
    31: op1_02_in13 = imem02_in[31:28];
    32: op1_02_in13 = reg_0809;
    33: op1_02_in13 = reg_0297;
    34: op1_02_in13 = reg_0351;
    35: op1_02_in13 = imem01_in[35:32];
    36: op1_02_in13 = reg_0541;
    37: op1_02_in13 = imem04_in[15:12];
    38: op1_02_in13 = reg_0008;
    39: op1_02_in13 = reg_0775;
    40: op1_02_in13 = reg_0489;
    41: op1_02_in13 = reg_0688;
    42: op1_02_in13 = reg_0660;
    43: op1_02_in13 = reg_0088;
    44: op1_02_in13 = reg_0278;
    45: op1_02_in13 = reg_0208;
    46: op1_02_in13 = reg_0000;
    47: op1_02_in13 = reg_0482;
    48: op1_02_in13 = reg_0450;
    49: op1_02_in13 = reg_0686;
    50: op1_02_in13 = reg_0170;
    51: op1_02_in13 = reg_0128;
    52: op1_02_in13 = reg_0776;
    53: op1_02_in13 = reg_0367;
    54: op1_02_in13 = reg_0725;
    55: op1_02_in13 = reg_0197;
    56: op1_02_in13 = imem02_in[75:72];
    57: op1_02_in13 = reg_0362;
    58: op1_02_in13 = reg_0214;
    59: op1_02_in13 = reg_0542;
    60: op1_02_in13 = reg_0098;
    61: op1_02_in13 = imem04_in[23:20];
    62: op1_02_in13 = imem07_in[83:80];
    64: op1_02_in13 = reg_0461;
    66: op1_02_in13 = reg_0481;
    67: op1_02_in13 = reg_0212;
    68: op1_02_in13 = reg_0793;
    69: op1_02_in13 = reg_0162;
    70: op1_02_in13 = reg_0676;
    71: op1_02_in13 = reg_0721;
    72: op1_02_in13 = reg_0470;
    73: op1_02_in13 = reg_0190;
    74: op1_02_in13 = reg_0254;
    75: op1_02_in13 = reg_0610;
    76: op1_02_in13 = reg_0429;
    77: op1_02_in13 = reg_0663;
    78: op1_02_in13 = reg_0478;
    79: op1_02_in13 = reg_0475;
    80: op1_02_in13 = reg_0353;
    81: op1_02_in13 = reg_0485;
    82: op1_02_in13 = reg_0784;
    83: op1_02_in13 = reg_0550;
    84: op1_02_in13 = reg_0196;
    85: op1_02_in13 = reg_0540;
    88: op1_02_in13 = imem03_in[95:92];
    89: op1_02_in13 = reg_0211;
    90: op1_02_in13 = reg_0479;
    91: op1_02_in13 = reg_0457;
    92: op1_02_in13 = reg_0641;
    94: op1_02_in13 = reg_0585;
    95: op1_02_in13 = imem05_in[31:28];
    96: op1_02_in13 = reg_0604;
    default: op1_02_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv13 = 1;
    7: op1_02_inv13 = 1;
    8: op1_02_inv13 = 1;
    9: op1_02_inv13 = 1;
    11: op1_02_inv13 = 1;
    12: op1_02_inv13 = 1;
    13: op1_02_inv13 = 1;
    16: op1_02_inv13 = 1;
    17: op1_02_inv13 = 1;
    21: op1_02_inv13 = 1;
    22: op1_02_inv13 = 1;
    24: op1_02_inv13 = 1;
    27: op1_02_inv13 = 1;
    28: op1_02_inv13 = 1;
    29: op1_02_inv13 = 1;
    32: op1_02_inv13 = 1;
    38: op1_02_inv13 = 1;
    42: op1_02_inv13 = 1;
    45: op1_02_inv13 = 1;
    47: op1_02_inv13 = 1;
    48: op1_02_inv13 = 1;
    51: op1_02_inv13 = 1;
    52: op1_02_inv13 = 1;
    53: op1_02_inv13 = 1;
    54: op1_02_inv13 = 1;
    56: op1_02_inv13 = 1;
    57: op1_02_inv13 = 1;
    58: op1_02_inv13 = 1;
    59: op1_02_inv13 = 1;
    64: op1_02_inv13 = 1;
    65: op1_02_inv13 = 1;
    67: op1_02_inv13 = 1;
    70: op1_02_inv13 = 1;
    73: op1_02_inv13 = 1;
    75: op1_02_inv13 = 1;
    76: op1_02_inv13 = 1;
    78: op1_02_inv13 = 1;
    81: op1_02_inv13 = 1;
    89: op1_02_inv13 = 1;
    90: op1_02_inv13 = 1;
    91: op1_02_inv13 = 1;
    92: op1_02_inv13 = 1;
    default: op1_02_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in14 = reg_0570;
    5: op1_02_in14 = reg_0211;
    6: op1_02_in14 = imem05_in[7:4];
    7: op1_02_in14 = reg_0459;
    90: op1_02_in14 = reg_0459;
    8: op1_02_in14 = reg_0598;
    9: op1_02_in14 = reg_0802;
    10: op1_02_in14 = reg_0275;
    11: op1_02_in14 = reg_0661;
    12: op1_02_in14 = reg_0809;
    13: op1_02_in14 = reg_0479;
    14: op1_02_in14 = reg_0573;
    15: op1_02_in14 = reg_0307;
    16: op1_02_in14 = reg_0158;
    17: op1_02_in14 = reg_0088;
    18: op1_02_in14 = reg_0692;
    19: op1_02_in14 = imem03_in[15:12];
    20: op1_02_in14 = reg_0039;
    21: op1_02_in14 = reg_0095;
    28: op1_02_in14 = reg_0095;
    22: op1_02_in14 = reg_0059;
    23: op1_02_in14 = reg_0496;
    24: op1_02_in14 = imem05_in[15:12];
    25: op1_02_in14 = reg_0029;
    26: op1_02_in14 = imem05_in[79:76];
    27: op1_02_in14 = reg_0706;
    29: op1_02_in14 = reg_0015;
    30: op1_02_in14 = reg_0419;
    31: op1_02_in14 = imem02_in[47:44];
    32: op1_02_in14 = imem04_in[7:4];
    33: op1_02_in14 = reg_0078;
    34: op1_02_in14 = reg_0355;
    35: op1_02_in14 = imem01_in[75:72];
    36: op1_02_in14 = reg_0314;
    37: op1_02_in14 = imem04_in[55:52];
    38: op1_02_in14 = reg_0009;
    39: op1_02_in14 = reg_0821;
    40: op1_02_in14 = reg_0736;
    41: op1_02_in14 = reg_0673;
    42: op1_02_in14 = reg_0651;
    43: op1_02_in14 = reg_0523;
    44: op1_02_in14 = reg_0577;
    45: op1_02_in14 = reg_0205;
    46: op1_02_in14 = reg_0019;
    47: op1_02_in14 = reg_0797;
    48: op1_02_in14 = reg_0464;
    49: op1_02_in14 = reg_0670;
    51: op1_02_in14 = reg_0142;
    52: op1_02_in14 = reg_0576;
    53: op1_02_in14 = imem07_in[19:16];
    54: op1_02_in14 = reg_0701;
    55: op1_02_in14 = imem01_in[31:28];
    56: op1_02_in14 = imem02_in[103:100];
    57: op1_02_in14 = reg_0345;
    58: op1_02_in14 = reg_0212;
    59: op1_02_in14 = reg_0055;
    60: op1_02_in14 = reg_0094;
    61: op1_02_in14 = imem04_in[39:36];
    62: op1_02_in14 = imem07_in[95:92];
    64: op1_02_in14 = reg_0481;
    65: op1_02_in14 = reg_0458;
    66: op1_02_in14 = reg_0470;
    67: op1_02_in14 = imem01_in[3:0];
    68: op1_02_in14 = reg_0227;
    69: op1_02_in14 = reg_0169;
    70: op1_02_in14 = reg_0126;
    71: op1_02_in14 = reg_0709;
    72: op1_02_in14 = reg_0452;
    73: op1_02_in14 = reg_0202;
    84: op1_02_in14 = reg_0202;
    74: op1_02_in14 = reg_0584;
    75: op1_02_in14 = imem05_in[55:52];
    76: op1_02_in14 = reg_0432;
    77: op1_02_in14 = reg_0484;
    78: op1_02_in14 = reg_0203;
    79: op1_02_in14 = reg_0199;
    80: op1_02_in14 = reg_0323;
    81: op1_02_in14 = reg_0359;
    82: op1_02_in14 = reg_0160;
    83: op1_02_in14 = reg_0246;
    85: op1_02_in14 = reg_0770;
    88: op1_02_in14 = imem03_in[119:116];
    89: op1_02_in14 = reg_0195;
    91: op1_02_in14 = reg_0476;
    92: op1_02_in14 = reg_0795;
    93: op1_02_in14 = imem05_in[19:16];
    94: op1_02_in14 = reg_0069;
    95: op1_02_in14 = imem05_in[39:36];
    96: op1_02_in14 = reg_0599;
    default: op1_02_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_02_inv14 = 1;
    10: op1_02_inv14 = 1;
    11: op1_02_inv14 = 1;
    12: op1_02_inv14 = 1;
    13: op1_02_inv14 = 1;
    19: op1_02_inv14 = 1;
    20: op1_02_inv14 = 1;
    22: op1_02_inv14 = 1;
    23: op1_02_inv14 = 1;
    25: op1_02_inv14 = 1;
    26: op1_02_inv14 = 1;
    29: op1_02_inv14 = 1;
    30: op1_02_inv14 = 1;
    31: op1_02_inv14 = 1;
    32: op1_02_inv14 = 1;
    33: op1_02_inv14 = 1;
    35: op1_02_inv14 = 1;
    41: op1_02_inv14 = 1;
    42: op1_02_inv14 = 1;
    45: op1_02_inv14 = 1;
    48: op1_02_inv14 = 1;
    49: op1_02_inv14 = 1;
    54: op1_02_inv14 = 1;
    58: op1_02_inv14 = 1;
    59: op1_02_inv14 = 1;
    60: op1_02_inv14 = 1;
    61: op1_02_inv14 = 1;
    62: op1_02_inv14 = 1;
    64: op1_02_inv14 = 1;
    66: op1_02_inv14 = 1;
    69: op1_02_inv14 = 1;
    70: op1_02_inv14 = 1;
    71: op1_02_inv14 = 1;
    74: op1_02_inv14 = 1;
    75: op1_02_inv14 = 1;
    78: op1_02_inv14 = 1;
    80: op1_02_inv14 = 1;
    82: op1_02_inv14 = 1;
    84: op1_02_inv14 = 1;
    89: op1_02_inv14 = 1;
    90: op1_02_inv14 = 1;
    91: op1_02_inv14 = 1;
    93: op1_02_inv14 = 1;
    95: op1_02_inv14 = 1;
    96: op1_02_inv14 = 1;
    default: op1_02_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in15 = reg_0321;
    5: op1_02_in15 = reg_0212;
    6: op1_02_in15 = imem05_in[23:20];
    7: op1_02_in15 = reg_0191;
    8: op1_02_in15 = reg_0586;
    9: op1_02_in15 = reg_0016;
    10: op1_02_in15 = reg_0061;
    11: op1_02_in15 = reg_0643;
    12: op1_02_in15 = imem04_in[103:100];
    13: op1_02_in15 = reg_0478;
    14: op1_02_in15 = reg_0596;
    15: op1_02_in15 = reg_0284;
    17: op1_02_in15 = reg_0081;
    18: op1_02_in15 = reg_0457;
    19: op1_02_in15 = imem03_in[35:32];
    20: op1_02_in15 = reg_0031;
    21: op1_02_in15 = reg_0535;
    36: op1_02_in15 = reg_0535;
    22: op1_02_in15 = reg_0560;
    23: op1_02_in15 = reg_0514;
    24: op1_02_in15 = imem05_in[55:52];
    25: op1_02_in15 = reg_0749;
    26: op1_02_in15 = imem05_in[111:108];
    27: op1_02_in15 = reg_0423;
    30: op1_02_in15 = reg_0423;
    28: op1_02_in15 = reg_0096;
    29: op1_02_in15 = reg_0799;
    96: op1_02_in15 = reg_0799;
    31: op1_02_in15 = imem02_in[51:48];
    32: op1_02_in15 = imem04_in[11:8];
    33: op1_02_in15 = imem05_in[11:8];
    34: op1_02_in15 = reg_0530;
    35: op1_02_in15 = reg_0336;
    37: op1_02_in15 = imem04_in[59:56];
    61: op1_02_in15 = imem04_in[59:56];
    38: op1_02_in15 = imem04_in[23:20];
    39: op1_02_in15 = reg_0404;
    40: op1_02_in15 = reg_0304;
    41: op1_02_in15 = reg_0453;
    42: op1_02_in15 = reg_0647;
    43: op1_02_in15 = reg_0558;
    59: op1_02_in15 = reg_0558;
    44: op1_02_in15 = reg_0377;
    45: op1_02_in15 = reg_0192;
    73: op1_02_in15 = reg_0192;
    46: op1_02_in15 = reg_0007;
    47: op1_02_in15 = reg_0488;
    48: op1_02_in15 = reg_0462;
    49: op1_02_in15 = reg_0677;
    51: op1_02_in15 = reg_0155;
    52: op1_02_in15 = reg_0621;
    53: op1_02_in15 = imem07_in[59:56];
    54: op1_02_in15 = reg_0706;
    55: op1_02_in15 = imem01_in[43:40];
    56: op1_02_in15 = reg_0655;
    57: op1_02_in15 = reg_0353;
    58: op1_02_in15 = imem01_in[15:12];
    60: op1_02_in15 = imem03_in[11:8];
    62: op1_02_in15 = imem07_in[123:120];
    64: op1_02_in15 = reg_0473;
    65: op1_02_in15 = reg_0188;
    66: op1_02_in15 = reg_0452;
    67: op1_02_in15 = imem01_in[47:44];
    68: op1_02_in15 = reg_0782;
    69: op1_02_in15 = reg_0182;
    70: op1_02_in15 = imem02_in[23:20];
    71: op1_02_in15 = reg_0441;
    72: op1_02_in15 = reg_0456;
    74: op1_02_in15 = reg_0753;
    75: op1_02_in15 = imem05_in[59:56];
    76: op1_02_in15 = reg_0052;
    77: op1_02_in15 = reg_0818;
    78: op1_02_in15 = reg_0207;
    79: op1_02_in15 = reg_0197;
    80: op1_02_in15 = reg_0533;
    81: op1_02_in15 = reg_0360;
    82: op1_02_in15 = reg_0708;
    83: op1_02_in15 = reg_0315;
    84: op1_02_in15 = imem01_in[23:20];
    85: op1_02_in15 = reg_0526;
    88: op1_02_in15 = reg_0186;
    89: op1_02_in15 = imem01_in[11:8];
    90: op1_02_in15 = reg_0214;
    91: op1_02_in15 = reg_0475;
    92: op1_02_in15 = reg_0090;
    93: op1_02_in15 = imem05_in[35:32];
    94: op1_02_in15 = reg_0513;
    95: op1_02_in15 = imem05_in[47:44];
    default: op1_02_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv15 = 1;
    6: op1_02_inv15 = 1;
    8: op1_02_inv15 = 1;
    9: op1_02_inv15 = 1;
    11: op1_02_inv15 = 1;
    12: op1_02_inv15 = 1;
    14: op1_02_inv15 = 1;
    15: op1_02_inv15 = 1;
    17: op1_02_inv15 = 1;
    20: op1_02_inv15 = 1;
    22: op1_02_inv15 = 1;
    23: op1_02_inv15 = 1;
    25: op1_02_inv15 = 1;
    26: op1_02_inv15 = 1;
    27: op1_02_inv15 = 1;
    28: op1_02_inv15 = 1;
    29: op1_02_inv15 = 1;
    30: op1_02_inv15 = 1;
    34: op1_02_inv15 = 1;
    35: op1_02_inv15 = 1;
    36: op1_02_inv15 = 1;
    37: op1_02_inv15 = 1;
    39: op1_02_inv15 = 1;
    41: op1_02_inv15 = 1;
    42: op1_02_inv15 = 1;
    44: op1_02_inv15 = 1;
    46: op1_02_inv15 = 1;
    47: op1_02_inv15 = 1;
    49: op1_02_inv15 = 1;
    52: op1_02_inv15 = 1;
    54: op1_02_inv15 = 1;
    55: op1_02_inv15 = 1;
    56: op1_02_inv15 = 1;
    57: op1_02_inv15 = 1;
    61: op1_02_inv15 = 1;
    62: op1_02_inv15 = 1;
    64: op1_02_inv15 = 1;
    67: op1_02_inv15 = 1;
    68: op1_02_inv15 = 1;
    71: op1_02_inv15 = 1;
    74: op1_02_inv15 = 1;
    75: op1_02_inv15 = 1;
    76: op1_02_inv15 = 1;
    78: op1_02_inv15 = 1;
    82: op1_02_inv15 = 1;
    89: op1_02_inv15 = 1;
    93: op1_02_inv15 = 1;
    94: op1_02_inv15 = 1;
    95: op1_02_inv15 = 1;
    96: op1_02_inv15 = 1;
    default: op1_02_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in16 = reg_0343;
    5: op1_02_in16 = imem01_in[27:24];
    84: op1_02_in16 = imem01_in[27:24];
    6: op1_02_in16 = imem05_in[43:40];
    7: op1_02_in16 = imem01_in[19:16];
    8: op1_02_in16 = reg_0571;
    9: op1_02_in16 = reg_0809;
    10: op1_02_in16 = reg_0046;
    11: op1_02_in16 = reg_0665;
    12: op1_02_in16 = imem04_in[115:112];
    13: op1_02_in16 = reg_0204;
    72: op1_02_in16 = reg_0204;
    14: op1_02_in16 = reg_0568;
    15: op1_02_in16 = reg_0054;
    17: op1_02_in16 = reg_0080;
    18: op1_02_in16 = reg_0469;
    41: op1_02_in16 = reg_0469;
    19: op1_02_in16 = imem03_in[47:44];
    60: op1_02_in16 = imem03_in[47:44];
    20: op1_02_in16 = reg_0753;
    21: op1_02_in16 = reg_0757;
    22: op1_02_in16 = reg_0087;
    23: op1_02_in16 = reg_0505;
    24: op1_02_in16 = imem05_in[67:64];
    25: op1_02_in16 = imem07_in[23:20];
    26: op1_02_in16 = imem05_in[115:112];
    27: op1_02_in16 = reg_0442;
    28: op1_02_in16 = reg_0097;
    29: op1_02_in16 = imem04_in[23:20];
    30: op1_02_in16 = reg_0428;
    31: op1_02_in16 = reg_0653;
    32: op1_02_in16 = imem04_in[31:28];
    33: op1_02_in16 = imem05_in[47:44];
    34: op1_02_in16 = reg_0096;
    35: op1_02_in16 = reg_0497;
    36: op1_02_in16 = reg_0756;
    37: op1_02_in16 = imem04_in[71:68];
    38: op1_02_in16 = imem04_in[71:68];
    39: op1_02_in16 = reg_0319;
    40: op1_02_in16 = reg_0279;
    42: op1_02_in16 = reg_0352;
    43: op1_02_in16 = reg_0433;
    76: op1_02_in16 = reg_0433;
    44: op1_02_in16 = reg_0621;
    45: op1_02_in16 = reg_0197;
    46: op1_02_in16 = reg_0806;
    47: op1_02_in16 = reg_0793;
    48: op1_02_in16 = reg_0481;
    91: op1_02_in16 = reg_0481;
    49: op1_02_in16 = reg_0691;
    51: op1_02_in16 = imem06_in[3:0];
    52: op1_02_in16 = reg_0632;
    53: op1_02_in16 = imem07_in[71:68];
    54: op1_02_in16 = reg_0053;
    71: op1_02_in16 = reg_0053;
    55: op1_02_in16 = imem01_in[59:56];
    56: op1_02_in16 = reg_0654;
    57: op1_02_in16 = reg_0527;
    58: op1_02_in16 = imem01_in[39:36];
    79: op1_02_in16 = imem01_in[39:36];
    59: op1_02_in16 = reg_0058;
    61: op1_02_in16 = imem04_in[67:64];
    62: op1_02_in16 = reg_0726;
    64: op1_02_in16 = reg_0471;
    65: op1_02_in16 = imem01_in[83:80];
    67: op1_02_in16 = imem01_in[83:80];
    66: op1_02_in16 = reg_0200;
    68: op1_02_in16 = reg_0322;
    69: op1_02_in16 = reg_0173;
    70: op1_02_in16 = imem02_in[39:36];
    73: op1_02_in16 = imem01_in[23:20];
    74: op1_02_in16 = reg_0607;
    75: op1_02_in16 = imem05_in[71:68];
    77: op1_02_in16 = reg_0661;
    78: op1_02_in16 = reg_0198;
    80: op1_02_in16 = reg_0081;
    81: op1_02_in16 = reg_0594;
    82: op1_02_in16 = reg_0713;
    83: op1_02_in16 = reg_0720;
    85: op1_02_in16 = reg_0532;
    88: op1_02_in16 = reg_0597;
    89: op1_02_in16 = imem01_in[47:44];
    90: op1_02_in16 = reg_0207;
    92: op1_02_in16 = reg_0027;
    93: op1_02_in16 = imem05_in[55:52];
    94: op1_02_in16 = reg_0371;
    95: op1_02_in16 = imem05_in[59:56];
    96: op1_02_in16 = reg_0600;
    default: op1_02_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv16 = 1;
    6: op1_02_inv16 = 1;
    7: op1_02_inv16 = 1;
    9: op1_02_inv16 = 1;
    10: op1_02_inv16 = 1;
    11: op1_02_inv16 = 1;
    12: op1_02_inv16 = 1;
    15: op1_02_inv16 = 1;
    17: op1_02_inv16 = 1;
    18: op1_02_inv16 = 1;
    23: op1_02_inv16 = 1;
    26: op1_02_inv16 = 1;
    27: op1_02_inv16 = 1;
    30: op1_02_inv16 = 1;
    31: op1_02_inv16 = 1;
    34: op1_02_inv16 = 1;
    35: op1_02_inv16 = 1;
    38: op1_02_inv16 = 1;
    40: op1_02_inv16 = 1;
    41: op1_02_inv16 = 1;
    42: op1_02_inv16 = 1;
    46: op1_02_inv16 = 1;
    55: op1_02_inv16 = 1;
    58: op1_02_inv16 = 1;
    59: op1_02_inv16 = 1;
    60: op1_02_inv16 = 1;
    65: op1_02_inv16 = 1;
    68: op1_02_inv16 = 1;
    71: op1_02_inv16 = 1;
    72: op1_02_inv16 = 1;
    75: op1_02_inv16 = 1;
    76: op1_02_inv16 = 1;
    78: op1_02_inv16 = 1;
    79: op1_02_inv16 = 1;
    83: op1_02_inv16 = 1;
    84: op1_02_inv16 = 1;
    85: op1_02_inv16 = 1;
    90: op1_02_inv16 = 1;
    91: op1_02_inv16 = 1;
    92: op1_02_inv16 = 1;
    94: op1_02_inv16 = 1;
    96: op1_02_inv16 = 1;
    default: op1_02_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in17 = reg_0331;
    5: op1_02_in17 = imem01_in[59:56];
    6: op1_02_in17 = imem05_in[47:44];
    7: op1_02_in17 = imem01_in[35:32];
    8: op1_02_in17 = reg_0599;
    9: op1_02_in17 = reg_0004;
    10: op1_02_in17 = reg_0078;
    11: op1_02_in17 = reg_0659;
    12: op1_02_in17 = imem04_in[127:124];
    13: op1_02_in17 = reg_0212;
    14: op1_02_in17 = reg_0591;
    15: op1_02_in17 = reg_0056;
    17: op1_02_in17 = reg_0082;
    18: op1_02_in17 = reg_0462;
    19: op1_02_in17 = imem03_in[71:68];
    20: op1_02_in17 = reg_0036;
    21: op1_02_in17 = reg_0094;
    36: op1_02_in17 = reg_0094;
    22: op1_02_in17 = reg_0057;
    23: op1_02_in17 = reg_0503;
    24: op1_02_in17 = imem05_in[75:72];
    25: op1_02_in17 = imem07_in[79:76];
    26: op1_02_in17 = reg_0792;
    27: op1_02_in17 = reg_0420;
    28: op1_02_in17 = reg_0769;
    29: op1_02_in17 = imem04_in[63:60];
    30: op1_02_in17 = reg_0172;
    31: op1_02_in17 = reg_0637;
    32: op1_02_in17 = imem04_in[71:68];
    33: op1_02_in17 = imem05_in[67:64];
    34: op1_02_in17 = reg_0539;
    35: op1_02_in17 = reg_0513;
    37: op1_02_in17 = imem04_in[95:92];
    38: op1_02_in17 = imem04_in[75:72];
    39: op1_02_in17 = reg_0242;
    40: op1_02_in17 = reg_0742;
    41: op1_02_in17 = reg_0466;
    42: op1_02_in17 = reg_0359;
    43: op1_02_in17 = reg_0615;
    44: op1_02_in17 = reg_0819;
    45: op1_02_in17 = imem01_in[23:20];
    46: op1_02_in17 = imem04_in[7:4];
    47: op1_02_in17 = reg_0794;
    48: op1_02_in17 = reg_0198;
    49: op1_02_in17 = reg_0674;
    51: op1_02_in17 = imem06_in[47:44];
    52: op1_02_in17 = imem07_in[27:24];
    53: op1_02_in17 = reg_0722;
    54: op1_02_in17 = reg_0175;
    55: op1_02_in17 = imem01_in[75:72];
    56: op1_02_in17 = reg_0548;
    57: op1_02_in17 = reg_0590;
    58: op1_02_in17 = imem01_in[47:44];
    59: op1_02_in17 = reg_0500;
    60: op1_02_in17 = imem03_in[119:116];
    61: op1_02_in17 = imem04_in[99:96];
    62: op1_02_in17 = reg_0729;
    64: op1_02_in17 = reg_0479;
    65: op1_02_in17 = imem01_in[107:104];
    66: op1_02_in17 = reg_0204;
    67: op1_02_in17 = imem01_in[95:92];
    68: op1_02_in17 = reg_0326;
    69: op1_02_in17 = reg_0171;
    70: op1_02_in17 = imem02_in[55:52];
    71: op1_02_in17 = reg_0051;
    72: op1_02_in17 = reg_0193;
    73: op1_02_in17 = imem01_in[31:28];
    74: op1_02_in17 = reg_0140;
    75: op1_02_in17 = imem05_in[87:84];
    76: op1_02_in17 = reg_0297;
    77: op1_02_in17 = imem07_in[3:0];
    78: op1_02_in17 = reg_0201;
    79: op1_02_in17 = imem01_in[67:64];
    80: op1_02_in17 = reg_0096;
    81: op1_02_in17 = reg_0353;
    82: op1_02_in17 = reg_0724;
    83: op1_02_in17 = reg_0276;
    84: op1_02_in17 = imem01_in[71:68];
    85: op1_02_in17 = imem03_in[11:8];
    88: op1_02_in17 = reg_0338;
    89: op1_02_in17 = imem01_in[79:76];
    90: op1_02_in17 = imem01_in[103:100];
    91: op1_02_in17 = reg_0191;
    92: op1_02_in17 = reg_0489;
    93: op1_02_in17 = imem05_in[59:56];
    94: op1_02_in17 = reg_0771;
    95: op1_02_in17 = imem05_in[63:60];
    96: op1_02_in17 = reg_0648;
    default: op1_02_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv17 = 1;
    7: op1_02_inv17 = 1;
    9: op1_02_inv17 = 1;
    10: op1_02_inv17 = 1;
    20: op1_02_inv17 = 1;
    21: op1_02_inv17 = 1;
    24: op1_02_inv17 = 1;
    26: op1_02_inv17 = 1;
    27: op1_02_inv17 = 1;
    29: op1_02_inv17 = 1;
    34: op1_02_inv17 = 1;
    35: op1_02_inv17 = 1;
    37: op1_02_inv17 = 1;
    38: op1_02_inv17 = 1;
    39: op1_02_inv17 = 1;
    40: op1_02_inv17 = 1;
    43: op1_02_inv17 = 1;
    44: op1_02_inv17 = 1;
    45: op1_02_inv17 = 1;
    46: op1_02_inv17 = 1;
    47: op1_02_inv17 = 1;
    48: op1_02_inv17 = 1;
    49: op1_02_inv17 = 1;
    52: op1_02_inv17 = 1;
    57: op1_02_inv17 = 1;
    58: op1_02_inv17 = 1;
    59: op1_02_inv17 = 1;
    61: op1_02_inv17 = 1;
    62: op1_02_inv17 = 1;
    66: op1_02_inv17 = 1;
    68: op1_02_inv17 = 1;
    70: op1_02_inv17 = 1;
    72: op1_02_inv17 = 1;
    75: op1_02_inv17 = 1;
    77: op1_02_inv17 = 1;
    80: op1_02_inv17 = 1;
    81: op1_02_inv17 = 1;
    82: op1_02_inv17 = 1;
    83: op1_02_inv17 = 1;
    88: op1_02_inv17 = 1;
    89: op1_02_inv17 = 1;
    90: op1_02_inv17 = 1;
    92: op1_02_inv17 = 1;
    93: op1_02_inv17 = 1;
    94: op1_02_inv17 = 1;
    96: op1_02_inv17 = 1;
    default: op1_02_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in18 = reg_0000;
    5: op1_02_in18 = imem01_in[103:100];
    6: op1_02_in18 = imem05_in[59:56];
    7: op1_02_in18 = imem01_in[43:40];
    8: op1_02_in18 = reg_0591;
    9: op1_02_in18 = imem04_in[79:76];
    10: op1_02_in18 = reg_0062;
    76: op1_02_in18 = reg_0062;
    11: op1_02_in18 = reg_0333;
    71: op1_02_in18 = reg_0333;
    12: op1_02_in18 = reg_0545;
    13: op1_02_in18 = reg_0197;
    14: op1_02_in18 = reg_0594;
    15: op1_02_in18 = reg_0053;
    17: op1_02_in18 = imem03_in[23:20];
    85: op1_02_in18 = imem03_in[23:20];
    18: op1_02_in18 = reg_0472;
    41: op1_02_in18 = reg_0472;
    19: op1_02_in18 = imem03_in[79:76];
    20: op1_02_in18 = reg_0750;
    21: op1_02_in18 = imem03_in[31:28];
    22: op1_02_in18 = reg_0303;
    59: op1_02_in18 = reg_0303;
    23: op1_02_in18 = reg_0243;
    24: op1_02_in18 = imem05_in[111:108];
    25: op1_02_in18 = reg_0719;
    53: op1_02_in18 = reg_0719;
    26: op1_02_in18 = reg_0798;
    27: op1_02_in18 = reg_0431;
    28: op1_02_in18 = imem03_in[3:0];
    29: op1_02_in18 = imem04_in[107:104];
    30: op1_02_in18 = reg_0157;
    31: op1_02_in18 = reg_0659;
    32: op1_02_in18 = imem04_in[95:92];
    33: op1_02_in18 = imem05_in[71:68];
    34: op1_02_in18 = imem03_in[91:88];
    35: op1_02_in18 = reg_0520;
    36: op1_02_in18 = imem03_in[87:84];
    37: op1_02_in18 = imem04_in[111:108];
    38: op1_02_in18 = imem04_in[99:96];
    39: op1_02_in18 = reg_0777;
    40: op1_02_in18 = reg_0260;
    42: op1_02_in18 = reg_0360;
    43: op1_02_in18 = reg_0529;
    44: op1_02_in18 = reg_0029;
    45: op1_02_in18 = imem01_in[63:60];
    46: op1_02_in18 = imem04_in[11:8];
    47: op1_02_in18 = reg_0784;
    48: op1_02_in18 = reg_0190;
    49: op1_02_in18 = reg_0671;
    51: op1_02_in18 = imem06_in[71:68];
    52: op1_02_in18 = imem07_in[43:40];
    54: op1_02_in18 = reg_0172;
    55: op1_02_in18 = imem01_in[87:84];
    56: op1_02_in18 = reg_0364;
    57: op1_02_in18 = reg_0533;
    58: op1_02_in18 = imem01_in[127:124];
    60: op1_02_in18 = reg_0599;
    61: op1_02_in18 = imem04_in[119:116];
    62: op1_02_in18 = reg_0253;
    64: op1_02_in18 = reg_0210;
    65: op1_02_in18 = reg_0820;
    66: op1_02_in18 = reg_0188;
    67: op1_02_in18 = reg_0497;
    90: op1_02_in18 = reg_0497;
    68: op1_02_in18 = reg_0215;
    70: op1_02_in18 = imem02_in[79:76];
    72: op1_02_in18 = reg_0194;
    73: op1_02_in18 = imem01_in[83:80];
    74: op1_02_in18 = reg_0361;
    75: op1_02_in18 = reg_0736;
    77: op1_02_in18 = imem07_in[11:8];
    78: op1_02_in18 = imem01_in[23:20];
    79: op1_02_in18 = imem01_in[95:92];
    80: op1_02_in18 = reg_0093;
    81: op1_02_in18 = reg_0406;
    82: op1_02_in18 = reg_0727;
    83: op1_02_in18 = reg_0138;
    84: op1_02_in18 = imem01_in[79:76];
    88: op1_02_in18 = reg_0494;
    89: op1_02_in18 = imem01_in[99:96];
    91: op1_02_in18 = reg_0199;
    92: op1_02_in18 = reg_0517;
    93: op1_02_in18 = imem05_in[107:104];
    94: op1_02_in18 = imem05_in[15:12];
    95: op1_02_in18 = imem05_in[67:64];
    96: op1_02_in18 = reg_0384;
    default: op1_02_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv18 = 1;
    5: op1_02_inv18 = 1;
    6: op1_02_inv18 = 1;
    7: op1_02_inv18 = 1;
    8: op1_02_inv18 = 1;
    9: op1_02_inv18 = 1;
    11: op1_02_inv18 = 1;
    12: op1_02_inv18 = 1;
    15: op1_02_inv18 = 1;
    18: op1_02_inv18 = 1;
    20: op1_02_inv18 = 1;
    21: op1_02_inv18 = 1;
    22: op1_02_inv18 = 1;
    25: op1_02_inv18 = 1;
    26: op1_02_inv18 = 1;
    28: op1_02_inv18 = 1;
    29: op1_02_inv18 = 1;
    30: op1_02_inv18 = 1;
    31: op1_02_inv18 = 1;
    32: op1_02_inv18 = 1;
    34: op1_02_inv18 = 1;
    35: op1_02_inv18 = 1;
    36: op1_02_inv18 = 1;
    37: op1_02_inv18 = 1;
    38: op1_02_inv18 = 1;
    39: op1_02_inv18 = 1;
    40: op1_02_inv18 = 1;
    41: op1_02_inv18 = 1;
    42: op1_02_inv18 = 1;
    46: op1_02_inv18 = 1;
    48: op1_02_inv18 = 1;
    53: op1_02_inv18 = 1;
    54: op1_02_inv18 = 1;
    57: op1_02_inv18 = 1;
    59: op1_02_inv18 = 1;
    60: op1_02_inv18 = 1;
    61: op1_02_inv18 = 1;
    65: op1_02_inv18 = 1;
    66: op1_02_inv18 = 1;
    67: op1_02_inv18 = 1;
    68: op1_02_inv18 = 1;
    72: op1_02_inv18 = 1;
    74: op1_02_inv18 = 1;
    76: op1_02_inv18 = 1;
    81: op1_02_inv18 = 1;
    82: op1_02_inv18 = 1;
    83: op1_02_inv18 = 1;
    84: op1_02_inv18 = 1;
    85: op1_02_inv18 = 1;
    88: op1_02_inv18 = 1;
    89: op1_02_inv18 = 1;
    90: op1_02_inv18 = 1;
    91: op1_02_inv18 = 1;
    92: op1_02_inv18 = 1;
    94: op1_02_inv18 = 1;
    default: op1_02_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in19 = reg_0001;
    5: op1_02_in19 = reg_0496;
    6: op1_02_in19 = imem05_in[79:76];
    7: op1_02_in19 = imem01_in[51:48];
    8: op1_02_in19 = reg_0589;
    9: op1_02_in19 = imem04_in[87:84];
    10: op1_02_in19 = reg_0065;
    11: op1_02_in19 = reg_0359;
    56: op1_02_in19 = reg_0359;
    12: op1_02_in19 = reg_0532;
    13: op1_02_in19 = imem01_in[11:8];
    14: op1_02_in19 = reg_0576;
    15: op1_02_in19 = reg_0063;
    17: op1_02_in19 = imem03_in[31:28];
    18: op1_02_in19 = reg_0214;
    19: op1_02_in19 = reg_0598;
    20: op1_02_in19 = reg_0751;
    21: op1_02_in19 = imem03_in[43:40];
    22: op1_02_in19 = reg_0283;
    23: op1_02_in19 = reg_0122;
    24: op1_02_in19 = reg_0791;
    25: op1_02_in19 = reg_0730;
    26: op1_02_in19 = reg_0483;
    27: op1_02_in19 = reg_0172;
    28: op1_02_in19 = imem03_in[51:48];
    29: op1_02_in19 = imem04_in[127:124];
    30: op1_02_in19 = reg_0171;
    31: op1_02_in19 = reg_0663;
    32: op1_02_in19 = imem04_in[107:104];
    33: op1_02_in19 = reg_0482;
    34: op1_02_in19 = imem03_in[103:100];
    35: op1_02_in19 = reg_0334;
    36: op1_02_in19 = imem03_in[111:108];
    37: op1_02_in19 = reg_0059;
    38: op1_02_in19 = imem04_in[103:100];
    39: op1_02_in19 = reg_0814;
    40: op1_02_in19 = reg_0277;
    41: op1_02_in19 = reg_0480;
    42: op1_02_in19 = reg_0324;
    43: op1_02_in19 = reg_0071;
    44: op1_02_in19 = imem07_in[3:0];
    45: op1_02_in19 = reg_0825;
    46: op1_02_in19 = imem04_in[71:68];
    47: op1_02_in19 = reg_0309;
    48: op1_02_in19 = imem01_in[23:20];
    49: op1_02_in19 = reg_0463;
    51: op1_02_in19 = imem06_in[119:116];
    52: op1_02_in19 = imem07_in[47:44];
    53: op1_02_in19 = reg_0061;
    54: op1_02_in19 = reg_0163;
    55: op1_02_in19 = imem01_in[95:92];
    57: op1_02_in19 = reg_0096;
    58: op1_02_in19 = reg_0085;
    59: op1_02_in19 = reg_0077;
    60: op1_02_in19 = reg_0319;
    61: op1_02_in19 = imem04_in[123:120];
    62: op1_02_in19 = reg_0067;
    64: op1_02_in19 = reg_0198;
    65: op1_02_in19 = reg_0322;
    66: op1_02_in19 = reg_0207;
    67: op1_02_in19 = reg_0668;
    68: op1_02_in19 = reg_0491;
    70: op1_02_in19 = imem02_in[119:116];
    71: op1_02_in19 = reg_0167;
    72: op1_02_in19 = reg_0213;
    73: op1_02_in19 = imem01_in[107:104];
    74: op1_02_in19 = reg_0343;
    75: op1_02_in19 = reg_0070;
    76: op1_02_in19 = reg_0776;
    77: op1_02_in19 = imem07_in[15:12];
    78: op1_02_in19 = imem01_in[27:24];
    79: op1_02_in19 = reg_0772;
    80: op1_02_in19 = imem03_in[7:4];
    81: op1_02_in19 = reg_0590;
    82: op1_02_in19 = reg_0441;
    83: op1_02_in19 = reg_0278;
    84: op1_02_in19 = imem01_in[115:112];
    85: op1_02_in19 = imem03_in[63:60];
    88: op1_02_in19 = reg_0575;
    96: op1_02_in19 = reg_0575;
    89: op1_02_in19 = reg_0376;
    90: op1_02_in19 = reg_0645;
    91: op1_02_in19 = imem01_in[19:16];
    92: op1_02_in19 = reg_0326;
    93: op1_02_in19 = reg_0736;
    94: op1_02_in19 = imem05_in[39:36];
    95: op1_02_in19 = imem05_in[103:100];
    default: op1_02_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv19 = 1;
    6: op1_02_inv19 = 1;
    8: op1_02_inv19 = 1;
    9: op1_02_inv19 = 1;
    14: op1_02_inv19 = 1;
    15: op1_02_inv19 = 1;
    20: op1_02_inv19 = 1;
    22: op1_02_inv19 = 1;
    23: op1_02_inv19 = 1;
    25: op1_02_inv19 = 1;
    28: op1_02_inv19 = 1;
    32: op1_02_inv19 = 1;
    33: op1_02_inv19 = 1;
    35: op1_02_inv19 = 1;
    36: op1_02_inv19 = 1;
    39: op1_02_inv19 = 1;
    41: op1_02_inv19 = 1;
    42: op1_02_inv19 = 1;
    45: op1_02_inv19 = 1;
    55: op1_02_inv19 = 1;
    57: op1_02_inv19 = 1;
    58: op1_02_inv19 = 1;
    59: op1_02_inv19 = 1;
    60: op1_02_inv19 = 1;
    62: op1_02_inv19 = 1;
    64: op1_02_inv19 = 1;
    68: op1_02_inv19 = 1;
    72: op1_02_inv19 = 1;
    75: op1_02_inv19 = 1;
    77: op1_02_inv19 = 1;
    78: op1_02_inv19 = 1;
    82: op1_02_inv19 = 1;
    83: op1_02_inv19 = 1;
    84: op1_02_inv19 = 1;
    85: op1_02_inv19 = 1;
    90: op1_02_inv19 = 1;
    92: op1_02_inv19 = 1;
    94: op1_02_inv19 = 1;
    default: op1_02_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in20 = reg_0002;
    5: op1_02_in20 = reg_0513;
    6: op1_02_in20 = imem05_in[115:112];
    7: op1_02_in20 = reg_0504;
    8: op1_02_in20 = reg_0594;
    9: op1_02_in20 = imem04_in[111:108];
    10: op1_02_in20 = reg_0058;
    11: op1_02_in20 = reg_0363;
    12: op1_02_in20 = reg_0301;
    13: op1_02_in20 = imem01_in[15:12];
    14: op1_02_in20 = reg_0384;
    15: op1_02_in20 = reg_0074;
    17: op1_02_in20 = imem03_in[63:60];
    18: op1_02_in20 = reg_0210;
    19: op1_02_in20 = reg_0579;
    20: op1_02_in20 = reg_0749;
    21: op1_02_in20 = imem03_in[47:44];
    22: op1_02_in20 = reg_0306;
    23: op1_02_in20 = reg_0124;
    24: op1_02_in20 = reg_0798;
    25: op1_02_in20 = reg_0721;
    26: op1_02_in20 = reg_0494;
    27: op1_02_in20 = reg_0169;
    28: op1_02_in20 = imem03_in[111:108];
    34: op1_02_in20 = imem03_in[111:108];
    29: op1_02_in20 = reg_0537;
    31: op1_02_in20 = reg_0362;
    32: op1_02_in20 = imem04_in[119:116];
    33: op1_02_in20 = reg_0492;
    35: op1_02_in20 = reg_0122;
    36: op1_02_in20 = reg_0601;
    37: op1_02_in20 = reg_0316;
    38: op1_02_in20 = imem04_in[123:120];
    39: op1_02_in20 = reg_0037;
    40: op1_02_in20 = reg_0734;
    41: op1_02_in20 = reg_0468;
    42: op1_02_in20 = reg_0073;
    43: op1_02_in20 = reg_0616;
    44: op1_02_in20 = imem07_in[43:40];
    45: op1_02_in20 = reg_0511;
    46: op1_02_in20 = imem04_in[83:80];
    47: op1_02_in20 = reg_0742;
    48: op1_02_in20 = imem01_in[47:44];
    49: op1_02_in20 = reg_0450;
    51: op1_02_in20 = imem06_in[127:124];
    52: op1_02_in20 = imem07_in[87:84];
    53: op1_02_in20 = reg_0239;
    54: op1_02_in20 = reg_0177;
    55: op1_02_in20 = imem01_in[99:96];
    56: op1_02_in20 = reg_0353;
    57: op1_02_in20 = reg_0757;
    58: op1_02_in20 = reg_0496;
    59: op1_02_in20 = reg_0050;
    60: op1_02_in20 = reg_0357;
    61: op1_02_in20 = reg_0262;
    62: op1_02_in20 = reg_0635;
    82: op1_02_in20 = reg_0635;
    64: op1_02_in20 = reg_0196;
    65: op1_02_in20 = reg_0100;
    66: op1_02_in20 = reg_0212;
    72: op1_02_in20 = reg_0212;
    67: op1_02_in20 = reg_0761;
    68: op1_02_in20 = reg_0040;
    70: op1_02_in20 = reg_0621;
    71: op1_02_in20 = reg_0159;
    73: op1_02_in20 = reg_0085;
    74: op1_02_in20 = reg_0314;
    75: op1_02_in20 = reg_0550;
    76: op1_02_in20 = reg_0109;
    77: op1_02_in20 = imem07_in[51:48];
    78: op1_02_in20 = imem01_in[31:28];
    79: op1_02_in20 = reg_0385;
    80: op1_02_in20 = imem03_in[55:52];
    81: op1_02_in20 = reg_0343;
    83: op1_02_in20 = reg_0288;
    84: op1_02_in20 = imem01_in[123:120];
    85: op1_02_in20 = imem03_in[71:68];
    88: op1_02_in20 = reg_0568;
    89: op1_02_in20 = reg_0112;
    90: op1_02_in20 = reg_0394;
    91: op1_02_in20 = reg_0653;
    92: op1_02_in20 = reg_0518;
    93: op1_02_in20 = reg_0135;
    94: op1_02_in20 = imem05_in[59:56];
    95: op1_02_in20 = reg_0337;
    96: op1_02_in20 = reg_0637;
    default: op1_02_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv20 = 1;
    7: op1_02_inv20 = 1;
    8: op1_02_inv20 = 1;
    9: op1_02_inv20 = 1;
    10: op1_02_inv20 = 1;
    11: op1_02_inv20 = 1;
    17: op1_02_inv20 = 1;
    18: op1_02_inv20 = 1;
    19: op1_02_inv20 = 1;
    20: op1_02_inv20 = 1;
    21: op1_02_inv20 = 1;
    22: op1_02_inv20 = 1;
    27: op1_02_inv20 = 1;
    32: op1_02_inv20 = 1;
    33: op1_02_inv20 = 1;
    35: op1_02_inv20 = 1;
    36: op1_02_inv20 = 1;
    37: op1_02_inv20 = 1;
    40: op1_02_inv20 = 1;
    41: op1_02_inv20 = 1;
    42: op1_02_inv20 = 1;
    43: op1_02_inv20 = 1;
    45: op1_02_inv20 = 1;
    49: op1_02_inv20 = 1;
    55: op1_02_inv20 = 1;
    57: op1_02_inv20 = 1;
    59: op1_02_inv20 = 1;
    62: op1_02_inv20 = 1;
    64: op1_02_inv20 = 1;
    71: op1_02_inv20 = 1;
    79: op1_02_inv20 = 1;
    80: op1_02_inv20 = 1;
    81: op1_02_inv20 = 1;
    84: op1_02_inv20 = 1;
    89: op1_02_inv20 = 1;
    90: op1_02_inv20 = 1;
    91: op1_02_inv20 = 1;
    93: op1_02_inv20 = 1;
    94: op1_02_inv20 = 1;
    95: op1_02_inv20 = 1;
    default: op1_02_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in21 = reg_0003;
    5: op1_02_in21 = reg_0499;
    6: op1_02_in21 = imem05_in[119:116];
    7: op1_02_in21 = reg_0501;
    8: op1_02_in21 = reg_0600;
    36: op1_02_in21 = reg_0600;
    9: op1_02_in21 = reg_0544;
    10: op1_02_in21 = reg_0074;
    11: op1_02_in21 = reg_0353;
    12: op1_02_in21 = reg_0283;
    13: op1_02_in21 = imem01_in[27:24];
    72: op1_02_in21 = imem01_in[27:24];
    14: op1_02_in21 = reg_0387;
    15: op1_02_in21 = imem05_in[15:12];
    17: op1_02_in21 = imem03_in[99:96];
    18: op1_02_in21 = reg_0209;
    19: op1_02_in21 = reg_0568;
    20: op1_02_in21 = imem07_in[7:4];
    21: op1_02_in21 = imem03_in[51:48];
    22: op1_02_in21 = reg_0297;
    23: op1_02_in21 = reg_0118;
    24: op1_02_in21 = reg_0788;
    25: op1_02_in21 = reg_0726;
    26: op1_02_in21 = reg_0495;
    83: op1_02_in21 = reg_0495;
    27: op1_02_in21 = reg_0166;
    28: op1_02_in21 = reg_0579;
    29: op1_02_in21 = reg_0554;
    31: op1_02_in21 = reg_0341;
    32: op1_02_in21 = reg_0553;
    37: op1_02_in21 = reg_0553;
    33: op1_02_in21 = reg_0780;
    34: op1_02_in21 = reg_0598;
    35: op1_02_in21 = reg_0103;
    45: op1_02_in21 = reg_0103;
    38: op1_02_in21 = imem04_in[127:124];
    39: op1_02_in21 = reg_0238;
    40: op1_02_in21 = reg_0285;
    41: op1_02_in21 = reg_0191;
    42: op1_02_in21 = reg_0518;
    43: op1_02_in21 = reg_0503;
    44: op1_02_in21 = imem07_in[47:44];
    46: op1_02_in21 = imem04_in[99:96];
    47: op1_02_in21 = reg_0275;
    48: op1_02_in21 = imem01_in[111:108];
    49: op1_02_in21 = reg_0457;
    51: op1_02_in21 = reg_0289;
    52: op1_02_in21 = imem07_in[119:116];
    53: op1_02_in21 = reg_0440;
    54: op1_02_in21 = reg_0170;
    55: op1_02_in21 = imem01_in[103:100];
    56: op1_02_in21 = reg_0351;
    57: op1_02_in21 = reg_0094;
    58: op1_02_in21 = reg_0652;
    59: op1_02_in21 = reg_0687;
    60: op1_02_in21 = reg_0383;
    61: op1_02_in21 = reg_0043;
    62: op1_02_in21 = reg_0061;
    64: op1_02_in21 = reg_0205;
    65: op1_02_in21 = reg_0321;
    66: op1_02_in21 = imem01_in[59:56];
    67: op1_02_in21 = reg_0765;
    68: op1_02_in21 = reg_0288;
    70: op1_02_in21 = reg_0753;
    71: op1_02_in21 = reg_0169;
    73: op1_02_in21 = reg_0385;
    74: op1_02_in21 = reg_0533;
    75: op1_02_in21 = reg_0231;
    93: op1_02_in21 = reg_0231;
    76: op1_02_in21 = imem05_in[95:92];
    77: op1_02_in21 = imem07_in[91:88];
    78: op1_02_in21 = imem01_in[47:44];
    79: op1_02_in21 = reg_0394;
    80: op1_02_in21 = imem03_in[103:100];
    81: op1_02_in21 = reg_0514;
    82: op1_02_in21 = reg_0445;
    84: op1_02_in21 = reg_0336;
    85: op1_02_in21 = imem03_in[107:104];
    88: op1_02_in21 = reg_0483;
    89: op1_02_in21 = reg_0114;
    90: op1_02_in21 = reg_0101;
    91: op1_02_in21 = reg_0111;
    92: op1_02_in21 = reg_0538;
    94: op1_02_in21 = imem05_in[87:84];
    95: op1_02_in21 = reg_0227;
    96: op1_02_in21 = reg_0396;
    default: op1_02_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv21 = 1;
    5: op1_02_inv21 = 1;
    6: op1_02_inv21 = 1;
    7: op1_02_inv21 = 1;
    8: op1_02_inv21 = 1;
    9: op1_02_inv21 = 1;
    11: op1_02_inv21 = 1;
    12: op1_02_inv21 = 1;
    13: op1_02_inv21 = 1;
    15: op1_02_inv21 = 1;
    17: op1_02_inv21 = 1;
    18: op1_02_inv21 = 1;
    19: op1_02_inv21 = 1;
    20: op1_02_inv21 = 1;
    25: op1_02_inv21 = 1;
    28: op1_02_inv21 = 1;
    31: op1_02_inv21 = 1;
    32: op1_02_inv21 = 1;
    35: op1_02_inv21 = 1;
    39: op1_02_inv21 = 1;
    41: op1_02_inv21 = 1;
    47: op1_02_inv21 = 1;
    48: op1_02_inv21 = 1;
    51: op1_02_inv21 = 1;
    53: op1_02_inv21 = 1;
    54: op1_02_inv21 = 1;
    57: op1_02_inv21 = 1;
    60: op1_02_inv21 = 1;
    61: op1_02_inv21 = 1;
    68: op1_02_inv21 = 1;
    70: op1_02_inv21 = 1;
    71: op1_02_inv21 = 1;
    74: op1_02_inv21 = 1;
    77: op1_02_inv21 = 1;
    78: op1_02_inv21 = 1;
    79: op1_02_inv21 = 1;
    83: op1_02_inv21 = 1;
    85: op1_02_inv21 = 1;
    88: op1_02_inv21 = 1;
    90: op1_02_inv21 = 1;
    91: op1_02_inv21 = 1;
    94: op1_02_inv21 = 1;
    96: op1_02_inv21 = 1;
    default: op1_02_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in22 = reg_0004;
    5: op1_02_in22 = reg_0518;
    6: op1_02_in22 = reg_0792;
    7: op1_02_in22 = reg_0500;
    8: op1_02_in22 = reg_0595;
    9: op1_02_in22 = reg_0545;
    10: op1_02_in22 = reg_0044;
    11: op1_02_in22 = reg_0355;
    12: op1_02_in22 = reg_0294;
    13: op1_02_in22 = imem01_in[95:92];
    14: op1_02_in22 = reg_0321;
    15: op1_02_in22 = imem05_in[19:16];
    17: op1_02_in22 = reg_0596;
    18: op1_02_in22 = reg_0186;
    96: op1_02_in22 = reg_0186;
    19: op1_02_in22 = reg_0569;
    20: op1_02_in22 = imem07_in[19:16];
    21: op1_02_in22 = imem03_in[67:64];
    22: op1_02_in22 = reg_0295;
    23: op1_02_in22 = reg_0125;
    24: op1_02_in22 = reg_0309;
    25: op1_02_in22 = reg_0729;
    26: op1_02_in22 = reg_0782;
    28: op1_02_in22 = reg_0580;
    36: op1_02_in22 = reg_0580;
    29: op1_02_in22 = reg_0057;
    31: op1_02_in22 = reg_0356;
    32: op1_02_in22 = reg_0552;
    33: op1_02_in22 = reg_0304;
    34: op1_02_in22 = reg_0039;
    35: op1_02_in22 = reg_0108;
    37: op1_02_in22 = reg_0083;
    38: op1_02_in22 = reg_0059;
    39: op1_02_in22 = imem07_in[99:96];
    40: op1_02_in22 = reg_0132;
    41: op1_02_in22 = reg_0187;
    42: op1_02_in22 = reg_0743;
    43: op1_02_in22 = reg_0629;
    44: op1_02_in22 = imem07_in[95:92];
    77: op1_02_in22 = imem07_in[95:92];
    45: op1_02_in22 = reg_0111;
    46: op1_02_in22 = imem04_in[123:120];
    47: op1_02_in22 = reg_0744;
    48: op1_02_in22 = reg_0567;
    49: op1_02_in22 = reg_0469;
    51: op1_02_in22 = reg_0624;
    52: op1_02_in22 = reg_0718;
    53: op1_02_in22 = reg_0443;
    62: op1_02_in22 = reg_0443;
    55: op1_02_in22 = imem01_in[111:108];
    56: op1_02_in22 = reg_0514;
    57: op1_02_in22 = imem03_in[31:28];
    58: op1_02_in22 = reg_0760;
    59: op1_02_in22 = reg_0771;
    60: op1_02_in22 = reg_0385;
    61: op1_02_in22 = reg_0556;
    64: op1_02_in22 = reg_0199;
    65: op1_02_in22 = reg_0422;
    66: op1_02_in22 = imem01_in[91:88];
    67: op1_02_in22 = reg_0778;
    68: op1_02_in22 = reg_0307;
    70: op1_02_in22 = reg_0655;
    71: op1_02_in22 = reg_0160;
    72: op1_02_in22 = imem01_in[47:44];
    73: op1_02_in22 = reg_0759;
    79: op1_02_in22 = reg_0759;
    89: op1_02_in22 = reg_0759;
    74: op1_02_in22 = reg_0080;
    75: op1_02_in22 = reg_0665;
    93: op1_02_in22 = reg_0665;
    76: op1_02_in22 = imem05_in[111:108];
    78: op1_02_in22 = imem01_in[67:64];
    80: op1_02_in22 = imem03_in[119:116];
    81: op1_02_in22 = reg_0323;
    82: op1_02_in22 = reg_0434;
    83: op1_02_in22 = reg_0314;
    84: op1_02_in22 = reg_0497;
    85: op1_02_in22 = reg_0317;
    88: op1_02_in22 = reg_0387;
    90: op1_02_in22 = reg_0237;
    91: op1_02_in22 = reg_0102;
    92: op1_02_in22 = reg_0563;
    94: op1_02_in22 = imem05_in[99:96];
    95: op1_02_in22 = reg_0666;
    default: op1_02_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv22 = 1;
    5: op1_02_inv22 = 1;
    7: op1_02_inv22 = 1;
    8: op1_02_inv22 = 1;
    10: op1_02_inv22 = 1;
    11: op1_02_inv22 = 1;
    12: op1_02_inv22 = 1;
    15: op1_02_inv22 = 1;
    17: op1_02_inv22 = 1;
    18: op1_02_inv22 = 1;
    19: op1_02_inv22 = 1;
    21: op1_02_inv22 = 1;
    23: op1_02_inv22 = 1;
    28: op1_02_inv22 = 1;
    29: op1_02_inv22 = 1;
    31: op1_02_inv22 = 1;
    33: op1_02_inv22 = 1;
    35: op1_02_inv22 = 1;
    36: op1_02_inv22 = 1;
    39: op1_02_inv22 = 1;
    40: op1_02_inv22 = 1;
    42: op1_02_inv22 = 1;
    43: op1_02_inv22 = 1;
    44: op1_02_inv22 = 1;
    45: op1_02_inv22 = 1;
    49: op1_02_inv22 = 1;
    52: op1_02_inv22 = 1;
    55: op1_02_inv22 = 1;
    57: op1_02_inv22 = 1;
    58: op1_02_inv22 = 1;
    64: op1_02_inv22 = 1;
    67: op1_02_inv22 = 1;
    70: op1_02_inv22 = 1;
    71: op1_02_inv22 = 1;
    73: op1_02_inv22 = 1;
    75: op1_02_inv22 = 1;
    78: op1_02_inv22 = 1;
    79: op1_02_inv22 = 1;
    80: op1_02_inv22 = 1;
    81: op1_02_inv22 = 1;
    83: op1_02_inv22 = 1;
    88: op1_02_inv22 = 1;
    89: op1_02_inv22 = 1;
    94: op1_02_inv22 = 1;
    96: op1_02_inv22 = 1;
    default: op1_02_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in23 = imem04_in[7:4];
    5: op1_02_in23 = reg_0507;
    6: op1_02_in23 = reg_0483;
    7: op1_02_in23 = reg_0521;
    8: op1_02_in23 = reg_0576;
    9: op1_02_in23 = reg_0530;
    10: op1_02_in23 = imem05_in[7:4];
    11: op1_02_in23 = reg_0328;
    12: op1_02_in23 = reg_0293;
    13: op1_02_in23 = reg_0517;
    14: op1_02_in23 = reg_0360;
    15: op1_02_in23 = imem05_in[87:84];
    17: op1_02_in23 = reg_0599;
    18: op1_02_in23 = reg_0195;
    19: op1_02_in23 = reg_0592;
    20: op1_02_in23 = imem07_in[27:24];
    21: op1_02_in23 = imem03_in[127:124];
    22: op1_02_in23 = reg_0257;
    23: op1_02_in23 = reg_0099;
    24: op1_02_in23 = reg_0275;
    25: op1_02_in23 = reg_0715;
    26: op1_02_in23 = reg_0783;
    28: op1_02_in23 = reg_0590;
    29: op1_02_in23 = reg_0510;
    31: op1_02_in23 = reg_0346;
    32: op1_02_in23 = reg_0537;
    33: op1_02_in23 = reg_0279;
    34: op1_02_in23 = reg_0589;
    85: op1_02_in23 = reg_0589;
    35: op1_02_in23 = reg_0114;
    36: op1_02_in23 = reg_0578;
    37: op1_02_in23 = reg_0057;
    38: op1_02_in23 = reg_0262;
    39: op1_02_in23 = imem07_in[119:116];
    40: op1_02_in23 = reg_0128;
    41: op1_02_in23 = imem01_in[19:16];
    64: op1_02_in23 = imem01_in[19:16];
    42: op1_02_in23 = reg_0757;
    43: op1_02_in23 = reg_0062;
    44: op1_02_in23 = imem07_in[111:108];
    45: op1_02_in23 = reg_0118;
    46: op1_02_in23 = reg_0316;
    47: op1_02_in23 = reg_0734;
    48: op1_02_in23 = reg_0123;
    49: op1_02_in23 = reg_0476;
    51: op1_02_in23 = reg_0817;
    52: op1_02_in23 = reg_0711;
    53: op1_02_in23 = reg_0161;
    55: op1_02_in23 = reg_0646;
    56: op1_02_in23 = reg_0541;
    57: op1_02_in23 = imem03_in[35:32];
    58: op1_02_in23 = reg_0225;
    59: op1_02_in23 = reg_0233;
    60: op1_02_in23 = reg_0569;
    61: op1_02_in23 = reg_0615;
    62: op1_02_in23 = reg_0435;
    65: op1_02_in23 = reg_0220;
    66: op1_02_in23 = imem01_in[107:104];
    67: op1_02_in23 = reg_0418;
    68: op1_02_in23 = reg_0142;
    70: op1_02_in23 = reg_0548;
    71: op1_02_in23 = reg_0168;
    72: op1_02_in23 = imem01_in[59:56];
    73: op1_02_in23 = reg_0778;
    74: op1_02_in23 = reg_0540;
    75: op1_02_in23 = reg_0226;
    76: op1_02_in23 = reg_0027;
    77: op1_02_in23 = imem07_in[99:96];
    78: op1_02_in23 = imem01_in[75:72];
    79: op1_02_in23 = reg_0737;
    80: op1_02_in23 = reg_0582;
    81: op1_02_in23 = reg_0096;
    82: op1_02_in23 = reg_0449;
    83: op1_02_in23 = reg_0277;
    84: op1_02_in23 = reg_0520;
    88: op1_02_in23 = reg_0396;
    89: op1_02_in23 = reg_0258;
    90: op1_02_in23 = reg_0388;
    91: op1_02_in23 = reg_0240;
    92: op1_02_in23 = reg_0495;
    93: op1_02_in23 = reg_0489;
    94: op1_02_in23 = imem05_in[103:100];
    95: op1_02_in23 = reg_0795;
    96: op1_02_in23 = reg_0002;
    default: op1_02_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv23 = 1;
    5: op1_02_inv23 = 1;
    7: op1_02_inv23 = 1;
    9: op1_02_inv23 = 1;
    12: op1_02_inv23 = 1;
    14: op1_02_inv23 = 1;
    17: op1_02_inv23 = 1;
    21: op1_02_inv23 = 1;
    22: op1_02_inv23 = 1;
    24: op1_02_inv23 = 1;
    26: op1_02_inv23 = 1;
    31: op1_02_inv23 = 1;
    32: op1_02_inv23 = 1;
    34: op1_02_inv23 = 1;
    36: op1_02_inv23 = 1;
    37: op1_02_inv23 = 1;
    38: op1_02_inv23 = 1;
    40: op1_02_inv23 = 1;
    43: op1_02_inv23 = 1;
    44: op1_02_inv23 = 1;
    45: op1_02_inv23 = 1;
    53: op1_02_inv23 = 1;
    58: op1_02_inv23 = 1;
    59: op1_02_inv23 = 1;
    60: op1_02_inv23 = 1;
    65: op1_02_inv23 = 1;
    66: op1_02_inv23 = 1;
    67: op1_02_inv23 = 1;
    68: op1_02_inv23 = 1;
    71: op1_02_inv23 = 1;
    72: op1_02_inv23 = 1;
    74: op1_02_inv23 = 1;
    75: op1_02_inv23 = 1;
    76: op1_02_inv23 = 1;
    78: op1_02_inv23 = 1;
    83: op1_02_inv23 = 1;
    84: op1_02_inv23 = 1;
    88: op1_02_inv23 = 1;
    92: op1_02_inv23 = 1;
    94: op1_02_inv23 = 1;
    95: op1_02_inv23 = 1;
    96: op1_02_inv23 = 1;
    default: op1_02_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in24 = imem04_in[11:8];
    5: op1_02_in24 = reg_0508;
    6: op1_02_in24 = reg_0484;
    7: op1_02_in24 = reg_0510;
    8: op1_02_in24 = reg_0321;
    9: op1_02_in24 = reg_0534;
    10: op1_02_in24 = imem05_in[75:72];
    11: op1_02_in24 = reg_0089;
    12: op1_02_in24 = reg_0285;
    13: op1_02_in24 = reg_0778;
    14: op1_02_in24 = reg_0385;
    15: op1_02_in24 = imem05_in[107:104];
    17: op1_02_in24 = reg_0572;
    18: op1_02_in24 = reg_0199;
    19: op1_02_in24 = reg_0563;
    20: op1_02_in24 = imem07_in[43:40];
    21: op1_02_in24 = reg_0586;
    22: op1_02_in24 = reg_0258;
    73: op1_02_in24 = reg_0258;
    23: op1_02_in24 = reg_0107;
    24: op1_02_in24 = reg_0732;
    25: op1_02_in24 = reg_0706;
    26: op1_02_in24 = reg_0090;
    28: op1_02_in24 = reg_0395;
    29: op1_02_in24 = reg_0280;
    31: op1_02_in24 = reg_0355;
    95: op1_02_in24 = reg_0355;
    32: op1_02_in24 = reg_0056;
    33: op1_02_in24 = reg_0735;
    34: op1_02_in24 = reg_0593;
    35: op1_02_in24 = reg_0127;
    36: op1_02_in24 = reg_0595;
    37: op1_02_in24 = reg_0523;
    38: op1_02_in24 = reg_0316;
    39: op1_02_in24 = reg_0719;
    40: op1_02_in24 = reg_0142;
    41: op1_02_in24 = imem01_in[43:40];
    42: op1_02_in24 = reg_0740;
    43: op1_02_in24 = reg_0296;
    44: op1_02_in24 = reg_0720;
    45: op1_02_in24 = reg_0099;
    46: op1_02_in24 = reg_0303;
    47: op1_02_in24 = reg_0136;
    48: op1_02_in24 = reg_0103;
    49: op1_02_in24 = reg_0470;
    51: op1_02_in24 = reg_0286;
    52: op1_02_in24 = reg_0700;
    53: op1_02_in24 = reg_0162;
    55: op1_02_in24 = reg_0772;
    56: op1_02_in24 = reg_0096;
    57: op1_02_in24 = imem03_in[39:36];
    58: op1_02_in24 = reg_0235;
    89: op1_02_in24 = reg_0235;
    59: op1_02_in24 = reg_0644;
    60: op1_02_in24 = reg_0570;
    88: op1_02_in24 = reg_0570;
    61: op1_02_in24 = reg_0302;
    62: op1_02_in24 = reg_0180;
    64: op1_02_in24 = imem01_in[23:20];
    65: op1_02_in24 = reg_0290;
    66: op1_02_in24 = reg_0100;
    67: op1_02_in24 = reg_0424;
    68: op1_02_in24 = reg_0146;
    70: op1_02_in24 = reg_0358;
    72: op1_02_in24 = imem01_in[75:72];
    74: op1_02_in24 = reg_0535;
    75: op1_02_in24 = reg_0326;
    76: op1_02_in24 = reg_0489;
    77: op1_02_in24 = reg_0722;
    78: op1_02_in24 = imem01_in[79:76];
    79: op1_02_in24 = reg_0241;
    80: op1_02_in24 = reg_0579;
    81: op1_02_in24 = reg_0540;
    82: op1_02_in24 = reg_0444;
    83: op1_02_in24 = reg_0383;
    84: op1_02_in24 = reg_0759;
    85: op1_02_in24 = reg_0599;
    90: op1_02_in24 = reg_0422;
    91: op1_02_in24 = reg_0504;
    92: op1_02_in24 = reg_0560;
    93: op1_02_in24 = reg_0552;
    94: op1_02_in24 = imem05_in[119:116];
    96: op1_02_in24 = reg_0418;
    default: op1_02_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv24 = 1;
    7: op1_02_inv24 = 1;
    9: op1_02_inv24 = 1;
    10: op1_02_inv24 = 1;
    12: op1_02_inv24 = 1;
    14: op1_02_inv24 = 1;
    17: op1_02_inv24 = 1;
    18: op1_02_inv24 = 1;
    20: op1_02_inv24 = 1;
    21: op1_02_inv24 = 1;
    23: op1_02_inv24 = 1;
    25: op1_02_inv24 = 1;
    26: op1_02_inv24 = 1;
    32: op1_02_inv24 = 1;
    37: op1_02_inv24 = 1;
    40: op1_02_inv24 = 1;
    41: op1_02_inv24 = 1;
    43: op1_02_inv24 = 1;
    45: op1_02_inv24 = 1;
    49: op1_02_inv24 = 1;
    51: op1_02_inv24 = 1;
    52: op1_02_inv24 = 1;
    53: op1_02_inv24 = 1;
    58: op1_02_inv24 = 1;
    64: op1_02_inv24 = 1;
    65: op1_02_inv24 = 1;
    67: op1_02_inv24 = 1;
    70: op1_02_inv24 = 1;
    75: op1_02_inv24 = 1;
    76: op1_02_inv24 = 1;
    77: op1_02_inv24 = 1;
    78: op1_02_inv24 = 1;
    80: op1_02_inv24 = 1;
    84: op1_02_inv24 = 1;
    85: op1_02_inv24 = 1;
    88: op1_02_inv24 = 1;
    89: op1_02_inv24 = 1;
    91: op1_02_inv24 = 1;
    94: op1_02_inv24 = 1;
    default: op1_02_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in25 = imem04_in[23:20];
    5: op1_02_in25 = reg_0232;
    6: op1_02_in25 = reg_0495;
    7: op1_02_in25 = reg_0226;
    8: op1_02_in25 = reg_0373;
    9: op1_02_in25 = reg_0529;
    10: op1_02_in25 = imem05_in[79:76];
    11: op1_02_in25 = reg_0084;
    12: op1_02_in25 = reg_0286;
    13: op1_02_in25 = reg_0525;
    14: op1_02_in25 = reg_0323;
    15: op1_02_in25 = imem05_in[123:120];
    94: op1_02_in25 = imem05_in[123:120];
    17: op1_02_in25 = reg_0576;
    18: op1_02_in25 = imem01_in[67:64];
    19: op1_02_in25 = reg_0597;
    20: op1_02_in25 = imem07_in[47:44];
    21: op1_02_in25 = reg_0582;
    22: op1_02_in25 = reg_0281;
    23: op1_02_in25 = reg_0127;
    24: op1_02_in25 = reg_0744;
    33: op1_02_in25 = reg_0744;
    25: op1_02_in25 = reg_0727;
    26: op1_02_in25 = reg_0224;
    28: op1_02_in25 = reg_0517;
    29: op1_02_in25 = reg_0268;
    31: op1_02_in25 = reg_0321;
    66: op1_02_in25 = reg_0321;
    32: op1_02_in25 = reg_0536;
    34: op1_02_in25 = reg_0588;
    35: op1_02_in25 = imem02_in[39:36];
    36: op1_02_in25 = reg_0569;
    37: op1_02_in25 = reg_0558;
    38: op1_02_in25 = reg_0060;
    39: op1_02_in25 = reg_0723;
    40: op1_02_in25 = reg_0153;
    41: op1_02_in25 = imem01_in[55:52];
    42: op1_02_in25 = imem03_in[23:20];
    43: op1_02_in25 = reg_0070;
    44: op1_02_in25 = reg_0721;
    45: op1_02_in25 = reg_0108;
    46: op1_02_in25 = reg_0308;
    47: op1_02_in25 = reg_0128;
    48: op1_02_in25 = reg_0104;
    49: op1_02_in25 = reg_0193;
    51: op1_02_in25 = reg_0608;
    52: op1_02_in25 = reg_0064;
    53: op1_02_in25 = reg_0160;
    55: op1_02_in25 = reg_0322;
    56: op1_02_in25 = reg_0770;
    57: op1_02_in25 = imem03_in[47:44];
    58: op1_02_in25 = reg_0241;
    59: op1_02_in25 = reg_0416;
    60: op1_02_in25 = reg_0001;
    88: op1_02_in25 = reg_0001;
    61: op1_02_in25 = reg_0430;
    62: op1_02_in25 = reg_0177;
    64: op1_02_in25 = imem01_in[39:36];
    65: op1_02_in25 = reg_0234;
    67: op1_02_in25 = reg_0073;
    68: op1_02_in25 = imem06_in[31:28];
    70: op1_02_in25 = reg_0362;
    72: op1_02_in25 = imem01_in[79:76];
    73: op1_02_in25 = reg_0421;
    74: op1_02_in25 = reg_0082;
    75: op1_02_in25 = reg_0215;
    76: op1_02_in25 = reg_0099;
    77: op1_02_in25 = reg_0382;
    78: op1_02_in25 = imem01_in[87:84];
    79: op1_02_in25 = reg_0216;
    80: op1_02_in25 = reg_0319;
    81: op1_02_in25 = reg_0538;
    82: op1_02_in25 = reg_0442;
    83: op1_02_in25 = reg_0389;
    84: op1_02_in25 = reg_0397;
    85: op1_02_in25 = reg_0329;
    89: op1_02_in25 = reg_0567;
    90: op1_02_in25 = reg_0603;
    91: op1_02_in25 = reg_0119;
    92: op1_02_in25 = reg_0812;
    93: op1_02_in25 = reg_0797;
    95: op1_02_in25 = reg_0489;
    96: op1_02_in25 = reg_0368;
    default: op1_02_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv25 = 1;
    6: op1_02_inv25 = 1;
    7: op1_02_inv25 = 1;
    9: op1_02_inv25 = 1;
    10: op1_02_inv25 = 1;
    11: op1_02_inv25 = 1;
    13: op1_02_inv25 = 1;
    14: op1_02_inv25 = 1;
    15: op1_02_inv25 = 1;
    17: op1_02_inv25 = 1;
    19: op1_02_inv25 = 1;
    20: op1_02_inv25 = 1;
    22: op1_02_inv25 = 1;
    23: op1_02_inv25 = 1;
    24: op1_02_inv25 = 1;
    33: op1_02_inv25 = 1;
    35: op1_02_inv25 = 1;
    38: op1_02_inv25 = 1;
    39: op1_02_inv25 = 1;
    41: op1_02_inv25 = 1;
    43: op1_02_inv25 = 1;
    46: op1_02_inv25 = 1;
    49: op1_02_inv25 = 1;
    52: op1_02_inv25 = 1;
    55: op1_02_inv25 = 1;
    56: op1_02_inv25 = 1;
    57: op1_02_inv25 = 1;
    60: op1_02_inv25 = 1;
    62: op1_02_inv25 = 1;
    64: op1_02_inv25 = 1;
    65: op1_02_inv25 = 1;
    66: op1_02_inv25 = 1;
    68: op1_02_inv25 = 1;
    70: op1_02_inv25 = 1;
    73: op1_02_inv25 = 1;
    77: op1_02_inv25 = 1;
    79: op1_02_inv25 = 1;
    84: op1_02_inv25 = 1;
    85: op1_02_inv25 = 1;
    89: op1_02_inv25 = 1;
    90: op1_02_inv25 = 1;
    91: op1_02_inv25 = 1;
    92: op1_02_inv25 = 1;
    93: op1_02_inv25 = 1;
    95: op1_02_inv25 = 1;
    96: op1_02_inv25 = 1;
    default: op1_02_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in26 = imem04_in[71:68];
    5: op1_02_in26 = reg_0218;
    6: op1_02_in26 = reg_0783;
    7: op1_02_in26 = reg_0239;
    8: op1_02_in26 = reg_0377;
    9: op1_02_in26 = reg_0548;
    10: op1_02_in26 = reg_0791;
    11: op1_02_in26 = reg_0087;
    12: op1_02_in26 = reg_0307;
    13: op1_02_in26 = reg_0507;
    14: op1_02_in26 = reg_0393;
    15: op1_02_in26 = reg_0482;
    17: op1_02_in26 = reg_0322;
    18: op1_02_in26 = imem01_in[79:76];
    19: op1_02_in26 = reg_0319;
    96: op1_02_in26 = reg_0319;
    20: op1_02_in26 = imem07_in[79:76];
    21: op1_02_in26 = reg_0573;
    22: op1_02_in26 = reg_0078;
    23: op1_02_in26 = reg_0121;
    24: op1_02_in26 = reg_0734;
    55: op1_02_in26 = reg_0734;
    25: op1_02_in26 = reg_0438;
    26: op1_02_in26 = reg_0272;
    28: op1_02_in26 = reg_0562;
    29: op1_02_in26 = reg_0050;
    31: op1_02_in26 = reg_0323;
    32: op1_02_in26 = reg_0516;
    33: op1_02_in26 = reg_0138;
    34: op1_02_in26 = reg_0590;
    35: op1_02_in26 = imem02_in[95:92];
    36: op1_02_in26 = reg_0572;
    37: op1_02_in26 = reg_0556;
    38: op1_02_in26 = reg_0523;
    39: op1_02_in26 = reg_0708;
    40: op1_02_in26 = reg_0137;
    41: op1_02_in26 = reg_0336;
    42: op1_02_in26 = imem03_in[47:44];
    43: op1_02_in26 = imem05_in[3:0];
    59: op1_02_in26 = imem05_in[3:0];
    44: op1_02_in26 = reg_0713;
    45: op1_02_in26 = reg_0109;
    46: op1_02_in26 = reg_0529;
    47: op1_02_in26 = reg_0152;
    48: op1_02_in26 = reg_0117;
    49: op1_02_in26 = reg_0202;
    51: op1_02_in26 = reg_0339;
    52: op1_02_in26 = reg_0266;
    53: op1_02_in26 = reg_0164;
    56: op1_02_in26 = reg_0498;
    57: op1_02_in26 = imem03_in[51:48];
    58: op1_02_in26 = reg_0240;
    60: op1_02_in26 = reg_0003;
    61: op1_02_in26 = reg_0074;
    62: op1_02_in26 = reg_0178;
    64: op1_02_in26 = imem01_in[59:56];
    65: op1_02_in26 = reg_0243;
    66: op1_02_in26 = reg_0241;
    67: op1_02_in26 = reg_0670;
    68: op1_02_in26 = imem06_in[71:68];
    70: op1_02_in26 = reg_0341;
    72: op1_02_in26 = imem01_in[87:84];
    73: op1_02_in26 = reg_0418;
    74: op1_02_in26 = reg_0098;
    75: op1_02_in26 = reg_0786;
    76: op1_02_in26 = reg_0309;
    77: op1_02_in26 = reg_0158;
    78: op1_02_in26 = imem01_in[127:124];
    79: op1_02_in26 = reg_0234;
    90: op1_02_in26 = reg_0234;
    80: op1_02_in26 = reg_0116;
    81: op1_02_in26 = reg_0093;
    82: op1_02_in26 = reg_0139;
    83: op1_02_in26 = reg_0285;
    84: op1_02_in26 = reg_0423;
    85: op1_02_in26 = reg_0600;
    88: op1_02_in26 = reg_0002;
    89: op1_02_in26 = reg_0419;
    91: op1_02_in26 = reg_0106;
    92: op1_02_in26 = reg_0148;
    93: op1_02_in26 = reg_0580;
    94: op1_02_in26 = imem05_in[127:124];
    95: op1_02_in26 = reg_0538;
    default: op1_02_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_02_inv26 = 1;
    9: op1_02_inv26 = 1;
    11: op1_02_inv26 = 1;
    13: op1_02_inv26 = 1;
    14: op1_02_inv26 = 1;
    15: op1_02_inv26 = 1;
    19: op1_02_inv26 = 1;
    25: op1_02_inv26 = 1;
    28: op1_02_inv26 = 1;
    31: op1_02_inv26 = 1;
    32: op1_02_inv26 = 1;
    33: op1_02_inv26 = 1;
    34: op1_02_inv26 = 1;
    37: op1_02_inv26 = 1;
    40: op1_02_inv26 = 1;
    44: op1_02_inv26 = 1;
    45: op1_02_inv26 = 1;
    46: op1_02_inv26 = 1;
    47: op1_02_inv26 = 1;
    48: op1_02_inv26 = 1;
    49: op1_02_inv26 = 1;
    51: op1_02_inv26 = 1;
    52: op1_02_inv26 = 1;
    56: op1_02_inv26 = 1;
    57: op1_02_inv26 = 1;
    58: op1_02_inv26 = 1;
    64: op1_02_inv26 = 1;
    65: op1_02_inv26 = 1;
    66: op1_02_inv26 = 1;
    67: op1_02_inv26 = 1;
    70: op1_02_inv26 = 1;
    72: op1_02_inv26 = 1;
    73: op1_02_inv26 = 1;
    74: op1_02_inv26 = 1;
    75: op1_02_inv26 = 1;
    80: op1_02_inv26 = 1;
    81: op1_02_inv26 = 1;
    84: op1_02_inv26 = 1;
    85: op1_02_inv26 = 1;
    93: op1_02_inv26 = 1;
    94: op1_02_inv26 = 1;
    96: op1_02_inv26 = 1;
    default: op1_02_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in27 = reg_0543;
    5: op1_02_in27 = reg_0242;
    6: op1_02_in27 = reg_0790;
    7: op1_02_in27 = reg_0227;
    8: op1_02_in27 = reg_0006;
    9: op1_02_in27 = reg_0555;
    10: op1_02_in27 = reg_0792;
    11: op1_02_in27 = imem03_in[7:4];
    12: op1_02_in27 = reg_0063;
    13: op1_02_in27 = reg_0232;
    14: op1_02_in27 = reg_0396;
    15: op1_02_in27 = reg_0797;
    17: op1_02_in27 = reg_0374;
    18: op1_02_in27 = imem01_in[111:108];
    19: op1_02_in27 = reg_0019;
    20: op1_02_in27 = imem07_in[91:88];
    21: op1_02_in27 = reg_0587;
    22: op1_02_in27 = reg_0255;
    23: op1_02_in27 = reg_0126;
    24: op1_02_in27 = reg_0135;
    94: op1_02_in27 = reg_0135;
    25: op1_02_in27 = reg_0175;
    26: op1_02_in27 = reg_0089;
    28: op1_02_in27 = reg_0747;
    29: op1_02_in27 = reg_0051;
    52: op1_02_in27 = reg_0051;
    31: op1_02_in27 = reg_0092;
    32: op1_02_in27 = reg_0500;
    33: op1_02_in27 = reg_0140;
    34: op1_02_in27 = reg_0384;
    35: op1_02_in27 = imem02_in[99:96];
    36: op1_02_in27 = reg_0376;
    37: op1_02_in27 = reg_0280;
    38: op1_02_in27 = reg_0558;
    39: op1_02_in27 = reg_0425;
    40: op1_02_in27 = reg_0134;
    41: op1_02_in27 = reg_0497;
    42: op1_02_in27 = imem03_in[91:88];
    43: op1_02_in27 = imem05_in[39:36];
    44: op1_02_in27 = reg_0701;
    45: op1_02_in27 = imem02_in[19:16];
    46: op1_02_in27 = reg_0292;
    47: op1_02_in27 = reg_0156;
    48: op1_02_in27 = imem02_in[51:48];
    49: op1_02_in27 = imem01_in[3:0];
    51: op1_02_in27 = reg_0622;
    55: op1_02_in27 = reg_0737;
    56: op1_02_in27 = reg_0526;
    57: op1_02_in27 = imem03_in[103:100];
    58: op1_02_in27 = reg_0506;
    59: op1_02_in27 = imem05_in[19:16];
    60: op1_02_in27 = reg_0803;
    61: op1_02_in27 = reg_0627;
    62: op1_02_in27 = reg_0158;
    64: op1_02_in27 = imem01_in[67:64];
    65: op1_02_in27 = reg_0125;
    66: op1_02_in27 = reg_0567;
    67: op1_02_in27 = reg_0660;
    68: op1_02_in27 = reg_0815;
    70: op1_02_in27 = reg_0345;
    72: op1_02_in27 = imem01_in[103:100];
    73: op1_02_in27 = reg_0217;
    74: op1_02_in27 = imem03_in[3:0];
    75: op1_02_in27 = reg_0486;
    76: op1_02_in27 = reg_0229;
    77: op1_02_in27 = reg_0334;
    78: op1_02_in27 = reg_0085;
    79: op1_02_in27 = reg_0124;
    80: op1_02_in27 = reg_0350;
    81: op1_02_in27 = imem03_in[55:52];
    82: op1_02_in27 = reg_0116;
    83: op1_02_in27 = reg_0148;
    84: op1_02_in27 = reg_0422;
    85: op1_02_in27 = reg_0488;
    88: op1_02_in27 = reg_0014;
    89: op1_02_in27 = reg_0243;
    90: op1_02_in27 = reg_0504;
    91: op1_02_in27 = imem02_in[31:28];
    92: op1_02_in27 = reg_0781;
    93: op1_02_in27 = reg_0751;
    95: op1_02_in27 = reg_0563;
    96: op1_02_in27 = reg_0306;
    default: op1_02_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv27 = 1;
    5: op1_02_inv27 = 1;
    6: op1_02_inv27 = 1;
    7: op1_02_inv27 = 1;
    9: op1_02_inv27 = 1;
    11: op1_02_inv27 = 1;
    12: op1_02_inv27 = 1;
    20: op1_02_inv27 = 1;
    33: op1_02_inv27 = 1;
    35: op1_02_inv27 = 1;
    37: op1_02_inv27 = 1;
    40: op1_02_inv27 = 1;
    44: op1_02_inv27 = 1;
    46: op1_02_inv27 = 1;
    49: op1_02_inv27 = 1;
    52: op1_02_inv27 = 1;
    55: op1_02_inv27 = 1;
    59: op1_02_inv27 = 1;
    64: op1_02_inv27 = 1;
    65: op1_02_inv27 = 1;
    66: op1_02_inv27 = 1;
    67: op1_02_inv27 = 1;
    73: op1_02_inv27 = 1;
    76: op1_02_inv27 = 1;
    77: op1_02_inv27 = 1;
    78: op1_02_inv27 = 1;
    80: op1_02_inv27 = 1;
    81: op1_02_inv27 = 1;
    82: op1_02_inv27 = 1;
    83: op1_02_inv27 = 1;
    84: op1_02_inv27 = 1;
    85: op1_02_inv27 = 1;
    89: op1_02_inv27 = 1;
    90: op1_02_inv27 = 1;
    91: op1_02_inv27 = 1;
    93: op1_02_inv27 = 1;
    default: op1_02_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in28 = reg_0544;
    5: op1_02_in28 = reg_0240;
    6: op1_02_in28 = reg_0251;
    7: op1_02_in28 = reg_0105;
    8: op1_02_in28 = reg_0019;
    9: op1_02_in28 = reg_0531;
    10: op1_02_in28 = reg_0789;
    11: op1_02_in28 = imem03_in[87:84];
    12: op1_02_in28 = reg_0070;
    13: op1_02_in28 = reg_0217;
    14: op1_02_in28 = reg_0309;
    15: op1_02_in28 = reg_0780;
    17: op1_02_in28 = reg_0331;
    18: op1_02_in28 = reg_0501;
    19: op1_02_in28 = reg_0811;
    20: op1_02_in28 = imem07_in[95:92];
    21: op1_02_in28 = reg_0594;
    22: op1_02_in28 = reg_0071;
    23: op1_02_in28 = imem02_in[55:52];
    24: op1_02_in28 = reg_0142;
    25: op1_02_in28 = reg_0179;
    26: op1_02_in28 = reg_0128;
    28: op1_02_in28 = reg_0374;
    29: op1_02_in28 = reg_0278;
    31: op1_02_in28 = reg_0314;
    32: op1_02_in28 = reg_0556;
    33: op1_02_in28 = imem06_in[27:24];
    34: op1_02_in28 = reg_0389;
    35: op1_02_in28 = imem02_in[103:100];
    36: op1_02_in28 = reg_0397;
    37: op1_02_in28 = reg_0297;
    38: op1_02_in28 = reg_0058;
    39: op1_02_in28 = reg_0423;
    40: op1_02_in28 = reg_0144;
    41: op1_02_in28 = reg_0513;
    42: op1_02_in28 = imem03_in[99:96];
    43: op1_02_in28 = imem05_in[63:60];
    44: op1_02_in28 = reg_0239;
    45: op1_02_in28 = imem02_in[23:20];
    46: op1_02_in28 = reg_0626;
    47: op1_02_in28 = reg_0130;
    48: op1_02_in28 = imem02_in[71:68];
    49: op1_02_in28 = imem01_in[19:16];
    51: op1_02_in28 = reg_0318;
    52: op1_02_in28 = reg_0175;
    55: op1_02_in28 = reg_0550;
    56: op1_02_in28 = reg_0093;
    57: op1_02_in28 = imem03_in[111:108];
    58: op1_02_in28 = reg_0424;
    90: op1_02_in28 = reg_0424;
    59: op1_02_in28 = imem05_in[43:40];
    60: op1_02_in28 = reg_0013;
    61: op1_02_in28 = reg_0585;
    62: op1_02_in28 = reg_0184;
    64: op1_02_in28 = imem01_in[71:68];
    65: op1_02_in28 = reg_0108;
    66: op1_02_in28 = reg_0603;
    67: op1_02_in28 = reg_0107;
    68: op1_02_in28 = reg_0409;
    70: op1_02_in28 = reg_0356;
    72: op1_02_in28 = reg_0085;
    73: op1_02_in28 = reg_0122;
    74: op1_02_in28 = imem03_in[39:36];
    75: op1_02_in28 = reg_0154;
    76: op1_02_in28 = reg_0288;
    77: op1_02_in28 = reg_0442;
    78: op1_02_in28 = reg_0772;
    79: op1_02_in28 = reg_0673;
    80: op1_02_in28 = reg_0281;
    81: op1_02_in28 = imem03_in[91:88];
    82: op1_02_in28 = reg_0110;
    83: op1_02_in28 = reg_0785;
    84: op1_02_in28 = reg_0504;
    85: op1_02_in28 = reg_0403;
    88: op1_02_in28 = reg_0806;
    89: op1_02_in28 = reg_0601;
    91: op1_02_in28 = imem02_in[79:76];
    92: op1_02_in28 = reg_0150;
    93: op1_02_in28 = reg_0254;
    94: op1_02_in28 = reg_0793;
    95: op1_02_in28 = reg_0245;
    96: op1_02_in28 = reg_0294;
    default: op1_02_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv28 = 1;
    7: op1_02_inv28 = 1;
    8: op1_02_inv28 = 1;
    9: op1_02_inv28 = 1;
    11: op1_02_inv28 = 1;
    19: op1_02_inv28 = 1;
    26: op1_02_inv28 = 1;
    29: op1_02_inv28 = 1;
    31: op1_02_inv28 = 1;
    32: op1_02_inv28 = 1;
    37: op1_02_inv28 = 1;
    38: op1_02_inv28 = 1;
    39: op1_02_inv28 = 1;
    40: op1_02_inv28 = 1;
    41: op1_02_inv28 = 1;
    47: op1_02_inv28 = 1;
    49: op1_02_inv28 = 1;
    52: op1_02_inv28 = 1;
    56: op1_02_inv28 = 1;
    57: op1_02_inv28 = 1;
    58: op1_02_inv28 = 1;
    59: op1_02_inv28 = 1;
    61: op1_02_inv28 = 1;
    62: op1_02_inv28 = 1;
    65: op1_02_inv28 = 1;
    74: op1_02_inv28 = 1;
    75: op1_02_inv28 = 1;
    81: op1_02_inv28 = 1;
    84: op1_02_inv28 = 1;
    91: op1_02_inv28 = 1;
    96: op1_02_inv28 = 1;
    default: op1_02_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in29 = reg_0545;
    5: op1_02_in29 = reg_0227;
    6: op1_02_in29 = reg_0223;
    7: op1_02_in29 = reg_0124;
    58: op1_02_in29 = reg_0124;
    8: op1_02_in29 = imem04_in[7:4];
    9: op1_02_in29 = reg_0556;
    10: op1_02_in29 = reg_0793;
    11: op1_02_in29 = imem03_in[91:88];
    12: op1_02_in29 = imem05_in[15:12];
    13: op1_02_in29 = reg_0248;
    14: op1_02_in29 = reg_0374;
    15: op1_02_in29 = reg_0495;
    17: op1_02_in29 = reg_0001;
    18: op1_02_in29 = reg_0825;
    19: op1_02_in29 = reg_0002;
    20: op1_02_in29 = imem07_in[107:104];
    21: op1_02_in29 = reg_0387;
    22: op1_02_in29 = reg_0296;
    23: op1_02_in29 = imem02_in[103:100];
    24: op1_02_in29 = reg_0144;
    25: op1_02_in29 = reg_0161;
    26: op1_02_in29 = imem06_in[7:4];
    75: op1_02_in29 = imem06_in[7:4];
    28: op1_02_in29 = reg_0803;
    29: op1_02_in29 = reg_0258;
    31: op1_02_in29 = reg_0096;
    32: op1_02_in29 = reg_0547;
    33: op1_02_in29 = imem06_in[99:96];
    34: op1_02_in29 = reg_0805;
    35: op1_02_in29 = reg_0637;
    36: op1_02_in29 = reg_0396;
    37: op1_02_in29 = reg_0298;
    38: op1_02_in29 = reg_0516;
    39: op1_02_in29 = reg_0445;
    40: op1_02_in29 = imem06_in[3:0];
    41: op1_02_in29 = reg_0820;
    42: op1_02_in29 = imem03_in[107:104];
    43: op1_02_in29 = imem05_in[87:84];
    44: op1_02_in29 = reg_0438;
    45: op1_02_in29 = imem02_in[67:64];
    46: op1_02_in29 = reg_0512;
    47: op1_02_in29 = imem06_in[59:56];
    48: op1_02_in29 = imem02_in[87:84];
    49: op1_02_in29 = imem01_in[51:48];
    51: op1_02_in29 = reg_0407;
    52: op1_02_in29 = reg_0180;
    55: op1_02_in29 = reg_0574;
    56: op1_02_in29 = imem03_in[3:0];
    57: op1_02_in29 = reg_0599;
    59: op1_02_in29 = imem05_in[63:60];
    60: op1_02_in29 = reg_0800;
    61: op1_02_in29 = reg_0598;
    64: op1_02_in29 = imem01_in[111:108];
    65: op1_02_in29 = reg_0660;
    66: op1_02_in29 = reg_0219;
    67: op1_02_in29 = imem02_in[23:20];
    68: op1_02_in29 = reg_0242;
    70: op1_02_in29 = reg_0566;
    72: op1_02_in29 = reg_0497;
    73: op1_02_in29 = reg_0672;
    74: op1_02_in29 = imem03_in[47:44];
    76: op1_02_in29 = reg_0249;
    77: op1_02_in29 = reg_0175;
    78: op1_02_in29 = reg_0101;
    79: op1_02_in29 = reg_0675;
    80: op1_02_in29 = reg_0588;
    81: op1_02_in29 = imem03_in[103:100];
    82: op1_02_in29 = reg_0182;
    83: op1_02_in29 = reg_0742;
    84: op1_02_in29 = reg_0506;
    85: op1_02_in29 = reg_0808;
    88: op1_02_in29 = reg_0810;
    89: op1_02_in29 = reg_0671;
    90: op1_02_in29 = reg_0505;
    91: op1_02_in29 = imem02_in[115:112];
    92: op1_02_in29 = reg_0257;
    93: op1_02_in29 = reg_0277;
    94: op1_02_in29 = reg_0499;
    95: op1_02_in29 = reg_0491;
    96: op1_02_in29 = reg_0290;
    default: op1_02_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_02_inv29 = 1;
    6: op1_02_inv29 = 1;
    7: op1_02_inv29 = 1;
    9: op1_02_inv29 = 1;
    11: op1_02_inv29 = 1;
    12: op1_02_inv29 = 1;
    14: op1_02_inv29 = 1;
    15: op1_02_inv29 = 1;
    17: op1_02_inv29 = 1;
    18: op1_02_inv29 = 1;
    19: op1_02_inv29 = 1;
    22: op1_02_inv29 = 1;
    25: op1_02_inv29 = 1;
    26: op1_02_inv29 = 1;
    28: op1_02_inv29 = 1;
    31: op1_02_inv29 = 1;
    32: op1_02_inv29 = 1;
    34: op1_02_inv29 = 1;
    36: op1_02_inv29 = 1;
    38: op1_02_inv29 = 1;
    40: op1_02_inv29 = 1;
    43: op1_02_inv29 = 1;
    49: op1_02_inv29 = 1;
    52: op1_02_inv29 = 1;
    55: op1_02_inv29 = 1;
    57: op1_02_inv29 = 1;
    58: op1_02_inv29 = 1;
    61: op1_02_inv29 = 1;
    64: op1_02_inv29 = 1;
    72: op1_02_inv29 = 1;
    73: op1_02_inv29 = 1;
    74: op1_02_inv29 = 1;
    75: op1_02_inv29 = 1;
    77: op1_02_inv29 = 1;
    84: op1_02_inv29 = 1;
    89: op1_02_inv29 = 1;
    92: op1_02_inv29 = 1;
    93: op1_02_inv29 = 1;
    94: op1_02_inv29 = 1;
    default: op1_02_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_02_in30 = reg_0546;
    5: op1_02_in30 = reg_0219;
    6: op1_02_in30 = reg_0147;
    93: op1_02_in30 = reg_0147;
    7: op1_02_in30 = reg_0111;
    8: op1_02_in30 = imem04_in[67:64];
    9: op1_02_in30 = reg_0547;
    10: op1_02_in30 = reg_0494;
    11: op1_02_in30 = imem03_in[107:104];
    12: op1_02_in30 = imem05_in[39:36];
    13: op1_02_in30 = reg_0245;
    14: op1_02_in30 = reg_0001;
    15: op1_02_in30 = reg_0273;
    17: op1_02_in30 = reg_0807;
    28: op1_02_in30 = reg_0807;
    18: op1_02_in30 = reg_0516;
    19: op1_02_in30 = reg_0808;
    20: op1_02_in30 = reg_0720;
    21: op1_02_in30 = reg_0317;
    22: op1_02_in30 = reg_0256;
    23: op1_02_in30 = reg_0654;
    24: op1_02_in30 = reg_0791;
    25: op1_02_in30 = reg_0169;
    52: op1_02_in30 = reg_0169;
    26: op1_02_in30 = imem06_in[59:56];
    29: op1_02_in30 = reg_0255;
    31: op1_02_in30 = reg_0535;
    32: op1_02_in30 = reg_0303;
    33: op1_02_in30 = reg_0617;
    34: op1_02_in30 = reg_0004;
    88: op1_02_in30 = reg_0004;
    35: op1_02_in30 = reg_0657;
    36: op1_02_in30 = reg_0570;
    37: op1_02_in30 = reg_0278;
    38: op1_02_in30 = reg_0053;
    39: op1_02_in30 = reg_0427;
    40: op1_02_in30 = imem06_in[39:36];
    41: op1_02_in30 = reg_0227;
    42: op1_02_in30 = reg_0579;
    57: op1_02_in30 = reg_0579;
    43: op1_02_in30 = imem05_in[127:124];
    44: op1_02_in30 = reg_0167;
    45: op1_02_in30 = imem02_in[75:72];
    46: op1_02_in30 = reg_0513;
    47: op1_02_in30 = imem06_in[67:64];
    48: op1_02_in30 = imem02_in[107:104];
    49: op1_02_in30 = imem01_in[55:52];
    51: op1_02_in30 = reg_0405;
    55: op1_02_in30 = reg_0054;
    56: op1_02_in30 = imem03_in[63:60];
    58: op1_02_in30 = reg_0670;
    59: op1_02_in30 = imem05_in[71:68];
    60: op1_02_in30 = reg_0806;
    96: op1_02_in30 = reg_0806;
    61: op1_02_in30 = imem05_in[23:20];
    64: op1_02_in30 = reg_0653;
    65: op1_02_in30 = reg_0106;
    66: op1_02_in30 = reg_0124;
    67: op1_02_in30 = imem02_in[51:48];
    68: op1_02_in30 = reg_0031;
    70: op1_02_in30 = reg_0518;
    72: op1_02_in30 = reg_0102;
    73: op1_02_in30 = reg_0675;
    74: op1_02_in30 = imem03_in[59:56];
    75: op1_02_in30 = imem06_in[11:8];
    76: op1_02_in30 = reg_0307;
    77: op1_02_in30 = reg_0172;
    78: op1_02_in30 = reg_0237;
    79: op1_02_in30 = reg_0126;
    80: op1_02_in30 = reg_0331;
    81: op1_02_in30 = imem03_in[115:112];
    82: op1_02_in30 = reg_0183;
    83: op1_02_in30 = reg_0152;
    84: op1_02_in30 = reg_0123;
    85: op1_02_in30 = reg_0800;
    89: op1_02_in30 = imem02_in[15:12];
    90: op1_02_in30 = reg_0673;
    91: op1_02_in30 = reg_0704;
    92: op1_02_in30 = reg_0783;
    94: op1_02_in30 = reg_0144;
    95: op1_02_in30 = reg_0138;
    default: op1_02_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_02_inv30 = 1;
    5: op1_02_inv30 = 1;
    7: op1_02_inv30 = 1;
    8: op1_02_inv30 = 1;
    9: op1_02_inv30 = 1;
    10: op1_02_inv30 = 1;
    14: op1_02_inv30 = 1;
    17: op1_02_inv30 = 1;
    18: op1_02_inv30 = 1;
    22: op1_02_inv30 = 1;
    23: op1_02_inv30 = 1;
    26: op1_02_inv30 = 1;
    33: op1_02_inv30 = 1;
    34: op1_02_inv30 = 1;
    36: op1_02_inv30 = 1;
    40: op1_02_inv30 = 1;
    41: op1_02_inv30 = 1;
    47: op1_02_inv30 = 1;
    49: op1_02_inv30 = 1;
    52: op1_02_inv30 = 1;
    59: op1_02_inv30 = 1;
    66: op1_02_inv30 = 1;
    68: op1_02_inv30 = 1;
    70: op1_02_inv30 = 1;
    72: op1_02_inv30 = 1;
    73: op1_02_inv30 = 1;
    74: op1_02_inv30 = 1;
    76: op1_02_inv30 = 1;
    77: op1_02_inv30 = 1;
    78: op1_02_inv30 = 1;
    81: op1_02_inv30 = 1;
    83: op1_02_inv30 = 1;
    89: op1_02_inv30 = 1;
    92: op1_02_inv30 = 1;
    96: op1_02_inv30 = 1;
    default: op1_02_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_02_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_02_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in00 = reg_0547;
    5: op1_03_in00 = reg_0122;
    6: op1_03_in00 = reg_0149;
    7: op1_03_in00 = reg_0125;
    8: op1_03_in00 = imem04_in[91:88];
    9: op1_03_in00 = reg_0281;
    3: op1_03_in00 = imem07_in[27:24];
    2: op1_03_in00 = imem07_in[47:44];
    10: op1_03_in00 = reg_0780;
    43: op1_03_in00 = reg_0780;
    11: op1_03_in00 = imem03_in[127:124];
    12: op1_03_in00 = imem05_in[47:44];
    13: op1_03_in00 = reg_0249;
    14: op1_03_in00 = reg_0003;
    19: op1_03_in00 = reg_0003;
    15: op1_03_in00 = reg_0226;
    94: op1_03_in00 = reg_0226;
    16: op1_03_in00 = imem00_in[27:24];
    17: op1_03_in00 = reg_0283;
    18: op1_03_in00 = reg_0235;
    1: op1_03_in00 = imem07_in[91:88];
    20: op1_03_in00 = imem00_in[59:56];
    21: op1_03_in00 = reg_0319;
    22: op1_03_in00 = imem05_in[31:28];
    23: op1_03_in00 = reg_0647;
    24: op1_03_in00 = imem06_in[39:36];
    25: op1_03_in00 = imem00_in[3:0];
    26: op1_03_in00 = imem06_in[71:68];
    27: op1_03_in00 = imem00_in[11:8];
    30: op1_03_in00 = imem00_in[11:8];
    62: op1_03_in00 = imem00_in[11:8];
    28: op1_03_in00 = reg_0806;
    29: op1_03_in00 = reg_0077;
    31: op1_03_in00 = reg_0538;
    32: op1_03_in00 = reg_0054;
    33: op1_03_in00 = reg_0619;
    34: op1_03_in00 = imem04_in[11:8];
    35: op1_03_in00 = reg_0665;
    36: op1_03_in00 = reg_0803;
    37: op1_03_in00 = reg_0257;
    38: op1_03_in00 = reg_0290;
    39: op1_03_in00 = reg_0437;
    40: op1_03_in00 = imem06_in[51:48];
    41: op1_03_in00 = reg_0548;
    42: op1_03_in00 = reg_0585;
    44: op1_03_in00 = imem00_in[55:52];
    45: op1_03_in00 = imem02_in[79:76];
    46: op1_03_in00 = imem05_in[11:8];
    47: op1_03_in00 = imem06_in[87:84];
    48: op1_03_in00 = imem02_in[123:120];
    49: op1_03_in00 = imem01_in[63:60];
    50: op1_03_in00 = imem00_in[83:80];
    51: op1_03_in00 = reg_0776;
    52: op1_03_in00 = reg_0160;
    53: op1_03_in00 = imem00_in[15:12];
    69: op1_03_in00 = imem00_in[15:12];
    54: op1_03_in00 = imem00_in[123:120];
    63: op1_03_in00 = imem00_in[123:120];
    55: op1_03_in00 = reg_0294;
    56: op1_03_in00 = imem03_in[79:76];
    57: op1_03_in00 = reg_0596;
    58: op1_03_in00 = reg_0104;
    59: op1_03_in00 = imem05_in[79:76];
    60: op1_03_in00 = reg_0004;
    61: op1_03_in00 = imem05_in[27:24];
    64: op1_03_in00 = reg_0765;
    65: op1_03_in00 = reg_0671;
    66: op1_03_in00 = reg_0673;
    67: op1_03_in00 = imem02_in[103:100];
    68: op1_03_in00 = reg_0608;
    70: op1_03_in00 = reg_0314;
    71: op1_03_in00 = imem00_in[7:4];
    72: op1_03_in00 = reg_0101;
    73: op1_03_in00 = imem02_in[23:20];
    74: op1_03_in00 = imem03_in[83:80];
    75: op1_03_in00 = imem06_in[43:40];
    76: op1_03_in00 = reg_0790;
    77: op1_03_in00 = reg_0169;
    78: op1_03_in00 = reg_0241;
    79: op1_03_in00 = imem02_in[3:0];
    80: op1_03_in00 = reg_0755;
    81: op1_03_in00 = reg_0347;
    82: op1_03_in00 = reg_0141;
    83: op1_03_in00 = reg_0829;
    84: op1_03_in00 = reg_0677;
    85: op1_03_in00 = imem04_in[15:12];
    86: op1_03_in00 = imem00_in[35:32];
    87: op1_03_in00 = imem00_in[99:96];
    88: op1_03_in00 = imem04_in[39:36];
    89: op1_03_in00 = imem02_in[19:16];
    90: op1_03_in00 = reg_0118;
    91: op1_03_in00 = reg_0753;
    92: op1_03_in00 = reg_0155;
    93: op1_03_in00 = reg_0822;
    95: op1_03_in00 = reg_0148;
    96: op1_03_in00 = reg_0809;
    default: op1_03_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv00 = 1;
    3: op1_03_inv00 = 1;
    14: op1_03_inv00 = 1;
    15: op1_03_inv00 = 1;
    16: op1_03_inv00 = 1;
    17: op1_03_inv00 = 1;
    18: op1_03_inv00 = 1;
    1: op1_03_inv00 = 1;
    21: op1_03_inv00 = 1;
    30: op1_03_inv00 = 1;
    31: op1_03_inv00 = 1;
    34: op1_03_inv00 = 1;
    40: op1_03_inv00 = 1;
    41: op1_03_inv00 = 1;
    43: op1_03_inv00 = 1;
    46: op1_03_inv00 = 1;
    47: op1_03_inv00 = 1;
    50: op1_03_inv00 = 1;
    56: op1_03_inv00 = 1;
    57: op1_03_inv00 = 1;
    59: op1_03_inv00 = 1;
    60: op1_03_inv00 = 1;
    61: op1_03_inv00 = 1;
    62: op1_03_inv00 = 1;
    63: op1_03_inv00 = 1;
    64: op1_03_inv00 = 1;
    67: op1_03_inv00 = 1;
    68: op1_03_inv00 = 1;
    69: op1_03_inv00 = 1;
    70: op1_03_inv00 = 1;
    72: op1_03_inv00 = 1;
    76: op1_03_inv00 = 1;
    78: op1_03_inv00 = 1;
    79: op1_03_inv00 = 1;
    81: op1_03_inv00 = 1;
    85: op1_03_inv00 = 1;
    87: op1_03_inv00 = 1;
    88: op1_03_inv00 = 1;
    91: op1_03_inv00 = 1;
    92: op1_03_inv00 = 1;
    93: op1_03_inv00 = 1;
    95: op1_03_inv00 = 1;
    default: op1_03_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in01 = reg_0301;
    5: op1_03_in01 = reg_0114;
    6: op1_03_in01 = reg_0134;
    7: op1_03_in01 = reg_0116;
    8: op1_03_in01 = imem04_in[107:104];
    9: op1_03_in01 = reg_0283;
    3: op1_03_in01 = imem07_in[51:48];
    2: op1_03_in01 = imem07_in[63:60];
    10: op1_03_in01 = reg_0271;
    11: op1_03_in01 = reg_0596;
    12: op1_03_in01 = imem05_in[71:68];
    13: op1_03_in01 = reg_0127;
    14: op1_03_in01 = reg_0802;
    15: op1_03_in01 = reg_0133;
    16: op1_03_in01 = imem00_in[115:112];
    62: op1_03_in01 = imem00_in[115:112];
    17: op1_03_in01 = reg_0055;
    18: op1_03_in01 = reg_0236;
    19: op1_03_in01 = reg_0807;
    20: op1_03_in01 = imem00_in[119:116];
    21: op1_03_in01 = reg_0377;
    22: op1_03_in01 = imem05_in[35:32];
    61: op1_03_in01 = imem05_in[35:32];
    23: op1_03_in01 = reg_0334;
    24: op1_03_in01 = reg_0625;
    25: op1_03_in01 = imem00_in[19:16];
    69: op1_03_in01 = imem00_in[19:16];
    71: op1_03_in01 = imem00_in[19:16];
    26: op1_03_in01 = imem06_in[75:72];
    40: op1_03_in01 = imem06_in[75:72];
    27: op1_03_in01 = imem00_in[43:40];
    28: op1_03_in01 = reg_0809;
    29: op1_03_in01 = reg_0064;
    30: op1_03_in01 = imem00_in[35:32];
    31: op1_03_in01 = imem03_in[19:16];
    32: op1_03_in01 = reg_0305;
    33: op1_03_in01 = reg_0618;
    34: op1_03_in01 = imem04_in[15:12];
    35: op1_03_in01 = reg_0094;
    36: op1_03_in01 = imem04_in[55:52];
    37: op1_03_in01 = reg_0289;
    38: op1_03_in01 = reg_0267;
    39: op1_03_in01 = reg_0435;
    41: op1_03_in01 = reg_0559;
    42: op1_03_in01 = reg_0578;
    43: op1_03_in01 = reg_0785;
    44: op1_03_in01 = imem00_in[59:56];
    45: op1_03_in01 = imem02_in[107:104];
    67: op1_03_in01 = imem02_in[107:104];
    46: op1_03_in01 = imem05_in[27:24];
    47: op1_03_in01 = imem06_in[115:112];
    48: op1_03_in01 = reg_0664;
    49: op1_03_in01 = imem01_in[75:72];
    50: op1_03_in01 = imem00_in[91:88];
    51: op1_03_in01 = reg_0038;
    52: op1_03_in01 = reg_0166;
    77: op1_03_in01 = reg_0166;
    53: op1_03_in01 = imem00_in[63:60];
    54: op1_03_in01 = reg_0472;
    55: op1_03_in01 = reg_0243;
    56: op1_03_in01 = reg_0319;
    57: op1_03_in01 = reg_0329;
    58: op1_03_in01 = reg_0592;
    59: op1_03_in01 = imem05_in[107:104];
    60: op1_03_in01 = imem04_in[19:16];
    63: op1_03_in01 = reg_0612;
    64: op1_03_in01 = reg_0322;
    65: op1_03_in01 = reg_0107;
    66: op1_03_in01 = reg_0073;
    68: op1_03_in01 = reg_0549;
    70: op1_03_in01 = reg_0095;
    72: op1_03_in01 = reg_0130;
    73: op1_03_in01 = imem02_in[47:44];
    74: op1_03_in01 = reg_0579;
    75: op1_03_in01 = imem06_in[83:80];
    76: op1_03_in01 = reg_0822;
    78: op1_03_in01 = reg_0220;
    79: op1_03_in01 = imem02_in[119:116];
    80: op1_03_in01 = reg_0483;
    81: op1_03_in01 = reg_0604;
    82: op1_03_in01 = reg_0091;
    83: op1_03_in01 = reg_0796;
    84: op1_03_in01 = reg_0675;
    85: op1_03_in01 = imem04_in[51:48];
    86: op1_03_in01 = imem00_in[39:36];
    87: op1_03_in01 = reg_0685;
    88: op1_03_in01 = imem04_in[59:56];
    89: op1_03_in01 = imem02_in[91:88];
    90: op1_03_in01 = reg_0125;
    91: op1_03_in01 = reg_0274;
    92: op1_03_in01 = reg_0824;
    93: op1_03_in01 = reg_0156;
    94: op1_03_in01 = reg_0583;
    95: op1_03_in01 = reg_0827;
    96: op1_03_in01 = reg_0004;
    default: op1_03_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv01 = 1;
    5: op1_03_inv01 = 1;
    7: op1_03_inv01 = 1;
    9: op1_03_inv01 = 1;
    10: op1_03_inv01 = 1;
    11: op1_03_inv01 = 1;
    12: op1_03_inv01 = 1;
    13: op1_03_inv01 = 1;
    16: op1_03_inv01 = 1;
    18: op1_03_inv01 = 1;
    19: op1_03_inv01 = 1;
    20: op1_03_inv01 = 1;
    22: op1_03_inv01 = 1;
    23: op1_03_inv01 = 1;
    24: op1_03_inv01 = 1;
    25: op1_03_inv01 = 1;
    26: op1_03_inv01 = 1;
    27: op1_03_inv01 = 1;
    31: op1_03_inv01 = 1;
    33: op1_03_inv01 = 1;
    34: op1_03_inv01 = 1;
    38: op1_03_inv01 = 1;
    40: op1_03_inv01 = 1;
    43: op1_03_inv01 = 1;
    45: op1_03_inv01 = 1;
    50: op1_03_inv01 = 1;
    52: op1_03_inv01 = 1;
    54: op1_03_inv01 = 1;
    56: op1_03_inv01 = 1;
    57: op1_03_inv01 = 1;
    58: op1_03_inv01 = 1;
    59: op1_03_inv01 = 1;
    60: op1_03_inv01 = 1;
    64: op1_03_inv01 = 1;
    65: op1_03_inv01 = 1;
    66: op1_03_inv01 = 1;
    68: op1_03_inv01 = 1;
    71: op1_03_inv01 = 1;
    72: op1_03_inv01 = 1;
    73: op1_03_inv01 = 1;
    75: op1_03_inv01 = 1;
    80: op1_03_inv01 = 1;
    83: op1_03_inv01 = 1;
    84: op1_03_inv01 = 1;
    90: op1_03_inv01 = 1;
    92: op1_03_inv01 = 1;
    95: op1_03_inv01 = 1;
    default: op1_03_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in02 = reg_0302;
    5: op1_03_in02 = reg_0113;
    6: op1_03_in02 = imem06_in[27:24];
    7: op1_03_in02 = reg_0117;
    8: op1_03_in02 = imem04_in[111:108];
    9: op1_03_in02 = reg_0282;
    3: op1_03_in02 = imem07_in[79:76];
    2: op1_03_in02 = imem07_in[79:76];
    10: op1_03_in02 = reg_0273;
    11: op1_03_in02 = reg_0578;
    12: op1_03_in02 = reg_0786;
    13: op1_03_in02 = reg_0110;
    14: op1_03_in02 = reg_0810;
    15: op1_03_in02 = reg_0151;
    16: op1_03_in02 = reg_0693;
    17: op1_03_in02 = reg_0285;
    18: op1_03_in02 = reg_0245;
    19: op1_03_in02 = reg_0802;
    20: op1_03_in02 = reg_0672;
    66: op1_03_in02 = reg_0672;
    21: op1_03_in02 = reg_0397;
    72: op1_03_in02 = reg_0397;
    22: op1_03_in02 = imem05_in[51:48];
    23: op1_03_in02 = reg_0333;
    24: op1_03_in02 = reg_0613;
    25: op1_03_in02 = imem00_in[35:32];
    26: op1_03_in02 = imem06_in[95:92];
    40: op1_03_in02 = imem06_in[95:92];
    27: op1_03_in02 = imem00_in[127:124];
    28: op1_03_in02 = imem04_in[55:52];
    29: op1_03_in02 = imem05_in[67:64];
    30: op1_03_in02 = imem00_in[71:68];
    31: op1_03_in02 = imem03_in[43:40];
    35: op1_03_in02 = imem03_in[43:40];
    32: op1_03_in02 = reg_0294;
    33: op1_03_in02 = reg_0632;
    34: op1_03_in02 = imem04_in[19:16];
    36: op1_03_in02 = imem04_in[87:84];
    37: op1_03_in02 = reg_0254;
    38: op1_03_in02 = reg_0065;
    39: op1_03_in02 = reg_0179;
    41: op1_03_in02 = reg_0241;
    42: op1_03_in02 = reg_0384;
    43: op1_03_in02 = reg_0783;
    83: op1_03_in02 = reg_0783;
    93: op1_03_in02 = reg_0783;
    44: op1_03_in02 = imem00_in[63:60];
    45: op1_03_in02 = reg_0664;
    46: op1_03_in02 = imem05_in[71:68];
    47: op1_03_in02 = reg_0630;
    48: op1_03_in02 = reg_0301;
    49: op1_03_in02 = imem01_in[83:80];
    50: op1_03_in02 = imem00_in[95:92];
    69: op1_03_in02 = imem00_in[95:92];
    51: op1_03_in02 = reg_0028;
    52: op1_03_in02 = reg_0177;
    53: op1_03_in02 = imem00_in[67:64];
    54: op1_03_in02 = imem01_in[19:16];
    55: op1_03_in02 = reg_0592;
    56: op1_03_in02 = reg_0350;
    57: op1_03_in02 = reg_0751;
    58: op1_03_in02 = reg_0120;
    59: op1_03_in02 = reg_0781;
    60: op1_03_in02 = imem04_in[35:32];
    61: op1_03_in02 = imem05_in[75:72];
    62: op1_03_in02 = reg_0697;
    63: op1_03_in02 = reg_0463;
    64: op1_03_in02 = reg_0232;
    65: op1_03_in02 = reg_0678;
    67: op1_03_in02 = reg_0639;
    68: op1_03_in02 = imem07_in[63:60];
    70: op1_03_in02 = reg_0097;
    71: op1_03_in02 = imem00_in[75:72];
    73: op1_03_in02 = imem02_in[51:48];
    74: op1_03_in02 = reg_0319;
    75: op1_03_in02 = imem06_in[99:96];
    76: op1_03_in02 = reg_0150;
    95: op1_03_in02 = reg_0150;
    77: op1_03_in02 = reg_0173;
    78: op1_03_in02 = reg_0504;
    79: op1_03_in02 = reg_0141;
    80: op1_03_in02 = reg_0562;
    81: op1_03_in02 = reg_0596;
    82: op1_03_in02 = reg_0176;
    84: op1_03_in02 = reg_0107;
    85: op1_03_in02 = imem04_in[99:96];
    86: op1_03_in02 = imem00_in[47:44];
    87: op1_03_in02 = reg_0686;
    88: op1_03_in02 = imem04_in[127:124];
    89: op1_03_in02 = imem02_in[127:124];
    90: op1_03_in02 = reg_0126;
    91: op1_03_in02 = reg_0059;
    92: op1_03_in02 = imem06_in[59:56];
    94: op1_03_in02 = reg_0491;
    96: op1_03_in02 = imem04_in[23:20];
    default: op1_03_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_03_inv02 = 1;
    8: op1_03_inv02 = 1;
    9: op1_03_inv02 = 1;
    3: op1_03_inv02 = 1;
    11: op1_03_inv02 = 1;
    13: op1_03_inv02 = 1;
    18: op1_03_inv02 = 1;
    19: op1_03_inv02 = 1;
    21: op1_03_inv02 = 1;
    23: op1_03_inv02 = 1;
    24: op1_03_inv02 = 1;
    29: op1_03_inv02 = 1;
    30: op1_03_inv02 = 1;
    33: op1_03_inv02 = 1;
    35: op1_03_inv02 = 1;
    39: op1_03_inv02 = 1;
    43: op1_03_inv02 = 1;
    49: op1_03_inv02 = 1;
    50: op1_03_inv02 = 1;
    51: op1_03_inv02 = 1;
    52: op1_03_inv02 = 1;
    53: op1_03_inv02 = 1;
    54: op1_03_inv02 = 1;
    55: op1_03_inv02 = 1;
    59: op1_03_inv02 = 1;
    61: op1_03_inv02 = 1;
    62: op1_03_inv02 = 1;
    64: op1_03_inv02 = 1;
    66: op1_03_inv02 = 1;
    68: op1_03_inv02 = 1;
    70: op1_03_inv02 = 1;
    71: op1_03_inv02 = 1;
    72: op1_03_inv02 = 1;
    74: op1_03_inv02 = 1;
    76: op1_03_inv02 = 1;
    77: op1_03_inv02 = 1;
    78: op1_03_inv02 = 1;
    79: op1_03_inv02 = 1;
    81: op1_03_inv02 = 1;
    82: op1_03_inv02 = 1;
    83: op1_03_inv02 = 1;
    86: op1_03_inv02 = 1;
    88: op1_03_inv02 = 1;
    91: op1_03_inv02 = 1;
    92: op1_03_inv02 = 1;
    93: op1_03_inv02 = 1;
    95: op1_03_inv02 = 1;
    default: op1_03_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in03 = reg_0276;
    5: op1_03_in03 = imem02_in[7:4];
    65: op1_03_in03 = imem02_in[7:4];
    6: op1_03_in03 = imem06_in[43:40];
    7: op1_03_in03 = imem02_in[27:24];
    8: op1_03_in03 = imem04_in[115:112];
    9: op1_03_in03 = reg_0293;
    3: op1_03_in03 = imem07_in[87:84];
    2: op1_03_in03 = imem07_in[107:104];
    10: op1_03_in03 = reg_0260;
    11: op1_03_in03 = reg_0384;
    12: op1_03_in03 = reg_0498;
    13: op1_03_in03 = imem02_in[11:8];
    14: op1_03_in03 = imem04_in[67:64];
    15: op1_03_in03 = reg_0128;
    16: op1_03_in03 = reg_0683;
    62: op1_03_in03 = reg_0683;
    17: op1_03_in03 = reg_0050;
    18: op1_03_in03 = reg_0111;
    19: op1_03_in03 = reg_0810;
    20: op1_03_in03 = reg_0684;
    21: op1_03_in03 = reg_0361;
    22: op1_03_in03 = imem05_in[55:52];
    23: op1_03_in03 = reg_0345;
    24: op1_03_in03 = reg_0609;
    25: op1_03_in03 = imem00_in[39:36];
    26: op1_03_in03 = reg_0610;
    27: op1_03_in03 = reg_0690;
    28: op1_03_in03 = imem04_in[63:60];
    34: op1_03_in03 = imem04_in[63:60];
    29: op1_03_in03 = imem05_in[91:88];
    30: op1_03_in03 = imem00_in[75:72];
    31: op1_03_in03 = imem03_in[51:48];
    35: op1_03_in03 = imem03_in[51:48];
    32: op1_03_in03 = reg_0274;
    33: op1_03_in03 = reg_0762;
    36: op1_03_in03 = reg_0556;
    37: op1_03_in03 = reg_0069;
    38: op1_03_in03 = reg_0255;
    39: op1_03_in03 = reg_0163;
    40: op1_03_in03 = imem06_in[127:124];
    41: op1_03_in03 = reg_0418;
    42: op1_03_in03 = reg_0755;
    43: op1_03_in03 = reg_0790;
    44: op1_03_in03 = imem00_in[91:88];
    45: op1_03_in03 = reg_0661;
    46: op1_03_in03 = reg_0792;
    47: op1_03_in03 = reg_0218;
    48: op1_03_in03 = reg_0641;
    49: op1_03_in03 = reg_0563;
    50: op1_03_in03 = imem00_in[127:124];
    51: op1_03_in03 = reg_0607;
    52: op1_03_in03 = reg_0168;
    53: op1_03_in03 = imem00_in[111:108];
    54: op1_03_in03 = imem01_in[23:20];
    55: op1_03_in03 = reg_0660;
    56: op1_03_in03 = reg_0281;
    57: op1_03_in03 = reg_0571;
    58: op1_03_in03 = reg_0108;
    66: op1_03_in03 = reg_0108;
    59: op1_03_in03 = reg_0495;
    60: op1_03_in03 = imem04_in[51:48];
    61: op1_03_in03 = imem05_in[111:108];
    63: op1_03_in03 = reg_0465;
    64: op1_03_in03 = reg_0423;
    67: op1_03_in03 = reg_0753;
    68: op1_03_in03 = imem07_in[111:108];
    69: op1_03_in03 = imem00_in[123:120];
    70: op1_03_in03 = reg_0531;
    71: op1_03_in03 = imem00_in[79:76];
    86: op1_03_in03 = imem00_in[79:76];
    72: op1_03_in03 = reg_0235;
    73: op1_03_in03 = imem02_in[79:76];
    74: op1_03_in03 = reg_0600;
    75: op1_03_in03 = imem06_in[123:120];
    76: op1_03_in03 = reg_0152;
    78: op1_03_in03 = reg_0424;
    79: op1_03_in03 = reg_0548;
    80: op1_03_in03 = reg_0019;
    81: op1_03_in03 = reg_0591;
    82: op1_03_in03 = reg_0279;
    83: op1_03_in03 = reg_0765;
    93: op1_03_in03 = reg_0765;
    84: op1_03_in03 = reg_0676;
    85: op1_03_in03 = imem04_in[103:100];
    87: op1_03_in03 = reg_0680;
    88: op1_03_in03 = reg_0544;
    89: op1_03_in03 = reg_0057;
    90: op1_03_in03 = imem02_in[99:96];
    91: op1_03_in03 = reg_0320;
    92: op1_03_in03 = imem06_in[83:80];
    94: op1_03_in03 = reg_0579;
    95: op1_03_in03 = reg_0143;
    96: op1_03_in03 = imem04_in[31:28];
    default: op1_03_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv03 = 1;
    5: op1_03_inv03 = 1;
    9: op1_03_inv03 = 1;
    2: op1_03_inv03 = 1;
    12: op1_03_inv03 = 1;
    14: op1_03_inv03 = 1;
    16: op1_03_inv03 = 1;
    18: op1_03_inv03 = 1;
    19: op1_03_inv03 = 1;
    21: op1_03_inv03 = 1;
    22: op1_03_inv03 = 1;
    26: op1_03_inv03 = 1;
    28: op1_03_inv03 = 1;
    29: op1_03_inv03 = 1;
    30: op1_03_inv03 = 1;
    32: op1_03_inv03 = 1;
    33: op1_03_inv03 = 1;
    34: op1_03_inv03 = 1;
    35: op1_03_inv03 = 1;
    38: op1_03_inv03 = 1;
    39: op1_03_inv03 = 1;
    43: op1_03_inv03 = 1;
    44: op1_03_inv03 = 1;
    45: op1_03_inv03 = 1;
    46: op1_03_inv03 = 1;
    47: op1_03_inv03 = 1;
    49: op1_03_inv03 = 1;
    50: op1_03_inv03 = 1;
    52: op1_03_inv03 = 1;
    53: op1_03_inv03 = 1;
    55: op1_03_inv03 = 1;
    56: op1_03_inv03 = 1;
    58: op1_03_inv03 = 1;
    59: op1_03_inv03 = 1;
    60: op1_03_inv03 = 1;
    61: op1_03_inv03 = 1;
    62: op1_03_inv03 = 1;
    64: op1_03_inv03 = 1;
    66: op1_03_inv03 = 1;
    67: op1_03_inv03 = 1;
    70: op1_03_inv03 = 1;
    71: op1_03_inv03 = 1;
    73: op1_03_inv03 = 1;
    76: op1_03_inv03 = 1;
    78: op1_03_inv03 = 1;
    80: op1_03_inv03 = 1;
    82: op1_03_inv03 = 1;
    83: op1_03_inv03 = 1;
    85: op1_03_inv03 = 1;
    86: op1_03_inv03 = 1;
    89: op1_03_inv03 = 1;
    90: op1_03_inv03 = 1;
    93: op1_03_inv03 = 1;
    96: op1_03_inv03 = 1;
    default: op1_03_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in04 = reg_0288;
    5: op1_03_in04 = reg_0653;
    6: op1_03_in04 = imem06_in[79:76];
    7: op1_03_in04 = imem02_in[51:48];
    8: op1_03_in04 = reg_0550;
    9: op1_03_in04 = reg_0285;
    3: op1_03_in04 = imem07_in[95:92];
    2: op1_03_in04 = imem07_in[111:108];
    10: op1_03_in04 = reg_0272;
    11: op1_03_in04 = reg_0388;
    42: op1_03_in04 = reg_0388;
    12: op1_03_in04 = reg_0735;
    13: op1_03_in04 = imem02_in[27:24];
    65: op1_03_in04 = imem02_in[27:24];
    14: op1_03_in04 = imem04_in[83:80];
    15: op1_03_in04 = reg_0129;
    16: op1_03_in04 = reg_0672;
    17: op1_03_in04 = reg_0542;
    18: op1_03_in04 = reg_0119;
    19: op1_03_in04 = reg_0004;
    20: op1_03_in04 = reg_0481;
    21: op1_03_in04 = reg_0331;
    22: op1_03_in04 = imem05_in[67:64];
    23: op1_03_in04 = reg_0355;
    48: op1_03_in04 = reg_0355;
    24: op1_03_in04 = reg_0618;
    25: op1_03_in04 = imem00_in[47:44];
    26: op1_03_in04 = reg_0631;
    27: op1_03_in04 = reg_0678;
    28: op1_03_in04 = imem04_in[79:76];
    34: op1_03_in04 = imem04_in[79:76];
    29: op1_03_in04 = imem05_in[95:92];
    30: op1_03_in04 = imem00_in[107:104];
    31: op1_03_in04 = imem03_in[59:56];
    35: op1_03_in04 = imem03_in[59:56];
    32: op1_03_in04 = reg_0291;
    33: op1_03_in04 = reg_0405;
    36: op1_03_in04 = reg_0054;
    37: op1_03_in04 = reg_0256;
    38: op1_03_in04 = imem05_in[15:12];
    39: op1_03_in04 = reg_0166;
    40: op1_03_in04 = reg_0625;
    41: op1_03_in04 = reg_0240;
    43: op1_03_in04 = reg_0784;
    44: op1_03_in04 = imem00_in[103:100];
    45: op1_03_in04 = reg_0656;
    46: op1_03_in04 = reg_0494;
    47: op1_03_in04 = reg_0020;
    49: op1_03_in04 = reg_0734;
    50: op1_03_in04 = reg_0682;
    69: op1_03_in04 = reg_0682;
    51: op1_03_in04 = reg_0620;
    52: op1_03_in04 = reg_0158;
    53: op1_03_in04 = imem00_in[123:120];
    54: op1_03_in04 = imem01_in[59:56];
    55: op1_03_in04 = reg_0106;
    66: op1_03_in04 = reg_0106;
    56: op1_03_in04 = reg_0595;
    57: op1_03_in04 = reg_0389;
    58: op1_03_in04 = reg_0669;
    59: op1_03_in04 = reg_0091;
    60: op1_03_in04 = imem04_in[67:64];
    61: op1_03_in04 = imem05_in[127:124];
    62: op1_03_in04 = reg_0689;
    63: op1_03_in04 = reg_0455;
    64: op1_03_in04 = reg_0511;
    72: op1_03_in04 = reg_0511;
    67: op1_03_in04 = reg_0417;
    68: op1_03_in04 = imem07_in[119:116];
    70: op1_03_in04 = reg_0532;
    71: op1_03_in04 = reg_0683;
    73: op1_03_in04 = imem02_in[87:84];
    74: op1_03_in04 = reg_0571;
    75: op1_03_in04 = reg_0624;
    76: op1_03_in04 = reg_0824;
    78: op1_03_in04 = reg_0673;
    79: op1_03_in04 = reg_0702;
    80: op1_03_in04 = reg_0800;
    81: op1_03_in04 = reg_0751;
    82: op1_03_in04 = reg_0184;
    83: op1_03_in04 = imem06_in[15:12];
    84: op1_03_in04 = reg_0518;
    85: op1_03_in04 = reg_0262;
    86: op1_03_in04 = imem00_in[83:80];
    87: op1_03_in04 = reg_0469;
    88: op1_03_in04 = reg_0058;
    89: op1_03_in04 = reg_0088;
    90: op1_03_in04 = reg_0264;
    91: op1_03_in04 = reg_0594;
    92: op1_03_in04 = imem06_in[91:88];
    93: op1_03_in04 = reg_0155;
    94: op1_03_in04 = reg_0147;
    95: op1_03_in04 = imem06_in[11:8];
    96: op1_03_in04 = imem04_in[71:68];
    default: op1_03_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv04 = 1;
    9: op1_03_inv04 = 1;
    3: op1_03_inv04 = 1;
    2: op1_03_inv04 = 1;
    10: op1_03_inv04 = 1;
    13: op1_03_inv04 = 1;
    15: op1_03_inv04 = 1;
    21: op1_03_inv04 = 1;
    24: op1_03_inv04 = 1;
    25: op1_03_inv04 = 1;
    26: op1_03_inv04 = 1;
    28: op1_03_inv04 = 1;
    30: op1_03_inv04 = 1;
    31: op1_03_inv04 = 1;
    32: op1_03_inv04 = 1;
    33: op1_03_inv04 = 1;
    35: op1_03_inv04 = 1;
    36: op1_03_inv04 = 1;
    38: op1_03_inv04 = 1;
    39: op1_03_inv04 = 1;
    42: op1_03_inv04 = 1;
    44: op1_03_inv04 = 1;
    45: op1_03_inv04 = 1;
    48: op1_03_inv04 = 1;
    50: op1_03_inv04 = 1;
    51: op1_03_inv04 = 1;
    52: op1_03_inv04 = 1;
    55: op1_03_inv04 = 1;
    58: op1_03_inv04 = 1;
    60: op1_03_inv04 = 1;
    61: op1_03_inv04 = 1;
    65: op1_03_inv04 = 1;
    66: op1_03_inv04 = 1;
    69: op1_03_inv04 = 1;
    71: op1_03_inv04 = 1;
    72: op1_03_inv04 = 1;
    76: op1_03_inv04 = 1;
    78: op1_03_inv04 = 1;
    79: op1_03_inv04 = 1;
    85: op1_03_inv04 = 1;
    87: op1_03_inv04 = 1;
    88: op1_03_inv04 = 1;
    89: op1_03_inv04 = 1;
    91: op1_03_inv04 = 1;
    92: op1_03_inv04 = 1;
    95: op1_03_inv04 = 1;
    96: op1_03_inv04 = 1;
    default: op1_03_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in05 = reg_0061;
    5: op1_03_in05 = reg_0638;
    6: op1_03_in05 = imem06_in[103:100];
    7: op1_03_in05 = imem02_in[55:52];
    8: op1_03_in05 = reg_0555;
    9: op1_03_in05 = reg_0292;
    3: op1_03_in05 = imem07_in[103:100];
    2: op1_03_in05 = imem07_in[115:112];
    10: op1_03_in05 = reg_0261;
    11: op1_03_in05 = reg_0393;
    12: op1_03_in05 = reg_0526;
    13: op1_03_in05 = imem02_in[47:44];
    14: op1_03_in05 = imem04_in[91:88];
    15: op1_03_in05 = reg_0153;
    16: op1_03_in05 = reg_0676;
    58: op1_03_in05 = reg_0676;
    17: op1_03_in05 = reg_0534;
    18: op1_03_in05 = reg_0120;
    19: op1_03_in05 = imem04_in[11:8];
    20: op1_03_in05 = reg_0470;
    21: op1_03_in05 = reg_0013;
    22: op1_03_in05 = imem05_in[95:92];
    23: op1_03_in05 = reg_0335;
    24: op1_03_in05 = reg_0402;
    25: op1_03_in05 = imem00_in[75:72];
    26: op1_03_in05 = reg_0577;
    27: op1_03_in05 = reg_0688;
    28: op1_03_in05 = reg_0043;
    29: op1_03_in05 = imem05_in[115:112];
    30: op1_03_in05 = reg_0678;
    31: op1_03_in05 = imem03_in[99:96];
    32: op1_03_in05 = reg_0051;
    33: op1_03_in05 = reg_0319;
    34: op1_03_in05 = reg_0262;
    35: op1_03_in05 = imem03_in[63:60];
    36: op1_03_in05 = reg_0280;
    37: op1_03_in05 = imem05_in[7:4];
    38: op1_03_in05 = imem05_in[31:28];
    39: op1_03_in05 = reg_0164;
    40: op1_03_in05 = reg_0331;
    41: op1_03_in05 = reg_0290;
    42: op1_03_in05 = reg_0383;
    43: op1_03_in05 = reg_0787;
    46: op1_03_in05 = reg_0787;
    44: op1_03_in05 = imem00_in[107:104];
    45: op1_03_in05 = reg_0662;
    47: op1_03_in05 = reg_0606;
    48: op1_03_in05 = reg_0659;
    49: op1_03_in05 = reg_0652;
    50: op1_03_in05 = reg_0693;
    86: op1_03_in05 = reg_0693;
    51: op1_03_in05 = reg_0040;
    53: op1_03_in05 = reg_0696;
    54: op1_03_in05 = imem01_in[95:92];
    55: op1_03_in05 = reg_0669;
    78: op1_03_in05 = reg_0669;
    56: op1_03_in05 = reg_0588;
    57: op1_03_in05 = reg_0003;
    59: op1_03_in05 = reg_0246;
    60: op1_03_in05 = imem04_in[103:100];
    61: op1_03_in05 = reg_0337;
    62: op1_03_in05 = reg_0494;
    63: op1_03_in05 = reg_0466;
    64: op1_03_in05 = reg_0502;
    65: op1_03_in05 = imem02_in[43:40];
    66: op1_03_in05 = reg_0601;
    67: op1_03_in05 = reg_0114;
    68: op1_03_in05 = reg_0720;
    69: op1_03_in05 = reg_0697;
    70: op1_03_in05 = imem03_in[47:44];
    71: op1_03_in05 = reg_0117;
    72: op1_03_in05 = reg_0422;
    73: op1_03_in05 = imem02_in[99:96];
    74: op1_03_in05 = reg_0568;
    81: op1_03_in05 = reg_0568;
    75: op1_03_in05 = reg_0409;
    76: op1_03_in05 = imem06_in[11:8];
    79: op1_03_in05 = reg_0587;
    80: op1_03_in05 = reg_0008;
    83: op1_03_in05 = imem06_in[31:28];
    84: op1_03_in05 = reg_0655;
    85: op1_03_in05 = reg_0553;
    87: op1_03_in05 = reg_0460;
    88: op1_03_in05 = reg_0516;
    89: op1_03_in05 = reg_0081;
    90: op1_03_in05 = reg_0086;
    91: op1_03_in05 = reg_0365;
    92: op1_03_in05 = imem06_in[99:96];
    93: op1_03_in05 = reg_0824;
    94: op1_03_in05 = reg_0828;
    95: op1_03_in05 = imem06_in[51:48];
    96: op1_03_in05 = imem04_in[119:116];
    default: op1_03_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv05 = 1;
    5: op1_03_inv05 = 1;
    7: op1_03_inv05 = 1;
    8: op1_03_inv05 = 1;
    9: op1_03_inv05 = 1;
    10: op1_03_inv05 = 1;
    11: op1_03_inv05 = 1;
    12: op1_03_inv05 = 1;
    14: op1_03_inv05 = 1;
    15: op1_03_inv05 = 1;
    20: op1_03_inv05 = 1;
    24: op1_03_inv05 = 1;
    26: op1_03_inv05 = 1;
    28: op1_03_inv05 = 1;
    30: op1_03_inv05 = 1;
    31: op1_03_inv05 = 1;
    32: op1_03_inv05 = 1;
    34: op1_03_inv05 = 1;
    35: op1_03_inv05 = 1;
    36: op1_03_inv05 = 1;
    37: op1_03_inv05 = 1;
    39: op1_03_inv05 = 1;
    41: op1_03_inv05 = 1;
    44: op1_03_inv05 = 1;
    45: op1_03_inv05 = 1;
    46: op1_03_inv05 = 1;
    48: op1_03_inv05 = 1;
    49: op1_03_inv05 = 1;
    50: op1_03_inv05 = 1;
    51: op1_03_inv05 = 1;
    56: op1_03_inv05 = 1;
    59: op1_03_inv05 = 1;
    60: op1_03_inv05 = 1;
    61: op1_03_inv05 = 1;
    62: op1_03_inv05 = 1;
    63: op1_03_inv05 = 1;
    64: op1_03_inv05 = 1;
    66: op1_03_inv05 = 1;
    67: op1_03_inv05 = 1;
    68: op1_03_inv05 = 1;
    70: op1_03_inv05 = 1;
    71: op1_03_inv05 = 1;
    73: op1_03_inv05 = 1;
    74: op1_03_inv05 = 1;
    76: op1_03_inv05 = 1;
    78: op1_03_inv05 = 1;
    79: op1_03_inv05 = 1;
    80: op1_03_inv05 = 1;
    81: op1_03_inv05 = 1;
    84: op1_03_inv05 = 1;
    85: op1_03_inv05 = 1;
    88: op1_03_inv05 = 1;
    89: op1_03_inv05 = 1;
    90: op1_03_inv05 = 1;
    92: op1_03_inv05 = 1;
    94: op1_03_inv05 = 1;
    95: op1_03_inv05 = 1;
    96: op1_03_inv05 = 1;
    default: op1_03_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in06 = reg_0062;
    5: op1_03_in06 = reg_0643;
    6: op1_03_in06 = reg_0629;
    7: op1_03_in06 = imem02_in[111:108];
    8: op1_03_in06 = reg_0546;
    9: op1_03_in06 = reg_0286;
    3: op1_03_in06 = imem07_in[111:108];
    2: op1_03_in06 = reg_0174;
    10: op1_03_in06 = reg_0263;
    11: op1_03_in06 = reg_0007;
    12: op1_03_in06 = reg_0148;
    13: op1_03_in06 = imem02_in[71:68];
    14: op1_03_in06 = reg_0543;
    15: op1_03_in06 = reg_0140;
    16: op1_03_in06 = reg_0671;
    78: op1_03_in06 = reg_0671;
    17: op1_03_in06 = reg_0304;
    18: op1_03_in06 = reg_0101;
    19: op1_03_in06 = imem04_in[23:20];
    20: op1_03_in06 = reg_0474;
    21: op1_03_in06 = reg_0805;
    22: op1_03_in06 = imem05_in[115:112];
    23: op1_03_in06 = reg_0743;
    24: op1_03_in06 = reg_0344;
    25: op1_03_in06 = imem00_in[127:124];
    26: op1_03_in06 = reg_0627;
    27: op1_03_in06 = reg_0699;
    28: op1_03_in06 = reg_0088;
    29: op1_03_in06 = reg_0789;
    30: op1_03_in06 = reg_0463;
    31: op1_03_in06 = imem03_in[119:116];
    32: op1_03_in06 = reg_0070;
    33: op1_03_in06 = reg_0381;
    34: op1_03_in06 = reg_0087;
    35: op1_03_in06 = imem03_in[67:64];
    36: op1_03_in06 = reg_0265;
    37: op1_03_in06 = imem05_in[19:16];
    38: op1_03_in06 = reg_0488;
    39: op1_03_in06 = reg_0176;
    40: op1_03_in06 = reg_0370;
    41: op1_03_in06 = reg_0425;
    64: op1_03_in06 = reg_0425;
    42: op1_03_in06 = reg_0389;
    43: op1_03_in06 = reg_0091;
    46: op1_03_in06 = reg_0091;
    44: op1_03_in06 = reg_0695;
    45: op1_03_in06 = reg_0659;
    47: op1_03_in06 = reg_0577;
    48: op1_03_in06 = reg_0349;
    49: op1_03_in06 = reg_0217;
    50: op1_03_in06 = reg_0676;
    51: op1_03_in06 = reg_0368;
    81: op1_03_in06 = reg_0368;
    53: op1_03_in06 = reg_0691;
    54: op1_03_in06 = imem01_in[99:96];
    55: op1_03_in06 = reg_0674;
    56: op1_03_in06 = reg_0391;
    57: op1_03_in06 = reg_0803;
    58: op1_03_in06 = imem02_in[43:40];
    59: op1_03_in06 = reg_0309;
    60: op1_03_in06 = reg_0545;
    61: op1_03_in06 = reg_0113;
    62: op1_03_in06 = reg_0680;
    63: op1_03_in06 = reg_0456;
    65: op1_03_in06 = imem02_in[87:84];
    66: op1_03_in06 = reg_0121;
    67: op1_03_in06 = reg_0372;
    68: op1_03_in06 = reg_0708;
    69: op1_03_in06 = reg_0694;
    70: op1_03_in06 = imem03_in[51:48];
    71: op1_03_in06 = reg_0494;
    72: op1_03_in06 = reg_0502;
    73: op1_03_in06 = reg_0534;
    74: op1_03_in06 = reg_0403;
    75: op1_03_in06 = reg_0619;
    76: op1_03_in06 = imem06_in[67:64];
    79: op1_03_in06 = reg_0363;
    80: op1_03_in06 = imem04_in[15:12];
    83: op1_03_in06 = imem06_in[51:48];
    84: op1_03_in06 = reg_0538;
    85: op1_03_in06 = reg_0275;
    86: op1_03_in06 = reg_0697;
    87: op1_03_in06 = reg_0473;
    88: op1_03_in06 = reg_0556;
    89: op1_03_in06 = reg_0322;
    90: op1_03_in06 = reg_0352;
    91: op1_03_in06 = reg_0590;
    92: op1_03_in06 = imem06_in[103:100];
    93: op1_03_in06 = imem06_in[23:20];
    94: op1_03_in06 = imem06_in[75:72];
    95: op1_03_in06 = imem06_in[55:52];
    96: op1_03_in06 = imem04_in[123:120];
    default: op1_03_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv06 = 1;
    8: op1_03_inv06 = 1;
    3: op1_03_inv06 = 1;
    12: op1_03_inv06 = 1;
    13: op1_03_inv06 = 1;
    19: op1_03_inv06 = 1;
    21: op1_03_inv06 = 1;
    23: op1_03_inv06 = 1;
    27: op1_03_inv06 = 1;
    30: op1_03_inv06 = 1;
    36: op1_03_inv06 = 1;
    37: op1_03_inv06 = 1;
    38: op1_03_inv06 = 1;
    40: op1_03_inv06 = 1;
    41: op1_03_inv06 = 1;
    44: op1_03_inv06 = 1;
    49: op1_03_inv06 = 1;
    53: op1_03_inv06 = 1;
    55: op1_03_inv06 = 1;
    56: op1_03_inv06 = 1;
    57: op1_03_inv06 = 1;
    58: op1_03_inv06 = 1;
    59: op1_03_inv06 = 1;
    60: op1_03_inv06 = 1;
    64: op1_03_inv06 = 1;
    65: op1_03_inv06 = 1;
    67: op1_03_inv06 = 1;
    68: op1_03_inv06 = 1;
    69: op1_03_inv06 = 1;
    70: op1_03_inv06 = 1;
    71: op1_03_inv06 = 1;
    74: op1_03_inv06 = 1;
    76: op1_03_inv06 = 1;
    80: op1_03_inv06 = 1;
    81: op1_03_inv06 = 1;
    84: op1_03_inv06 = 1;
    85: op1_03_inv06 = 1;
    89: op1_03_inv06 = 1;
    91: op1_03_inv06 = 1;
    93: op1_03_inv06 = 1;
    94: op1_03_inv06 = 1;
    95: op1_03_inv06 = 1;
    default: op1_03_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in07 = reg_0048;
    5: op1_03_in07 = reg_0325;
    6: op1_03_in07 = reg_0620;
    7: op1_03_in07 = imem02_in[115:112];
    8: op1_03_in07 = reg_0303;
    9: op1_03_in07 = reg_0062;
    3: op1_03_in07 = imem07_in[115:112];
    2: op1_03_in07 = reg_0158;
    10: op1_03_in07 = reg_0151;
    11: op1_03_in07 = reg_0807;
    12: op1_03_in07 = reg_0156;
    13: op1_03_in07 = imem02_in[75:72];
    14: op1_03_in07 = reg_0544;
    15: op1_03_in07 = reg_0137;
    16: op1_03_in07 = reg_0688;
    17: op1_03_in07 = imem04_in[31:28];
    18: op1_03_in07 = reg_0126;
    66: op1_03_in07 = reg_0126;
    19: op1_03_in07 = imem04_in[27:24];
    20: op1_03_in07 = reg_0191;
    21: op1_03_in07 = reg_0009;
    22: op1_03_in07 = imem05_in[127:124];
    23: op1_03_in07 = reg_0095;
    24: op1_03_in07 = reg_0381;
    25: op1_03_in07 = reg_0697;
    44: op1_03_in07 = reg_0697;
    26: op1_03_in07 = reg_0402;
    27: op1_03_in07 = reg_0463;
    71: op1_03_in07 = reg_0463;
    28: op1_03_in07 = reg_0083;
    29: op1_03_in07 = reg_0495;
    30: op1_03_in07 = reg_0464;
    31: op1_03_in07 = reg_0583;
    32: op1_03_in07 = imem05_in[7:4];
    33: op1_03_in07 = reg_0817;
    34: op1_03_in07 = reg_0555;
    35: op1_03_in07 = reg_0598;
    36: op1_03_in07 = reg_0051;
    37: op1_03_in07 = imem05_in[27:24];
    38: op1_03_in07 = reg_0484;
    40: op1_03_in07 = reg_0377;
    41: op1_03_in07 = reg_0506;
    42: op1_03_in07 = reg_0006;
    43: op1_03_in07 = reg_0277;
    45: op1_03_in07 = reg_0667;
    46: op1_03_in07 = reg_0090;
    47: op1_03_in07 = reg_0408;
    48: op1_03_in07 = reg_0362;
    49: op1_03_in07 = reg_0504;
    64: op1_03_in07 = reg_0504;
    50: op1_03_in07 = reg_0686;
    51: op1_03_in07 = reg_0375;
    53: op1_03_in07 = reg_0450;
    54: op1_03_in07 = reg_0735;
    55: op1_03_in07 = imem02_in[19:16];
    56: op1_03_in07 = reg_0573;
    57: op1_03_in07 = reg_0013;
    58: op1_03_in07 = reg_0639;
    59: op1_03_in07 = reg_0102;
    60: op1_03_in07 = reg_0552;
    61: op1_03_in07 = reg_0307;
    62: op1_03_in07 = reg_0633;
    63: op1_03_in07 = reg_0478;
    65: op1_03_in07 = imem02_in[95:92];
    67: op1_03_in07 = reg_0427;
    68: op1_03_in07 = reg_0707;
    69: op1_03_in07 = reg_0494;
    70: op1_03_in07 = reg_0582;
    72: op1_03_in07 = reg_0290;
    73: op1_03_in07 = reg_0139;
    74: op1_03_in07 = reg_0557;
    75: op1_03_in07 = reg_0766;
    76: op1_03_in07 = imem06_in[99:96];
    78: op1_03_in07 = reg_0676;
    79: op1_03_in07 = reg_0594;
    80: op1_03_in07 = imem04_in[63:60];
    81: op1_03_in07 = reg_0649;
    83: op1_03_in07 = imem06_in[67:64];
    84: op1_03_in07 = reg_0642;
    85: op1_03_in07 = reg_0534;
    86: op1_03_in07 = reg_0758;
    87: op1_03_in07 = reg_0467;
    88: op1_03_in07 = reg_0615;
    89: op1_03_in07 = reg_0274;
    90: op1_03_in07 = reg_0344;
    91: op1_03_in07 = reg_0343;
    92: op1_03_in07 = reg_0625;
    93: op1_03_in07 = imem06_in[39:36];
    94: op1_03_in07 = imem06_in[83:80];
    95: op1_03_in07 = imem06_in[59:56];
    96: op1_03_in07 = reg_0545;
    default: op1_03_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv07 = 1;
    6: op1_03_inv07 = 1;
    8: op1_03_inv07 = 1;
    3: op1_03_inv07 = 1;
    11: op1_03_inv07 = 1;
    13: op1_03_inv07 = 1;
    17: op1_03_inv07 = 1;
    19: op1_03_inv07 = 1;
    20: op1_03_inv07 = 1;
    22: op1_03_inv07 = 1;
    28: op1_03_inv07 = 1;
    30: op1_03_inv07 = 1;
    32: op1_03_inv07 = 1;
    34: op1_03_inv07 = 1;
    36: op1_03_inv07 = 1;
    38: op1_03_inv07 = 1;
    41: op1_03_inv07 = 1;
    47: op1_03_inv07 = 1;
    48: op1_03_inv07 = 1;
    50: op1_03_inv07 = 1;
    58: op1_03_inv07 = 1;
    59: op1_03_inv07 = 1;
    60: op1_03_inv07 = 1;
    61: op1_03_inv07 = 1;
    64: op1_03_inv07 = 1;
    68: op1_03_inv07 = 1;
    69: op1_03_inv07 = 1;
    71: op1_03_inv07 = 1;
    72: op1_03_inv07 = 1;
    76: op1_03_inv07 = 1;
    80: op1_03_inv07 = 1;
    81: op1_03_inv07 = 1;
    83: op1_03_inv07 = 1;
    85: op1_03_inv07 = 1;
    86: op1_03_inv07 = 1;
    87: op1_03_inv07 = 1;
    89: op1_03_inv07 = 1;
    90: op1_03_inv07 = 1;
    93: op1_03_inv07 = 1;
    94: op1_03_inv07 = 1;
    96: op1_03_inv07 = 1;
    default: op1_03_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in08 = reg_0063;
    5: op1_03_in08 = reg_0326;
    6: op1_03_in08 = reg_0616;
    7: op1_03_in08 = reg_0660;
    8: op1_03_in08 = reg_0290;
    9: op1_03_in08 = reg_0056;
    3: op1_03_in08 = imem07_in[127:124];
    2: op1_03_in08 = reg_0171;
    10: op1_03_in08 = reg_0153;
    11: op1_03_in08 = reg_0801;
    12: op1_03_in08 = reg_0154;
    13: op1_03_in08 = imem02_in[83:80];
    14: op1_03_in08 = reg_0530;
    15: op1_03_in08 = reg_0134;
    16: op1_03_in08 = reg_0453;
    27: op1_03_in08 = reg_0453;
    17: op1_03_in08 = imem04_in[51:48];
    18: op1_03_in08 = reg_0110;
    19: op1_03_in08 = imem04_in[67:64];
    20: op1_03_in08 = reg_0203;
    21: op1_03_in08 = imem04_in[39:36];
    22: op1_03_in08 = reg_0792;
    23: op1_03_in08 = reg_0757;
    24: op1_03_in08 = reg_0392;
    25: op1_03_in08 = reg_0685;
    26: op1_03_in08 = reg_0379;
    28: op1_03_in08 = reg_0060;
    85: op1_03_in08 = reg_0060;
    29: op1_03_in08 = reg_0309;
    30: op1_03_in08 = reg_0472;
    31: op1_03_in08 = reg_0592;
    32: op1_03_in08 = imem05_in[11:8];
    33: op1_03_in08 = reg_0338;
    34: op1_03_in08 = reg_0551;
    35: op1_03_in08 = reg_0601;
    36: op1_03_in08 = reg_0074;
    37: op1_03_in08 = imem05_in[71:68];
    38: op1_03_in08 = reg_0788;
    40: op1_03_in08 = reg_0406;
    41: op1_03_in08 = reg_0219;
    42: op1_03_in08 = reg_0015;
    43: op1_03_in08 = reg_0128;
    44: op1_03_in08 = reg_0694;
    45: op1_03_in08 = reg_0344;
    46: op1_03_in08 = reg_0225;
    47: op1_03_in08 = reg_0377;
    48: op1_03_in08 = reg_0320;
    49: op1_03_in08 = reg_0419;
    50: op1_03_in08 = reg_0691;
    51: op1_03_in08 = reg_0238;
    76: op1_03_in08 = reg_0238;
    53: op1_03_in08 = reg_0477;
    71: op1_03_in08 = reg_0477;
    54: op1_03_in08 = reg_0237;
    55: op1_03_in08 = imem02_in[35:32];
    56: op1_03_in08 = reg_0385;
    57: op1_03_in08 = reg_0007;
    58: op1_03_in08 = reg_0651;
    59: op1_03_in08 = reg_0249;
    60: op1_03_in08 = reg_0055;
    61: op1_03_in08 = reg_0257;
    62: op1_03_in08 = reg_0465;
    63: op1_03_in08 = reg_0200;
    64: op1_03_in08 = reg_0678;
    65: op1_03_in08 = reg_0089;
    66: op1_03_in08 = imem02_in[11:8];
    67: op1_03_in08 = reg_0586;
    68: op1_03_in08 = reg_0295;
    69: op1_03_in08 = reg_0634;
    70: op1_03_in08 = reg_0319;
    72: op1_03_in08 = reg_0425;
    73: op1_03_in08 = reg_0704;
    74: op1_03_in08 = reg_0623;
    75: op1_03_in08 = reg_0339;
    78: op1_03_in08 = reg_0674;
    79: op1_03_in08 = reg_0353;
    80: op1_03_in08 = imem04_in[79:76];
    81: op1_03_in08 = reg_0570;
    83: op1_03_in08 = imem06_in[71:68];
    84: op1_03_in08 = reg_0541;
    86: op1_03_in08 = reg_0494;
    87: op1_03_in08 = reg_0471;
    88: op1_03_in08 = reg_0077;
    89: op1_03_in08 = reg_0362;
    90: op1_03_in08 = reg_0341;
    91: op1_03_in08 = reg_0743;
    92: op1_03_in08 = reg_0605;
    93: op1_03_in08 = imem06_in[79:76];
    94: op1_03_in08 = imem06_in[91:88];
    95: op1_03_in08 = reg_0577;
    96: op1_03_in08 = reg_0058;
    default: op1_03_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_03_inv08 = 1;
    3: op1_03_inv08 = 1;
    11: op1_03_inv08 = 1;
    12: op1_03_inv08 = 1;
    13: op1_03_inv08 = 1;
    14: op1_03_inv08 = 1;
    16: op1_03_inv08 = 1;
    19: op1_03_inv08 = 1;
    20: op1_03_inv08 = 1;
    23: op1_03_inv08 = 1;
    24: op1_03_inv08 = 1;
    25: op1_03_inv08 = 1;
    27: op1_03_inv08 = 1;
    28: op1_03_inv08 = 1;
    30: op1_03_inv08 = 1;
    32: op1_03_inv08 = 1;
    33: op1_03_inv08 = 1;
    34: op1_03_inv08 = 1;
    35: op1_03_inv08 = 1;
    36: op1_03_inv08 = 1;
    38: op1_03_inv08 = 1;
    40: op1_03_inv08 = 1;
    43: op1_03_inv08 = 1;
    47: op1_03_inv08 = 1;
    49: op1_03_inv08 = 1;
    50: op1_03_inv08 = 1;
    55: op1_03_inv08 = 1;
    56: op1_03_inv08 = 1;
    57: op1_03_inv08 = 1;
    58: op1_03_inv08 = 1;
    59: op1_03_inv08 = 1;
    62: op1_03_inv08 = 1;
    65: op1_03_inv08 = 1;
    66: op1_03_inv08 = 1;
    71: op1_03_inv08 = 1;
    72: op1_03_inv08 = 1;
    73: op1_03_inv08 = 1;
    74: op1_03_inv08 = 1;
    75: op1_03_inv08 = 1;
    76: op1_03_inv08 = 1;
    79: op1_03_inv08 = 1;
    80: op1_03_inv08 = 1;
    81: op1_03_inv08 = 1;
    84: op1_03_inv08 = 1;
    86: op1_03_inv08 = 1;
    88: op1_03_inv08 = 1;
    92: op1_03_inv08 = 1;
    94: op1_03_inv08 = 1;
    default: op1_03_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in09 = reg_0064;
    5: op1_03_in09 = reg_0354;
    6: op1_03_in09 = reg_0631;
    7: op1_03_in09 = reg_0353;
    8: op1_03_in09 = reg_0296;
    9: op1_03_in09 = reg_0043;
    3: op1_03_in09 = reg_0424;
    49: op1_03_in09 = reg_0424;
    10: op1_03_in09 = reg_0141;
    12: op1_03_in09 = reg_0141;
    11: op1_03_in09 = reg_0800;
    57: op1_03_in09 = reg_0800;
    13: op1_03_in09 = imem02_in[103:100];
    14: op1_03_in09 = reg_0542;
    15: op1_03_in09 = imem06_in[7:4];
    16: op1_03_in09 = reg_0476;
    53: op1_03_in09 = reg_0476;
    69: op1_03_in09 = reg_0476;
    17: op1_03_in09 = imem04_in[63:60];
    18: op1_03_in09 = imem02_in[7:4];
    19: op1_03_in09 = imem04_in[75:72];
    20: op1_03_in09 = reg_0186;
    21: op1_03_in09 = imem04_in[79:76];
    22: op1_03_in09 = reg_0780;
    23: op1_03_in09 = reg_0094;
    24: op1_03_in09 = reg_0351;
    25: op1_03_in09 = reg_0676;
    26: op1_03_in09 = reg_0381;
    27: op1_03_in09 = reg_0451;
    28: op1_03_in09 = reg_0551;
    29: op1_03_in09 = reg_0084;
    30: op1_03_in09 = reg_0470;
    31: op1_03_in09 = reg_0591;
    35: op1_03_in09 = reg_0591;
    32: op1_03_in09 = imem05_in[27:24];
    33: op1_03_in09 = reg_0339;
    34: op1_03_in09 = reg_0274;
    36: op1_03_in09 = imem05_in[19:16];
    37: op1_03_in09 = imem05_in[99:96];
    38: op1_03_in09 = reg_0493;
    40: op1_03_in09 = reg_0038;
    41: op1_03_in09 = reg_0120;
    42: op1_03_in09 = reg_0799;
    43: op1_03_in09 = reg_0129;
    44: op1_03_in09 = reg_0691;
    45: op1_03_in09 = reg_0341;
    46: op1_03_in09 = reg_0272;
    47: op1_03_in09 = reg_0403;
    48: op1_03_in09 = reg_0342;
    79: op1_03_in09 = reg_0342;
    50: op1_03_in09 = reg_0674;
    51: op1_03_in09 = reg_0029;
    54: op1_03_in09 = reg_0557;
    55: op1_03_in09 = imem02_in[75:72];
    56: op1_03_in09 = reg_0562;
    58: op1_03_in09 = reg_0427;
    59: op1_03_in09 = reg_0066;
    60: op1_03_in09 = reg_0536;
    61: op1_03_in09 = reg_0148;
    62: op1_03_in09 = reg_0457;
    63: op1_03_in09 = reg_0203;
    64: op1_03_in09 = imem02_in[3:0];
    65: op1_03_in09 = reg_0584;
    66: op1_03_in09 = imem02_in[35:32];
    67: op1_03_in09 = reg_0565;
    68: op1_03_in09 = reg_0447;
    70: op1_03_in09 = reg_0350;
    71: op1_03_in09 = reg_0462;
    72: op1_03_in09 = reg_0123;
    73: op1_03_in09 = reg_0138;
    74: op1_03_in09 = reg_0649;
    75: op1_03_in09 = reg_0265;
    76: op1_03_in09 = reg_0580;
    78: op1_03_in09 = imem02_in[11:8];
    80: op1_03_in09 = imem04_in[95:92];
    81: op1_03_in09 = reg_0001;
    83: op1_03_in09 = imem06_in[79:76];
    84: op1_03_in09 = reg_0704;
    85: op1_03_in09 = reg_0331;
    86: op1_03_in09 = reg_0450;
    87: op1_03_in09 = reg_0208;
    88: op1_03_in09 = reg_0071;
    89: op1_03_in09 = reg_0364;
    90: op1_03_in09 = reg_0324;
    91: op1_03_in09 = reg_0487;
    92: op1_03_in09 = reg_0409;
    93: op1_03_in09 = reg_0291;
    94: op1_03_in09 = imem06_in[107:104];
    95: op1_03_in09 = reg_0817;
    96: op1_03_in09 = reg_0179;
    default: op1_03_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv09 = 1;
    5: op1_03_inv09 = 1;
    10: op1_03_inv09 = 1;
    13: op1_03_inv09 = 1;
    14: op1_03_inv09 = 1;
    17: op1_03_inv09 = 1;
    18: op1_03_inv09 = 1;
    19: op1_03_inv09 = 1;
    20: op1_03_inv09 = 1;
    22: op1_03_inv09 = 1;
    23: op1_03_inv09 = 1;
    24: op1_03_inv09 = 1;
    26: op1_03_inv09 = 1;
    28: op1_03_inv09 = 1;
    29: op1_03_inv09 = 1;
    30: op1_03_inv09 = 1;
    31: op1_03_inv09 = 1;
    33: op1_03_inv09 = 1;
    36: op1_03_inv09 = 1;
    37: op1_03_inv09 = 1;
    38: op1_03_inv09 = 1;
    40: op1_03_inv09 = 1;
    41: op1_03_inv09 = 1;
    44: op1_03_inv09 = 1;
    45: op1_03_inv09 = 1;
    46: op1_03_inv09 = 1;
    51: op1_03_inv09 = 1;
    53: op1_03_inv09 = 1;
    54: op1_03_inv09 = 1;
    55: op1_03_inv09 = 1;
    56: op1_03_inv09 = 1;
    63: op1_03_inv09 = 1;
    64: op1_03_inv09 = 1;
    66: op1_03_inv09 = 1;
    68: op1_03_inv09 = 1;
    71: op1_03_inv09 = 1;
    72: op1_03_inv09 = 1;
    73: op1_03_inv09 = 1;
    74: op1_03_inv09 = 1;
    75: op1_03_inv09 = 1;
    76: op1_03_inv09 = 1;
    79: op1_03_inv09 = 1;
    83: op1_03_inv09 = 1;
    84: op1_03_inv09 = 1;
    85: op1_03_inv09 = 1;
    86: op1_03_inv09 = 1;
    94: op1_03_inv09 = 1;
    95: op1_03_inv09 = 1;
    default: op1_03_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in10 = imem05_in[23:20];
    5: op1_03_in10 = reg_0355;
    6: op1_03_in10 = reg_0632;
    7: op1_03_in10 = reg_0350;
    8: op1_03_in10 = reg_0298;
    9: op1_03_in10 = reg_0053;
    3: op1_03_in10 = reg_0446;
    10: op1_03_in10 = reg_0140;
    11: op1_03_in10 = reg_0799;
    12: op1_03_in10 = reg_0130;
    13: op1_03_in10 = reg_0660;
    14: op1_03_in10 = reg_0548;
    15: op1_03_in10 = imem06_in[47:44];
    16: op1_03_in10 = reg_0470;
    53: op1_03_in10 = reg_0470;
    17: op1_03_in10 = imem04_in[67:64];
    18: op1_03_in10 = imem02_in[11:8];
    19: op1_03_in10 = imem04_in[91:88];
    20: op1_03_in10 = imem01_in[59:56];
    21: op1_03_in10 = imem04_in[83:80];
    22: op1_03_in10 = reg_0786;
    23: op1_03_in10 = reg_0740;
    24: op1_03_in10 = reg_0375;
    25: op1_03_in10 = reg_0466;
    26: op1_03_in10 = reg_0408;
    27: op1_03_in10 = reg_0455;
    86: op1_03_in10 = reg_0455;
    28: op1_03_in10 = reg_0500;
    29: op1_03_in10 = reg_0142;
    30: op1_03_in10 = reg_0474;
    31: op1_03_in10 = reg_0589;
    32: op1_03_in10 = imem05_in[67:64];
    33: op1_03_in10 = imem07_in[23:20];
    34: op1_03_in10 = reg_0050;
    88: op1_03_in10 = reg_0050;
    35: op1_03_in10 = reg_0600;
    36: op1_03_in10 = imem05_in[35:32];
    37: op1_03_in10 = reg_0798;
    38: op1_03_in10 = reg_0495;
    40: op1_03_in10 = reg_0311;
    41: op1_03_in10 = reg_0117;
    42: op1_03_in10 = reg_0009;
    43: op1_03_in10 = reg_0153;
    44: op1_03_in10 = reg_0673;
    45: op1_03_in10 = reg_0348;
    46: op1_03_in10 = reg_0744;
    47: op1_03_in10 = reg_0776;
    48: op1_03_in10 = reg_0314;
    49: op1_03_in10 = reg_0219;
    50: op1_03_in10 = reg_0692;
    51: op1_03_in10 = reg_0752;
    54: op1_03_in10 = reg_0652;
    55: op1_03_in10 = imem02_in[111:108];
    56: op1_03_in10 = reg_0001;
    57: op1_03_in10 = reg_0805;
    58: op1_03_in10 = reg_0336;
    59: op1_03_in10 = reg_0101;
    60: op1_03_in10 = reg_0429;
    85: op1_03_in10 = reg_0429;
    61: op1_03_in10 = reg_0135;
    62: op1_03_in10 = reg_0464;
    63: op1_03_in10 = reg_0213;
    64: op1_03_in10 = imem02_in[55:52];
    65: op1_03_in10 = reg_0621;
    66: op1_03_in10 = reg_0045;
    67: op1_03_in10 = reg_0530;
    68: op1_03_in10 = reg_0445;
    69: op1_03_in10 = reg_0187;
    70: op1_03_in10 = reg_0571;
    71: op1_03_in10 = reg_0472;
    72: op1_03_in10 = reg_0125;
    73: op1_03_in10 = reg_0586;
    74: op1_03_in10 = reg_0013;
    75: op1_03_in10 = reg_0369;
    76: op1_03_in10 = reg_0664;
    78: op1_03_in10 = imem02_in[71:68];
    79: op1_03_in10 = reg_0590;
    80: op1_03_in10 = reg_0316;
    81: op1_03_in10 = reg_0003;
    83: op1_03_in10 = imem06_in[87:84];
    84: op1_03_in10 = reg_0075;
    87: op1_03_in10 = reg_0207;
    89: op1_03_in10 = reg_0320;
    90: op1_03_in10 = reg_0527;
    91: op1_03_in10 = reg_0055;
    92: op1_03_in10 = reg_0238;
    93: op1_03_in10 = reg_0814;
    95: op1_03_in10 = reg_0814;
    94: op1_03_in10 = reg_0289;
    96: op1_03_in10 = reg_0539;
    default: op1_03_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv10 = 1;
    7: op1_03_inv10 = 1;
    8: op1_03_inv10 = 1;
    3: op1_03_inv10 = 1;
    10: op1_03_inv10 = 1;
    12: op1_03_inv10 = 1;
    14: op1_03_inv10 = 1;
    16: op1_03_inv10 = 1;
    17: op1_03_inv10 = 1;
    18: op1_03_inv10 = 1;
    19: op1_03_inv10 = 1;
    20: op1_03_inv10 = 1;
    21: op1_03_inv10 = 1;
    22: op1_03_inv10 = 1;
    24: op1_03_inv10 = 1;
    28: op1_03_inv10 = 1;
    29: op1_03_inv10 = 1;
    31: op1_03_inv10 = 1;
    34: op1_03_inv10 = 1;
    37: op1_03_inv10 = 1;
    38: op1_03_inv10 = 1;
    42: op1_03_inv10 = 1;
    44: op1_03_inv10 = 1;
    46: op1_03_inv10 = 1;
    51: op1_03_inv10 = 1;
    54: op1_03_inv10 = 1;
    56: op1_03_inv10 = 1;
    57: op1_03_inv10 = 1;
    59: op1_03_inv10 = 1;
    60: op1_03_inv10 = 1;
    62: op1_03_inv10 = 1;
    64: op1_03_inv10 = 1;
    65: op1_03_inv10 = 1;
    67: op1_03_inv10 = 1;
    69: op1_03_inv10 = 1;
    70: op1_03_inv10 = 1;
    71: op1_03_inv10 = 1;
    72: op1_03_inv10 = 1;
    73: op1_03_inv10 = 1;
    74: op1_03_inv10 = 1;
    75: op1_03_inv10 = 1;
    85: op1_03_inv10 = 1;
    87: op1_03_inv10 = 1;
    88: op1_03_inv10 = 1;
    94: op1_03_inv10 = 1;
    95: op1_03_inv10 = 1;
    96: op1_03_inv10 = 1;
    default: op1_03_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in11 = reg_0482;
    5: op1_03_in11 = reg_0335;
    6: op1_03_in11 = reg_0351;
    7: op1_03_in11 = reg_0083;
    80: op1_03_in11 = reg_0083;
    8: op1_03_in11 = reg_0307;
    9: op1_03_in11 = reg_0063;
    3: op1_03_in11 = reg_0174;
    10: op1_03_in11 = reg_0131;
    11: op1_03_in11 = reg_0810;
    12: op1_03_in11 = reg_0137;
    13: op1_03_in11 = reg_0661;
    14: op1_03_in11 = reg_0558;
    15: op1_03_in11 = imem06_in[115:112];
    16: op1_03_in11 = reg_0456;
    71: op1_03_in11 = reg_0456;
    17: op1_03_in11 = imem04_in[79:76];
    18: op1_03_in11 = imem02_in[91:88];
    64: op1_03_in11 = imem02_in[91:88];
    19: op1_03_in11 = reg_0557;
    20: op1_03_in11 = imem01_in[67:64];
    21: op1_03_in11 = imem04_in[95:92];
    22: op1_03_in11 = reg_0485;
    23: op1_03_in11 = imem03_in[59:56];
    91: op1_03_in11 = imem03_in[59:56];
    24: op1_03_in11 = reg_0390;
    25: op1_03_in11 = reg_0475;
    26: op1_03_in11 = reg_0386;
    27: op1_03_in11 = reg_0476;
    28: op1_03_in11 = reg_0298;
    95: op1_03_in11 = reg_0298;
    29: op1_03_in11 = reg_0156;
    30: op1_03_in11 = reg_0459;
    31: op1_03_in11 = reg_0600;
    32: op1_03_in11 = reg_0797;
    37: op1_03_in11 = reg_0797;
    33: op1_03_in11 = imem07_in[27:24];
    34: op1_03_in11 = reg_0061;
    35: op1_03_in11 = reg_0387;
    36: op1_03_in11 = imem05_in[51:48];
    38: op1_03_in11 = reg_0794;
    40: op1_03_in11 = reg_0242;
    41: op1_03_in11 = reg_0126;
    42: op1_03_in11 = imem04_in[47:44];
    43: op1_03_in11 = imem06_in[31:28];
    44: op1_03_in11 = reg_0699;
    45: op1_03_in11 = reg_0322;
    84: op1_03_in11 = reg_0322;
    46: op1_03_in11 = reg_0285;
    47: op1_03_in11 = reg_0404;
    48: op1_03_in11 = reg_0533;
    49: op1_03_in11 = reg_0111;
    50: op1_03_in11 = reg_0465;
    51: op1_03_in11 = imem07_in[23:20];
    53: op1_03_in11 = reg_0207;
    54: op1_03_in11 = reg_0737;
    55: op1_03_in11 = imem02_in[123:120];
    56: op1_03_in11 = reg_0803;
    57: op1_03_in11 = reg_0016;
    58: op1_03_in11 = reg_0565;
    59: op1_03_in11 = reg_0136;
    60: op1_03_in11 = reg_0280;
    61: op1_03_in11 = reg_0138;
    62: op1_03_in11 = reg_0477;
    63: op1_03_in11 = reg_0205;
    65: op1_03_in11 = reg_0651;
    66: op1_03_in11 = reg_0666;
    67: op1_03_in11 = reg_0096;
    68: op1_03_in11 = reg_0439;
    69: op1_03_in11 = reg_0193;
    70: op1_03_in11 = reg_0417;
    72: op1_03_in11 = reg_0120;
    73: op1_03_in11 = reg_0345;
    74: op1_03_in11 = reg_0805;
    75: op1_03_in11 = reg_0630;
    76: op1_03_in11 = reg_0501;
    78: op1_03_in11 = imem02_in[75:72];
    79: op1_03_in11 = reg_0092;
    81: op1_03_in11 = reg_0801;
    83: op1_03_in11 = imem06_in[103:100];
    85: op1_03_in11 = reg_0079;
    86: op1_03_in11 = reg_0469;
    87: op1_03_in11 = reg_0211;
    88: op1_03_in11 = reg_0585;
    89: op1_03_in11 = reg_0594;
    90: op1_03_in11 = reg_0770;
    92: op1_03_in11 = reg_0265;
    93: op1_03_in11 = reg_0766;
    94: op1_03_in11 = reg_0291;
    96: op1_03_in11 = reg_0261;
    default: op1_03_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv11 = 1;
    9: op1_03_inv11 = 1;
    10: op1_03_inv11 = 1;
    11: op1_03_inv11 = 1;
    13: op1_03_inv11 = 1;
    14: op1_03_inv11 = 1;
    16: op1_03_inv11 = 1;
    18: op1_03_inv11 = 1;
    19: op1_03_inv11 = 1;
    23: op1_03_inv11 = 1;
    25: op1_03_inv11 = 1;
    29: op1_03_inv11 = 1;
    30: op1_03_inv11 = 1;
    32: op1_03_inv11 = 1;
    35: op1_03_inv11 = 1;
    36: op1_03_inv11 = 1;
    38: op1_03_inv11 = 1;
    40: op1_03_inv11 = 1;
    42: op1_03_inv11 = 1;
    44: op1_03_inv11 = 1;
    45: op1_03_inv11 = 1;
    46: op1_03_inv11 = 1;
    48: op1_03_inv11 = 1;
    49: op1_03_inv11 = 1;
    50: op1_03_inv11 = 1;
    53: op1_03_inv11 = 1;
    56: op1_03_inv11 = 1;
    58: op1_03_inv11 = 1;
    59: op1_03_inv11 = 1;
    61: op1_03_inv11 = 1;
    62: op1_03_inv11 = 1;
    63: op1_03_inv11 = 1;
    65: op1_03_inv11 = 1;
    67: op1_03_inv11 = 1;
    68: op1_03_inv11 = 1;
    70: op1_03_inv11 = 1;
    71: op1_03_inv11 = 1;
    73: op1_03_inv11 = 1;
    75: op1_03_inv11 = 1;
    78: op1_03_inv11 = 1;
    79: op1_03_inv11 = 1;
    80: op1_03_inv11 = 1;
    81: op1_03_inv11 = 1;
    83: op1_03_inv11 = 1;
    88: op1_03_inv11 = 1;
    89: op1_03_inv11 = 1;
    90: op1_03_inv11 = 1;
    91: op1_03_inv11 = 1;
    default: op1_03_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in12 = reg_0483;
    5: op1_03_in12 = reg_0042;
    7: op1_03_in12 = reg_0042;
    6: op1_03_in12 = reg_0025;
    8: op1_03_in12 = reg_0284;
    9: op1_03_in12 = imem05_in[7:4];
    3: op1_03_in12 = reg_0180;
    10: op1_03_in12 = reg_0134;
    11: op1_03_in12 = reg_0009;
    12: op1_03_in12 = imem06_in[39:36];
    13: op1_03_in12 = reg_0636;
    14: op1_03_in12 = reg_0533;
    15: op1_03_in12 = reg_0628;
    92: op1_03_in12 = reg_0628;
    16: op1_03_in12 = reg_0200;
    17: op1_03_in12 = imem05_in[91:88];
    18: op1_03_in12 = reg_0655;
    19: op1_03_in12 = reg_0552;
    20: op1_03_in12 = imem01_in[75:72];
    21: op1_03_in12 = reg_0305;
    22: op1_03_in12 = reg_0787;
    23: op1_03_in12 = imem03_in[123:120];
    24: op1_03_in12 = reg_0039;
    25: op1_03_in12 = reg_0472;
    26: op1_03_in12 = reg_0382;
    27: op1_03_in12 = reg_0471;
    28: op1_03_in12 = reg_0299;
    29: op1_03_in12 = reg_0139;
    30: op1_03_in12 = reg_0214;
    71: op1_03_in12 = reg_0214;
    31: op1_03_in12 = reg_0580;
    32: op1_03_in12 = reg_0795;
    33: op1_03_in12 = imem07_in[35:32];
    34: op1_03_in12 = reg_0067;
    35: op1_03_in12 = reg_0755;
    36: op1_03_in12 = imem05_in[75:72];
    37: op1_03_in12 = reg_0484;
    38: op1_03_in12 = reg_0485;
    40: op1_03_in12 = reg_0815;
    41: op1_03_in12 = reg_0110;
    42: op1_03_in12 = imem04_in[55:52];
    43: op1_03_in12 = reg_0218;
    44: op1_03_in12 = reg_0463;
    45: op1_03_in12 = reg_0321;
    46: op1_03_in12 = reg_0149;
    47: op1_03_in12 = reg_0329;
    48: op1_03_in12 = reg_0540;
    49: op1_03_in12 = reg_0108;
    50: op1_03_in12 = reg_0481;
    51: op1_03_in12 = imem07_in[51:48];
    53: op1_03_in12 = reg_0198;
    69: op1_03_in12 = reg_0198;
    54: op1_03_in12 = reg_0235;
    55: op1_03_in12 = reg_0642;
    56: op1_03_in12 = reg_0015;
    57: op1_03_in12 = reg_0004;
    58: op1_03_in12 = reg_0361;
    59: op1_03_in12 = reg_0144;
    60: op1_03_in12 = reg_0615;
    61: op1_03_in12 = reg_0140;
    62: op1_03_in12 = reg_0475;
    63: op1_03_in12 = imem01_in[27:24];
    64: op1_03_in12 = reg_0657;
    65: op1_03_in12 = reg_0548;
    66: op1_03_in12 = reg_0637;
    67: op1_03_in12 = imem03_in[127:124];
    68: op1_03_in12 = reg_0175;
    70: op1_03_in12 = reg_0490;
    72: op1_03_in12 = reg_0660;
    73: op1_03_in12 = reg_0365;
    74: op1_03_in12 = reg_0809;
    75: op1_03_in12 = reg_0408;
    76: op1_03_in12 = reg_0632;
    78: op1_03_in12 = imem02_in[99:96];
    79: op1_03_in12 = reg_0081;
    80: op1_03_in12 = reg_0554;
    81: op1_03_in12 = reg_0008;
    83: op1_03_in12 = reg_0289;
    84: op1_03_in12 = reg_0251;
    85: op1_03_in12 = reg_0631;
    86: op1_03_in12 = reg_0460;
    87: op1_03_in12 = reg_0213;
    88: op1_03_in12 = reg_0780;
    89: op1_03_in12 = reg_0342;
    90: op1_03_in12 = imem03_in[31:28];
    91: op1_03_in12 = imem03_in[83:80];
    93: op1_03_in12 = reg_0578;
    94: op1_03_in12 = reg_0409;
    95: op1_03_in12 = reg_0354;
    96: op1_03_in12 = reg_0331;
    default: op1_03_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv12 = 1;
    6: op1_03_inv12 = 1;
    7: op1_03_inv12 = 1;
    8: op1_03_inv12 = 1;
    9: op1_03_inv12 = 1;
    3: op1_03_inv12 = 1;
    12: op1_03_inv12 = 1;
    17: op1_03_inv12 = 1;
    19: op1_03_inv12 = 1;
    26: op1_03_inv12 = 1;
    29: op1_03_inv12 = 1;
    31: op1_03_inv12 = 1;
    32: op1_03_inv12 = 1;
    33: op1_03_inv12 = 1;
    34: op1_03_inv12 = 1;
    36: op1_03_inv12 = 1;
    38: op1_03_inv12 = 1;
    40: op1_03_inv12 = 1;
    45: op1_03_inv12 = 1;
    46: op1_03_inv12 = 1;
    47: op1_03_inv12 = 1;
    48: op1_03_inv12 = 1;
    50: op1_03_inv12 = 1;
    51: op1_03_inv12 = 1;
    53: op1_03_inv12 = 1;
    54: op1_03_inv12 = 1;
    55: op1_03_inv12 = 1;
    57: op1_03_inv12 = 1;
    58: op1_03_inv12 = 1;
    59: op1_03_inv12 = 1;
    61: op1_03_inv12 = 1;
    62: op1_03_inv12 = 1;
    66: op1_03_inv12 = 1;
    67: op1_03_inv12 = 1;
    68: op1_03_inv12 = 1;
    73: op1_03_inv12 = 1;
    74: op1_03_inv12 = 1;
    76: op1_03_inv12 = 1;
    80: op1_03_inv12 = 1;
    81: op1_03_inv12 = 1;
    83: op1_03_inv12 = 1;
    84: op1_03_inv12 = 1;
    85: op1_03_inv12 = 1;
    86: op1_03_inv12 = 1;
    88: op1_03_inv12 = 1;
    90: op1_03_inv12 = 1;
    91: op1_03_inv12 = 1;
    92: op1_03_inv12 = 1;
    94: op1_03_inv12 = 1;
    default: op1_03_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in13 = reg_0484;
    5: op1_03_in13 = reg_0088;
    6: op1_03_in13 = reg_0030;
    7: op1_03_in13 = reg_0089;
    8: op1_03_in13 = reg_0074;
    9: op1_03_in13 = imem05_in[27:24];
    3: op1_03_in13 = reg_0169;
    10: op1_03_in13 = reg_0144;
    11: op1_03_in13 = imem04_in[27:24];
    12: op1_03_in13 = imem06_in[79:76];
    13: op1_03_in13 = reg_0667;
    14: op1_03_in13 = reg_0541;
    15: op1_03_in13 = reg_0610;
    16: op1_03_in13 = reg_0194;
    17: op1_03_in13 = imem05_in[95:92];
    18: op1_03_in13 = reg_0661;
    64: op1_03_in13 = reg_0661;
    19: op1_03_in13 = reg_0539;
    20: op1_03_in13 = imem01_in[79:76];
    21: op1_03_in13 = reg_0290;
    22: op1_03_in13 = reg_0136;
    23: op1_03_in13 = reg_0598;
    24: op1_03_in13 = reg_0753;
    25: op1_03_in13 = reg_0213;
    26: op1_03_in13 = reg_0383;
    27: op1_03_in13 = reg_0209;
    28: op1_03_in13 = reg_0067;
    29: op1_03_in13 = reg_0137;
    30: op1_03_in13 = reg_0210;
    31: op1_03_in13 = reg_0395;
    32: op1_03_in13 = reg_0780;
    33: op1_03_in13 = imem07_in[47:44];
    34: op1_03_in13 = reg_0068;
    35: op1_03_in13 = reg_0373;
    36: op1_03_in13 = reg_0796;
    37: op1_03_in13 = reg_0493;
    38: op1_03_in13 = reg_0741;
    40: op1_03_in13 = reg_0621;
    41: op1_03_in13 = imem02_in[19:16];
    42: op1_03_in13 = imem04_in[59:56];
    43: op1_03_in13 = reg_0298;
    44: op1_03_in13 = reg_0451;
    45: op1_03_in13 = reg_0743;
    46: op1_03_in13 = reg_0151;
    47: op1_03_in13 = reg_0311;
    48: op1_03_in13 = reg_0535;
    49: op1_03_in13 = reg_0106;
    50: op1_03_in13 = reg_0470;
    51: op1_03_in13 = imem07_in[63:60];
    53: op1_03_in13 = reg_0201;
    69: op1_03_in13 = reg_0201;
    54: op1_03_in13 = reg_0306;
    55: op1_03_in13 = reg_0650;
    56: op1_03_in13 = reg_0016;
    57: op1_03_in13 = imem04_in[11:8];
    58: op1_03_in13 = reg_0092;
    59: op1_03_in13 = imem06_in[31:28];
    60: op1_03_in13 = reg_0077;
    61: op1_03_in13 = reg_0155;
    62: op1_03_in13 = reg_0460;
    63: op1_03_in13 = imem01_in[35:32];
    65: op1_03_in13 = reg_0237;
    66: op1_03_in13 = reg_0563;
    67: op1_03_in13 = reg_0319;
    68: op1_03_in13 = reg_0162;
    70: op1_03_in13 = reg_0570;
    71: op1_03_in13 = reg_0208;
    72: op1_03_in13 = reg_0674;
    73: op1_03_in13 = reg_0323;
    74: op1_03_in13 = imem04_in[3:0];
    75: op1_03_in13 = reg_0608;
    76: op1_03_in13 = reg_0367;
    78: op1_03_in13 = reg_0739;
    79: op1_03_in13 = reg_0095;
    80: op1_03_in13 = reg_0558;
    81: op1_03_in13 = reg_0802;
    83: op1_03_in13 = reg_0299;
    84: op1_03_in13 = reg_0594;
    85: op1_03_in13 = reg_0302;
    86: op1_03_in13 = reg_0471;
    87: op1_03_in13 = reg_0190;
    88: op1_03_in13 = reg_0643;
    89: op1_03_in13 = reg_0527;
    90: op1_03_in13 = imem03_in[47:44];
    91: op1_03_in13 = imem03_in[87:84];
    92: op1_03_in13 = reg_0654;
    93: op1_03_in13 = reg_0246;
    94: op1_03_in13 = reg_0038;
    95: op1_03_in13 = reg_0402;
    96: op1_03_in13 = reg_0516;
    default: op1_03_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv13 = 1;
    6: op1_03_inv13 = 1;
    3: op1_03_inv13 = 1;
    13: op1_03_inv13 = 1;
    14: op1_03_inv13 = 1;
    15: op1_03_inv13 = 1;
    16: op1_03_inv13 = 1;
    17: op1_03_inv13 = 1;
    18: op1_03_inv13 = 1;
    19: op1_03_inv13 = 1;
    21: op1_03_inv13 = 1;
    24: op1_03_inv13 = 1;
    25: op1_03_inv13 = 1;
    26: op1_03_inv13 = 1;
    29: op1_03_inv13 = 1;
    32: op1_03_inv13 = 1;
    33: op1_03_inv13 = 1;
    35: op1_03_inv13 = 1;
    41: op1_03_inv13 = 1;
    42: op1_03_inv13 = 1;
    43: op1_03_inv13 = 1;
    45: op1_03_inv13 = 1;
    51: op1_03_inv13 = 1;
    53: op1_03_inv13 = 1;
    56: op1_03_inv13 = 1;
    57: op1_03_inv13 = 1;
    58: op1_03_inv13 = 1;
    61: op1_03_inv13 = 1;
    62: op1_03_inv13 = 1;
    63: op1_03_inv13 = 1;
    67: op1_03_inv13 = 1;
    69: op1_03_inv13 = 1;
    70: op1_03_inv13 = 1;
    74: op1_03_inv13 = 1;
    75: op1_03_inv13 = 1;
    76: op1_03_inv13 = 1;
    81: op1_03_inv13 = 1;
    84: op1_03_inv13 = 1;
    85: op1_03_inv13 = 1;
    88: op1_03_inv13 = 1;
    89: op1_03_inv13 = 1;
    90: op1_03_inv13 = 1;
    91: op1_03_inv13 = 1;
    95: op1_03_inv13 = 1;
    default: op1_03_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in14 = reg_0485;
    5: op1_03_in14 = reg_0084;
    38: op1_03_in14 = reg_0084;
    6: op1_03_in14 = imem07_in[11:8];
    7: op1_03_in14 = reg_0097;
    8: op1_03_in14 = reg_0072;
    9: op1_03_in14 = imem05_in[51:48];
    3: op1_03_in14 = reg_0164;
    10: op1_03_in14 = imem06_in[19:16];
    11: op1_03_in14 = imem04_in[51:48];
    12: op1_03_in14 = imem06_in[111:108];
    13: op1_03_in14 = reg_0352;
    14: op1_03_in14 = reg_0547;
    15: op1_03_in14 = reg_0608;
    16: op1_03_in14 = imem01_in[3:0];
    17: op1_03_in14 = imem05_in[103:100];
    18: op1_03_in14 = reg_0648;
    19: op1_03_in14 = reg_0551;
    20: op1_03_in14 = imem01_in[107:104];
    21: op1_03_in14 = reg_0291;
    22: op1_03_in14 = reg_0154;
    23: op1_03_in14 = reg_0569;
    24: op1_03_in14 = reg_0036;
    25: op1_03_in14 = reg_0196;
    26: op1_03_in14 = reg_0403;
    27: op1_03_in14 = reg_0211;
    28: op1_03_in14 = reg_0077;
    29: op1_03_in14 = imem06_in[7:4];
    30: op1_03_in14 = reg_0190;
    31: op1_03_in14 = reg_0384;
    32: op1_03_in14 = reg_0790;
    33: op1_03_in14 = reg_0720;
    34: op1_03_in14 = reg_0075;
    35: op1_03_in14 = reg_0385;
    36: op1_03_in14 = reg_0492;
    37: op1_03_in14 = reg_0785;
    40: op1_03_in14 = reg_0819;
    41: op1_03_in14 = imem02_in[71:68];
    42: op1_03_in14 = imem04_in[63:60];
    43: op1_03_in14 = reg_0618;
    44: op1_03_in14 = reg_0473;
    45: op1_03_in14 = reg_0533;
    58: op1_03_in14 = reg_0533;
    46: op1_03_in14 = reg_0153;
    47: op1_03_in14 = reg_0614;
    48: op1_03_in14 = reg_0539;
    49: op1_03_in14 = reg_0115;
    50: op1_03_in14 = reg_0478;
    51: op1_03_in14 = imem07_in[75:72];
    53: op1_03_in14 = reg_0195;
    69: op1_03_in14 = reg_0195;
    54: op1_03_in14 = reg_0511;
    55: op1_03_in14 = reg_0666;
    56: op1_03_in14 = imem04_in[71:68];
    57: op1_03_in14 = imem04_in[31:28];
    59: op1_03_in14 = imem06_in[75:72];
    60: op1_03_in14 = reg_0617;
    61: op1_03_in14 = imem06_in[11:8];
    62: op1_03_in14 = reg_0462;
    63: op1_03_in14 = imem01_in[71:68];
    64: op1_03_in14 = reg_0483;
    65: op1_03_in14 = reg_0581;
    66: op1_03_in14 = reg_0661;
    67: op1_03_in14 = reg_0116;
    68: op1_03_in14 = reg_0169;
    70: op1_03_in14 = reg_0808;
    71: op1_03_in14 = reg_0193;
    72: op1_03_in14 = reg_0121;
    73: op1_03_in14 = reg_0541;
    74: op1_03_in14 = imem04_in[19:16];
    75: op1_03_in14 = reg_0593;
    76: op1_03_in14 = reg_0256;
    78: op1_03_in14 = reg_0548;
    79: op1_03_in14 = reg_0532;
    80: op1_03_in14 = reg_0556;
    96: op1_03_in14 = reg_0556;
    81: op1_03_in14 = reg_0799;
    83: op1_03_in14 = reg_0625;
    84: op1_03_in14 = reg_0342;
    85: op1_03_in14 = reg_0071;
    86: op1_03_in14 = reg_0214;
    87: op1_03_in14 = reg_0197;
    88: op1_03_in14 = reg_0771;
    89: op1_03_in14 = reg_0030;
    90: op1_03_in14 = imem03_in[71:68];
    91: op1_03_in14 = reg_0602;
    92: op1_03_in14 = reg_0763;
    93: op1_03_in14 = reg_0750;
    94: op1_03_in14 = reg_0654;
    95: op1_03_in14 = reg_0659;
    default: op1_03_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv14 = 1;
    6: op1_03_inv14 = 1;
    7: op1_03_inv14 = 1;
    8: op1_03_inv14 = 1;
    3: op1_03_inv14 = 1;
    12: op1_03_inv14 = 1;
    13: op1_03_inv14 = 1;
    14: op1_03_inv14 = 1;
    15: op1_03_inv14 = 1;
    16: op1_03_inv14 = 1;
    17: op1_03_inv14 = 1;
    20: op1_03_inv14 = 1;
    22: op1_03_inv14 = 1;
    26: op1_03_inv14 = 1;
    28: op1_03_inv14 = 1;
    30: op1_03_inv14 = 1;
    31: op1_03_inv14 = 1;
    34: op1_03_inv14 = 1;
    35: op1_03_inv14 = 1;
    37: op1_03_inv14 = 1;
    38: op1_03_inv14 = 1;
    41: op1_03_inv14 = 1;
    43: op1_03_inv14 = 1;
    46: op1_03_inv14 = 1;
    47: op1_03_inv14 = 1;
    49: op1_03_inv14 = 1;
    50: op1_03_inv14 = 1;
    51: op1_03_inv14 = 1;
    58: op1_03_inv14 = 1;
    63: op1_03_inv14 = 1;
    64: op1_03_inv14 = 1;
    66: op1_03_inv14 = 1;
    67: op1_03_inv14 = 1;
    69: op1_03_inv14 = 1;
    71: op1_03_inv14 = 1;
    74: op1_03_inv14 = 1;
    78: op1_03_inv14 = 1;
    79: op1_03_inv14 = 1;
    81: op1_03_inv14 = 1;
    85: op1_03_inv14 = 1;
    91: op1_03_inv14 = 1;
    95: op1_03_inv14 = 1;
    default: op1_03_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in15 = reg_0486;
    5: op1_03_in15 = reg_0093;
    6: op1_03_in15 = imem07_in[23:20];
    76: op1_03_in15 = imem07_in[23:20];
    7: op1_03_in15 = reg_0073;
    8: op1_03_in15 = imem05_in[19:16];
    9: op1_03_in15 = imem05_in[55:52];
    10: op1_03_in15 = imem06_in[43:40];
    11: op1_03_in15 = imem04_in[107:104];
    12: op1_03_in15 = reg_0606;
    13: op1_03_in15 = reg_0334;
    14: op1_03_in15 = reg_0281;
    15: op1_03_in15 = reg_0618;
    16: op1_03_in15 = imem01_in[11:8];
    17: op1_03_in15 = imem05_in[107:104];
    18: op1_03_in15 = reg_0638;
    19: op1_03_in15 = reg_0054;
    20: op1_03_in15 = reg_0523;
    21: op1_03_in15 = reg_0268;
    22: op1_03_in15 = reg_0139;
    23: op1_03_in15 = reg_0592;
    24: op1_03_in15 = reg_0037;
    25: op1_03_in15 = imem01_in[31:28];
    26: op1_03_in15 = reg_0390;
    27: op1_03_in15 = reg_0194;
    28: op1_03_in15 = reg_0072;
    29: op1_03_in15 = imem06_in[11:8];
    30: op1_03_in15 = reg_0199;
    31: op1_03_in15 = reg_0564;
    32: op1_03_in15 = reg_0304;
    33: op1_03_in15 = reg_0708;
    34: op1_03_in15 = reg_0070;
    35: op1_03_in15 = reg_0397;
    36: op1_03_in15 = reg_0780;
    60: op1_03_in15 = reg_0780;
    37: op1_03_in15 = reg_0783;
    38: op1_03_in15 = reg_0285;
    40: op1_03_in15 = reg_0814;
    47: op1_03_in15 = reg_0814;
    41: op1_03_in15 = reg_0657;
    42: op1_03_in15 = imem04_in[95:92];
    43: op1_03_in15 = reg_0622;
    44: op1_03_in15 = reg_0471;
    45: op1_03_in15 = reg_0095;
    46: op1_03_in15 = imem06_in[7:4];
    48: op1_03_in15 = imem03_in[15:12];
    49: op1_03_in15 = reg_0107;
    50: op1_03_in15 = reg_0214;
    51: op1_03_in15 = imem07_in[83:80];
    53: op1_03_in15 = reg_0192;
    54: op1_03_in15 = reg_0603;
    55: op1_03_in15 = reg_0637;
    56: op1_03_in15 = imem04_in[119:116];
    57: op1_03_in15 = imem04_in[43:40];
    58: op1_03_in15 = reg_0098;
    59: op1_03_in15 = imem06_in[83:80];
    61: op1_03_in15 = imem06_in[15:12];
    62: op1_03_in15 = reg_0456;
    63: op1_03_in15 = imem01_in[107:104];
    64: op1_03_in15 = reg_0345;
    65: op1_03_in15 = reg_0360;
    66: op1_03_in15 = reg_0483;
    67: op1_03_in15 = reg_0509;
    91: op1_03_in15 = reg_0509;
    68: op1_03_in15 = reg_0182;
    69: op1_03_in15 = imem01_in[63:60];
    70: op1_03_in15 = reg_0015;
    71: op1_03_in15 = reg_0198;
    72: op1_03_in15 = imem02_in[19:16];
    73: op1_03_in15 = reg_0530;
    74: op1_03_in15 = imem04_in[59:56];
    75: op1_03_in15 = reg_0663;
    78: op1_03_in15 = reg_0426;
    79: op1_03_in15 = imem03_in[11:8];
    80: op1_03_in15 = reg_0432;
    81: op1_03_in15 = reg_0016;
    83: op1_03_in15 = reg_0291;
    84: op1_03_in15 = imem02_in[35:32];
    85: op1_03_in15 = reg_0617;
    86: op1_03_in15 = reg_0200;
    87: op1_03_in15 = imem01_in[75:72];
    88: op1_03_in15 = imem05_in[3:0];
    89: op1_03_in15 = reg_0743;
    90: op1_03_in15 = imem03_in[87:84];
    92: op1_03_in15 = reg_0215;
    93: op1_03_in15 = reg_0608;
    94: op1_03_in15 = reg_0750;
    95: op1_03_in15 = reg_0512;
    96: op1_03_in15 = reg_0305;
    default: op1_03_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv15 = 1;
    10: op1_03_inv15 = 1;
    12: op1_03_inv15 = 1;
    13: op1_03_inv15 = 1;
    17: op1_03_inv15 = 1;
    18: op1_03_inv15 = 1;
    20: op1_03_inv15 = 1;
    22: op1_03_inv15 = 1;
    23: op1_03_inv15 = 1;
    24: op1_03_inv15 = 1;
    26: op1_03_inv15 = 1;
    27: op1_03_inv15 = 1;
    28: op1_03_inv15 = 1;
    29: op1_03_inv15 = 1;
    30: op1_03_inv15 = 1;
    34: op1_03_inv15 = 1;
    36: op1_03_inv15 = 1;
    37: op1_03_inv15 = 1;
    40: op1_03_inv15 = 1;
    42: op1_03_inv15 = 1;
    43: op1_03_inv15 = 1;
    46: op1_03_inv15 = 1;
    47: op1_03_inv15 = 1;
    54: op1_03_inv15 = 1;
    55: op1_03_inv15 = 1;
    57: op1_03_inv15 = 1;
    63: op1_03_inv15 = 1;
    64: op1_03_inv15 = 1;
    65: op1_03_inv15 = 1;
    67: op1_03_inv15 = 1;
    70: op1_03_inv15 = 1;
    71: op1_03_inv15 = 1;
    72: op1_03_inv15 = 1;
    73: op1_03_inv15 = 1;
    74: op1_03_inv15 = 1;
    75: op1_03_inv15 = 1;
    76: op1_03_inv15 = 1;
    78: op1_03_inv15 = 1;
    79: op1_03_inv15 = 1;
    84: op1_03_inv15 = 1;
    88: op1_03_inv15 = 1;
    92: op1_03_inv15 = 1;
    96: op1_03_inv15 = 1;
    default: op1_03_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in16 = reg_0259;
    5: op1_03_in16 = reg_0740;
    6: op1_03_in16 = imem07_in[47:44];
    7: op1_03_in16 = imem03_in[115:112];
    8: op1_03_in16 = imem05_in[63:60];
    9: op1_03_in16 = imem05_in[63:60];
    10: op1_03_in16 = imem06_in[87:84];
    11: op1_03_in16 = reg_0545;
    12: op1_03_in16 = reg_0619;
    13: op1_03_in16 = reg_0341;
    14: op1_03_in16 = reg_0285;
    15: op1_03_in16 = reg_0622;
    16: op1_03_in16 = imem01_in[47:44];
    53: op1_03_in16 = imem01_in[47:44];
    17: op1_03_in16 = imem05_in[111:108];
    18: op1_03_in16 = reg_0644;
    41: op1_03_in16 = reg_0644;
    19: op1_03_in16 = reg_0298;
    20: op1_03_in16 = reg_0522;
    21: op1_03_in16 = reg_0061;
    22: op1_03_in16 = reg_0138;
    23: op1_03_in16 = reg_0585;
    24: op1_03_in16 = reg_0750;
    25: op1_03_in16 = imem01_in[63:60];
    26: op1_03_in16 = reg_0380;
    27: op1_03_in16 = reg_0206;
    28: op1_03_in16 = imem05_in[39:36];
    29: op1_03_in16 = imem06_in[35:32];
    30: op1_03_in16 = imem01_in[7:4];
    31: op1_03_in16 = reg_0392;
    32: op1_03_in16 = reg_0309;
    33: op1_03_in16 = reg_0709;
    34: op1_03_in16 = imem05_in[15:12];
    35: op1_03_in16 = reg_0747;
    36: op1_03_in16 = reg_0787;
    37: op1_03_in16 = reg_0786;
    38: op1_03_in16 = reg_0145;
    40: op1_03_in16 = imem07_in[23:20];
    42: op1_03_in16 = reg_0316;
    43: op1_03_in16 = reg_0278;
    44: op1_03_in16 = reg_0479;
    45: op1_03_in16 = reg_0770;
    46: op1_03_in16 = reg_0289;
    47: op1_03_in16 = imem07_in[11:8];
    75: op1_03_in16 = imem07_in[11:8];
    48: op1_03_in16 = imem03_in[39:36];
    49: op1_03_in16 = reg_0126;
    50: op1_03_in16 = reg_0209;
    86: op1_03_in16 = reg_0209;
    51: op1_03_in16 = imem07_in[91:88];
    54: op1_03_in16 = reg_0234;
    55: op1_03_in16 = reg_0638;
    56: op1_03_in16 = imem04_in[127:124];
    57: op1_03_in16 = imem04_in[83:80];
    58: op1_03_in16 = imem03_in[3:0];
    59: op1_03_in16 = reg_0115;
    60: op1_03_in16 = reg_0774;
    61: op1_03_in16 = imem06_in[71:68];
    62: op1_03_in16 = reg_0210;
    63: op1_03_in16 = reg_0085;
    64: op1_03_in16 = reg_0324;
    65: op1_03_in16 = reg_0324;
    66: op1_03_in16 = reg_0647;
    67: op1_03_in16 = reg_0755;
    68: op1_03_in16 = reg_0185;
    69: op1_03_in16 = imem01_in[83:80];
    70: op1_03_in16 = reg_0806;
    71: op1_03_in16 = imem01_in[51:48];
    72: op1_03_in16 = imem02_in[55:52];
    73: op1_03_in16 = reg_0535;
    74: op1_03_in16 = imem04_in[99:96];
    76: op1_03_in16 = imem07_in[95:92];
    78: op1_03_in16 = reg_0358;
    79: op1_03_in16 = imem03_in[35:32];
    80: op1_03_in16 = reg_0283;
    81: op1_03_in16 = imem04_in[35:32];
    83: op1_03_in16 = reg_0370;
    84: op1_03_in16 = imem02_in[51:48];
    85: op1_03_in16 = reg_0687;
    87: op1_03_in16 = imem01_in[79:76];
    88: op1_03_in16 = imem05_in[79:76];
    89: op1_03_in16 = reg_0132;
    90: op1_03_in16 = imem03_in[91:88];
    91: op1_03_in16 = reg_0559;
    92: op1_03_in16 = reg_0515;
    93: op1_03_in16 = reg_0242;
    94: op1_03_in16 = reg_0242;
    95: op1_03_in16 = reg_0663;
    96: op1_03_in16 = reg_0071;
    default: op1_03_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv16 = 1;
    5: op1_03_inv16 = 1;
    10: op1_03_inv16 = 1;
    11: op1_03_inv16 = 1;
    14: op1_03_inv16 = 1;
    19: op1_03_inv16 = 1;
    22: op1_03_inv16 = 1;
    23: op1_03_inv16 = 1;
    24: op1_03_inv16 = 1;
    26: op1_03_inv16 = 1;
    28: op1_03_inv16 = 1;
    31: op1_03_inv16 = 1;
    32: op1_03_inv16 = 1;
    34: op1_03_inv16 = 1;
    38: op1_03_inv16 = 1;
    40: op1_03_inv16 = 1;
    42: op1_03_inv16 = 1;
    43: op1_03_inv16 = 1;
    44: op1_03_inv16 = 1;
    47: op1_03_inv16 = 1;
    48: op1_03_inv16 = 1;
    53: op1_03_inv16 = 1;
    54: op1_03_inv16 = 1;
    55: op1_03_inv16 = 1;
    57: op1_03_inv16 = 1;
    60: op1_03_inv16 = 1;
    64: op1_03_inv16 = 1;
    66: op1_03_inv16 = 1;
    67: op1_03_inv16 = 1;
    68: op1_03_inv16 = 1;
    75: op1_03_inv16 = 1;
    76: op1_03_inv16 = 1;
    80: op1_03_inv16 = 1;
    85: op1_03_inv16 = 1;
    86: op1_03_inv16 = 1;
    87: op1_03_inv16 = 1;
    88: op1_03_inv16 = 1;
    91: op1_03_inv16 = 1;
    95: op1_03_inv16 = 1;
    96: op1_03_inv16 = 1;
    default: op1_03_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in17 = reg_0260;
    5: op1_03_in17 = reg_0568;
    6: op1_03_in17 = imem07_in[51:48];
    7: op1_03_in17 = reg_0573;
    8: op1_03_in17 = imem05_in[67:64];
    9: op1_03_in17 = imem05_in[75:72];
    10: op1_03_in17 = imem06_in[103:100];
    11: op1_03_in17 = reg_0550;
    12: op1_03_in17 = reg_0615;
    13: op1_03_in17 = reg_0330;
    14: op1_03_in17 = reg_0286;
    15: op1_03_in17 = reg_0407;
    16: op1_03_in17 = imem01_in[51:48];
    17: op1_03_in17 = imem05_in[119:116];
    18: op1_03_in17 = reg_0643;
    19: op1_03_in17 = reg_0266;
    20: op1_03_in17 = reg_0520;
    21: op1_03_in17 = reg_0281;
    22: op1_03_in17 = reg_0153;
    38: op1_03_in17 = reg_0153;
    23: op1_03_in17 = reg_0600;
    24: op1_03_in17 = reg_0029;
    25: op1_03_in17 = imem01_in[95:92];
    87: op1_03_in17 = imem01_in[95:92];
    26: op1_03_in17 = reg_0028;
    27: op1_03_in17 = reg_0197;
    28: op1_03_in17 = imem05_in[63:60];
    29: op1_03_in17 = imem06_in[95:92];
    30: op1_03_in17 = imem01_in[39:36];
    31: op1_03_in17 = reg_0376;
    32: op1_03_in17 = reg_0735;
    33: op1_03_in17 = reg_0718;
    34: op1_03_in17 = imem05_in[59:56];
    35: op1_03_in17 = reg_0003;
    36: op1_03_in17 = reg_0489;
    37: op1_03_in17 = reg_0787;
    40: op1_03_in17 = imem07_in[27:24];
    41: op1_03_in17 = reg_0652;
    42: op1_03_in17 = reg_0560;
    43: op1_03_in17 = reg_0778;
    44: op1_03_in17 = reg_0456;
    45: op1_03_in17 = reg_0093;
    46: op1_03_in17 = reg_0291;
    47: op1_03_in17 = imem07_in[59:56];
    48: op1_03_in17 = imem03_in[47:44];
    49: op1_03_in17 = imem02_in[51:48];
    50: op1_03_in17 = reg_0207;
    51: op1_03_in17 = imem07_in[95:92];
    53: op1_03_in17 = imem01_in[79:76];
    54: op1_03_in17 = reg_0504;
    55: op1_03_in17 = reg_0417;
    56: op1_03_in17 = reg_0059;
    57: op1_03_in17 = reg_0087;
    58: op1_03_in17 = imem03_in[19:16];
    59: op1_03_in17 = reg_0577;
    60: op1_03_in17 = reg_0233;
    61: op1_03_in17 = imem06_in[91:88];
    62: op1_03_in17 = reg_0189;
    63: op1_03_in17 = reg_0100;
    64: op1_03_in17 = reg_0518;
    65: op1_03_in17 = reg_0566;
    66: op1_03_in17 = reg_0753;
    67: op1_03_in17 = reg_0002;
    69: op1_03_in17 = imem01_in[87:84];
    71: op1_03_in17 = imem01_in[87:84];
    70: op1_03_in17 = imem04_in[43:40];
    72: op1_03_in17 = imem02_in[59:56];
    73: op1_03_in17 = reg_0098;
    74: op1_03_in17 = reg_0088;
    75: op1_03_in17 = imem07_in[19:16];
    76: op1_03_in17 = imem07_in[123:120];
    78: op1_03_in17 = reg_0364;
    79: op1_03_in17 = imem03_in[83:80];
    80: op1_03_in17 = reg_0529;
    81: op1_03_in17 = imem04_in[51:48];
    83: op1_03_in17 = reg_0619;
    84: op1_03_in17 = imem02_in[75:72];
    85: op1_03_in17 = reg_0068;
    86: op1_03_in17 = reg_0193;
    88: op1_03_in17 = imem05_in[115:112];
    89: op1_03_in17 = reg_0584;
    90: op1_03_in17 = imem03_in[103:100];
    91: op1_03_in17 = reg_0389;
    92: op1_03_in17 = reg_0655;
    93: op1_03_in17 = reg_0661;
    94: op1_03_in17 = reg_0576;
    95: op1_03_in17 = reg_0612;
    96: op1_03_in17 = reg_0629;
    default: op1_03_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv17 = 1;
    6: op1_03_inv17 = 1;
    7: op1_03_inv17 = 1;
    8: op1_03_inv17 = 1;
    10: op1_03_inv17 = 1;
    11: op1_03_inv17 = 1;
    12: op1_03_inv17 = 1;
    13: op1_03_inv17 = 1;
    15: op1_03_inv17 = 1;
    16: op1_03_inv17 = 1;
    18: op1_03_inv17 = 1;
    23: op1_03_inv17 = 1;
    24: op1_03_inv17 = 1;
    25: op1_03_inv17 = 1;
    26: op1_03_inv17 = 1;
    28: op1_03_inv17 = 1;
    29: op1_03_inv17 = 1;
    31: op1_03_inv17 = 1;
    32: op1_03_inv17 = 1;
    35: op1_03_inv17 = 1;
    36: op1_03_inv17 = 1;
    37: op1_03_inv17 = 1;
    40: op1_03_inv17 = 1;
    41: op1_03_inv17 = 1;
    46: op1_03_inv17 = 1;
    50: op1_03_inv17 = 1;
    51: op1_03_inv17 = 1;
    53: op1_03_inv17 = 1;
    54: op1_03_inv17 = 1;
    55: op1_03_inv17 = 1;
    57: op1_03_inv17 = 1;
    58: op1_03_inv17 = 1;
    59: op1_03_inv17 = 1;
    62: op1_03_inv17 = 1;
    69: op1_03_inv17 = 1;
    71: op1_03_inv17 = 1;
    72: op1_03_inv17 = 1;
    73: op1_03_inv17 = 1;
    75: op1_03_inv17 = 1;
    76: op1_03_inv17 = 1;
    79: op1_03_inv17 = 1;
    80: op1_03_inv17 = 1;
    84: op1_03_inv17 = 1;
    86: op1_03_inv17 = 1;
    87: op1_03_inv17 = 1;
    88: op1_03_inv17 = 1;
    89: op1_03_inv17 = 1;
    91: op1_03_inv17 = 1;
    92: op1_03_inv17 = 1;
    93: op1_03_inv17 = 1;
    94: op1_03_inv17 = 1;
    default: op1_03_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in18 = reg_0132;
    5: op1_03_in18 = reg_0589;
    6: op1_03_in18 = imem07_in[67:64];
    7: op1_03_in18 = reg_0579;
    8: op1_03_in18 = imem05_in[75:72];
    34: op1_03_in18 = imem05_in[75:72];
    9: op1_03_in18 = imem05_in[83:80];
    10: op1_03_in18 = reg_0614;
    11: op1_03_in18 = reg_0529;
    12: op1_03_in18 = reg_0379;
    13: op1_03_in18 = reg_0324;
    14: op1_03_in18 = reg_0307;
    15: op1_03_in18 = reg_0371;
    16: op1_03_in18 = imem01_in[67:64];
    17: op1_03_in18 = reg_0789;
    18: op1_03_in18 = reg_0652;
    19: op1_03_in18 = reg_0284;
    20: op1_03_in18 = reg_0778;
    21: op1_03_in18 = reg_0253;
    22: op1_03_in18 = reg_0144;
    23: op1_03_in18 = reg_0597;
    24: op1_03_in18 = imem07_in[23:20];
    75: op1_03_in18 = imem07_in[23:20];
    25: op1_03_in18 = imem01_in[103:100];
    26: op1_03_in18 = reg_0815;
    27: op1_03_in18 = imem01_in[15:12];
    28: op1_03_in18 = imem05_in[91:88];
    29: op1_03_in18 = reg_0628;
    30: op1_03_in18 = imem01_in[55:52];
    31: op1_03_in18 = reg_0499;
    32: op1_03_in18 = reg_0147;
    33: op1_03_in18 = reg_0422;
    35: op1_03_in18 = reg_0008;
    36: op1_03_in18 = reg_0736;
    88: op1_03_in18 = reg_0736;
    37: op1_03_in18 = reg_0486;
    38: op1_03_in18 = reg_0140;
    40: op1_03_in18 = imem07_in[55:52];
    41: op1_03_in18 = reg_0349;
    42: op1_03_in18 = reg_0043;
    43: op1_03_in18 = reg_0620;
    44: op1_03_in18 = reg_0214;
    45: op1_03_in18 = imem03_in[3:0];
    46: op1_03_in18 = reg_0624;
    47: op1_03_in18 = imem07_in[87:84];
    48: op1_03_in18 = imem03_in[59:56];
    49: op1_03_in18 = imem02_in[67:64];
    50: op1_03_in18 = reg_0211;
    51: op1_03_in18 = imem07_in[111:108];
    53: op1_03_in18 = reg_0497;
    54: op1_03_in18 = reg_0118;
    55: op1_03_in18 = reg_0426;
    56: op1_03_in18 = reg_0316;
    57: op1_03_in18 = reg_0060;
    58: op1_03_in18 = imem03_in[43:40];
    59: op1_03_in18 = reg_0038;
    60: op1_03_in18 = imem05_in[7:4];
    61: op1_03_in18 = imem06_in[107:104];
    62: op1_03_in18 = reg_0201;
    63: op1_03_in18 = reg_0321;
    64: op1_03_in18 = reg_0092;
    65: op1_03_in18 = reg_0097;
    66: op1_03_in18 = reg_0417;
    67: op1_03_in18 = reg_0003;
    69: op1_03_in18 = reg_0385;
    70: op1_03_in18 = imem04_in[103:100];
    71: op1_03_in18 = imem01_in[95:92];
    72: op1_03_in18 = imem02_in[107:104];
    73: op1_03_in18 = imem03_in[67:64];
    74: op1_03_in18 = reg_0554;
    76: op1_03_in18 = imem07_in[127:124];
    78: op1_03_in18 = reg_0345;
    79: op1_03_in18 = imem03_in[99:96];
    80: op1_03_in18 = reg_0071;
    81: op1_03_in18 = imem04_in[83:80];
    83: op1_03_in18 = reg_0618;
    84: op1_03_in18 = imem02_in[111:108];
    85: op1_03_in18 = reg_0780;
    86: op1_03_in18 = reg_0192;
    87: op1_03_in18 = imem01_in[119:116];
    89: op1_03_in18 = reg_0136;
    90: op1_03_in18 = reg_0507;
    91: op1_03_in18 = reg_0572;
    92: op1_03_in18 = reg_0651;
    93: op1_03_in18 = imem07_in[39:36];
    94: op1_03_in18 = reg_0612;
    95: op1_03_in18 = reg_0351;
    96: op1_03_in18 = reg_0627;
    default: op1_03_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv18 = 1;
    5: op1_03_inv18 = 1;
    6: op1_03_inv18 = 1;
    7: op1_03_inv18 = 1;
    10: op1_03_inv18 = 1;
    11: op1_03_inv18 = 1;
    13: op1_03_inv18 = 1;
    14: op1_03_inv18 = 1;
    17: op1_03_inv18 = 1;
    19: op1_03_inv18 = 1;
    20: op1_03_inv18 = 1;
    21: op1_03_inv18 = 1;
    23: op1_03_inv18 = 1;
    27: op1_03_inv18 = 1;
    28: op1_03_inv18 = 1;
    29: op1_03_inv18 = 1;
    30: op1_03_inv18 = 1;
    32: op1_03_inv18 = 1;
    33: op1_03_inv18 = 1;
    34: op1_03_inv18 = 1;
    35: op1_03_inv18 = 1;
    36: op1_03_inv18 = 1;
    38: op1_03_inv18 = 1;
    42: op1_03_inv18 = 1;
    46: op1_03_inv18 = 1;
    48: op1_03_inv18 = 1;
    53: op1_03_inv18 = 1;
    55: op1_03_inv18 = 1;
    56: op1_03_inv18 = 1;
    57: op1_03_inv18 = 1;
    58: op1_03_inv18 = 1;
    60: op1_03_inv18 = 1;
    64: op1_03_inv18 = 1;
    67: op1_03_inv18 = 1;
    69: op1_03_inv18 = 1;
    72: op1_03_inv18 = 1;
    73: op1_03_inv18 = 1;
    75: op1_03_inv18 = 1;
    78: op1_03_inv18 = 1;
    80: op1_03_inv18 = 1;
    81: op1_03_inv18 = 1;
    83: op1_03_inv18 = 1;
    84: op1_03_inv18 = 1;
    87: op1_03_inv18 = 1;
    89: op1_03_inv18 = 1;
    90: op1_03_inv18 = 1;
    91: op1_03_inv18 = 1;
    92: op1_03_inv18 = 1;
    93: op1_03_inv18 = 1;
    default: op1_03_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in19 = reg_0136;
    5: op1_03_in19 = reg_0580;
    6: op1_03_in19 = imem07_in[71:68];
    7: op1_03_in19 = reg_0597;
    8: op1_03_in19 = imem05_in[91:88];
    9: op1_03_in19 = imem05_in[119:116];
    10: op1_03_in19 = reg_0604;
    11: op1_03_in19 = reg_0556;
    12: op1_03_in19 = reg_0390;
    13: op1_03_in19 = reg_0365;
    14: op1_03_in19 = reg_0061;
    19: op1_03_in19 = reg_0061;
    15: op1_03_in19 = reg_0382;
    16: op1_03_in19 = imem01_in[119:116];
    17: op1_03_in19 = reg_0780;
    18: op1_03_in19 = reg_0357;
    20: op1_03_in19 = reg_0515;
    21: op1_03_in19 = reg_0068;
    22: op1_03_in19 = imem06_in[15:12];
    23: op1_03_in19 = reg_0391;
    24: op1_03_in19 = imem07_in[31:28];
    25: op1_03_in19 = reg_0761;
    26: op1_03_in19 = reg_0749;
    27: op1_03_in19 = imem01_in[31:28];
    28: op1_03_in19 = reg_0788;
    29: op1_03_in19 = reg_0621;
    72: op1_03_in19 = reg_0621;
    30: op1_03_in19 = imem01_in[87:84];
    31: op1_03_in19 = reg_0374;
    32: op1_03_in19 = reg_0139;
    33: op1_03_in19 = reg_0421;
    34: op1_03_in19 = imem05_in[99:96];
    35: op1_03_in19 = imem04_in[11:8];
    36: op1_03_in19 = reg_0741;
    37: op1_03_in19 = reg_0090;
    38: op1_03_in19 = reg_0155;
    40: op1_03_in19 = imem07_in[59:56];
    93: op1_03_in19 = imem07_in[59:56];
    41: op1_03_in19 = reg_0359;
    42: op1_03_in19 = reg_0555;
    43: op1_03_in19 = reg_0037;
    44: op1_03_in19 = reg_0189;
    45: op1_03_in19 = imem03_in[71:68];
    46: op1_03_in19 = reg_0613;
    47: op1_03_in19 = imem07_in[115:112];
    48: op1_03_in19 = imem03_in[127:124];
    49: op1_03_in19 = imem02_in[119:116];
    50: op1_03_in19 = reg_0192;
    51: op1_03_in19 = reg_0722;
    76: op1_03_in19 = reg_0722;
    53: op1_03_in19 = reg_0496;
    54: op1_03_in19 = reg_0106;
    55: op1_03_in19 = reg_0485;
    56: op1_03_in19 = reg_0553;
    57: op1_03_in19 = reg_0308;
    58: op1_03_in19 = imem03_in[95:92];
    59: op1_03_in19 = reg_0260;
    60: op1_03_in19 = imem05_in[23:20];
    61: op1_03_in19 = reg_0346;
    62: op1_03_in19 = reg_0213;
    63: op1_03_in19 = reg_0225;
    64: op1_03_in19 = reg_0770;
    65: op1_03_in19 = reg_0535;
    66: op1_03_in19 = reg_0587;
    67: op1_03_in19 = reg_0807;
    69: op1_03_in19 = reg_0131;
    70: op1_03_in19 = imem04_in[111:108];
    71: op1_03_in19 = imem01_in[99:96];
    73: op1_03_in19 = imem03_in[91:88];
    74: op1_03_in19 = reg_0631;
    75: op1_03_in19 = imem07_in[39:36];
    78: op1_03_in19 = reg_0356;
    79: op1_03_in19 = imem03_in[111:108];
    80: op1_03_in19 = reg_0050;
    81: op1_03_in19 = imem04_in[103:100];
    83: op1_03_in19 = reg_0766;
    84: op1_03_in19 = imem03_in[7:4];
    85: op1_03_in19 = reg_0311;
    86: op1_03_in19 = imem01_in[35:32];
    87: op1_03_in19 = imem01_in[127:124];
    88: op1_03_in19 = reg_0135;
    89: op1_03_in19 = reg_0703;
    90: op1_03_in19 = reg_0755;
    91: op1_03_in19 = reg_0571;
    92: op1_03_in19 = reg_0681;
    94: op1_03_in19 = reg_0620;
    95: op1_03_in19 = reg_0501;
    96: op1_03_in19 = reg_0078;
    default: op1_03_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_03_inv19 = 1;
    8: op1_03_inv19 = 1;
    13: op1_03_inv19 = 1;
    15: op1_03_inv19 = 1;
    17: op1_03_inv19 = 1;
    18: op1_03_inv19 = 1;
    19: op1_03_inv19 = 1;
    20: op1_03_inv19 = 1;
    23: op1_03_inv19 = 1;
    25: op1_03_inv19 = 1;
    30: op1_03_inv19 = 1;
    32: op1_03_inv19 = 1;
    34: op1_03_inv19 = 1;
    36: op1_03_inv19 = 1;
    40: op1_03_inv19 = 1;
    41: op1_03_inv19 = 1;
    43: op1_03_inv19 = 1;
    44: op1_03_inv19 = 1;
    45: op1_03_inv19 = 1;
    46: op1_03_inv19 = 1;
    50: op1_03_inv19 = 1;
    51: op1_03_inv19 = 1;
    54: op1_03_inv19 = 1;
    56: op1_03_inv19 = 1;
    59: op1_03_inv19 = 1;
    63: op1_03_inv19 = 1;
    64: op1_03_inv19 = 1;
    74: op1_03_inv19 = 1;
    80: op1_03_inv19 = 1;
    81: op1_03_inv19 = 1;
    83: op1_03_inv19 = 1;
    84: op1_03_inv19 = 1;
    88: op1_03_inv19 = 1;
    89: op1_03_inv19 = 1;
    90: op1_03_inv19 = 1;
    92: op1_03_inv19 = 1;
    94: op1_03_inv19 = 1;
    95: op1_03_inv19 = 1;
    96: op1_03_inv19 = 1;
    default: op1_03_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in20 = reg_0137;
    5: op1_03_in20 = reg_0590;
    7: op1_03_in20 = reg_0590;
    6: op1_03_in20 = imem07_in[79:76];
    8: op1_03_in20 = reg_0798;
    9: op1_03_in20 = reg_0798;
    10: op1_03_in20 = reg_0607;
    11: op1_03_in20 = reg_0308;
    12: op1_03_in20 = reg_0035;
    13: op1_03_in20 = reg_0336;
    14: op1_03_in20 = reg_0062;
    15: op1_03_in20 = reg_0368;
    16: op1_03_in20 = imem01_in[127:124];
    17: op1_03_in20 = reg_0783;
    18: op1_03_in20 = reg_0341;
    19: op1_03_in20 = reg_0079;
    20: op1_03_in20 = reg_0525;
    21: op1_03_in20 = reg_0064;
    22: op1_03_in20 = imem06_in[91:88];
    23: op1_03_in20 = reg_0360;
    78: op1_03_in20 = reg_0360;
    24: op1_03_in20 = imem07_in[39:36];
    25: op1_03_in20 = reg_0217;
    26: op1_03_in20 = imem07_in[35:32];
    27: op1_03_in20 = imem01_in[39:36];
    86: op1_03_in20 = imem01_in[39:36];
    28: op1_03_in20 = reg_0491;
    29: op1_03_in20 = reg_0626;
    30: op1_03_in20 = imem01_in[111:108];
    31: op1_03_in20 = reg_0001;
    32: op1_03_in20 = reg_0131;
    33: op1_03_in20 = reg_0426;
    34: op1_03_in20 = imem05_in[119:116];
    35: op1_03_in20 = imem04_in[39:36];
    36: op1_03_in20 = reg_0304;
    37: op1_03_in20 = reg_0304;
    38: op1_03_in20 = imem06_in[79:76];
    40: op1_03_in20 = reg_0703;
    72: op1_03_in20 = reg_0703;
    41: op1_03_in20 = reg_0323;
    42: op1_03_in20 = reg_0523;
    43: op1_03_in20 = reg_0632;
    44: op1_03_in20 = reg_0203;
    45: op1_03_in20 = imem03_in[99:96];
    46: op1_03_in20 = reg_0608;
    47: op1_03_in20 = reg_0726;
    48: op1_03_in20 = reg_0591;
    49: op1_03_in20 = reg_0650;
    50: op1_03_in20 = imem01_in[47:44];
    51: op1_03_in20 = reg_0731;
    76: op1_03_in20 = reg_0731;
    53: op1_03_in20 = reg_0765;
    54: op1_03_in20 = reg_0601;
    55: op1_03_in20 = reg_0363;
    56: op1_03_in20 = reg_0056;
    57: op1_03_in20 = reg_0615;
    58: op1_03_in20 = imem03_in[103:100];
    59: op1_03_in20 = reg_0519;
    60: op1_03_in20 = imem05_in[31:28];
    61: op1_03_in20 = reg_0815;
    62: op1_03_in20 = reg_0206;
    63: op1_03_in20 = reg_0418;
    64: op1_03_in20 = imem03_in[11:8];
    65: op1_03_in20 = reg_0756;
    66: op1_03_in20 = reg_0320;
    67: op1_03_in20 = reg_0014;
    69: op1_03_in20 = reg_0237;
    70: op1_03_in20 = reg_0262;
    71: op1_03_in20 = imem01_in[119:116];
    73: op1_03_in20 = imem03_in[95:92];
    74: op1_03_in20 = reg_0292;
    75: op1_03_in20 = imem07_in[47:44];
    79: op1_03_in20 = imem03_in[119:116];
    80: op1_03_in20 = reg_0622;
    81: op1_03_in20 = imem04_in[119:116];
    83: op1_03_in20 = reg_0260;
    84: op1_03_in20 = imem03_in[19:16];
    85: op1_03_in20 = reg_0371;
    87: op1_03_in20 = reg_0111;
    88: op1_03_in20 = reg_0227;
    89: op1_03_in20 = reg_0803;
    90: op1_03_in20 = reg_0646;
    91: op1_03_in20 = reg_0321;
    92: op1_03_in20 = reg_0612;
    93: op1_03_in20 = imem07_in[83:80];
    94: op1_03_in20 = reg_0609;
    95: op1_03_in20 = reg_0037;
    96: op1_03_in20 = reg_0065;
    default: op1_03_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv20 = 1;
    5: op1_03_inv20 = 1;
    6: op1_03_inv20 = 1;
    7: op1_03_inv20 = 1;
    9: op1_03_inv20 = 1;
    12: op1_03_inv20 = 1;
    13: op1_03_inv20 = 1;
    14: op1_03_inv20 = 1;
    16: op1_03_inv20 = 1;
    18: op1_03_inv20 = 1;
    20: op1_03_inv20 = 1;
    22: op1_03_inv20 = 1;
    23: op1_03_inv20 = 1;
    24: op1_03_inv20 = 1;
    25: op1_03_inv20 = 1;
    29: op1_03_inv20 = 1;
    35: op1_03_inv20 = 1;
    36: op1_03_inv20 = 1;
    40: op1_03_inv20 = 1;
    41: op1_03_inv20 = 1;
    42: op1_03_inv20 = 1;
    44: op1_03_inv20 = 1;
    46: op1_03_inv20 = 1;
    47: op1_03_inv20 = 1;
    50: op1_03_inv20 = 1;
    54: op1_03_inv20 = 1;
    55: op1_03_inv20 = 1;
    56: op1_03_inv20 = 1;
    57: op1_03_inv20 = 1;
    58: op1_03_inv20 = 1;
    62: op1_03_inv20 = 1;
    63: op1_03_inv20 = 1;
    64: op1_03_inv20 = 1;
    65: op1_03_inv20 = 1;
    70: op1_03_inv20 = 1;
    74: op1_03_inv20 = 1;
    79: op1_03_inv20 = 1;
    80: op1_03_inv20 = 1;
    84: op1_03_inv20 = 1;
    89: op1_03_inv20 = 1;
    91: op1_03_inv20 = 1;
    92: op1_03_inv20 = 1;
    95: op1_03_inv20 = 1;
    default: op1_03_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in21 = reg_0144;
    5: op1_03_in21 = reg_0387;
    6: op1_03_in21 = reg_0719;
    7: op1_03_in21 = reg_0360;
    8: op1_03_in21 = reg_0781;
    9: op1_03_in21 = reg_0796;
    10: op1_03_in21 = reg_0624;
    11: op1_03_in21 = reg_0301;
    12: op1_03_in21 = reg_0040;
    13: op1_03_in21 = reg_0081;
    14: op1_03_in21 = reg_0065;
    15: op1_03_in21 = reg_0033;
    16: op1_03_in21 = reg_0497;
    30: op1_03_in21 = reg_0497;
    17: op1_03_in21 = reg_0486;
    18: op1_03_in21 = reg_0359;
    19: op1_03_in21 = reg_0064;
    20: op1_03_in21 = reg_0516;
    21: op1_03_in21 = imem05_in[3:0];
    22: op1_03_in21 = reg_0625;
    23: op1_03_in21 = reg_0369;
    59: op1_03_in21 = reg_0369;
    24: op1_03_in21 = imem07_in[87:84];
    26: op1_03_in21 = imem07_in[87:84];
    93: op1_03_in21 = imem07_in[87:84];
    25: op1_03_in21 = reg_0504;
    27: op1_03_in21 = imem01_in[67:64];
    28: op1_03_in21 = reg_0794;
    29: op1_03_in21 = reg_0601;
    31: op1_03_in21 = reg_0003;
    32: op1_03_in21 = imem06_in[39:36];
    33: op1_03_in21 = reg_0434;
    34: op1_03_in21 = reg_0780;
    35: op1_03_in21 = imem04_in[51:48];
    36: op1_03_in21 = reg_0279;
    37: op1_03_in21 = reg_0226;
    38: op1_03_in21 = imem06_in[119:116];
    40: op1_03_in21 = reg_0712;
    41: op1_03_in21 = reg_0092;
    42: op1_03_in21 = reg_0547;
    43: op1_03_in21 = imem07_in[3:0];
    44: op1_03_in21 = reg_0186;
    45: op1_03_in21 = reg_0579;
    46: op1_03_in21 = reg_0766;
    47: op1_03_in21 = reg_0714;
    48: op1_03_in21 = reg_0573;
    49: op1_03_in21 = reg_0654;
    50: op1_03_in21 = imem01_in[99:96];
    51: op1_03_in21 = reg_0726;
    53: op1_03_in21 = reg_0778;
    54: op1_03_in21 = reg_0674;
    55: op1_03_in21 = reg_0406;
    56: op1_03_in21 = reg_0057;
    57: op1_03_in21 = reg_0050;
    58: op1_03_in21 = imem03_in[107:104];
    73: op1_03_in21 = imem03_in[107:104];
    60: op1_03_in21 = imem05_in[55:52];
    61: op1_03_in21 = reg_0404;
    62: op1_03_in21 = imem01_in[31:28];
    63: op1_03_in21 = reg_0306;
    64: op1_03_in21 = imem03_in[43:40];
    65: op1_03_in21 = reg_0094;
    66: op1_03_in21 = reg_0586;
    67: op1_03_in21 = imem04_in[23:20];
    69: op1_03_in21 = reg_0110;
    70: op1_03_in21 = reg_0088;
    71: op1_03_in21 = reg_0520;
    72: op1_03_in21 = reg_0426;
    74: op1_03_in21 = reg_0598;
    75: op1_03_in21 = reg_0720;
    76: op1_03_in21 = reg_0277;
    78: op1_03_in21 = reg_0351;
    79: op1_03_in21 = reg_0599;
    80: op1_03_in21 = reg_0069;
    81: op1_03_in21 = imem04_in[127:124];
    83: op1_03_in21 = reg_0628;
    84: op1_03_in21 = imem03_in[39:36];
    85: op1_03_in21 = reg_0296;
    86: op1_03_in21 = imem01_in[51:48];
    87: op1_03_in21 = reg_0741;
    88: op1_03_in21 = reg_0788;
    89: op1_03_in21 = reg_0805;
    90: op1_03_in21 = reg_0562;
    91: op1_03_in21 = reg_0755;
    92: op1_03_in21 = reg_0218;
    94: op1_03_in21 = reg_0037;
    95: op1_03_in21 = reg_0633;
    96: op1_03_in21 = reg_0233;
    default: op1_03_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv21 = 1;
    9: op1_03_inv21 = 1;
    12: op1_03_inv21 = 1;
    14: op1_03_inv21 = 1;
    18: op1_03_inv21 = 1;
    20: op1_03_inv21 = 1;
    21: op1_03_inv21 = 1;
    22: op1_03_inv21 = 1;
    23: op1_03_inv21 = 1;
    25: op1_03_inv21 = 1;
    29: op1_03_inv21 = 1;
    32: op1_03_inv21 = 1;
    36: op1_03_inv21 = 1;
    37: op1_03_inv21 = 1;
    40: op1_03_inv21 = 1;
    42: op1_03_inv21 = 1;
    43: op1_03_inv21 = 1;
    47: op1_03_inv21 = 1;
    48: op1_03_inv21 = 1;
    49: op1_03_inv21 = 1;
    50: op1_03_inv21 = 1;
    51: op1_03_inv21 = 1;
    55: op1_03_inv21 = 1;
    56: op1_03_inv21 = 1;
    58: op1_03_inv21 = 1;
    59: op1_03_inv21 = 1;
    60: op1_03_inv21 = 1;
    61: op1_03_inv21 = 1;
    63: op1_03_inv21 = 1;
    64: op1_03_inv21 = 1;
    65: op1_03_inv21 = 1;
    69: op1_03_inv21 = 1;
    70: op1_03_inv21 = 1;
    73: op1_03_inv21 = 1;
    75: op1_03_inv21 = 1;
    79: op1_03_inv21 = 1;
    80: op1_03_inv21 = 1;
    81: op1_03_inv21 = 1;
    83: op1_03_inv21 = 1;
    87: op1_03_inv21 = 1;
    90: op1_03_inv21 = 1;
    92: op1_03_inv21 = 1;
    94: op1_03_inv21 = 1;
    95: op1_03_inv21 = 1;
    default: op1_03_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in22 = imem06_in[35:32];
    5: op1_03_in22 = reg_0388;
    6: op1_03_in22 = reg_0712;
    7: op1_03_in22 = reg_0311;
    8: op1_03_in22 = reg_0488;
    9: op1_03_in22 = reg_0483;
    10: op1_03_in22 = reg_0631;
    11: op1_03_in22 = reg_0289;
    12: op1_03_in22 = reg_0750;
    13: op1_03_in22 = reg_0095;
    41: op1_03_in22 = reg_0095;
    14: op1_03_in22 = reg_0070;
    15: op1_03_in22 = reg_0039;
    16: op1_03_in22 = reg_0825;
    17: op1_03_in22 = reg_0268;
    18: op1_03_in22 = reg_0353;
    19: op1_03_in22 = reg_0498;
    20: op1_03_in22 = reg_0821;
    21: op1_03_in22 = imem05_in[7:4];
    22: op1_03_in22 = reg_0604;
    23: op1_03_in22 = reg_0385;
    24: op1_03_in22 = imem07_in[107:104];
    25: op1_03_in22 = reg_0238;
    26: op1_03_in22 = imem07_in[95:92];
    27: op1_03_in22 = imem01_in[99:96];
    28: op1_03_in22 = reg_0085;
    29: op1_03_in22 = reg_0775;
    30: op1_03_in22 = reg_0496;
    31: op1_03_in22 = reg_0801;
    32: op1_03_in22 = imem06_in[63:60];
    33: op1_03_in22 = reg_0449;
    34: op1_03_in22 = reg_0783;
    35: op1_03_in22 = imem04_in[87:84];
    36: op1_03_in22 = reg_0742;
    37: op1_03_in22 = reg_0272;
    38: op1_03_in22 = imem06_in[127:124];
    40: op1_03_in22 = reg_0701;
    42: op1_03_in22 = reg_0305;
    43: op1_03_in22 = imem07_in[19:16];
    44: op1_03_in22 = reg_0194;
    45: op1_03_in22 = reg_0565;
    46: op1_03_in22 = reg_0339;
    47: op1_03_in22 = reg_0709;
    48: op1_03_in22 = reg_0562;
    49: op1_03_in22 = reg_0656;
    50: op1_03_in22 = imem01_in[127:124];
    51: op1_03_in22 = reg_0702;
    53: op1_03_in22 = reg_0237;
    54: op1_03_in22 = imem02_in[3:0];
    55: op1_03_in22 = reg_0323;
    56: op1_03_in22 = reg_0516;
    57: op1_03_in22 = reg_0513;
    58: op1_03_in22 = reg_0599;
    59: op1_03_in22 = reg_0654;
    60: op1_03_in22 = imem05_in[63:60];
    96: op1_03_in22 = imem05_in[63:60];
    61: op1_03_in22 = reg_0293;
    62: op1_03_in22 = imem01_in[39:36];
    63: op1_03_in22 = reg_0217;
    64: op1_03_in22 = imem03_in[75:72];
    65: op1_03_in22 = imem03_in[23:20];
    66: op1_03_in22 = reg_0341;
    67: op1_03_in22 = imem04_in[91:88];
    69: op1_03_in22 = reg_0422;
    70: op1_03_in22 = reg_0555;
    71: op1_03_in22 = reg_0741;
    72: op1_03_in22 = reg_0352;
    73: op1_03_in22 = imem03_in[123:120];
    74: op1_03_in22 = imem05_in[27:24];
    75: op1_03_in22 = reg_0726;
    76: op1_03_in22 = reg_0729;
    78: op1_03_in22 = reg_0518;
    79: op1_03_in22 = reg_0579;
    80: op1_03_in22 = reg_0068;
    81: op1_03_in22 = reg_0316;
    83: op1_03_in22 = reg_0580;
    84: op1_03_in22 = imem03_in[55:52];
    85: op1_03_in22 = reg_0233;
    86: op1_03_in22 = imem01_in[71:68];
    87: op1_03_in22 = reg_0224;
    88: op1_03_in22 = reg_0782;
    89: op1_03_in22 = reg_0350;
    90: op1_03_in22 = reg_0549;
    91: op1_03_in22 = reg_0733;
    92: op1_03_in22 = reg_0664;
    93: op1_03_in22 = imem07_in[119:116];
    94: op1_03_in22 = imem07_in[27:24];
    95: op1_03_in22 = reg_0650;
    default: op1_03_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv22 = 1;
    5: op1_03_inv22 = 1;
    6: op1_03_inv22 = 1;
    8: op1_03_inv22 = 1;
    10: op1_03_inv22 = 1;
    11: op1_03_inv22 = 1;
    12: op1_03_inv22 = 1;
    13: op1_03_inv22 = 1;
    15: op1_03_inv22 = 1;
    16: op1_03_inv22 = 1;
    18: op1_03_inv22 = 1;
    19: op1_03_inv22 = 1;
    21: op1_03_inv22 = 1;
    23: op1_03_inv22 = 1;
    24: op1_03_inv22 = 1;
    25: op1_03_inv22 = 1;
    27: op1_03_inv22 = 1;
    28: op1_03_inv22 = 1;
    30: op1_03_inv22 = 1;
    31: op1_03_inv22 = 1;
    32: op1_03_inv22 = 1;
    33: op1_03_inv22 = 1;
    35: op1_03_inv22 = 1;
    37: op1_03_inv22 = 1;
    40: op1_03_inv22 = 1;
    41: op1_03_inv22 = 1;
    42: op1_03_inv22 = 1;
    43: op1_03_inv22 = 1;
    44: op1_03_inv22 = 1;
    45: op1_03_inv22 = 1;
    51: op1_03_inv22 = 1;
    54: op1_03_inv22 = 1;
    56: op1_03_inv22 = 1;
    57: op1_03_inv22 = 1;
    58: op1_03_inv22 = 1;
    59: op1_03_inv22 = 1;
    63: op1_03_inv22 = 1;
    65: op1_03_inv22 = 1;
    66: op1_03_inv22 = 1;
    67: op1_03_inv22 = 1;
    70: op1_03_inv22 = 1;
    71: op1_03_inv22 = 1;
    73: op1_03_inv22 = 1;
    75: op1_03_inv22 = 1;
    79: op1_03_inv22 = 1;
    81: op1_03_inv22 = 1;
    88: op1_03_inv22 = 1;
    89: op1_03_inv22 = 1;
    90: op1_03_inv22 = 1;
    92: op1_03_inv22 = 1;
    93: op1_03_inv22 = 1;
    94: op1_03_inv22 = 1;
    95: op1_03_inv22 = 1;
    default: op1_03_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in23 = imem06_in[63:60];
    5: op1_03_in23 = reg_0323;
    6: op1_03_in23 = reg_0708;
    7: op1_03_in23 = reg_0369;
    8: op1_03_in23 = reg_0491;
    9: op1_03_in23 = reg_0781;
    10: op1_03_in23 = reg_0622;
    46: op1_03_in23 = reg_0622;
    11: op1_03_in23 = reg_0306;
    12: op1_03_in23 = reg_0029;
    13: op1_03_in23 = reg_0086;
    14: op1_03_in23 = imem05_in[27:24];
    85: op1_03_in23 = imem05_in[27:24];
    15: op1_03_in23 = reg_0747;
    16: op1_03_in23 = reg_0515;
    17: op1_03_in23 = reg_0527;
    18: op1_03_in23 = reg_0347;
    19: op1_03_in23 = reg_0526;
    20: op1_03_in23 = reg_0235;
    21: op1_03_in23 = imem05_in[83:80];
    22: op1_03_in23 = reg_0611;
    23: op1_03_in23 = reg_0376;
    24: op1_03_in23 = imem07_in[115:112];
    25: op1_03_in23 = reg_0243;
    26: op1_03_in23 = imem07_in[119:116];
    27: op1_03_in23 = imem01_in[115:112];
    28: op1_03_in23 = reg_0733;
    29: op1_03_in23 = reg_0403;
    30: op1_03_in23 = reg_0513;
    31: op1_03_in23 = reg_0009;
    32: op1_03_in23 = imem06_in[67:64];
    33: op1_03_in23 = reg_0444;
    34: op1_03_in23 = reg_0786;
    35: op1_03_in23 = imem04_in[107:104];
    36: op1_03_in23 = reg_0275;
    37: op1_03_in23 = reg_0285;
    38: op1_03_in23 = reg_0402;
    40: op1_03_in23 = reg_0430;
    41: op1_03_in23 = reg_0096;
    42: op1_03_in23 = reg_0615;
    43: op1_03_in23 = imem07_in[127:124];
    44: op1_03_in23 = reg_0206;
    45: op1_03_in23 = reg_0592;
    47: op1_03_in23 = reg_0711;
    48: op1_03_in23 = reg_0572;
    49: op1_03_in23 = reg_0346;
    50: op1_03_in23 = reg_0085;
    51: op1_03_in23 = reg_0334;
    53: op1_03_in23 = reg_0734;
    54: op1_03_in23 = imem02_in[27:24];
    55: op1_03_in23 = reg_0541;
    78: op1_03_in23 = reg_0541;
    56: op1_03_in23 = reg_0303;
    57: op1_03_in23 = reg_0078;
    58: op1_03_in23 = reg_0750;
    59: op1_03_in23 = reg_0375;
    60: op1_03_in23 = imem05_in[79:76];
    61: op1_03_in23 = reg_0628;
    62: op1_03_in23 = imem01_in[55:52];
    63: op1_03_in23 = reg_0244;
    64: op1_03_in23 = imem03_in[83:80];
    65: op1_03_in23 = imem03_in[27:24];
    66: op1_03_in23 = reg_0356;
    67: op1_03_in23 = reg_0083;
    69: op1_03_in23 = reg_0220;
    70: op1_03_in23 = reg_0536;
    71: op1_03_in23 = reg_0385;
    72: op1_03_in23 = reg_0344;
    73: op1_03_in23 = reg_0317;
    74: op1_03_in23 = imem05_in[31:28];
    75: op1_03_in23 = reg_0717;
    76: op1_03_in23 = reg_0295;
    79: op1_03_in23 = reg_0338;
    80: op1_03_in23 = reg_0259;
    81: op1_03_in23 = reg_0544;
    83: op1_03_in23 = reg_0620;
    84: op1_03_in23 = imem03_in[59:56];
    86: op1_03_in23 = imem01_in[95:92];
    87: op1_03_in23 = reg_0102;
    88: op1_03_in23 = reg_0517;
    89: op1_03_in23 = reg_0016;
    90: op1_03_in23 = reg_0496;
    91: op1_03_in23 = reg_0007;
    92: op1_03_in23 = imem07_in[43:40];
    93: op1_03_in23 = imem07_in[123:120];
    94: op1_03_in23 = imem07_in[31:28];
    95: op1_03_in23 = imem07_in[39:36];
    96: op1_03_in23 = imem05_in[71:68];
    default: op1_03_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv23 = 1;
    5: op1_03_inv23 = 1;
    6: op1_03_inv23 = 1;
    7: op1_03_inv23 = 1;
    8: op1_03_inv23 = 1;
    11: op1_03_inv23 = 1;
    13: op1_03_inv23 = 1;
    17: op1_03_inv23 = 1;
    18: op1_03_inv23 = 1;
    23: op1_03_inv23 = 1;
    25: op1_03_inv23 = 1;
    28: op1_03_inv23 = 1;
    31: op1_03_inv23 = 1;
    35: op1_03_inv23 = 1;
    37: op1_03_inv23 = 1;
    38: op1_03_inv23 = 1;
    40: op1_03_inv23 = 1;
    41: op1_03_inv23 = 1;
    43: op1_03_inv23 = 1;
    46: op1_03_inv23 = 1;
    50: op1_03_inv23 = 1;
    53: op1_03_inv23 = 1;
    54: op1_03_inv23 = 1;
    58: op1_03_inv23 = 1;
    59: op1_03_inv23 = 1;
    63: op1_03_inv23 = 1;
    64: op1_03_inv23 = 1;
    66: op1_03_inv23 = 1;
    67: op1_03_inv23 = 1;
    69: op1_03_inv23 = 1;
    70: op1_03_inv23 = 1;
    73: op1_03_inv23 = 1;
    74: op1_03_inv23 = 1;
    76: op1_03_inv23 = 1;
    78: op1_03_inv23 = 1;
    83: op1_03_inv23 = 1;
    84: op1_03_inv23 = 1;
    86: op1_03_inv23 = 1;
    87: op1_03_inv23 = 1;
    89: op1_03_inv23 = 1;
    90: op1_03_inv23 = 1;
    92: op1_03_inv23 = 1;
    93: op1_03_inv23 = 1;
    95: op1_03_inv23 = 1;
    96: op1_03_inv23 = 1;
    default: op1_03_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in24 = imem06_in[111:108];
    5: op1_03_in24 = reg_0389;
    6: op1_03_in24 = reg_0445;
    7: op1_03_in24 = reg_0323;
    8: op1_03_in24 = reg_0493;
    9: op1_03_in24 = reg_0490;
    10: op1_03_in24 = reg_0381;
    11: op1_03_in24 = reg_0292;
    12: op1_03_in24 = reg_0005;
    13: op1_03_in24 = reg_0094;
    14: op1_03_in24 = imem05_in[47:44];
    15: op1_03_in24 = reg_0819;
    16: op1_03_in24 = reg_0505;
    17: op1_03_in24 = reg_0266;
    18: op1_03_in24 = reg_0086;
    19: op1_03_in24 = reg_0791;
    20: op1_03_in24 = reg_0506;
    21: op1_03_in24 = imem05_in[103:100];
    22: op1_03_in24 = reg_0332;
    23: op1_03_in24 = reg_0331;
    24: op1_03_in24 = reg_0730;
    25: op1_03_in24 = reg_0122;
    26: op1_03_in24 = imem07_in[123:120];
    27: op1_03_in24 = reg_0758;
    28: op1_03_in24 = reg_0282;
    29: op1_03_in24 = reg_0311;
    30: op1_03_in24 = reg_0822;
    31: op1_03_in24 = imem04_in[11:8];
    32: op1_03_in24 = imem06_in[95:92];
    33: op1_03_in24 = reg_0443;
    34: op1_03_in24 = reg_0486;
    35: op1_03_in24 = reg_0316;
    36: op1_03_in24 = reg_0260;
    37: op1_03_in24 = reg_0148;
    38: op1_03_in24 = reg_0748;
    40: op1_03_in24 = reg_0432;
    56: op1_03_in24 = reg_0432;
    41: op1_03_in24 = reg_0540;
    42: op1_03_in24 = reg_0430;
    43: op1_03_in24 = reg_0703;
    44: op1_03_in24 = imem01_in[39:36];
    45: op1_03_in24 = reg_0600;
    46: op1_03_in24 = reg_0407;
    47: op1_03_in24 = reg_0053;
    48: op1_03_in24 = reg_0014;
    49: op1_03_in24 = reg_0417;
    50: op1_03_in24 = reg_0497;
    51: op1_03_in24 = reg_0636;
    53: op1_03_in24 = reg_0737;
    54: op1_03_in24 = imem02_in[115:112];
    55: op1_03_in24 = reg_0314;
    57: op1_03_in24 = reg_0643;
    58: op1_03_in24 = reg_0350;
    59: op1_03_in24 = reg_0593;
    60: op1_03_in24 = reg_0215;
    61: op1_03_in24 = reg_0031;
    62: op1_03_in24 = imem01_in[79:76];
    63: op1_03_in24 = reg_0419;
    64: op1_03_in24 = reg_0602;
    65: op1_03_in24 = imem03_in[39:36];
    66: op1_03_in24 = reg_0360;
    67: op1_03_in24 = reg_0554;
    69: op1_03_in24 = reg_0234;
    70: op1_03_in24 = reg_0308;
    71: op1_03_in24 = reg_0224;
    72: op1_03_in24 = reg_0361;
    73: op1_03_in24 = reg_0589;
    74: op1_03_in24 = imem05_in[75:72];
    75: op1_03_in24 = reg_0276;
    76: op1_03_in24 = reg_0436;
    78: op1_03_in24 = reg_0770;
    79: op1_03_in24 = reg_0028;
    80: op1_03_in24 = reg_0233;
    81: op1_03_in24 = reg_0542;
    83: op1_03_in24 = reg_0787;
    84: op1_03_in24 = reg_0604;
    85: op1_03_in24 = imem05_in[43:40];
    86: op1_03_in24 = imem01_in[107:104];
    87: op1_03_in24 = reg_0388;
    88: op1_03_in24 = reg_0552;
    89: op1_03_in24 = reg_0130;
    90: op1_03_in24 = reg_0637;
    91: op1_03_in24 = reg_0306;
    92: op1_03_in24 = imem07_in[79:76];
    93: op1_03_in24 = reg_0728;
    94: op1_03_in24 = imem07_in[63:60];
    95: op1_03_in24 = imem07_in[43:40];
    96: op1_03_in24 = imem05_in[79:76];
    default: op1_03_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_03_inv24 = 1;
    8: op1_03_inv24 = 1;
    9: op1_03_inv24 = 1;
    11: op1_03_inv24 = 1;
    13: op1_03_inv24 = 1;
    14: op1_03_inv24 = 1;
    17: op1_03_inv24 = 1;
    23: op1_03_inv24 = 1;
    24: op1_03_inv24 = 1;
    27: op1_03_inv24 = 1;
    29: op1_03_inv24 = 1;
    30: op1_03_inv24 = 1;
    31: op1_03_inv24 = 1;
    34: op1_03_inv24 = 1;
    35: op1_03_inv24 = 1;
    38: op1_03_inv24 = 1;
    40: op1_03_inv24 = 1;
    42: op1_03_inv24 = 1;
    43: op1_03_inv24 = 1;
    45: op1_03_inv24 = 1;
    46: op1_03_inv24 = 1;
    48: op1_03_inv24 = 1;
    50: op1_03_inv24 = 1;
    53: op1_03_inv24 = 1;
    59: op1_03_inv24 = 1;
    60: op1_03_inv24 = 1;
    61: op1_03_inv24 = 1;
    62: op1_03_inv24 = 1;
    63: op1_03_inv24 = 1;
    64: op1_03_inv24 = 1;
    65: op1_03_inv24 = 1;
    72: op1_03_inv24 = 1;
    73: op1_03_inv24 = 1;
    75: op1_03_inv24 = 1;
    78: op1_03_inv24 = 1;
    83: op1_03_inv24 = 1;
    86: op1_03_inv24 = 1;
    87: op1_03_inv24 = 1;
    89: op1_03_inv24 = 1;
    90: op1_03_inv24 = 1;
    95: op1_03_inv24 = 1;
    96: op1_03_inv24 = 1;
    default: op1_03_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in25 = reg_0620;
    5: op1_03_in25 = imem03_in[3:0];
    6: op1_03_in25 = reg_0435;
    7: op1_03_in25 = reg_0397;
    8: op1_03_in25 = reg_0782;
    9: op1_03_in25 = reg_0488;
    10: op1_03_in25 = reg_0372;
    11: op1_03_in25 = reg_0286;
    12: op1_03_in25 = reg_0038;
    13: op1_03_in25 = reg_0093;
    14: op1_03_in25 = imem05_in[95:92];
    15: op1_03_in25 = imem07_in[3:0];
    16: op1_03_in25 = reg_0240;
    17: op1_03_in25 = reg_0150;
    18: op1_03_in25 = reg_0090;
    19: op1_03_in25 = reg_0798;
    20: op1_03_in25 = reg_0239;
    21: op1_03_in25 = imem05_in[111:108];
    22: op1_03_in25 = reg_0356;
    23: op1_03_in25 = reg_0002;
    24: op1_03_in25 = reg_0709;
    25: op1_03_in25 = reg_0113;
    26: op1_03_in25 = reg_0716;
    94: op1_03_in25 = reg_0716;
    27: op1_03_in25 = reg_0501;
    28: op1_03_in25 = reg_0272;
    29: op1_03_in25 = reg_0753;
    30: op1_03_in25 = reg_0549;
    31: op1_03_in25 = imem04_in[35:32];
    32: op1_03_in25 = imem06_in[103:100];
    33: op1_03_in25 = reg_0420;
    34: op1_03_in25 = reg_0275;
    35: op1_03_in25 = reg_0553;
    36: op1_03_in25 = reg_0732;
    37: op1_03_in25 = reg_0146;
    38: op1_03_in25 = reg_0776;
    40: op1_03_in25 = reg_0426;
    41: op1_03_in25 = reg_0535;
    42: op1_03_in25 = reg_0258;
    71: op1_03_in25 = reg_0258;
    43: op1_03_in25 = reg_0729;
    44: op1_03_in25 = imem01_in[71:68];
    45: op1_03_in25 = reg_0751;
    88: op1_03_in25 = reg_0751;
    46: op1_03_in25 = reg_0773;
    47: op1_03_in25 = reg_0445;
    76: op1_03_in25 = reg_0445;
    48: op1_03_in25 = reg_0015;
    49: op1_03_in25 = reg_0548;
    50: op1_03_in25 = reg_0645;
    51: op1_03_in25 = reg_0333;
    53: op1_03_in25 = reg_0421;
    54: op1_03_in25 = imem02_in[119:116];
    55: op1_03_in25 = reg_0530;
    56: op1_03_in25 = reg_0305;
    57: op1_03_in25 = reg_0296;
    58: op1_03_in25 = reg_0399;
    59: op1_03_in25 = reg_0580;
    60: op1_03_in25 = reg_0103;
    61: op1_03_in25 = reg_0775;
    62: op1_03_in25 = imem01_in[87:84];
    63: op1_03_in25 = reg_0123;
    64: op1_03_in25 = reg_0582;
    65: op1_03_in25 = imem03_in[67:64];
    66: op1_03_in25 = reg_0095;
    67: op1_03_in25 = reg_0551;
    69: op1_03_in25 = reg_0424;
    70: op1_03_in25 = reg_0052;
    72: op1_03_in25 = reg_0363;
    73: op1_03_in25 = reg_0596;
    74: op1_03_in25 = imem05_in[87:84];
    75: op1_03_in25 = reg_0295;
    78: op1_03_in25 = reg_0498;
    79: op1_03_in25 = reg_0564;
    80: op1_03_in25 = imem05_in[63:60];
    81: op1_03_in25 = reg_0555;
    83: op1_03_in25 = reg_0767;
    84: op1_03_in25 = reg_0319;
    85: op1_03_in25 = imem05_in[103:100];
    86: op1_03_in25 = reg_0085;
    87: op1_03_in25 = reg_0130;
    89: op1_03_in25 = reg_0357;
    90: op1_03_in25 = reg_0557;
    91: op1_03_in25 = reg_0802;
    92: op1_03_in25 = imem07_in[111:108];
    93: op1_03_in25 = reg_0159;
    95: op1_03_in25 = imem07_in[115:112];
    96: op1_03_in25 = imem05_in[123:120];
    default: op1_03_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv25 = 1;
    5: op1_03_inv25 = 1;
    6: op1_03_inv25 = 1;
    8: op1_03_inv25 = 1;
    14: op1_03_inv25 = 1;
    20: op1_03_inv25 = 1;
    22: op1_03_inv25 = 1;
    23: op1_03_inv25 = 1;
    29: op1_03_inv25 = 1;
    30: op1_03_inv25 = 1;
    36: op1_03_inv25 = 1;
    37: op1_03_inv25 = 1;
    40: op1_03_inv25 = 1;
    42: op1_03_inv25 = 1;
    43: op1_03_inv25 = 1;
    44: op1_03_inv25 = 1;
    48: op1_03_inv25 = 1;
    53: op1_03_inv25 = 1;
    54: op1_03_inv25 = 1;
    57: op1_03_inv25 = 1;
    59: op1_03_inv25 = 1;
    61: op1_03_inv25 = 1;
    62: op1_03_inv25 = 1;
    63: op1_03_inv25 = 1;
    64: op1_03_inv25 = 1;
    67: op1_03_inv25 = 1;
    69: op1_03_inv25 = 1;
    70: op1_03_inv25 = 1;
    71: op1_03_inv25 = 1;
    74: op1_03_inv25 = 1;
    76: op1_03_inv25 = 1;
    78: op1_03_inv25 = 1;
    81: op1_03_inv25 = 1;
    83: op1_03_inv25 = 1;
    84: op1_03_inv25 = 1;
    87: op1_03_inv25 = 1;
    88: op1_03_inv25 = 1;
    89: op1_03_inv25 = 1;
    93: op1_03_inv25 = 1;
    94: op1_03_inv25 = 1;
    default: op1_03_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in26 = reg_0621;
    5: op1_03_in26 = imem03_in[75:72];
    6: op1_03_in26 = reg_0175;
    7: op1_03_in26 = reg_0393;
    8: op1_03_in26 = reg_0783;
    9: op1_03_in26 = reg_0795;
    10: op1_03_in26 = reg_0405;
    11: op1_03_in26 = reg_0275;
    12: op1_03_in26 = imem07_in[31:28];
    13: op1_03_in26 = imem03_in[3:0];
    14: op1_03_in26 = imem05_in[127:124];
    15: op1_03_in26 = imem07_in[39:36];
    16: op1_03_in26 = reg_0238;
    17: op1_03_in26 = reg_0151;
    18: op1_03_in26 = reg_0087;
    19: op1_03_in26 = reg_0793;
    20: op1_03_in26 = reg_0240;
    21: op1_03_in26 = reg_0798;
    22: op1_03_in26 = reg_0372;
    23: op1_03_in26 = reg_0807;
    24: op1_03_in26 = reg_0718;
    25: op1_03_in26 = reg_0270;
    26: op1_03_in26 = reg_0704;
    27: op1_03_in26 = reg_0520;
    28: op1_03_in26 = reg_0744;
    29: op1_03_in26 = reg_0812;
    30: op1_03_in26 = reg_0557;
    31: op1_03_in26 = imem04_in[43:40];
    32: op1_03_in26 = imem06_in[115:112];
    33: op1_03_in26 = reg_0180;
    34: op1_03_in26 = reg_0085;
    35: op1_03_in26 = reg_0328;
    36: op1_03_in26 = reg_0277;
    37: op1_03_in26 = reg_0130;
    38: op1_03_in26 = reg_0815;
    40: op1_03_in26 = reg_0428;
    41: op1_03_in26 = reg_0526;
    78: op1_03_in26 = reg_0526;
    42: op1_03_in26 = reg_0063;
    43: op1_03_in26 = reg_0711;
    44: op1_03_in26 = imem01_in[83:80];
    45: op1_03_in26 = reg_0590;
    46: op1_03_in26 = reg_0821;
    47: op1_03_in26 = reg_0446;
    48: op1_03_in26 = reg_0806;
    49: op1_03_in26 = reg_0665;
    50: op1_03_in26 = reg_0496;
    51: op1_03_in26 = reg_0442;
    53: op1_03_in26 = reg_0574;
    54: op1_03_in26 = reg_0642;
    55: op1_03_in26 = reg_0498;
    56: op1_03_in26 = reg_0433;
    57: op1_03_in26 = reg_0233;
    58: op1_03_in26 = reg_0331;
    59: op1_03_in26 = reg_0028;
    60: op1_03_in26 = reg_0279;
    61: op1_03_in26 = reg_0748;
    62: op1_03_in26 = reg_0646;
    63: op1_03_in26 = reg_0105;
    64: op1_03_in26 = reg_0600;
    73: op1_03_in26 = reg_0600;
    65: op1_03_in26 = reg_0493;
    66: op1_03_in26 = reg_0769;
    67: op1_03_in26 = reg_0510;
    69: op1_03_in26 = reg_0505;
    70: op1_03_in26 = reg_0611;
    71: op1_03_in26 = reg_0511;
    87: op1_03_in26 = reg_0511;
    72: op1_03_in26 = reg_0360;
    74: op1_03_in26 = reg_0337;
    75: op1_03_in26 = reg_0051;
    76: op1_03_in26 = reg_0449;
    79: op1_03_in26 = reg_0549;
    80: op1_03_in26 = imem05_in[67:64];
    81: op1_03_in26 = reg_0060;
    83: op1_03_in26 = reg_0367;
    84: op1_03_in26 = reg_0488;
    85: op1_03_in26 = reg_0791;
    86: op1_03_in26 = reg_0385;
    88: op1_03_in26 = reg_0579;
    89: op1_03_in26 = reg_0573;
    90: op1_03_in26 = reg_0290;
    91: op1_03_in26 = reg_0278;
    92: op1_03_in26 = reg_0710;
    93: op1_03_in26 = reg_0784;
    94: op1_03_in26 = reg_0784;
    95: op1_03_in26 = reg_0722;
    96: op1_03_in26 = reg_0666;
    default: op1_03_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_03_inv26 = 1;
    6: op1_03_inv26 = 1;
    9: op1_03_inv26 = 1;
    10: op1_03_inv26 = 1;
    11: op1_03_inv26 = 1;
    17: op1_03_inv26 = 1;
    18: op1_03_inv26 = 1;
    19: op1_03_inv26 = 1;
    20: op1_03_inv26 = 1;
    21: op1_03_inv26 = 1;
    24: op1_03_inv26 = 1;
    26: op1_03_inv26 = 1;
    27: op1_03_inv26 = 1;
    28: op1_03_inv26 = 1;
    30: op1_03_inv26 = 1;
    31: op1_03_inv26 = 1;
    32: op1_03_inv26 = 1;
    34: op1_03_inv26 = 1;
    36: op1_03_inv26 = 1;
    38: op1_03_inv26 = 1;
    41: op1_03_inv26 = 1;
    43: op1_03_inv26 = 1;
    46: op1_03_inv26 = 1;
    53: op1_03_inv26 = 1;
    55: op1_03_inv26 = 1;
    61: op1_03_inv26 = 1;
    65: op1_03_inv26 = 1;
    66: op1_03_inv26 = 1;
    70: op1_03_inv26 = 1;
    71: op1_03_inv26 = 1;
    74: op1_03_inv26 = 1;
    75: op1_03_inv26 = 1;
    79: op1_03_inv26 = 1;
    81: op1_03_inv26 = 1;
    83: op1_03_inv26 = 1;
    85: op1_03_inv26 = 1;
    86: op1_03_inv26 = 1;
    87: op1_03_inv26 = 1;
    89: op1_03_inv26 = 1;
    90: op1_03_inv26 = 1;
    92: op1_03_inv26 = 1;
    93: op1_03_inv26 = 1;
    94: op1_03_inv26 = 1;
    95: op1_03_inv26 = 1;
    96: op1_03_inv26 = 1;
    default: op1_03_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in27 = reg_0622;
    5: op1_03_in27 = imem04_in[3:0];
    90: op1_03_in27 = imem04_in[3:0];
    6: op1_03_in27 = reg_0172;
    47: op1_03_in27 = reg_0172;
    7: op1_03_in27 = reg_0000;
    8: op1_03_in27 = reg_0485;
    9: op1_03_in27 = reg_0793;
    10: op1_03_in27 = reg_0375;
    11: op1_03_in27 = reg_0288;
    12: op1_03_in27 = imem07_in[75:72];
    13: op1_03_in27 = imem03_in[11:8];
    14: op1_03_in27 = reg_0482;
    15: op1_03_in27 = imem07_in[43:40];
    16: op1_03_in27 = reg_0243;
    17: op1_03_in27 = reg_0146;
    18: op1_03_in27 = reg_0094;
    19: op1_03_in27 = reg_0794;
    20: op1_03_in27 = reg_0504;
    21: op1_03_in27 = reg_0797;
    22: op1_03_in27 = reg_0407;
    23: op1_03_in27 = reg_0270;
    24: op1_03_in27 = reg_0706;
    25: op1_03_in27 = reg_0319;
    26: op1_03_in27 = reg_0726;
    27: op1_03_in27 = reg_0549;
    28: op1_03_in27 = reg_0285;
    29: op1_03_in27 = reg_0813;
    30: op1_03_in27 = reg_0761;
    50: op1_03_in27 = reg_0761;
    31: op1_03_in27 = imem04_in[59:56];
    32: op1_03_in27 = reg_0609;
    33: op1_03_in27 = reg_0161;
    34: op1_03_in27 = reg_0226;
    35: op1_03_in27 = reg_0056;
    36: op1_03_in27 = reg_0156;
    88: op1_03_in27 = reg_0156;
    37: op1_03_in27 = reg_0144;
    38: op1_03_in27 = reg_0368;
    40: op1_03_in27 = reg_0443;
    41: op1_03_in27 = reg_0740;
    78: op1_03_in27 = reg_0740;
    42: op1_03_in27 = reg_0296;
    43: op1_03_in27 = reg_0700;
    44: op1_03_in27 = imem01_in[99:96];
    45: op1_03_in27 = reg_0569;
    46: op1_03_in27 = reg_0776;
    48: op1_03_in27 = reg_0810;
    49: op1_03_in27 = reg_0352;
    51: op1_03_in27 = reg_0175;
    53: op1_03_in27 = reg_0054;
    54: op1_03_in27 = reg_0650;
    55: op1_03_in27 = reg_0526;
    56: op1_03_in27 = reg_0529;
    57: op1_03_in27 = reg_0644;
    58: op1_03_in27 = reg_0383;
    59: op1_03_in27 = reg_0367;
    60: op1_03_in27 = reg_0224;
    61: op1_03_in27 = reg_0593;
    62: op1_03_in27 = reg_0735;
    63: op1_03_in27 = reg_0126;
    64: op1_03_in27 = reg_0331;
    65: op1_03_in27 = reg_0357;
    84: op1_03_in27 = reg_0357;
    66: op1_03_in27 = reg_0757;
    67: op1_03_in27 = reg_0779;
    69: op1_03_in27 = reg_0420;
    70: op1_03_in27 = reg_0629;
    71: op1_03_in27 = reg_0422;
    87: op1_03_in27 = reg_0422;
    72: op1_03_in27 = reg_0097;
    73: op1_03_in27 = reg_0595;
    74: op1_03_in27 = reg_0736;
    75: op1_03_in27 = reg_0447;
    76: op1_03_in27 = reg_0440;
    79: op1_03_in27 = reg_0733;
    80: op1_03_in27 = imem05_in[119:116];
    81: op1_03_in27 = reg_0558;
    83: op1_03_in27 = imem07_in[19:16];
    85: op1_03_in27 = reg_0499;
    86: op1_03_in27 = reg_0820;
    89: op1_03_in27 = reg_0799;
    91: op1_03_in27 = reg_0216;
    92: op1_03_in27 = reg_0391;
    95: op1_03_in27 = reg_0391;
    93: op1_03_in27 = reg_0725;
    94: op1_03_in27 = reg_0166;
    96: op1_03_in27 = reg_0788;
    default: op1_03_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv27 = 1;
    5: op1_03_inv27 = 1;
    9: op1_03_inv27 = 1;
    10: op1_03_inv27 = 1;
    11: op1_03_inv27 = 1;
    13: op1_03_inv27 = 1;
    15: op1_03_inv27 = 1;
    16: op1_03_inv27 = 1;
    24: op1_03_inv27 = 1;
    26: op1_03_inv27 = 1;
    28: op1_03_inv27 = 1;
    33: op1_03_inv27 = 1;
    34: op1_03_inv27 = 1;
    35: op1_03_inv27 = 1;
    36: op1_03_inv27 = 1;
    37: op1_03_inv27 = 1;
    38: op1_03_inv27 = 1;
    40: op1_03_inv27 = 1;
    41: op1_03_inv27 = 1;
    42: op1_03_inv27 = 1;
    43: op1_03_inv27 = 1;
    46: op1_03_inv27 = 1;
    50: op1_03_inv27 = 1;
    54: op1_03_inv27 = 1;
    55: op1_03_inv27 = 1;
    57: op1_03_inv27 = 1;
    59: op1_03_inv27 = 1;
    61: op1_03_inv27 = 1;
    62: op1_03_inv27 = 1;
    64: op1_03_inv27 = 1;
    67: op1_03_inv27 = 1;
    72: op1_03_inv27 = 1;
    75: op1_03_inv27 = 1;
    76: op1_03_inv27 = 1;
    84: op1_03_inv27 = 1;
    89: op1_03_inv27 = 1;
    91: op1_03_inv27 = 1;
    default: op1_03_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in28 = reg_0623;
    5: op1_03_in28 = imem04_in[23:20];
    6: op1_03_in28 = reg_0181;
    7: op1_03_in28 = reg_0004;
    8: op1_03_in28 = reg_0267;
    76: op1_03_in28 = reg_0267;
    9: op1_03_in28 = reg_0494;
    10: op1_03_in28 = reg_0404;
    11: op1_03_in28 = reg_0307;
    12: op1_03_in28 = imem07_in[83:80];
    13: op1_03_in28 = imem03_in[15:12];
    14: op1_03_in28 = reg_0488;
    15: op1_03_in28 = imem07_in[47:44];
    16: op1_03_in28 = reg_0105;
    17: op1_03_in28 = reg_0138;
    18: op1_03_in28 = imem03_in[11:8];
    41: op1_03_in28 = imem03_in[11:8];
    55: op1_03_in28 = imem03_in[11:8];
    19: op1_03_in28 = reg_0783;
    20: op1_03_in28 = reg_0245;
    21: op1_03_in28 = reg_0789;
    22: op1_03_in28 = reg_0337;
    54: op1_03_in28 = reg_0337;
    23: op1_03_in28 = reg_0318;
    25: op1_03_in28 = reg_0318;
    24: op1_03_in28 = reg_0425;
    26: op1_03_in28 = reg_0725;
    27: op1_03_in28 = reg_0487;
    28: op1_03_in28 = reg_0147;
    29: op1_03_in28 = reg_0035;
    30: op1_03_in28 = reg_0760;
    31: op1_03_in28 = imem04_in[71:68];
    32: op1_03_in28 = reg_0622;
    33: op1_03_in28 = reg_0182;
    34: op1_03_in28 = reg_0732;
    35: op1_03_in28 = reg_0043;
    36: op1_03_in28 = reg_0032;
    37: op1_03_in28 = imem06_in[23:20];
    38: op1_03_in28 = reg_0037;
    40: op1_03_in28 = reg_0175;
    42: op1_03_in28 = reg_0075;
    43: op1_03_in28 = reg_0441;
    44: op1_03_in28 = reg_0758;
    45: op1_03_in28 = reg_0499;
    46: op1_03_in28 = reg_0614;
    47: op1_03_in28 = reg_0167;
    48: op1_03_in28 = reg_0009;
    49: op1_03_in28 = reg_0349;
    50: op1_03_in28 = reg_0649;
    51: op1_03_in28 = reg_0180;
    53: op1_03_in28 = reg_0244;
    56: op1_03_in28 = reg_0503;
    57: op1_03_in28 = imem05_in[27:24];
    58: op1_03_in28 = reg_0385;
    59: op1_03_in28 = imem07_in[3:0];
    60: op1_03_in28 = reg_0249;
    61: op1_03_in28 = reg_0819;
    62: op1_03_in28 = reg_0741;
    63: op1_03_in28 = imem02_in[47:44];
    64: op1_03_in28 = reg_0395;
    65: op1_03_in28 = reg_0561;
    66: op1_03_in28 = imem03_in[23:20];
    67: op1_03_in28 = reg_0679;
    69: op1_03_in28 = reg_0124;
    70: op1_03_in28 = reg_0508;
    71: op1_03_in28 = reg_0420;
    72: op1_03_in28 = reg_0757;
    73: op1_03_in28 = reg_0751;
    74: op1_03_in28 = reg_0788;
    75: op1_03_in28 = reg_0635;
    78: op1_03_in28 = imem03_in[19:16];
    79: op1_03_in28 = reg_0387;
    80: op1_03_in28 = imem05_in[123:120];
    81: op1_03_in28 = reg_0283;
    83: op1_03_in28 = imem07_in[59:56];
    84: op1_03_in28 = reg_0384;
    85: op1_03_in28 = reg_0326;
    86: op1_03_in28 = reg_0507;
    87: op1_03_in28 = reg_0217;
    88: op1_03_in28 = reg_0154;
    89: op1_03_in28 = reg_0600;
    90: op1_03_in28 = imem04_in[19:16];
    91: op1_03_in28 = imem04_in[59:56];
    92: op1_03_in28 = reg_0723;
    93: op1_03_in28 = reg_0709;
    94: op1_03_in28 = reg_0731;
    95: op1_03_in28 = reg_0166;
    96: op1_03_in28 = reg_0782;
    default: op1_03_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv28 = 1;
    9: op1_03_inv28 = 1;
    11: op1_03_inv28 = 1;
    12: op1_03_inv28 = 1;
    13: op1_03_inv28 = 1;
    15: op1_03_inv28 = 1;
    16: op1_03_inv28 = 1;
    17: op1_03_inv28 = 1;
    18: op1_03_inv28 = 1;
    19: op1_03_inv28 = 1;
    25: op1_03_inv28 = 1;
    27: op1_03_inv28 = 1;
    28: op1_03_inv28 = 1;
    31: op1_03_inv28 = 1;
    32: op1_03_inv28 = 1;
    36: op1_03_inv28 = 1;
    40: op1_03_inv28 = 1;
    44: op1_03_inv28 = 1;
    46: op1_03_inv28 = 1;
    49: op1_03_inv28 = 1;
    56: op1_03_inv28 = 1;
    57: op1_03_inv28 = 1;
    58: op1_03_inv28 = 1;
    59: op1_03_inv28 = 1;
    60: op1_03_inv28 = 1;
    61: op1_03_inv28 = 1;
    62: op1_03_inv28 = 1;
    65: op1_03_inv28 = 1;
    67: op1_03_inv28 = 1;
    69: op1_03_inv28 = 1;
    72: op1_03_inv28 = 1;
    73: op1_03_inv28 = 1;
    74: op1_03_inv28 = 1;
    76: op1_03_inv28 = 1;
    78: op1_03_inv28 = 1;
    79: op1_03_inv28 = 1;
    81: op1_03_inv28 = 1;
    85: op1_03_inv28 = 1;
    86: op1_03_inv28 = 1;
    88: op1_03_inv28 = 1;
    91: op1_03_inv28 = 1;
    92: op1_03_inv28 = 1;
    93: op1_03_inv28 = 1;
    94: op1_03_inv28 = 1;
    96: op1_03_inv28 = 1;
    default: op1_03_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in29 = reg_0332;
    5: op1_03_in29 = imem04_in[71:68];
    6: op1_03_in29 = reg_0169;
    7: op1_03_in29 = imem04_in[3:0];
    8: op1_03_in29 = reg_0268;
    9: op1_03_in29 = reg_0785;
    10: op1_03_in29 = reg_0315;
    11: op1_03_in29 = reg_0062;
    12: op1_03_in29 = imem07_in[107:104];
    13: op1_03_in29 = imem03_in[55:52];
    14: op1_03_in29 = reg_0788;
    15: op1_03_in29 = imem07_in[63:60];
    16: op1_03_in29 = reg_0122;
    17: op1_03_in29 = reg_0129;
    18: op1_03_in29 = imem03_in[15:12];
    19: op1_03_in29 = imem05_in[59:56];
    20: op1_03_in29 = reg_0219;
    21: op1_03_in29 = reg_0491;
    22: op1_03_in29 = reg_0753;
    46: op1_03_in29 = reg_0753;
    60: op1_03_in29 = reg_0753;
    23: op1_03_in29 = reg_0559;
    24: op1_03_in29 = reg_0436;
    25: op1_03_in29 = reg_0339;
    26: op1_03_in29 = reg_0712;
    27: op1_03_in29 = reg_0760;
    28: op1_03_in29 = reg_0136;
    29: op1_03_in29 = reg_0752;
    30: op1_03_in29 = reg_0241;
    31: op1_03_in29 = imem04_in[99:96];
    32: op1_03_in29 = reg_0331;
    33: op1_03_in29 = reg_0170;
    34: op1_03_in29 = reg_0277;
    35: op1_03_in29 = reg_0555;
    36: op1_03_in29 = reg_0616;
    37: op1_03_in29 = imem06_in[91:88];
    38: op1_03_in29 = imem07_in[15:12];
    40: op1_03_in29 = reg_0167;
    41: op1_03_in29 = imem03_in[23:20];
    42: op1_03_in29 = imem05_in[11:8];
    43: op1_03_in29 = reg_0067;
    44: op1_03_in29 = reg_0512;
    45: op1_03_in29 = reg_0396;
    47: op1_03_in29 = reg_0160;
    51: op1_03_in29 = reg_0160;
    48: op1_03_in29 = reg_0258;
    49: op1_03_in29 = reg_0358;
    50: op1_03_in29 = reg_0322;
    53: op1_03_in29 = reg_0216;
    54: op1_03_in29 = reg_0661;
    55: op1_03_in29 = imem03_in[43:40];
    56: op1_03_in29 = reg_0431;
    57: op1_03_in29 = imem05_in[51:48];
    58: op1_03_in29 = reg_0747;
    59: op1_03_in29 = imem07_in[47:44];
    61: op1_03_in29 = reg_0507;
    62: op1_03_in29 = reg_0778;
    63: op1_03_in29 = imem02_in[55:52];
    64: op1_03_in29 = reg_0391;
    65: op1_03_in29 = reg_0564;
    66: op1_03_in29 = imem03_in[27:24];
    78: op1_03_in29 = imem03_in[27:24];
    67: op1_03_in29 = reg_0223;
    70: op1_03_in29 = reg_0223;
    69: op1_03_in29 = reg_0125;
    71: op1_03_in29 = reg_0105;
    72: op1_03_in29 = reg_0094;
    73: op1_03_in29 = reg_0028;
    74: op1_03_in29 = reg_0641;
    75: op1_03_in29 = reg_0439;
    76: op1_03_in29 = reg_0435;
    79: op1_03_in29 = reg_0013;
    80: op1_03_in29 = imem05_in[127:124];
    81: op1_03_in29 = reg_0305;
    83: op1_03_in29 = imem07_in[71:68];
    84: op1_03_in29 = reg_0568;
    85: op1_03_in29 = reg_0245;
    86: op1_03_in29 = reg_0235;
    87: op1_03_in29 = reg_0240;
    88: op1_03_in29 = reg_0137;
    89: op1_03_in29 = reg_0486;
    90: op1_03_in29 = imem04_in[23:20];
    91: op1_03_in29 = imem04_in[119:116];
    92: op1_03_in29 = reg_0166;
    93: op1_03_in29 = reg_0266;
    94: op1_03_in29 = reg_0444;
    95: op1_03_in29 = reg_0158;
    96: op1_03_in29 = reg_0517;
    default: op1_03_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv29 = 1;
    6: op1_03_inv29 = 1;
    7: op1_03_inv29 = 1;
    9: op1_03_inv29 = 1;
    13: op1_03_inv29 = 1;
    14: op1_03_inv29 = 1;
    16: op1_03_inv29 = 1;
    17: op1_03_inv29 = 1;
    18: op1_03_inv29 = 1;
    22: op1_03_inv29 = 1;
    23: op1_03_inv29 = 1;
    26: op1_03_inv29 = 1;
    27: op1_03_inv29 = 1;
    28: op1_03_inv29 = 1;
    29: op1_03_inv29 = 1;
    30: op1_03_inv29 = 1;
    31: op1_03_inv29 = 1;
    33: op1_03_inv29 = 1;
    36: op1_03_inv29 = 1;
    37: op1_03_inv29 = 1;
    40: op1_03_inv29 = 1;
    45: op1_03_inv29 = 1;
    49: op1_03_inv29 = 1;
    54: op1_03_inv29 = 1;
    56: op1_03_inv29 = 1;
    57: op1_03_inv29 = 1;
    62: op1_03_inv29 = 1;
    67: op1_03_inv29 = 1;
    69: op1_03_inv29 = 1;
    70: op1_03_inv29 = 1;
    72: op1_03_inv29 = 1;
    73: op1_03_inv29 = 1;
    74: op1_03_inv29 = 1;
    79: op1_03_inv29 = 1;
    80: op1_03_inv29 = 1;
    81: op1_03_inv29 = 1;
    83: op1_03_inv29 = 1;
    85: op1_03_inv29 = 1;
    89: op1_03_inv29 = 1;
    93: op1_03_inv29 = 1;
    94: op1_03_inv29 = 1;
    96: op1_03_inv29 = 1;
    default: op1_03_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_03_in30 = reg_0344;
    5: op1_03_in30 = reg_0543;
    6: op1_03_in30 = reg_0176;
    7: op1_03_in30 = imem04_in[7:4];
    8: op1_03_in30 = reg_0259;
    9: op1_03_in30 = reg_0495;
    10: op1_03_in30 = reg_0406;
    11: op1_03_in30 = reg_0065;
    12: op1_03_in30 = reg_0722;
    13: op1_03_in30 = imem03_in[107:104];
    14: op1_03_in30 = reg_0492;
    15: op1_03_in30 = imem07_in[91:88];
    16: op1_03_in30 = reg_0116;
    17: op1_03_in30 = reg_0153;
    18: op1_03_in30 = imem03_in[31:28];
    78: op1_03_in30 = imem03_in[31:28];
    19: op1_03_in30 = imem05_in[67:64];
    20: op1_03_in30 = reg_0123;
    21: op1_03_in30 = reg_0494;
    22: op1_03_in30 = reg_0040;
    23: op1_03_in30 = imem04_in[39:36];
    24: op1_03_in30 = reg_0423;
    25: op1_03_in30 = reg_0338;
    26: op1_03_in30 = reg_0709;
    27: op1_03_in30 = reg_0232;
    28: op1_03_in30 = reg_0133;
    29: op1_03_in30 = reg_0751;
    30: op1_03_in30 = reg_0511;
    31: op1_03_in30 = reg_0315;
    32: op1_03_in30 = reg_0577;
    33: op1_03_in30 = reg_0157;
    34: op1_03_in30 = reg_0135;
    35: op1_03_in30 = reg_0060;
    36: op1_03_in30 = reg_0608;
    37: op1_03_in30 = reg_0628;
    38: op1_03_in30 = imem07_in[51:48];
    40: op1_03_in30 = reg_0177;
    41: op1_03_in30 = imem03_in[99:96];
    42: op1_03_in30 = imem05_in[23:20];
    43: op1_03_in30 = reg_0053;
    44: op1_03_in30 = reg_0549;
    61: op1_03_in30 = reg_0549;
    45: op1_03_in30 = reg_0374;
    46: op1_03_in30 = reg_0620;
    47: op1_03_in30 = reg_0183;
    48: op1_03_in30 = reg_0249;
    49: op1_03_in30 = reg_0361;
    50: op1_03_in30 = reg_0100;
    51: op1_03_in30 = imem07_in[75:72];
    53: op1_03_in30 = reg_0290;
    54: op1_03_in30 = reg_0656;
    55: op1_03_in30 = imem03_in[59:56];
    56: op1_03_in30 = reg_0508;
    57: op1_03_in30 = reg_0798;
    58: op1_03_in30 = reg_0000;
    59: op1_03_in30 = imem07_in[59:56];
    60: op1_03_in30 = reg_0372;
    62: op1_03_in30 = reg_0652;
    63: op1_03_in30 = imem02_in[87:84];
    64: op1_03_in30 = reg_0755;
    65: op1_03_in30 = reg_0499;
    66: op1_03_in30 = imem03_in[39:36];
    67: op1_03_in30 = reg_0416;
    69: op1_03_in30 = reg_0104;
    70: op1_03_in30 = reg_0078;
    71: op1_03_in30 = reg_0670;
    72: op1_03_in30 = imem03_in[27:24];
    73: op1_03_in30 = reg_0568;
    74: op1_03_in30 = reg_0793;
    75: op1_03_in30 = reg_0239;
    76: op1_03_in30 = reg_0268;
    79: op1_03_in30 = reg_0804;
    80: op1_03_in30 = reg_0667;
    81: op1_03_in30 = reg_0280;
    83: op1_03_in30 = reg_0721;
    84: op1_03_in30 = reg_0398;
    85: op1_03_in30 = reg_0252;
    86: op1_03_in30 = reg_0241;
    87: op1_03_in30 = reg_0244;
    88: op1_03_in30 = reg_0165;
    89: op1_03_in30 = reg_0389;
    90: op1_03_in30 = imem04_in[47:44];
    91: op1_03_in30 = reg_0173;
    92: op1_03_in30 = reg_0164;
    93: op1_03_in30 = reg_0436;
    94: op1_03_in30 = reg_0084;
    95: op1_03_in30 = reg_0266;
    96: op1_03_in30 = reg_0797;
    default: op1_03_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_03_inv30 = 1;
    7: op1_03_inv30 = 1;
    8: op1_03_inv30 = 1;
    12: op1_03_inv30 = 1;
    13: op1_03_inv30 = 1;
    16: op1_03_inv30 = 1;
    17: op1_03_inv30 = 1;
    18: op1_03_inv30 = 1;
    19: op1_03_inv30 = 1;
    20: op1_03_inv30 = 1;
    22: op1_03_inv30 = 1;
    25: op1_03_inv30 = 1;
    26: op1_03_inv30 = 1;
    28: op1_03_inv30 = 1;
    29: op1_03_inv30 = 1;
    30: op1_03_inv30 = 1;
    32: op1_03_inv30 = 1;
    34: op1_03_inv30 = 1;
    37: op1_03_inv30 = 1;
    38: op1_03_inv30 = 1;
    40: op1_03_inv30 = 1;
    42: op1_03_inv30 = 1;
    43: op1_03_inv30 = 1;
    44: op1_03_inv30 = 1;
    47: op1_03_inv30 = 1;
    50: op1_03_inv30 = 1;
    51: op1_03_inv30 = 1;
    54: op1_03_inv30 = 1;
    55: op1_03_inv30 = 1;
    58: op1_03_inv30 = 1;
    59: op1_03_inv30 = 1;
    60: op1_03_inv30 = 1;
    61: op1_03_inv30 = 1;
    63: op1_03_inv30 = 1;
    65: op1_03_inv30 = 1;
    67: op1_03_inv30 = 1;
    69: op1_03_inv30 = 1;
    70: op1_03_inv30 = 1;
    73: op1_03_inv30 = 1;
    74: op1_03_inv30 = 1;
    83: op1_03_inv30 = 1;
    84: op1_03_inv30 = 1;
    88: op1_03_inv30 = 1;
    89: op1_03_inv30 = 1;
    92: op1_03_inv30 = 1;
    94: op1_03_inv30 = 1;
    95: op1_03_inv30 = 1;
    96: op1_03_inv30 = 1;
    default: op1_03_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_03_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_03_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in00 = reg_0401;
    5: op1_04_in00 = reg_0552;
    6: op1_04_in00 = imem00_in[11:8];
    7: op1_04_in00 = imem04_in[15:12];
    8: op1_04_in00 = reg_0256;
    9: op1_04_in00 = reg_0786;
    10: op1_04_in00 = reg_0367;
    3: op1_04_in00 = imem07_in[39:36];
    2: op1_04_in00 = imem07_in[39:36];
    11: op1_04_in00 = reg_0043;
    12: op1_04_in00 = imem00_in[3:0];
    52: op1_04_in00 = imem00_in[3:0];
    13: op1_04_in00 = reg_0598;
    41: op1_04_in00 = reg_0598;
    14: op1_04_in00 = reg_0493;
    15: op1_04_in00 = imem00_in[7:4];
    68: op1_04_in00 = imem00_in[7:4];
    16: op1_04_in00 = reg_0119;
    17: op1_04_in00 = imem06_in[27:24];
    18: op1_04_in00 = imem03_in[43:40];
    19: op1_04_in00 = imem05_in[95:92];
    20: op1_04_in00 = reg_0127;
    21: op1_04_in00 = reg_0785;
    22: op1_04_in00 = reg_0817;
    1: op1_04_in00 = imem07_in[35:32];
    23: op1_04_in00 = imem04_in[67:64];
    24: op1_04_in00 = imem00_in[67:64];
    25: op1_04_in00 = reg_0658;
    26: op1_04_in00 = reg_0697;
    27: op1_04_in00 = reg_0241;
    28: op1_04_in00 = reg_0152;
    29: op1_04_in00 = imem07_in[27:24];
    30: op1_04_in00 = reg_0506;
    31: op1_04_in00 = reg_0558;
    32: op1_04_in00 = reg_0762;
    33: op1_04_in00 = imem00_in[19:16];
    77: op1_04_in00 = imem00_in[19:16];
    34: op1_04_in00 = reg_0133;
    80: op1_04_in00 = reg_0133;
    35: op1_04_in00 = reg_0057;
    36: op1_04_in00 = reg_0237;
    37: op1_04_in00 = reg_0630;
    38: op1_04_in00 = imem07_in[75:72];
    39: op1_04_in00 = imem00_in[27:24];
    40: op1_04_in00 = reg_0171;
    42: op1_04_in00 = imem05_in[39:36];
    43: op1_04_in00 = reg_0447;
    93: op1_04_in00 = reg_0447;
    44: op1_04_in00 = reg_0515;
    45: op1_04_in00 = reg_0003;
    46: op1_04_in00 = reg_0231;
    47: op1_04_in00 = imem00_in[15:12];
    82: op1_04_in00 = imem00_in[15:12];
    48: op1_04_in00 = reg_0063;
    49: op1_04_in00 = reg_0324;
    50: op1_04_in00 = reg_0825;
    51: op1_04_in00 = reg_0183;
    53: op1_04_in00 = reg_0425;
    54: op1_04_in00 = reg_0346;
    55: op1_04_in00 = imem03_in[71:68];
    56: op1_04_in00 = reg_0050;
    57: op1_04_in00 = reg_0112;
    58: op1_04_in00 = reg_0006;
    59: op1_04_in00 = imem07_in[71:68];
    60: op1_04_in00 = reg_0227;
    61: op1_04_in00 = reg_0767;
    62: op1_04_in00 = reg_0760;
    63: op1_04_in00 = reg_0403;
    64: op1_04_in00 = reg_0376;
    65: op1_04_in00 = reg_0396;
    66: op1_04_in00 = imem03_in[51:48];
    67: op1_04_in00 = reg_0109;
    69: op1_04_in00 = reg_0121;
    70: op1_04_in00 = reg_0780;
    71: op1_04_in00 = reg_0108;
    72: op1_04_in00 = imem03_in[39:36];
    73: op1_04_in00 = reg_0368;
    74: op1_04_in00 = reg_0732;
    75: op1_04_in00 = reg_0449;
    76: op1_04_in00 = reg_0165;
    78: op1_04_in00 = imem03_in[47:44];
    79: op1_04_in00 = reg_0805;
    81: op1_04_in00 = reg_0076;
    83: op1_04_in00 = reg_0723;
    84: op1_04_in00 = reg_0747;
    85: op1_04_in00 = reg_0491;
    86: op1_04_in00 = reg_0567;
    87: op1_04_in00 = reg_0248;
    88: op1_04_in00 = reg_0794;
    89: op1_04_in00 = reg_0395;
    90: op1_04_in00 = imem04_in[51:48];
    91: op1_04_in00 = reg_0537;
    92: op1_04_in00 = reg_0064;
    94: op1_04_in00 = reg_0139;
    95: op1_04_in00 = reg_0295;
    96: op1_04_in00 = reg_0583;
    default: op1_04_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv00 = 1;
    5: op1_04_inv00 = 1;
    6: op1_04_inv00 = 1;
    12: op1_04_inv00 = 1;
    14: op1_04_inv00 = 1;
    15: op1_04_inv00 = 1;
    2: op1_04_inv00 = 1;
    17: op1_04_inv00 = 1;
    19: op1_04_inv00 = 1;
    20: op1_04_inv00 = 1;
    22: op1_04_inv00 = 1;
    23: op1_04_inv00 = 1;
    26: op1_04_inv00 = 1;
    31: op1_04_inv00 = 1;
    34: op1_04_inv00 = 1;
    35: op1_04_inv00 = 1;
    36: op1_04_inv00 = 1;
    37: op1_04_inv00 = 1;
    38: op1_04_inv00 = 1;
    39: op1_04_inv00 = 1;
    41: op1_04_inv00 = 1;
    43: op1_04_inv00 = 1;
    48: op1_04_inv00 = 1;
    51: op1_04_inv00 = 1;
    54: op1_04_inv00 = 1;
    55: op1_04_inv00 = 1;
    56: op1_04_inv00 = 1;
    57: op1_04_inv00 = 1;
    61: op1_04_inv00 = 1;
    62: op1_04_inv00 = 1;
    63: op1_04_inv00 = 1;
    66: op1_04_inv00 = 1;
    67: op1_04_inv00 = 1;
    72: op1_04_inv00 = 1;
    73: op1_04_inv00 = 1;
    74: op1_04_inv00 = 1;
    75: op1_04_inv00 = 1;
    76: op1_04_inv00 = 1;
    79: op1_04_inv00 = 1;
    82: op1_04_inv00 = 1;
    84: op1_04_inv00 = 1;
    86: op1_04_inv00 = 1;
    88: op1_04_inv00 = 1;
    92: op1_04_inv00 = 1;
    93: op1_04_inv00 = 1;
    94: op1_04_inv00 = 1;
    95: op1_04_inv00 = 1;
    default: op1_04_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in01 = reg_0028;
    10: op1_04_in01 = reg_0028;
    5: op1_04_in01 = reg_0532;
    6: op1_04_in01 = imem00_in[39:36];
    7: op1_04_in01 = imem04_in[19:16];
    8: op1_04_in01 = reg_0243;
    9: op1_04_in01 = reg_0790;
    3: op1_04_in01 = imem07_in[51:48];
    1: op1_04_in01 = imem07_in[51:48];
    11: op1_04_in01 = reg_0044;
    12: op1_04_in01 = imem00_in[27:24];
    82: op1_04_in01 = imem00_in[27:24];
    13: op1_04_in01 = reg_0572;
    14: op1_04_in01 = reg_0259;
    15: op1_04_in01 = imem00_in[23:20];
    16: op1_04_in01 = reg_0108;
    2: op1_04_in01 = imem07_in[63:60];
    17: op1_04_in01 = imem06_in[35:32];
    18: op1_04_in01 = imem03_in[51:48];
    19: op1_04_in01 = imem05_in[103:100];
    20: op1_04_in01 = reg_0121;
    21: op1_04_in01 = reg_0486;
    22: op1_04_in01 = reg_0816;
    23: op1_04_in01 = imem04_in[83:80];
    24: op1_04_in01 = imem00_in[83:80];
    25: op1_04_in01 = reg_0666;
    26: op1_04_in01 = reg_0683;
    27: op1_04_in01 = reg_0503;
    28: op1_04_in01 = reg_0146;
    29: op1_04_in01 = imem07_in[75:72];
    30: op1_04_in01 = reg_0104;
    31: op1_04_in01 = reg_0551;
    32: op1_04_in01 = reg_0405;
    33: op1_04_in01 = imem00_in[47:44];
    34: op1_04_in01 = reg_0151;
    35: op1_04_in01 = reg_0536;
    91: op1_04_in01 = reg_0536;
    36: op1_04_in01 = reg_0293;
    37: op1_04_in01 = reg_0613;
    38: op1_04_in01 = reg_0720;
    39: op1_04_in01 = imem00_in[43:40];
    41: op1_04_in01 = reg_0589;
    42: op1_04_in01 = imem05_in[47:44];
    43: op1_04_in01 = reg_0635;
    44: op1_04_in01 = reg_0557;
    45: op1_04_in01 = reg_0008;
    46: op1_04_in01 = reg_0632;
    47: op1_04_in01 = imem00_in[19:16];
    52: op1_04_in01 = imem00_in[19:16];
    68: op1_04_in01 = imem00_in[19:16];
    48: op1_04_in01 = reg_0090;
    49: op1_04_in01 = reg_0351;
    50: op1_04_in01 = reg_0321;
    51: op1_04_in01 = reg_0177;
    53: op1_04_in01 = reg_0234;
    54: op1_04_in01 = reg_0587;
    55: op1_04_in01 = imem03_in[119:116];
    56: op1_04_in01 = reg_0512;
    57: op1_04_in01 = reg_0793;
    58: op1_04_in01 = reg_0811;
    59: op1_04_in01 = reg_0708;
    60: op1_04_in01 = reg_0236;
    61: op1_04_in01 = imem07_in[11:8];
    62: op1_04_in01 = reg_0054;
    63: op1_04_in01 = reg_0563;
    64: op1_04_in01 = reg_0397;
    65: op1_04_in01 = reg_0808;
    66: op1_04_in01 = imem03_in[75:72];
    78: op1_04_in01 = imem03_in[75:72];
    67: op1_04_in01 = reg_0110;
    69: op1_04_in01 = imem02_in[55:52];
    70: op1_04_in01 = reg_0771;
    71: op1_04_in01 = reg_0601;
    72: op1_04_in01 = reg_0559;
    73: op1_04_in01 = reg_0496;
    74: op1_04_in01 = reg_0517;
    75: op1_04_in01 = reg_0443;
    76: op1_04_in01 = reg_0167;
    77: op1_04_in01 = imem00_in[99:96];
    79: op1_04_in01 = reg_0015;
    80: op1_04_in01 = reg_0227;
    81: op1_04_in01 = reg_0302;
    83: op1_04_in01 = reg_0161;
    84: op1_04_in01 = reg_0396;
    85: op1_04_in01 = reg_0229;
    96: op1_04_in01 = reg_0229;
    86: op1_04_in01 = reg_0240;
    87: op1_04_in01 = reg_0506;
    88: op1_04_in01 = reg_0278;
    89: op1_04_in01 = reg_0384;
    90: op1_04_in01 = imem04_in[67:64];
    92: op1_04_in01 = reg_0434;
    93: op1_04_in01 = reg_0239;
    94: op1_04_in01 = reg_0175;
    95: op1_04_in01 = reg_0436;
    default: op1_04_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv01 = 1;
    7: op1_04_inv01 = 1;
    10: op1_04_inv01 = 1;
    11: op1_04_inv01 = 1;
    12: op1_04_inv01 = 1;
    13: op1_04_inv01 = 1;
    17: op1_04_inv01 = 1;
    21: op1_04_inv01 = 1;
    1: op1_04_inv01 = 1;
    24: op1_04_inv01 = 1;
    25: op1_04_inv01 = 1;
    26: op1_04_inv01 = 1;
    27: op1_04_inv01 = 1;
    28: op1_04_inv01 = 1;
    29: op1_04_inv01 = 1;
    33: op1_04_inv01 = 1;
    34: op1_04_inv01 = 1;
    35: op1_04_inv01 = 1;
    36: op1_04_inv01 = 1;
    37: op1_04_inv01 = 1;
    41: op1_04_inv01 = 1;
    44: op1_04_inv01 = 1;
    45: op1_04_inv01 = 1;
    46: op1_04_inv01 = 1;
    48: op1_04_inv01 = 1;
    52: op1_04_inv01 = 1;
    53: op1_04_inv01 = 1;
    54: op1_04_inv01 = 1;
    56: op1_04_inv01 = 1;
    57: op1_04_inv01 = 1;
    59: op1_04_inv01 = 1;
    60: op1_04_inv01 = 1;
    61: op1_04_inv01 = 1;
    62: op1_04_inv01 = 1;
    63: op1_04_inv01 = 1;
    66: op1_04_inv01 = 1;
    69: op1_04_inv01 = 1;
    70: op1_04_inv01 = 1;
    72: op1_04_inv01 = 1;
    75: op1_04_inv01 = 1;
    76: op1_04_inv01 = 1;
    77: op1_04_inv01 = 1;
    80: op1_04_inv01 = 1;
    81: op1_04_inv01 = 1;
    83: op1_04_inv01 = 1;
    84: op1_04_inv01 = 1;
    85: op1_04_inv01 = 1;
    89: op1_04_inv01 = 1;
    90: op1_04_inv01 = 1;
    91: op1_04_inv01 = 1;
    92: op1_04_inv01 = 1;
    default: op1_04_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in02 = reg_0025;
    5: op1_04_in02 = reg_0301;
    6: op1_04_in02 = imem00_in[55:52];
    15: op1_04_in02 = imem00_in[55:52];
    52: op1_04_in02 = imem00_in[55:52];
    7: op1_04_in02 = imem04_in[59:56];
    8: op1_04_in02 = reg_0253;
    9: op1_04_in02 = reg_0485;
    10: op1_04_in02 = reg_0039;
    3: op1_04_in02 = imem07_in[75:72];
    11: op1_04_in02 = reg_0252;
    12: op1_04_in02 = imem00_in[75:72];
    13: op1_04_in02 = reg_0587;
    14: op1_04_in02 = reg_0224;
    16: op1_04_in02 = imem02_in[3:0];
    2: op1_04_in02 = imem07_in[95:92];
    17: op1_04_in02 = reg_0610;
    36: op1_04_in02 = reg_0610;
    18: op1_04_in02 = imem03_in[59:56];
    19: op1_04_in02 = imem05_in[115:112];
    20: op1_04_in02 = reg_0057;
    21: op1_04_in02 = reg_0225;
    22: op1_04_in02 = reg_0037;
    1: op1_04_in02 = imem07_in[59:56];
    23: op1_04_in02 = imem04_in[103:100];
    24: op1_04_in02 = imem00_in[87:84];
    25: op1_04_in02 = reg_0655;
    26: op1_04_in02 = reg_0698;
    27: op1_04_in02 = reg_0234;
    28: op1_04_in02 = reg_0156;
    29: op1_04_in02 = imem07_in[99:96];
    30: op1_04_in02 = reg_0119;
    31: op1_04_in02 = reg_0280;
    32: op1_04_in02 = reg_0404;
    33: op1_04_in02 = imem00_in[91:88];
    34: op1_04_in02 = reg_0128;
    80: op1_04_in02 = reg_0128;
    35: op1_04_in02 = reg_0523;
    37: op1_04_in02 = reg_0371;
    38: op1_04_in02 = reg_0730;
    39: op1_04_in02 = imem00_in[59:56];
    47: op1_04_in02 = imem00_in[59:56];
    41: op1_04_in02 = reg_0597;
    42: op1_04_in02 = imem05_in[55:52];
    43: op1_04_in02 = reg_0440;
    93: op1_04_in02 = reg_0440;
    44: op1_04_in02 = reg_0244;
    62: op1_04_in02 = reg_0244;
    45: op1_04_in02 = reg_0799;
    46: op1_04_in02 = imem07_in[7:4];
    48: op1_04_in02 = reg_0256;
    49: op1_04_in02 = reg_0073;
    50: op1_04_in02 = reg_0306;
    51: op1_04_in02 = reg_0168;
    53: op1_04_in02 = reg_0419;
    54: op1_04_in02 = reg_0358;
    55: op1_04_in02 = imem03_in[123:120];
    56: op1_04_in02 = reg_0078;
    57: op1_04_in02 = reg_0785;
    58: op1_04_in02 = reg_0003;
    65: op1_04_in02 = reg_0003;
    59: op1_04_in02 = reg_0709;
    60: op1_04_in02 = reg_0624;
    61: op1_04_in02 = imem07_in[67:64];
    63: op1_04_in02 = reg_0657;
    64: op1_04_in02 = reg_0386;
    66: op1_04_in02 = imem03_in[83:80];
    67: op1_04_in02 = reg_0111;
    68: op1_04_in02 = imem00_in[31:28];
    69: op1_04_in02 = imem02_in[99:96];
    70: op1_04_in02 = imem05_in[11:8];
    71: op1_04_in02 = reg_0678;
    72: op1_04_in02 = reg_0596;
    73: op1_04_in02 = reg_0387;
    74: op1_04_in02 = reg_0326;
    75: op1_04_in02 = reg_0084;
    76: op1_04_in02 = reg_0163;
    77: op1_04_in02 = imem00_in[127:124];
    78: op1_04_in02 = imem03_in[103:100];
    79: op1_04_in02 = reg_0806;
    81: op1_04_in02 = reg_0071;
    82: op1_04_in02 = imem00_in[47:44];
    83: op1_04_in02 = reg_0167;
    84: op1_04_in02 = reg_0570;
    85: op1_04_in02 = reg_0393;
    86: op1_04_in02 = reg_0216;
    87: op1_04_in02 = reg_0219;
    88: op1_04_in02 = reg_0289;
    89: op1_04_in02 = reg_0483;
    90: op1_04_in02 = imem04_in[91:88];
    91: op1_04_in02 = reg_0433;
    92: op1_04_in02 = reg_0446;
    94: op1_04_in02 = reg_0116;
    95: op1_04_in02 = reg_0333;
    96: op1_04_in02 = reg_0580;
    default: op1_04_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_04_inv02 = 1;
    3: op1_04_inv02 = 1;
    16: op1_04_inv02 = 1;
    2: op1_04_inv02 = 1;
    17: op1_04_inv02 = 1;
    20: op1_04_inv02 = 1;
    21: op1_04_inv02 = 1;
    22: op1_04_inv02 = 1;
    23: op1_04_inv02 = 1;
    27: op1_04_inv02 = 1;
    28: op1_04_inv02 = 1;
    32: op1_04_inv02 = 1;
    35: op1_04_inv02 = 1;
    42: op1_04_inv02 = 1;
    43: op1_04_inv02 = 1;
    45: op1_04_inv02 = 1;
    46: op1_04_inv02 = 1;
    47: op1_04_inv02 = 1;
    50: op1_04_inv02 = 1;
    51: op1_04_inv02 = 1;
    55: op1_04_inv02 = 1;
    58: op1_04_inv02 = 1;
    59: op1_04_inv02 = 1;
    60: op1_04_inv02 = 1;
    61: op1_04_inv02 = 1;
    64: op1_04_inv02 = 1;
    65: op1_04_inv02 = 1;
    66: op1_04_inv02 = 1;
    68: op1_04_inv02 = 1;
    69: op1_04_inv02 = 1;
    70: op1_04_inv02 = 1;
    72: op1_04_inv02 = 1;
    78: op1_04_inv02 = 1;
    79: op1_04_inv02 = 1;
    80: op1_04_inv02 = 1;
    83: op1_04_inv02 = 1;
    85: op1_04_inv02 = 1;
    86: op1_04_inv02 = 1;
    88: op1_04_inv02 = 1;
    90: op1_04_inv02 = 1;
    92: op1_04_inv02 = 1;
    93: op1_04_inv02 = 1;
    96: op1_04_inv02 = 1;
    default: op1_04_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in03 = reg_0029;
    5: op1_04_in03 = reg_0291;
    6: op1_04_in03 = imem00_in[71:68];
    7: op1_04_in03 = imem04_in[79:76];
    8: op1_04_in03 = reg_0147;
    9: op1_04_in03 = reg_0787;
    10: op1_04_in03 = reg_0812;
    3: op1_04_in03 = imem07_in[127:124];
    11: op1_04_in03 = reg_0253;
    12: op1_04_in03 = imem00_in[79:76];
    13: op1_04_in03 = reg_0319;
    72: op1_04_in03 = reg_0319;
    14: op1_04_in03 = reg_0744;
    15: op1_04_in03 = imem00_in[63:60];
    52: op1_04_in03 = imem00_in[63:60];
    16: op1_04_in03 = imem02_in[47:44];
    2: op1_04_in03 = imem07_in[123:120];
    17: op1_04_in03 = reg_0626;
    18: op1_04_in03 = imem03_in[63:60];
    19: op1_04_in03 = imem05_in[123:120];
    42: op1_04_in03 = imem05_in[123:120];
    20: op1_04_in03 = reg_0088;
    21: op1_04_in03 = reg_0741;
    22: op1_04_in03 = imem07_in[3:0];
    23: op1_04_in03 = imem04_in[111:108];
    24: op1_04_in03 = reg_0693;
    47: op1_04_in03 = reg_0693;
    25: op1_04_in03 = reg_0653;
    26: op1_04_in03 = reg_0686;
    27: op1_04_in03 = reg_0508;
    28: op1_04_in03 = reg_0372;
    29: op1_04_in03 = reg_0720;
    30: op1_04_in03 = reg_0120;
    31: op1_04_in03 = reg_0267;
    32: op1_04_in03 = reg_0329;
    33: op1_04_in03 = reg_0677;
    34: op1_04_in03 = reg_0138;
    35: op1_04_in03 = reg_0058;
    36: op1_04_in03 = reg_0629;
    37: op1_04_in03 = reg_0622;
    38: op1_04_in03 = reg_0702;
    39: op1_04_in03 = imem00_in[87:84];
    41: op1_04_in03 = reg_0391;
    43: op1_04_in03 = reg_0437;
    75: op1_04_in03 = reg_0437;
    44: op1_04_in03 = reg_0603;
    45: op1_04_in03 = reg_0016;
    46: op1_04_in03 = imem07_in[19:16];
    48: op1_04_in03 = reg_0091;
    49: op1_04_in03 = reg_0347;
    50: op1_04_in03 = reg_0240;
    51: op1_04_in03 = reg_0173;
    53: op1_04_in03 = reg_0219;
    54: op1_04_in03 = reg_0341;
    55: op1_04_in03 = reg_0599;
    56: op1_04_in03 = reg_0585;
    57: op1_04_in03 = reg_0246;
    58: op1_04_in03 = reg_0807;
    59: op1_04_in03 = reg_0705;
    60: op1_04_in03 = reg_0605;
    61: op1_04_in03 = reg_0703;
    62: op1_04_in03 = reg_0425;
    63: op1_04_in03 = reg_0548;
    64: op1_04_in03 = reg_0389;
    65: op1_04_in03 = reg_0007;
    66: op1_04_in03 = imem03_in[99:96];
    67: op1_04_in03 = reg_0490;
    68: op1_04_in03 = imem00_in[59:56];
    69: op1_04_in03 = reg_0501;
    70: op1_04_in03 = imem05_in[51:48];
    71: op1_04_in03 = reg_0070;
    73: op1_04_in03 = reg_0747;
    74: op1_04_in03 = reg_0075;
    76: op1_04_in03 = reg_0185;
    77: op1_04_in03 = reg_0695;
    78: op1_04_in03 = reg_0063;
    79: op1_04_in03 = reg_0809;
    80: op1_04_in03 = reg_0146;
    81: op1_04_in03 = reg_0627;
    82: op1_04_in03 = imem00_in[83:80];
    83: op1_04_in03 = reg_0158;
    84: op1_04_in03 = reg_0006;
    85: op1_04_in03 = reg_0719;
    86: op1_04_in03 = reg_0290;
    87: op1_04_in03 = reg_0670;
    88: op1_04_in03 = reg_0625;
    89: op1_04_in03 = reg_0387;
    90: op1_04_in03 = reg_0555;
    91: op1_04_in03 = reg_0615;
    92: op1_04_in03 = reg_0440;
    93: op1_04_in03 = reg_0444;
    94: op1_04_in03 = reg_0110;
    95: op1_04_in03 = reg_0439;
    96: op1_04_in03 = reg_0495;
    default: op1_04_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv03 = 1;
    5: op1_04_inv03 = 1;
    8: op1_04_inv03 = 1;
    9: op1_04_inv03 = 1;
    10: op1_04_inv03 = 1;
    11: op1_04_inv03 = 1;
    14: op1_04_inv03 = 1;
    16: op1_04_inv03 = 1;
    2: op1_04_inv03 = 1;
    20: op1_04_inv03 = 1;
    22: op1_04_inv03 = 1;
    24: op1_04_inv03 = 1;
    25: op1_04_inv03 = 1;
    26: op1_04_inv03 = 1;
    27: op1_04_inv03 = 1;
    28: op1_04_inv03 = 1;
    29: op1_04_inv03 = 1;
    32: op1_04_inv03 = 1;
    33: op1_04_inv03 = 1;
    37: op1_04_inv03 = 1;
    38: op1_04_inv03 = 1;
    39: op1_04_inv03 = 1;
    44: op1_04_inv03 = 1;
    47: op1_04_inv03 = 1;
    48: op1_04_inv03 = 1;
    49: op1_04_inv03 = 1;
    50: op1_04_inv03 = 1;
    53: op1_04_inv03 = 1;
    56: op1_04_inv03 = 1;
    57: op1_04_inv03 = 1;
    59: op1_04_inv03 = 1;
    61: op1_04_inv03 = 1;
    62: op1_04_inv03 = 1;
    63: op1_04_inv03 = 1;
    64: op1_04_inv03 = 1;
    65: op1_04_inv03 = 1;
    66: op1_04_inv03 = 1;
    73: op1_04_inv03 = 1;
    74: op1_04_inv03 = 1;
    77: op1_04_inv03 = 1;
    78: op1_04_inv03 = 1;
    80: op1_04_inv03 = 1;
    81: op1_04_inv03 = 1;
    83: op1_04_inv03 = 1;
    84: op1_04_inv03 = 1;
    86: op1_04_inv03 = 1;
    87: op1_04_inv03 = 1;
    90: op1_04_inv03 = 1;
    92: op1_04_inv03 = 1;
    93: op1_04_inv03 = 1;
    94: op1_04_inv03 = 1;
    95: op1_04_inv03 = 1;
    96: op1_04_inv03 = 1;
    default: op1_04_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in04 = reg_0005;
    5: op1_04_in04 = reg_0053;
    6: op1_04_in04 = imem00_in[83:80];
    7: op1_04_in04 = imem04_in[127:124];
    8: op1_04_in04 = reg_0136;
    9: op1_04_in04 = reg_0268;
    10: op1_04_in04 = reg_0037;
    3: op1_04_in04 = reg_0430;
    11: op1_04_in04 = reg_0251;
    12: op1_04_in04 = imem00_in[123:120];
    13: op1_04_in04 = reg_0012;
    14: op1_04_in04 = reg_0263;
    15: op1_04_in04 = imem00_in[71:68];
    16: op1_04_in04 = imem02_in[95:92];
    2: op1_04_in04 = reg_0172;
    17: op1_04_in04 = reg_0632;
    18: op1_04_in04 = imem03_in[79:76];
    19: op1_04_in04 = reg_0133;
    20: op1_04_in04 = reg_0055;
    21: op1_04_in04 = reg_0226;
    22: op1_04_in04 = imem07_in[7:4];
    23: op1_04_in04 = imem04_in[119:116];
    24: op1_04_in04 = reg_0697;
    47: op1_04_in04 = reg_0697;
    77: op1_04_in04 = reg_0697;
    25: op1_04_in04 = reg_0640;
    26: op1_04_in04 = reg_0680;
    27: op1_04_in04 = reg_0120;
    87: op1_04_in04 = reg_0120;
    28: op1_04_in04 = reg_0020;
    29: op1_04_in04 = reg_0726;
    30: op1_04_in04 = reg_0112;
    31: op1_04_in04 = reg_0295;
    32: op1_04_in04 = reg_0038;
    33: op1_04_in04 = reg_0191;
    34: op1_04_in04 = reg_0153;
    35: op1_04_in04 = reg_0308;
    36: op1_04_in04 = reg_0617;
    37: op1_04_in04 = reg_0380;
    38: op1_04_in04 = reg_0708;
    39: op1_04_in04 = imem00_in[119:116];
    41: op1_04_in04 = reg_0564;
    42: op1_04_in04 = reg_0792;
    43: op1_04_in04 = reg_0267;
    44: op1_04_in04 = reg_0505;
    45: op1_04_in04 = reg_0010;
    46: op1_04_in04 = imem07_in[75:72];
    48: op1_04_in04 = reg_0560;
    49: op1_04_in04 = reg_0080;
    50: op1_04_in04 = reg_0216;
    52: op1_04_in04 = imem00_in[107:104];
    53: op1_04_in04 = reg_0673;
    54: op1_04_in04 = reg_0365;
    55: op1_04_in04 = reg_0596;
    56: op1_04_in04 = reg_0075;
    57: op1_04_in04 = reg_0099;
    58: op1_04_in04 = reg_0014;
    59: op1_04_in04 = reg_0707;
    60: op1_04_in04 = reg_0814;
    61: op1_04_in04 = reg_0334;
    62: op1_04_in04 = reg_0420;
    63: op1_04_in04 = reg_0355;
    64: op1_04_in04 = reg_0006;
    65: op1_04_in04 = reg_0806;
    66: op1_04_in04 = imem03_in[123:120];
    67: op1_04_in04 = reg_0085;
    68: op1_04_in04 = reg_0695;
    69: op1_04_in04 = reg_0666;
    70: op1_04_in04 = imem05_in[75:72];
    71: op1_04_in04 = reg_0641;
    72: op1_04_in04 = reg_0591;
    73: op1_04_in04 = reg_0649;
    74: op1_04_in04 = reg_0246;
    75: op1_04_in04 = reg_0175;
    76: op1_04_in04 = reg_0173;
    78: op1_04_in04 = reg_0582;
    79: op1_04_in04 = imem04_in[3:0];
    80: op1_04_in04 = reg_0113;
    81: op1_04_in04 = reg_0050;
    82: op1_04_in04 = imem00_in[91:88];
    83: op1_04_in04 = reg_0711;
    84: op1_04_in04 = reg_0811;
    85: op1_04_in04 = reg_0285;
    86: op1_04_in04 = reg_0506;
    88: op1_04_in04 = reg_0115;
    89: op1_04_in04 = reg_0747;
    90: op1_04_in04 = reg_0536;
    91: op1_04_in04 = reg_0529;
    92: op1_04_in04 = reg_0084;
    93: op1_04_in04 = reg_0116;
    94: op1_04_in04 = reg_0327;
    95: op1_04_in04 = reg_0066;
    96: op1_04_in04 = reg_0579;
    default: op1_04_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv04 = 1;
    5: op1_04_inv04 = 1;
    10: op1_04_inv04 = 1;
    14: op1_04_inv04 = 1;
    15: op1_04_inv04 = 1;
    2: op1_04_inv04 = 1;
    21: op1_04_inv04 = 1;
    26: op1_04_inv04 = 1;
    28: op1_04_inv04 = 1;
    30: op1_04_inv04 = 1;
    32: op1_04_inv04 = 1;
    33: op1_04_inv04 = 1;
    34: op1_04_inv04 = 1;
    35: op1_04_inv04 = 1;
    36: op1_04_inv04 = 1;
    39: op1_04_inv04 = 1;
    42: op1_04_inv04 = 1;
    44: op1_04_inv04 = 1;
    54: op1_04_inv04 = 1;
    58: op1_04_inv04 = 1;
    60: op1_04_inv04 = 1;
    62: op1_04_inv04 = 1;
    63: op1_04_inv04 = 1;
    64: op1_04_inv04 = 1;
    65: op1_04_inv04 = 1;
    67: op1_04_inv04 = 1;
    71: op1_04_inv04 = 1;
    72: op1_04_inv04 = 1;
    73: op1_04_inv04 = 1;
    74: op1_04_inv04 = 1;
    78: op1_04_inv04 = 1;
    79: op1_04_inv04 = 1;
    80: op1_04_inv04 = 1;
    81: op1_04_inv04 = 1;
    83: op1_04_inv04 = 1;
    85: op1_04_inv04 = 1;
    86: op1_04_inv04 = 1;
    92: op1_04_inv04 = 1;
    default: op1_04_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in05 = imem07_in[7:4];
    5: op1_04_in05 = reg_0071;
    6: op1_04_in05 = imem00_in[107:104];
    7: op1_04_in05 = reg_0530;
    8: op1_04_in05 = reg_0133;
    9: op1_04_in05 = reg_0259;
    10: op1_04_in05 = reg_0818;
    3: op1_04_in05 = reg_0436;
    11: op1_04_in05 = reg_0490;
    12: op1_04_in05 = reg_0681;
    13: op1_04_in05 = reg_0002;
    14: op1_04_in05 = reg_0150;
    96: op1_04_in05 = reg_0150;
    15: op1_04_in05 = imem00_in[79:76];
    16: op1_04_in05 = imem02_in[111:108];
    2: op1_04_in05 = reg_0169;
    17: op1_04_in05 = reg_0622;
    18: op1_04_in05 = reg_0583;
    19: op1_04_in05 = reg_0142;
    93: op1_04_in05 = reg_0142;
    20: op1_04_in05 = reg_0087;
    21: op1_04_in05 = reg_0307;
    22: op1_04_in05 = imem07_in[35:32];
    23: op1_04_in05 = reg_0529;
    24: op1_04_in05 = reg_0696;
    25: op1_04_in05 = reg_0636;
    26: op1_04_in05 = reg_0687;
    27: op1_04_in05 = reg_0108;
    53: op1_04_in05 = reg_0108;
    28: op1_04_in05 = reg_0368;
    29: op1_04_in05 = reg_0705;
    30: op1_04_in05 = imem02_in[7:4];
    31: op1_04_in05 = reg_0061;
    32: op1_04_in05 = reg_0764;
    33: op1_04_in05 = reg_0188;
    34: op1_04_in05 = imem06_in[15:12];
    35: op1_04_in05 = reg_0283;
    36: op1_04_in05 = reg_0631;
    37: op1_04_in05 = reg_0331;
    38: op1_04_in05 = reg_0709;
    39: op1_04_in05 = imem00_in[123:120];
    41: op1_04_in05 = reg_0568;
    42: op1_04_in05 = reg_0494;
    43: op1_04_in05 = reg_0175;
    92: op1_04_in05 = reg_0175;
    44: op1_04_in05 = reg_0123;
    45: op1_04_in05 = reg_0063;
    46: op1_04_in05 = imem07_in[119:116];
    47: op1_04_in05 = reg_0689;
    52: op1_04_in05 = reg_0689;
    48: op1_04_in05 = reg_0554;
    49: op1_04_in05 = reg_0756;
    50: op1_04_in05 = reg_0603;
    54: op1_04_in05 = reg_0342;
    55: op1_04_in05 = reg_0600;
    56: op1_04_in05 = imem05_in[19:16];
    57: op1_04_in05 = reg_0249;
    58: op1_04_in05 = reg_0809;
    59: op1_04_in05 = reg_0447;
    60: op1_04_in05 = reg_0619;
    61: op1_04_in05 = reg_0053;
    62: op1_04_in05 = reg_0104;
    63: op1_04_in05 = reg_0426;
    64: op1_04_in05 = reg_0811;
    65: op1_04_in05 = reg_0810;
    66: op1_04_in05 = reg_0597;
    67: op1_04_in05 = reg_0090;
    68: op1_04_in05 = reg_0682;
    69: op1_04_in05 = reg_0647;
    70: op1_04_in05 = imem05_in[91:88];
    71: op1_04_in05 = reg_0665;
    72: op1_04_in05 = reg_0116;
    73: op1_04_in05 = reg_0004;
    74: op1_04_in05 = reg_0309;
    75: op1_04_in05 = reg_0172;
    77: op1_04_in05 = reg_0492;
    78: op1_04_in05 = reg_0604;
    79: op1_04_in05 = imem04_in[27:24];
    80: op1_04_in05 = reg_0782;
    81: op1_04_in05 = reg_0598;
    82: op1_04_in05 = imem00_in[119:116];
    83: op1_04_in05 = reg_0157;
    84: op1_04_in05 = reg_0001;
    85: op1_04_in05 = reg_0149;
    86: op1_04_in05 = reg_0424;
    87: op1_04_in05 = reg_0677;
    88: op1_04_in05 = reg_0815;
    89: op1_04_in05 = reg_0623;
    90: op1_04_in05 = reg_0551;
    91: op1_04_in05 = reg_0302;
    94: op1_04_in05 = reg_0066;
    95: op1_04_in05 = reg_0178;
    default: op1_04_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv05 = 1;
    7: op1_04_inv05 = 1;
    14: op1_04_inv05 = 1;
    15: op1_04_inv05 = 1;
    16: op1_04_inv05 = 1;
    2: op1_04_inv05 = 1;
    17: op1_04_inv05 = 1;
    19: op1_04_inv05 = 1;
    20: op1_04_inv05 = 1;
    22: op1_04_inv05 = 1;
    25: op1_04_inv05 = 1;
    26: op1_04_inv05 = 1;
    27: op1_04_inv05 = 1;
    32: op1_04_inv05 = 1;
    33: op1_04_inv05 = 1;
    34: op1_04_inv05 = 1;
    44: op1_04_inv05 = 1;
    46: op1_04_inv05 = 1;
    47: op1_04_inv05 = 1;
    49: op1_04_inv05 = 1;
    50: op1_04_inv05 = 1;
    52: op1_04_inv05 = 1;
    53: op1_04_inv05 = 1;
    54: op1_04_inv05 = 1;
    56: op1_04_inv05 = 1;
    58: op1_04_inv05 = 1;
    59: op1_04_inv05 = 1;
    60: op1_04_inv05 = 1;
    61: op1_04_inv05 = 1;
    62: op1_04_inv05 = 1;
    63: op1_04_inv05 = 1;
    64: op1_04_inv05 = 1;
    67: op1_04_inv05 = 1;
    68: op1_04_inv05 = 1;
    70: op1_04_inv05 = 1;
    71: op1_04_inv05 = 1;
    72: op1_04_inv05 = 1;
    74: op1_04_inv05 = 1;
    78: op1_04_inv05 = 1;
    79: op1_04_inv05 = 1;
    82: op1_04_inv05 = 1;
    83: op1_04_inv05 = 1;
    84: op1_04_inv05 = 1;
    85: op1_04_inv05 = 1;
    87: op1_04_inv05 = 1;
    95: op1_04_inv05 = 1;
    default: op1_04_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in06 = imem07_in[31:28];
    5: op1_04_in06 = reg_0070;
    6: op1_04_in06 = reg_0695;
    7: op1_04_in06 = reg_0553;
    8: op1_04_in06 = reg_0139;
    9: op1_04_in06 = reg_0273;
    10: op1_04_in06 = reg_0030;
    3: op1_04_in06 = reg_0442;
    11: op1_04_in06 = reg_0484;
    12: op1_04_in06 = reg_0685;
    13: op1_04_in06 = reg_0803;
    14: op1_04_in06 = reg_0142;
    15: op1_04_in06 = imem00_in[91:88];
    16: op1_04_in06 = imem02_in[115:112];
    2: op1_04_in06 = reg_0157;
    17: op1_04_in06 = reg_0348;
    18: op1_04_in06 = reg_0587;
    19: op1_04_in06 = reg_0156;
    20: op1_04_in06 = reg_0650;
    21: op1_04_in06 = reg_0084;
    22: op1_04_in06 = imem07_in[59:56];
    23: op1_04_in06 = reg_0306;
    24: op1_04_in06 = reg_0689;
    25: op1_04_in06 = reg_0667;
    71: op1_04_in06 = reg_0667;
    26: op1_04_in06 = reg_0453;
    27: op1_04_in06 = reg_0101;
    28: op1_04_in06 = reg_0399;
    29: op1_04_in06 = reg_0707;
    30: op1_04_in06 = imem02_in[35:32];
    31: op1_04_in06 = reg_0253;
    32: op1_04_in06 = reg_0040;
    33: op1_04_in06 = reg_0203;
    34: op1_04_in06 = imem06_in[51:48];
    35: op1_04_in06 = reg_0295;
    83: op1_04_in06 = reg_0295;
    36: op1_04_in06 = reg_0626;
    37: op1_04_in06 = reg_0407;
    38: op1_04_in06 = reg_0705;
    39: op1_04_in06 = reg_0679;
    41: op1_04_in06 = reg_0383;
    42: op1_04_in06 = reg_0736;
    43: op1_04_in06 = reg_0180;
    44: op1_04_in06 = reg_0118;
    45: op1_04_in06 = reg_0075;
    46: op1_04_in06 = reg_0722;
    47: op1_04_in06 = reg_0684;
    52: op1_04_in06 = reg_0684;
    48: op1_04_in06 = reg_0071;
    91: op1_04_in06 = reg_0071;
    49: op1_04_in06 = imem03_in[3:0];
    50: op1_04_in06 = reg_0506;
    53: op1_04_in06 = reg_0106;
    87: op1_04_in06 = reg_0106;
    54: op1_04_in06 = reg_0514;
    55: op1_04_in06 = reg_0488;
    56: op1_04_in06 = imem05_in[67:64];
    57: op1_04_in06 = reg_0086;
    58: op1_04_in06 = reg_0520;
    59: op1_04_in06 = reg_0635;
    60: op1_04_in06 = reg_0618;
    61: op1_04_in06 = reg_0444;
    62: op1_04_in06 = reg_0675;
    63: op1_04_in06 = reg_0427;
    64: op1_04_in06 = imem04_in[11:8];
    65: op1_04_in06 = imem04_in[7:4];
    66: op1_04_in06 = reg_0493;
    67: op1_04_in06 = reg_0112;
    68: op1_04_in06 = reg_0697;
    69: op1_04_in06 = reg_0355;
    80: op1_04_in06 = reg_0355;
    70: op1_04_in06 = imem05_in[95:92];
    72: op1_04_in06 = reg_0329;
    73: op1_04_in06 = imem04_in[99:96];
    74: op1_04_in06 = reg_0236;
    75: op1_04_in06 = reg_0161;
    77: op1_04_in06 = reg_0658;
    78: op1_04_in06 = reg_0528;
    79: op1_04_in06 = imem04_in[43:40];
    81: op1_04_in06 = reg_0640;
    82: op1_04_in06 = reg_0696;
    84: op1_04_in06 = reg_0003;
    85: op1_04_in06 = reg_0781;
    86: op1_04_in06 = reg_0673;
    88: op1_04_in06 = reg_0370;
    89: op1_04_in06 = reg_0570;
    90: op1_04_in06 = reg_0174;
    92: op1_04_in06 = reg_0730;
    93: op1_04_in06 = reg_0185;
    96: op1_04_in06 = reg_0257;
    default: op1_04_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv06 = 1;
    6: op1_04_inv06 = 1;
    9: op1_04_inv06 = 1;
    3: op1_04_inv06 = 1;
    11: op1_04_inv06 = 1;
    12: op1_04_inv06 = 1;
    13: op1_04_inv06 = 1;
    14: op1_04_inv06 = 1;
    16: op1_04_inv06 = 1;
    2: op1_04_inv06 = 1;
    18: op1_04_inv06 = 1;
    20: op1_04_inv06 = 1;
    21: op1_04_inv06 = 1;
    22: op1_04_inv06 = 1;
    23: op1_04_inv06 = 1;
    25: op1_04_inv06 = 1;
    26: op1_04_inv06 = 1;
    29: op1_04_inv06 = 1;
    30: op1_04_inv06 = 1;
    31: op1_04_inv06 = 1;
    34: op1_04_inv06 = 1;
    35: op1_04_inv06 = 1;
    36: op1_04_inv06 = 1;
    37: op1_04_inv06 = 1;
    38: op1_04_inv06 = 1;
    41: op1_04_inv06 = 1;
    47: op1_04_inv06 = 1;
    48: op1_04_inv06 = 1;
    55: op1_04_inv06 = 1;
    56: op1_04_inv06 = 1;
    57: op1_04_inv06 = 1;
    58: op1_04_inv06 = 1;
    60: op1_04_inv06 = 1;
    61: op1_04_inv06 = 1;
    65: op1_04_inv06 = 1;
    66: op1_04_inv06 = 1;
    67: op1_04_inv06 = 1;
    69: op1_04_inv06 = 1;
    70: op1_04_inv06 = 1;
    71: op1_04_inv06 = 1;
    72: op1_04_inv06 = 1;
    73: op1_04_inv06 = 1;
    74: op1_04_inv06 = 1;
    78: op1_04_inv06 = 1;
    88: op1_04_inv06 = 1;
    90: op1_04_inv06 = 1;
    91: op1_04_inv06 = 1;
    92: op1_04_inv06 = 1;
    93: op1_04_inv06 = 1;
    96: op1_04_inv06 = 1;
    default: op1_04_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in07 = imem07_in[99:96];
    5: op1_04_in07 = reg_0741;
    6: op1_04_in07 = reg_0696;
    7: op1_04_in07 = reg_0554;
    8: op1_04_in07 = reg_0141;
    9: op1_04_in07 = reg_0256;
    10: op1_04_in07 = reg_0029;
    3: op1_04_in07 = reg_0427;
    11: op1_04_in07 = reg_0795;
    12: op1_04_in07 = reg_0698;
    13: op1_04_in07 = reg_0801;
    14: op1_04_in07 = reg_0140;
    15: op1_04_in07 = imem00_in[115:112];
    16: op1_04_in07 = imem02_in[123:120];
    17: op1_04_in07 = reg_0372;
    18: op1_04_in07 = reg_0589;
    19: op1_04_in07 = reg_0155;
    96: op1_04_in07 = reg_0155;
    20: op1_04_in07 = reg_0665;
    21: op1_04_in07 = reg_0089;
    57: op1_04_in07 = reg_0089;
    22: op1_04_in07 = imem07_in[95:92];
    23: op1_04_in07 = reg_0297;
    24: op1_04_in07 = reg_0679;
    25: op1_04_in07 = imem02_in[11:8];
    26: op1_04_in07 = reg_0450;
    27: op1_04_in07 = reg_0121;
    28: op1_04_in07 = reg_0390;
    29: op1_04_in07 = reg_0430;
    30: op1_04_in07 = imem02_in[67:64];
    31: op1_04_in07 = reg_0065;
    32: op1_04_in07 = reg_0338;
    33: op1_04_in07 = reg_0199;
    34: op1_04_in07 = imem06_in[67:64];
    35: op1_04_in07 = reg_0066;
    36: op1_04_in07 = reg_0232;
    37: op1_04_in07 = reg_0377;
    38: op1_04_in07 = reg_0701;
    39: op1_04_in07 = reg_0680;
    41: op1_04_in07 = reg_0499;
    42: op1_04_in07 = reg_0085;
    43: op1_04_in07 = reg_0183;
    92: op1_04_in07 = reg_0183;
    44: op1_04_in07 = reg_0125;
    86: op1_04_in07 = reg_0125;
    45: op1_04_in07 = reg_0068;
    46: op1_04_in07 = reg_0720;
    47: op1_04_in07 = reg_0686;
    48: op1_04_in07 = reg_0074;
    49: op1_04_in07 = imem03_in[27:24];
    50: op1_04_in07 = reg_0419;
    52: op1_04_in07 = reg_0687;
    53: op1_04_in07 = reg_0678;
    54: op1_04_in07 = reg_0081;
    55: op1_04_in07 = reg_0573;
    56: op1_04_in07 = imem05_in[75:72];
    58: op1_04_in07 = reg_0227;
    59: op1_04_in07 = reg_0061;
    60: op1_04_in07 = reg_0265;
    61: op1_04_in07 = reg_0437;
    62: op1_04_in07 = reg_0111;
    63: op1_04_in07 = reg_0275;
    64: op1_04_in07 = imem04_in[15:12];
    65: op1_04_in07 = imem04_in[79:76];
    66: op1_04_in07 = reg_0591;
    67: op1_04_in07 = reg_0784;
    68: op1_04_in07 = reg_0683;
    69: op1_04_in07 = reg_0587;
    70: op1_04_in07 = imem05_in[127:124];
    71: op1_04_in07 = imem02_in[35:32];
    72: op1_04_in07 = reg_0595;
    73: op1_04_in07 = reg_0262;
    74: op1_04_in07 = reg_0285;
    75: op1_04_in07 = reg_0164;
    77: op1_04_in07 = reg_0691;
    78: op1_04_in07 = reg_0350;
    79: op1_04_in07 = imem04_in[71:68];
    80: op1_04_in07 = reg_0144;
    81: op1_04_in07 = reg_0776;
    82: op1_04_in07 = reg_0684;
    83: op1_04_in07 = reg_0636;
    84: op1_04_in07 = reg_0007;
    85: op1_04_in07 = reg_0150;
    87: op1_04_in07 = imem02_in[75:72];
    88: op1_04_in07 = reg_0404;
    89: op1_04_in07 = imem03_in[31:28];
    90: op1_04_in07 = reg_0429;
    91: op1_04_in07 = reg_0292;
    93: op1_04_in07 = reg_0091;
    default: op1_04_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv07 = 1;
    7: op1_04_inv07 = 1;
    8: op1_04_inv07 = 1;
    10: op1_04_inv07 = 1;
    12: op1_04_inv07 = 1;
    15: op1_04_inv07 = 1;
    18: op1_04_inv07 = 1;
    22: op1_04_inv07 = 1;
    23: op1_04_inv07 = 1;
    25: op1_04_inv07 = 1;
    26: op1_04_inv07 = 1;
    33: op1_04_inv07 = 1;
    35: op1_04_inv07 = 1;
    38: op1_04_inv07 = 1;
    39: op1_04_inv07 = 1;
    42: op1_04_inv07 = 1;
    43: op1_04_inv07 = 1;
    44: op1_04_inv07 = 1;
    47: op1_04_inv07 = 1;
    49: op1_04_inv07 = 1;
    53: op1_04_inv07 = 1;
    54: op1_04_inv07 = 1;
    55: op1_04_inv07 = 1;
    57: op1_04_inv07 = 1;
    59: op1_04_inv07 = 1;
    64: op1_04_inv07 = 1;
    65: op1_04_inv07 = 1;
    66: op1_04_inv07 = 1;
    67: op1_04_inv07 = 1;
    68: op1_04_inv07 = 1;
    69: op1_04_inv07 = 1;
    70: op1_04_inv07 = 1;
    72: op1_04_inv07 = 1;
    74: op1_04_inv07 = 1;
    79: op1_04_inv07 = 1;
    80: op1_04_inv07 = 1;
    81: op1_04_inv07 = 1;
    86: op1_04_inv07 = 1;
    87: op1_04_inv07 = 1;
    88: op1_04_inv07 = 1;
    89: op1_04_inv07 = 1;
    91: op1_04_inv07 = 1;
    92: op1_04_inv07 = 1;
    93: op1_04_inv07 = 1;
    default: op1_04_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in08 = imem07_in[103:100];
    5: op1_04_in08 = reg_0742;
    6: op1_04_in08 = reg_0463;
    77: op1_04_in08 = reg_0463;
    7: op1_04_in08 = reg_0532;
    8: op1_04_in08 = reg_0025;
    9: op1_04_in08 = reg_0274;
    10: op1_04_in08 = imem07_in[3:0];
    3: op1_04_in08 = reg_0437;
    11: op1_04_in08 = reg_0780;
    12: op1_04_in08 = reg_0467;
    13: op1_04_in08 = reg_0799;
    14: op1_04_in08 = reg_0155;
    15: op1_04_in08 = imem00_in[127:124];
    16: op1_04_in08 = reg_0654;
    17: op1_04_in08 = reg_0392;
    18: op1_04_in08 = reg_0600;
    19: op1_04_in08 = reg_0134;
    20: op1_04_in08 = reg_0341;
    69: op1_04_in08 = reg_0341;
    21: op1_04_in08 = reg_0132;
    22: op1_04_in08 = imem07_in[107:104];
    23: op1_04_in08 = reg_0298;
    24: op1_04_in08 = reg_0677;
    25: op1_04_in08 = imem02_in[27:24];
    26: op1_04_in08 = reg_0468;
    27: op1_04_in08 = imem02_in[51:48];
    28: op1_04_in08 = reg_0380;
    29: op1_04_in08 = reg_0432;
    30: op1_04_in08 = imem02_in[71:68];
    31: op1_04_in08 = reg_0299;
    32: op1_04_in08 = reg_0371;
    33: op1_04_in08 = imem01_in[11:8];
    34: op1_04_in08 = imem06_in[75:72];
    35: op1_04_in08 = reg_0256;
    36: op1_04_in08 = reg_0774;
    37: op1_04_in08 = reg_0821;
    38: op1_04_in08 = reg_0706;
    39: op1_04_in08 = reg_0692;
    41: op1_04_in08 = reg_0396;
    42: op1_04_in08 = reg_0277;
    43: op1_04_in08 = reg_0158;
    44: op1_04_in08 = reg_0104;
    45: op1_04_in08 = reg_0227;
    46: op1_04_in08 = reg_0714;
    47: op1_04_in08 = reg_0679;
    48: op1_04_in08 = reg_0627;
    49: op1_04_in08 = imem03_in[39:36];
    50: op1_04_in08 = reg_0424;
    52: op1_04_in08 = reg_0453;
    53: op1_04_in08 = imem02_in[11:8];
    54: op1_04_in08 = reg_0095;
    55: op1_04_in08 = reg_0755;
    56: op1_04_in08 = imem05_in[79:76];
    57: op1_04_in08 = reg_0142;
    58: op1_04_in08 = reg_0482;
    59: op1_04_in08 = reg_0440;
    83: op1_04_in08 = reg_0440;
    60: op1_04_in08 = reg_0401;
    61: op1_04_in08 = reg_0182;
    62: op1_04_in08 = reg_0112;
    63: op1_04_in08 = reg_0345;
    64: op1_04_in08 = imem04_in[31:28];
    65: op1_04_in08 = reg_0542;
    66: op1_04_in08 = reg_0329;
    67: op1_04_in08 = reg_0101;
    68: op1_04_in08 = reg_0685;
    70: op1_04_in08 = reg_0781;
    71: op1_04_in08 = imem02_in[95:92];
    72: op1_04_in08 = reg_0751;
    73: op1_04_in08 = reg_0544;
    74: op1_04_in08 = reg_0812;
    78: op1_04_in08 = reg_0281;
    79: op1_04_in08 = imem04_in[99:96];
    80: op1_04_in08 = reg_0517;
    81: op1_04_in08 = imem05_in[39:36];
    82: op1_04_in08 = reg_0744;
    84: op1_04_in08 = reg_0008;
    85: op1_04_in08 = reg_0377;
    86: op1_04_in08 = reg_0670;
    87: op1_04_in08 = reg_0057;
    88: op1_04_in08 = reg_0402;
    89: op1_04_in08 = imem03_in[47:44];
    90: op1_04_in08 = reg_0433;
    91: op1_04_in08 = reg_0617;
    92: op1_04_in08 = reg_0141;
    96: op1_04_in08 = imem06_in[3:0];
    default: op1_04_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv08 = 1;
    7: op1_04_inv08 = 1;
    3: op1_04_inv08 = 1;
    14: op1_04_inv08 = 1;
    15: op1_04_inv08 = 1;
    16: op1_04_inv08 = 1;
    17: op1_04_inv08 = 1;
    18: op1_04_inv08 = 1;
    19: op1_04_inv08 = 1;
    21: op1_04_inv08 = 1;
    22: op1_04_inv08 = 1;
    23: op1_04_inv08 = 1;
    26: op1_04_inv08 = 1;
    29: op1_04_inv08 = 1;
    30: op1_04_inv08 = 1;
    34: op1_04_inv08 = 1;
    38: op1_04_inv08 = 1;
    39: op1_04_inv08 = 1;
    41: op1_04_inv08 = 1;
    43: op1_04_inv08 = 1;
    46: op1_04_inv08 = 1;
    50: op1_04_inv08 = 1;
    52: op1_04_inv08 = 1;
    54: op1_04_inv08 = 1;
    60: op1_04_inv08 = 1;
    64: op1_04_inv08 = 1;
    67: op1_04_inv08 = 1;
    74: op1_04_inv08 = 1;
    78: op1_04_inv08 = 1;
    82: op1_04_inv08 = 1;
    84: op1_04_inv08 = 1;
    85: op1_04_inv08 = 1;
    86: op1_04_inv08 = 1;
    87: op1_04_inv08 = 1;
    88: op1_04_inv08 = 1;
    90: op1_04_inv08 = 1;
    91: op1_04_inv08 = 1;
    92: op1_04_inv08 = 1;
    default: op1_04_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in09 = imem07_in[115:112];
    5: op1_04_in09 = reg_0743;
    6: op1_04_in09 = reg_0465;
    7: op1_04_in09 = reg_0559;
    8: op1_04_in09 = reg_0027;
    9: op1_04_in09 = reg_0264;
    10: op1_04_in09 = imem07_in[7:4];
    3: op1_04_in09 = reg_0180;
    11: op1_04_in09 = imem05_in[23:20];
    12: op1_04_in09 = reg_0195;
    13: op1_04_in09 = reg_0016;
    14: op1_04_in09 = imem06_in[7:4];
    15: op1_04_in09 = reg_0682;
    16: op1_04_in09 = reg_0333;
    17: op1_04_in09 = reg_0407;
    18: op1_04_in09 = reg_0360;
    19: op1_04_in09 = imem06_in[11:8];
    20: op1_04_in09 = reg_0353;
    21: op1_04_in09 = reg_0142;
    22: op1_04_in09 = imem07_in[123:120];
    23: op1_04_in09 = reg_0266;
    24: op1_04_in09 = reg_0678;
    25: op1_04_in09 = imem02_in[111:108];
    26: op1_04_in09 = reg_0189;
    27: op1_04_in09 = imem02_in[55:52];
    28: op1_04_in09 = reg_0612;
    29: op1_04_in09 = reg_0426;
    30: op1_04_in09 = imem02_in[79:76];
    31: op1_04_in09 = reg_0070;
    32: op1_04_in09 = reg_0368;
    33: op1_04_in09 = imem01_in[31:28];
    34: op1_04_in09 = imem06_in[119:116];
    35: op1_04_in09 = imem05_in[63:60];
    36: op1_04_in09 = reg_0762;
    37: op1_04_in09 = reg_0270;
    38: op1_04_in09 = reg_0727;
    39: op1_04_in09 = reg_0451;
    41: op1_04_in09 = reg_0019;
    42: op1_04_in09 = reg_0744;
    44: op1_04_in09 = reg_0106;
    45: op1_04_in09 = reg_0296;
    46: op1_04_in09 = reg_0713;
    47: op1_04_in09 = reg_0680;
    48: op1_04_in09 = reg_0626;
    49: op1_04_in09 = imem03_in[71:68];
    50: op1_04_in09 = reg_0420;
    52: op1_04_in09 = reg_0455;
    53: op1_04_in09 = imem02_in[35:32];
    54: op1_04_in09 = reg_0757;
    55: op1_04_in09 = reg_0385;
    56: op1_04_in09 = imem05_in[87:84];
    57: op1_04_in09 = reg_0146;
    58: op1_04_in09 = reg_0075;
    59: op1_04_in09 = reg_0448;
    60: op1_04_in09 = reg_0821;
    61: op1_04_in09 = reg_0160;
    62: op1_04_in09 = reg_0665;
    63: op1_04_in09 = reg_0565;
    64: op1_04_in09 = imem04_in[63:60];
    65: op1_04_in09 = reg_0088;
    66: op1_04_in09 = reg_0561;
    67: op1_04_in09 = imem05_in[19:16];
    68: op1_04_in09 = reg_0684;
    69: op1_04_in09 = reg_0092;
    70: op1_04_in09 = reg_0252;
    71: op1_04_in09 = imem02_in[99:96];
    72: op1_04_in09 = reg_0331;
    73: op1_04_in09 = reg_0553;
    74: op1_04_in09 = reg_0149;
    77: op1_04_in09 = reg_0453;
    78: op1_04_in09 = reg_0417;
    79: op1_04_in09 = imem04_in[111:108];
    80: op1_04_in09 = reg_0386;
    85: op1_04_in09 = reg_0386;
    81: op1_04_in09 = imem05_in[59:56];
    82: op1_04_in09 = reg_0749;
    83: op1_04_in09 = reg_0444;
    84: op1_04_in09 = reg_0802;
    86: op1_04_in09 = reg_0119;
    87: op1_04_in09 = reg_0081;
    88: op1_04_in09 = reg_0608;
    89: op1_04_in09 = imem03_in[75:72];
    90: op1_04_in09 = reg_0611;
    91: op1_04_in09 = reg_0610;
    92: op1_04_in09 = reg_0091;
    96: op1_04_in09 = imem06_in[19:16];
    default: op1_04_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv09 = 1;
    8: op1_04_inv09 = 1;
    10: op1_04_inv09 = 1;
    12: op1_04_inv09 = 1;
    13: op1_04_inv09 = 1;
    14: op1_04_inv09 = 1;
    15: op1_04_inv09 = 1;
    20: op1_04_inv09 = 1;
    22: op1_04_inv09 = 1;
    28: op1_04_inv09 = 1;
    31: op1_04_inv09 = 1;
    32: op1_04_inv09 = 1;
    33: op1_04_inv09 = 1;
    35: op1_04_inv09 = 1;
    36: op1_04_inv09 = 1;
    47: op1_04_inv09 = 1;
    49: op1_04_inv09 = 1;
    50: op1_04_inv09 = 1;
    53: op1_04_inv09 = 1;
    57: op1_04_inv09 = 1;
    58: op1_04_inv09 = 1;
    59: op1_04_inv09 = 1;
    60: op1_04_inv09 = 1;
    65: op1_04_inv09 = 1;
    67: op1_04_inv09 = 1;
    71: op1_04_inv09 = 1;
    77: op1_04_inv09 = 1;
    79: op1_04_inv09 = 1;
    80: op1_04_inv09 = 1;
    81: op1_04_inv09 = 1;
    83: op1_04_inv09 = 1;
    85: op1_04_inv09 = 1;
    90: op1_04_inv09 = 1;
    92: op1_04_inv09 = 1;
    96: op1_04_inv09 = 1;
    default: op1_04_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in10 = reg_0704;
    22: op1_04_in10 = reg_0704;
    5: op1_04_in10 = reg_0744;
    6: op1_04_in10 = reg_0457;
    7: op1_04_in10 = reg_0308;
    8: op1_04_in10 = reg_0219;
    9: op1_04_in10 = reg_0251;
    10: op1_04_in10 = imem07_in[75:72];
    3: op1_04_in10 = reg_0162;
    11: op1_04_in10 = imem05_in[115:112];
    56: op1_04_in10 = imem05_in[115:112];
    12: op1_04_in10 = imem01_in[11:8];
    13: op1_04_in10 = imem04_in[99:96];
    14: op1_04_in10 = imem06_in[31:28];
    15: op1_04_in10 = reg_0672;
    16: op1_04_in10 = reg_0358;
    17: op1_04_in10 = reg_0390;
    18: op1_04_in10 = reg_0370;
    19: op1_04_in10 = imem06_in[39:36];
    96: op1_04_in10 = imem06_in[39:36];
    20: op1_04_in10 = imem02_in[3:0];
    21: op1_04_in10 = reg_0146;
    23: op1_04_in10 = reg_0299;
    24: op1_04_in10 = reg_0688;
    25: op1_04_in10 = imem02_in[119:116];
    26: op1_04_in10 = reg_0190;
    27: op1_04_in10 = imem02_in[59:56];
    28: op1_04_in10 = imem06_in[15:12];
    29: op1_04_in10 = reg_0419;
    30: op1_04_in10 = imem02_in[87:84];
    31: op1_04_in10 = imem05_in[95:92];
    32: op1_04_in10 = reg_0375;
    33: op1_04_in10 = imem01_in[59:56];
    34: op1_04_in10 = reg_0628;
    35: op1_04_in10 = imem05_in[103:100];
    36: op1_04_in10 = reg_0773;
    85: op1_04_in10 = reg_0773;
    37: op1_04_in10 = reg_0403;
    38: op1_04_in10 = reg_0436;
    39: op1_04_in10 = reg_0469;
    41: op1_04_in10 = reg_0811;
    42: op1_04_in10 = reg_0285;
    44: op1_04_in10 = reg_0648;
    45: op1_04_in10 = reg_0233;
    46: op1_04_in10 = reg_0701;
    47: op1_04_in10 = reg_0699;
    48: op1_04_in10 = imem04_in[23:20];
    49: op1_04_in10 = imem03_in[83:80];
    50: op1_04_in10 = reg_0124;
    52: op1_04_in10 = reg_0460;
    53: op1_04_in10 = imem02_in[75:72];
    54: op1_04_in10 = reg_0348;
    55: op1_04_in10 = reg_0376;
    57: op1_04_in10 = reg_0143;
    58: op1_04_in10 = reg_0549;
    59: op1_04_in10 = reg_0168;
    60: op1_04_in10 = reg_0763;
    61: op1_04_in10 = reg_0184;
    62: op1_04_in10 = reg_0224;
    63: op1_04_in10 = reg_0365;
    64: op1_04_in10 = imem04_in[87:84];
    65: op1_04_in10 = reg_0500;
    66: op1_04_in10 = reg_0568;
    67: op1_04_in10 = imem05_in[23:20];
    68: op1_04_in10 = reg_0117;
    69: op1_04_in10 = reg_0541;
    70: op1_04_in10 = reg_0392;
    71: op1_04_in10 = reg_0485;
    72: op1_04_in10 = reg_0321;
    73: op1_04_in10 = reg_0043;
    74: op1_04_in10 = reg_0827;
    77: op1_04_in10 = reg_0462;
    78: op1_04_in10 = reg_0572;
    79: op1_04_in10 = reg_0262;
    80: op1_04_in10 = reg_0246;
    81: op1_04_in10 = imem05_in[119:116];
    82: op1_04_in10 = reg_0255;
    83: op1_04_in10 = reg_0442;
    84: op1_04_in10 = reg_0016;
    86: op1_04_in10 = reg_0669;
    87: op1_04_in10 = reg_0705;
    88: op1_04_in10 = reg_0593;
    89: op1_04_in10 = reg_0247;
    90: op1_04_in10 = reg_0629;
    91: op1_04_in10 = reg_0614;
    default: op1_04_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv10 = 1;
    10: op1_04_inv10 = 1;
    14: op1_04_inv10 = 1;
    15: op1_04_inv10 = 1;
    16: op1_04_inv10 = 1;
    17: op1_04_inv10 = 1;
    18: op1_04_inv10 = 1;
    20: op1_04_inv10 = 1;
    21: op1_04_inv10 = 1;
    23: op1_04_inv10 = 1;
    24: op1_04_inv10 = 1;
    25: op1_04_inv10 = 1;
    26: op1_04_inv10 = 1;
    27: op1_04_inv10 = 1;
    30: op1_04_inv10 = 1;
    32: op1_04_inv10 = 1;
    34: op1_04_inv10 = 1;
    35: op1_04_inv10 = 1;
    37: op1_04_inv10 = 1;
    38: op1_04_inv10 = 1;
    41: op1_04_inv10 = 1;
    42: op1_04_inv10 = 1;
    46: op1_04_inv10 = 1;
    49: op1_04_inv10 = 1;
    50: op1_04_inv10 = 1;
    52: op1_04_inv10 = 1;
    53: op1_04_inv10 = 1;
    56: op1_04_inv10 = 1;
    59: op1_04_inv10 = 1;
    60: op1_04_inv10 = 1;
    61: op1_04_inv10 = 1;
    62: op1_04_inv10 = 1;
    63: op1_04_inv10 = 1;
    68: op1_04_inv10 = 1;
    69: op1_04_inv10 = 1;
    70: op1_04_inv10 = 1;
    71: op1_04_inv10 = 1;
    73: op1_04_inv10 = 1;
    79: op1_04_inv10 = 1;
    83: op1_04_inv10 = 1;
    88: op1_04_inv10 = 1;
    89: op1_04_inv10 = 1;
    96: op1_04_inv10 = 1;
    default: op1_04_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in11 = reg_0717;
    5: op1_04_in11 = imem05_in[59:56];
    6: op1_04_in11 = reg_0477;
    7: op1_04_in11 = reg_0283;
    8: op1_04_in11 = reg_0613;
    9: op1_04_in11 = reg_0257;
    10: op1_04_in11 = imem07_in[87:84];
    3: op1_04_in11 = reg_0169;
    11: op1_04_in11 = reg_0132;
    12: op1_04_in11 = imem01_in[19:16];
    13: op1_04_in11 = imem04_in[111:108];
    14: op1_04_in11 = imem06_in[95:92];
    15: op1_04_in11 = reg_0461;
    16: op1_04_in11 = reg_0341;
    17: op1_04_in11 = reg_0005;
    18: op1_04_in11 = reg_0319;
    19: op1_04_in11 = imem06_in[71:68];
    96: op1_04_in11 = imem06_in[71:68];
    20: op1_04_in11 = imem02_in[19:16];
    21: op1_04_in11 = reg_0138;
    22: op1_04_in11 = reg_0719;
    23: op1_04_in11 = reg_0071;
    24: op1_04_in11 = reg_0673;
    25: op1_04_in11 = imem02_in[127:124];
    26: op1_04_in11 = imem01_in[79:76];
    27: op1_04_in11 = imem02_in[91:88];
    28: op1_04_in11 = imem06_in[39:36];
    29: op1_04_in11 = reg_0440;
    30: op1_04_in11 = imem02_in[95:92];
    53: op1_04_in11 = imem02_in[95:92];
    31: op1_04_in11 = imem05_in[111:108];
    35: op1_04_in11 = imem05_in[111:108];
    32: op1_04_in11 = reg_0779;
    33: op1_04_in11 = imem01_in[87:84];
    34: op1_04_in11 = reg_0621;
    36: op1_04_in11 = reg_0763;
    37: op1_04_in11 = reg_0406;
    38: op1_04_in11 = reg_0439;
    39: op1_04_in11 = reg_0475;
    41: op1_04_in11 = reg_0001;
    42: op1_04_in11 = reg_0136;
    44: op1_04_in11 = reg_0652;
    45: op1_04_in11 = reg_0237;
    46: op1_04_in11 = reg_0706;
    47: op1_04_in11 = reg_0450;
    48: op1_04_in11 = imem04_in[47:44];
    49: op1_04_in11 = imem03_in[91:88];
    50: op1_04_in11 = reg_0111;
    52: op1_04_in11 = reg_0456;
    54: op1_04_in11 = reg_0583;
    55: op1_04_in11 = reg_0570;
    56: op1_04_in11 = imem05_in[123:120];
    57: op1_04_in11 = reg_0139;
    58: op1_04_in11 = reg_0483;
    60: op1_04_in11 = reg_0638;
    62: op1_04_in11 = reg_0336;
    63: op1_04_in11 = reg_0527;
    64: op1_04_in11 = imem04_in[95:92];
    65: op1_04_in11 = reg_0432;
    66: op1_04_in11 = reg_0517;
    67: op1_04_in11 = imem05_in[43:40];
    68: op1_04_in11 = reg_0634;
    69: op1_04_in11 = reg_0743;
    70: op1_04_in11 = reg_0282;
    71: op1_04_in11 = reg_0359;
    72: op1_04_in11 = reg_0368;
    78: op1_04_in11 = reg_0368;
    73: op1_04_in11 = reg_0055;
    74: op1_04_in11 = reg_0151;
    77: op1_04_in11 = reg_0458;
    79: op1_04_in11 = reg_0558;
    80: op1_04_in11 = reg_0245;
    81: op1_04_in11 = reg_0135;
    82: op1_04_in11 = reg_0457;
    83: op1_04_in11 = reg_0443;
    84: op1_04_in11 = reg_0810;
    85: op1_04_in11 = reg_0632;
    86: op1_04_in11 = reg_0107;
    87: op1_04_in11 = reg_0587;
    88: op1_04_in11 = reg_0328;
    89: op1_04_in11 = reg_0536;
    90: op1_04_in11 = reg_0074;
    91: op1_04_in11 = reg_0687;
    default: op1_04_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv11 = 1;
    5: op1_04_inv11 = 1;
    8: op1_04_inv11 = 1;
    3: op1_04_inv11 = 1;
    16: op1_04_inv11 = 1;
    18: op1_04_inv11 = 1;
    20: op1_04_inv11 = 1;
    22: op1_04_inv11 = 1;
    23: op1_04_inv11 = 1;
    24: op1_04_inv11 = 1;
    26: op1_04_inv11 = 1;
    29: op1_04_inv11 = 1;
    34: op1_04_inv11 = 1;
    37: op1_04_inv11 = 1;
    45: op1_04_inv11 = 1;
    49: op1_04_inv11 = 1;
    53: op1_04_inv11 = 1;
    56: op1_04_inv11 = 1;
    63: op1_04_inv11 = 1;
    66: op1_04_inv11 = 1;
    71: op1_04_inv11 = 1;
    73: op1_04_inv11 = 1;
    74: op1_04_inv11 = 1;
    78: op1_04_inv11 = 1;
    81: op1_04_inv11 = 1;
    84: op1_04_inv11 = 1;
    85: op1_04_inv11 = 1;
    87: op1_04_inv11 = 1;
    88: op1_04_inv11 = 1;
    89: op1_04_inv11 = 1;
    90: op1_04_inv11 = 1;
    default: op1_04_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in12 = reg_0718;
    5: op1_04_in12 = imem05_in[99:96];
    6: op1_04_in12 = reg_0466;
    7: op1_04_in12 = reg_0293;
    8: op1_04_in12 = reg_0617;
    9: op1_04_in12 = reg_0272;
    10: op1_04_in12 = imem07_in[103:100];
    3: op1_04_in12 = reg_0166;
    11: op1_04_in12 = reg_0152;
    12: op1_04_in12 = imem01_in[99:96];
    13: op1_04_in12 = reg_0552;
    14: op1_04_in12 = imem06_in[115:112];
    19: op1_04_in12 = imem06_in[115:112];
    15: op1_04_in12 = reg_0469;
    16: op1_04_in12 = reg_0330;
    17: op1_04_in12 = reg_0038;
    18: op1_04_in12 = reg_0322;
    20: op1_04_in12 = imem02_in[87:84];
    21: op1_04_in12 = reg_0140;
    22: op1_04_in12 = reg_0720;
    23: op1_04_in12 = reg_0296;
    24: op1_04_in12 = reg_0461;
    25: op1_04_in12 = reg_0314;
    26: op1_04_in12 = imem01_in[107:104];
    27: op1_04_in12 = imem02_in[103:100];
    28: op1_04_in12 = imem06_in[103:100];
    29: op1_04_in12 = reg_0442;
    30: op1_04_in12 = reg_0642;
    31: op1_04_in12 = reg_0792;
    32: op1_04_in12 = imem07_in[3:0];
    33: op1_04_in12 = reg_0758;
    34: op1_04_in12 = reg_0631;
    35: op1_04_in12 = imem05_in[119:116];
    36: op1_04_in12 = reg_0404;
    37: op1_04_in12 = reg_0401;
    38: op1_04_in12 = reg_0167;
    39: op1_04_in12 = reg_0470;
    41: op1_04_in12 = reg_0002;
    42: op1_04_in12 = reg_0150;
    44: op1_04_in12 = reg_0065;
    45: op1_04_in12 = reg_0560;
    46: op1_04_in12 = reg_0061;
    47: op1_04_in12 = reg_0451;
    48: op1_04_in12 = imem04_in[63:60];
    49: op1_04_in12 = imem03_in[127:124];
    50: op1_04_in12 = reg_0116;
    52: op1_04_in12 = reg_0186;
    53: op1_04_in12 = reg_0337;
    54: op1_04_in12 = reg_0349;
    55: op1_04_in12 = reg_0006;
    56: op1_04_in12 = imem05_in[127:124];
    57: op1_04_in12 = reg_0131;
    58: op1_04_in12 = reg_0545;
    60: op1_04_in12 = reg_0035;
    62: op1_04_in12 = imem02_in[35:32];
    63: op1_04_in12 = reg_0590;
    64: op1_04_in12 = imem04_in[99:96];
    65: op1_04_in12 = reg_0283;
    66: op1_04_in12 = reg_0001;
    67: op1_04_in12 = imem05_in[47:44];
    68: op1_04_in12 = reg_0477;
    69: op1_04_in12 = reg_0531;
    70: op1_04_in12 = reg_0393;
    71: op1_04_in12 = reg_0565;
    72: op1_04_in12 = reg_0496;
    73: op1_04_in12 = reg_0083;
    74: op1_04_in12 = reg_0154;
    77: op1_04_in12 = reg_0200;
    78: op1_04_in12 = reg_0372;
    79: op1_04_in12 = reg_0556;
    80: op1_04_in12 = reg_0735;
    81: op1_04_in12 = reg_0128;
    82: op1_04_in12 = reg_0476;
    83: op1_04_in12 = reg_0448;
    84: op1_04_in12 = imem04_in[15:12];
    85: op1_04_in12 = reg_0764;
    86: op1_04_in12 = reg_0678;
    87: op1_04_in12 = reg_0586;
    88: op1_04_in12 = reg_0512;
    89: op1_04_in12 = reg_0523;
    90: op1_04_in12 = reg_0311;
    91: op1_04_in12 = reg_0598;
    96: op1_04_in12 = imem06_in[91:88];
    default: op1_04_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv12 = 1;
    6: op1_04_inv12 = 1;
    7: op1_04_inv12 = 1;
    8: op1_04_inv12 = 1;
    9: op1_04_inv12 = 1;
    3: op1_04_inv12 = 1;
    11: op1_04_inv12 = 1;
    14: op1_04_inv12 = 1;
    16: op1_04_inv12 = 1;
    17: op1_04_inv12 = 1;
    18: op1_04_inv12 = 1;
    20: op1_04_inv12 = 1;
    21: op1_04_inv12 = 1;
    25: op1_04_inv12 = 1;
    28: op1_04_inv12 = 1;
    34: op1_04_inv12 = 1;
    35: op1_04_inv12 = 1;
    37: op1_04_inv12 = 1;
    41: op1_04_inv12 = 1;
    42: op1_04_inv12 = 1;
    44: op1_04_inv12 = 1;
    45: op1_04_inv12 = 1;
    47: op1_04_inv12 = 1;
    49: op1_04_inv12 = 1;
    53: op1_04_inv12 = 1;
    54: op1_04_inv12 = 1;
    55: op1_04_inv12 = 1;
    57: op1_04_inv12 = 1;
    60: op1_04_inv12 = 1;
    62: op1_04_inv12 = 1;
    64: op1_04_inv12 = 1;
    65: op1_04_inv12 = 1;
    70: op1_04_inv12 = 1;
    71: op1_04_inv12 = 1;
    72: op1_04_inv12 = 1;
    73: op1_04_inv12 = 1;
    78: op1_04_inv12 = 1;
    79: op1_04_inv12 = 1;
    81: op1_04_inv12 = 1;
    82: op1_04_inv12 = 1;
    87: op1_04_inv12 = 1;
    88: op1_04_inv12 = 1;
    89: op1_04_inv12 = 1;
    91: op1_04_inv12 = 1;
    default: op1_04_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in13 = reg_0706;
    5: op1_04_in13 = reg_0267;
    6: op1_04_in13 = reg_0474;
    7: op1_04_in13 = reg_0046;
    8: op1_04_in13 = reg_0606;
    9: op1_04_in13 = reg_0261;
    10: op1_04_in13 = reg_0704;
    3: op1_04_in13 = reg_0185;
    11: op1_04_in13 = reg_0153;
    12: op1_04_in13 = imem01_in[115:112];
    13: op1_04_in13 = reg_0555;
    14: op1_04_in13 = reg_0630;
    15: op1_04_in13 = reg_0472;
    16: op1_04_in13 = reg_0363;
    17: op1_04_in13 = imem07_in[75:72];
    18: op1_04_in13 = reg_0396;
    19: op1_04_in13 = imem06_in[119:116];
    20: op1_04_in13 = imem03_in[7:4];
    21: op1_04_in13 = imem06_in[35:32];
    22: op1_04_in13 = reg_0730;
    23: op1_04_in13 = imem05_in[39:36];
    24: op1_04_in13 = reg_0462;
    82: op1_04_in13 = reg_0462;
    25: op1_04_in13 = reg_0533;
    26: op1_04_in13 = reg_0501;
    27: op1_04_in13 = reg_0650;
    30: op1_04_in13 = reg_0650;
    28: op1_04_in13 = imem06_in[107:104];
    29: op1_04_in13 = reg_0180;
    31: op1_04_in13 = reg_0796;
    32: op1_04_in13 = imem07_in[23:20];
    33: op1_04_in13 = reg_0820;
    34: op1_04_in13 = reg_0626;
    35: op1_04_in13 = reg_0788;
    81: op1_04_in13 = reg_0788;
    36: op1_04_in13 = reg_0329;
    37: op1_04_in13 = reg_0028;
    39: op1_04_in13 = reg_0468;
    41: op1_04_in13 = reg_0805;
    42: op1_04_in13 = reg_0152;
    44: op1_04_in13 = imem02_in[63:60];
    45: op1_04_in13 = reg_0328;
    46: op1_04_in13 = reg_0442;
    47: op1_04_in13 = reg_0455;
    48: op1_04_in13 = imem04_in[75:72];
    49: op1_04_in13 = reg_0259;
    56: op1_04_in13 = reg_0259;
    50: op1_04_in13 = reg_0115;
    85: op1_04_in13 = reg_0115;
    52: op1_04_in13 = reg_0199;
    53: op1_04_in13 = reg_0656;
    54: op1_04_in13 = reg_0354;
    55: op1_04_in13 = reg_0007;
    57: op1_04_in13 = reg_0144;
    58: op1_04_in13 = reg_0087;
    60: op1_04_in13 = reg_0512;
    62: op1_04_in13 = imem02_in[47:44];
    63: op1_04_in13 = reg_0343;
    64: op1_04_in13 = reg_0547;
    65: op1_04_in13 = reg_0297;
    66: op1_04_in13 = reg_0801;
    67: op1_04_in13 = imem05_in[51:48];
    68: op1_04_in13 = reg_0459;
    69: op1_04_in13 = reg_0740;
    70: op1_04_in13 = reg_0277;
    71: op1_04_in13 = reg_0414;
    72: op1_04_in13 = reg_0387;
    73: op1_04_in13 = reg_0611;
    74: op1_04_in13 = reg_0137;
    77: op1_04_in13 = reg_0193;
    78: op1_04_in13 = reg_0646;
    79: op1_04_in13 = reg_0077;
    80: op1_04_in13 = reg_0229;
    83: op1_04_in13 = reg_0268;
    84: op1_04_in13 = imem04_in[19:16];
    86: op1_04_in13 = imem02_in[3:0];
    87: op1_04_in13 = reg_0566;
    88: op1_04_in13 = imem06_in[63:60];
    89: op1_04_in13 = reg_0331;
    90: op1_04_in13 = reg_0371;
    91: op1_04_in13 = reg_0771;
    96: op1_04_in13 = imem06_in[111:108];
    default: op1_04_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv13 = 1;
    5: op1_04_inv13 = 1;
    6: op1_04_inv13 = 1;
    7: op1_04_inv13 = 1;
    8: op1_04_inv13 = 1;
    10: op1_04_inv13 = 1;
    12: op1_04_inv13 = 1;
    14: op1_04_inv13 = 1;
    17: op1_04_inv13 = 1;
    18: op1_04_inv13 = 1;
    19: op1_04_inv13 = 1;
    20: op1_04_inv13 = 1;
    21: op1_04_inv13 = 1;
    22: op1_04_inv13 = 1;
    23: op1_04_inv13 = 1;
    24: op1_04_inv13 = 1;
    25: op1_04_inv13 = 1;
    27: op1_04_inv13 = 1;
    29: op1_04_inv13 = 1;
    30: op1_04_inv13 = 1;
    31: op1_04_inv13 = 1;
    32: op1_04_inv13 = 1;
    41: op1_04_inv13 = 1;
    42: op1_04_inv13 = 1;
    45: op1_04_inv13 = 1;
    47: op1_04_inv13 = 1;
    53: op1_04_inv13 = 1;
    56: op1_04_inv13 = 1;
    63: op1_04_inv13 = 1;
    65: op1_04_inv13 = 1;
    66: op1_04_inv13 = 1;
    68: op1_04_inv13 = 1;
    71: op1_04_inv13 = 1;
    72: op1_04_inv13 = 1;
    73: op1_04_inv13 = 1;
    74: op1_04_inv13 = 1;
    77: op1_04_inv13 = 1;
    82: op1_04_inv13 = 1;
    83: op1_04_inv13 = 1;
    84: op1_04_inv13 = 1;
    85: op1_04_inv13 = 1;
    86: op1_04_inv13 = 1;
    96: op1_04_inv13 = 1;
    default: op1_04_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in14 = reg_0423;
    5: op1_04_in14 = reg_0268;
    6: op1_04_in14 = reg_0471;
    15: op1_04_in14 = reg_0471;
    7: op1_04_in14 = reg_0054;
    8: op1_04_in14 = reg_0577;
    9: op1_04_in14 = reg_0253;
    10: op1_04_in14 = reg_0719;
    3: op1_04_in14 = reg_0173;
    11: op1_04_in14 = reg_0130;
    12: op1_04_in14 = reg_0523;
    13: op1_04_in14 = reg_0547;
    14: op1_04_in14 = reg_0626;
    16: op1_04_in14 = reg_0092;
    17: op1_04_in14 = imem07_in[115:112];
    18: op1_04_in14 = reg_0803;
    19: op1_04_in14 = reg_0614;
    20: op1_04_in14 = imem03_in[27:24];
    21: op1_04_in14 = imem06_in[47:44];
    22: op1_04_in14 = reg_0723;
    23: op1_04_in14 = imem05_in[75:72];
    24: op1_04_in14 = reg_0480;
    25: op1_04_in14 = reg_0531;
    63: op1_04_in14 = reg_0531;
    26: op1_04_in14 = reg_0496;
    27: op1_04_in14 = reg_0645;
    28: op1_04_in14 = imem06_in[111:108];
    29: op1_04_in14 = reg_0163;
    30: op1_04_in14 = reg_0666;
    31: op1_04_in14 = reg_0490;
    32: op1_04_in14 = imem07_in[51:48];
    33: op1_04_in14 = reg_0334;
    34: op1_04_in14 = reg_0622;
    35: op1_04_in14 = reg_0789;
    36: op1_04_in14 = reg_0319;
    37: op1_04_in14 = reg_0031;
    39: op1_04_in14 = reg_0213;
    41: op1_04_in14 = reg_0806;
    42: op1_04_in14 = reg_0153;
    44: op1_04_in14 = imem02_in[99:96];
    45: op1_04_in14 = reg_0087;
    46: op1_04_in14 = reg_0175;
    47: op1_04_in14 = reg_0472;
    48: op1_04_in14 = imem04_in[115:112];
    49: op1_04_in14 = reg_0587;
    50: op1_04_in14 = reg_0110;
    52: op1_04_in14 = reg_0110;
    56: op1_04_in14 = reg_0110;
    53: op1_04_in14 = reg_0548;
    54: op1_04_in14 = reg_0593;
    55: op1_04_in14 = reg_0801;
    57: op1_04_in14 = reg_0062;
    58: op1_04_in14 = reg_0510;
    60: op1_04_in14 = imem06_in[11:8];
    62: op1_04_in14 = imem02_in[95:92];
    64: op1_04_in14 = reg_0429;
    65: op1_04_in14 = reg_0292;
    66: op1_04_in14 = reg_0014;
    67: op1_04_in14 = reg_0245;
    68: op1_04_in14 = reg_0214;
    69: op1_04_in14 = reg_0532;
    70: op1_04_in14 = reg_0257;
    71: op1_04_in14 = reg_0590;
    72: op1_04_in14 = reg_0000;
    73: op1_04_in14 = reg_0077;
    74: op1_04_in14 = reg_0734;
    77: op1_04_in14 = reg_0186;
    78: op1_04_in14 = reg_0562;
    79: op1_04_in14 = reg_0616;
    80: op1_04_in14 = reg_0276;
    81: op1_04_in14 = reg_0090;
    82: op1_04_in14 = reg_0474;
    83: op1_04_in14 = reg_0116;
    84: op1_04_in14 = imem04_in[23:20];
    85: op1_04_in14 = reg_0609;
    86: op1_04_in14 = imem02_in[11:8];
    87: op1_04_in14 = reg_0030;
    88: op1_04_in14 = imem06_in[75:72];
    89: op1_04_in14 = reg_0249;
    90: op1_04_in14 = reg_0640;
    91: op1_04_in14 = reg_0233;
    96: op1_04_in14 = reg_0605;
    default: op1_04_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv14 = 1;
    9: op1_04_inv14 = 1;
    10: op1_04_inv14 = 1;
    3: op1_04_inv14 = 1;
    11: op1_04_inv14 = 1;
    12: op1_04_inv14 = 1;
    13: op1_04_inv14 = 1;
    15: op1_04_inv14 = 1;
    17: op1_04_inv14 = 1;
    20: op1_04_inv14 = 1;
    21: op1_04_inv14 = 1;
    24: op1_04_inv14 = 1;
    25: op1_04_inv14 = 1;
    32: op1_04_inv14 = 1;
    33: op1_04_inv14 = 1;
    35: op1_04_inv14 = 1;
    36: op1_04_inv14 = 1;
    37: op1_04_inv14 = 1;
    41: op1_04_inv14 = 1;
    45: op1_04_inv14 = 1;
    46: op1_04_inv14 = 1;
    48: op1_04_inv14 = 1;
    49: op1_04_inv14 = 1;
    50: op1_04_inv14 = 1;
    53: op1_04_inv14 = 1;
    55: op1_04_inv14 = 1;
    57: op1_04_inv14 = 1;
    58: op1_04_inv14 = 1;
    62: op1_04_inv14 = 1;
    64: op1_04_inv14 = 1;
    67: op1_04_inv14 = 1;
    69: op1_04_inv14 = 1;
    73: op1_04_inv14 = 1;
    74: op1_04_inv14 = 1;
    77: op1_04_inv14 = 1;
    78: op1_04_inv14 = 1;
    80: op1_04_inv14 = 1;
    82: op1_04_inv14 = 1;
    84: op1_04_inv14 = 1;
    85: op1_04_inv14 = 1;
    86: op1_04_inv14 = 1;
    87: op1_04_inv14 = 1;
    89: op1_04_inv14 = 1;
    96: op1_04_inv14 = 1;
    default: op1_04_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in15 = reg_0180;
    5: op1_04_in15 = reg_0252;
    6: op1_04_in15 = reg_0478;
    7: op1_04_in15 = reg_0067;
    8: op1_04_in15 = reg_0402;
    9: op1_04_in15 = reg_0132;
    10: op1_04_in15 = reg_0726;
    3: op1_04_in15 = reg_0184;
    11: op1_04_in15 = reg_0155;
    12: op1_04_in15 = reg_0227;
    13: op1_04_in15 = reg_0308;
    89: op1_04_in15 = reg_0308;
    14: op1_04_in15 = reg_0349;
    44: op1_04_in15 = reg_0349;
    15: op1_04_in15 = reg_0458;
    16: op1_04_in15 = reg_0084;
    17: op1_04_in15 = reg_0714;
    18: op1_04_in15 = reg_0809;
    19: op1_04_in15 = reg_0617;
    20: op1_04_in15 = imem03_in[107:104];
    21: op1_04_in15 = imem06_in[119:116];
    22: op1_04_in15 = reg_0700;
    23: op1_04_in15 = imem05_in[103:100];
    24: op1_04_in15 = reg_0471;
    25: op1_04_in15 = reg_0498;
    26: op1_04_in15 = reg_0514;
    27: op1_04_in15 = reg_0655;
    28: op1_04_in15 = reg_0039;
    29: op1_04_in15 = reg_0185;
    30: op1_04_in15 = reg_0639;
    31: op1_04_in15 = reg_0789;
    32: op1_04_in15 = imem07_in[63:60];
    33: op1_04_in15 = reg_0825;
    34: op1_04_in15 = reg_0762;
    35: op1_04_in15 = reg_0492;
    36: op1_04_in15 = reg_0038;
    37: op1_04_in15 = reg_0037;
    39: op1_04_in15 = reg_0196;
    41: op1_04_in15 = reg_0810;
    42: op1_04_in15 = imem06_in[67:64];
    45: op1_04_in15 = reg_0542;
    46: op1_04_in15 = reg_0172;
    47: op1_04_in15 = reg_0480;
    48: op1_04_in15 = imem05_in[15:12];
    49: op1_04_in15 = reg_0594;
    50: op1_04_in15 = imem02_in[51:48];
    52: op1_04_in15 = reg_0114;
    53: op1_04_in15 = reg_0362;
    54: op1_04_in15 = reg_0580;
    55: op1_04_in15 = reg_0014;
    56: op1_04_in15 = reg_0270;
    57: op1_04_in15 = reg_0286;
    58: op1_04_in15 = reg_0516;
    60: op1_04_in15 = imem06_in[27:24];
    62: op1_04_in15 = imem02_in[103:100];
    63: op1_04_in15 = reg_0093;
    64: op1_04_in15 = reg_0076;
    65: op1_04_in15 = reg_0508;
    66: op1_04_in15 = reg_0799;
    67: op1_04_in15 = reg_0276;
    68: op1_04_in15 = reg_0208;
    69: op1_04_in15 = reg_0070;
    70: op1_04_in15 = reg_0285;
    71: op1_04_in15 = reg_0743;
    72: op1_04_in15 = reg_0006;
    73: op1_04_in15 = reg_0297;
    74: op1_04_in15 = imem06_in[23:20];
    77: op1_04_in15 = reg_0194;
    78: op1_04_in15 = reg_0637;
    79: op1_04_in15 = reg_0431;
    80: op1_04_in15 = reg_0138;
    81: op1_04_in15 = reg_0027;
    82: op1_04_in15 = reg_0209;
    83: op1_04_in15 = reg_0181;
    84: op1_04_in15 = imem04_in[35:32];
    85: op1_04_in15 = reg_0606;
    86: op1_04_in15 = imem02_in[47:44];
    87: op1_04_in15 = reg_0096;
    88: op1_04_in15 = imem06_in[115:112];
    90: op1_04_in15 = reg_0416;
    91: op1_04_in15 = imem05_in[43:40];
    96: op1_04_in15 = reg_0298;
    default: op1_04_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv15 = 1;
    8: op1_04_inv15 = 1;
    9: op1_04_inv15 = 1;
    10: op1_04_inv15 = 1;
    12: op1_04_inv15 = 1;
    13: op1_04_inv15 = 1;
    19: op1_04_inv15 = 1;
    20: op1_04_inv15 = 1;
    24: op1_04_inv15 = 1;
    25: op1_04_inv15 = 1;
    27: op1_04_inv15 = 1;
    28: op1_04_inv15 = 1;
    30: op1_04_inv15 = 1;
    31: op1_04_inv15 = 1;
    32: op1_04_inv15 = 1;
    33: op1_04_inv15 = 1;
    34: op1_04_inv15 = 1;
    46: op1_04_inv15 = 1;
    47: op1_04_inv15 = 1;
    48: op1_04_inv15 = 1;
    49: op1_04_inv15 = 1;
    50: op1_04_inv15 = 1;
    52: op1_04_inv15 = 1;
    53: op1_04_inv15 = 1;
    54: op1_04_inv15 = 1;
    58: op1_04_inv15 = 1;
    60: op1_04_inv15 = 1;
    62: op1_04_inv15 = 1;
    63: op1_04_inv15 = 1;
    64: op1_04_inv15 = 1;
    66: op1_04_inv15 = 1;
    67: op1_04_inv15 = 1;
    69: op1_04_inv15 = 1;
    70: op1_04_inv15 = 1;
    71: op1_04_inv15 = 1;
    72: op1_04_inv15 = 1;
    73: op1_04_inv15 = 1;
    74: op1_04_inv15 = 1;
    77: op1_04_inv15 = 1;
    78: op1_04_inv15 = 1;
    80: op1_04_inv15 = 1;
    81: op1_04_inv15 = 1;
    83: op1_04_inv15 = 1;
    84: op1_04_inv15 = 1;
    86: op1_04_inv15 = 1;
    87: op1_04_inv15 = 1;
    89: op1_04_inv15 = 1;
    90: op1_04_inv15 = 1;
    91: op1_04_inv15 = 1;
    default: op1_04_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in16 = reg_0166;
    5: op1_04_in16 = reg_0243;
    6: op1_04_in16 = reg_0210;
    15: op1_04_in16 = reg_0210;
    7: op1_04_in16 = reg_0043;
    8: op1_04_in16 = reg_0372;
    9: op1_04_in16 = reg_0147;
    10: op1_04_in16 = reg_0713;
    11: op1_04_in16 = reg_0144;
    12: op1_04_in16 = reg_0505;
    13: op1_04_in16 = reg_0301;
    14: op1_04_in16 = reg_0407;
    16: op1_04_in16 = reg_0073;
    17: op1_04_in16 = reg_0709;
    18: op1_04_in16 = reg_0056;
    19: op1_04_in16 = reg_0615;
    20: op1_04_in16 = reg_0598;
    21: op1_04_in16 = reg_0610;
    73: op1_04_in16 = reg_0610;
    22: op1_04_in16 = reg_0727;
    23: op1_04_in16 = reg_0483;
    24: op1_04_in16 = reg_0458;
    25: op1_04_in16 = imem03_in[15:12];
    26: op1_04_in16 = reg_0559;
    27: op1_04_in16 = reg_0661;
    28: op1_04_in16 = reg_0040;
    29: op1_04_in16 = reg_0168;
    30: op1_04_in16 = reg_0652;
    31: op1_04_in16 = reg_0795;
    32: op1_04_in16 = imem07_in[71:68];
    33: op1_04_in16 = reg_0759;
    34: op1_04_in16 = reg_0763;
    35: op1_04_in16 = reg_0790;
    36: op1_04_in16 = reg_0576;
    37: op1_04_in16 = reg_0238;
    39: op1_04_in16 = reg_0054;
    41: op1_04_in16 = reg_0267;
    42: op1_04_in16 = reg_0289;
    44: op1_04_in16 = reg_0364;
    45: op1_04_in16 = reg_0060;
    46: op1_04_in16 = reg_0159;
    47: op1_04_in16 = reg_0468;
    48: op1_04_in16 = imem05_in[23:20];
    49: op1_04_in16 = reg_0581;
    50: op1_04_in16 = reg_0639;
    52: op1_04_in16 = reg_0824;
    53: op1_04_in16 = reg_0341;
    54: op1_04_in16 = imem03_in[51:48];
    55: op1_04_in16 = reg_0016;
    56: op1_04_in16 = reg_0788;
    57: op1_04_in16 = reg_0068;
    58: op1_04_in16 = reg_0303;
    60: op1_04_in16 = imem06_in[63:60];
    62: op1_04_in16 = imem02_in[111:108];
    63: op1_04_in16 = reg_0532;
    64: op1_04_in16 = reg_0529;
    65: op1_04_in16 = reg_0617;
    66: op1_04_in16 = reg_0010;
    67: op1_04_in16 = reg_0149;
    68: op1_04_in16 = reg_0211;
    69: op1_04_in16 = reg_0090;
    70: op1_04_in16 = reg_0486;
    71: op1_04_in16 = reg_0095;
    72: op1_04_in16 = reg_0806;
    74: op1_04_in16 = imem06_in[59:56];
    77: op1_04_in16 = reg_0190;
    78: op1_04_in16 = reg_0623;
    79: op1_04_in16 = reg_0508;
    80: op1_04_in16 = reg_0719;
    81: op1_04_in16 = reg_0732;
    82: op1_04_in16 = reg_0213;
    83: op1_04_in16 = reg_0236;
    84: op1_04_in16 = imem04_in[43:40];
    85: op1_04_in16 = reg_0766;
    86: op1_04_in16 = imem02_in[59:56];
    87: op1_04_in16 = reg_0136;
    88: op1_04_in16 = imem07_in[31:28];
    89: op1_04_in16 = reg_0283;
    90: op1_04_in16 = imem05_in[7:4];
    91: op1_04_in16 = imem05_in[51:48];
    96: op1_04_in16 = reg_0404;
    default: op1_04_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_04_inv16 = 1;
    7: op1_04_inv16 = 1;
    8: op1_04_inv16 = 1;
    9: op1_04_inv16 = 1;
    10: op1_04_inv16 = 1;
    11: op1_04_inv16 = 1;
    12: op1_04_inv16 = 1;
    14: op1_04_inv16 = 1;
    15: op1_04_inv16 = 1;
    16: op1_04_inv16 = 1;
    18: op1_04_inv16 = 1;
    20: op1_04_inv16 = 1;
    22: op1_04_inv16 = 1;
    25: op1_04_inv16 = 1;
    27: op1_04_inv16 = 1;
    28: op1_04_inv16 = 1;
    29: op1_04_inv16 = 1;
    30: op1_04_inv16 = 1;
    33: op1_04_inv16 = 1;
    34: op1_04_inv16 = 1;
    35: op1_04_inv16 = 1;
    36: op1_04_inv16 = 1;
    37: op1_04_inv16 = 1;
    42: op1_04_inv16 = 1;
    45: op1_04_inv16 = 1;
    46: op1_04_inv16 = 1;
    50: op1_04_inv16 = 1;
    56: op1_04_inv16 = 1;
    57: op1_04_inv16 = 1;
    58: op1_04_inv16 = 1;
    62: op1_04_inv16 = 1;
    63: op1_04_inv16 = 1;
    65: op1_04_inv16 = 1;
    67: op1_04_inv16 = 1;
    70: op1_04_inv16 = 1;
    71: op1_04_inv16 = 1;
    72: op1_04_inv16 = 1;
    74: op1_04_inv16 = 1;
    78: op1_04_inv16 = 1;
    82: op1_04_inv16 = 1;
    83: op1_04_inv16 = 1;
    85: op1_04_inv16 = 1;
    88: op1_04_inv16 = 1;
    90: op1_04_inv16 = 1;
    91: op1_04_inv16 = 1;
    default: op1_04_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_04_in17 = reg_0168;
    5: op1_04_in17 = reg_0269;
    6: op1_04_in17 = reg_0203;
    7: op1_04_in17 = reg_0068;
    8: op1_04_in17 = reg_0408;
    9: op1_04_in17 = reg_0148;
    10: op1_04_in17 = reg_0711;
    11: op1_04_in17 = imem06_in[3:0];
    12: op1_04_in17 = reg_0246;
    13: op1_04_in17 = reg_0283;
    14: op1_04_in17 = reg_0405;
    15: op1_04_in17 = reg_0187;
    47: op1_04_in17 = reg_0187;
    16: op1_04_in17 = imem03_in[3:0];
    17: op1_04_in17 = reg_0715;
    18: op1_04_in17 = reg_0055;
    19: op1_04_in17 = reg_0349;
    20: op1_04_in17 = reg_0573;
    21: op1_04_in17 = reg_0617;
    22: op1_04_in17 = reg_0424;
    23: op1_04_in17 = reg_0488;
    24: op1_04_in17 = reg_0200;
    25: op1_04_in17 = imem03_in[23:20];
    26: op1_04_in17 = reg_0235;
    27: op1_04_in17 = reg_0656;
    28: op1_04_in17 = reg_0819;
    29: op1_04_in17 = reg_0158;
    30: op1_04_in17 = reg_0663;
    31: op1_04_in17 = reg_0793;
    32: op1_04_in17 = imem07_in[123:120];
    33: op1_04_in17 = reg_0771;
    34: op1_04_in17 = reg_0270;
    35: op1_04_in17 = reg_0784;
    36: op1_04_in17 = imem06_in[15:12];
    85: op1_04_in17 = imem06_in[15:12];
    37: op1_04_in17 = reg_0029;
    39: op1_04_in17 = reg_0233;
    41: op1_04_in17 = reg_0266;
    42: op1_04_in17 = reg_0218;
    44: op1_04_in17 = reg_0359;
    45: op1_04_in17 = reg_0510;
    46: op1_04_in17 = reg_0169;
    48: op1_04_in17 = imem05_in[27:24];
    49: op1_04_in17 = reg_0749;
    50: op1_04_in17 = reg_0651;
    52: op1_04_in17 = reg_0116;
    53: op1_04_in17 = reg_0360;
    54: op1_04_in17 = imem03_in[59:56];
    55: op1_04_in17 = imem04_in[23:20];
    56: op1_04_in17 = reg_0795;
    57: op1_04_in17 = reg_0624;
    58: op1_04_in17 = reg_0432;
    60: op1_04_in17 = imem06_in[71:68];
    62: op1_04_in17 = reg_0362;
    63: op1_04_in17 = imem03_in[79:76];
    64: op1_04_in17 = reg_0071;
    65: op1_04_in17 = reg_0598;
    66: op1_04_in17 = imem04_in[7:4];
    67: op1_04_in17 = reg_0142;
    83: op1_04_in17 = reg_0142;
    68: op1_04_in17 = reg_0206;
    69: op1_04_in17 = reg_0599;
    70: op1_04_in17 = reg_0143;
    71: op1_04_in17 = reg_0530;
    72: op1_04_in17 = reg_0009;
    73: op1_04_in17 = reg_0223;
    74: op1_04_in17 = imem06_in[87:84];
    77: op1_04_in17 = imem01_in[39:36];
    78: op1_04_in17 = reg_0003;
    79: op1_04_in17 = reg_0065;
    80: op1_04_in17 = reg_0742;
    81: op1_04_in17 = reg_0486;
    82: op1_04_in17 = imem01_in[43:40];
    84: op1_04_in17 = imem04_in[91:88];
    86: op1_04_in17 = reg_0088;
    87: op1_04_in17 = reg_0756;
    88: op1_04_in17 = imem07_in[51:48];
    89: op1_04_in17 = reg_0077;
    90: op1_04_in17 = imem05_in[59:56];
    91: op1_04_in17 = imem05_in[103:100];
    96: op1_04_in17 = reg_0339;
    default: op1_04_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv17 = 1;
    7: op1_04_inv17 = 1;
    8: op1_04_inv17 = 1;
    10: op1_04_inv17 = 1;
    13: op1_04_inv17 = 1;
    15: op1_04_inv17 = 1;
    16: op1_04_inv17 = 1;
    18: op1_04_inv17 = 1;
    21: op1_04_inv17 = 1;
    23: op1_04_inv17 = 1;
    24: op1_04_inv17 = 1;
    26: op1_04_inv17 = 1;
    27: op1_04_inv17 = 1;
    30: op1_04_inv17 = 1;
    33: op1_04_inv17 = 1;
    34: op1_04_inv17 = 1;
    39: op1_04_inv17 = 1;
    44: op1_04_inv17 = 1;
    46: op1_04_inv17 = 1;
    47: op1_04_inv17 = 1;
    48: op1_04_inv17 = 1;
    50: op1_04_inv17 = 1;
    53: op1_04_inv17 = 1;
    54: op1_04_inv17 = 1;
    55: op1_04_inv17 = 1;
    56: op1_04_inv17 = 1;
    57: op1_04_inv17 = 1;
    62: op1_04_inv17 = 1;
    63: op1_04_inv17 = 1;
    65: op1_04_inv17 = 1;
    68: op1_04_inv17 = 1;
    74: op1_04_inv17 = 1;
    78: op1_04_inv17 = 1;
    81: op1_04_inv17 = 1;
    82: op1_04_inv17 = 1;
    85: op1_04_inv17 = 1;
    88: op1_04_inv17 = 1;
    89: op1_04_inv17 = 1;
    91: op1_04_inv17 = 1;
    96: op1_04_inv17 = 1;
    default: op1_04_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in18 = reg_0244;
    6: op1_04_in18 = reg_0186;
    7: op1_04_in18 = reg_0075;
    8: op1_04_in18 = reg_0392;
    9: op1_04_in18 = reg_0145;
    10: op1_04_in18 = reg_0424;
    11: op1_04_in18 = imem06_in[7:4];
    12: op1_04_in18 = reg_0041;
    13: op1_04_in18 = reg_0279;
    14: op1_04_in18 = reg_0375;
    19: op1_04_in18 = reg_0375;
    15: op1_04_in18 = reg_0193;
    16: op1_04_in18 = imem03_in[19:16];
    17: op1_04_in18 = reg_0707;
    18: op1_04_in18 = reg_0276;
    20: op1_04_in18 = reg_0568;
    21: op1_04_in18 = reg_0605;
    57: op1_04_in18 = reg_0605;
    22: op1_04_in18 = reg_0430;
    23: op1_04_in18 = reg_0741;
    24: op1_04_in18 = reg_0204;
    47: op1_04_in18 = reg_0204;
    25: op1_04_in18 = imem03_in[47:44];
    26: op1_04_in18 = reg_0215;
    33: op1_04_in18 = reg_0215;
    27: op1_04_in18 = reg_0651;
    28: op1_04_in18 = imem07_in[23:20];
    37: op1_04_in18 = imem07_in[23:20];
    30: op1_04_in18 = reg_0540;
    71: op1_04_in18 = reg_0540;
    31: op1_04_in18 = reg_0309;
    32: op1_04_in18 = reg_0719;
    34: op1_04_in18 = reg_0038;
    35: op1_04_in18 = reg_0486;
    36: op1_04_in18 = imem06_in[63:60];
    39: op1_04_in18 = reg_0237;
    41: op1_04_in18 = reg_0053;
    42: op1_04_in18 = reg_0020;
    44: op1_04_in18 = reg_0361;
    45: op1_04_in18 = reg_0283;
    46: op1_04_in18 = reg_0163;
    48: op1_04_in18 = imem05_in[43:40];
    49: op1_04_in18 = reg_0387;
    54: op1_04_in18 = reg_0387;
    50: op1_04_in18 = reg_0301;
    52: op1_04_in18 = reg_0115;
    53: op1_04_in18 = reg_0594;
    55: op1_04_in18 = imem04_in[35:32];
    56: op1_04_in18 = reg_0790;
    58: op1_04_in18 = reg_0631;
    60: op1_04_in18 = imem07_in[19:16];
    62: op1_04_in18 = reg_0360;
    63: op1_04_in18 = reg_0338;
    69: op1_04_in18 = reg_0338;
    64: op1_04_in18 = reg_0503;
    65: op1_04_in18 = reg_0622;
    66: op1_04_in18 = imem04_in[51:48];
    67: op1_04_in18 = reg_0146;
    68: op1_04_in18 = reg_0199;
    70: op1_04_in18 = reg_0139;
    72: op1_04_in18 = imem04_in[7:4];
    73: op1_04_in18 = reg_0078;
    74: op1_04_in18 = reg_0298;
    77: op1_04_in18 = imem01_in[55:52];
    82: op1_04_in18 = imem01_in[55:52];
    78: op1_04_in18 = reg_0013;
    79: op1_04_in18 = reg_0371;
    80: op1_04_in18 = reg_0830;
    81: op1_04_in18 = reg_0500;
    83: op1_04_in18 = reg_0327;
    84: op1_04_in18 = imem04_in[95:92];
    85: op1_04_in18 = imem06_in[23:20];
    86: op1_04_in18 = reg_0533;
    87: op1_04_in18 = reg_0063;
    88: op1_04_in18 = reg_0725;
    89: op1_04_in18 = reg_0626;
    90: op1_04_in18 = imem05_in[63:60];
    91: op1_04_in18 = reg_0133;
    96: op1_04_in18 = reg_0628;
    default: op1_04_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv18 = 1;
    8: op1_04_inv18 = 1;
    9: op1_04_inv18 = 1;
    12: op1_04_inv18 = 1;
    16: op1_04_inv18 = 1;
    18: op1_04_inv18 = 1;
    21: op1_04_inv18 = 1;
    26: op1_04_inv18 = 1;
    34: op1_04_inv18 = 1;
    37: op1_04_inv18 = 1;
    42: op1_04_inv18 = 1;
    45: op1_04_inv18 = 1;
    48: op1_04_inv18 = 1;
    49: op1_04_inv18 = 1;
    53: op1_04_inv18 = 1;
    56: op1_04_inv18 = 1;
    57: op1_04_inv18 = 1;
    58: op1_04_inv18 = 1;
    60: op1_04_inv18 = 1;
    62: op1_04_inv18 = 1;
    63: op1_04_inv18 = 1;
    65: op1_04_inv18 = 1;
    70: op1_04_inv18 = 1;
    71: op1_04_inv18 = 1;
    72: op1_04_inv18 = 1;
    74: op1_04_inv18 = 1;
    77: op1_04_inv18 = 1;
    80: op1_04_inv18 = 1;
    81: op1_04_inv18 = 1;
    82: op1_04_inv18 = 1;
    86: op1_04_inv18 = 1;
    91: op1_04_inv18 = 1;
    96: op1_04_inv18 = 1;
    default: op1_04_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in19 = reg_0263;
    6: op1_04_in19 = reg_0212;
    15: op1_04_in19 = reg_0212;
    7: op1_04_in19 = reg_0044;
    8: op1_04_in19 = reg_0409;
    9: op1_04_in19 = reg_0136;
    10: op1_04_in19 = reg_0429;
    22: op1_04_in19 = reg_0429;
    11: op1_04_in19 = imem06_in[43:40];
    12: op1_04_in19 = reg_0124;
    13: op1_04_in19 = reg_0300;
    14: op1_04_in19 = reg_0383;
    16: op1_04_in19 = imem03_in[35:32];
    17: op1_04_in19 = reg_0436;
    18: op1_04_in19 = reg_0060;
    19: op1_04_in19 = reg_0406;
    20: op1_04_in19 = reg_0592;
    21: op1_04_in19 = reg_0632;
    23: op1_04_in19 = reg_0737;
    24: op1_04_in19 = reg_0207;
    25: op1_04_in19 = imem03_in[71:68];
    26: op1_04_in19 = reg_0246;
    27: op1_04_in19 = reg_0649;
    28: op1_04_in19 = imem07_in[71:68];
    30: op1_04_in19 = reg_0498;
    31: op1_04_in19 = reg_0735;
    81: op1_04_in19 = reg_0735;
    32: op1_04_in19 = reg_0717;
    33: op1_04_in19 = reg_0242;
    34: op1_04_in19 = reg_0381;
    35: op1_04_in19 = reg_0271;
    36: op1_04_in19 = imem06_in[75:72];
    37: op1_04_in19 = imem07_in[75:72];
    39: op1_04_in19 = reg_0508;
    41: op1_04_in19 = reg_0295;
    42: op1_04_in19 = reg_0371;
    44: op1_04_in19 = reg_0363;
    45: op1_04_in19 = reg_0280;
    46: op1_04_in19 = reg_0178;
    47: op1_04_in19 = reg_0188;
    48: op1_04_in19 = imem05_in[51:48];
    49: op1_04_in19 = reg_0392;
    50: op1_04_in19 = reg_0548;
    52: op1_04_in19 = reg_0112;
    53: op1_04_in19 = reg_0514;
    54: op1_04_in19 = reg_0391;
    55: op1_04_in19 = imem04_in[91:88];
    56: op1_04_in19 = reg_0486;
    57: op1_04_in19 = reg_0814;
    58: op1_04_in19 = reg_0430;
    60: op1_04_in19 = imem07_in[27:24];
    62: op1_04_in19 = reg_0594;
    63: op1_04_in19 = reg_0350;
    64: op1_04_in19 = reg_0223;
    65: op1_04_in19 = reg_0513;
    66: op1_04_in19 = imem04_in[55:52];
    67: op1_04_in19 = reg_0129;
    68: op1_04_in19 = reg_0192;
    69: op1_04_in19 = reg_0596;
    70: op1_04_in19 = reg_0153;
    71: op1_04_in19 = reg_0531;
    72: op1_04_in19 = imem04_in[19:16];
    73: op1_04_in19 = reg_0598;
    89: op1_04_in19 = reg_0598;
    74: op1_04_in19 = reg_0038;
    77: op1_04_in19 = imem01_in[115:112];
    78: op1_04_in19 = reg_0004;
    79: op1_04_in19 = reg_0771;
    80: op1_04_in19 = reg_0829;
    82: op1_04_in19 = imem01_in[63:60];
    83: op1_04_in19 = reg_0066;
    84: op1_04_in19 = imem04_in[119:116];
    85: op1_04_in19 = imem06_in[63:60];
    86: op1_04_in19 = reg_0530;
    87: op1_04_in19 = reg_0317;
    88: op1_04_in19 = reg_0709;
    90: op1_04_in19 = imem05_in[99:96];
    91: op1_04_in19 = reg_0788;
    96: op1_04_in19 = reg_0307;
    default: op1_04_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_04_inv19 = 1;
    9: op1_04_inv19 = 1;
    10: op1_04_inv19 = 1;
    12: op1_04_inv19 = 1;
    14: op1_04_inv19 = 1;
    15: op1_04_inv19 = 1;
    16: op1_04_inv19 = 1;
    19: op1_04_inv19 = 1;
    20: op1_04_inv19 = 1;
    21: op1_04_inv19 = 1;
    22: op1_04_inv19 = 1;
    24: op1_04_inv19 = 1;
    25: op1_04_inv19 = 1;
    34: op1_04_inv19 = 1;
    35: op1_04_inv19 = 1;
    36: op1_04_inv19 = 1;
    42: op1_04_inv19 = 1;
    45: op1_04_inv19 = 1;
    46: op1_04_inv19 = 1;
    48: op1_04_inv19 = 1;
    50: op1_04_inv19 = 1;
    57: op1_04_inv19 = 1;
    58: op1_04_inv19 = 1;
    62: op1_04_inv19 = 1;
    63: op1_04_inv19 = 1;
    66: op1_04_inv19 = 1;
    67: op1_04_inv19 = 1;
    69: op1_04_inv19 = 1;
    70: op1_04_inv19 = 1;
    72: op1_04_inv19 = 1;
    74: op1_04_inv19 = 1;
    79: op1_04_inv19 = 1;
    84: op1_04_inv19 = 1;
    86: op1_04_inv19 = 1;
    87: op1_04_inv19 = 1;
    88: op1_04_inv19 = 1;
    89: op1_04_inv19 = 1;
    90: op1_04_inv19 = 1;
    91: op1_04_inv19 = 1;
    96: op1_04_inv19 = 1;
    default: op1_04_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in20 = reg_0145;
    6: op1_04_in20 = reg_0197;
    68: op1_04_in20 = reg_0197;
    7: op1_04_in20 = imem05_in[3:0];
    8: op1_04_in20 = reg_0371;
    9: op1_04_in20 = reg_0128;
    10: op1_04_in20 = reg_0423;
    11: op1_04_in20 = imem06_in[47:44];
    12: op1_04_in20 = reg_0125;
    13: op1_04_in20 = reg_0295;
    14: op1_04_in20 = reg_0404;
    15: op1_04_in20 = reg_0202;
    16: op1_04_in20 = imem03_in[55:52];
    17: op1_04_in20 = reg_0419;
    18: op1_04_in20 = reg_0224;
    19: op1_04_in20 = reg_0039;
    20: op1_04_in20 = reg_0591;
    21: op1_04_in20 = reg_0386;
    22: op1_04_in20 = reg_0443;
    23: op1_04_in20 = reg_0276;
    24: op1_04_in20 = reg_0073;
    25: op1_04_in20 = imem03_in[87:84];
    26: op1_04_in20 = reg_0218;
    27: op1_04_in20 = reg_0229;
    28: op1_04_in20 = imem07_in[111:108];
    30: op1_04_in20 = reg_0028;
    31: op1_04_in20 = reg_0085;
    77: op1_04_in20 = reg_0085;
    32: op1_04_in20 = reg_0706;
    33: op1_04_in20 = reg_0502;
    34: op1_04_in20 = reg_0817;
    35: op1_04_in20 = reg_0275;
    36: op1_04_in20 = imem06_in[83:80];
    37: op1_04_in20 = imem07_in[95:92];
    39: op1_04_in20 = reg_0758;
    41: op1_04_in20 = reg_0051;
    42: op1_04_in20 = reg_0609;
    44: op1_04_in20 = reg_0324;
    45: op1_04_in20 = imem04_in[39:36];
    46: op1_04_in20 = reg_0173;
    47: op1_04_in20 = reg_0193;
    48: op1_04_in20 = imem05_in[95:92];
    49: op1_04_in20 = reg_0499;
    50: op1_04_in20 = reg_0426;
    52: op1_04_in20 = reg_0559;
    53: op1_04_in20 = reg_0092;
    54: op1_04_in20 = reg_0755;
    55: op1_04_in20 = imem04_in[107:104];
    56: op1_04_in20 = reg_0091;
    57: op1_04_in20 = reg_0298;
    58: op1_04_in20 = reg_0292;
    60: op1_04_in20 = imem07_in[55:52];
    62: op1_04_in20 = reg_0530;
    63: op1_04_in20 = reg_0488;
    69: op1_04_in20 = reg_0488;
    64: op1_04_in20 = reg_0062;
    65: op1_04_in20 = reg_0233;
    66: op1_04_in20 = imem04_in[59:56];
    67: op1_04_in20 = reg_0130;
    70: op1_04_in20 = reg_0141;
    71: op1_04_in20 = imem03_in[15:12];
    72: op1_04_in20 = imem04_in[67:64];
    73: op1_04_in20 = reg_0311;
    74: op1_04_in20 = reg_0401;
    78: op1_04_in20 = imem04_in[51:48];
    79: op1_04_in20 = reg_0640;
    80: op1_04_in20 = imem06_in[71:68];
    81: op1_04_in20 = reg_0278;
    82: op1_04_in20 = imem01_in[71:68];
    83: op1_04_in20 = reg_0184;
    84: op1_04_in20 = reg_0316;
    85: op1_04_in20 = imem06_in[111:108];
    86: op1_04_in20 = reg_0031;
    87: op1_04_in20 = reg_0596;
    88: op1_04_in20 = reg_0158;
    89: op1_04_in20 = imem05_in[55:52];
    90: op1_04_in20 = reg_0027;
    91: op1_04_in20 = reg_0231;
    96: op1_04_in20 = reg_0638;
    default: op1_04_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv20 = 1;
    12: op1_04_inv20 = 1;
    13: op1_04_inv20 = 1;
    14: op1_04_inv20 = 1;
    15: op1_04_inv20 = 1;
    16: op1_04_inv20 = 1;
    17: op1_04_inv20 = 1;
    19: op1_04_inv20 = 1;
    21: op1_04_inv20 = 1;
    24: op1_04_inv20 = 1;
    26: op1_04_inv20 = 1;
    31: op1_04_inv20 = 1;
    33: op1_04_inv20 = 1;
    35: op1_04_inv20 = 1;
    36: op1_04_inv20 = 1;
    41: op1_04_inv20 = 1;
    48: op1_04_inv20 = 1;
    52: op1_04_inv20 = 1;
    53: op1_04_inv20 = 1;
    54: op1_04_inv20 = 1;
    58: op1_04_inv20 = 1;
    60: op1_04_inv20 = 1;
    62: op1_04_inv20 = 1;
    64: op1_04_inv20 = 1;
    70: op1_04_inv20 = 1;
    72: op1_04_inv20 = 1;
    73: op1_04_inv20 = 1;
    74: op1_04_inv20 = 1;
    78: op1_04_inv20 = 1;
    79: op1_04_inv20 = 1;
    80: op1_04_inv20 = 1;
    81: op1_04_inv20 = 1;
    82: op1_04_inv20 = 1;
    88: op1_04_inv20 = 1;
    89: op1_04_inv20 = 1;
    90: op1_04_inv20 = 1;
    91: op1_04_inv20 = 1;
    default: op1_04_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in21 = reg_0140;
    70: op1_04_in21 = reg_0140;
    6: op1_04_in21 = imem01_in[107:104];
    7: op1_04_in21 = imem05_in[15:12];
    8: op1_04_in21 = reg_0382;
    9: op1_04_in21 = reg_0142;
    10: op1_04_in21 = reg_0439;
    11: op1_04_in21 = imem06_in[71:68];
    12: op1_04_in21 = reg_0102;
    82: op1_04_in21 = reg_0102;
    13: op1_04_in21 = reg_0065;
    14: op1_04_in21 = reg_0315;
    15: op1_04_in21 = imem01_in[11:8];
    16: op1_04_in21 = imem03_in[83:80];
    17: op1_04_in21 = reg_0431;
    18: op1_04_in21 = reg_0275;
    19: op1_04_in21 = reg_0752;
    20: op1_04_in21 = reg_0580;
    21: op1_04_in21 = reg_0399;
    63: op1_04_in21 = reg_0399;
    22: op1_04_in21 = reg_0175;
    23: op1_04_in21 = reg_0282;
    24: op1_04_in21 = reg_0229;
    25: op1_04_in21 = imem03_in[91:88];
    26: op1_04_in21 = reg_0242;
    74: op1_04_in21 = reg_0242;
    27: op1_04_in21 = reg_0356;
    28: op1_04_in21 = imem07_in[119:116];
    30: op1_04_in21 = reg_0371;
    31: op1_04_in21 = reg_0744;
    32: op1_04_in21 = reg_0700;
    33: op1_04_in21 = reg_0503;
    34: op1_04_in21 = reg_0819;
    35: op1_04_in21 = reg_0260;
    36: op1_04_in21 = imem06_in[95:92];
    37: op1_04_in21 = imem07_in[99:96];
    39: op1_04_in21 = reg_0501;
    41: op1_04_in21 = reg_0544;
    42: op1_04_in21 = reg_0317;
    44: op1_04_in21 = reg_0342;
    45: op1_04_in21 = imem04_in[91:88];
    47: op1_04_in21 = reg_0199;
    48: op1_04_in21 = imem05_in[99:96];
    49: op1_04_in21 = reg_0019;
    50: op1_04_in21 = reg_0359;
    52: op1_04_in21 = reg_0497;
    53: op1_04_in21 = reg_0530;
    54: op1_04_in21 = reg_0568;
    55: op1_04_in21 = imem04_in[119:116];
    56: op1_04_in21 = reg_0309;
    57: op1_04_in21 = reg_0618;
    58: op1_04_in21 = reg_0627;
    60: op1_04_in21 = imem07_in[75:72];
    62: op1_04_in21 = reg_0082;
    64: op1_04_in21 = reg_0585;
    65: op1_04_in21 = reg_0070;
    66: op1_04_in21 = imem04_in[107:104];
    67: op1_04_in21 = reg_0131;
    68: op1_04_in21 = reg_0646;
    69: op1_04_in21 = reg_0331;
    71: op1_04_in21 = imem03_in[43:40];
    72: op1_04_in21 = imem04_in[75:72];
    73: op1_04_in21 = reg_0771;
    77: op1_04_in21 = reg_0759;
    78: op1_04_in21 = imem04_in[59:56];
    79: op1_04_in21 = reg_0233;
    80: op1_04_in21 = imem06_in[75:72];
    81: op1_04_in21 = reg_0719;
    84: op1_04_in21 = reg_0060;
    85: op1_04_in21 = imem06_in[123:120];
    86: op1_04_in21 = reg_0753;
    87: op1_04_in21 = imem03_in[7:4];
    88: op1_04_in21 = reg_0711;
    89: op1_04_in21 = imem05_in[75:72];
    90: op1_04_in21 = reg_0665;
    91: op1_04_in21 = reg_0355;
    96: op1_04_in21 = reg_0328;
    default: op1_04_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv21 = 1;
    8: op1_04_inv21 = 1;
    9: op1_04_inv21 = 1;
    10: op1_04_inv21 = 1;
    12: op1_04_inv21 = 1;
    13: op1_04_inv21 = 1;
    14: op1_04_inv21 = 1;
    15: op1_04_inv21 = 1;
    16: op1_04_inv21 = 1;
    17: op1_04_inv21 = 1;
    18: op1_04_inv21 = 1;
    20: op1_04_inv21 = 1;
    23: op1_04_inv21 = 1;
    24: op1_04_inv21 = 1;
    25: op1_04_inv21 = 1;
    27: op1_04_inv21 = 1;
    30: op1_04_inv21 = 1;
    32: op1_04_inv21 = 1;
    34: op1_04_inv21 = 1;
    37: op1_04_inv21 = 1;
    39: op1_04_inv21 = 1;
    44: op1_04_inv21 = 1;
    45: op1_04_inv21 = 1;
    49: op1_04_inv21 = 1;
    53: op1_04_inv21 = 1;
    55: op1_04_inv21 = 1;
    56: op1_04_inv21 = 1;
    58: op1_04_inv21 = 1;
    60: op1_04_inv21 = 1;
    63: op1_04_inv21 = 1;
    64: op1_04_inv21 = 1;
    68: op1_04_inv21 = 1;
    71: op1_04_inv21 = 1;
    74: op1_04_inv21 = 1;
    77: op1_04_inv21 = 1;
    78: op1_04_inv21 = 1;
    80: op1_04_inv21 = 1;
    82: op1_04_inv21 = 1;
    84: op1_04_inv21 = 1;
    87: op1_04_inv21 = 1;
    88: op1_04_inv21 = 1;
    89: op1_04_inv21 = 1;
    91: op1_04_inv21 = 1;
    default: op1_04_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in22 = imem06_in[47:44];
    6: op1_04_in22 = imem01_in[111:108];
    7: op1_04_in22 = imem05_in[75:72];
    8: op1_04_in22 = reg_0380;
    9: op1_04_in22 = reg_0146;
    10: op1_04_in22 = reg_0435;
    11: op1_04_in22 = imem06_in[79:76];
    12: op1_04_in22 = reg_0114;
    13: op1_04_in22 = reg_0056;
    14: op1_04_in22 = reg_0390;
    15: op1_04_in22 = imem01_in[23:20];
    16: op1_04_in22 = reg_0582;
    17: op1_04_in22 = reg_0172;
    18: op1_04_in22 = reg_0543;
    19: op1_04_in22 = imem07_in[11:8];
    20: op1_04_in22 = reg_0595;
    21: op1_04_in22 = reg_0753;
    22: op1_04_in22 = reg_0167;
    23: op1_04_in22 = reg_0260;
    24: op1_04_in22 = reg_0320;
    25: op1_04_in22 = imem03_in[95:92];
    26: op1_04_in22 = reg_0216;
    27: op1_04_in22 = reg_0363;
    28: op1_04_in22 = reg_0719;
    30: op1_04_in22 = reg_0338;
    31: op1_04_in22 = reg_0734;
    32: op1_04_in22 = reg_0432;
    33: op1_04_in22 = reg_0236;
    34: op1_04_in22 = reg_0605;
    35: op1_04_in22 = reg_0744;
    36: op1_04_in22 = imem06_in[99:96];
    37: op1_04_in22 = reg_0728;
    39: op1_04_in22 = reg_0497;
    41: op1_04_in22 = reg_0315;
    42: op1_04_in22 = reg_0408;
    44: op1_04_in22 = reg_0518;
    45: op1_04_in22 = imem04_in[103:100];
    47: op1_04_in22 = reg_0062;
    48: op1_04_in22 = reg_0781;
    49: op1_04_in22 = reg_0804;
    50: op1_04_in22 = reg_0361;
    52: op1_04_in22 = reg_0225;
    53: op1_04_in22 = reg_0063;
    54: op1_04_in22 = reg_0383;
    55: op1_04_in22 = imem04_in[127:124];
    56: op1_04_in22 = reg_0256;
    57: op1_04_in22 = reg_0339;
    58: op1_04_in22 = imem04_in[87:84];
    60: op1_04_in22 = imem07_in[91:88];
    62: op1_04_in22 = reg_0538;
    63: op1_04_in22 = reg_0281;
    64: op1_04_in22 = reg_0371;
    65: op1_04_in22 = reg_0102;
    66: op1_04_in22 = reg_0328;
    67: op1_04_in22 = imem06_in[55:52];
    68: op1_04_in22 = reg_0037;
    69: op1_04_in22 = imem03_in[23:20];
    70: op1_04_in22 = reg_0137;
    71: op1_04_in22 = imem03_in[107:104];
    72: op1_04_in22 = imem04_in[79:76];
    73: op1_04_in22 = reg_0233;
    74: op1_04_in22 = reg_0369;
    77: op1_04_in22 = reg_0778;
    78: op1_04_in22 = imem04_in[63:60];
    79: op1_04_in22 = reg_0109;
    80: op1_04_in22 = imem06_in[83:80];
    81: op1_04_in22 = reg_0277;
    82: op1_04_in22 = reg_0394;
    84: op1_04_in22 = reg_0554;
    85: op1_04_in22 = imem06_in[127:124];
    86: op1_04_in22 = reg_0075;
    87: op1_04_in22 = imem03_in[19:16];
    88: op1_04_in22 = reg_0724;
    89: op1_04_in22 = imem05_in[83:80];
    90: op1_04_in22 = reg_0517;
    91: op1_04_in22 = reg_0134;
    96: op1_04_in22 = reg_0655;
    default: op1_04_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_04_inv22 = 1;
    12: op1_04_inv22 = 1;
    13: op1_04_inv22 = 1;
    15: op1_04_inv22 = 1;
    18: op1_04_inv22 = 1;
    20: op1_04_inv22 = 1;
    21: op1_04_inv22 = 1;
    24: op1_04_inv22 = 1;
    28: op1_04_inv22 = 1;
    33: op1_04_inv22 = 1;
    34: op1_04_inv22 = 1;
    35: op1_04_inv22 = 1;
    36: op1_04_inv22 = 1;
    39: op1_04_inv22 = 1;
    45: op1_04_inv22 = 1;
    47: op1_04_inv22 = 1;
    49: op1_04_inv22 = 1;
    50: op1_04_inv22 = 1;
    52: op1_04_inv22 = 1;
    54: op1_04_inv22 = 1;
    55: op1_04_inv22 = 1;
    57: op1_04_inv22 = 1;
    58: op1_04_inv22 = 1;
    60: op1_04_inv22 = 1;
    62: op1_04_inv22 = 1;
    66: op1_04_inv22 = 1;
    67: op1_04_inv22 = 1;
    68: op1_04_inv22 = 1;
    69: op1_04_inv22 = 1;
    72: op1_04_inv22 = 1;
    77: op1_04_inv22 = 1;
    80: op1_04_inv22 = 1;
    81: op1_04_inv22 = 1;
    82: op1_04_inv22 = 1;
    84: op1_04_inv22 = 1;
    86: op1_04_inv22 = 1;
    88: op1_04_inv22 = 1;
    89: op1_04_inv22 = 1;
    96: op1_04_inv22 = 1;
    default: op1_04_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in23 = imem06_in[67:64];
    6: op1_04_in23 = reg_0499;
    7: op1_04_in23 = imem05_in[83:80];
    8: op1_04_in23 = imem06_in[71:68];
    9: op1_04_in23 = reg_0139;
    10: op1_04_in23 = reg_0175;
    11: op1_04_in23 = imem06_in[83:80];
    12: op1_04_in23 = reg_0107;
    13: op1_04_in23 = reg_0064;
    14: op1_04_in23 = reg_0028;
    15: op1_04_in23 = imem01_in[83:80];
    16: op1_04_in23 = reg_0573;
    18: op1_04_in23 = reg_0536;
    19: op1_04_in23 = imem07_in[31:28];
    20: op1_04_in23 = reg_0576;
    21: op1_04_in23 = imem07_in[55:52];
    22: op1_04_in23 = reg_0160;
    23: op1_04_in23 = reg_0277;
    24: op1_04_in23 = reg_0321;
    25: op1_04_in23 = reg_0583;
    53: op1_04_in23 = reg_0583;
    26: op1_04_in23 = reg_0220;
    27: op1_04_in23 = reg_0343;
    28: op1_04_in23 = reg_0731;
    30: op1_04_in23 = reg_0368;
    31: op1_04_in23 = reg_0285;
    32: op1_04_in23 = reg_0439;
    33: op1_04_in23 = reg_0248;
    34: op1_04_in23 = reg_0380;
    35: op1_04_in23 = reg_0734;
    36: op1_04_in23 = imem06_in[103:100];
    37: op1_04_in23 = reg_0719;
    39: op1_04_in23 = reg_0512;
    41: op1_04_in23 = reg_0328;
    42: op1_04_in23 = reg_0763;
    74: op1_04_in23 = reg_0763;
    44: op1_04_in23 = reg_0081;
    45: op1_04_in23 = imem05_in[7:4];
    79: op1_04_in23 = imem05_in[7:4];
    47: op1_04_in23 = reg_0246;
    48: op1_04_in23 = reg_0795;
    49: op1_04_in23 = reg_0801;
    50: op1_04_in23 = reg_0356;
    52: op1_04_in23 = reg_0574;
    54: op1_04_in23 = reg_0747;
    55: op1_04_in23 = reg_0262;
    56: op1_04_in23 = reg_0070;
    57: op1_04_in23 = imem06_in[59:56];
    58: op1_04_in23 = imem04_in[95:92];
    72: op1_04_in23 = imem04_in[95:92];
    60: op1_04_in23 = imem07_in[127:124];
    62: op1_04_in23 = reg_0094;
    63: op1_04_in23 = reg_0394;
    64: op1_04_in23 = reg_0233;
    65: op1_04_in23 = reg_0227;
    66: op1_04_in23 = reg_0055;
    67: op1_04_in23 = imem06_in[99:96];
    80: op1_04_in23 = imem06_in[99:96];
    68: op1_04_in23 = reg_0825;
    69: op1_04_in23 = imem03_in[31:28];
    70: op1_04_in23 = reg_0534;
    71: op1_04_in23 = reg_0317;
    73: op1_04_in23 = reg_0416;
    77: op1_04_in23 = reg_0110;
    78: op1_04_in23 = imem04_in[67:64];
    81: op1_04_in23 = reg_0389;
    82: op1_04_in23 = reg_0397;
    84: op1_04_in23 = reg_0629;
    85: op1_04_in23 = reg_0563;
    86: op1_04_in23 = reg_0256;
    87: op1_04_in23 = imem03_in[35:32];
    88: op1_04_in23 = reg_0253;
    89: op1_04_in23 = imem05_in[87:84];
    90: op1_04_in23 = reg_0386;
    91: op1_04_in23 = reg_0226;
    96: op1_04_in23 = reg_0681;
    default: op1_04_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv23 = 1;
    7: op1_04_inv23 = 1;
    8: op1_04_inv23 = 1;
    9: op1_04_inv23 = 1;
    11: op1_04_inv23 = 1;
    12: op1_04_inv23 = 1;
    13: op1_04_inv23 = 1;
    21: op1_04_inv23 = 1;
    24: op1_04_inv23 = 1;
    25: op1_04_inv23 = 1;
    26: op1_04_inv23 = 1;
    27: op1_04_inv23 = 1;
    30: op1_04_inv23 = 1;
    33: op1_04_inv23 = 1;
    35: op1_04_inv23 = 1;
    39: op1_04_inv23 = 1;
    41: op1_04_inv23 = 1;
    47: op1_04_inv23 = 1;
    49: op1_04_inv23 = 1;
    53: op1_04_inv23 = 1;
    56: op1_04_inv23 = 1;
    57: op1_04_inv23 = 1;
    58: op1_04_inv23 = 1;
    64: op1_04_inv23 = 1;
    68: op1_04_inv23 = 1;
    70: op1_04_inv23 = 1;
    77: op1_04_inv23 = 1;
    79: op1_04_inv23 = 1;
    82: op1_04_inv23 = 1;
    84: op1_04_inv23 = 1;
    85: op1_04_inv23 = 1;
    86: op1_04_inv23 = 1;
    88: op1_04_inv23 = 1;
    89: op1_04_inv23 = 1;
    90: op1_04_inv23 = 1;
    91: op1_04_inv23 = 1;
    default: op1_04_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in24 = imem06_in[95:92];
    6: op1_04_in24 = reg_0518;
    90: op1_04_in24 = reg_0518;
    7: op1_04_in24 = imem05_in[107:104];
    8: op1_04_in24 = imem06_in[99:96];
    11: op1_04_in24 = imem06_in[99:96];
    9: op1_04_in24 = reg_0137;
    10: op1_04_in24 = reg_0161;
    12: op1_04_in24 = reg_0127;
    13: op1_04_in24 = imem05_in[15:12];
    45: op1_04_in24 = imem05_in[15:12];
    79: op1_04_in24 = imem05_in[15:12];
    14: op1_04_in24 = reg_0039;
    65: op1_04_in24 = reg_0039;
    15: op1_04_in24 = imem01_in[103:100];
    16: op1_04_in24 = reg_0583;
    18: op1_04_in24 = reg_0548;
    19: op1_04_in24 = imem07_in[63:60];
    20: op1_04_in24 = reg_0321;
    21: op1_04_in24 = reg_0722;
    22: op1_04_in24 = reg_0183;
    23: op1_04_in24 = reg_0128;
    24: op1_04_in24 = imem01_in[15:12];
    25: op1_04_in24 = reg_0592;
    26: op1_04_in24 = reg_0237;
    47: op1_04_in24 = reg_0237;
    27: op1_04_in24 = reg_0323;
    28: op1_04_in24 = reg_0724;
    30: op1_04_in24 = reg_0372;
    31: op1_04_in24 = reg_0135;
    32: op1_04_in24 = reg_0427;
    33: op1_04_in24 = reg_0238;
    34: op1_04_in24 = imem07_in[19:16];
    35: op1_04_in24 = reg_0086;
    36: op1_04_in24 = imem07_in[27:24];
    37: op1_04_in24 = reg_0710;
    39: op1_04_in24 = reg_0333;
    41: op1_04_in24 = reg_0555;
    42: op1_04_in24 = reg_0270;
    74: op1_04_in24 = reg_0270;
    44: op1_04_in24 = reg_0539;
    48: op1_04_in24 = reg_0780;
    49: op1_04_in24 = reg_0799;
    50: op1_04_in24 = reg_0360;
    52: op1_04_in24 = reg_0505;
    53: op1_04_in24 = reg_0347;
    54: op1_04_in24 = reg_0374;
    55: op1_04_in24 = reg_0553;
    56: op1_04_in24 = reg_0229;
    57: op1_04_in24 = imem06_in[67:64];
    58: op1_04_in24 = imem05_in[39:36];
    60: op1_04_in24 = reg_0731;
    62: op1_04_in24 = reg_0532;
    63: op1_04_in24 = reg_0395;
    64: op1_04_in24 = reg_0288;
    66: op1_04_in24 = reg_0554;
    67: op1_04_in24 = imem06_in[107:104];
    68: op1_04_in24 = reg_0304;
    69: op1_04_in24 = imem03_in[43:40];
    70: op1_04_in24 = reg_0037;
    71: op1_04_in24 = reg_0116;
    72: op1_04_in24 = reg_0059;
    86: op1_04_in24 = reg_0059;
    73: op1_04_in24 = reg_0252;
    77: op1_04_in24 = reg_0423;
    78: op1_04_in24 = imem04_in[87:84];
    80: op1_04_in24 = imem06_in[127:124];
    81: op1_04_in24 = reg_0285;
    82: op1_04_in24 = reg_0241;
    84: op1_04_in24 = reg_0292;
    85: op1_04_in24 = reg_0218;
    96: op1_04_in24 = reg_0218;
    87: op1_04_in24 = imem03_in[75:72];
    88: op1_04_in24 = reg_0636;
    89: op1_04_in24 = imem05_in[91:88];
    91: op1_04_in24 = reg_0538;
    default: op1_04_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv24 = 1;
    9: op1_04_inv24 = 1;
    10: op1_04_inv24 = 1;
    11: op1_04_inv24 = 1;
    13: op1_04_inv24 = 1;
    14: op1_04_inv24 = 1;
    21: op1_04_inv24 = 1;
    23: op1_04_inv24 = 1;
    24: op1_04_inv24 = 1;
    25: op1_04_inv24 = 1;
    26: op1_04_inv24 = 1;
    27: op1_04_inv24 = 1;
    28: op1_04_inv24 = 1;
    36: op1_04_inv24 = 1;
    37: op1_04_inv24 = 1;
    41: op1_04_inv24 = 1;
    42: op1_04_inv24 = 1;
    44: op1_04_inv24 = 1;
    48: op1_04_inv24 = 1;
    49: op1_04_inv24 = 1;
    53: op1_04_inv24 = 1;
    54: op1_04_inv24 = 1;
    63: op1_04_inv24 = 1;
    64: op1_04_inv24 = 1;
    66: op1_04_inv24 = 1;
    68: op1_04_inv24 = 1;
    69: op1_04_inv24 = 1;
    70: op1_04_inv24 = 1;
    71: op1_04_inv24 = 1;
    78: op1_04_inv24 = 1;
    79: op1_04_inv24 = 1;
    84: op1_04_inv24 = 1;
    85: op1_04_inv24 = 1;
    86: op1_04_inv24 = 1;
    87: op1_04_inv24 = 1;
    89: op1_04_inv24 = 1;
    91: op1_04_inv24 = 1;
    96: op1_04_inv24 = 1;
    default: op1_04_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in25 = reg_0628;
    6: op1_04_in25 = reg_0515;
    39: op1_04_in25 = reg_0515;
    7: op1_04_in25 = imem05_in[115:112];
    8: op1_04_in25 = imem06_in[115:112];
    9: op1_04_in25 = imem06_in[15:12];
    10: op1_04_in25 = reg_0163;
    11: op1_04_in25 = imem06_in[119:116];
    12: op1_04_in25 = imem02_in[3:0];
    13: op1_04_in25 = imem05_in[39:36];
    14: op1_04_in25 = reg_0035;
    15: op1_04_in25 = imem01_in[107:104];
    16: op1_04_in25 = reg_0592;
    18: op1_04_in25 = reg_0555;
    19: op1_04_in25 = imem07_in[107:104];
    20: op1_04_in25 = reg_0397;
    21: op1_04_in25 = reg_0716;
    22: op1_04_in25 = reg_0177;
    23: op1_04_in25 = reg_0152;
    24: op1_04_in25 = imem01_in[39:36];
    25: op1_04_in25 = reg_0585;
    26: op1_04_in25 = reg_0234;
    27: op1_04_in25 = reg_0541;
    28: op1_04_in25 = reg_0715;
    30: op1_04_in25 = imem03_in[7:4];
    44: op1_04_in25 = imem03_in[7:4];
    31: op1_04_in25 = reg_0143;
    32: op1_04_in25 = reg_0448;
    33: op1_04_in25 = reg_0122;
    34: op1_04_in25 = imem07_in[59:56];
    35: op1_04_in25 = reg_0145;
    79: op1_04_in25 = reg_0145;
    36: op1_04_in25 = imem07_in[31:28];
    37: op1_04_in25 = reg_0729;
    41: op1_04_in25 = reg_0060;
    42: op1_04_in25 = reg_0403;
    45: op1_04_in25 = imem05_in[19:16];
    47: op1_04_in25 = imem01_in[47:44];
    48: op1_04_in25 = reg_0790;
    49: op1_04_in25 = reg_0010;
    50: op1_04_in25 = reg_0092;
    52: op1_04_in25 = imem01_in[15:12];
    53: op1_04_in25 = imem03_in[3:0];
    62: op1_04_in25 = imem03_in[3:0];
    54: op1_04_in25 = reg_0008;
    55: op1_04_in25 = reg_0554;
    56: op1_04_in25 = reg_0249;
    57: op1_04_in25 = imem06_in[75:72];
    58: op1_04_in25 = imem05_in[43:40];
    60: op1_04_in25 = reg_0705;
    63: op1_04_in25 = reg_0391;
    64: op1_04_in25 = reg_0040;
    65: op1_04_in25 = reg_0258;
    66: op1_04_in25 = reg_0523;
    67: op1_04_in25 = imem06_in[111:108];
    68: op1_04_in25 = reg_0321;
    69: op1_04_in25 = imem03_in[59:56];
    70: op1_04_in25 = reg_0100;
    71: op1_04_in25 = reg_0350;
    72: op1_04_in25 = reg_0262;
    73: op1_04_in25 = reg_0132;
    74: op1_04_in25 = reg_0608;
    77: op1_04_in25 = reg_0418;
    78: op1_04_in25 = imem04_in[119:116];
    80: op1_04_in25 = reg_0299;
    81: op1_04_in25 = reg_0148;
    82: op1_04_in25 = reg_0306;
    84: op1_04_in25 = reg_0627;
    85: op1_04_in25 = imem07_in[23:20];
    86: op1_04_in25 = reg_0320;
    87: op1_04_in25 = reg_0028;
    88: op1_04_in25 = reg_0442;
    89: op1_04_in25 = imem05_in[95:92];
    90: op1_04_in25 = reg_0538;
    91: op1_04_in25 = reg_0488;
    96: op1_04_in25 = reg_0621;
    default: op1_04_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv25 = 1;
    6: op1_04_inv25 = 1;
    7: op1_04_inv25 = 1;
    9: op1_04_inv25 = 1;
    11: op1_04_inv25 = 1;
    13: op1_04_inv25 = 1;
    18: op1_04_inv25 = 1;
    19: op1_04_inv25 = 1;
    20: op1_04_inv25 = 1;
    21: op1_04_inv25 = 1;
    22: op1_04_inv25 = 1;
    23: op1_04_inv25 = 1;
    25: op1_04_inv25 = 1;
    26: op1_04_inv25 = 1;
    27: op1_04_inv25 = 1;
    28: op1_04_inv25 = 1;
    33: op1_04_inv25 = 1;
    34: op1_04_inv25 = 1;
    35: op1_04_inv25 = 1;
    36: op1_04_inv25 = 1;
    37: op1_04_inv25 = 1;
    39: op1_04_inv25 = 1;
    41: op1_04_inv25 = 1;
    42: op1_04_inv25 = 1;
    47: op1_04_inv25 = 1;
    50: op1_04_inv25 = 1;
    52: op1_04_inv25 = 1;
    53: op1_04_inv25 = 1;
    54: op1_04_inv25 = 1;
    55: op1_04_inv25 = 1;
    56: op1_04_inv25 = 1;
    58: op1_04_inv25 = 1;
    60: op1_04_inv25 = 1;
    62: op1_04_inv25 = 1;
    64: op1_04_inv25 = 1;
    68: op1_04_inv25 = 1;
    70: op1_04_inv25 = 1;
    71: op1_04_inv25 = 1;
    72: op1_04_inv25 = 1;
    73: op1_04_inv25 = 1;
    74: op1_04_inv25 = 1;
    81: op1_04_inv25 = 1;
    86: op1_04_inv25 = 1;
    88: op1_04_inv25 = 1;
    91: op1_04_inv25 = 1;
    96: op1_04_inv25 = 1;
    default: op1_04_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in26 = reg_0613;
    6: op1_04_in26 = reg_0233;
    7: op1_04_in26 = reg_0488;
    90: op1_04_in26 = reg_0488;
    8: op1_04_in26 = imem07_in[39:36];
    85: op1_04_in26 = imem07_in[39:36];
    9: op1_04_in26 = imem06_in[39:36];
    10: op1_04_in26 = reg_0183;
    11: op1_04_in26 = reg_0628;
    12: op1_04_in26 = reg_0645;
    13: op1_04_in26 = imem05_in[43:40];
    14: op1_04_in26 = reg_0040;
    15: op1_04_in26 = reg_0227;
    79: op1_04_in26 = reg_0227;
    16: op1_04_in26 = reg_0578;
    18: op1_04_in26 = reg_0549;
    19: op1_04_in26 = reg_0721;
    20: op1_04_in26 = reg_0389;
    21: op1_04_in26 = reg_0712;
    22: op1_04_in26 = reg_0168;
    23: op1_04_in26 = reg_0146;
    24: op1_04_in26 = imem01_in[51:48];
    25: op1_04_in26 = reg_0593;
    26: op1_04_in26 = reg_0219;
    27: op1_04_in26 = reg_0533;
    28: op1_04_in26 = reg_0701;
    30: op1_04_in26 = imem03_in[15:12];
    31: op1_04_in26 = reg_0139;
    32: op1_04_in26 = reg_0435;
    33: op1_04_in26 = reg_0116;
    34: op1_04_in26 = imem07_in[103:100];
    35: op1_04_in26 = reg_0133;
    36: op1_04_in26 = imem07_in[47:44];
    37: op1_04_in26 = reg_0705;
    39: op1_04_in26 = reg_0557;
    41: op1_04_in26 = reg_0556;
    42: op1_04_in26 = reg_0614;
    44: op1_04_in26 = imem03_in[43:40];
    45: op1_04_in26 = imem05_in[27:24];
    47: op1_04_in26 = imem01_in[59:56];
    48: op1_04_in26 = reg_0489;
    49: op1_04_in26 = imem04_in[27:24];
    50: op1_04_in26 = reg_0530;
    52: op1_04_in26 = imem01_in[27:24];
    68: op1_04_in26 = imem01_in[27:24];
    53: op1_04_in26 = imem03_in[19:16];
    54: op1_04_in26 = reg_0015;
    55: op1_04_in26 = reg_0523;
    56: op1_04_in26 = reg_0066;
    57: op1_04_in26 = reg_0777;
    58: op1_04_in26 = imem05_in[47:44];
    60: op1_04_in26 = reg_0707;
    62: op1_04_in26 = imem03_in[7:4];
    63: op1_04_in26 = reg_0383;
    64: op1_04_in26 = reg_0269;
    65: op1_04_in26 = reg_0101;
    66: op1_04_in26 = reg_0547;
    67: op1_04_in26 = imem06_in[119:116];
    69: op1_04_in26 = imem03_in[63:60];
    70: op1_04_in26 = reg_0072;
    71: op1_04_in26 = reg_0329;
    72: op1_04_in26 = reg_0558;
    73: op1_04_in26 = reg_0277;
    74: op1_04_in26 = reg_0583;
    77: op1_04_in26 = reg_0240;
    78: op1_04_in26 = imem04_in[123:120];
    80: op1_04_in26 = reg_0265;
    81: op1_04_in26 = reg_0150;
    82: op1_04_in26 = reg_0567;
    84: op1_04_in26 = reg_0626;
    86: op1_04_in26 = reg_0341;
    87: op1_04_in26 = reg_0483;
    88: op1_04_in26 = reg_0437;
    89: op1_04_in26 = imem05_in[103:100];
    91: op1_04_in26 = reg_0229;
    96: op1_04_in26 = reg_0657;
    default: op1_04_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv26 = 1;
    8: op1_04_inv26 = 1;
    9: op1_04_inv26 = 1;
    10: op1_04_inv26 = 1;
    11: op1_04_inv26 = 1;
    12: op1_04_inv26 = 1;
    16: op1_04_inv26 = 1;
    18: op1_04_inv26 = 1;
    20: op1_04_inv26 = 1;
    23: op1_04_inv26 = 1;
    24: op1_04_inv26 = 1;
    25: op1_04_inv26 = 1;
    26: op1_04_inv26 = 1;
    28: op1_04_inv26 = 1;
    31: op1_04_inv26 = 1;
    32: op1_04_inv26 = 1;
    33: op1_04_inv26 = 1;
    35: op1_04_inv26 = 1;
    37: op1_04_inv26 = 1;
    45: op1_04_inv26 = 1;
    48: op1_04_inv26 = 1;
    50: op1_04_inv26 = 1;
    52: op1_04_inv26 = 1;
    54: op1_04_inv26 = 1;
    55: op1_04_inv26 = 1;
    58: op1_04_inv26 = 1;
    63: op1_04_inv26 = 1;
    65: op1_04_inv26 = 1;
    67: op1_04_inv26 = 1;
    70: op1_04_inv26 = 1;
    71: op1_04_inv26 = 1;
    73: op1_04_inv26 = 1;
    74: op1_04_inv26 = 1;
    79: op1_04_inv26 = 1;
    82: op1_04_inv26 = 1;
    84: op1_04_inv26 = 1;
    85: op1_04_inv26 = 1;
    86: op1_04_inv26 = 1;
    89: op1_04_inv26 = 1;
    91: op1_04_inv26 = 1;
    default: op1_04_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in27 = reg_0612;
    6: op1_04_in27 = reg_0246;
    7: op1_04_in27 = reg_0789;
    8: op1_04_in27 = imem07_in[47:44];
    85: op1_04_in27 = imem07_in[47:44];
    9: op1_04_in27 = imem06_in[67:64];
    11: op1_04_in27 = reg_0351;
    12: op1_04_in27 = reg_0666;
    13: op1_04_in27 = imem05_in[67:64];
    14: op1_04_in27 = reg_0036;
    15: op1_04_in27 = reg_0521;
    16: op1_04_in27 = reg_0360;
    18: op1_04_in27 = reg_0546;
    19: op1_04_in27 = reg_0729;
    20: op1_04_in27 = reg_0000;
    21: op1_04_in27 = reg_0709;
    22: op1_04_in27 = reg_0173;
    23: op1_04_in27 = reg_0138;
    24: op1_04_in27 = imem01_in[79:76];
    25: op1_04_in27 = reg_0597;
    26: op1_04_in27 = reg_0108;
    27: op1_04_in27 = reg_0081;
    28: op1_04_in27 = reg_0429;
    30: op1_04_in27 = imem03_in[35:32];
    31: op1_04_in27 = reg_0153;
    32: op1_04_in27 = reg_0180;
    33: op1_04_in27 = imem02_in[3:0];
    34: op1_04_in27 = reg_0728;
    35: op1_04_in27 = reg_0142;
    36: op1_04_in27 = reg_0717;
    37: op1_04_in27 = reg_0707;
    39: op1_04_in27 = reg_0507;
    41: op1_04_in27 = imem04_in[39:36];
    42: op1_04_in27 = reg_0040;
    44: op1_04_in27 = imem03_in[55:52];
    45: op1_04_in27 = imem05_in[87:84];
    47: op1_04_in27 = imem01_in[75:72];
    48: op1_04_in27 = reg_0282;
    49: op1_04_in27 = imem04_in[35:32];
    50: op1_04_in27 = reg_0540;
    52: op1_04_in27 = imem01_in[35:32];
    53: op1_04_in27 = imem03_in[39:36];
    54: op1_04_in27 = reg_0016;
    55: op1_04_in27 = reg_0510;
    56: op1_04_in27 = reg_0285;
    57: op1_04_in27 = reg_0620;
    58: op1_04_in27 = imem05_in[107:104];
    60: op1_04_in27 = reg_0706;
    62: op1_04_in27 = imem03_in[15:12];
    63: op1_04_in27 = reg_0385;
    64: op1_04_in27 = reg_0066;
    65: op1_04_in27 = reg_0277;
    66: op1_04_in27 = reg_0432;
    67: op1_04_in27 = imem06_in[123:120];
    68: op1_04_in27 = imem01_in[71:68];
    69: op1_04_in27 = imem03_in[83:80];
    70: op1_04_in27 = reg_0625;
    71: op1_04_in27 = reg_0357;
    72: op1_04_in27 = reg_0551;
    73: op1_04_in27 = reg_0135;
    74: op1_04_in27 = reg_0035;
    77: op1_04_in27 = reg_0244;
    78: op1_04_in27 = imem04_in[127:124];
    79: op1_04_in27 = reg_0070;
    80: op1_04_in27 = reg_0628;
    81: op1_04_in27 = reg_0829;
    82: op1_04_in27 = reg_0123;
    84: op1_04_in27 = reg_0078;
    86: op1_04_in27 = reg_0565;
    87: op1_04_in27 = reg_0569;
    88: op1_04_in27 = reg_0448;
    89: op1_04_in27 = imem05_in[111:108];
    90: op1_04_in27 = reg_0229;
    91: op1_04_in27 = reg_0751;
    96: op1_04_in27 = reg_0501;
    default: op1_04_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv27 = 1;
    7: op1_04_inv27 = 1;
    8: op1_04_inv27 = 1;
    12: op1_04_inv27 = 1;
    14: op1_04_inv27 = 1;
    15: op1_04_inv27 = 1;
    20: op1_04_inv27 = 1;
    22: op1_04_inv27 = 1;
    26: op1_04_inv27 = 1;
    30: op1_04_inv27 = 1;
    34: op1_04_inv27 = 1;
    36: op1_04_inv27 = 1;
    44: op1_04_inv27 = 1;
    49: op1_04_inv27 = 1;
    50: op1_04_inv27 = 1;
    52: op1_04_inv27 = 1;
    53: op1_04_inv27 = 1;
    55: op1_04_inv27 = 1;
    56: op1_04_inv27 = 1;
    57: op1_04_inv27 = 1;
    58: op1_04_inv27 = 1;
    60: op1_04_inv27 = 1;
    64: op1_04_inv27 = 1;
    65: op1_04_inv27 = 1;
    66: op1_04_inv27 = 1;
    69: op1_04_inv27 = 1;
    70: op1_04_inv27 = 1;
    73: op1_04_inv27 = 1;
    74: op1_04_inv27 = 1;
    77: op1_04_inv27 = 1;
    85: op1_04_inv27 = 1;
    86: op1_04_inv27 = 1;
    87: op1_04_inv27 = 1;
    88: op1_04_inv27 = 1;
    89: op1_04_inv27 = 1;
    90: op1_04_inv27 = 1;
    96: op1_04_inv27 = 1;
    default: op1_04_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in28 = reg_0348;
    6: op1_04_in28 = reg_0245;
    7: op1_04_in28 = reg_0793;
    8: op1_04_in28 = imem07_in[83:80];
    9: op1_04_in28 = imem06_in[71:68];
    11: op1_04_in28 = reg_0748;
    12: op1_04_in28 = reg_0639;
    13: op1_04_in28 = imem05_in[79:76];
    14: op1_04_in28 = reg_0037;
    96: op1_04_in28 = reg_0037;
    15: op1_04_in28 = reg_0499;
    16: op1_04_in28 = reg_0370;
    18: op1_04_in28 = reg_0540;
    27: op1_04_in28 = reg_0540;
    19: op1_04_in28 = reg_0709;
    20: op1_04_in28 = reg_0019;
    21: op1_04_in28 = reg_0718;
    22: op1_04_in28 = reg_0171;
    23: op1_04_in28 = reg_0144;
    24: op1_04_in28 = imem01_in[103:100];
    25: op1_04_in28 = reg_0570;
    26: op1_04_in28 = reg_0114;
    28: op1_04_in28 = reg_0174;
    30: op1_04_in28 = imem03_in[43:40];
    53: op1_04_in28 = imem03_in[43:40];
    31: op1_04_in28 = reg_0029;
    74: op1_04_in28 = reg_0029;
    32: op1_04_in28 = reg_0165;
    33: op1_04_in28 = imem02_in[11:8];
    34: op1_04_in28 = reg_0720;
    35: op1_04_in28 = reg_0138;
    36: op1_04_in28 = reg_0729;
    37: op1_04_in28 = reg_0428;
    39: op1_04_in28 = imem01_in[47:44];
    41: op1_04_in28 = imem04_in[55:52];
    42: op1_04_in28 = reg_0375;
    44: op1_04_in28 = imem03_in[111:108];
    45: op1_04_in28 = imem05_in[99:96];
    47: op1_04_in28 = imem01_in[83:80];
    48: op1_04_in28 = reg_0277;
    49: op1_04_in28 = imem04_in[39:36];
    50: op1_04_in28 = imem03_in[15:12];
    52: op1_04_in28 = imem01_in[67:64];
    54: op1_04_in28 = imem04_in[7:4];
    55: op1_04_in28 = reg_0429;
    56: op1_04_in28 = reg_0148;
    57: op1_04_in28 = reg_0040;
    58: op1_04_in28 = imem05_in[123:120];
    89: op1_04_in28 = imem05_in[123:120];
    60: op1_04_in28 = reg_0727;
    62: op1_04_in28 = imem03_in[27:24];
    63: op1_04_in28 = reg_0002;
    69: op1_04_in28 = reg_0002;
    64: op1_04_in28 = imem05_in[7:4];
    65: op1_04_in28 = reg_0784;
    66: op1_04_in28 = reg_0615;
    67: op1_04_in28 = reg_0618;
    68: op1_04_in28 = imem01_in[107:104];
    70: op1_04_in28 = reg_0349;
    71: op1_04_in28 = reg_0751;
    72: op1_04_in28 = reg_0433;
    73: op1_04_in28 = reg_0113;
    77: op1_04_in28 = reg_0425;
    78: op1_04_in28 = reg_0059;
    79: op1_04_in28 = reg_0231;
    80: op1_04_in28 = reg_0578;
    81: op1_04_in28 = reg_0257;
    82: op1_04_in28 = reg_0124;
    84: op1_04_in28 = reg_0062;
    85: op1_04_in28 = imem07_in[55:52];
    86: op1_04_in28 = reg_0356;
    87: op1_04_in28 = reg_0496;
    88: op1_04_in28 = reg_0091;
    90: op1_04_in28 = reg_0407;
    91: op1_04_in28 = reg_0495;
    default: op1_04_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_04_inv28 = 1;
    9: op1_04_inv28 = 1;
    11: op1_04_inv28 = 1;
    15: op1_04_inv28 = 1;
    20: op1_04_inv28 = 1;
    22: op1_04_inv28 = 1;
    24: op1_04_inv28 = 1;
    25: op1_04_inv28 = 1;
    28: op1_04_inv28 = 1;
    30: op1_04_inv28 = 1;
    35: op1_04_inv28 = 1;
    37: op1_04_inv28 = 1;
    45: op1_04_inv28 = 1;
    47: op1_04_inv28 = 1;
    48: op1_04_inv28 = 1;
    49: op1_04_inv28 = 1;
    52: op1_04_inv28 = 1;
    53: op1_04_inv28 = 1;
    57: op1_04_inv28 = 1;
    58: op1_04_inv28 = 1;
    60: op1_04_inv28 = 1;
    62: op1_04_inv28 = 1;
    63: op1_04_inv28 = 1;
    64: op1_04_inv28 = 1;
    65: op1_04_inv28 = 1;
    67: op1_04_inv28 = 1;
    69: op1_04_inv28 = 1;
    71: op1_04_inv28 = 1;
    77: op1_04_inv28 = 1;
    82: op1_04_inv28 = 1;
    86: op1_04_inv28 = 1;
    87: op1_04_inv28 = 1;
    88: op1_04_inv28 = 1;
    89: op1_04_inv28 = 1;
    90: op1_04_inv28 = 1;
    96: op1_04_inv28 = 1;
    default: op1_04_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in29 = reg_0356;
    6: op1_04_in29 = reg_0221;
    7: op1_04_in29 = reg_0494;
    8: op1_04_in29 = reg_0730;
    9: op1_04_in29 = imem06_in[87:84];
    11: op1_04_in29 = reg_0038;
    67: op1_04_in29 = reg_0038;
    12: op1_04_in29 = reg_0648;
    13: op1_04_in29 = imem05_in[95:92];
    14: op1_04_in29 = reg_0029;
    15: op1_04_in29 = reg_0219;
    16: op1_04_in29 = reg_0319;
    18: op1_04_in29 = imem04_in[15:12];
    19: op1_04_in29 = reg_0425;
    20: op1_04_in29 = reg_0811;
    21: op1_04_in29 = reg_0707;
    23: op1_04_in29 = imem06_in[7:4];
    24: op1_04_in29 = imem01_in[123:120];
    25: op1_04_in29 = reg_0373;
    26: op1_04_in29 = reg_0113;
    27: op1_04_in29 = reg_0770;
    28: op1_04_in29 = reg_0165;
    30: op1_04_in29 = imem03_in[55:52];
    31: op1_04_in29 = reg_0813;
    32: op1_04_in29 = reg_0183;
    33: op1_04_in29 = imem02_in[67:64];
    34: op1_04_in29 = reg_0721;
    35: op1_04_in29 = reg_0153;
    36: op1_04_in29 = reg_0713;
    37: op1_04_in29 = reg_0438;
    39: op1_04_in29 = imem01_in[55:52];
    41: op1_04_in29 = reg_0061;
    42: op1_04_in29 = reg_0818;
    44: op1_04_in29 = reg_0566;
    45: op1_04_in29 = reg_0791;
    47: op1_04_in29 = imem01_in[115:112];
    48: op1_04_in29 = reg_0744;
    49: op1_04_in29 = imem04_in[55:52];
    50: op1_04_in29 = imem03_in[79:76];
    53: op1_04_in29 = imem03_in[79:76];
    52: op1_04_in29 = imem01_in[75:72];
    54: op1_04_in29 = imem04_in[95:92];
    55: op1_04_in29 = reg_0076;
    56: op1_04_in29 = reg_0136;
    57: op1_04_in29 = reg_0621;
    58: op1_04_in29 = reg_0797;
    60: op1_04_in29 = reg_0253;
    62: op1_04_in29 = imem03_in[103:100];
    63: op1_04_in29 = reg_0803;
    64: op1_04_in29 = imem05_in[99:96];
    65: op1_04_in29 = imem05_in[23:20];
    66: op1_04_in29 = reg_0430;
    68: op1_04_in29 = reg_0422;
    69: op1_04_in29 = reg_0007;
    70: op1_04_in29 = reg_0619;
    71: op1_04_in29 = reg_0395;
    72: op1_04_in29 = reg_0615;
    73: op1_04_in29 = reg_0215;
    74: op1_04_in29 = reg_0787;
    77: op1_04_in29 = reg_0248;
    78: op1_04_in29 = reg_0316;
    79: op1_04_in29 = reg_0719;
    80: op1_04_in29 = reg_0659;
    81: op1_04_in29 = reg_0155;
    82: op1_04_in29 = reg_0592;
    84: op1_04_in29 = reg_0065;
    85: op1_04_in29 = imem07_in[111:108];
    86: op1_04_in29 = reg_0363;
    87: op1_04_in29 = reg_0006;
    89: op1_04_in29 = reg_0667;
    90: op1_04_in29 = reg_0531;
    91: op1_04_in29 = reg_0407;
    96: op1_04_in29 = reg_0680;
    default: op1_04_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_04_inv29 = 1;
    8: op1_04_inv29 = 1;
    9: op1_04_inv29 = 1;
    11: op1_04_inv29 = 1;
    12: op1_04_inv29 = 1;
    13: op1_04_inv29 = 1;
    16: op1_04_inv29 = 1;
    18: op1_04_inv29 = 1;
    19: op1_04_inv29 = 1;
    21: op1_04_inv29 = 1;
    25: op1_04_inv29 = 1;
    26: op1_04_inv29 = 1;
    28: op1_04_inv29 = 1;
    30: op1_04_inv29 = 1;
    33: op1_04_inv29 = 1;
    34: op1_04_inv29 = 1;
    36: op1_04_inv29 = 1;
    39: op1_04_inv29 = 1;
    42: op1_04_inv29 = 1;
    48: op1_04_inv29 = 1;
    49: op1_04_inv29 = 1;
    53: op1_04_inv29 = 1;
    54: op1_04_inv29 = 1;
    55: op1_04_inv29 = 1;
    58: op1_04_inv29 = 1;
    60: op1_04_inv29 = 1;
    62: op1_04_inv29 = 1;
    63: op1_04_inv29 = 1;
    64: op1_04_inv29 = 1;
    65: op1_04_inv29 = 1;
    66: op1_04_inv29 = 1;
    67: op1_04_inv29 = 1;
    69: op1_04_inv29 = 1;
    71: op1_04_inv29 = 1;
    72: op1_04_inv29 = 1;
    77: op1_04_inv29 = 1;
    78: op1_04_inv29 = 1;
    84: op1_04_inv29 = 1;
    86: op1_04_inv29 = 1;
    89: op1_04_inv29 = 1;
    90: op1_04_inv29 = 1;
    96: op1_04_inv29 = 1;
    default: op1_04_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_04_in30 = reg_0382;
    6: op1_04_in30 = reg_0123;
    7: op1_04_in30 = reg_0780;
    8: op1_04_in30 = reg_0731;
    9: op1_04_in30 = imem06_in[99:96];
    11: op1_04_in30 = imem07_in[31:28];
    12: op1_04_in30 = reg_0643;
    13: op1_04_in30 = imem05_in[107:104];
    14: op1_04_in30 = reg_0038;
    15: op1_04_in30 = reg_0249;
    16: op1_04_in30 = reg_0385;
    18: op1_04_in30 = imem04_in[35:32];
    19: op1_04_in30 = reg_0436;
    20: op1_04_in30 = reg_0003;
    21: op1_04_in30 = reg_0426;
    23: op1_04_in30 = imem06_in[95:92];
    24: op1_04_in30 = reg_0232;
    25: op1_04_in30 = reg_0804;
    26: op1_04_in30 = reg_0110;
    58: op1_04_in30 = reg_0110;
    27: op1_04_in30 = reg_0757;
    28: op1_04_in30 = reg_0162;
    30: op1_04_in30 = imem03_in[75:72];
    31: op1_04_in30 = reg_0005;
    32: op1_04_in30 = reg_0185;
    33: op1_04_in30 = imem02_in[83:80];
    34: op1_04_in30 = reg_0714;
    35: op1_04_in30 = reg_0614;
    36: op1_04_in30 = reg_0718;
    37: op1_04_in30 = reg_0448;
    39: op1_04_in30 = imem01_in[111:108];
    41: op1_04_in30 = reg_0253;
    42: op1_04_in30 = reg_0246;
    44: op1_04_in30 = reg_0587;
    45: op1_04_in30 = reg_0798;
    47: op1_04_in30 = imem01_in[119:116];
    48: op1_04_in30 = reg_0285;
    79: op1_04_in30 = reg_0285;
    49: op1_04_in30 = imem04_in[119:116];
    50: op1_04_in30 = imem03_in[111:108];
    52: op1_04_in30 = imem01_in[87:84];
    53: op1_04_in30 = imem03_in[87:84];
    54: op1_04_in30 = imem04_in[103:100];
    55: op1_04_in30 = reg_0529;
    56: op1_04_in30 = reg_0133;
    57: op1_04_in30 = reg_0029;
    60: op1_04_in30 = reg_0333;
    62: op1_04_in30 = reg_0559;
    63: op1_04_in30 = reg_0007;
    64: op1_04_in30 = imem05_in[123:120];
    65: op1_04_in30 = imem05_in[71:68];
    66: op1_04_in30 = reg_0617;
    67: op1_04_in30 = reg_0628;
    68: op1_04_in30 = reg_0219;
    69: op1_04_in30 = reg_0801;
    70: op1_04_in30 = reg_0238;
    71: op1_04_in30 = reg_0483;
    72: op1_04_in30 = reg_0611;
    73: op1_04_in30 = reg_0486;
    74: op1_04_in30 = reg_0767;
    77: op1_04_in30 = reg_0506;
    78: op1_04_in30 = reg_0544;
    80: op1_04_in30 = reg_0773;
    81: op1_04_in30 = reg_0137;
    82: op1_04_in30 = imem02_in[7:4];
    84: op1_04_in30 = reg_0622;
    85: op1_04_in30 = reg_0716;
    86: op1_04_in30 = reg_0594;
    87: op1_04_in30 = reg_0805;
    89: op1_04_in30 = reg_0788;
    90: op1_04_in30 = reg_0254;
    91: op1_04_in30 = reg_0393;
    96: op1_04_in30 = reg_0661;
    default: op1_04_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_04_inv30 = 1;
    7: op1_04_inv30 = 1;
    9: op1_04_inv30 = 1;
    13: op1_04_inv30 = 1;
    15: op1_04_inv30 = 1;
    16: op1_04_inv30 = 1;
    18: op1_04_inv30 = 1;
    19: op1_04_inv30 = 1;
    23: op1_04_inv30 = 1;
    25: op1_04_inv30 = 1;
    27: op1_04_inv30 = 1;
    28: op1_04_inv30 = 1;
    30: op1_04_inv30 = 1;
    31: op1_04_inv30 = 1;
    34: op1_04_inv30 = 1;
    36: op1_04_inv30 = 1;
    37: op1_04_inv30 = 1;
    39: op1_04_inv30 = 1;
    41: op1_04_inv30 = 1;
    42: op1_04_inv30 = 1;
    47: op1_04_inv30 = 1;
    49: op1_04_inv30 = 1;
    50: op1_04_inv30 = 1;
    52: op1_04_inv30 = 1;
    53: op1_04_inv30 = 1;
    54: op1_04_inv30 = 1;
    56: op1_04_inv30 = 1;
    57: op1_04_inv30 = 1;
    62: op1_04_inv30 = 1;
    64: op1_04_inv30 = 1;
    67: op1_04_inv30 = 1;
    68: op1_04_inv30 = 1;
    69: op1_04_inv30 = 1;
    71: op1_04_inv30 = 1;
    72: op1_04_inv30 = 1;
    74: op1_04_inv30 = 1;
    77: op1_04_inv30 = 1;
    78: op1_04_inv30 = 1;
    81: op1_04_inv30 = 1;
    82: op1_04_inv30 = 1;
    85: op1_04_inv30 = 1;
    86: op1_04_inv30 = 1;
    87: op1_04_inv30 = 1;
    96: op1_04_inv30 = 1;
    default: op1_04_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_04_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_04_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in00 = imem00_in[31:28];
    10: op1_05_in00 = imem00_in[31:28];
    94: op1_05_in00 = imem00_in[31:28];
    5: op1_05_in00 = reg_0315;
    6: op1_05_in00 = reg_0122;
    7: op1_05_in00 = reg_0495;
    8: op1_05_in00 = imem00_in[55:52];
    76: op1_05_in00 = imem00_in[55:52];
    9: op1_05_in00 = reg_0630;
    11: op1_05_in00 = imem07_in[75:72];
    3: op1_05_in00 = imem07_in[47:44];
    12: op1_05_in00 = reg_0667;
    13: op1_05_in00 = imem05_in[127:124];
    14: op1_05_in00 = imem07_in[7:4];
    2: op1_05_in00 = imem07_in[7:4];
    96: op1_05_in00 = imem07_in[7:4];
    15: op1_05_in00 = reg_0124;
    16: op1_05_in00 = reg_0377;
    17: op1_05_in00 = imem00_in[7:4];
    22: op1_05_in00 = imem00_in[7:4];
    29: op1_05_in00 = imem00_in[7:4];
    61: op1_05_in00 = imem00_in[7:4];
    18: op1_05_in00 = imem04_in[51:48];
    19: op1_05_in00 = imem00_in[27:24];
    21: op1_05_in00 = imem00_in[27:24];
    20: op1_05_in00 = reg_0004;
    23: op1_05_in00 = imem06_in[127:124];
    1: op1_05_in00 = imem07_in[63:60];
    24: op1_05_in00 = reg_0246;
    25: op1_05_in00 = reg_0802;
    26: op1_05_in00 = imem02_in[7:4];
    27: op1_05_in00 = reg_0038;
    28: op1_05_in00 = imem00_in[67:64];
    30: op1_05_in00 = reg_0391;
    31: op1_05_in00 = reg_0614;
    32: op1_05_in00 = imem00_in[3:0];
    92: op1_05_in00 = imem00_in[3:0];
    33: op1_05_in00 = imem02_in[99:96];
    34: op1_05_in00 = reg_0711;
    36: op1_05_in00 = reg_0711;
    35: op1_05_in00 = reg_0029;
    37: op1_05_in00 = reg_0172;
    38: op1_05_in00 = imem00_in[95:92];
    39: op1_05_in00 = reg_0116;
    40: op1_05_in00 = imem00_in[35:32];
    46: op1_05_in00 = imem00_in[35:32];
    88: op1_05_in00 = imem00_in[35:32];
    41: op1_05_in00 = reg_0066;
    42: op1_05_in00 = reg_0249;
    43: op1_05_in00 = imem00_in[47:44];
    44: op1_05_in00 = reg_0585;
    45: op1_05_in00 = reg_0483;
    47: op1_05_in00 = reg_0511;
    48: op1_05_in00 = reg_0152;
    49: op1_05_in00 = imem04_in[127:124];
    50: op1_05_in00 = imem03_in[127:124];
    51: op1_05_in00 = imem00_in[15:12];
    75: op1_05_in00 = imem00_in[15:12];
    83: op1_05_in00 = imem00_in[15:12];
    52: op1_05_in00 = imem01_in[95:92];
    53: op1_05_in00 = imem03_in[99:96];
    54: op1_05_in00 = imem04_in[111:108];
    55: op1_05_in00 = reg_0611;
    56: op1_05_in00 = reg_0142;
    57: op1_05_in00 = reg_0236;
    58: op1_05_in00 = reg_0111;
    59: op1_05_in00 = imem00_in[39:36];
    60: op1_05_in00 = reg_0434;
    62: op1_05_in00 = reg_0318;
    63: op1_05_in00 = reg_0799;
    64: op1_05_in00 = reg_0103;
    65: op1_05_in00 = imem05_in[83:80];
    66: op1_05_in00 = reg_0626;
    67: op1_05_in00 = reg_0369;
    90: op1_05_in00 = reg_0369;
    68: op1_05_in00 = reg_0673;
    69: op1_05_in00 = reg_0015;
    70: op1_05_in00 = reg_0293;
    71: op1_05_in00 = reg_0803;
    72: op1_05_in00 = reg_0302;
    73: op1_05_in00 = imem05_in[51:48];
    74: op1_05_in00 = reg_0661;
    77: op1_05_in00 = reg_0073;
    78: op1_05_in00 = reg_0553;
    79: op1_05_in00 = reg_0148;
    80: op1_05_in00 = reg_0821;
    81: op1_05_in00 = reg_0734;
    82: op1_05_in00 = imem02_in[35:32];
    84: op1_05_in00 = reg_0780;
    85: op1_05_in00 = reg_0163;
    86: op1_05_in00 = reg_0406;
    87: op1_05_in00 = reg_0016;
    89: op1_05_in00 = reg_0793;
    91: op1_05_in00 = reg_0579;
    93: op1_05_in00 = imem00_in[43:40];
    95: op1_05_in00 = imem00_in[103:100];
    default: op1_05_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv00 = 1;
    5: op1_05_inv00 = 1;
    6: op1_05_inv00 = 1;
    7: op1_05_inv00 = 1;
    8: op1_05_inv00 = 1;
    11: op1_05_inv00 = 1;
    14: op1_05_inv00 = 1;
    19: op1_05_inv00 = 1;
    20: op1_05_inv00 = 1;
    24: op1_05_inv00 = 1;
    25: op1_05_inv00 = 1;
    27: op1_05_inv00 = 1;
    28: op1_05_inv00 = 1;
    29: op1_05_inv00 = 1;
    30: op1_05_inv00 = 1;
    31: op1_05_inv00 = 1;
    34: op1_05_inv00 = 1;
    40: op1_05_inv00 = 1;
    42: op1_05_inv00 = 1;
    43: op1_05_inv00 = 1;
    45: op1_05_inv00 = 1;
    47: op1_05_inv00 = 1;
    49: op1_05_inv00 = 1;
    50: op1_05_inv00 = 1;
    51: op1_05_inv00 = 1;
    52: op1_05_inv00 = 1;
    54: op1_05_inv00 = 1;
    56: op1_05_inv00 = 1;
    57: op1_05_inv00 = 1;
    58: op1_05_inv00 = 1;
    59: op1_05_inv00 = 1;
    61: op1_05_inv00 = 1;
    63: op1_05_inv00 = 1;
    65: op1_05_inv00 = 1;
    67: op1_05_inv00 = 1;
    69: op1_05_inv00 = 1;
    70: op1_05_inv00 = 1;
    73: op1_05_inv00 = 1;
    76: op1_05_inv00 = 1;
    77: op1_05_inv00 = 1;
    79: op1_05_inv00 = 1;
    80: op1_05_inv00 = 1;
    83: op1_05_inv00 = 1;
    84: op1_05_inv00 = 1;
    85: op1_05_inv00 = 1;
    89: op1_05_inv00 = 1;
    90: op1_05_inv00 = 1;
    91: op1_05_inv00 = 1;
    96: op1_05_inv00 = 1;
    default: op1_05_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in01 = imem00_in[35:32];
    22: op1_05_in01 = imem00_in[35:32];
    5: op1_05_in01 = reg_0390;
    6: op1_05_in01 = imem02_in[3:0];
    7: op1_05_in01 = reg_0794;
    8: op1_05_in01 = imem00_in[79:76];
    9: op1_05_in01 = reg_0613;
    10: op1_05_in01 = imem00_in[47:44];
    46: op1_05_in01 = imem00_in[47:44];
    11: op1_05_in01 = imem07_in[123:120];
    3: op1_05_in01 = imem07_in[59:56];
    57: op1_05_in01 = imem07_in[59:56];
    12: op1_05_in01 = reg_0339;
    13: op1_05_in01 = reg_0482;
    14: op1_05_in01 = imem07_in[23:20];
    15: op1_05_in01 = reg_0125;
    77: op1_05_in01 = reg_0125;
    16: op1_05_in01 = reg_0361;
    17: op1_05_in01 = reg_0682;
    18: op1_05_in01 = imem04_in[59:56];
    2: op1_05_in01 = imem07_in[19:16];
    19: op1_05_in01 = imem00_in[99:96];
    38: op1_05_in01 = imem00_in[99:96];
    20: op1_05_in01 = imem04_in[35:32];
    21: op1_05_in01 = imem00_in[51:48];
    43: op1_05_in01 = imem00_in[51:48];
    88: op1_05_in01 = imem00_in[51:48];
    23: op1_05_in01 = reg_0607;
    1: op1_05_in01 = imem07_in[83:80];
    24: op1_05_in01 = reg_0218;
    25: op1_05_in01 = reg_0809;
    26: op1_05_in01 = imem02_in[11:8];
    27: op1_05_in01 = reg_0370;
    28: op1_05_in01 = imem00_in[75:72];
    29: op1_05_in01 = imem00_in[27:24];
    75: op1_05_in01 = imem00_in[27:24];
    30: op1_05_in01 = reg_0561;
    31: op1_05_in01 = reg_0628;
    70: op1_05_in01 = reg_0628;
    32: op1_05_in01 = imem00_in[19:16];
    51: op1_05_in01 = imem00_in[19:16];
    83: op1_05_in01 = imem00_in[19:16];
    33: op1_05_in01 = imem02_in[123:120];
    34: op1_05_in01 = reg_0426;
    35: op1_05_in01 = reg_0037;
    36: op1_05_in01 = reg_0424;
    37: op1_05_in01 = reg_0162;
    39: op1_05_in01 = reg_0100;
    40: op1_05_in01 = imem00_in[39:36];
    41: op1_05_in01 = imem05_in[79:76];
    42: op1_05_in01 = reg_0237;
    44: op1_05_in01 = reg_0600;
    45: op1_05_in01 = reg_0490;
    47: op1_05_in01 = reg_0422;
    48: op1_05_in01 = reg_0138;
    49: op1_05_in01 = reg_0544;
    54: op1_05_in01 = reg_0544;
    50: op1_05_in01 = reg_0602;
    52: op1_05_in01 = imem02_in[35:32];
    53: op1_05_in01 = imem03_in[107:104];
    55: op1_05_in01 = reg_0071;
    56: op1_05_in01 = reg_0139;
    58: op1_05_in01 = reg_0790;
    59: op1_05_in01 = imem00_in[43:40];
    60: op1_05_in01 = reg_0449;
    61: op1_05_in01 = reg_0693;
    62: op1_05_in01 = reg_0528;
    63: op1_05_in01 = imem04_in[55:52];
    64: op1_05_in01 = reg_0279;
    65: op1_05_in01 = imem05_in[127:124];
    66: op1_05_in01 = reg_0610;
    67: op1_05_in01 = reg_0659;
    68: op1_05_in01 = reg_0120;
    69: op1_05_in01 = reg_0016;
    71: op1_05_in01 = reg_0807;
    72: op1_05_in01 = reg_0616;
    73: op1_05_in01 = imem05_in[95:92];
    74: op1_05_in01 = reg_0716;
    76: op1_05_in01 = imem00_in[59:56];
    94: op1_05_in01 = imem00_in[59:56];
    78: op1_05_in01 = reg_0060;
    79: op1_05_in01 = reg_0827;
    80: op1_05_in01 = reg_0748;
    81: op1_05_in01 = imem06_in[7:4];
    82: op1_05_in01 = imem02_in[63:60];
    84: op1_05_in01 = reg_0513;
    85: op1_05_in01 = reg_0166;
    86: op1_05_in01 = reg_0514;
    87: op1_05_in01 = imem04_in[71:68];
    89: op1_05_in01 = reg_0090;
    90: op1_05_in01 = reg_0579;
    91: op1_05_in01 = reg_0150;
    92: op1_05_in01 = imem00_in[11:8];
    93: op1_05_in01 = imem00_in[87:84];
    95: op1_05_in01 = reg_0112;
    96: op1_05_in01 = imem07_in[39:36];
    default: op1_05_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv01 = 1;
    9: op1_05_inv01 = 1;
    11: op1_05_inv01 = 1;
    12: op1_05_inv01 = 1;
    13: op1_05_inv01 = 1;
    14: op1_05_inv01 = 1;
    15: op1_05_inv01 = 1;
    16: op1_05_inv01 = 1;
    18: op1_05_inv01 = 1;
    21: op1_05_inv01 = 1;
    23: op1_05_inv01 = 1;
    1: op1_05_inv01 = 1;
    24: op1_05_inv01 = 1;
    25: op1_05_inv01 = 1;
    27: op1_05_inv01 = 1;
    28: op1_05_inv01 = 1;
    29: op1_05_inv01 = 1;
    30: op1_05_inv01 = 1;
    31: op1_05_inv01 = 1;
    35: op1_05_inv01 = 1;
    39: op1_05_inv01 = 1;
    41: op1_05_inv01 = 1;
    42: op1_05_inv01 = 1;
    45: op1_05_inv01 = 1;
    46: op1_05_inv01 = 1;
    47: op1_05_inv01 = 1;
    48: op1_05_inv01 = 1;
    53: op1_05_inv01 = 1;
    57: op1_05_inv01 = 1;
    58: op1_05_inv01 = 1;
    59: op1_05_inv01 = 1;
    61: op1_05_inv01 = 1;
    62: op1_05_inv01 = 1;
    63: op1_05_inv01 = 1;
    64: op1_05_inv01 = 1;
    65: op1_05_inv01 = 1;
    67: op1_05_inv01 = 1;
    70: op1_05_inv01 = 1;
    71: op1_05_inv01 = 1;
    72: op1_05_inv01 = 1;
    74: op1_05_inv01 = 1;
    76: op1_05_inv01 = 1;
    79: op1_05_inv01 = 1;
    83: op1_05_inv01 = 1;
    85: op1_05_inv01 = 1;
    86: op1_05_inv01 = 1;
    88: op1_05_inv01 = 1;
    89: op1_05_inv01 = 1;
    90: op1_05_inv01 = 1;
    93: op1_05_inv01 = 1;
    94: op1_05_inv01 = 1;
    96: op1_05_inv01 = 1;
    default: op1_05_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in02 = imem00_in[51:48];
    5: op1_05_in02 = reg_0034;
    6: op1_05_in02 = imem02_in[11:8];
    7: op1_05_in02 = reg_0267;
    8: op1_05_in02 = imem00_in[123:120];
    9: op1_05_in02 = reg_0620;
    10: op1_05_in02 = imem00_in[59:56];
    11: op1_05_in02 = reg_0729;
    3: op1_05_in02 = imem07_in[95:92];
    12: op1_05_in02 = reg_0324;
    13: op1_05_in02 = reg_0484;
    14: op1_05_in02 = imem07_in[31:28];
    15: op1_05_in02 = reg_0115;
    16: op1_05_in02 = reg_0396;
    17: op1_05_in02 = reg_0696;
    76: op1_05_in02 = reg_0696;
    18: op1_05_in02 = imem04_in[63:60];
    2: op1_05_in02 = imem07_in[35:32];
    19: op1_05_in02 = reg_0684;
    20: op1_05_in02 = imem04_in[47:44];
    21: op1_05_in02 = imem00_in[55:52];
    43: op1_05_in02 = imem00_in[55:52];
    22: op1_05_in02 = imem00_in[39:36];
    23: op1_05_in02 = reg_0624;
    31: op1_05_in02 = reg_0624;
    24: op1_05_in02 = reg_0220;
    25: op1_05_in02 = imem04_in[15:12];
    26: op1_05_in02 = imem02_in[15:12];
    27: op1_05_in02 = reg_0369;
    28: op1_05_in02 = imem00_in[95:92];
    29: op1_05_in02 = imem00_in[87:84];
    30: op1_05_in02 = reg_0755;
    32: op1_05_in02 = imem00_in[43:40];
    33: op1_05_in02 = reg_0642;
    34: op1_05_in02 = reg_0443;
    35: op1_05_in02 = imem06_in[27:24];
    36: op1_05_in02 = reg_0429;
    37: op1_05_in02 = reg_0167;
    38: op1_05_in02 = reg_0693;
    39: op1_05_in02 = imem02_in[87:84];
    40: op1_05_in02 = imem00_in[115:112];
    41: op1_05_in02 = imem05_in[115:112];
    73: op1_05_in02 = imem05_in[115:112];
    42: op1_05_in02 = reg_0427;
    44: op1_05_in02 = reg_0597;
    45: op1_05_in02 = reg_0491;
    46: op1_05_in02 = imem00_in[67:64];
    94: op1_05_in02 = imem00_in[67:64];
    47: op1_05_in02 = reg_0504;
    48: op1_05_in02 = reg_0153;
    49: op1_05_in02 = reg_0553;
    50: op1_05_in02 = reg_0599;
    51: op1_05_in02 = imem00_in[91:88];
    52: op1_05_in02 = imem02_in[91:88];
    53: op1_05_in02 = reg_0391;
    54: op1_05_in02 = reg_0542;
    55: op1_05_in02 = reg_0508;
    56: op1_05_in02 = reg_0131;
    57: op1_05_in02 = reg_0441;
    58: op1_05_in02 = reg_0218;
    59: op1_05_in02 = imem00_in[83:80];
    60: op1_05_in02 = reg_0437;
    61: op1_05_in02 = reg_0683;
    62: op1_05_in02 = reg_0331;
    63: op1_05_in02 = imem04_in[67:64];
    64: op1_05_in02 = reg_0249;
    65: op1_05_in02 = reg_0152;
    66: op1_05_in02 = reg_0779;
    67: op1_05_in02 = reg_0816;
    68: op1_05_in02 = reg_0660;
    69: op1_05_in02 = imem04_in[3:0];
    70: op1_05_in02 = imem06_in[3:0];
    71: op1_05_in02 = reg_0805;
    72: op1_05_in02 = reg_0629;
    74: op1_05_in02 = reg_0089;
    75: op1_05_in02 = imem00_in[63:60];
    77: op1_05_in02 = reg_0670;
    78: op1_05_in02 = reg_0510;
    79: op1_05_in02 = reg_0785;
    80: op1_05_in02 = reg_0270;
    81: op1_05_in02 = imem06_in[11:8];
    82: op1_05_in02 = imem02_in[67:64];
    83: op1_05_in02 = imem00_in[27:24];
    84: op1_05_in02 = imem05_in[3:0];
    85: op1_05_in02 = reg_0713;
    86: op1_05_in02 = reg_0323;
    87: op1_05_in02 = imem04_in[91:88];
    88: op1_05_in02 = imem00_in[75:72];
    89: op1_05_in02 = reg_0027;
    90: op1_05_in02 = reg_0560;
    91: op1_05_in02 = reg_0765;
    92: op1_05_in02 = imem00_in[19:16];
    93: op1_05_in02 = reg_0689;
    95: op1_05_in02 = reg_0686;
    96: op1_05_in02 = imem07_in[103:100];
    default: op1_05_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv02 = 1;
    10: op1_05_inv02 = 1;
    12: op1_05_inv02 = 1;
    15: op1_05_inv02 = 1;
    16: op1_05_inv02 = 1;
    17: op1_05_inv02 = 1;
    18: op1_05_inv02 = 1;
    19: op1_05_inv02 = 1;
    21: op1_05_inv02 = 1;
    22: op1_05_inv02 = 1;
    23: op1_05_inv02 = 1;
    25: op1_05_inv02 = 1;
    26: op1_05_inv02 = 1;
    27: op1_05_inv02 = 1;
    28: op1_05_inv02 = 1;
    29: op1_05_inv02 = 1;
    30: op1_05_inv02 = 1;
    34: op1_05_inv02 = 1;
    37: op1_05_inv02 = 1;
    39: op1_05_inv02 = 1;
    40: op1_05_inv02 = 1;
    42: op1_05_inv02 = 1;
    43: op1_05_inv02 = 1;
    44: op1_05_inv02 = 1;
    45: op1_05_inv02 = 1;
    48: op1_05_inv02 = 1;
    49: op1_05_inv02 = 1;
    51: op1_05_inv02 = 1;
    52: op1_05_inv02 = 1;
    53: op1_05_inv02 = 1;
    54: op1_05_inv02 = 1;
    55: op1_05_inv02 = 1;
    58: op1_05_inv02 = 1;
    59: op1_05_inv02 = 1;
    62: op1_05_inv02 = 1;
    63: op1_05_inv02 = 1;
    65: op1_05_inv02 = 1;
    67: op1_05_inv02 = 1;
    69: op1_05_inv02 = 1;
    70: op1_05_inv02 = 1;
    71: op1_05_inv02 = 1;
    73: op1_05_inv02 = 1;
    74: op1_05_inv02 = 1;
    76: op1_05_inv02 = 1;
    77: op1_05_inv02 = 1;
    78: op1_05_inv02 = 1;
    81: op1_05_inv02 = 1;
    82: op1_05_inv02 = 1;
    85: op1_05_inv02 = 1;
    88: op1_05_inv02 = 1;
    90: op1_05_inv02 = 1;
    91: op1_05_inv02 = 1;
    92: op1_05_inv02 = 1;
    94: op1_05_inv02 = 1;
    96: op1_05_inv02 = 1;
    default: op1_05_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in03 = imem00_in[55:52];
    83: op1_05_in03 = imem00_in[55:52];
    5: op1_05_in03 = reg_0035;
    6: op1_05_in03 = imem02_in[19:16];
    7: op1_05_in03 = reg_0271;
    8: op1_05_in03 = reg_0681;
    9: op1_05_in03 = reg_0617;
    55: op1_05_in03 = reg_0617;
    10: op1_05_in03 = imem00_in[99:96];
    11: op1_05_in03 = reg_0713;
    3: op1_05_in03 = reg_0424;
    12: op1_05_in03 = reg_0083;
    13: op1_05_in03 = reg_0788;
    14: op1_05_in03 = imem07_in[39:36];
    15: op1_05_in03 = reg_0113;
    16: op1_05_in03 = reg_0374;
    17: op1_05_in03 = reg_0672;
    18: op1_05_in03 = imem04_in[95:92];
    87: op1_05_in03 = imem04_in[95:92];
    2: op1_05_in03 = imem07_in[59:56];
    19: op1_05_in03 = reg_0690;
    88: op1_05_in03 = reg_0690;
    95: op1_05_in03 = reg_0690;
    20: op1_05_in03 = imem04_in[67:64];
    21: op1_05_in03 = imem00_in[91:88];
    22: op1_05_in03 = imem00_in[43:40];
    23: op1_05_in03 = reg_0620;
    24: op1_05_in03 = reg_0116;
    25: op1_05_in03 = imem04_in[19:16];
    26: op1_05_in03 = imem02_in[51:48];
    27: op1_05_in03 = reg_0264;
    28: op1_05_in03 = imem00_in[103:100];
    29: op1_05_in03 = imem00_in[127:124];
    30: op1_05_in03 = reg_0373;
    31: op1_05_in03 = reg_0613;
    32: op1_05_in03 = imem00_in[47:44];
    33: op1_05_in03 = reg_0656;
    34: op1_05_in03 = reg_0181;
    35: op1_05_in03 = imem06_in[55:52];
    36: op1_05_in03 = reg_0432;
    37: op1_05_in03 = reg_0163;
    38: op1_05_in03 = reg_0697;
    39: op1_05_in03 = imem02_in[111:108];
    40: op1_05_in03 = reg_0696;
    41: op1_05_in03 = imem05_in[123:120];
    42: op1_05_in03 = reg_0717;
    43: op1_05_in03 = imem00_in[67:64];
    44: op1_05_in03 = reg_0395;
    45: op1_05_in03 = reg_0492;
    61: op1_05_in03 = reg_0492;
    46: op1_05_in03 = imem00_in[83:80];
    47: op1_05_in03 = reg_0103;
    48: op1_05_in03 = reg_0141;
    49: op1_05_in03 = reg_0552;
    50: op1_05_in03 = reg_0583;
    67: op1_05_in03 = reg_0583;
    80: op1_05_in03 = reg_0583;
    51: op1_05_in03 = reg_0682;
    52: op1_05_in03 = imem02_in[103:100];
    53: op1_05_in03 = reg_0572;
    54: op1_05_in03 = reg_0088;
    56: op1_05_in03 = imem06_in[47:44];
    57: op1_05_in03 = reg_0266;
    58: op1_05_in03 = reg_0486;
    59: op1_05_in03 = imem00_in[107:104];
    60: op1_05_in03 = reg_0267;
    62: op1_05_in03 = reg_0387;
    63: op1_05_in03 = imem04_in[111:108];
    64: op1_05_in03 = reg_0307;
    65: op1_05_in03 = reg_0156;
    66: op1_05_in03 = reg_0622;
    68: op1_05_in03 = reg_0676;
    69: op1_05_in03 = imem04_in[31:28];
    70: op1_05_in03 = imem06_in[31:28];
    71: op1_05_in03 = reg_0008;
    72: op1_05_in03 = reg_0078;
    73: op1_05_in03 = imem06_in[7:4];
    74: op1_05_in03 = reg_0391;
    75: op1_05_in03 = reg_0685;
    76: op1_05_in03 = reg_0686;
    77: op1_05_in03 = reg_0108;
    78: op1_05_in03 = reg_0556;
    79: op1_05_in03 = reg_0742;
    81: op1_05_in03 = imem06_in[23:20];
    82: op1_05_in03 = imem02_in[115:112];
    84: op1_05_in03 = imem05_in[11:8];
    85: op1_05_in03 = reg_0334;
    86: op1_05_in03 = reg_0092;
    89: op1_05_in03 = reg_0488;
    90: op1_05_in03 = reg_0149;
    91: op1_05_in03 = reg_0824;
    92: op1_05_in03 = imem00_in[31:28];
    93: op1_05_in03 = reg_0130;
    94: op1_05_in03 = imem00_in[79:76];
    96: op1_05_in03 = imem07_in[107:104];
    default: op1_05_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv03 = 1;
    6: op1_05_inv03 = 1;
    7: op1_05_inv03 = 1;
    8: op1_05_inv03 = 1;
    9: op1_05_inv03 = 1;
    10: op1_05_inv03 = 1;
    11: op1_05_inv03 = 1;
    13: op1_05_inv03 = 1;
    15: op1_05_inv03 = 1;
    17: op1_05_inv03 = 1;
    20: op1_05_inv03 = 1;
    22: op1_05_inv03 = 1;
    25: op1_05_inv03 = 1;
    26: op1_05_inv03 = 1;
    30: op1_05_inv03 = 1;
    32: op1_05_inv03 = 1;
    37: op1_05_inv03 = 1;
    40: op1_05_inv03 = 1;
    47: op1_05_inv03 = 1;
    48: op1_05_inv03 = 1;
    50: op1_05_inv03 = 1;
    51: op1_05_inv03 = 1;
    52: op1_05_inv03 = 1;
    54: op1_05_inv03 = 1;
    57: op1_05_inv03 = 1;
    59: op1_05_inv03 = 1;
    60: op1_05_inv03 = 1;
    62: op1_05_inv03 = 1;
    63: op1_05_inv03 = 1;
    64: op1_05_inv03 = 1;
    66: op1_05_inv03 = 1;
    68: op1_05_inv03 = 1;
    69: op1_05_inv03 = 1;
    71: op1_05_inv03 = 1;
    72: op1_05_inv03 = 1;
    73: op1_05_inv03 = 1;
    74: op1_05_inv03 = 1;
    78: op1_05_inv03 = 1;
    82: op1_05_inv03 = 1;
    83: op1_05_inv03 = 1;
    85: op1_05_inv03 = 1;
    87: op1_05_inv03 = 1;
    88: op1_05_inv03 = 1;
    89: op1_05_inv03 = 1;
    90: op1_05_inv03 = 1;
    92: op1_05_inv03 = 1;
    93: op1_05_inv03 = 1;
    96: op1_05_inv03 = 1;
    default: op1_05_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in04 = imem00_in[107:104];
    5: op1_05_in04 = reg_0036;
    6: op1_05_in04 = imem02_in[111:108];
    7: op1_05_in04 = reg_0264;
    8: op1_05_in04 = reg_0696;
    9: op1_05_in04 = reg_0621;
    10: op1_05_in04 = imem00_in[123:120];
    11: op1_05_in04 = reg_0433;
    3: op1_05_in04 = reg_0429;
    12: op1_05_in04 = reg_0096;
    13: op1_05_in04 = reg_0789;
    14: op1_05_in04 = imem07_in[79:76];
    15: op1_05_in04 = imem02_in[7:4];
    16: op1_05_in04 = reg_0389;
    17: op1_05_in04 = reg_0687;
    18: op1_05_in04 = imem04_in[119:116];
    2: op1_05_in04 = imem07_in[75:72];
    19: op1_05_in04 = reg_0691;
    20: op1_05_in04 = imem04_in[71:68];
    21: op1_05_in04 = imem00_in[111:108];
    22: op1_05_in04 = imem00_in[47:44];
    23: op1_05_in04 = reg_0606;
    24: op1_05_in04 = imem02_in[51:48];
    25: op1_05_in04 = imem04_in[83:80];
    26: op1_05_in04 = imem02_in[71:68];
    27: op1_05_in04 = reg_0270;
    28: op1_05_in04 = reg_0695;
    83: op1_05_in04 = reg_0695;
    29: op1_05_in04 = reg_0690;
    30: op1_05_in04 = reg_0562;
    31: op1_05_in04 = reg_0617;
    32: op1_05_in04 = imem00_in[51:48];
    33: op1_05_in04 = reg_0647;
    34: op1_05_in04 = reg_0161;
    35: op1_05_in04 = imem06_in[91:88];
    36: op1_05_in04 = reg_0436;
    37: op1_05_in04 = reg_0168;
    38: op1_05_in04 = reg_0676;
    39: op1_05_in04 = imem02_in[127:124];
    40: op1_05_in04 = reg_0672;
    41: op1_05_in04 = imem05_in[127:124];
    42: op1_05_in04 = reg_0708;
    43: op1_05_in04 = imem00_in[71:68];
    44: op1_05_in04 = reg_0387;
    45: op1_05_in04 = reg_0780;
    46: op1_05_in04 = imem00_in[119:116];
    59: op1_05_in04 = imem00_in[119:116];
    47: op1_05_in04 = reg_0116;
    48: op1_05_in04 = reg_0131;
    49: op1_05_in04 = reg_0555;
    50: op1_05_in04 = reg_0578;
    51: op1_05_in04 = reg_0683;
    52: op1_05_in04 = reg_0655;
    53: op1_05_in04 = reg_0499;
    54: op1_05_in04 = reg_0430;
    55: op1_05_in04 = reg_0520;
    56: op1_05_in04 = imem06_in[59:56];
    57: op1_05_in04 = reg_0053;
    58: op1_05_in04 = reg_0256;
    60: op1_05_in04 = reg_0448;
    61: op1_05_in04 = reg_0698;
    62: op1_05_in04 = reg_0564;
    63: op1_05_in04 = reg_0059;
    64: op1_05_in04 = reg_0086;
    65: op1_05_in04 = reg_0154;
    66: op1_05_in04 = reg_0774;
    67: op1_05_in04 = reg_0580;
    80: op1_05_in04 = reg_0580;
    68: op1_05_in04 = reg_0121;
    69: op1_05_in04 = imem04_in[55:52];
    70: op1_05_in04 = imem06_in[55:52];
    71: op1_05_in04 = reg_0809;
    72: op1_05_in04 = reg_0062;
    73: op1_05_in04 = imem06_in[11:8];
    74: op1_05_in04 = reg_0100;
    75: op1_05_in04 = reg_0492;
    89: op1_05_in04 = reg_0492;
    76: op1_05_in04 = reg_0749;
    77: op1_05_in04 = reg_0601;
    78: op1_05_in04 = reg_0547;
    79: op1_05_in04 = reg_0152;
    81: op1_05_in04 = imem06_in[31:28];
    82: op1_05_in04 = reg_0705;
    84: op1_05_in04 = imem05_in[27:24];
    85: op1_05_in04 = reg_0064;
    86: op1_05_in04 = reg_0281;
    87: op1_05_in04 = reg_0262;
    88: op1_05_in04 = reg_0658;
    90: op1_05_in04 = reg_0153;
    91: op1_05_in04 = reg_0734;
    92: op1_05_in04 = imem00_in[43:40];
    93: op1_05_in04 = reg_0688;
    94: op1_05_in04 = imem00_in[83:80];
    95: op1_05_in04 = reg_0699;
    96: op1_05_in04 = reg_0784;
    default: op1_05_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv04 = 1;
    7: op1_05_inv04 = 1;
    8: op1_05_inv04 = 1;
    9: op1_05_inv04 = 1;
    12: op1_05_inv04 = 1;
    14: op1_05_inv04 = 1;
    17: op1_05_inv04 = 1;
    18: op1_05_inv04 = 1;
    19: op1_05_inv04 = 1;
    20: op1_05_inv04 = 1;
    24: op1_05_inv04 = 1;
    25: op1_05_inv04 = 1;
    26: op1_05_inv04 = 1;
    30: op1_05_inv04 = 1;
    31: op1_05_inv04 = 1;
    33: op1_05_inv04 = 1;
    37: op1_05_inv04 = 1;
    38: op1_05_inv04 = 1;
    40: op1_05_inv04 = 1;
    41: op1_05_inv04 = 1;
    42: op1_05_inv04 = 1;
    43: op1_05_inv04 = 1;
    46: op1_05_inv04 = 1;
    47: op1_05_inv04 = 1;
    51: op1_05_inv04 = 1;
    52: op1_05_inv04 = 1;
    54: op1_05_inv04 = 1;
    58: op1_05_inv04 = 1;
    60: op1_05_inv04 = 1;
    61: op1_05_inv04 = 1;
    62: op1_05_inv04 = 1;
    63: op1_05_inv04 = 1;
    64: op1_05_inv04 = 1;
    67: op1_05_inv04 = 1;
    69: op1_05_inv04 = 1;
    77: op1_05_inv04 = 1;
    78: op1_05_inv04 = 1;
    81: op1_05_inv04 = 1;
    84: op1_05_inv04 = 1;
    87: op1_05_inv04 = 1;
    88: op1_05_inv04 = 1;
    91: op1_05_inv04 = 1;
    92: op1_05_inv04 = 1;
    94: op1_05_inv04 = 1;
    95: op1_05_inv04 = 1;
    96: op1_05_inv04 = 1;
    default: op1_05_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in05 = imem00_in[115:112];
    21: op1_05_in05 = imem00_in[115:112];
    94: op1_05_in05 = imem00_in[115:112];
    5: op1_05_in05 = reg_0021;
    6: op1_05_in05 = imem02_in[115:112];
    7: op1_05_in05 = reg_0229;
    8: op1_05_in05 = reg_0689;
    61: op1_05_in05 = reg_0689;
    9: op1_05_in05 = reg_0616;
    31: op1_05_in05 = reg_0616;
    10: op1_05_in05 = reg_0675;
    11: op1_05_in05 = reg_0426;
    3: op1_05_in05 = reg_0436;
    12: op1_05_in05 = reg_0090;
    13: op1_05_in05 = reg_0491;
    14: op1_05_in05 = imem07_in[87:84];
    15: op1_05_in05 = imem02_in[35:32];
    16: op1_05_in05 = reg_0000;
    17: op1_05_in05 = reg_0699;
    18: op1_05_in05 = reg_0078;
    2: op1_05_in05 = imem07_in[127:124];
    19: op1_05_in05 = reg_0688;
    20: op1_05_in05 = imem04_in[127:124];
    22: op1_05_in05 = imem00_in[55:52];
    23: op1_05_in05 = reg_0609;
    24: op1_05_in05 = imem02_in[55:52];
    25: op1_05_in05 = imem04_in[99:96];
    26: op1_05_in05 = imem02_in[103:100];
    27: op1_05_in05 = reg_0331;
    28: op1_05_in05 = reg_0682;
    29: op1_05_in05 = reg_0454;
    30: op1_05_in05 = reg_0376;
    32: op1_05_in05 = imem00_in[83:80];
    33: op1_05_in05 = reg_0636;
    34: op1_05_in05 = reg_0183;
    35: op1_05_in05 = imem06_in[95:92];
    36: op1_05_in05 = reg_0422;
    37: op1_05_in05 = reg_0157;
    38: op1_05_in05 = reg_0686;
    39: op1_05_in05 = reg_0653;
    40: op1_05_in05 = reg_0694;
    41: op1_05_in05 = reg_0798;
    42: op1_05_in05 = reg_0715;
    43: op1_05_in05 = imem00_in[99:96];
    44: op1_05_in05 = reg_0564;
    45: op1_05_in05 = reg_0785;
    46: op1_05_in05 = reg_0693;
    47: op1_05_in05 = reg_0117;
    48: op1_05_in05 = imem06_in[11:8];
    49: op1_05_in05 = reg_0060;
    50: op1_05_in05 = reg_0394;
    51: op1_05_in05 = reg_0469;
    52: op1_05_in05 = reg_0661;
    53: op1_05_in05 = reg_0396;
    54: op1_05_in05 = reg_0503;
    55: op1_05_in05 = reg_0296;
    56: op1_05_in05 = imem06_in[71:68];
    57: op1_05_in05 = reg_0449;
    58: op1_05_in05 = reg_0102;
    59: op1_05_in05 = reg_0612;
    60: op1_05_in05 = reg_0435;
    62: op1_05_in05 = reg_0562;
    63: op1_05_in05 = reg_0537;
    64: op1_05_in05 = reg_0150;
    65: op1_05_in05 = reg_0155;
    66: op1_05_in05 = reg_0644;
    67: op1_05_in05 = reg_0035;
    68: op1_05_in05 = imem02_in[75:72];
    69: op1_05_in05 = imem04_in[119:116];
    70: op1_05_in05 = imem06_in[83:80];
    71: op1_05_in05 = reg_0004;
    72: op1_05_in05 = reg_0771;
    73: op1_05_in05 = imem06_in[43:40];
    74: op1_05_in05 = reg_0709;
    75: op1_05_in05 = reg_0690;
    76: op1_05_in05 = reg_0494;
    77: op1_05_in05 = reg_0674;
    78: op1_05_in05 = reg_0077;
    79: op1_05_in05 = reg_0783;
    80: op1_05_in05 = reg_0777;
    81: op1_05_in05 = imem06_in[103:100];
    82: op1_05_in05 = reg_0362;
    83: op1_05_in05 = reg_0492;
    84: op1_05_in05 = imem05_in[35:32];
    85: op1_05_in05 = reg_0053;
    86: op1_05_in05 = reg_0136;
    87: op1_05_in05 = reg_0553;
    88: op1_05_in05 = reg_0691;
    89: op1_05_in05 = reg_0285;
    90: op1_05_in05 = reg_0828;
    91: op1_05_in05 = imem06_in[3:0];
    92: op1_05_in05 = imem00_in[71:68];
    93: op1_05_in05 = reg_0455;
    95: op1_05_in05 = reg_0465;
    96: op1_05_in05 = reg_0382;
    default: op1_05_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv05 = 1;
    9: op1_05_inv05 = 1;
    11: op1_05_inv05 = 1;
    3: op1_05_inv05 = 1;
    12: op1_05_inv05 = 1;
    13: op1_05_inv05 = 1;
    14: op1_05_inv05 = 1;
    15: op1_05_inv05 = 1;
    16: op1_05_inv05 = 1;
    2: op1_05_inv05 = 1;
    19: op1_05_inv05 = 1;
    23: op1_05_inv05 = 1;
    24: op1_05_inv05 = 1;
    27: op1_05_inv05 = 1;
    29: op1_05_inv05 = 1;
    33: op1_05_inv05 = 1;
    34: op1_05_inv05 = 1;
    35: op1_05_inv05 = 1;
    40: op1_05_inv05 = 1;
    42: op1_05_inv05 = 1;
    43: op1_05_inv05 = 1;
    49: op1_05_inv05 = 1;
    50: op1_05_inv05 = 1;
    52: op1_05_inv05 = 1;
    55: op1_05_inv05 = 1;
    58: op1_05_inv05 = 1;
    63: op1_05_inv05 = 1;
    64: op1_05_inv05 = 1;
    69: op1_05_inv05 = 1;
    71: op1_05_inv05 = 1;
    72: op1_05_inv05 = 1;
    74: op1_05_inv05 = 1;
    79: op1_05_inv05 = 1;
    80: op1_05_inv05 = 1;
    81: op1_05_inv05 = 1;
    87: op1_05_inv05 = 1;
    88: op1_05_inv05 = 1;
    89: op1_05_inv05 = 1;
    94: op1_05_inv05 = 1;
    default: op1_05_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in06 = reg_0674;
    5: op1_05_in06 = reg_0029;
    6: op1_05_in06 = imem02_in[119:116];
    7: op1_05_in06 = reg_0260;
    8: op1_05_in06 = reg_0671;
    9: op1_05_in06 = reg_0626;
    10: op1_05_in06 = reg_0687;
    11: op1_05_in06 = reg_0447;
    3: op1_05_in06 = reg_0447;
    12: op1_05_in06 = reg_0051;
    13: op1_05_in06 = reg_0785;
    41: op1_05_in06 = reg_0785;
    14: op1_05_in06 = imem07_in[95:92];
    15: op1_05_in06 = imem02_in[43:40];
    16: op1_05_in06 = reg_0001;
    17: op1_05_in06 = reg_0463;
    18: op1_05_in06 = reg_0067;
    2: op1_05_in06 = reg_0180;
    19: op1_05_in06 = reg_0673;
    20: op1_05_in06 = reg_0545;
    21: op1_05_in06 = reg_0682;
    22: op1_05_in06 = imem00_in[63:60];
    23: op1_05_in06 = reg_0632;
    24: op1_05_in06 = imem02_in[67:64];
    25: op1_05_in06 = imem04_in[103:100];
    26: op1_05_in06 = reg_0658;
    27: op1_05_in06 = reg_0582;
    28: op1_05_in06 = reg_0698;
    59: op1_05_in06 = reg_0698;
    29: op1_05_in06 = reg_0450;
    30: op1_05_in06 = reg_0396;
    31: op1_05_in06 = reg_0631;
    32: op1_05_in06 = imem00_in[87:84];
    33: op1_05_in06 = reg_0667;
    34: op1_05_in06 = reg_0171;
    35: op1_05_in06 = imem06_in[99:96];
    36: op1_05_in06 = reg_0433;
    38: op1_05_in06 = reg_0670;
    39: op1_05_in06 = reg_0654;
    40: op1_05_in06 = reg_0668;
    42: op1_05_in06 = reg_0701;
    43: op1_05_in06 = imem00_in[119:116];
    44: op1_05_in06 = reg_0517;
    45: op1_05_in06 = reg_0786;
    46: op1_05_in06 = reg_0681;
    47: op1_05_in06 = reg_0126;
    48: op1_05_in06 = imem06_in[55:52];
    73: op1_05_in06 = imem06_in[55:52];
    49: op1_05_in06 = reg_0556;
    50: op1_05_in06 = reg_0575;
    51: op1_05_in06 = reg_0473;
    52: op1_05_in06 = reg_0647;
    53: op1_05_in06 = reg_0374;
    54: op1_05_in06 = reg_0062;
    55: op1_05_in06 = reg_0115;
    56: op1_05_in06 = imem06_in[87:84];
    57: op1_05_in06 = reg_0440;
    58: op1_05_in06 = reg_0226;
    60: op1_05_in06 = reg_0174;
    61: op1_05_in06 = reg_0407;
    62: op1_05_in06 = reg_0393;
    63: op1_05_in06 = reg_0555;
    64: op1_05_in06 = reg_0146;
    65: op1_05_in06 = reg_0144;
    66: op1_05_in06 = imem05_in[19:16];
    67: op1_05_in06 = reg_0534;
    87: op1_05_in06 = reg_0534;
    68: op1_05_in06 = imem02_in[107:104];
    69: op1_05_in06 = reg_0262;
    70: op1_05_in06 = imem06_in[103:100];
    71: op1_05_in06 = imem04_in[7:4];
    72: op1_05_in06 = reg_0136;
    74: op1_05_in06 = reg_0711;
    75: op1_05_in06 = reg_0691;
    76: op1_05_in06 = reg_0247;
    77: op1_05_in06 = reg_0121;
    78: op1_05_in06 = reg_0071;
    79: op1_05_in06 = imem06_in[19:16];
    80: op1_05_in06 = reg_0011;
    81: op1_05_in06 = imem06_in[107:104];
    82: op1_05_in06 = reg_0356;
    83: op1_05_in06 = reg_0694;
    84: op1_05_in06 = imem05_in[79:76];
    85: op1_05_in06 = reg_0239;
    86: op1_05_in06 = reg_0094;
    88: op1_05_in06 = reg_0480;
    89: op1_05_in06 = reg_0822;
    90: op1_05_in06 = reg_0824;
    91: op1_05_in06 = imem06_in[71:68];
    92: op1_05_in06 = imem00_in[83:80];
    93: op1_05_in06 = reg_0464;
    94: op1_05_in06 = imem00_in[127:124];
    95: op1_05_in06 = reg_0469;
    96: op1_05_in06 = reg_0166;
    default: op1_05_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv06 = 1;
    5: op1_05_inv06 = 1;
    6: op1_05_inv06 = 1;
    8: op1_05_inv06 = 1;
    10: op1_05_inv06 = 1;
    3: op1_05_inv06 = 1;
    12: op1_05_inv06 = 1;
    15: op1_05_inv06 = 1;
    17: op1_05_inv06 = 1;
    19: op1_05_inv06 = 1;
    20: op1_05_inv06 = 1;
    24: op1_05_inv06 = 1;
    26: op1_05_inv06 = 1;
    30: op1_05_inv06 = 1;
    31: op1_05_inv06 = 1;
    32: op1_05_inv06 = 1;
    33: op1_05_inv06 = 1;
    34: op1_05_inv06 = 1;
    38: op1_05_inv06 = 1;
    42: op1_05_inv06 = 1;
    44: op1_05_inv06 = 1;
    46: op1_05_inv06 = 1;
    50: op1_05_inv06 = 1;
    53: op1_05_inv06 = 1;
    55: op1_05_inv06 = 1;
    57: op1_05_inv06 = 1;
    59: op1_05_inv06 = 1;
    61: op1_05_inv06 = 1;
    62: op1_05_inv06 = 1;
    63: op1_05_inv06 = 1;
    65: op1_05_inv06 = 1;
    68: op1_05_inv06 = 1;
    70: op1_05_inv06 = 1;
    74: op1_05_inv06 = 1;
    76: op1_05_inv06 = 1;
    80: op1_05_inv06 = 1;
    87: op1_05_inv06 = 1;
    89: op1_05_inv06 = 1;
    91: op1_05_inv06 = 1;
    92: op1_05_inv06 = 1;
    94: op1_05_inv06 = 1;
    95: op1_05_inv06 = 1;
    default: op1_05_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in07 = reg_0475;
    5: op1_05_in07 = reg_0022;
    6: op1_05_in07 = reg_0357;
    7: op1_05_in07 = reg_0265;
    8: op1_05_in07 = reg_0680;
    75: op1_05_in07 = reg_0680;
    9: op1_05_in07 = reg_0615;
    10: op1_05_in07 = reg_0692;
    76: op1_05_in07 = reg_0692;
    11: op1_05_in07 = reg_0419;
    3: op1_05_in07 = reg_0418;
    12: op1_05_in07 = reg_0094;
    13: op1_05_in07 = reg_0782;
    14: op1_05_in07 = imem07_in[107:104];
    15: op1_05_in07 = imem02_in[51:48];
    16: op1_05_in07 = reg_0002;
    17: op1_05_in07 = reg_0464;
    18: op1_05_in07 = reg_0289;
    2: op1_05_in07 = reg_0172;
    19: op1_05_in07 = reg_0687;
    20: op1_05_in07 = reg_0557;
    21: op1_05_in07 = reg_0683;
    22: op1_05_in07 = imem00_in[67:64];
    23: op1_05_in07 = reg_0402;
    24: op1_05_in07 = imem02_in[87:84];
    25: op1_05_in07 = imem04_in[111:108];
    26: op1_05_in07 = reg_0660;
    27: op1_05_in07 = reg_0593;
    28: op1_05_in07 = reg_0679;
    29: op1_05_in07 = reg_0455;
    30: op1_05_in07 = reg_0001;
    31: op1_05_in07 = reg_0331;
    32: op1_05_in07 = imem00_in[91:88];
    33: op1_05_in07 = reg_0663;
    35: op1_05_in07 = imem06_in[115:112];
    36: op1_05_in07 = reg_0421;
    38: op1_05_in07 = reg_0690;
    39: op1_05_in07 = reg_0639;
    40: op1_05_in07 = reg_0465;
    41: op1_05_in07 = reg_0794;
    42: op1_05_in07 = imem07_in[3:0];
    70: op1_05_in07 = imem07_in[3:0];
    74: op1_05_in07 = imem07_in[3:0];
    43: op1_05_in07 = imem00_in[123:120];
    44: op1_05_in07 = reg_0572;
    45: op1_05_in07 = reg_0736;
    46: op1_05_in07 = reg_0672;
    47: op1_05_in07 = imem02_in[55:52];
    48: op1_05_in07 = imem06_in[87:84];
    49: op1_05_in07 = reg_0429;
    50: op1_05_in07 = reg_0499;
    51: op1_05_in07 = reg_0474;
    52: op1_05_in07 = reg_0659;
    53: op1_05_in07 = reg_0389;
    54: op1_05_in07 = reg_0068;
    55: op1_05_in07 = reg_0491;
    56: op1_05_in07 = reg_0408;
    57: op1_05_in07 = reg_0180;
    58: op1_05_in07 = reg_0279;
    59: op1_05_in07 = reg_0689;
    60: op1_05_in07 = reg_0175;
    61: op1_05_in07 = reg_0494;
    62: op1_05_in07 = reg_0747;
    63: op1_05_in07 = reg_0060;
    64: op1_05_in07 = reg_0139;
    65: op1_05_in07 = imem06_in[15:12];
    66: op1_05_in07 = imem05_in[59:56];
    67: op1_05_in07 = reg_0777;
    68: op1_05_in07 = reg_0785;
    69: op1_05_in07 = reg_0552;
    71: op1_05_in07 = imem04_in[63:60];
    72: op1_05_in07 = reg_0781;
    73: op1_05_in07 = imem06_in[103:100];
    77: op1_05_in07 = reg_0678;
    78: op1_05_in07 = reg_0078;
    79: op1_05_in07 = imem06_in[23:20];
    80: op1_05_in07 = reg_0256;
    81: op1_05_in07 = imem06_in[111:108];
    82: op1_05_in07 = reg_0360;
    83: op1_05_in07 = reg_0612;
    84: op1_05_in07 = imem05_in[91:88];
    85: op1_05_in07 = reg_0449;
    86: op1_05_in07 = reg_0532;
    87: op1_05_in07 = reg_0179;
    88: op1_05_in07 = reg_0467;
    89: op1_05_in07 = reg_0742;
    90: op1_05_in07 = imem06_in[31:28];
    91: op1_05_in07 = reg_0349;
    92: op1_05_in07 = imem00_in[115:112];
    93: op1_05_in07 = reg_0462;
    94: op1_05_in07 = reg_0695;
    95: op1_05_in07 = reg_0466;
    96: op1_05_in07 = reg_0708;
    default: op1_05_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv07 = 1;
    6: op1_05_inv07 = 1;
    8: op1_05_inv07 = 1;
    10: op1_05_inv07 = 1;
    11: op1_05_inv07 = 1;
    13: op1_05_inv07 = 1;
    17: op1_05_inv07 = 1;
    18: op1_05_inv07 = 1;
    20: op1_05_inv07 = 1;
    23: op1_05_inv07 = 1;
    27: op1_05_inv07 = 1;
    28: op1_05_inv07 = 1;
    31: op1_05_inv07 = 1;
    36: op1_05_inv07 = 1;
    39: op1_05_inv07 = 1;
    40: op1_05_inv07 = 1;
    43: op1_05_inv07 = 1;
    44: op1_05_inv07 = 1;
    47: op1_05_inv07 = 1;
    50: op1_05_inv07 = 1;
    51: op1_05_inv07 = 1;
    53: op1_05_inv07 = 1;
    55: op1_05_inv07 = 1;
    56: op1_05_inv07 = 1;
    58: op1_05_inv07 = 1;
    59: op1_05_inv07 = 1;
    64: op1_05_inv07 = 1;
    66: op1_05_inv07 = 1;
    67: op1_05_inv07 = 1;
    70: op1_05_inv07 = 1;
    71: op1_05_inv07 = 1;
    73: op1_05_inv07 = 1;
    80: op1_05_inv07 = 1;
    81: op1_05_inv07 = 1;
    83: op1_05_inv07 = 1;
    84: op1_05_inv07 = 1;
    86: op1_05_inv07 = 1;
    87: op1_05_inv07 = 1;
    93: op1_05_inv07 = 1;
    94: op1_05_inv07 = 1;
    default: op1_05_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in08 = reg_0452;
    5: op1_05_in08 = imem07_in[11:8];
    6: op1_05_in08 = reg_0330;
    7: op1_05_in08 = reg_0255;
    18: op1_05_in08 = reg_0255;
    8: op1_05_in08 = reg_0669;
    19: op1_05_in08 = reg_0669;
    9: op1_05_in08 = reg_0332;
    10: op1_05_in08 = reg_0463;
    11: op1_05_in08 = reg_0444;
    3: op1_05_in08 = reg_0437;
    12: op1_05_in08 = imem03_in[27:24];
    13: op1_05_in08 = reg_0485;
    14: op1_05_in08 = reg_0728;
    15: op1_05_in08 = reg_0650;
    16: op1_05_in08 = reg_0003;
    17: op1_05_in08 = reg_0466;
    2: op1_05_in08 = reg_0165;
    60: op1_05_in08 = reg_0165;
    20: op1_05_in08 = reg_0548;
    21: op1_05_in08 = reg_0676;
    43: op1_05_in08 = reg_0676;
    46: op1_05_in08 = reg_0676;
    22: op1_05_in08 = imem00_in[87:84];
    23: op1_05_in08 = reg_0372;
    24: op1_05_in08 = reg_0665;
    25: op1_05_in08 = reg_0262;
    26: op1_05_in08 = reg_0639;
    27: op1_05_in08 = reg_0576;
    28: op1_05_in08 = reg_0691;
    59: op1_05_in08 = reg_0691;
    29: op1_05_in08 = reg_0461;
    40: op1_05_in08 = reg_0461;
    30: op1_05_in08 = reg_0002;
    31: op1_05_in08 = reg_0270;
    32: op1_05_in08 = imem00_in[111:108];
    33: op1_05_in08 = reg_0349;
    35: op1_05_in08 = reg_0775;
    56: op1_05_in08 = reg_0775;
    36: op1_05_in08 = reg_0419;
    38: op1_05_in08 = reg_0677;
    39: op1_05_in08 = reg_0648;
    41: op1_05_in08 = reg_0786;
    42: op1_05_in08 = imem07_in[51:48];
    44: op1_05_in08 = reg_0396;
    45: op1_05_in08 = reg_0085;
    47: op1_05_in08 = imem02_in[71:68];
    48: op1_05_in08 = imem06_in[103:100];
    49: op1_05_in08 = reg_0079;
    50: op1_05_in08 = reg_0747;
    51: op1_05_in08 = reg_0187;
    52: op1_05_in08 = reg_0352;
    53: op1_05_in08 = reg_0570;
    54: op1_05_in08 = reg_0275;
    55: op1_05_in08 = reg_0260;
    57: op1_05_in08 = reg_0185;
    58: op1_05_in08 = reg_0257;
    89: op1_05_in08 = reg_0257;
    61: op1_05_in08 = reg_0699;
    62: op1_05_in08 = reg_0389;
    63: op1_05_in08 = reg_0516;
    64: op1_05_in08 = reg_0137;
    65: op1_05_in08 = imem06_in[31:28];
    79: op1_05_in08 = imem06_in[31:28];
    66: op1_05_in08 = imem05_in[87:84];
    67: op1_05_in08 = reg_0368;
    68: op1_05_in08 = reg_0657;
    69: op1_05_in08 = reg_0554;
    70: op1_05_in08 = imem07_in[15:12];
    71: op1_05_in08 = imem04_in[75:72];
    72: op1_05_in08 = reg_0391;
    73: op1_05_in08 = imem06_in[127:124];
    74: op1_05_in08 = imem07_in[63:60];
    75: op1_05_in08 = reg_0688;
    76: op1_05_in08 = reg_0453;
    77: op1_05_in08 = imem02_in[15:12];
    78: op1_05_in08 = reg_0296;
    80: op1_05_in08 = reg_0057;
    81: op1_05_in08 = imem06_in[119:116];
    82: op1_05_in08 = reg_0590;
    83: op1_05_in08 = reg_0686;
    84: op1_05_in08 = reg_0337;
    85: op1_05_in08 = reg_0438;
    86: op1_05_in08 = imem03_in[15:12];
    87: op1_05_in08 = reg_0536;
    88: op1_05_in08 = reg_0456;
    90: op1_05_in08 = imem06_in[35:32];
    91: op1_05_in08 = reg_0409;
    92: op1_05_in08 = reg_0000;
    93: op1_05_in08 = reg_0474;
    94: op1_05_in08 = reg_0744;
    95: op1_05_in08 = reg_0473;
    96: op1_05_in08 = reg_0158;
    default: op1_05_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv08 = 1;
    6: op1_05_inv08 = 1;
    8: op1_05_inv08 = 1;
    9: op1_05_inv08 = 1;
    10: op1_05_inv08 = 1;
    11: op1_05_inv08 = 1;
    3: op1_05_inv08 = 1;
    12: op1_05_inv08 = 1;
    20: op1_05_inv08 = 1;
    22: op1_05_inv08 = 1;
    24: op1_05_inv08 = 1;
    28: op1_05_inv08 = 1;
    38: op1_05_inv08 = 1;
    39: op1_05_inv08 = 1;
    46: op1_05_inv08 = 1;
    49: op1_05_inv08 = 1;
    54: op1_05_inv08 = 1;
    55: op1_05_inv08 = 1;
    56: op1_05_inv08 = 1;
    57: op1_05_inv08 = 1;
    58: op1_05_inv08 = 1;
    59: op1_05_inv08 = 1;
    62: op1_05_inv08 = 1;
    66: op1_05_inv08 = 1;
    67: op1_05_inv08 = 1;
    71: op1_05_inv08 = 1;
    72: op1_05_inv08 = 1;
    73: op1_05_inv08 = 1;
    76: op1_05_inv08 = 1;
    84: op1_05_inv08 = 1;
    85: op1_05_inv08 = 1;
    86: op1_05_inv08 = 1;
    89: op1_05_inv08 = 1;
    91: op1_05_inv08 = 1;
    93: op1_05_inv08 = 1;
    96: op1_05_inv08 = 1;
    default: op1_05_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in09 = reg_0208;
    5: op1_05_in09 = imem07_in[15:12];
    6: op1_05_in09 = reg_0310;
    7: op1_05_in09 = reg_0145;
    8: op1_05_in09 = reg_0454;
    9: op1_05_in09 = reg_0381;
    10: op1_05_in09 = reg_0460;
    29: op1_05_in09 = reg_0460;
    11: op1_05_in09 = reg_0437;
    3: op1_05_in09 = reg_0175;
    12: op1_05_in09 = imem03_in[51:48];
    13: op1_05_in09 = reg_0267;
    14: op1_05_in09 = reg_0719;
    15: op1_05_in09 = reg_0656;
    16: op1_05_in09 = reg_0801;
    17: op1_05_in09 = reg_0473;
    18: op1_05_in09 = reg_0068;
    2: op1_05_in09 = reg_0162;
    19: op1_05_in09 = reg_0475;
    20: op1_05_in09 = reg_0554;
    21: op1_05_in09 = reg_0687;
    22: op1_05_in09 = imem00_in[91:88];
    23: op1_05_in09 = reg_0033;
    24: op1_05_in09 = reg_0663;
    25: op1_05_in09 = reg_0544;
    26: op1_05_in09 = reg_0638;
    27: op1_05_in09 = imem03_in[19:16];
    28: op1_05_in09 = reg_0674;
    30: op1_05_in09 = reg_0807;
    31: op1_05_in09 = reg_0776;
    32: op1_05_in09 = imem00_in[123:120];
    33: op1_05_in09 = reg_0357;
    35: op1_05_in09 = reg_0773;
    36: op1_05_in09 = reg_0439;
    38: op1_05_in09 = reg_0691;
    39: op1_05_in09 = reg_0641;
    40: op1_05_in09 = reg_0477;
    41: op1_05_in09 = reg_0787;
    67: op1_05_in09 = reg_0787;
    42: op1_05_in09 = imem07_in[75:72];
    43: op1_05_in09 = reg_0684;
    44: op1_05_in09 = reg_0389;
    45: op1_05_in09 = reg_0224;
    46: op1_05_in09 = reg_0686;
    47: op1_05_in09 = imem02_in[95:92];
    48: op1_05_in09 = imem06_in[115:112];
    90: op1_05_in09 = imem06_in[115:112];
    49: op1_05_in09 = reg_0052;
    50: op1_05_in09 = reg_0396;
    51: op1_05_in09 = reg_0209;
    52: op1_05_in09 = reg_0341;
    53: op1_05_in09 = reg_0019;
    54: op1_05_in09 = imem05_in[23:20];
    55: op1_05_in09 = reg_0265;
    56: op1_05_in09 = reg_0748;
    57: op1_05_in09 = reg_0170;
    58: op1_05_in09 = reg_0086;
    59: op1_05_in09 = reg_0407;
    60: op1_05_in09 = reg_0161;
    61: op1_05_in09 = reg_0464;
    62: op1_05_in09 = reg_0811;
    63: op1_05_in09 = reg_0283;
    64: op1_05_in09 = imem06_in[11:8];
    65: op1_05_in09 = imem06_in[35:32];
    79: op1_05_in09 = imem06_in[35:32];
    66: op1_05_in09 = imem05_in[111:108];
    68: op1_05_in09 = reg_0417;
    69: op1_05_in09 = reg_0058;
    70: op1_05_in09 = imem07_in[39:36];
    71: op1_05_in09 = imem04_in[103:100];
    72: op1_05_in09 = reg_0393;
    73: op1_05_in09 = reg_0348;
    74: op1_05_in09 = imem07_in[91:88];
    75: op1_05_in09 = reg_0457;
    76: op1_05_in09 = reg_0469;
    77: op1_05_in09 = imem02_in[35:32];
    78: op1_05_in09 = reg_0136;
    80: op1_05_in09 = reg_0165;
    81: op1_05_in09 = reg_0289;
    82: op1_05_in09 = reg_0566;
    83: op1_05_in09 = reg_0255;
    84: op1_05_in09 = reg_0070;
    92: op1_05_in09 = reg_0070;
    85: op1_05_in09 = reg_0141;
    86: op1_05_in09 = imem03_in[59:56];
    87: op1_05_in09 = reg_0510;
    88: op1_05_in09 = reg_0214;
    89: op1_05_in09 = reg_0765;
    91: op1_05_in09 = reg_0038;
    93: op1_05_in09 = reg_0479;
    94: op1_05_in09 = reg_0131;
    95: op1_05_in09 = reg_0467;
    96: op1_05_in09 = reg_0731;
    default: op1_05_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv09 = 1;
    10: op1_05_inv09 = 1;
    3: op1_05_inv09 = 1;
    13: op1_05_inv09 = 1;
    16: op1_05_inv09 = 1;
    17: op1_05_inv09 = 1;
    2: op1_05_inv09 = 1;
    20: op1_05_inv09 = 1;
    21: op1_05_inv09 = 1;
    22: op1_05_inv09 = 1;
    23: op1_05_inv09 = 1;
    24: op1_05_inv09 = 1;
    25: op1_05_inv09 = 1;
    26: op1_05_inv09 = 1;
    27: op1_05_inv09 = 1;
    32: op1_05_inv09 = 1;
    35: op1_05_inv09 = 1;
    40: op1_05_inv09 = 1;
    45: op1_05_inv09 = 1;
    47: op1_05_inv09 = 1;
    48: op1_05_inv09 = 1;
    52: op1_05_inv09 = 1;
    55: op1_05_inv09 = 1;
    57: op1_05_inv09 = 1;
    58: op1_05_inv09 = 1;
    59: op1_05_inv09 = 1;
    60: op1_05_inv09 = 1;
    61: op1_05_inv09 = 1;
    63: op1_05_inv09 = 1;
    66: op1_05_inv09 = 1;
    67: op1_05_inv09 = 1;
    69: op1_05_inv09 = 1;
    71: op1_05_inv09 = 1;
    73: op1_05_inv09 = 1;
    74: op1_05_inv09 = 1;
    77: op1_05_inv09 = 1;
    78: op1_05_inv09 = 1;
    80: op1_05_inv09 = 1;
    81: op1_05_inv09 = 1;
    82: op1_05_inv09 = 1;
    84: op1_05_inv09 = 1;
    85: op1_05_inv09 = 1;
    89: op1_05_inv09 = 1;
    91: op1_05_inv09 = 1;
    93: op1_05_inv09 = 1;
    96: op1_05_inv09 = 1;
    default: op1_05_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in10 = reg_0191;
    5: op1_05_in10 = imem07_in[71:68];
    6: op1_05_in10 = reg_0083;
    7: op1_05_in10 = reg_0136;
    8: op1_05_in10 = reg_0466;
    9: op1_05_in10 = reg_0392;
    10: op1_05_in10 = reg_0480;
    11: op1_05_in10 = reg_0448;
    3: op1_05_in10 = reg_0162;
    12: op1_05_in10 = imem03_in[63:60];
    13: op1_05_in10 = reg_0736;
    41: op1_05_in10 = reg_0736;
    14: op1_05_in10 = reg_0726;
    15: op1_05_in10 = reg_0649;
    16: op1_05_in10 = imem04_in[7:4];
    17: op1_05_in10 = reg_0470;
    18: op1_05_in10 = imem05_in[15:12];
    2: op1_05_in10 = reg_0167;
    19: op1_05_in10 = reg_0468;
    20: op1_05_in10 = reg_0546;
    21: op1_05_in10 = reg_0669;
    22: op1_05_in10 = reg_0672;
    23: op1_05_in10 = reg_0040;
    24: op1_05_in10 = reg_0364;
    25: op1_05_in10 = reg_0553;
    26: op1_05_in10 = reg_0659;
    27: op1_05_in10 = imem03_in[39:36];
    28: op1_05_in10 = reg_0678;
    29: op1_05_in10 = reg_0462;
    83: op1_05_in10 = reg_0462;
    30: op1_05_in10 = reg_0804;
    31: op1_05_in10 = reg_0404;
    32: op1_05_in10 = reg_0694;
    33: op1_05_in10 = reg_0362;
    35: op1_05_in10 = reg_0748;
    36: op1_05_in10 = reg_0446;
    38: op1_05_in10 = reg_0671;
    39: op1_05_in10 = reg_0665;
    40: op1_05_in10 = reg_0469;
    42: op1_05_in10 = imem07_in[119:116];
    43: op1_05_in10 = reg_0670;
    46: op1_05_in10 = reg_0670;
    44: op1_05_in10 = reg_0012;
    45: op1_05_in10 = reg_0089;
    47: op1_05_in10 = reg_0651;
    48: op1_05_in10 = imem06_in[127:124];
    49: op1_05_in10 = reg_0074;
    50: op1_05_in10 = reg_0386;
    51: op1_05_in10 = reg_0186;
    52: op1_05_in10 = reg_0345;
    53: op1_05_in10 = reg_0811;
    54: op1_05_in10 = imem05_in[51:48];
    55: op1_05_in10 = reg_0787;
    56: op1_05_in10 = reg_0403;
    58: op1_05_in10 = reg_0146;
    59: op1_05_in10 = reg_0494;
    60: op1_05_in10 = reg_0183;
    61: op1_05_in10 = reg_0477;
    62: op1_05_in10 = reg_0803;
    63: op1_05_in10 = reg_0077;
    64: op1_05_in10 = imem06_in[23:20];
    65: op1_05_in10 = imem06_in[71:68];
    66: op1_05_in10 = reg_0337;
    67: op1_05_in10 = reg_0623;
    68: op1_05_in10 = reg_0655;
    69: op1_05_in10 = reg_0052;
    70: op1_05_in10 = imem07_in[59:56];
    71: op1_05_in10 = imem04_in[119:116];
    72: op1_05_in10 = imem05_in[23:20];
    73: op1_05_in10 = reg_0346;
    74: op1_05_in10 = imem07_in[115:112];
    75: op1_05_in10 = reg_0464;
    76: op1_05_in10 = reg_0452;
    77: op1_05_in10 = imem02_in[51:48];
    78: op1_05_in10 = reg_0099;
    79: op1_05_in10 = imem06_in[43:40];
    80: op1_05_in10 = reg_0066;
    81: op1_05_in10 = reg_0624;
    82: op1_05_in10 = reg_0514;
    84: op1_05_in10 = reg_0793;
    86: op1_05_in10 = imem03_in[75:72];
    87: op1_05_in10 = reg_0283;
    88: op1_05_in10 = reg_0189;
    89: op1_05_in10 = imem06_in[39:36];
    90: op1_05_in10 = imem06_in[123:120];
    91: op1_05_in10 = reg_0168;
    92: op1_05_in10 = reg_0461;
    93: op1_05_in10 = reg_0201;
    94: op1_05_in10 = reg_0463;
    95: op1_05_in10 = reg_0474;
    96: op1_05_in10 = reg_0334;
    default: op1_05_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv10 = 1;
    7: op1_05_inv10 = 1;
    9: op1_05_inv10 = 1;
    13: op1_05_inv10 = 1;
    17: op1_05_inv10 = 1;
    18: op1_05_inv10 = 1;
    20: op1_05_inv10 = 1;
    21: op1_05_inv10 = 1;
    22: op1_05_inv10 = 1;
    23: op1_05_inv10 = 1;
    24: op1_05_inv10 = 1;
    26: op1_05_inv10 = 1;
    29: op1_05_inv10 = 1;
    30: op1_05_inv10 = 1;
    35: op1_05_inv10 = 1;
    36: op1_05_inv10 = 1;
    39: op1_05_inv10 = 1;
    42: op1_05_inv10 = 1;
    45: op1_05_inv10 = 1;
    46: op1_05_inv10 = 1;
    48: op1_05_inv10 = 1;
    53: op1_05_inv10 = 1;
    54: op1_05_inv10 = 1;
    58: op1_05_inv10 = 1;
    59: op1_05_inv10 = 1;
    60: op1_05_inv10 = 1;
    61: op1_05_inv10 = 1;
    64: op1_05_inv10 = 1;
    65: op1_05_inv10 = 1;
    67: op1_05_inv10 = 1;
    68: op1_05_inv10 = 1;
    69: op1_05_inv10 = 1;
    70: op1_05_inv10 = 1;
    73: op1_05_inv10 = 1;
    76: op1_05_inv10 = 1;
    83: op1_05_inv10 = 1;
    86: op1_05_inv10 = 1;
    87: op1_05_inv10 = 1;
    88: op1_05_inv10 = 1;
    91: op1_05_inv10 = 1;
    92: op1_05_inv10 = 1;
    93: op1_05_inv10 = 1;
    94: op1_05_inv10 = 1;
    95: op1_05_inv10 = 1;
    default: op1_05_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in11 = reg_0209;
    5: op1_05_in11 = reg_0722;
    6: op1_05_in11 = reg_0042;
    7: op1_05_in11 = reg_0151;
    8: op1_05_in11 = reg_0471;
    9: op1_05_in11 = reg_0351;
    10: op1_05_in11 = reg_0473;
    11: op1_05_in11 = reg_0174;
    3: op1_05_in11 = reg_0167;
    12: op1_05_in11 = imem03_in[95:92];
    13: op1_05_in11 = reg_0265;
    14: op1_05_in11 = reg_0425;
    15: op1_05_in11 = reg_0644;
    16: op1_05_in11 = imem04_in[39:36];
    17: op1_05_in11 = reg_0479;
    18: op1_05_in11 = imem05_in[47:44];
    72: op1_05_in11 = imem05_in[47:44];
    2: op1_05_in11 = reg_0182;
    19: op1_05_in11 = reg_0478;
    20: op1_05_in11 = reg_0558;
    21: op1_05_in11 = reg_0477;
    22: op1_05_in11 = reg_0699;
    23: op1_05_in11 = reg_0748;
    24: op1_05_in11 = reg_0359;
    39: op1_05_in11 = reg_0359;
    25: op1_05_in11 = reg_0328;
    26: op1_05_in11 = reg_0349;
    27: op1_05_in11 = imem03_in[47:44];
    28: op1_05_in11 = reg_0673;
    29: op1_05_in11 = reg_0474;
    30: op1_05_in11 = reg_0008;
    31: op1_05_in11 = reg_0406;
    52: op1_05_in11 = reg_0406;
    32: op1_05_in11 = reg_0676;
    33: op1_05_in11 = reg_0361;
    35: op1_05_in11 = reg_0814;
    36: op1_05_in11 = reg_0440;
    38: op1_05_in11 = reg_0675;
    40: op1_05_in11 = reg_0476;
    41: op1_05_in11 = reg_0304;
    43: op1_05_in11 = reg_0679;
    44: op1_05_in11 = reg_0001;
    45: op1_05_in11 = reg_0155;
    46: op1_05_in11 = reg_0668;
    47: op1_05_in11 = reg_0667;
    48: op1_05_in11 = reg_0613;
    49: op1_05_in11 = reg_0627;
    50: op1_05_in11 = reg_0389;
    51: op1_05_in11 = reg_0194;
    53: op1_05_in11 = reg_0806;
    54: op1_05_in11 = imem05_in[79:76];
    55: op1_05_in11 = imem05_in[31:28];
    56: op1_05_in11 = reg_0776;
    58: op1_05_in11 = reg_0129;
    59: op1_05_in11 = reg_0688;
    60: op1_05_in11 = reg_0168;
    61: op1_05_in11 = reg_0469;
    62: op1_05_in11 = reg_0013;
    63: op1_05_in11 = reg_0292;
    64: op1_05_in11 = imem06_in[55:52];
    65: op1_05_in11 = imem06_in[75:72];
    66: op1_05_in11 = reg_0227;
    67: op1_05_in11 = imem07_in[31:28];
    68: op1_05_in11 = reg_0485;
    69: op1_05_in11 = reg_0617;
    70: op1_05_in11 = imem07_in[107:104];
    71: op1_05_in11 = imem04_in[127:124];
    73: op1_05_in11 = reg_0291;
    74: op1_05_in11 = reg_0441;
    75: op1_05_in11 = reg_0460;
    76: op1_05_in11 = reg_0200;
    77: op1_05_in11 = imem02_in[59:56];
    78: op1_05_in11 = reg_0797;
    79: op1_05_in11 = imem06_in[71:68];
    80: op1_05_in11 = reg_0729;
    81: op1_05_in11 = reg_0370;
    82: op1_05_in11 = reg_0081;
    83: op1_05_in11 = reg_0480;
    84: op1_05_in11 = reg_0113;
    86: op1_05_in11 = imem03_in[83:80];
    87: op1_05_in11 = reg_0305;
    88: op1_05_in11 = reg_0206;
    89: op1_05_in11 = imem06_in[63:60];
    90: op1_05_in11 = reg_0624;
    91: op1_05_in11 = reg_0276;
    92: op1_05_in11 = reg_0475;
    93: op1_05_in11 = reg_0195;
    94: op1_05_in11 = reg_0466;
    95: op1_05_in11 = reg_0468;
    96: op1_05_in11 = reg_0436;
    default: op1_05_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv11 = 1;
    6: op1_05_inv11 = 1;
    7: op1_05_inv11 = 1;
    8: op1_05_inv11 = 1;
    10: op1_05_inv11 = 1;
    11: op1_05_inv11 = 1;
    3: op1_05_inv11 = 1;
    12: op1_05_inv11 = 1;
    14: op1_05_inv11 = 1;
    16: op1_05_inv11 = 1;
    18: op1_05_inv11 = 1;
    2: op1_05_inv11 = 1;
    21: op1_05_inv11 = 1;
    23: op1_05_inv11 = 1;
    26: op1_05_inv11 = 1;
    27: op1_05_inv11 = 1;
    29: op1_05_inv11 = 1;
    30: op1_05_inv11 = 1;
    32: op1_05_inv11 = 1;
    38: op1_05_inv11 = 1;
    39: op1_05_inv11 = 1;
    40: op1_05_inv11 = 1;
    41: op1_05_inv11 = 1;
    46: op1_05_inv11 = 1;
    48: op1_05_inv11 = 1;
    50: op1_05_inv11 = 1;
    51: op1_05_inv11 = 1;
    52: op1_05_inv11 = 1;
    55: op1_05_inv11 = 1;
    56: op1_05_inv11 = 1;
    59: op1_05_inv11 = 1;
    60: op1_05_inv11 = 1;
    62: op1_05_inv11 = 1;
    65: op1_05_inv11 = 1;
    68: op1_05_inv11 = 1;
    72: op1_05_inv11 = 1;
    73: op1_05_inv11 = 1;
    79: op1_05_inv11 = 1;
    80: op1_05_inv11 = 1;
    83: op1_05_inv11 = 1;
    84: op1_05_inv11 = 1;
    86: op1_05_inv11 = 1;
    89: op1_05_inv11 = 1;
    90: op1_05_inv11 = 1;
    default: op1_05_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in12 = reg_0203;
    76: op1_05_in12 = reg_0203;
    95: op1_05_in12 = reg_0203;
    5: op1_05_in12 = reg_0726;
    6: op1_05_in12 = reg_0095;
    7: op1_05_in12 = reg_0142;
    8: op1_05_in12 = reg_0468;
    38: op1_05_in12 = reg_0468;
    9: op1_05_in12 = reg_0409;
    10: op1_05_in12 = reg_0467;
    11: op1_05_in12 = reg_0165;
    3: op1_05_in12 = reg_0177;
    12: op1_05_in12 = reg_0582;
    13: op1_05_in12 = reg_0732;
    14: op1_05_in12 = reg_0430;
    15: op1_05_in12 = reg_0358;
    16: op1_05_in12 = imem04_in[43:40];
    17: op1_05_in12 = reg_0478;
    18: op1_05_in12 = imem05_in[59:56];
    2: op1_05_in12 = reg_0160;
    19: op1_05_in12 = imem01_in[19:16];
    20: op1_05_in12 = reg_0551;
    21: op1_05_in12 = reg_0462;
    22: op1_05_in12 = reg_0461;
    23: op1_05_in12 = imem07_in[47:44];
    24: op1_05_in12 = reg_0345;
    25: op1_05_in12 = reg_0552;
    26: op1_05_in12 = reg_0348;
    27: op1_05_in12 = imem03_in[59:56];
    28: op1_05_in12 = reg_0463;
    29: op1_05_in12 = reg_0194;
    30: op1_05_in12 = reg_0010;
    31: op1_05_in12 = reg_0038;
    32: op1_05_in12 = reg_0670;
    33: op1_05_in12 = reg_0363;
    35: op1_05_in12 = reg_0339;
    36: op1_05_in12 = reg_0437;
    39: op1_05_in12 = reg_0356;
    40: op1_05_in12 = reg_0480;
    41: op1_05_in12 = reg_0309;
    43: op1_05_in12 = reg_0690;
    44: op1_05_in12 = reg_0803;
    45: op1_05_in12 = imem06_in[31:28];
    46: op1_05_in12 = reg_0477;
    47: op1_05_in12 = reg_0336;
    48: op1_05_in12 = reg_0605;
    49: op1_05_in12 = reg_0507;
    50: op1_05_in12 = reg_0007;
    51: op1_05_in12 = reg_0195;
    52: op1_05_in12 = reg_0590;
    53: op1_05_in12 = imem04_in[7:4];
    54: op1_05_in12 = imem05_in[87:84];
    55: op1_05_in12 = imem05_in[35:32];
    56: op1_05_in12 = reg_0242;
    91: op1_05_in12 = reg_0242;
    58: op1_05_in12 = reg_0131;
    59: op1_05_in12 = reg_0247;
    60: op1_05_in12 = reg_0171;
    61: op1_05_in12 = reg_0466;
    62: op1_05_in12 = reg_0804;
    63: op1_05_in12 = reg_0627;
    64: op1_05_in12 = imem06_in[115:112];
    65: op1_05_in12 = imem06_in[119:116];
    66: op1_05_in12 = reg_0075;
    67: op1_05_in12 = imem07_in[39:36];
    68: op1_05_in12 = reg_0565;
    69: op1_05_in12 = reg_0679;
    70: op1_05_in12 = reg_0704;
    71: op1_05_in12 = reg_0315;
    72: op1_05_in12 = imem05_in[55:52];
    73: op1_05_in12 = reg_0654;
    74: op1_05_in12 = reg_0333;
    75: op1_05_in12 = reg_0187;
    77: op1_05_in12 = imem02_in[75:72];
    78: op1_05_in12 = reg_0249;
    79: op1_05_in12 = imem06_in[75:72];
    80: op1_05_in12 = reg_0176;
    81: op1_05_in12 = reg_0814;
    82: op1_05_in12 = reg_0096;
    83: op1_05_in12 = reg_0474;
    84: op1_05_in12 = reg_0499;
    86: op1_05_in12 = imem03_in[107:104];
    87: op1_05_in12 = reg_0050;
    88: op1_05_in12 = imem01_in[71:68];
    89: op1_05_in12 = imem06_in[67:64];
    90: op1_05_in12 = reg_0817;
    92: op1_05_in12 = reg_0459;
    93: op1_05_in12 = reg_0199;
    94: op1_05_in12 = reg_0475;
    96: op1_05_in12 = reg_0636;
    default: op1_05_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv12 = 1;
    7: op1_05_inv12 = 1;
    8: op1_05_inv12 = 1;
    10: op1_05_inv12 = 1;
    14: op1_05_inv12 = 1;
    16: op1_05_inv12 = 1;
    17: op1_05_inv12 = 1;
    18: op1_05_inv12 = 1;
    2: op1_05_inv12 = 1;
    19: op1_05_inv12 = 1;
    20: op1_05_inv12 = 1;
    23: op1_05_inv12 = 1;
    24: op1_05_inv12 = 1;
    25: op1_05_inv12 = 1;
    27: op1_05_inv12 = 1;
    29: op1_05_inv12 = 1;
    30: op1_05_inv12 = 1;
    32: op1_05_inv12 = 1;
    39: op1_05_inv12 = 1;
    40: op1_05_inv12 = 1;
    43: op1_05_inv12 = 1;
    45: op1_05_inv12 = 1;
    47: op1_05_inv12 = 1;
    48: op1_05_inv12 = 1;
    50: op1_05_inv12 = 1;
    52: op1_05_inv12 = 1;
    53: op1_05_inv12 = 1;
    56: op1_05_inv12 = 1;
    60: op1_05_inv12 = 1;
    62: op1_05_inv12 = 1;
    63: op1_05_inv12 = 1;
    64: op1_05_inv12 = 1;
    65: op1_05_inv12 = 1;
    67: op1_05_inv12 = 1;
    68: op1_05_inv12 = 1;
    72: op1_05_inv12 = 1;
    74: op1_05_inv12 = 1;
    79: op1_05_inv12 = 1;
    82: op1_05_inv12 = 1;
    84: op1_05_inv12 = 1;
    88: op1_05_inv12 = 1;
    91: op1_05_inv12 = 1;
    92: op1_05_inv12 = 1;
    95: op1_05_inv12 = 1;
    default: op1_05_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in13 = reg_0190;
    5: op1_05_in13 = reg_0711;
    6: op1_05_in13 = reg_0096;
    7: op1_05_in13 = reg_0146;
    8: op1_05_in13 = reg_0479;
    10: op1_05_in13 = reg_0479;
    9: op1_05_in13 = reg_0371;
    3: op1_05_in13 = reg_0157;
    12: op1_05_in13 = reg_0572;
    13: op1_05_in13 = reg_0266;
    14: op1_05_in13 = reg_0447;
    15: op1_05_in13 = reg_0320;
    16: op1_05_in13 = imem04_in[119:116];
    17: op1_05_in13 = reg_0212;
    29: op1_05_in13 = reg_0212;
    18: op1_05_in13 = imem05_in[71:68];
    2: op1_05_in13 = reg_0176;
    19: op1_05_in13 = imem01_in[23:20];
    20: op1_05_in13 = reg_0559;
    21: op1_05_in13 = reg_0472;
    22: op1_05_in13 = reg_0476;
    23: op1_05_in13 = imem07_in[55:52];
    24: op1_05_in13 = reg_0353;
    25: op1_05_in13 = reg_0087;
    26: op1_05_in13 = reg_0361;
    68: op1_05_in13 = reg_0361;
    27: op1_05_in13 = imem03_in[63:60];
    28: op1_05_in13 = reg_0454;
    30: op1_05_in13 = imem04_in[7:4];
    31: op1_05_in13 = reg_0764;
    32: op1_05_in13 = reg_0677;
    33: op1_05_in13 = reg_0322;
    35: op1_05_in13 = reg_0367;
    36: op1_05_in13 = reg_0173;
    38: op1_05_in13 = reg_0187;
    39: op1_05_in13 = reg_0756;
    40: op1_05_in13 = reg_0468;
    41: op1_05_in13 = reg_0527;
    43: op1_05_in13 = reg_0455;
    44: op1_05_in13 = reg_0804;
    50: op1_05_in13 = reg_0804;
    45: op1_05_in13 = imem06_in[87:84];
    46: op1_05_in13 = reg_0469;
    47: op1_05_in13 = reg_0341;
    48: op1_05_in13 = reg_0762;
    49: op1_05_in13 = reg_0068;
    51: op1_05_in13 = reg_0199;
    52: op1_05_in13 = reg_0314;
    53: op1_05_in13 = imem04_in[51:48];
    54: op1_05_in13 = reg_0798;
    55: op1_05_in13 = imem05_in[51:48];
    56: op1_05_in13 = reg_0819;
    58: op1_05_in13 = reg_0144;
    59: op1_05_in13 = reg_0692;
    61: op1_05_in13 = reg_0480;
    62: op1_05_in13 = imem04_in[23:20];
    63: op1_05_in13 = reg_0508;
    64: op1_05_in13 = imem06_in[127:124];
    65: op1_05_in13 = reg_0624;
    66: op1_05_in13 = reg_0246;
    67: op1_05_in13 = imem07_in[51:48];
    69: op1_05_in13 = reg_0687;
    70: op1_05_in13 = reg_0719;
    71: op1_05_in13 = reg_0560;
    72: op1_05_in13 = reg_0307;
    73: op1_05_in13 = reg_0775;
    74: op1_05_in13 = reg_0438;
    75: op1_05_in13 = reg_0193;
    76: op1_05_in13 = reg_0201;
    77: op1_05_in13 = imem02_in[95:92];
    78: op1_05_in13 = reg_0786;
    79: op1_05_in13 = reg_0289;
    80: op1_05_in13 = reg_0712;
    81: op1_05_in13 = reg_0298;
    90: op1_05_in13 = reg_0298;
    82: op1_05_in13 = reg_0740;
    83: op1_05_in13 = reg_0478;
    84: op1_05_in13 = reg_0782;
    86: op1_05_in13 = imem03_in[119:116];
    87: op1_05_in13 = reg_0626;
    88: op1_05_in13 = imem01_in[123:120];
    89: op1_05_in13 = imem06_in[75:72];
    91: op1_05_in13 = reg_0576;
    92: op1_05_in13 = reg_0452;
    93: op1_05_in13 = reg_0422;
    94: op1_05_in13 = reg_0462;
    95: op1_05_in13 = reg_0211;
    96: op1_05_in13 = reg_0434;
    default: op1_05_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv13 = 1;
    6: op1_05_inv13 = 1;
    7: op1_05_inv13 = 1;
    8: op1_05_inv13 = 1;
    10: op1_05_inv13 = 1;
    12: op1_05_inv13 = 1;
    13: op1_05_inv13 = 1;
    14: op1_05_inv13 = 1;
    16: op1_05_inv13 = 1;
    18: op1_05_inv13 = 1;
    22: op1_05_inv13 = 1;
    25: op1_05_inv13 = 1;
    26: op1_05_inv13 = 1;
    35: op1_05_inv13 = 1;
    40: op1_05_inv13 = 1;
    41: op1_05_inv13 = 1;
    43: op1_05_inv13 = 1;
    46: op1_05_inv13 = 1;
    52: op1_05_inv13 = 1;
    53: op1_05_inv13 = 1;
    55: op1_05_inv13 = 1;
    58: op1_05_inv13 = 1;
    59: op1_05_inv13 = 1;
    61: op1_05_inv13 = 1;
    62: op1_05_inv13 = 1;
    64: op1_05_inv13 = 1;
    68: op1_05_inv13 = 1;
    71: op1_05_inv13 = 1;
    77: op1_05_inv13 = 1;
    78: op1_05_inv13 = 1;
    79: op1_05_inv13 = 1;
    81: op1_05_inv13 = 1;
    84: op1_05_inv13 = 1;
    86: op1_05_inv13 = 1;
    87: op1_05_inv13 = 1;
    93: op1_05_inv13 = 1;
    94: op1_05_inv13 = 1;
    default: op1_05_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in14 = reg_0202;
    5: op1_05_in14 = reg_0727;
    6: op1_05_in14 = reg_0086;
    7: op1_05_in14 = reg_0139;
    8: op1_05_in14 = reg_0187;
    9: op1_05_in14 = reg_0375;
    10: op1_05_in14 = reg_0208;
    3: op1_05_in14 = reg_0173;
    12: op1_05_in14 = reg_0588;
    13: op1_05_in14 = reg_0149;
    14: op1_05_in14 = reg_0419;
    15: op1_05_in14 = reg_0341;
    16: op1_05_in14 = reg_0552;
    71: op1_05_in14 = reg_0552;
    17: op1_05_in14 = reg_0205;
    18: op1_05_in14 = imem05_in[119:116];
    19: op1_05_in14 = imem01_in[39:36];
    20: op1_05_in14 = reg_0547;
    21: op1_05_in14 = reg_0473;
    22: op1_05_in14 = reg_0475;
    23: op1_05_in14 = imem07_in[59:56];
    24: op1_05_in14 = reg_0350;
    25: op1_05_in14 = reg_0056;
    26: op1_05_in14 = reg_0363;
    27: op1_05_in14 = imem03_in[71:68];
    28: op1_05_in14 = reg_0481;
    29: op1_05_in14 = reg_0197;
    30: op1_05_in14 = imem04_in[11:8];
    31: op1_05_in14 = reg_0576;
    32: op1_05_in14 = reg_0678;
    33: op1_05_in14 = reg_0355;
    35: op1_05_in14 = imem07_in[43:40];
    38: op1_05_in14 = reg_0204;
    39: op1_05_in14 = reg_0538;
    40: op1_05_in14 = reg_0478;
    41: op1_05_in14 = reg_0733;
    43: op1_05_in14 = reg_0472;
    94: op1_05_in14 = reg_0472;
    44: op1_05_in14 = imem04_in[31:28];
    45: op1_05_in14 = reg_0299;
    46: op1_05_in14 = reg_0462;
    47: op1_05_in14 = reg_0345;
    48: op1_05_in14 = reg_0377;
    49: op1_05_in14 = reg_0640;
    50: op1_05_in14 = reg_0801;
    51: op1_05_in14 = reg_0192;
    52: op1_05_in14 = reg_0535;
    53: op1_05_in14 = imem04_in[59:56];
    54: op1_05_in14 = reg_0483;
    55: op1_05_in14 = imem05_in[63:60];
    56: op1_05_in14 = reg_0236;
    58: op1_05_in14 = imem06_in[51:48];
    59: op1_05_in14 = reg_0453;
    61: op1_05_in14 = reg_0474;
    62: op1_05_in14 = imem04_in[51:48];
    63: op1_05_in14 = reg_0679;
    64: op1_05_in14 = reg_0238;
    65: op1_05_in14 = reg_0349;
    66: op1_05_in14 = reg_0797;
    67: op1_05_in14 = imem07_in[95:92];
    68: op1_05_in14 = reg_0351;
    69: op1_05_in14 = reg_0296;
    70: op1_05_in14 = reg_0717;
    72: op1_05_in14 = reg_0066;
    78: op1_05_in14 = reg_0066;
    73: op1_05_in14 = reg_0821;
    74: op1_05_in14 = reg_0268;
    75: op1_05_in14 = reg_0186;
    76: op1_05_in14 = imem01_in[19:16];
    77: op1_05_in14 = imem02_in[107:104];
    79: op1_05_in14 = reg_0348;
    80: op1_05_in14 = reg_0713;
    81: op1_05_in14 = reg_0766;
    82: op1_05_in14 = imem03_in[43:40];
    83: op1_05_in14 = reg_0210;
    84: op1_05_in14 = reg_0732;
    86: op1_05_in14 = imem03_in[123:120];
    87: op1_05_in14 = reg_0065;
    88: op1_05_in14 = reg_0653;
    89: op1_05_in14 = imem06_in[83:80];
    90: op1_05_in14 = reg_0619;
    91: op1_05_in14 = reg_0515;
    92: op1_05_in14 = reg_0456;
    93: op1_05_in14 = reg_0152;
    95: op1_05_in14 = reg_0201;
    96: op1_05_in14 = reg_0444;
    default: op1_05_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv14 = 1;
    6: op1_05_inv14 = 1;
    8: op1_05_inv14 = 1;
    9: op1_05_inv14 = 1;
    10: op1_05_inv14 = 1;
    16: op1_05_inv14 = 1;
    21: op1_05_inv14 = 1;
    23: op1_05_inv14 = 1;
    24: op1_05_inv14 = 1;
    25: op1_05_inv14 = 1;
    26: op1_05_inv14 = 1;
    28: op1_05_inv14 = 1;
    31: op1_05_inv14 = 1;
    32: op1_05_inv14 = 1;
    35: op1_05_inv14 = 1;
    38: op1_05_inv14 = 1;
    39: op1_05_inv14 = 1;
    40: op1_05_inv14 = 1;
    44: op1_05_inv14 = 1;
    45: op1_05_inv14 = 1;
    46: op1_05_inv14 = 1;
    47: op1_05_inv14 = 1;
    48: op1_05_inv14 = 1;
    53: op1_05_inv14 = 1;
    58: op1_05_inv14 = 1;
    61: op1_05_inv14 = 1;
    62: op1_05_inv14 = 1;
    64: op1_05_inv14 = 1;
    65: op1_05_inv14 = 1;
    66: op1_05_inv14 = 1;
    68: op1_05_inv14 = 1;
    69: op1_05_inv14 = 1;
    70: op1_05_inv14 = 1;
    72: op1_05_inv14 = 1;
    77: op1_05_inv14 = 1;
    78: op1_05_inv14 = 1;
    79: op1_05_inv14 = 1;
    80: op1_05_inv14 = 1;
    82: op1_05_inv14 = 1;
    87: op1_05_inv14 = 1;
    89: op1_05_inv14 = 1;
    91: op1_05_inv14 = 1;
    94: op1_05_inv14 = 1;
    95: op1_05_inv14 = 1;
    96: op1_05_inv14 = 1;
    default: op1_05_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in15 = imem01_in[19:16];
    5: op1_05_in15 = reg_0424;
    6: op1_05_in15 = imem03_in[31:28];
    7: op1_05_in15 = reg_0141;
    8: op1_05_in15 = reg_0188;
    93: op1_05_in15 = reg_0188;
    9: op1_05_in15 = reg_0382;
    10: op1_05_in15 = reg_0191;
    12: op1_05_in15 = reg_0384;
    13: op1_05_in15 = reg_0128;
    14: op1_05_in15 = reg_0442;
    15: op1_05_in15 = reg_0359;
    16: op1_05_in15 = reg_0542;
    17: op1_05_in15 = reg_0190;
    18: op1_05_in15 = imem05_in[123:120];
    19: op1_05_in15 = reg_0522;
    20: op1_05_in15 = reg_0079;
    21: op1_05_in15 = reg_0470;
    22: op1_05_in15 = reg_0474;
    23: op1_05_in15 = imem07_in[67:64];
    24: op1_05_in15 = reg_0347;
    25: op1_05_in15 = reg_0555;
    26: op1_05_in15 = reg_0350;
    27: op1_05_in15 = imem03_in[75:72];
    28: op1_05_in15 = reg_0471;
    61: op1_05_in15 = reg_0471;
    29: op1_05_in15 = imem01_in[3:0];
    30: op1_05_in15 = imem04_in[83:80];
    31: op1_05_in15 = imem06_in[11:8];
    32: op1_05_in15 = reg_0675;
    33: op1_05_in15 = reg_0073;
    35: op1_05_in15 = imem07_in[47:44];
    38: op1_05_in15 = reg_0211;
    39: op1_05_in15 = imem03_in[35:32];
    40: op1_05_in15 = reg_0204;
    41: op1_05_in15 = reg_0224;
    43: op1_05_in15 = reg_0452;
    44: op1_05_in15 = imem04_in[55:52];
    45: op1_05_in15 = reg_0625;
    46: op1_05_in15 = reg_0481;
    47: op1_05_in15 = reg_0324;
    48: op1_05_in15 = reg_0319;
    49: op1_05_in15 = reg_0260;
    50: op1_05_in15 = reg_0809;
    51: op1_05_in15 = imem01_in[39:36];
    52: op1_05_in15 = reg_0770;
    53: op1_05_in15 = imem04_in[75:72];
    54: op1_05_in15 = reg_0793;
    55: op1_05_in15 = imem05_in[75:72];
    56: op1_05_in15 = reg_0623;
    58: op1_05_in15 = reg_0289;
    59: op1_05_in15 = reg_0469;
    62: op1_05_in15 = imem04_in[67:64];
    63: op1_05_in15 = reg_0078;
    64: op1_05_in15 = reg_0766;
    65: op1_05_in15 = reg_0605;
    66: op1_05_in15 = reg_0309;
    67: op1_05_in15 = imem07_in[115:112];
    68: op1_05_in15 = reg_0414;
    69: op1_05_in15 = imem05_in[35:32];
    70: op1_05_in15 = reg_0713;
    71: op1_05_in15 = reg_0523;
    72: op1_05_in15 = reg_0149;
    73: op1_05_in15 = reg_0748;
    74: op1_05_in15 = reg_0175;
    75: op1_05_in15 = reg_0205;
    76: op1_05_in15 = imem01_in[23:20];
    77: op1_05_in15 = imem02_in[111:108];
    78: op1_05_in15 = reg_0795;
    79: op1_05_in15 = reg_0115;
    80: op1_05_in15 = reg_0711;
    81: op1_05_in15 = reg_0401;
    90: op1_05_in15 = reg_0401;
    82: op1_05_in15 = imem03_in[71:68];
    83: op1_05_in15 = reg_0209;
    92: op1_05_in15 = reg_0209;
    84: op1_05_in15 = reg_0326;
    86: op1_05_in15 = reg_0582;
    87: op1_05_in15 = reg_0371;
    88: op1_05_in15 = reg_0759;
    89: op1_05_in15 = imem06_in[95:92];
    91: op1_05_in15 = reg_0612;
    94: op1_05_in15 = reg_0459;
    95: op1_05_in15 = reg_0206;
    96: op1_05_in15 = reg_0443;
    default: op1_05_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv15 = 1;
    9: op1_05_inv15 = 1;
    13: op1_05_inv15 = 1;
    17: op1_05_inv15 = 1;
    20: op1_05_inv15 = 1;
    22: op1_05_inv15 = 1;
    23: op1_05_inv15 = 1;
    27: op1_05_inv15 = 1;
    28: op1_05_inv15 = 1;
    30: op1_05_inv15 = 1;
    32: op1_05_inv15 = 1;
    33: op1_05_inv15 = 1;
    41: op1_05_inv15 = 1;
    43: op1_05_inv15 = 1;
    45: op1_05_inv15 = 1;
    46: op1_05_inv15 = 1;
    47: op1_05_inv15 = 1;
    48: op1_05_inv15 = 1;
    50: op1_05_inv15 = 1;
    51: op1_05_inv15 = 1;
    52: op1_05_inv15 = 1;
    53: op1_05_inv15 = 1;
    54: op1_05_inv15 = 1;
    55: op1_05_inv15 = 1;
    56: op1_05_inv15 = 1;
    61: op1_05_inv15 = 1;
    62: op1_05_inv15 = 1;
    63: op1_05_inv15 = 1;
    65: op1_05_inv15 = 1;
    68: op1_05_inv15 = 1;
    69: op1_05_inv15 = 1;
    70: op1_05_inv15 = 1;
    72: op1_05_inv15 = 1;
    74: op1_05_inv15 = 1;
    75: op1_05_inv15 = 1;
    80: op1_05_inv15 = 1;
    81: op1_05_inv15 = 1;
    83: op1_05_inv15 = 1;
    84: op1_05_inv15 = 1;
    87: op1_05_inv15 = 1;
    89: op1_05_inv15 = 1;
    90: op1_05_inv15 = 1;
    92: op1_05_inv15 = 1;
    94: op1_05_inv15 = 1;
    95: op1_05_inv15 = 1;
    default: op1_05_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in16 = imem01_in[63:60];
    5: op1_05_in16 = reg_0419;
    6: op1_05_in16 = imem03_in[35:32];
    7: op1_05_in16 = reg_0137;
    8: op1_05_in16 = reg_0203;
    9: op1_05_in16 = reg_0406;
    10: op1_05_in16 = reg_0188;
    43: op1_05_in16 = reg_0188;
    12: op1_05_in16 = reg_0388;
    13: op1_05_in16 = reg_0154;
    14: op1_05_in16 = reg_0427;
    15: op1_05_in16 = reg_0318;
    16: op1_05_in16 = reg_0549;
    17: op1_05_in16 = reg_0197;
    18: op1_05_in16 = reg_0798;
    19: op1_05_in16 = reg_0497;
    20: op1_05_in16 = reg_0253;
    21: op1_05_in16 = reg_0452;
    22: op1_05_in16 = reg_0471;
    23: op1_05_in16 = imem07_in[87:84];
    24: op1_05_in16 = reg_0533;
    25: op1_05_in16 = reg_0283;
    26: op1_05_in16 = reg_0530;
    27: op1_05_in16 = imem03_in[83:80];
    28: op1_05_in16 = reg_0479;
    29: op1_05_in16 = imem01_in[15:12];
    30: op1_05_in16 = imem04_in[87:84];
    31: op1_05_in16 = imem06_in[23:20];
    32: op1_05_in16 = reg_0669;
    33: op1_05_in16 = reg_0347;
    35: op1_05_in16 = imem07_in[59:56];
    38: op1_05_in16 = reg_0198;
    39: op1_05_in16 = imem03_in[43:40];
    40: op1_05_in16 = reg_0503;
    41: op1_05_in16 = reg_0260;
    44: op1_05_in16 = imem04_in[63:60];
    45: op1_05_in16 = reg_0604;
    86: op1_05_in16 = reg_0604;
    46: op1_05_in16 = reg_0472;
    47: op1_05_in16 = reg_0323;
    48: op1_05_in16 = reg_0038;
    49: op1_05_in16 = reg_0527;
    68: op1_05_in16 = reg_0527;
    50: op1_05_in16 = reg_0004;
    51: op1_05_in16 = imem01_in[59:56];
    52: op1_05_in16 = imem03_in[51:48];
    53: op1_05_in16 = imem04_in[91:88];
    54: op1_05_in16 = reg_0794;
    55: op1_05_in16 = imem05_in[87:84];
    56: op1_05_in16 = imem07_in[15:12];
    58: op1_05_in16 = reg_0299;
    59: op1_05_in16 = reg_0470;
    61: op1_05_in16 = reg_0189;
    62: op1_05_in16 = imem04_in[99:96];
    63: op1_05_in16 = reg_0622;
    64: op1_05_in16 = reg_0339;
    65: op1_05_in16 = reg_0817;
    66: op1_05_in16 = reg_0279;
    67: op1_05_in16 = reg_0725;
    69: op1_05_in16 = imem05_in[51:48];
    70: op1_05_in16 = reg_0715;
    71: op1_05_in16 = reg_0076;
    72: op1_05_in16 = reg_0155;
    73: op1_05_in16 = reg_0593;
    74: op1_05_in16 = reg_0161;
    75: op1_05_in16 = reg_0206;
    76: op1_05_in16 = imem01_in[27:24];
    77: op1_05_in16 = reg_0739;
    78: op1_05_in16 = reg_0793;
    79: op1_05_in16 = reg_0624;
    80: op1_05_in16 = reg_0103;
    81: op1_05_in16 = reg_0031;
    82: op1_05_in16 = imem03_in[91:88];
    83: op1_05_in16 = imem01_in[55:52];
    84: op1_05_in16 = reg_0245;
    87: op1_05_in16 = reg_0774;
    88: op1_05_in16 = reg_0235;
    89: op1_05_in16 = imem06_in[107:104];
    90: op1_05_in16 = reg_0402;
    91: op1_05_in16 = reg_0777;
    92: op1_05_in16 = reg_0211;
    93: op1_05_in16 = reg_0243;
    94: op1_05_in16 = reg_0208;
    95: op1_05_in16 = reg_0422;
    96: op1_05_in16 = reg_0089;
    default: op1_05_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv16 = 1;
    9: op1_05_inv16 = 1;
    15: op1_05_inv16 = 1;
    16: op1_05_inv16 = 1;
    17: op1_05_inv16 = 1;
    19: op1_05_inv16 = 1;
    20: op1_05_inv16 = 1;
    21: op1_05_inv16 = 1;
    24: op1_05_inv16 = 1;
    26: op1_05_inv16 = 1;
    27: op1_05_inv16 = 1;
    29: op1_05_inv16 = 1;
    33: op1_05_inv16 = 1;
    39: op1_05_inv16 = 1;
    40: op1_05_inv16 = 1;
    43: op1_05_inv16 = 1;
    46: op1_05_inv16 = 1;
    48: op1_05_inv16 = 1;
    49: op1_05_inv16 = 1;
    51: op1_05_inv16 = 1;
    53: op1_05_inv16 = 1;
    54: op1_05_inv16 = 1;
    58: op1_05_inv16 = 1;
    63: op1_05_inv16 = 1;
    65: op1_05_inv16 = 1;
    70: op1_05_inv16 = 1;
    73: op1_05_inv16 = 1;
    76: op1_05_inv16 = 1;
    77: op1_05_inv16 = 1;
    78: op1_05_inv16 = 1;
    81: op1_05_inv16 = 1;
    83: op1_05_inv16 = 1;
    84: op1_05_inv16 = 1;
    88: op1_05_inv16 = 1;
    90: op1_05_inv16 = 1;
    92: op1_05_inv16 = 1;
    94: op1_05_inv16 = 1;
    95: op1_05_inv16 = 1;
    default: op1_05_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in17 = imem01_in[91:88];
    5: op1_05_in17 = reg_0439;
    6: op1_05_in17 = imem03_in[63:60];
    7: op1_05_in17 = imem06_in[19:16];
    8: op1_05_in17 = reg_0207;
    61: op1_05_in17 = reg_0207;
    9: op1_05_in17 = reg_0028;
    10: op1_05_in17 = reg_0203;
    12: op1_05_in17 = reg_0373;
    13: op1_05_in17 = reg_0153;
    14: op1_05_in17 = reg_0172;
    15: op1_05_in17 = reg_0092;
    33: op1_05_in17 = reg_0092;
    16: op1_05_in17 = reg_0546;
    17: op1_05_in17 = imem01_in[67:64];
    18: op1_05_in17 = reg_0488;
    19: op1_05_in17 = reg_0229;
    66: op1_05_in17 = reg_0229;
    20: op1_05_in17 = reg_0299;
    21: op1_05_in17 = reg_0458;
    22: op1_05_in17 = reg_0186;
    23: op1_05_in17 = imem07_in[95:92];
    24: op1_05_in17 = reg_0080;
    25: op1_05_in17 = reg_0280;
    26: op1_05_in17 = reg_0769;
    27: op1_05_in17 = imem03_in[87:84];
    28: op1_05_in17 = reg_0478;
    29: op1_05_in17 = imem01_in[35:32];
    30: op1_05_in17 = imem04_in[107:104];
    31: op1_05_in17 = imem06_in[67:64];
    32: op1_05_in17 = reg_0461;
    35: op1_05_in17 = imem07_in[127:124];
    38: op1_05_in17 = reg_0195;
    39: op1_05_in17 = imem03_in[103:100];
    40: op1_05_in17 = reg_0233;
    41: op1_05_in17 = reg_0744;
    43: op1_05_in17 = imem01_in[51:48];
    75: op1_05_in17 = imem01_in[51:48];
    44: op1_05_in17 = imem04_in[67:64];
    45: op1_05_in17 = reg_0291;
    46: op1_05_in17 = reg_0208;
    47: op1_05_in17 = reg_0518;
    48: op1_05_in17 = reg_0401;
    49: op1_05_in17 = reg_0272;
    50: op1_05_in17 = imem04_in[3:0];
    51: op1_05_in17 = imem01_in[83:80];
    83: op1_05_in17 = imem01_in[83:80];
    52: op1_05_in17 = imem03_in[59:56];
    53: op1_05_in17 = imem04_in[95:92];
    54: op1_05_in17 = reg_0090;
    55: op1_05_in17 = imem05_in[103:100];
    56: op1_05_in17 = imem07_in[23:20];
    58: op1_05_in17 = reg_0605;
    59: op1_05_in17 = reg_0479;
    62: op1_05_in17 = imem04_in[115:112];
    63: op1_05_in17 = reg_0644;
    64: op1_05_in17 = reg_0578;
    65: op1_05_in17 = reg_0609;
    67: op1_05_in17 = reg_0729;
    68: op1_05_in17 = reg_0406;
    69: op1_05_in17 = imem05_in[91:88];
    70: op1_05_in17 = reg_0727;
    80: op1_05_in17 = reg_0727;
    71: op1_05_in17 = reg_0292;
    72: op1_05_in17 = imem06_in[39:36];
    73: op1_05_in17 = reg_0576;
    74: op1_05_in17 = reg_0167;
    76: op1_05_in17 = imem01_in[55:52];
    77: op1_05_in17 = reg_0392;
    78: op1_05_in17 = reg_0665;
    79: op1_05_in17 = reg_0817;
    81: op1_05_in17 = reg_0748;
    82: op1_05_in17 = reg_0582;
    84: op1_05_in17 = reg_0389;
    86: op1_05_in17 = reg_0559;
    87: op1_05_in17 = reg_0640;
    88: op1_05_in17 = reg_0306;
    89: op1_05_in17 = imem06_in[115:112];
    90: op1_05_in17 = reg_0628;
    91: op1_05_in17 = reg_0664;
    92: op1_05_in17 = reg_0198;
    93: op1_05_in17 = imem01_in[7:4];
    94: op1_05_in17 = reg_0210;
    95: op1_05_in17 = reg_0114;
    96: op1_05_in17 = reg_0181;
    default: op1_05_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv17 = 1;
    7: op1_05_inv17 = 1;
    8: op1_05_inv17 = 1;
    13: op1_05_inv17 = 1;
    17: op1_05_inv17 = 1;
    18: op1_05_inv17 = 1;
    19: op1_05_inv17 = 1;
    20: op1_05_inv17 = 1;
    25: op1_05_inv17 = 1;
    28: op1_05_inv17 = 1;
    29: op1_05_inv17 = 1;
    30: op1_05_inv17 = 1;
    32: op1_05_inv17 = 1;
    35: op1_05_inv17 = 1;
    39: op1_05_inv17 = 1;
    43: op1_05_inv17 = 1;
    44: op1_05_inv17 = 1;
    48: op1_05_inv17 = 1;
    49: op1_05_inv17 = 1;
    50: op1_05_inv17 = 1;
    51: op1_05_inv17 = 1;
    53: op1_05_inv17 = 1;
    56: op1_05_inv17 = 1;
    59: op1_05_inv17 = 1;
    65: op1_05_inv17 = 1;
    66: op1_05_inv17 = 1;
    67: op1_05_inv17 = 1;
    68: op1_05_inv17 = 1;
    69: op1_05_inv17 = 1;
    70: op1_05_inv17 = 1;
    71: op1_05_inv17 = 1;
    72: op1_05_inv17 = 1;
    74: op1_05_inv17 = 1;
    75: op1_05_inv17 = 1;
    76: op1_05_inv17 = 1;
    77: op1_05_inv17 = 1;
    78: op1_05_inv17 = 1;
    79: op1_05_inv17 = 1;
    80: op1_05_inv17 = 1;
    81: op1_05_inv17 = 1;
    83: op1_05_inv17 = 1;
    87: op1_05_inv17 = 1;
    88: op1_05_inv17 = 1;
    89: op1_05_inv17 = 1;
    90: op1_05_inv17 = 1;
    92: op1_05_inv17 = 1;
    94: op1_05_inv17 = 1;
    96: op1_05_inv17 = 1;
    default: op1_05_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in18 = reg_0504;
    5: op1_05_in18 = reg_0440;
    6: op1_05_in18 = imem03_in[91:88];
    7: op1_05_in18 = imem06_in[23:20];
    8: op1_05_in18 = reg_0186;
    9: op1_05_in18 = reg_0813;
    10: op1_05_in18 = reg_0207;
    12: op1_05_in18 = reg_0398;
    13: op1_05_in18 = reg_0130;
    14: op1_05_in18 = reg_0167;
    15: op1_05_in18 = reg_0091;
    16: op1_05_in18 = reg_0308;
    17: op1_05_in18 = imem01_in[83:80];
    18: op1_05_in18 = reg_0788;
    19: op1_05_in18 = reg_0820;
    20: op1_05_in18 = reg_0296;
    21: op1_05_in18 = reg_0191;
    22: op1_05_in18 = reg_0199;
    38: op1_05_in18 = reg_0199;
    23: op1_05_in18 = reg_0728;
    24: op1_05_in18 = reg_0530;
    25: op1_05_in18 = reg_0291;
    26: op1_05_in18 = reg_0098;
    27: op1_05_in18 = imem03_in[99:96];
    52: op1_05_in18 = imem03_in[99:96];
    28: op1_05_in18 = reg_0200;
    59: op1_05_in18 = reg_0200;
    29: op1_05_in18 = imem01_in[63:60];
    30: op1_05_in18 = imem04_in[111:108];
    31: op1_05_in18 = imem06_in[71:68];
    32: op1_05_in18 = reg_0462;
    33: op1_05_in18 = reg_0533;
    35: op1_05_in18 = reg_0704;
    39: op1_05_in18 = reg_0582;
    40: op1_05_in18 = reg_0237;
    41: op1_05_in18 = reg_0137;
    43: op1_05_in18 = imem01_in[111:108];
    44: op1_05_in18 = imem04_in[79:76];
    45: op1_05_in18 = reg_0613;
    46: op1_05_in18 = reg_0190;
    61: op1_05_in18 = reg_0190;
    47: op1_05_in18 = imem03_in[31:28];
    48: op1_05_in18 = reg_0368;
    49: op1_05_in18 = reg_0039;
    50: op1_05_in18 = imem04_in[11:8];
    51: op1_05_in18 = reg_0772;
    53: op1_05_in18 = imem04_in[107:104];
    54: op1_05_in18 = reg_0309;
    55: op1_05_in18 = imem05_in[119:116];
    56: op1_05_in18 = imem07_in[39:36];
    58: op1_05_in18 = reg_0298;
    65: op1_05_in18 = reg_0298;
    62: op1_05_in18 = reg_0315;
    63: op1_05_in18 = reg_0416;
    64: op1_05_in18 = reg_0659;
    66: op1_05_in18 = reg_0132;
    67: op1_05_in18 = reg_0713;
    68: op1_05_in18 = reg_0514;
    69: op1_05_in18 = imem05_in[115:112];
    70: op1_05_in18 = reg_0441;
    71: op1_05_in18 = reg_0431;
    72: op1_05_in18 = imem06_in[47:44];
    73: op1_05_in18 = reg_0563;
    74: op1_05_in18 = reg_0163;
    75: op1_05_in18 = imem01_in[67:64];
    76: op1_05_in18 = imem01_in[67:64];
    77: op1_05_in18 = reg_0139;
    78: op1_05_in18 = reg_0134;
    79: op1_05_in18 = reg_0370;
    80: op1_05_in18 = reg_0635;
    81: op1_05_in18 = reg_0270;
    82: op1_05_in18 = reg_0588;
    83: op1_05_in18 = imem01_in[91:88];
    84: op1_05_in18 = reg_0781;
    86: op1_05_in18 = reg_0319;
    87: op1_05_in18 = reg_0233;
    88: op1_05_in18 = reg_0422;
    89: op1_05_in18 = reg_0814;
    90: op1_05_in18 = reg_0405;
    91: op1_05_in18 = reg_0037;
    92: op1_05_in18 = reg_0196;
    93: op1_05_in18 = imem01_in[47:44];
    94: op1_05_in18 = reg_0241;
    95: op1_05_in18 = reg_0506;
    96: op1_05_in18 = reg_0327;
    default: op1_05_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv18 = 1;
    5: op1_05_inv18 = 1;
    6: op1_05_inv18 = 1;
    8: op1_05_inv18 = 1;
    9: op1_05_inv18 = 1;
    10: op1_05_inv18 = 1;
    12: op1_05_inv18 = 1;
    13: op1_05_inv18 = 1;
    14: op1_05_inv18 = 1;
    15: op1_05_inv18 = 1;
    17: op1_05_inv18 = 1;
    23: op1_05_inv18 = 1;
    24: op1_05_inv18 = 1;
    27: op1_05_inv18 = 1;
    28: op1_05_inv18 = 1;
    29: op1_05_inv18 = 1;
    30: op1_05_inv18 = 1;
    33: op1_05_inv18 = 1;
    38: op1_05_inv18 = 1;
    39: op1_05_inv18 = 1;
    43: op1_05_inv18 = 1;
    44: op1_05_inv18 = 1;
    45: op1_05_inv18 = 1;
    48: op1_05_inv18 = 1;
    49: op1_05_inv18 = 1;
    51: op1_05_inv18 = 1;
    53: op1_05_inv18 = 1;
    54: op1_05_inv18 = 1;
    55: op1_05_inv18 = 1;
    58: op1_05_inv18 = 1;
    59: op1_05_inv18 = 1;
    61: op1_05_inv18 = 1;
    63: op1_05_inv18 = 1;
    65: op1_05_inv18 = 1;
    67: op1_05_inv18 = 1;
    68: op1_05_inv18 = 1;
    71: op1_05_inv18 = 1;
    74: op1_05_inv18 = 1;
    75: op1_05_inv18 = 1;
    76: op1_05_inv18 = 1;
    77: op1_05_inv18 = 1;
    78: op1_05_inv18 = 1;
    79: op1_05_inv18 = 1;
    80: op1_05_inv18 = 1;
    83: op1_05_inv18 = 1;
    84: op1_05_inv18 = 1;
    89: op1_05_inv18 = 1;
    95: op1_05_inv18 = 1;
    default: op1_05_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in19 = reg_0515;
    5: op1_05_in19 = reg_0427;
    6: op1_05_in19 = imem03_in[115:112];
    7: op1_05_in19 = imem06_in[35:32];
    8: op1_05_in19 = reg_0192;
    38: op1_05_in19 = reg_0192;
    9: op1_05_in19 = reg_0040;
    10: op1_05_in19 = reg_0212;
    12: op1_05_in19 = reg_0012;
    27: op1_05_in19 = reg_0012;
    13: op1_05_in19 = reg_0131;
    14: op1_05_in19 = reg_0169;
    15: op1_05_in19 = reg_0084;
    16: op1_05_in19 = reg_0305;
    17: op1_05_in19 = imem01_in[127:124];
    18: op1_05_in19 = reg_0494;
    19: op1_05_in19 = reg_0227;
    20: op1_05_in19 = reg_0074;
    21: op1_05_in19 = reg_0210;
    22: op1_05_in19 = imem01_in[3:0];
    23: op1_05_in19 = reg_0704;
    24: op1_05_in19 = reg_0539;
    25: op1_05_in19 = reg_0266;
    26: op1_05_in19 = reg_0740;
    28: op1_05_in19 = reg_0189;
    29: op1_05_in19 = imem01_in[67:64];
    30: op1_05_in19 = reg_0059;
    31: op1_05_in19 = imem06_in[75:72];
    32: op1_05_in19 = reg_0472;
    33: op1_05_in19 = reg_0097;
    35: op1_05_in19 = reg_0723;
    39: op1_05_in19 = reg_0599;
    40: op1_05_in19 = reg_0758;
    41: op1_05_in19 = reg_0134;
    43: op1_05_in19 = reg_0336;
    44: op1_05_in19 = reg_0316;
    45: op1_05_in19 = reg_0608;
    46: op1_05_in19 = reg_0197;
    47: op1_05_in19 = imem03_in[35:32];
    48: op1_05_in19 = imem07_in[39:36];
    49: op1_05_in19 = reg_0323;
    50: op1_05_in19 = imem04_in[59:56];
    51: op1_05_in19 = reg_0820;
    52: op1_05_in19 = imem03_in[127:124];
    53: op1_05_in19 = imem04_in[115:112];
    54: op1_05_in19 = reg_0226;
    55: op1_05_in19 = reg_0307;
    56: op1_05_in19 = imem07_in[91:88];
    58: op1_05_in19 = reg_0038;
    59: op1_05_in19 = reg_0208;
    61: op1_05_in19 = reg_0206;
    62: op1_05_in19 = reg_0560;
    63: op1_05_in19 = imem05_in[27:24];
    64: op1_05_in19 = reg_0405;
    65: op1_05_in19 = reg_0619;
    66: op1_05_in19 = reg_0154;
    67: op1_05_in19 = reg_0441;
    68: op1_05_in19 = reg_0541;
    69: op1_05_in19 = imem05_in[127:124];
    70: op1_05_in19 = reg_0253;
    71: op1_05_in19 = reg_0614;
    72: op1_05_in19 = imem06_in[51:48];
    73: op1_05_in19 = reg_0620;
    74: op1_05_in19 = reg_0183;
    96: op1_05_in19 = reg_0183;
    75: op1_05_in19 = imem01_in[71:68];
    76: op1_05_in19 = imem01_in[91:88];
    77: op1_05_in19 = reg_0656;
    78: op1_05_in19 = imem05_in[15:12];
    79: op1_05_in19 = reg_0766;
    80: op1_05_in19 = reg_0439;
    81: op1_05_in19 = reg_0777;
    82: op1_05_in19 = reg_0751;
    83: op1_05_in19 = imem01_in[99:96];
    84: op1_05_in19 = reg_0151;
    86: op1_05_in19 = reg_0509;
    87: op1_05_in19 = imem05_in[43:40];
    88: op1_05_in19 = reg_0244;
    89: op1_05_in19 = reg_0606;
    90: op1_05_in19 = reg_0270;
    91: op1_05_in19 = reg_0632;
    92: op1_05_in19 = reg_0202;
    93: op1_05_in19 = imem01_in[51:48];
    94: op1_05_in19 = reg_0761;
    95: op1_05_in19 = reg_0188;
    default: op1_05_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv19 = 1;
    8: op1_05_inv19 = 1;
    10: op1_05_inv19 = 1;
    13: op1_05_inv19 = 1;
    14: op1_05_inv19 = 1;
    15: op1_05_inv19 = 1;
    16: op1_05_inv19 = 1;
    18: op1_05_inv19 = 1;
    21: op1_05_inv19 = 1;
    23: op1_05_inv19 = 1;
    30: op1_05_inv19 = 1;
    31: op1_05_inv19 = 1;
    33: op1_05_inv19 = 1;
    39: op1_05_inv19 = 1;
    47: op1_05_inv19 = 1;
    48: op1_05_inv19 = 1;
    50: op1_05_inv19 = 1;
    52: op1_05_inv19 = 1;
    53: op1_05_inv19 = 1;
    54: op1_05_inv19 = 1;
    55: op1_05_inv19 = 1;
    56: op1_05_inv19 = 1;
    63: op1_05_inv19 = 1;
    66: op1_05_inv19 = 1;
    68: op1_05_inv19 = 1;
    71: op1_05_inv19 = 1;
    75: op1_05_inv19 = 1;
    76: op1_05_inv19 = 1;
    78: op1_05_inv19 = 1;
    79: op1_05_inv19 = 1;
    81: op1_05_inv19 = 1;
    84: op1_05_inv19 = 1;
    88: op1_05_inv19 = 1;
    92: op1_05_inv19 = 1;
    93: op1_05_inv19 = 1;
    94: op1_05_inv19 = 1;
    96: op1_05_inv19 = 1;
    default: op1_05_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in20 = reg_0487;
    5: op1_05_in20 = reg_0167;
    6: op1_05_in20 = reg_0571;
    7: op1_05_in20 = imem06_in[63:60];
    8: op1_05_in20 = imem01_in[91:88];
    9: op1_05_in20 = reg_0817;
    10: op1_05_in20 = reg_0733;
    12: op1_05_in20 = reg_0014;
    13: op1_05_in20 = imem06_in[39:36];
    14: op1_05_in20 = reg_0177;
    15: op1_05_in20 = reg_0098;
    16: op1_05_in20 = reg_0293;
    58: op1_05_in20 = reg_0293;
    17: op1_05_in20 = reg_0522;
    18: op1_05_in20 = reg_0780;
    19: op1_05_in20 = reg_0519;
    20: op1_05_in20 = imem05_in[19:16];
    21: op1_05_in20 = reg_0187;
    22: op1_05_in20 = imem01_in[39:36];
    46: op1_05_in20 = imem01_in[39:36];
    23: op1_05_in20 = reg_0723;
    24: op1_05_in20 = reg_0526;
    25: op1_05_in20 = reg_0289;
    26: op1_05_in20 = imem03_in[23:20];
    27: op1_05_in20 = reg_0808;
    28: op1_05_in20 = reg_0211;
    29: op1_05_in20 = imem01_in[99:96];
    30: op1_05_in20 = reg_0545;
    31: op1_05_in20 = imem06_in[95:92];
    32: op1_05_in20 = reg_0474;
    33: op1_05_in20 = reg_0535;
    35: op1_05_in20 = reg_0717;
    38: op1_05_in20 = imem01_in[7:4];
    39: op1_05_in20 = reg_0750;
    52: op1_05_in20 = reg_0750;
    40: op1_05_in20 = reg_0333;
    41: op1_05_in20 = imem06_in[23:20];
    43: op1_05_in20 = reg_0772;
    44: op1_05_in20 = reg_0560;
    45: op1_05_in20 = reg_0618;
    47: op1_05_in20 = imem03_in[39:36];
    48: op1_05_in20 = imem07_in[63:60];
    49: op1_05_in20 = reg_0255;
    50: op1_05_in20 = imem04_in[71:68];
    51: op1_05_in20 = reg_0563;
    53: op1_05_in20 = imem04_in[119:116];
    54: op1_05_in20 = reg_0269;
    55: op1_05_in20 = reg_0277;
    56: op1_05_in20 = imem07_in[107:104];
    59: op1_05_in20 = reg_0207;
    61: op1_05_in20 = reg_0192;
    62: op1_05_in20 = reg_0056;
    63: op1_05_in20 = imem05_in[67:64];
    64: op1_05_in20 = reg_0763;
    65: op1_05_in20 = reg_0404;
    66: op1_05_in20 = imem06_in[3:0];
    67: op1_05_in20 = reg_0446;
    68: op1_05_in20 = reg_0540;
    69: op1_05_in20 = reg_0231;
    70: op1_05_in20 = reg_0437;
    71: op1_05_in20 = reg_0774;
    72: op1_05_in20 = imem06_in[75:72];
    73: op1_05_in20 = reg_0787;
    75: op1_05_in20 = reg_0497;
    76: op1_05_in20 = imem01_in[103:100];
    83: op1_05_in20 = imem01_in[103:100];
    77: op1_05_in20 = reg_0703;
    78: op1_05_in20 = imem05_in[39:36];
    79: op1_05_in20 = reg_0265;
    80: op1_05_in20 = reg_0442;
    81: op1_05_in20 = reg_0651;
    82: op1_05_in20 = reg_0648;
    84: op1_05_in20 = imem06_in[115:112];
    86: op1_05_in20 = reg_0572;
    87: op1_05_in20 = imem05_in[47:44];
    88: op1_05_in20 = reg_0248;
    89: op1_05_in20 = reg_0619;
    90: op1_05_in20 = reg_0215;
    91: op1_05_in20 = imem07_in[11:8];
    92: op1_05_in20 = reg_0217;
    93: op1_05_in20 = imem01_in[63:60];
    94: op1_05_in20 = reg_0152;
    95: op1_05_in20 = reg_0505;
    96: op1_05_in20 = reg_0325;
    default: op1_05_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv20 = 1;
    7: op1_05_inv20 = 1;
    10: op1_05_inv20 = 1;
    12: op1_05_inv20 = 1;
    13: op1_05_inv20 = 1;
    14: op1_05_inv20 = 1;
    15: op1_05_inv20 = 1;
    17: op1_05_inv20 = 1;
    19: op1_05_inv20 = 1;
    21: op1_05_inv20 = 1;
    26: op1_05_inv20 = 1;
    28: op1_05_inv20 = 1;
    30: op1_05_inv20 = 1;
    31: op1_05_inv20 = 1;
    32: op1_05_inv20 = 1;
    41: op1_05_inv20 = 1;
    45: op1_05_inv20 = 1;
    47: op1_05_inv20 = 1;
    48: op1_05_inv20 = 1;
    51: op1_05_inv20 = 1;
    54: op1_05_inv20 = 1;
    55: op1_05_inv20 = 1;
    56: op1_05_inv20 = 1;
    59: op1_05_inv20 = 1;
    62: op1_05_inv20 = 1;
    64: op1_05_inv20 = 1;
    71: op1_05_inv20 = 1;
    72: op1_05_inv20 = 1;
    77: op1_05_inv20 = 1;
    78: op1_05_inv20 = 1;
    80: op1_05_inv20 = 1;
    81: op1_05_inv20 = 1;
    82: op1_05_inv20 = 1;
    83: op1_05_inv20 = 1;
    84: op1_05_inv20 = 1;
    86: op1_05_inv20 = 1;
    88: op1_05_inv20 = 1;
    91: op1_05_inv20 = 1;
    92: op1_05_inv20 = 1;
    94: op1_05_inv20 = 1;
    default: op1_05_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in21 = reg_0516;
    5: op1_05_in21 = reg_0182;
    6: op1_05_in21 = reg_0594;
    7: op1_05_in21 = imem06_in[79:76];
    8: op1_05_in21 = imem01_in[95:92];
    9: op1_05_in21 = reg_0037;
    10: op1_05_in21 = reg_0230;
    12: op1_05_in21 = reg_0805;
    13: op1_05_in21 = imem06_in[103:100];
    15: op1_05_in21 = reg_0077;
    16: op1_05_in21 = reg_0290;
    17: op1_05_in21 = reg_0514;
    18: op1_05_in21 = reg_0785;
    19: op1_05_in21 = reg_0507;
    20: op1_05_in21 = reg_0488;
    21: op1_05_in21 = reg_0213;
    22: op1_05_in21 = imem01_in[83:80];
    23: op1_05_in21 = reg_0729;
    24: op1_05_in21 = reg_0093;
    25: op1_05_in21 = reg_0071;
    26: op1_05_in21 = imem03_in[27:24];
    27: op1_05_in21 = reg_0014;
    28: op1_05_in21 = reg_0190;
    29: op1_05_in21 = imem01_in[119:116];
    30: op1_05_in21 = reg_0553;
    31: op1_05_in21 = imem07_in[23:20];
    32: op1_05_in21 = reg_0203;
    33: op1_05_in21 = reg_0756;
    35: op1_05_in21 = reg_0725;
    38: op1_05_in21 = imem01_in[43:40];
    39: op1_05_in21 = reg_0597;
    52: op1_05_in21 = reg_0597;
    40: op1_05_in21 = imem01_in[27:24];
    41: op1_05_in21 = imem06_in[63:60];
    43: op1_05_in21 = reg_0227;
    44: op1_05_in21 = reg_0429;
    45: op1_05_in21 = reg_0370;
    46: op1_05_in21 = imem01_in[47:44];
    47: op1_05_in21 = imem03_in[43:40];
    48: op1_05_in21 = imem07_in[75:72];
    49: op1_05_in21 = reg_0792;
    50: op1_05_in21 = imem04_in[75:72];
    51: op1_05_in21 = reg_0759;
    53: op1_05_in21 = reg_0059;
    54: op1_05_in21 = reg_0307;
    55: op1_05_in21 = reg_0149;
    56: op1_05_in21 = imem07_in[119:116];
    58: op1_05_in21 = reg_0242;
    79: op1_05_in21 = reg_0242;
    59: op1_05_in21 = reg_0196;
    61: op1_05_in21 = imem01_in[19:16];
    62: op1_05_in21 = reg_0303;
    63: op1_05_in21 = imem05_in[111:108];
    64: op1_05_in21 = reg_0270;
    65: op1_05_in21 = reg_0618;
    66: op1_05_in21 = reg_0291;
    67: op1_05_in21 = reg_0444;
    68: op1_05_in21 = reg_0535;
    69: op1_05_in21 = reg_0391;
    70: op1_05_in21 = reg_0435;
    71: op1_05_in21 = reg_0416;
    72: op1_05_in21 = imem06_in[123:120];
    73: op1_05_in21 = reg_0752;
    75: op1_05_in21 = reg_0388;
    76: op1_05_in21 = reg_0376;
    77: op1_05_in21 = reg_0548;
    78: op1_05_in21 = imem05_in[55:52];
    80: op1_05_in21 = reg_0437;
    81: op1_05_in21 = reg_0664;
    82: op1_05_in21 = reg_0571;
    83: op1_05_in21 = imem01_in[123:120];
    84: op1_05_in21 = reg_0289;
    86: op1_05_in21 = reg_0398;
    87: op1_05_in21 = imem05_in[51:48];
    88: op1_05_in21 = reg_0506;
    89: op1_05_in21 = reg_0354;
    90: op1_05_in21 = reg_0169;
    91: op1_05_in21 = imem07_in[19:16];
    92: op1_05_in21 = reg_0115;
    94: op1_05_in21 = reg_0115;
    93: op1_05_in21 = imem01_in[67:64];
    95: op1_05_in21 = imem01_in[35:32];
    96: op1_05_in21 = reg_0178;
    default: op1_05_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv21 = 1;
    6: op1_05_inv21 = 1;
    8: op1_05_inv21 = 1;
    17: op1_05_inv21 = 1;
    20: op1_05_inv21 = 1;
    23: op1_05_inv21 = 1;
    24: op1_05_inv21 = 1;
    25: op1_05_inv21 = 1;
    27: op1_05_inv21 = 1;
    28: op1_05_inv21 = 1;
    29: op1_05_inv21 = 1;
    30: op1_05_inv21 = 1;
    32: op1_05_inv21 = 1;
    33: op1_05_inv21 = 1;
    39: op1_05_inv21 = 1;
    40: op1_05_inv21 = 1;
    41: op1_05_inv21 = 1;
    43: op1_05_inv21 = 1;
    44: op1_05_inv21 = 1;
    48: op1_05_inv21 = 1;
    49: op1_05_inv21 = 1;
    58: op1_05_inv21 = 1;
    61: op1_05_inv21 = 1;
    68: op1_05_inv21 = 1;
    70: op1_05_inv21 = 1;
    71: op1_05_inv21 = 1;
    72: op1_05_inv21 = 1;
    75: op1_05_inv21 = 1;
    82: op1_05_inv21 = 1;
    88: op1_05_inv21 = 1;
    89: op1_05_inv21 = 1;
    90: op1_05_inv21 = 1;
    92: op1_05_inv21 = 1;
    93: op1_05_inv21 = 1;
    94: op1_05_inv21 = 1;
    default: op1_05_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in22 = reg_0505;
    88: op1_05_in22 = reg_0505;
    5: op1_05_in22 = reg_0160;
    6: op1_05_in22 = reg_0580;
    7: op1_05_in22 = reg_0606;
    8: op1_05_in22 = imem01_in[119:116];
    9: op1_05_in22 = reg_0029;
    10: op1_05_in22 = reg_0741;
    12: op1_05_in22 = imem04_in[55:52];
    13: op1_05_in22 = imem06_in[111:108];
    15: op1_05_in22 = reg_0079;
    44: op1_05_in22 = reg_0079;
    16: op1_05_in22 = reg_0296;
    17: op1_05_in22 = reg_0227;
    18: op1_05_in22 = reg_0784;
    19: op1_05_in22 = reg_0246;
    20: op1_05_in22 = reg_0788;
    21: op1_05_in22 = reg_0212;
    22: op1_05_in22 = imem01_in[95:92];
    23: op1_05_in22 = reg_0427;
    96: op1_05_in22 = reg_0427;
    24: op1_05_in22 = imem03_in[19:16];
    25: op1_05_in22 = imem05_in[11:8];
    26: op1_05_in22 = imem03_in[47:44];
    27: op1_05_in22 = reg_0802;
    28: op1_05_in22 = reg_0202;
    29: op1_05_in22 = reg_0519;
    30: op1_05_in22 = reg_0328;
    31: op1_05_in22 = imem07_in[39:36];
    32: op1_05_in22 = reg_0198;
    33: op1_05_in22 = reg_0740;
    35: op1_05_in22 = reg_0703;
    38: op1_05_in22 = imem01_in[71:68];
    39: op1_05_in22 = reg_0595;
    40: op1_05_in22 = imem01_in[55:52];
    41: op1_05_in22 = imem06_in[99:96];
    43: op1_05_in22 = reg_0760;
    45: op1_05_in22 = reg_0377;
    79: op1_05_in22 = reg_0377;
    46: op1_05_in22 = imem01_in[67:64];
    95: op1_05_in22 = imem01_in[67:64];
    47: op1_05_in22 = imem03_in[67:64];
    48: op1_05_in22 = imem07_in[83:80];
    49: op1_05_in22 = reg_0789;
    50: op1_05_in22 = imem04_in[95:92];
    51: op1_05_in22 = reg_0423;
    52: op1_05_in22 = reg_0751;
    53: op1_05_in22 = reg_0560;
    54: op1_05_in22 = reg_0148;
    55: op1_05_in22 = reg_0150;
    56: op1_05_in22 = imem07_in[123:120];
    58: op1_05_in22 = reg_0630;
    59: op1_05_in22 = imem01_in[3:0];
    61: op1_05_in22 = imem01_in[75:72];
    62: op1_05_in22 = reg_0052;
    63: op1_05_in22 = reg_0337;
    64: op1_05_in22 = reg_0375;
    65: op1_05_in22 = reg_0038;
    66: op1_05_in22 = reg_0624;
    67: op1_05_in22 = reg_0438;
    68: op1_05_in22 = reg_0756;
    69: op1_05_in22 = reg_0256;
    73: op1_05_in22 = reg_0256;
    70: op1_05_in22 = reg_0167;
    71: op1_05_in22 = imem05_in[39:36];
    72: op1_05_in22 = reg_0115;
    75: op1_05_in22 = reg_0397;
    76: op1_05_in22 = reg_0668;
    77: op1_05_in22 = reg_0705;
    78: op1_05_in22 = imem05_in[95:92];
    80: op1_05_in22 = reg_0448;
    81: op1_05_in22 = reg_0752;
    82: op1_05_in22 = reg_0568;
    83: op1_05_in22 = reg_0388;
    84: op1_05_in22 = reg_0299;
    86: op1_05_in22 = reg_0396;
    87: op1_05_in22 = imem05_in[75:72];
    89: op1_05_in22 = reg_0339;
    90: op1_05_in22 = reg_0242;
    91: op1_05_in22 = imem07_in[43:40];
    92: op1_05_in22 = reg_0225;
    93: op1_05_in22 = imem01_in[99:96];
    94: op1_05_in22 = reg_0234;
    default: op1_05_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_05_inv22 = 1;
    17: op1_05_inv22 = 1;
    19: op1_05_inv22 = 1;
    21: op1_05_inv22 = 1;
    23: op1_05_inv22 = 1;
    24: op1_05_inv22 = 1;
    25: op1_05_inv22 = 1;
    27: op1_05_inv22 = 1;
    29: op1_05_inv22 = 1;
    30: op1_05_inv22 = 1;
    31: op1_05_inv22 = 1;
    33: op1_05_inv22 = 1;
    38: op1_05_inv22 = 1;
    40: op1_05_inv22 = 1;
    43: op1_05_inv22 = 1;
    48: op1_05_inv22 = 1;
    49: op1_05_inv22 = 1;
    53: op1_05_inv22 = 1;
    55: op1_05_inv22 = 1;
    56: op1_05_inv22 = 1;
    58: op1_05_inv22 = 1;
    59: op1_05_inv22 = 1;
    61: op1_05_inv22 = 1;
    63: op1_05_inv22 = 1;
    65: op1_05_inv22 = 1;
    66: op1_05_inv22 = 1;
    67: op1_05_inv22 = 1;
    72: op1_05_inv22 = 1;
    75: op1_05_inv22 = 1;
    76: op1_05_inv22 = 1;
    79: op1_05_inv22 = 1;
    82: op1_05_inv22 = 1;
    84: op1_05_inv22 = 1;
    86: op1_05_inv22 = 1;
    93: op1_05_inv22 = 1;
    94: op1_05_inv22 = 1;
    default: op1_05_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in23 = reg_0235;
    43: op1_05_in23 = reg_0235;
    5: op1_05_in23 = reg_0168;
    6: op1_05_in23 = reg_0595;
    7: op1_05_in23 = reg_0402;
    8: op1_05_in23 = reg_0512;
    9: op1_05_in23 = reg_0038;
    10: op1_05_in23 = reg_0742;
    12: op1_05_in23 = imem04_in[59:56];
    13: op1_05_in23 = reg_0629;
    15: op1_05_in23 = imem03_in[35:32];
    16: op1_05_in23 = reg_0292;
    17: op1_05_in23 = reg_0776;
    18: op1_05_in23 = reg_0787;
    19: op1_05_in23 = reg_0218;
    20: op1_05_in23 = reg_0491;
    63: op1_05_in23 = reg_0491;
    21: op1_05_in23 = imem01_in[11:8];
    22: op1_05_in23 = reg_0523;
    23: op1_05_in23 = reg_0420;
    24: op1_05_in23 = imem03_in[47:44];
    25: op1_05_in23 = imem05_in[39:36];
    26: op1_05_in23 = imem03_in[83:80];
    27: op1_05_in23 = reg_0015;
    28: op1_05_in23 = imem01_in[63:60];
    29: op1_05_in23 = reg_0549;
    30: op1_05_in23 = reg_0542;
    53: op1_05_in23 = reg_0542;
    31: op1_05_in23 = imem07_in[43:40];
    32: op1_05_in23 = reg_0195;
    33: op1_05_in23 = imem03_in[59:56];
    35: op1_05_in23 = reg_0729;
    38: op1_05_in23 = imem01_in[79:76];
    39: op1_05_in23 = reg_0394;
    52: op1_05_in23 = reg_0394;
    40: op1_05_in23 = imem01_in[75:72];
    95: op1_05_in23 = imem01_in[75:72];
    41: op1_05_in23 = imem06_in[123:120];
    44: op1_05_in23 = reg_0433;
    62: op1_05_in23 = reg_0433;
    45: op1_05_in23 = reg_0405;
    46: op1_05_in23 = imem01_in[87:84];
    47: op1_05_in23 = imem03_in[99:96];
    48: op1_05_in23 = reg_0716;
    49: op1_05_in23 = reg_0493;
    50: op1_05_in23 = imem04_in[107:104];
    51: op1_05_in23 = reg_0054;
    54: op1_05_in23 = reg_0135;
    55: op1_05_in23 = reg_0151;
    56: op1_05_in23 = reg_0722;
    58: op1_05_in23 = reg_0270;
    59: op1_05_in23 = imem01_in[43:40];
    61: op1_05_in23 = imem01_in[91:88];
    64: op1_05_in23 = reg_0035;
    65: op1_05_in23 = reg_0242;
    66: op1_05_in23 = reg_0609;
    67: op1_05_in23 = reg_0182;
    68: op1_05_in23 = reg_0093;
    69: op1_05_in23 = reg_0550;
    70: op1_05_in23 = reg_0160;
    71: op1_05_in23 = imem05_in[67:64];
    72: op1_05_in23 = reg_0404;
    73: op1_05_in23 = imem07_in[51:48];
    75: op1_05_in23 = reg_0258;
    76: op1_05_in23 = reg_0772;
    77: op1_05_in23 = reg_0138;
    78: op1_05_in23 = imem05_in[99:96];
    79: op1_05_in23 = reg_0816;
    80: op1_05_in23 = reg_0435;
    81: op1_05_in23 = reg_0169;
    82: op1_05_in23 = reg_0572;
    83: op1_05_in23 = reg_0225;
    84: op1_05_in23 = reg_0291;
    86: op1_05_in23 = reg_0557;
    87: op1_05_in23 = imem05_in[87:84];
    88: op1_05_in23 = reg_0124;
    89: op1_05_in23 = reg_0265;
    90: op1_05_in23 = reg_0650;
    91: op1_05_in23 = imem07_in[47:44];
    92: op1_05_in23 = reg_0336;
    93: op1_05_in23 = imem01_in[107:104];
    94: op1_05_in23 = reg_0188;
    96: op1_05_in23 = reg_0184;
    default: op1_05_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv23 = 1;
    5: op1_05_inv23 = 1;
    6: op1_05_inv23 = 1;
    7: op1_05_inv23 = 1;
    8: op1_05_inv23 = 1;
    12: op1_05_inv23 = 1;
    19: op1_05_inv23 = 1;
    20: op1_05_inv23 = 1;
    21: op1_05_inv23 = 1;
    23: op1_05_inv23 = 1;
    27: op1_05_inv23 = 1;
    31: op1_05_inv23 = 1;
    32: op1_05_inv23 = 1;
    35: op1_05_inv23 = 1;
    38: op1_05_inv23 = 1;
    39: op1_05_inv23 = 1;
    40: op1_05_inv23 = 1;
    41: op1_05_inv23 = 1;
    44: op1_05_inv23 = 1;
    45: op1_05_inv23 = 1;
    46: op1_05_inv23 = 1;
    47: op1_05_inv23 = 1;
    48: op1_05_inv23 = 1;
    50: op1_05_inv23 = 1;
    51: op1_05_inv23 = 1;
    52: op1_05_inv23 = 1;
    53: op1_05_inv23 = 1;
    58: op1_05_inv23 = 1;
    63: op1_05_inv23 = 1;
    67: op1_05_inv23 = 1;
    75: op1_05_inv23 = 1;
    76: op1_05_inv23 = 1;
    77: op1_05_inv23 = 1;
    79: op1_05_inv23 = 1;
    81: op1_05_inv23 = 1;
    82: op1_05_inv23 = 1;
    89: op1_05_inv23 = 1;
    90: op1_05_inv23 = 1;
    93: op1_05_inv23 = 1;
    94: op1_05_inv23 = 1;
    default: op1_05_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in24 = reg_0227;
    5: op1_05_in24 = reg_0157;
    67: op1_05_in24 = reg_0157;
    6: op1_05_in24 = reg_0394;
    7: op1_05_in24 = reg_0356;
    8: op1_05_in24 = reg_0503;
    9: op1_05_in24 = imem07_in[3:0];
    10: op1_05_in24 = reg_0224;
    12: op1_05_in24 = imem04_in[111:108];
    13: op1_05_in24 = reg_0624;
    15: op1_05_in24 = imem03_in[55:52];
    16: op1_05_in24 = reg_0295;
    17: op1_05_in24 = reg_0507;
    18: op1_05_in24 = reg_0260;
    66: op1_05_in24 = reg_0260;
    89: op1_05_in24 = reg_0260;
    19: op1_05_in24 = reg_0502;
    20: op1_05_in24 = reg_0493;
    21: op1_05_in24 = imem01_in[35:32];
    22: op1_05_in24 = reg_0501;
    23: op1_05_in24 = reg_0175;
    24: op1_05_in24 = imem03_in[51:48];
    25: op1_05_in24 = imem05_in[67:64];
    26: op1_05_in24 = imem03_in[91:88];
    27: op1_05_in24 = reg_0016;
    28: op1_05_in24 = imem01_in[79:76];
    29: op1_05_in24 = reg_0759;
    30: op1_05_in24 = reg_0043;
    31: op1_05_in24 = imem07_in[63:60];
    32: op1_05_in24 = reg_0199;
    33: op1_05_in24 = imem03_in[79:76];
    35: op1_05_in24 = reg_0418;
    38: op1_05_in24 = imem01_in[87:84];
    39: op1_05_in24 = reg_0384;
    40: op1_05_in24 = reg_0100;
    41: op1_05_in24 = reg_0604;
    43: op1_05_in24 = reg_0425;
    44: op1_05_in24 = reg_0302;
    45: op1_05_in24 = reg_0776;
    46: op1_05_in24 = imem01_in[103:100];
    47: op1_05_in24 = imem03_in[107:104];
    48: op1_05_in24 = reg_0726;
    49: op1_05_in24 = reg_0793;
    63: op1_05_in24 = reg_0793;
    50: op1_05_in24 = imem04_in[115:112];
    51: op1_05_in24 = reg_0244;
    52: op1_05_in24 = reg_0395;
    53: op1_05_in24 = reg_0056;
    54: op1_05_in24 = reg_0128;
    55: op1_05_in24 = reg_0128;
    56: op1_05_in24 = reg_0719;
    58: op1_05_in24 = reg_0515;
    59: op1_05_in24 = imem01_in[55:52];
    61: op1_05_in24 = reg_0497;
    62: op1_05_in24 = reg_0631;
    64: op1_05_in24 = reg_0534;
    65: op1_05_in24 = reg_0748;
    68: op1_05_in24 = imem03_in[75:72];
    69: op1_05_in24 = reg_0489;
    70: op1_05_in24 = reg_0185;
    71: op1_05_in24 = imem05_in[91:88];
    72: op1_05_in24 = reg_0031;
    73: op1_05_in24 = imem07_in[79:76];
    75: op1_05_in24 = reg_0760;
    76: op1_05_in24 = reg_0741;
    77: op1_05_in24 = reg_0341;
    78: op1_05_in24 = reg_0827;
    79: op1_05_in24 = reg_0580;
    80: op1_05_in24 = reg_0268;
    81: op1_05_in24 = reg_0714;
    82: op1_05_in24 = reg_0372;
    83: op1_05_in24 = reg_0235;
    84: op1_05_in24 = reg_0618;
    86: op1_05_in24 = reg_0649;
    87: op1_05_in24 = reg_0337;
    88: op1_05_in24 = reg_0592;
    90: op1_05_in24 = imem07_in[15:12];
    91: op1_05_in24 = imem07_in[55:52];
    92: op1_05_in24 = reg_0102;
    93: op1_05_in24 = imem01_in[123:120];
    94: op1_05_in24 = reg_0243;
    95: op1_05_in24 = reg_0124;
    default: op1_05_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_05_inv24 = 1;
    10: op1_05_inv24 = 1;
    13: op1_05_inv24 = 1;
    20: op1_05_inv24 = 1;
    22: op1_05_inv24 = 1;
    23: op1_05_inv24 = 1;
    24: op1_05_inv24 = 1;
    26: op1_05_inv24 = 1;
    28: op1_05_inv24 = 1;
    29: op1_05_inv24 = 1;
    30: op1_05_inv24 = 1;
    31: op1_05_inv24 = 1;
    38: op1_05_inv24 = 1;
    43: op1_05_inv24 = 1;
    44: op1_05_inv24 = 1;
    46: op1_05_inv24 = 1;
    51: op1_05_inv24 = 1;
    53: op1_05_inv24 = 1;
    54: op1_05_inv24 = 1;
    55: op1_05_inv24 = 1;
    58: op1_05_inv24 = 1;
    63: op1_05_inv24 = 1;
    64: op1_05_inv24 = 1;
    68: op1_05_inv24 = 1;
    71: op1_05_inv24 = 1;
    72: op1_05_inv24 = 1;
    73: op1_05_inv24 = 1;
    76: op1_05_inv24 = 1;
    77: op1_05_inv24 = 1;
    78: op1_05_inv24 = 1;
    82: op1_05_inv24 = 1;
    83: op1_05_inv24 = 1;
    87: op1_05_inv24 = 1;
    89: op1_05_inv24 = 1;
    92: op1_05_inv24 = 1;
    94: op1_05_inv24 = 1;
    default: op1_05_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in25 = reg_0220;
    51: op1_05_in25 = reg_0220;
    6: op1_05_in25 = reg_0384;
    7: op1_05_in25 = reg_0405;
    72: op1_05_in25 = reg_0405;
    8: op1_05_in25 = reg_0506;
    9: op1_05_in25 = imem07_in[27:24];
    10: op1_05_in25 = reg_0743;
    12: op1_05_in25 = imem04_in[119:116];
    13: op1_05_in25 = reg_0618;
    15: op1_05_in25 = imem03_in[71:68];
    16: op1_05_in25 = reg_0307;
    17: op1_05_in25 = reg_0821;
    18: op1_05_in25 = reg_0149;
    19: op1_05_in25 = reg_0244;
    20: op1_05_in25 = reg_0787;
    21: op1_05_in25 = imem01_in[47:44];
    22: op1_05_in25 = reg_0497;
    23: op1_05_in25 = reg_0165;
    24: op1_05_in25 = imem03_in[55:52];
    25: op1_05_in25 = imem05_in[107:104];
    26: op1_05_in25 = imem03_in[115:112];
    27: op1_05_in25 = reg_0010;
    28: op1_05_in25 = imem01_in[107:104];
    59: op1_05_in25 = imem01_in[107:104];
    29: op1_05_in25 = reg_0233;
    30: op1_05_in25 = reg_0555;
    53: op1_05_in25 = reg_0555;
    31: op1_05_in25 = reg_0719;
    32: op1_05_in25 = reg_0197;
    33: op1_05_in25 = imem03_in[111:108];
    35: op1_05_in25 = reg_0434;
    38: op1_05_in25 = imem01_in[95:92];
    39: op1_05_in25 = reg_0575;
    40: op1_05_in25 = reg_0126;
    41: op1_05_in25 = reg_0291;
    43: op1_05_in25 = reg_0504;
    44: op1_05_in25 = reg_0297;
    45: op1_05_in25 = reg_0404;
    46: op1_05_in25 = imem01_in[111:108];
    47: op1_05_in25 = reg_0583;
    48: op1_05_in25 = reg_0717;
    49: op1_05_in25 = reg_0485;
    50: op1_05_in25 = reg_0542;
    52: op1_05_in25 = reg_0383;
    54: op1_05_in25 = reg_0152;
    55: op1_05_in25 = reg_0142;
    56: op1_05_in25 = reg_0729;
    58: op1_05_in25 = reg_0777;
    61: op1_05_in25 = reg_0653;
    62: op1_05_in25 = reg_0077;
    63: op1_05_in25 = reg_0113;
    64: op1_05_in25 = reg_0607;
    65: op1_05_in25 = reg_0638;
    66: op1_05_in25 = reg_0628;
    68: op1_05_in25 = imem03_in[87:84];
    69: op1_05_in25 = reg_0797;
    70: op1_05_in25 = reg_0176;
    71: op1_05_in25 = imem05_in[119:116];
    73: op1_05_in25 = imem07_in[119:116];
    75: op1_05_in25 = reg_0054;
    76: op1_05_in25 = reg_0645;
    77: op1_05_in25 = reg_0342;
    78: op1_05_in25 = reg_0825;
    79: op1_05_in25 = reg_0764;
    80: op1_05_in25 = imem07_in[31:28];
    90: op1_05_in25 = imem07_in[31:28];
    81: op1_05_in25 = reg_0161;
    82: op1_05_in25 = reg_0569;
    83: op1_05_in25 = reg_0421;
    84: op1_05_in25 = reg_0401;
    86: op1_05_in25 = reg_0000;
    87: op1_05_in25 = reg_0145;
    88: op1_05_in25 = reg_0119;
    89: op1_05_in25 = reg_0168;
    91: op1_05_in25 = imem07_in[67:64];
    92: op1_05_in25 = imem01_in[39:36];
    93: op1_05_in25 = reg_0376;
    94: op1_05_in25 = reg_0235;
    95: op1_05_in25 = reg_0111;
    default: op1_05_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv25 = 1;
    10: op1_05_inv25 = 1;
    12: op1_05_inv25 = 1;
    13: op1_05_inv25 = 1;
    15: op1_05_inv25 = 1;
    16: op1_05_inv25 = 1;
    17: op1_05_inv25 = 1;
    18: op1_05_inv25 = 1;
    19: op1_05_inv25 = 1;
    20: op1_05_inv25 = 1;
    21: op1_05_inv25 = 1;
    22: op1_05_inv25 = 1;
    23: op1_05_inv25 = 1;
    25: op1_05_inv25 = 1;
    29: op1_05_inv25 = 1;
    30: op1_05_inv25 = 1;
    31: op1_05_inv25 = 1;
    32: op1_05_inv25 = 1;
    33: op1_05_inv25 = 1;
    35: op1_05_inv25 = 1;
    39: op1_05_inv25 = 1;
    40: op1_05_inv25 = 1;
    49: op1_05_inv25 = 1;
    50: op1_05_inv25 = 1;
    51: op1_05_inv25 = 1;
    52: op1_05_inv25 = 1;
    53: op1_05_inv25 = 1;
    54: op1_05_inv25 = 1;
    56: op1_05_inv25 = 1;
    58: op1_05_inv25 = 1;
    61: op1_05_inv25 = 1;
    63: op1_05_inv25 = 1;
    64: op1_05_inv25 = 1;
    65: op1_05_inv25 = 1;
    66: op1_05_inv25 = 1;
    68: op1_05_inv25 = 1;
    70: op1_05_inv25 = 1;
    72: op1_05_inv25 = 1;
    75: op1_05_inv25 = 1;
    77: op1_05_inv25 = 1;
    78: op1_05_inv25 = 1;
    80: op1_05_inv25 = 1;
    81: op1_05_inv25 = 1;
    86: op1_05_inv25 = 1;
    87: op1_05_inv25 = 1;
    89: op1_05_inv25 = 1;
    91: op1_05_inv25 = 1;
    92: op1_05_inv25 = 1;
    94: op1_05_inv25 = 1;
    default: op1_05_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in26 = reg_0236;
    6: op1_05_in26 = reg_0388;
    7: op1_05_in26 = reg_0371;
    41: op1_05_in26 = reg_0371;
    8: op1_05_in26 = reg_0510;
    9: op1_05_in26 = imem07_in[31:28];
    10: op1_05_in26 = reg_0498;
    12: op1_05_in26 = reg_0530;
    13: op1_05_in26 = reg_0379;
    15: op1_05_in26 = imem03_in[107:104];
    68: op1_05_in26 = imem03_in[107:104];
    16: op1_05_in26 = reg_0078;
    17: op1_05_in26 = reg_0244;
    18: op1_05_in26 = reg_0154;
    54: op1_05_in26 = reg_0154;
    19: op1_05_in26 = reg_0216;
    20: op1_05_in26 = reg_0486;
    21: op1_05_in26 = imem01_in[95:92];
    22: op1_05_in26 = reg_0822;
    23: op1_05_in26 = reg_0166;
    24: op1_05_in26 = imem03_in[59:56];
    25: op1_05_in26 = imem05_in[127:124];
    26: op1_05_in26 = reg_0582;
    27: op1_05_in26 = imem04_in[43:40];
    28: op1_05_in26 = imem01_in[111:108];
    59: op1_05_in26 = imem01_in[111:108];
    29: op1_05_in26 = reg_0502;
    30: op1_05_in26 = reg_0280;
    31: op1_05_in26 = reg_0726;
    81: op1_05_in26 = reg_0726;
    32: op1_05_in26 = imem01_in[19:16];
    33: op1_05_in26 = imem03_in[123:120];
    35: op1_05_in26 = reg_0443;
    38: op1_05_in26 = imem01_in[103:100];
    39: op1_05_in26 = reg_0398;
    40: op1_05_in26 = imem02_in[59:56];
    43: op1_05_in26 = reg_0505;
    75: op1_05_in26 = reg_0505;
    44: op1_05_in26 = reg_0050;
    45: op1_05_in26 = reg_0242;
    46: op1_05_in26 = reg_0497;
    47: op1_05_in26 = reg_0597;
    48: op1_05_in26 = reg_0725;
    49: op1_05_in26 = reg_0787;
    50: op1_05_in26 = reg_0537;
    51: op1_05_in26 = reg_0425;
    52: op1_05_in26 = reg_0572;
    53: op1_05_in26 = reg_0060;
    55: op1_05_in26 = reg_0140;
    56: op1_05_in26 = reg_0715;
    58: op1_05_in26 = reg_0368;
    61: op1_05_in26 = reg_0668;
    62: op1_05_in26 = reg_0071;
    63: op1_05_in26 = reg_0278;
    64: op1_05_in26 = reg_0794;
    65: op1_05_in26 = reg_0593;
    66: op1_05_in26 = reg_0578;
    69: op1_05_in26 = reg_0229;
    70: op1_05_in26 = reg_0171;
    71: op1_05_in26 = reg_0550;
    72: op1_05_in26 = reg_0620;
    73: op1_05_in26 = reg_0730;
    76: op1_05_in26 = reg_0224;
    77: op1_05_in26 = reg_0414;
    78: op1_05_in26 = reg_0829;
    79: op1_05_in26 = reg_0576;
    80: op1_05_in26 = imem07_in[43:40];
    82: op1_05_in26 = reg_0747;
    83: op1_05_in26 = reg_0511;
    84: op1_05_in26 = reg_0260;
    86: op1_05_in26 = reg_0012;
    87: op1_05_in26 = reg_0538;
    88: op1_05_in26 = reg_0669;
    89: op1_05_in26 = reg_0405;
    90: op1_05_in26 = imem07_in[39:36];
    91: op1_05_in26 = imem07_in[75:72];
    92: op1_05_in26 = imem01_in[63:60];
    93: op1_05_in26 = reg_0085;
    94: op1_05_in26 = reg_0013;
    95: op1_05_in26 = reg_0007;
    default: op1_05_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_05_inv26 = 1;
    8: op1_05_inv26 = 1;
    9: op1_05_inv26 = 1;
    10: op1_05_inv26 = 1;
    13: op1_05_inv26 = 1;
    15: op1_05_inv26 = 1;
    16: op1_05_inv26 = 1;
    17: op1_05_inv26 = 1;
    19: op1_05_inv26 = 1;
    20: op1_05_inv26 = 1;
    21: op1_05_inv26 = 1;
    22: op1_05_inv26 = 1;
    24: op1_05_inv26 = 1;
    26: op1_05_inv26 = 1;
    28: op1_05_inv26 = 1;
    31: op1_05_inv26 = 1;
    32: op1_05_inv26 = 1;
    33: op1_05_inv26 = 1;
    35: op1_05_inv26 = 1;
    39: op1_05_inv26 = 1;
    41: op1_05_inv26 = 1;
    43: op1_05_inv26 = 1;
    47: op1_05_inv26 = 1;
    48: op1_05_inv26 = 1;
    51: op1_05_inv26 = 1;
    52: op1_05_inv26 = 1;
    58: op1_05_inv26 = 1;
    59: op1_05_inv26 = 1;
    61: op1_05_inv26 = 1;
    65: op1_05_inv26 = 1;
    68: op1_05_inv26 = 1;
    70: op1_05_inv26 = 1;
    71: op1_05_inv26 = 1;
    77: op1_05_inv26 = 1;
    78: op1_05_inv26 = 1;
    79: op1_05_inv26 = 1;
    80: op1_05_inv26 = 1;
    81: op1_05_inv26 = 1;
    84: op1_05_inv26 = 1;
    90: op1_05_inv26 = 1;
    92: op1_05_inv26 = 1;
    95: op1_05_inv26 = 1;
    default: op1_05_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in27 = reg_0237;
    6: op1_05_in27 = reg_0323;
    7: op1_05_in27 = reg_0375;
    8: op1_05_in27 = reg_0507;
    9: op1_05_in27 = imem07_in[39:36];
    10: op1_05_in27 = reg_0735;
    12: op1_05_in27 = reg_0542;
    13: op1_05_in27 = reg_0351;
    15: op1_05_in27 = reg_0602;
    16: op1_05_in27 = reg_0062;
    17: op1_05_in27 = reg_0123;
    18: op1_05_in27 = reg_0138;
    19: op1_05_in27 = reg_0503;
    20: op1_05_in27 = reg_0090;
    21: op1_05_in27 = imem01_in[115:112];
    22: op1_05_in27 = reg_0229;
    23: op1_05_in27 = reg_0177;
    24: op1_05_in27 = imem03_in[127:124];
    25: op1_05_in27 = reg_0785;
    26: op1_05_in27 = reg_0571;
    27: op1_05_in27 = imem04_in[51:48];
    28: op1_05_in27 = reg_0501;
    29: op1_05_in27 = reg_0245;
    30: op1_05_in27 = reg_0052;
    31: op1_05_in27 = reg_0715;
    32: op1_05_in27 = imem01_in[43:40];
    33: op1_05_in27 = reg_0565;
    35: op1_05_in27 = reg_0420;
    38: op1_05_in27 = reg_0822;
    39: op1_05_in27 = reg_0376;
    52: op1_05_in27 = reg_0376;
    40: op1_05_in27 = imem02_in[79:76];
    41: op1_05_in27 = reg_0298;
    43: op1_05_in27 = reg_0122;
    44: op1_05_in27 = reg_0078;
    45: op1_05_in27 = reg_0621;
    46: op1_05_in27 = reg_0825;
    47: op1_05_in27 = reg_0562;
    48: op1_05_in27 = reg_0709;
    49: op1_05_in27 = imem05_in[47:44];
    50: op1_05_in27 = reg_0088;
    51: op1_05_in27 = reg_0505;
    53: op1_05_in27 = reg_0057;
    54: op1_05_in27 = imem06_in[3:0];
    78: op1_05_in27 = imem06_in[3:0];
    55: op1_05_in27 = imem06_in[71:68];
    56: op1_05_in27 = reg_0253;
    58: op1_05_in27 = imem07_in[7:4];
    59: op1_05_in27 = imem01_in[119:116];
    61: op1_05_in27 = reg_0820;
    62: op1_05_in27 = reg_0074;
    63: op1_05_in27 = reg_0790;
    64: op1_05_in27 = reg_0656;
    65: op1_05_in27 = reg_0812;
    66: op1_05_in27 = reg_0638;
    68: op1_05_in27 = reg_0493;
    69: op1_05_in27 = reg_0307;
    71: op1_05_in27 = reg_0782;
    72: op1_05_in27 = reg_0651;
    73: op1_05_in27 = reg_0726;
    75: op1_05_in27 = reg_0124;
    76: op1_05_in27 = reg_0131;
    77: op1_05_in27 = reg_0590;
    79: op1_05_in27 = imem07_in[51:48];
    80: op1_05_in27 = imem07_in[67:64];
    81: op1_05_in27 = reg_0711;
    82: op1_05_in27 = reg_0007;
    83: op1_05_in27 = reg_0054;
    84: op1_05_in27 = reg_0613;
    86: op1_05_in27 = reg_0801;
    87: op1_05_in27 = reg_0751;
    88: op1_05_in27 = imem02_in[3:0];
    89: op1_05_in27 = reg_0484;
    90: op1_05_in27 = reg_0159;
    91: op1_05_in27 = imem07_in[83:80];
    92: op1_05_in27 = imem01_in[111:108];
    93: op1_05_in27 = reg_0111;
    94: op1_05_in27 = reg_0778;
    95: op1_05_in27 = reg_0101;
    default: op1_05_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv27 = 1;
    6: op1_05_inv27 = 1;
    7: op1_05_inv27 = 1;
    8: op1_05_inv27 = 1;
    15: op1_05_inv27 = 1;
    16: op1_05_inv27 = 1;
    17: op1_05_inv27 = 1;
    22: op1_05_inv27 = 1;
    25: op1_05_inv27 = 1;
    26: op1_05_inv27 = 1;
    27: op1_05_inv27 = 1;
    28: op1_05_inv27 = 1;
    29: op1_05_inv27 = 1;
    32: op1_05_inv27 = 1;
    33: op1_05_inv27 = 1;
    38: op1_05_inv27 = 1;
    40: op1_05_inv27 = 1;
    44: op1_05_inv27 = 1;
    45: op1_05_inv27 = 1;
    46: op1_05_inv27 = 1;
    48: op1_05_inv27 = 1;
    50: op1_05_inv27 = 1;
    52: op1_05_inv27 = 1;
    53: op1_05_inv27 = 1;
    54: op1_05_inv27 = 1;
    56: op1_05_inv27 = 1;
    59: op1_05_inv27 = 1;
    64: op1_05_inv27 = 1;
    76: op1_05_inv27 = 1;
    78: op1_05_inv27 = 1;
    81: op1_05_inv27 = 1;
    86: op1_05_inv27 = 1;
    90: op1_05_inv27 = 1;
    91: op1_05_inv27 = 1;
    92: op1_05_inv27 = 1;
    94: op1_05_inv27 = 1;
    default: op1_05_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in28 = reg_0238;
    6: op1_05_in28 = reg_0312;
    7: op1_05_in28 = reg_0383;
    8: op1_05_in28 = reg_0505;
    9: op1_05_in28 = imem07_in[59:56];
    79: op1_05_in28 = imem07_in[59:56];
    10: op1_05_in28 = imem01_in[115:112];
    12: op1_05_in28 = reg_0529;
    13: op1_05_in28 = reg_0337;
    15: op1_05_in28 = reg_0573;
    26: op1_05_in28 = reg_0573;
    16: op1_05_in28 = reg_0065;
    17: op1_05_in28 = imem02_in[19:16];
    18: op1_05_in28 = reg_0129;
    19: op1_05_in28 = reg_0234;
    20: op1_05_in28 = reg_0304;
    82: op1_05_in28 = reg_0304;
    21: op1_05_in28 = reg_0229;
    22: op1_05_in28 = reg_0514;
    23: op1_05_in28 = reg_0158;
    24: op1_05_in28 = reg_0582;
    25: op1_05_in28 = reg_0495;
    27: op1_05_in28 = imem04_in[71:68];
    28: op1_05_in28 = reg_0772;
    29: op1_05_in28 = reg_0243;
    30: op1_05_in28 = reg_0290;
    31: op1_05_in28 = reg_0707;
    48: op1_05_in28 = reg_0707;
    32: op1_05_in28 = imem01_in[59:56];
    33: op1_05_in28 = reg_0581;
    35: op1_05_in28 = reg_0431;
    38: op1_05_in28 = reg_0487;
    39: op1_05_in28 = reg_0396;
    40: op1_05_in28 = reg_0642;
    41: op1_05_in28 = reg_0215;
    43: op1_05_in28 = imem02_in[31:28];
    44: op1_05_in28 = reg_0066;
    45: op1_05_in28 = reg_0623;
    46: op1_05_in28 = reg_0759;
    47: op1_05_in28 = reg_0013;
    49: op1_05_in28 = imem05_in[67:64];
    50: op1_05_in28 = reg_0060;
    51: op1_05_in28 = reg_0122;
    52: op1_05_in28 = reg_0000;
    53: op1_05_in28 = reg_0516;
    54: op1_05_in28 = imem06_in[27:24];
    55: op1_05_in28 = reg_0299;
    56: op1_05_in28 = reg_0635;
    58: op1_05_in28 = imem07_in[11:8];
    59: op1_05_in28 = reg_0497;
    61: op1_05_in28 = reg_0563;
    62: op1_05_in28 = reg_0508;
    63: op1_05_in28 = reg_0742;
    64: op1_05_in28 = reg_0496;
    65: op1_05_in28 = reg_0368;
    66: op1_05_in28 = reg_0593;
    68: op1_05_in28 = reg_0588;
    69: op1_05_in28 = reg_0147;
    71: op1_05_in28 = reg_0489;
    72: op1_05_in28 = reg_0819;
    73: op1_05_in28 = reg_0718;
    75: op1_05_in28 = reg_0672;
    76: op1_05_in28 = reg_0101;
    77: op1_05_in28 = reg_0092;
    78: op1_05_in28 = imem06_in[7:4];
    80: op1_05_in28 = imem07_in[107:104];
    81: op1_05_in28 = reg_0731;
    83: op1_05_in28 = reg_0217;
    84: op1_05_in28 = reg_0659;
    86: op1_05_in28 = imem04_in[11:8];
    87: op1_05_in28 = reg_0285;
    88: op1_05_in28 = imem02_in[27:24];
    89: op1_05_in28 = reg_0750;
    90: op1_05_in28 = reg_0166;
    91: op1_05_in28 = imem07_in[119:116];
    92: op1_05_in28 = imem01_in[119:116];
    93: op1_05_in28 = reg_0511;
    94: op1_05_in28 = reg_0324;
    95: op1_05_in28 = reg_0425;
    default: op1_05_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_05_inv28 = 1;
    7: op1_05_inv28 = 1;
    8: op1_05_inv28 = 1;
    9: op1_05_inv28 = 1;
    12: op1_05_inv28 = 1;
    13: op1_05_inv28 = 1;
    15: op1_05_inv28 = 1;
    17: op1_05_inv28 = 1;
    18: op1_05_inv28 = 1;
    19: op1_05_inv28 = 1;
    20: op1_05_inv28 = 1;
    22: op1_05_inv28 = 1;
    24: op1_05_inv28 = 1;
    26: op1_05_inv28 = 1;
    29: op1_05_inv28 = 1;
    30: op1_05_inv28 = 1;
    32: op1_05_inv28 = 1;
    43: op1_05_inv28 = 1;
    44: op1_05_inv28 = 1;
    45: op1_05_inv28 = 1;
    46: op1_05_inv28 = 1;
    47: op1_05_inv28 = 1;
    49: op1_05_inv28 = 1;
    53: op1_05_inv28 = 1;
    55: op1_05_inv28 = 1;
    56: op1_05_inv28 = 1;
    59: op1_05_inv28 = 1;
    62: op1_05_inv28 = 1;
    63: op1_05_inv28 = 1;
    69: op1_05_inv28 = 1;
    72: op1_05_inv28 = 1;
    75: op1_05_inv28 = 1;
    78: op1_05_inv28 = 1;
    79: op1_05_inv28 = 1;
    80: op1_05_inv28 = 1;
    81: op1_05_inv28 = 1;
    82: op1_05_inv28 = 1;
    83: op1_05_inv28 = 1;
    86: op1_05_inv28 = 1;
    89: op1_05_inv28 = 1;
    92: op1_05_inv28 = 1;
    93: op1_05_inv28 = 1;
    default: op1_05_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in29 = reg_0119;
    6: op1_05_in29 = reg_0393;
    7: op1_05_in29 = reg_0404;
    8: op1_05_in29 = reg_0238;
    9: op1_05_in29 = imem07_in[83:80];
    10: op1_05_in29 = reg_0241;
    12: op1_05_in29 = reg_0539;
    13: op1_05_in29 = reg_0812;
    15: op1_05_in29 = reg_0568;
    16: op1_05_in29 = reg_0067;
    17: op1_05_in29 = imem02_in[35:32];
    18: op1_05_in29 = reg_0134;
    19: op1_05_in29 = reg_0508;
    20: op1_05_in29 = reg_0742;
    21: op1_05_in29 = reg_0517;
    71: op1_05_in29 = reg_0517;
    22: op1_05_in29 = reg_0776;
    23: op1_05_in29 = reg_0173;
    24: op1_05_in29 = reg_0571;
    25: op1_05_in29 = reg_0786;
    26: op1_05_in29 = reg_0583;
    27: op1_05_in29 = imem04_in[95:92];
    28: op1_05_in29 = reg_0232;
    29: op1_05_in29 = reg_0249;
    30: op1_05_in29 = reg_0284;
    31: op1_05_in29 = reg_0434;
    32: op1_05_in29 = reg_0772;
    33: op1_05_in29 = reg_0595;
    35: op1_05_in29 = reg_0162;
    38: op1_05_in29 = reg_0235;
    39: op1_05_in29 = reg_0389;
    40: op1_05_in29 = reg_0653;
    59: op1_05_in29 = reg_0653;
    41: op1_05_in29 = reg_0406;
    43: op1_05_in29 = imem02_in[43:40];
    44: op1_05_in29 = reg_0255;
    45: op1_05_in29 = imem07_in[23:20];
    46: op1_05_in29 = reg_0771;
    47: op1_05_in29 = reg_0004;
    48: op1_05_in29 = reg_0441;
    49: op1_05_in29 = reg_0147;
    50: op1_05_in29 = reg_0057;
    51: op1_05_in29 = reg_0124;
    52: op1_05_in29 = reg_0019;
    53: op1_05_in29 = reg_0432;
    54: op1_05_in29 = imem06_in[47:44];
    55: op1_05_in29 = reg_0291;
    56: op1_05_in29 = reg_0438;
    58: op1_05_in29 = imem07_in[15:12];
    61: op1_05_in29 = reg_0237;
    62: op1_05_in29 = imem05_in[7:4];
    63: op1_05_in29 = reg_0258;
    64: op1_05_in29 = reg_0495;
    65: op1_05_in29 = reg_0767;
    66: op1_05_in29 = reg_0512;
    68: op1_05_in29 = reg_0384;
    69: op1_05_in29 = reg_0148;
    72: op1_05_in29 = reg_0501;
    73: op1_05_in29 = reg_0727;
    75: op1_05_in29 = reg_0677;
    76: op1_05_in29 = reg_0054;
    77: op1_05_in29 = reg_0081;
    78: op1_05_in29 = imem06_in[55:52];
    79: op1_05_in29 = imem07_in[103:100];
    80: op1_05_in29 = imem07_in[115:112];
    81: op1_05_in29 = reg_0253;
    82: op1_05_in29 = reg_0560;
    83: op1_05_in29 = reg_0567;
    84: op1_05_in29 = reg_0654;
    86: op1_05_in29 = imem04_in[23:20];
    87: op1_05_in29 = reg_0152;
    88: op1_05_in29 = imem02_in[87:84];
    89: op1_05_in29 = reg_0593;
    90: op1_05_in29 = reg_0164;
    91: op1_05_in29 = imem07_in[127:124];
    92: op1_05_in29 = imem01_in[127:124];
    93: op1_05_in29 = reg_0051;
    94: op1_05_in29 = reg_0510;
    95: op1_05_in29 = reg_0504;
    default: op1_05_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_05_inv29 = 1;
    7: op1_05_inv29 = 1;
    12: op1_05_inv29 = 1;
    16: op1_05_inv29 = 1;
    17: op1_05_inv29 = 1;
    19: op1_05_inv29 = 1;
    20: op1_05_inv29 = 1;
    21: op1_05_inv29 = 1;
    22: op1_05_inv29 = 1;
    23: op1_05_inv29 = 1;
    24: op1_05_inv29 = 1;
    25: op1_05_inv29 = 1;
    26: op1_05_inv29 = 1;
    32: op1_05_inv29 = 1;
    39: op1_05_inv29 = 1;
    40: op1_05_inv29 = 1;
    43: op1_05_inv29 = 1;
    49: op1_05_inv29 = 1;
    50: op1_05_inv29 = 1;
    58: op1_05_inv29 = 1;
    59: op1_05_inv29 = 1;
    61: op1_05_inv29 = 1;
    62: op1_05_inv29 = 1;
    66: op1_05_inv29 = 1;
    68: op1_05_inv29 = 1;
    69: op1_05_inv29 = 1;
    71: op1_05_inv29 = 1;
    72: op1_05_inv29 = 1;
    75: op1_05_inv29 = 1;
    78: op1_05_inv29 = 1;
    80: op1_05_inv29 = 1;
    83: op1_05_inv29 = 1;
    84: op1_05_inv29 = 1;
    87: op1_05_inv29 = 1;
    88: op1_05_inv29 = 1;
    89: op1_05_inv29 = 1;
    90: op1_05_inv29 = 1;
    91: op1_05_inv29 = 1;
    94: op1_05_inv29 = 1;
    default: op1_05_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_05_in30 = reg_0120;
    8: op1_05_in30 = reg_0120;
    6: op1_05_in30 = reg_0389;
    7: op1_05_in30 = reg_0337;
    9: op1_05_in30 = reg_0719;
    10: op1_05_in30 = reg_0511;
    12: op1_05_in30 = reg_0281;
    13: op1_05_in30 = reg_0819;
    15: op1_05_in30 = reg_0584;
    16: op1_05_in30 = reg_0068;
    17: op1_05_in30 = imem02_in[67:64];
    18: op1_05_in30 = imem06_in[15:12];
    19: op1_05_in30 = reg_0103;
    20: op1_05_in30 = reg_0282;
    21: op1_05_in30 = reg_0776;
    22: op1_05_in30 = reg_0755;
    68: op1_05_in30 = reg_0755;
    24: op1_05_in30 = reg_0599;
    25: op1_05_in30 = reg_0304;
    26: op1_05_in30 = reg_0568;
    27: op1_05_in30 = imem04_in[127:124];
    28: op1_05_in30 = reg_0505;
    38: op1_05_in30 = reg_0505;
    29: op1_05_in30 = reg_0127;
    30: op1_05_in30 = reg_0062;
    31: op1_05_in30 = reg_0435;
    32: op1_05_in30 = reg_0520;
    33: op1_05_in30 = reg_0384;
    35: op1_05_in30 = reg_0173;
    39: op1_05_in30 = reg_0000;
    40: op1_05_in30 = reg_0646;
    41: op1_05_in30 = reg_0028;
    43: op1_05_in30 = imem02_in[71:68];
    44: op1_05_in30 = imem05_in[3:0];
    45: op1_05_in30 = imem07_in[63:60];
    46: op1_05_in30 = reg_0761;
    47: op1_05_in30 = imem04_in[51:48];
    48: op1_05_in30 = reg_0064;
    49: op1_05_in30 = reg_0145;
    69: op1_05_in30 = reg_0145;
    50: op1_05_in30 = reg_0551;
    51: op1_05_in30 = reg_0125;
    52: op1_05_in30 = reg_0002;
    53: op1_05_in30 = reg_0079;
    54: op1_05_in30 = imem06_in[79:76];
    55: op1_05_in30 = reg_0624;
    56: op1_05_in30 = reg_0268;
    58: op1_05_in30 = imem07_in[19:16];
    59: op1_05_in30 = reg_0772;
    61: op1_05_in30 = reg_0232;
    62: op1_05_in30 = imem05_in[59:56];
    63: op1_05_in30 = reg_0249;
    64: op1_05_in30 = imem07_in[47:44];
    65: op1_05_in30 = reg_0752;
    72: op1_05_in30 = reg_0752;
    66: op1_05_in30 = reg_0032;
    71: op1_05_in30 = reg_0326;
    73: op1_05_in30 = reg_0439;
    75: op1_05_in30 = reg_0678;
    76: op1_05_in30 = reg_0567;
    77: op1_05_in30 = reg_0535;
    78: op1_05_in30 = imem06_in[87:84];
    79: op1_05_in30 = reg_0716;
    81: op1_05_in30 = reg_0053;
    82: op1_05_in30 = reg_0080;
    83: op1_05_in30 = reg_0240;
    84: op1_05_in30 = reg_0583;
    86: op1_05_in30 = imem04_in[43:40];
    87: op1_05_in30 = reg_0143;
    88: op1_05_in30 = imem02_in[115:112];
    89: op1_05_in30 = reg_0335;
    90: op1_05_in30 = reg_0789;
    91: op1_05_in30 = reg_0160;
    92: op1_05_in30 = reg_0105;
    93: op1_05_in30 = reg_0220;
    94: op1_05_in30 = reg_0225;
    95: op1_05_in30 = reg_0420;
    default: op1_05_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_05_inv30 = 1;
    15: op1_05_inv30 = 1;
    17: op1_05_inv30 = 1;
    19: op1_05_inv30 = 1;
    20: op1_05_inv30 = 1;
    22: op1_05_inv30 = 1;
    24: op1_05_inv30 = 1;
    25: op1_05_inv30 = 1;
    26: op1_05_inv30 = 1;
    28: op1_05_inv30 = 1;
    29: op1_05_inv30 = 1;
    30: op1_05_inv30 = 1;
    32: op1_05_inv30 = 1;
    35: op1_05_inv30 = 1;
    41: op1_05_inv30 = 1;
    43: op1_05_inv30 = 1;
    44: op1_05_inv30 = 1;
    47: op1_05_inv30 = 1;
    48: op1_05_inv30 = 1;
    50: op1_05_inv30 = 1;
    51: op1_05_inv30 = 1;
    52: op1_05_inv30 = 1;
    54: op1_05_inv30 = 1;
    58: op1_05_inv30 = 1;
    61: op1_05_inv30 = 1;
    62: op1_05_inv30 = 1;
    66: op1_05_inv30 = 1;
    68: op1_05_inv30 = 1;
    69: op1_05_inv30 = 1;
    71: op1_05_inv30 = 1;
    73: op1_05_inv30 = 1;
    76: op1_05_inv30 = 1;
    79: op1_05_inv30 = 1;
    82: op1_05_inv30 = 1;
    86: op1_05_inv30 = 1;
    89: op1_05_inv30 = 1;
    93: op1_05_inv30 = 1;
    94: op1_05_inv30 = 1;
    default: op1_05_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_05_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_05_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in00 = reg_0121;
    5: op1_06_in00 = imem00_in[55:52];
    6: op1_06_in00 = reg_0001;
    7: op1_06_in00 = reg_0033;
    8: op1_06_in00 = reg_0112;
    9: op1_06_in00 = imem00_in[3:0];
    36: op1_06_in00 = imem00_in[3:0];
    42: op1_06_in00 = imem00_in[3:0];
    10: op1_06_in00 = reg_0502;
    83: op1_06_in00 = reg_0502;
    11: op1_06_in00 = imem00_in[23:20];
    3: op1_06_in00 = imem07_in[23:20];
    65: op1_06_in00 = imem07_in[23:20];
    12: op1_06_in00 = reg_0283;
    13: op1_06_in00 = reg_0816;
    14: op1_06_in00 = imem00_in[35:32];
    15: op1_06_in00 = reg_0585;
    16: op1_06_in00 = reg_0071;
    17: op1_06_in00 = imem02_in[95:92];
    18: op1_06_in00 = imem06_in[19:16];
    2: op1_06_in00 = imem07_in[47:44];
    19: op1_06_in00 = reg_0119;
    51: op1_06_in00 = reg_0119;
    20: op1_06_in00 = reg_0269;
    21: op1_06_in00 = reg_0234;
    22: op1_06_in00 = reg_0821;
    23: op1_06_in00 = reg_0694;
    24: op1_06_in00 = reg_0578;
    1: op1_06_in00 = imem07_in[115:112];
    25: op1_06_in00 = reg_0309;
    26: op1_06_in00 = reg_0592;
    27: op1_06_in00 = reg_0556;
    28: op1_06_in00 = reg_0233;
    29: op1_06_in00 = imem02_in[7:4];
    30: op1_06_in00 = reg_0254;
    31: op1_06_in00 = imem00_in[7:4];
    34: op1_06_in00 = imem00_in[7:4];
    67: op1_06_in00 = imem00_in[7:4];
    85: op1_06_in00 = imem00_in[7:4];
    96: op1_06_in00 = imem00_in[7:4];
    32: op1_06_in00 = reg_0519;
    33: op1_06_in00 = reg_0575;
    35: op1_06_in00 = reg_0184;
    37: op1_06_in00 = imem00_in[11:8];
    38: op1_06_in00 = reg_0239;
    39: op1_06_in00 = reg_0002;
    40: op1_06_in00 = reg_0660;
    41: op1_06_in00 = reg_0753;
    43: op1_06_in00 = imem02_in[83:80];
    44: op1_06_in00 = imem05_in[51:48];
    45: op1_06_in00 = imem07_in[71:68];
    46: op1_06_in00 = reg_0507;
    47: op1_06_in00 = imem04_in[127:124];
    48: op1_06_in00 = reg_0439;
    49: op1_06_in00 = reg_0142;
    50: op1_06_in00 = reg_0547;
    52: op1_06_in00 = reg_0013;
    53: op1_06_in00 = reg_0052;
    54: op1_06_in00 = imem06_in[83:80];
    55: op1_06_in00 = reg_0605;
    56: op1_06_in00 = reg_0161;
    57: op1_06_in00 = imem00_in[15:12];
    58: op1_06_in00 = imem07_in[59:56];
    59: op1_06_in00 = reg_0496;
    60: op1_06_in00 = imem00_in[83:80];
    61: op1_06_in00 = reg_0243;
    62: op1_06_in00 = imem05_in[79:76];
    63: op1_06_in00 = reg_0732;
    64: op1_06_in00 = reg_0713;
    66: op1_06_in00 = reg_0620;
    68: op1_06_in00 = reg_0747;
    69: op1_06_in00 = reg_0143;
    70: op1_06_in00 = imem00_in[19:16];
    71: op1_06_in00 = reg_0147;
    72: op1_06_in00 = imem07_in[3:0];
    73: op1_06_in00 = reg_0434;
    74: op1_06_in00 = imem00_in[43:40];
    75: op1_06_in00 = imem02_in[23:20];
    76: op1_06_in00 = reg_0505;
    77: op1_06_in00 = reg_0539;
    78: op1_06_in00 = imem06_in[91:88];
    79: op1_06_in00 = reg_0160;
    80: op1_06_in00 = imem00_in[27:24];
    81: op1_06_in00 = reg_0333;
    82: op1_06_in00 = reg_0056;
    84: op1_06_in00 = reg_0638;
    86: op1_06_in00 = imem04_in[47:44];
    87: op1_06_in00 = reg_0761;
    88: op1_06_in00 = imem02_in[127:124];
    89: op1_06_in00 = reg_0612;
    90: op1_06_in00 = reg_0158;
    91: op1_06_in00 = reg_0164;
    92: op1_06_in00 = reg_0118;
    93: op1_06_in00 = reg_0101;
    94: op1_06_in00 = imem01_in[7:4];
    95: op1_06_in00 = reg_0122;
    default: op1_06_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv00 = 1;
    5: op1_06_inv00 = 1;
    6: op1_06_inv00 = 1;
    8: op1_06_inv00 = 1;
    10: op1_06_inv00 = 1;
    14: op1_06_inv00 = 1;
    16: op1_06_inv00 = 1;
    17: op1_06_inv00 = 1;
    20: op1_06_inv00 = 1;
    23: op1_06_inv00 = 1;
    1: op1_06_inv00 = 1;
    25: op1_06_inv00 = 1;
    27: op1_06_inv00 = 1;
    28: op1_06_inv00 = 1;
    30: op1_06_inv00 = 1;
    32: op1_06_inv00 = 1;
    34: op1_06_inv00 = 1;
    37: op1_06_inv00 = 1;
    38: op1_06_inv00 = 1;
    40: op1_06_inv00 = 1;
    41: op1_06_inv00 = 1;
    43: op1_06_inv00 = 1;
    45: op1_06_inv00 = 1;
    46: op1_06_inv00 = 1;
    48: op1_06_inv00 = 1;
    50: op1_06_inv00 = 1;
    51: op1_06_inv00 = 1;
    52: op1_06_inv00 = 1;
    53: op1_06_inv00 = 1;
    57: op1_06_inv00 = 1;
    58: op1_06_inv00 = 1;
    60: op1_06_inv00 = 1;
    62: op1_06_inv00 = 1;
    66: op1_06_inv00 = 1;
    67: op1_06_inv00 = 1;
    68: op1_06_inv00 = 1;
    71: op1_06_inv00 = 1;
    73: op1_06_inv00 = 1;
    74: op1_06_inv00 = 1;
    76: op1_06_inv00 = 1;
    77: op1_06_inv00 = 1;
    79: op1_06_inv00 = 1;
    80: op1_06_inv00 = 1;
    81: op1_06_inv00 = 1;
    86: op1_06_inv00 = 1;
    87: op1_06_inv00 = 1;
    88: op1_06_inv00 = 1;
    90: op1_06_inv00 = 1;
    93: op1_06_inv00 = 1;
    95: op1_06_inv00 = 1;
    96: op1_06_inv00 = 1;
    default: op1_06_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in01 = reg_0110;
    5: op1_06_in01 = imem00_in[75:72];
    6: op1_06_in01 = reg_0808;
    7: op1_06_in01 = reg_0028;
    8: op1_06_in01 = reg_0113;
    9: op1_06_in01 = imem00_in[23:20];
    34: op1_06_in01 = imem00_in[23:20];
    70: op1_06_in01 = imem00_in[23:20];
    10: op1_06_in01 = reg_0244;
    11: op1_06_in01 = imem00_in[43:40];
    96: op1_06_in01 = imem00_in[43:40];
    3: op1_06_in01 = imem07_in[39:36];
    12: op1_06_in01 = reg_0300;
    13: op1_06_in01 = reg_0036;
    14: op1_06_in01 = imem00_in[39:36];
    42: op1_06_in01 = imem00_in[39:36];
    15: op1_06_in01 = reg_0600;
    16: op1_06_in01 = imem05_in[3:0];
    17: op1_06_in01 = reg_0653;
    18: op1_06_in01 = imem06_in[43:40];
    2: op1_06_in01 = imem07_in[71:68];
    19: op1_06_in01 = reg_0112;
    20: op1_06_in01 = reg_0084;
    21: op1_06_in01 = reg_0504;
    22: op1_06_in01 = reg_0217;
    23: op1_06_in01 = reg_0676;
    24: op1_06_in01 = reg_0597;
    25: op1_06_in01 = reg_0742;
    26: op1_06_in01 = reg_0589;
    27: op1_06_in01 = reg_0547;
    28: op1_06_in01 = reg_0245;
    29: op1_06_in01 = imem02_in[67:64];
    30: op1_06_in01 = reg_0069;
    31: op1_06_in01 = imem00_in[31:28];
    57: op1_06_in01 = imem00_in[31:28];
    32: op1_06_in01 = reg_0563;
    33: op1_06_in01 = reg_0568;
    36: op1_06_in01 = imem00_in[55:52];
    37: op1_06_in01 = imem00_in[59:56];
    38: op1_06_in01 = reg_0220;
    39: op1_06_in01 = reg_0003;
    40: op1_06_in01 = reg_0639;
    41: op1_06_in01 = reg_0372;
    43: op1_06_in01 = imem02_in[87:84];
    44: op1_06_in01 = imem05_in[63:60];
    45: op1_06_in01 = imem07_in[99:96];
    46: op1_06_in01 = reg_0421;
    47: op1_06_in01 = reg_0055;
    48: op1_06_in01 = reg_0180;
    49: op1_06_in01 = reg_0140;
    50: op1_06_in01 = reg_0305;
    51: op1_06_in01 = reg_0127;
    52: op1_06_in01 = reg_0007;
    53: op1_06_in01 = reg_0520;
    54: op1_06_in01 = imem06_in[99:96];
    55: op1_06_in01 = reg_0609;
    56: op1_06_in01 = reg_0167;
    58: op1_06_in01 = imem07_in[63:60];
    59: op1_06_in01 = reg_0778;
    60: op1_06_in01 = imem00_in[87:84];
    61: op1_06_in01 = reg_0118;
    95: op1_06_in01 = reg_0118;
    62: op1_06_in01 = imem05_in[111:108];
    63: op1_06_in01 = reg_0101;
    64: op1_06_in01 = reg_0707;
    65: op1_06_in01 = imem07_in[43:40];
    66: op1_06_in01 = reg_0794;
    67: op1_06_in01 = imem00_in[47:44];
    68: op1_06_in01 = reg_0396;
    69: op1_06_in01 = reg_0137;
    71: op1_06_in01 = reg_0149;
    72: op1_06_in01 = imem07_in[27:24];
    73: op1_06_in01 = reg_0440;
    74: op1_06_in01 = imem00_in[123:120];
    75: op1_06_in01 = imem02_in[99:96];
    76: op1_06_in01 = reg_0108;
    77: op1_06_in01 = reg_0756;
    78: op1_06_in01 = imem06_in[95:92];
    79: op1_06_in01 = reg_0103;
    80: op1_06_in01 = reg_0682;
    81: op1_06_in01 = reg_0449;
    82: op1_06_in01 = reg_0087;
    83: op1_06_in01 = reg_0294;
    84: op1_06_in01 = reg_0593;
    85: op1_06_in01 = imem00_in[11:8];
    86: op1_06_in01 = imem04_in[75:72];
    87: op1_06_in01 = reg_0765;
    88: op1_06_in01 = reg_0056;
    89: op1_06_in01 = reg_0777;
    90: op1_06_in01 = reg_0157;
    91: op1_06_in01 = reg_0709;
    92: op1_06_in01 = reg_0104;
    93: op1_06_in01 = reg_0388;
    94: op1_06_in01 = imem01_in[11:8];
    default: op1_06_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv01 = 1;
    5: op1_06_inv01 = 1;
    9: op1_06_inv01 = 1;
    13: op1_06_inv01 = 1;
    15: op1_06_inv01 = 1;
    16: op1_06_inv01 = 1;
    18: op1_06_inv01 = 1;
    19: op1_06_inv01 = 1;
    21: op1_06_inv01 = 1;
    24: op1_06_inv01 = 1;
    27: op1_06_inv01 = 1;
    28: op1_06_inv01 = 1;
    31: op1_06_inv01 = 1;
    32: op1_06_inv01 = 1;
    37: op1_06_inv01 = 1;
    38: op1_06_inv01 = 1;
    39: op1_06_inv01 = 1;
    45: op1_06_inv01 = 1;
    49: op1_06_inv01 = 1;
    51: op1_06_inv01 = 1;
    52: op1_06_inv01 = 1;
    53: op1_06_inv01 = 1;
    55: op1_06_inv01 = 1;
    56: op1_06_inv01 = 1;
    57: op1_06_inv01 = 1;
    58: op1_06_inv01 = 1;
    61: op1_06_inv01 = 1;
    62: op1_06_inv01 = 1;
    63: op1_06_inv01 = 1;
    66: op1_06_inv01 = 1;
    71: op1_06_inv01 = 1;
    74: op1_06_inv01 = 1;
    77: op1_06_inv01 = 1;
    80: op1_06_inv01 = 1;
    83: op1_06_inv01 = 1;
    84: op1_06_inv01 = 1;
    87: op1_06_inv01 = 1;
    90: op1_06_inv01 = 1;
    91: op1_06_inv01 = 1;
    93: op1_06_inv01 = 1;
    94: op1_06_inv01 = 1;
    default: op1_06_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in02 = imem02_in[3:0];
    5: op1_06_in02 = imem00_in[123:120];
    6: op1_06_in02 = reg_0804;
    7: op1_06_in02 = reg_0039;
    8: op1_06_in02 = imem02_in[23:20];
    9: op1_06_in02 = imem00_in[27:24];
    10: op1_06_in02 = reg_0248;
    11: op1_06_in02 = imem00_in[75:72];
    3: op1_06_in02 = imem07_in[83:80];
    12: op1_06_in02 = reg_0299;
    13: op1_06_in02 = reg_0752;
    14: op1_06_in02 = imem00_in[83:80];
    15: op1_06_in02 = reg_0576;
    84: op1_06_in02 = reg_0576;
    16: op1_06_in02 = imem05_in[15:12];
    30: op1_06_in02 = imem05_in[15:12];
    17: op1_06_in02 = reg_0662;
    18: op1_06_in02 = imem06_in[67:64];
    2: op1_06_in02 = imem07_in[87:84];
    19: op1_06_in02 = imem02_in[75:72];
    20: op1_06_in02 = reg_0277;
    21: op1_06_in02 = reg_0243;
    22: op1_06_in02 = reg_0243;
    23: op1_06_in02 = reg_0677;
    24: op1_06_in02 = reg_0581;
    25: op1_06_in02 = reg_0307;
    26: op1_06_in02 = reg_0580;
    27: op1_06_in02 = reg_0053;
    28: op1_06_in02 = reg_0123;
    29: op1_06_in02 = imem02_in[123:120];
    75: op1_06_in02 = imem02_in[123:120];
    31: op1_06_in02 = imem00_in[55:52];
    67: op1_06_in02 = imem00_in[55:52];
    70: op1_06_in02 = imem00_in[55:52];
    32: op1_06_in02 = reg_0515;
    33: op1_06_in02 = reg_0373;
    34: op1_06_in02 = imem00_in[35:32];
    36: op1_06_in02 = imem00_in[67:64];
    96: op1_06_in02 = imem00_in[67:64];
    37: op1_06_in02 = imem00_in[63:60];
    57: op1_06_in02 = imem00_in[63:60];
    38: op1_06_in02 = reg_0504;
    39: op1_06_in02 = reg_0014;
    52: op1_06_in02 = reg_0014;
    40: op1_06_in02 = reg_0652;
    41: op1_06_in02 = reg_0620;
    42: op1_06_in02 = imem00_in[99:96];
    43: op1_06_in02 = imem02_in[119:116];
    44: op1_06_in02 = reg_0796;
    45: op1_06_in02 = reg_0726;
    46: op1_06_in02 = reg_0216;
    47: op1_06_in02 = reg_0510;
    48: op1_06_in02 = reg_0182;
    49: op1_06_in02 = imem06_in[11:8];
    50: op1_06_in02 = reg_0503;
    51: op1_06_in02 = reg_0126;
    53: op1_06_in02 = reg_0227;
    54: op1_06_in02 = reg_0628;
    55: op1_06_in02 = reg_0619;
    56: op1_06_in02 = reg_0183;
    58: op1_06_in02 = reg_0704;
    59: op1_06_in02 = reg_0734;
    60: op1_06_in02 = reg_0492;
    61: op1_06_in02 = reg_0125;
    62: op1_06_in02 = reg_0797;
    63: op1_06_in02 = reg_0285;
    64: op1_06_in02 = reg_0706;
    65: op1_06_in02 = imem07_in[59:56];
    66: op1_06_in02 = reg_0549;
    68: op1_06_in02 = reg_0570;
    69: op1_06_in02 = reg_0134;
    71: op1_06_in02 = reg_0146;
    72: op1_06_in02 = imem07_in[43:40];
    73: op1_06_in02 = reg_0267;
    74: op1_06_in02 = reg_0695;
    76: op1_06_in02 = reg_0674;
    77: op1_06_in02 = imem03_in[11:8];
    78: op1_06_in02 = imem06_in[103:100];
    79: op1_06_in02 = reg_0253;
    80: op1_06_in02 = reg_0683;
    81: op1_06_in02 = reg_0268;
    82: op1_06_in02 = reg_0075;
    83: op1_06_in02 = reg_0506;
    85: op1_06_in02 = imem00_in[19:16];
    86: op1_06_in02 = imem04_in[119:116];
    87: op1_06_in02 = imem06_in[47:44];
    88: op1_06_in02 = reg_0639;
    89: op1_06_in02 = reg_0621;
    90: op1_06_in02 = reg_0334;
    91: op1_06_in02 = reg_0157;
    92: op1_06_in02 = reg_0120;
    93: op1_06_in02 = reg_0424;
    94: op1_06_in02 = imem01_in[47:44];
    95: op1_06_in02 = reg_0675;
    default: op1_06_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv02 = 1;
    5: op1_06_inv02 = 1;
    6: op1_06_inv02 = 1;
    7: op1_06_inv02 = 1;
    8: op1_06_inv02 = 1;
    11: op1_06_inv02 = 1;
    14: op1_06_inv02 = 1;
    16: op1_06_inv02 = 1;
    17: op1_06_inv02 = 1;
    18: op1_06_inv02 = 1;
    2: op1_06_inv02 = 1;
    20: op1_06_inv02 = 1;
    21: op1_06_inv02 = 1;
    23: op1_06_inv02 = 1;
    24: op1_06_inv02 = 1;
    25: op1_06_inv02 = 1;
    26: op1_06_inv02 = 1;
    27: op1_06_inv02 = 1;
    29: op1_06_inv02 = 1;
    34: op1_06_inv02 = 1;
    37: op1_06_inv02 = 1;
    38: op1_06_inv02 = 1;
    39: op1_06_inv02 = 1;
    40: op1_06_inv02 = 1;
    41: op1_06_inv02 = 1;
    42: op1_06_inv02 = 1;
    43: op1_06_inv02 = 1;
    44: op1_06_inv02 = 1;
    45: op1_06_inv02 = 1;
    46: op1_06_inv02 = 1;
    48: op1_06_inv02 = 1;
    49: op1_06_inv02 = 1;
    51: op1_06_inv02 = 1;
    52: op1_06_inv02 = 1;
    54: op1_06_inv02 = 1;
    55: op1_06_inv02 = 1;
    59: op1_06_inv02 = 1;
    60: op1_06_inv02 = 1;
    63: op1_06_inv02 = 1;
    66: op1_06_inv02 = 1;
    68: op1_06_inv02 = 1;
    69: op1_06_inv02 = 1;
    71: op1_06_inv02 = 1;
    72: op1_06_inv02 = 1;
    73: op1_06_inv02 = 1;
    74: op1_06_inv02 = 1;
    75: op1_06_inv02 = 1;
    76: op1_06_inv02 = 1;
    80: op1_06_inv02 = 1;
    81: op1_06_inv02 = 1;
    82: op1_06_inv02 = 1;
    83: op1_06_inv02 = 1;
    86: op1_06_inv02 = 1;
    90: op1_06_inv02 = 1;
    94: op1_06_inv02 = 1;
    96: op1_06_inv02 = 1;
    default: op1_06_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in03 = imem02_in[7:4];
    5: op1_06_in03 = reg_0681;
    6: op1_06_in03 = reg_0802;
    52: op1_06_in03 = reg_0802;
    7: op1_06_in03 = reg_0031;
    8: op1_06_in03 = imem02_in[31:28];
    9: op1_06_in03 = imem00_in[31:28];
    10: op1_06_in03 = reg_0237;
    11: op1_06_in03 = imem00_in[103:100];
    3: op1_06_in03 = imem07_in[99:96];
    12: op1_06_in03 = reg_0302;
    13: op1_06_in03 = reg_0005;
    14: op1_06_in03 = imem00_in[107:104];
    15: op1_06_in03 = reg_0395;
    16: op1_06_in03 = imem05_in[19:16];
    17: op1_06_in03 = reg_0352;
    18: op1_06_in03 = imem06_in[99:96];
    2: op1_06_in03 = imem07_in[91:88];
    19: op1_06_in03 = imem02_in[115:112];
    20: op1_06_in03 = reg_0086;
    21: op1_06_in03 = reg_0107;
    22: op1_06_in03 = reg_0123;
    23: op1_06_in03 = reg_0680;
    60: op1_06_in03 = reg_0680;
    89: op1_06_in03 = reg_0680;
    24: op1_06_in03 = reg_0595;
    25: op1_06_in03 = reg_0277;
    26: op1_06_in03 = reg_0590;
    27: op1_06_in03 = reg_0297;
    28: op1_06_in03 = reg_0100;
    29: op1_06_in03 = imem02_in[127:124];
    43: op1_06_in03 = imem02_in[127:124];
    30: op1_06_in03 = imem05_in[59:56];
    31: op1_06_in03 = imem00_in[79:76];
    32: op1_06_in03 = reg_0559;
    33: op1_06_in03 = reg_0569;
    34: op1_06_in03 = imem00_in[39:36];
    36: op1_06_in03 = imem00_in[95:92];
    37: op1_06_in03 = imem00_in[67:64];
    57: op1_06_in03 = imem00_in[67:64];
    38: op1_06_in03 = reg_0243;
    39: op1_06_in03 = reg_0016;
    40: op1_06_in03 = reg_0667;
    41: op1_06_in03 = reg_0819;
    42: op1_06_in03 = imem00_in[123:120];
    44: op1_06_in03 = reg_0488;
    45: op1_06_in03 = reg_0703;
    46: op1_06_in03 = reg_0220;
    47: op1_06_in03 = reg_0071;
    48: op1_06_in03 = reg_0177;
    49: op1_06_in03 = imem06_in[55:52];
    50: op1_06_in03 = reg_0074;
    51: op1_06_in03 = reg_0354;
    53: op1_06_in03 = reg_0296;
    54: op1_06_in03 = reg_0624;
    55: op1_06_in03 = reg_0293;
    56: op1_06_in03 = reg_0164;
    58: op1_06_in03 = reg_0724;
    59: op1_06_in03 = reg_0487;
    61: op1_06_in03 = reg_0670;
    62: op1_06_in03 = reg_0795;
    63: op1_06_in03 = reg_0133;
    64: op1_06_in03 = reg_0441;
    65: op1_06_in03 = imem07_in[79:76];
    66: op1_06_in03 = reg_0787;
    67: op1_06_in03 = reg_0694;
    68: op1_06_in03 = reg_0807;
    69: op1_06_in03 = imem06_in[7:4];
    70: op1_06_in03 = imem00_in[63:60];
    71: op1_06_in03 = imem06_in[91:88];
    72: op1_06_in03 = imem07_in[59:56];
    73: op1_06_in03 = reg_0173;
    74: op1_06_in03 = reg_0492;
    75: op1_06_in03 = reg_0325;
    76: op1_06_in03 = imem02_in[23:20];
    77: op1_06_in03 = imem03_in[127:124];
    78: op1_06_in03 = imem06_in[115:112];
    79: op1_06_in03 = reg_0295;
    80: op1_06_in03 = reg_0696;
    81: op1_06_in03 = imem07_in[3:0];
    82: op1_06_in03 = reg_0059;
    83: op1_06_in03 = reg_0073;
    84: op1_06_in03 = reg_0039;
    85: op1_06_in03 = imem00_in[35:32];
    86: op1_06_in03 = imem04_in[123:120];
    87: op1_06_in03 = imem06_in[59:56];
    88: op1_06_in03 = reg_0647;
    90: op1_06_in03 = reg_0064;
    91: op1_06_in03 = reg_0334;
    92: op1_06_in03 = reg_0106;
    93: op1_06_in03 = reg_0105;
    94: op1_06_in03 = imem01_in[51:48];
    95: op1_06_in03 = reg_0127;
    96: op1_06_in03 = imem00_in[75:72];
    default: op1_06_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv03 = 1;
    6: op1_06_inv03 = 1;
    8: op1_06_inv03 = 1;
    9: op1_06_inv03 = 1;
    10: op1_06_inv03 = 1;
    11: op1_06_inv03 = 1;
    12: op1_06_inv03 = 1;
    14: op1_06_inv03 = 1;
    17: op1_06_inv03 = 1;
    19: op1_06_inv03 = 1;
    20: op1_06_inv03 = 1;
    22: op1_06_inv03 = 1;
    23: op1_06_inv03 = 1;
    25: op1_06_inv03 = 1;
    29: op1_06_inv03 = 1;
    30: op1_06_inv03 = 1;
    33: op1_06_inv03 = 1;
    34: op1_06_inv03 = 1;
    38: op1_06_inv03 = 1;
    39: op1_06_inv03 = 1;
    40: op1_06_inv03 = 1;
    41: op1_06_inv03 = 1;
    46: op1_06_inv03 = 1;
    47: op1_06_inv03 = 1;
    50: op1_06_inv03 = 1;
    53: op1_06_inv03 = 1;
    54: op1_06_inv03 = 1;
    56: op1_06_inv03 = 1;
    58: op1_06_inv03 = 1;
    60: op1_06_inv03 = 1;
    61: op1_06_inv03 = 1;
    66: op1_06_inv03 = 1;
    68: op1_06_inv03 = 1;
    69: op1_06_inv03 = 1;
    71: op1_06_inv03 = 1;
    72: op1_06_inv03 = 1;
    74: op1_06_inv03 = 1;
    79: op1_06_inv03 = 1;
    81: op1_06_inv03 = 1;
    83: op1_06_inv03 = 1;
    89: op1_06_inv03 = 1;
    91: op1_06_inv03 = 1;
    93: op1_06_inv03 = 1;
    default: op1_06_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in04 = imem02_in[47:44];
    5: op1_06_in04 = reg_0686;
    67: op1_06_in04 = reg_0686;
    6: op1_06_in04 = imem04_in[11:8];
    7: op1_06_in04 = reg_0034;
    8: op1_06_in04 = imem02_in[51:48];
    9: op1_06_in04 = imem00_in[35:32];
    10: op1_06_in04 = reg_0504;
    11: op1_06_in04 = reg_0697;
    3: op1_06_in04 = reg_0424;
    12: op1_06_in04 = reg_0298;
    13: op1_06_in04 = imem07_in[15:12];
    14: op1_06_in04 = reg_0693;
    42: op1_06_in04 = reg_0693;
    15: op1_06_in04 = reg_0376;
    33: op1_06_in04 = reg_0376;
    16: op1_06_in04 = imem05_in[27:24];
    17: op1_06_in04 = reg_0357;
    18: op1_06_in04 = imem06_in[103:100];
    2: op1_06_in04 = imem07_in[107:104];
    19: op1_06_in04 = reg_0650;
    20: op1_06_in04 = reg_0149;
    21: op1_06_in04 = reg_0117;
    22: op1_06_in04 = reg_0103;
    23: op1_06_in04 = reg_0453;
    24: op1_06_in04 = reg_0590;
    25: op1_06_in04 = reg_0147;
    26: op1_06_in04 = reg_0395;
    27: op1_06_in04 = reg_0292;
    28: op1_06_in04 = imem02_in[3:0];
    29: op1_06_in04 = reg_0658;
    30: op1_06_in04 = imem05_in[79:76];
    31: op1_06_in04 = imem00_in[111:108];
    96: op1_06_in04 = imem00_in[111:108];
    32: op1_06_in04 = reg_0232;
    34: op1_06_in04 = imem00_in[43:40];
    36: op1_06_in04 = imem00_in[107:104];
    37: op1_06_in04 = imem00_in[115:112];
    38: op1_06_in04 = reg_0104;
    39: op1_06_in04 = imem04_in[7:4];
    68: op1_06_in04 = imem04_in[7:4];
    40: op1_06_in04 = reg_0344;
    41: op1_06_in04 = reg_0037;
    43: op1_06_in04 = reg_0660;
    44: op1_06_in04 = reg_0492;
    80: op1_06_in04 = reg_0492;
    45: op1_06_in04 = reg_0729;
    46: op1_06_in04 = reg_0603;
    47: op1_06_in04 = reg_0616;
    49: op1_06_in04 = imem06_in[67:64];
    50: op1_06_in04 = reg_0343;
    51: op1_06_in04 = reg_0105;
    52: op1_06_in04 = imem04_in[99:96];
    53: op1_06_in04 = reg_0519;
    54: op1_06_in04 = reg_0020;
    55: op1_06_in04 = reg_0577;
    56: op1_06_in04 = reg_0168;
    57: op1_06_in04 = imem00_in[99:96];
    58: op1_06_in04 = reg_0709;
    59: op1_06_in04 = reg_0235;
    60: op1_06_in04 = reg_0454;
    61: op1_06_in04 = reg_0592;
    62: op1_06_in04 = reg_0288;
    63: op1_06_in04 = reg_0152;
    64: op1_06_in04 = reg_0436;
    65: op1_06_in04 = imem07_in[95:92];
    66: op1_06_in04 = imem07_in[75:72];
    69: op1_06_in04 = imem06_in[39:36];
    70: op1_06_in04 = imem00_in[67:64];
    71: op1_06_in04 = imem06_in[107:104];
    72: op1_06_in04 = imem07_in[63:60];
    73: op1_06_in04 = reg_0171;
    74: op1_06_in04 = reg_0749;
    75: op1_06_in04 = reg_0739;
    76: op1_06_in04 = imem02_in[59:56];
    77: op1_06_in04 = reg_0493;
    78: op1_06_in04 = reg_0625;
    79: op1_06_in04 = reg_0434;
    81: op1_06_in04 = imem07_in[23:20];
    82: op1_06_in04 = reg_0256;
    83: op1_06_in04 = reg_0670;
    84: op1_06_in04 = reg_0700;
    85: op1_06_in04 = imem00_in[127:124];
    86: op1_06_in04 = reg_0544;
    87: op1_06_in04 = imem06_in[75:72];
    88: op1_06_in04 = reg_0087;
    89: op1_06_in04 = reg_0224;
    90: op1_06_in04 = reg_0253;
    91: op1_06_in04 = reg_0636;
    92: op1_06_in04 = imem02_in[11:8];
    93: op1_06_in04 = reg_0122;
    94: op1_06_in04 = imem01_in[63:60];
    95: op1_06_in04 = reg_0121;
    default: op1_06_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv04 = 1;
    7: op1_06_inv04 = 1;
    8: op1_06_inv04 = 1;
    10: op1_06_inv04 = 1;
    13: op1_06_inv04 = 1;
    14: op1_06_inv04 = 1;
    16: op1_06_inv04 = 1;
    19: op1_06_inv04 = 1;
    20: op1_06_inv04 = 1;
    23: op1_06_inv04 = 1;
    25: op1_06_inv04 = 1;
    28: op1_06_inv04 = 1;
    30: op1_06_inv04 = 1;
    31: op1_06_inv04 = 1;
    32: op1_06_inv04 = 1;
    33: op1_06_inv04 = 1;
    36: op1_06_inv04 = 1;
    37: op1_06_inv04 = 1;
    39: op1_06_inv04 = 1;
    40: op1_06_inv04 = 1;
    41: op1_06_inv04 = 1;
    42: op1_06_inv04 = 1;
    43: op1_06_inv04 = 1;
    49: op1_06_inv04 = 1;
    50: op1_06_inv04 = 1;
    55: op1_06_inv04 = 1;
    56: op1_06_inv04 = 1;
    57: op1_06_inv04 = 1;
    58: op1_06_inv04 = 1;
    59: op1_06_inv04 = 1;
    60: op1_06_inv04 = 1;
    61: op1_06_inv04 = 1;
    62: op1_06_inv04 = 1;
    63: op1_06_inv04 = 1;
    66: op1_06_inv04 = 1;
    68: op1_06_inv04 = 1;
    69: op1_06_inv04 = 1;
    71: op1_06_inv04 = 1;
    72: op1_06_inv04 = 1;
    74: op1_06_inv04 = 1;
    75: op1_06_inv04 = 1;
    76: op1_06_inv04 = 1;
    77: op1_06_inv04 = 1;
    80: op1_06_inv04 = 1;
    81: op1_06_inv04 = 1;
    82: op1_06_inv04 = 1;
    83: op1_06_inv04 = 1;
    84: op1_06_inv04 = 1;
    87: op1_06_inv04 = 1;
    88: op1_06_inv04 = 1;
    89: op1_06_inv04 = 1;
    91: op1_06_inv04 = 1;
    93: op1_06_inv04 = 1;
    default: op1_06_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in05 = imem02_in[71:68];
    8: op1_06_in05 = imem02_in[71:68];
    5: op1_06_in05 = reg_0691;
    6: op1_06_in05 = imem04_in[87:84];
    7: op1_06_in05 = reg_0035;
    9: op1_06_in05 = imem00_in[39:36];
    10: op1_06_in05 = reg_0041;
    11: op1_06_in05 = reg_0686;
    31: op1_06_in05 = reg_0686;
    3: op1_06_in05 = reg_0428;
    12: op1_06_in05 = reg_0278;
    13: op1_06_in05 = imem07_in[51:48];
    14: op1_06_in05 = reg_0683;
    15: op1_06_in05 = reg_0309;
    16: op1_06_in05 = imem05_in[51:48];
    17: op1_06_in05 = reg_0345;
    18: op1_06_in05 = imem06_in[111:108];
    2: op1_06_in05 = imem07_in[123:120];
    65: op1_06_in05 = imem07_in[123:120];
    66: op1_06_in05 = imem07_in[123:120];
    19: op1_06_in05 = reg_0655;
    20: op1_06_in05 = reg_0145;
    21: op1_06_in05 = reg_0113;
    22: op1_06_in05 = reg_0100;
    23: op1_06_in05 = reg_0476;
    24: op1_06_in05 = reg_0391;
    25: op1_06_in05 = reg_0135;
    26: op1_06_in05 = reg_0384;
    27: op1_06_in05 = reg_0079;
    28: op1_06_in05 = imem02_in[27:24];
    29: op1_06_in05 = reg_0640;
    30: op1_06_in05 = imem05_in[107:104];
    32: op1_06_in05 = reg_0505;
    33: op1_06_in05 = reg_0389;
    34: op1_06_in05 = imem00_in[51:48];
    36: op1_06_in05 = imem00_in[119:116];
    37: op1_06_in05 = imem00_in[119:116];
    38: op1_06_in05 = reg_0099;
    39: op1_06_in05 = imem04_in[31:28];
    40: op1_06_in05 = reg_0354;
    41: op1_06_in05 = reg_0818;
    42: op1_06_in05 = reg_0676;
    43: op1_06_in05 = reg_0662;
    44: op1_06_in05 = reg_0493;
    45: op1_06_in05 = reg_0718;
    46: op1_06_in05 = reg_0119;
    61: op1_06_in05 = reg_0119;
    47: op1_06_in05 = reg_0503;
    49: op1_06_in05 = imem06_in[75:72];
    50: op1_06_in05 = reg_0062;
    51: op1_06_in05 = reg_0104;
    52: op1_06_in05 = imem04_in[111:108];
    53: op1_06_in05 = reg_0644;
    54: op1_06_in05 = reg_0609;
    55: op1_06_in05 = reg_0762;
    78: op1_06_in05 = reg_0762;
    56: op1_06_in05 = reg_0170;
    57: op1_06_in05 = imem00_in[103:100];
    58: op1_06_in05 = reg_0635;
    59: op1_06_in05 = reg_0423;
    60: op1_06_in05 = reg_0450;
    62: op1_06_in05 = reg_0783;
    63: op1_06_in05 = reg_0156;
    64: op1_06_in05 = reg_0268;
    67: op1_06_in05 = reg_0749;
    68: op1_06_in05 = imem04_in[43:40];
    69: op1_06_in05 = imem06_in[59:56];
    70: op1_06_in05 = imem00_in[75:72];
    71: op1_06_in05 = reg_0619;
    72: op1_06_in05 = imem07_in[71:68];
    74: op1_06_in05 = reg_0407;
    75: op1_06_in05 = reg_0304;
    76: op1_06_in05 = imem02_in[91:88];
    77: op1_06_in05 = reg_0318;
    79: op1_06_in05 = reg_0443;
    80: op1_06_in05 = reg_0690;
    81: op1_06_in05 = imem07_in[27:24];
    82: op1_06_in05 = imem04_in[75:72];
    83: op1_06_in05 = reg_0592;
    84: op1_06_in05 = reg_0620;
    85: op1_06_in05 = reg_0697;
    86: op1_06_in05 = reg_0171;
    87: op1_06_in05 = imem06_in[83:80];
    88: op1_06_in05 = reg_0374;
    89: op1_06_in05 = reg_0764;
    90: op1_06_in05 = reg_0295;
    91: op1_06_in05 = reg_0061;
    92: op1_06_in05 = imem02_in[35:32];
    93: op1_06_in05 = reg_0660;
    94: op1_06_in05 = imem01_in[87:84];
    95: op1_06_in05 = reg_0126;
    96: op1_06_in05 = reg_0744;
    default: op1_06_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv05 = 1;
    10: op1_06_inv05 = 1;
    14: op1_06_inv05 = 1;
    17: op1_06_inv05 = 1;
    20: op1_06_inv05 = 1;
    21: op1_06_inv05 = 1;
    22: op1_06_inv05 = 1;
    23: op1_06_inv05 = 1;
    24: op1_06_inv05 = 1;
    27: op1_06_inv05 = 1;
    29: op1_06_inv05 = 1;
    31: op1_06_inv05 = 1;
    36: op1_06_inv05 = 1;
    37: op1_06_inv05 = 1;
    40: op1_06_inv05 = 1;
    41: op1_06_inv05 = 1;
    44: op1_06_inv05 = 1;
    45: op1_06_inv05 = 1;
    50: op1_06_inv05 = 1;
    52: op1_06_inv05 = 1;
    53: op1_06_inv05 = 1;
    54: op1_06_inv05 = 1;
    59: op1_06_inv05 = 1;
    61: op1_06_inv05 = 1;
    62: op1_06_inv05 = 1;
    64: op1_06_inv05 = 1;
    65: op1_06_inv05 = 1;
    66: op1_06_inv05 = 1;
    68: op1_06_inv05 = 1;
    70: op1_06_inv05 = 1;
    72: op1_06_inv05 = 1;
    74: op1_06_inv05 = 1;
    78: op1_06_inv05 = 1;
    82: op1_06_inv05 = 1;
    83: op1_06_inv05 = 1;
    84: op1_06_inv05 = 1;
    87: op1_06_inv05 = 1;
    91: op1_06_inv05 = 1;
    94: op1_06_inv05 = 1;
    96: op1_06_inv05 = 1;
    default: op1_06_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in06 = imem02_in[103:100];
    5: op1_06_in06 = reg_0680;
    6: op1_06_in06 = reg_0536;
    7: op1_06_in06 = reg_0040;
    8: op1_06_in06 = imem02_in[107:104];
    76: op1_06_in06 = imem02_in[107:104];
    9: op1_06_in06 = imem00_in[55:52];
    10: op1_06_in06 = reg_0122;
    11: op1_06_in06 = reg_0673;
    3: op1_06_in06 = reg_0434;
    12: op1_06_in06 = reg_0062;
    13: op1_06_in06 = imem07_in[79:76];
    72: op1_06_in06 = imem07_in[79:76];
    14: op1_06_in06 = reg_0685;
    85: op1_06_in06 = reg_0685;
    15: op1_06_in06 = reg_0012;
    16: op1_06_in06 = imem05_in[71:68];
    17: op1_06_in06 = reg_0363;
    18: op1_06_in06 = imem06_in[127:124];
    2: op1_06_in06 = imem07_in[127:124];
    19: op1_06_in06 = reg_0647;
    20: op1_06_in06 = reg_0151;
    21: op1_06_in06 = imem02_in[3:0];
    22: op1_06_in06 = reg_0110;
    23: op1_06_in06 = reg_0475;
    24: op1_06_in06 = reg_0397;
    25: op1_06_in06 = reg_0143;
    26: op1_06_in06 = reg_0388;
    27: op1_06_in06 = reg_0067;
    28: op1_06_in06 = imem02_in[67:64];
    29: op1_06_in06 = reg_0344;
    30: op1_06_in06 = imem05_in[119:116];
    31: op1_06_in06 = reg_0670;
    32: op1_06_in06 = reg_0242;
    33: op1_06_in06 = reg_0007;
    34: op1_06_in06 = imem00_in[79:76];
    36: op1_06_in06 = imem00_in[123:120];
    37: op1_06_in06 = reg_0697;
    38: op1_06_in06 = reg_0114;
    39: op1_06_in06 = imem04_in[39:36];
    40: op1_06_in06 = reg_0092;
    41: op1_06_in06 = reg_0231;
    42: op1_06_in06 = reg_0679;
    43: op1_06_in06 = reg_0665;
    44: op1_06_in06 = reg_0784;
    45: op1_06_in06 = reg_0701;
    46: op1_06_in06 = reg_0100;
    47: op1_06_in06 = reg_0292;
    49: op1_06_in06 = imem06_in[79:76];
    50: op1_06_in06 = reg_0585;
    51: op1_06_in06 = reg_0347;
    52: op1_06_in06 = reg_0262;
    53: op1_06_in06 = imem05_in[23:20];
    54: op1_06_in06 = reg_0618;
    55: op1_06_in06 = reg_0763;
    56: op1_06_in06 = reg_0171;
    57: op1_06_in06 = reg_0693;
    58: op1_06_in06 = reg_0160;
    59: op1_06_in06 = reg_0567;
    60: op1_06_in06 = reg_0451;
    61: op1_06_in06 = reg_0676;
    93: op1_06_in06 = reg_0676;
    62: op1_06_in06 = reg_0786;
    63: op1_06_in06 = reg_0138;
    64: op1_06_in06 = reg_0175;
    65: op1_06_in06 = reg_0722;
    66: op1_06_in06 = reg_0707;
    67: op1_06_in06 = reg_0658;
    68: op1_06_in06 = imem04_in[55:52];
    69: op1_06_in06 = imem06_in[107:104];
    70: op1_06_in06 = imem00_in[111:108];
    71: op1_06_in06 = reg_0339;
    74: op1_06_in06 = reg_0633;
    75: op1_06_in06 = reg_0655;
    77: op1_06_in06 = reg_0357;
    78: op1_06_in06 = reg_0815;
    79: op1_06_in06 = reg_0437;
    80: op1_06_in06 = reg_0463;
    81: op1_06_in06 = imem07_in[31:28];
    82: op1_06_in06 = imem04_in[79:76];
    83: op1_06_in06 = reg_0108;
    84: op1_06_in06 = reg_0367;
    86: op1_06_in06 = reg_0275;
    87: op1_06_in06 = imem06_in[99:96];
    88: op1_06_in06 = reg_0705;
    89: op1_06_in06 = imem07_in[19:16];
    90: op1_06_in06 = reg_0449;
    91: op1_06_in06 = reg_0445;
    92: op1_06_in06 = imem02_in[91:88];
    94: op1_06_in06 = imem01_in[95:92];
    95: op1_06_in06 = imem02_in[39:36];
    96: op1_06_in06 = reg_0145;
    default: op1_06_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv06 = 1;
    7: op1_06_inv06 = 1;
    9: op1_06_inv06 = 1;
    10: op1_06_inv06 = 1;
    11: op1_06_inv06 = 1;
    12: op1_06_inv06 = 1;
    13: op1_06_inv06 = 1;
    15: op1_06_inv06 = 1;
    16: op1_06_inv06 = 1;
    2: op1_06_inv06 = 1;
    22: op1_06_inv06 = 1;
    23: op1_06_inv06 = 1;
    25: op1_06_inv06 = 1;
    28: op1_06_inv06 = 1;
    32: op1_06_inv06 = 1;
    33: op1_06_inv06 = 1;
    36: op1_06_inv06 = 1;
    37: op1_06_inv06 = 1;
    38: op1_06_inv06 = 1;
    39: op1_06_inv06 = 1;
    41: op1_06_inv06 = 1;
    43: op1_06_inv06 = 1;
    44: op1_06_inv06 = 1;
    45: op1_06_inv06 = 1;
    49: op1_06_inv06 = 1;
    51: op1_06_inv06 = 1;
    52: op1_06_inv06 = 1;
    54: op1_06_inv06 = 1;
    58: op1_06_inv06 = 1;
    62: op1_06_inv06 = 1;
    64: op1_06_inv06 = 1;
    65: op1_06_inv06 = 1;
    66: op1_06_inv06 = 1;
    67: op1_06_inv06 = 1;
    68: op1_06_inv06 = 1;
    69: op1_06_inv06 = 1;
    74: op1_06_inv06 = 1;
    75: op1_06_inv06 = 1;
    81: op1_06_inv06 = 1;
    86: op1_06_inv06 = 1;
    89: op1_06_inv06 = 1;
    90: op1_06_inv06 = 1;
    93: op1_06_inv06 = 1;
    95: op1_06_inv06 = 1;
    96: op1_06_inv06 = 1;
    default: op1_06_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in07 = imem02_in[111:108];
    92: op1_06_in07 = imem02_in[111:108];
    5: op1_06_in07 = reg_0687;
    11: op1_06_in07 = reg_0687;
    6: op1_06_in07 = reg_0550;
    7: op1_06_in07 = reg_0030;
    8: op1_06_in07 = imem02_in[115:112];
    9: op1_06_in07 = reg_0463;
    67: op1_06_in07 = reg_0463;
    10: op1_06_in07 = reg_0120;
    3: op1_06_in07 = reg_0435;
    12: op1_06_in07 = reg_0065;
    50: op1_06_in07 = reg_0065;
    13: op1_06_in07 = imem07_in[99:96];
    14: op1_06_in07 = reg_0698;
    15: op1_06_in07 = reg_0807;
    16: op1_06_in07 = imem05_in[99:96];
    17: op1_06_in07 = reg_0338;
    18: op1_06_in07 = reg_0614;
    2: op1_06_in07 = reg_0174;
    19: op1_06_in07 = reg_0643;
    20: op1_06_in07 = reg_0129;
    63: op1_06_in07 = reg_0129;
    21: op1_06_in07 = imem02_in[11:8];
    22: op1_06_in07 = imem02_in[23:20];
    23: op1_06_in07 = reg_0472;
    60: op1_06_in07 = reg_0472;
    24: op1_06_in07 = reg_0393;
    25: op1_06_in07 = imem06_in[7:4];
    26: op1_06_in07 = reg_0385;
    27: op1_06_in07 = reg_0071;
    28: op1_06_in07 = imem02_in[75:72];
    29: op1_06_in07 = reg_0354;
    30: op1_06_in07 = reg_0789;
    31: op1_06_in07 = reg_0679;
    32: op1_06_in07 = reg_0216;
    33: op1_06_in07 = reg_0805;
    34: op1_06_in07 = imem00_in[87:84];
    36: op1_06_in07 = reg_0697;
    57: op1_06_in07 = reg_0697;
    70: op1_06_in07 = reg_0697;
    37: op1_06_in07 = reg_0685;
    38: op1_06_in07 = imem02_in[47:44];
    39: op1_06_in07 = imem04_in[75:72];
    40: op1_06_in07 = reg_0498;
    41: op1_06_in07 = reg_0029;
    42: op1_06_in07 = reg_0674;
    93: op1_06_in07 = reg_0674;
    43: op1_06_in07 = reg_0667;
    44: op1_06_in07 = reg_0279;
    45: op1_06_in07 = reg_0295;
    46: op1_06_in07 = reg_0110;
    47: op1_06_in07 = reg_0512;
    49: op1_06_in07 = imem06_in[103:100];
    51: op1_06_in07 = reg_0650;
    52: op1_06_in07 = reg_0544;
    53: op1_06_in07 = imem05_in[43:40];
    54: op1_06_in07 = reg_0622;
    55: op1_06_in07 = reg_0753;
    58: op1_06_in07 = reg_0183;
    59: op1_06_in07 = reg_0425;
    61: op1_06_in07 = reg_0678;
    62: op1_06_in07 = reg_0070;
    64: op1_06_in07 = reg_0167;
    65: op1_06_in07 = reg_0721;
    66: op1_06_in07 = reg_0727;
    68: op1_06_in07 = imem04_in[63:60];
    69: op1_06_in07 = reg_0299;
    71: op1_06_in07 = reg_0293;
    72: op1_06_in07 = imem07_in[83:80];
    74: op1_06_in07 = reg_0450;
    75: op1_06_in07 = reg_0702;
    76: op1_06_in07 = imem02_in[123:120];
    77: op1_06_in07 = reg_0395;
    78: op1_06_in07 = reg_0409;
    79: op1_06_in07 = reg_0448;
    80: op1_06_in07 = reg_0457;
    81: op1_06_in07 = imem07_in[43:40];
    82: op1_06_in07 = imem04_in[123:120];
    83: op1_06_in07 = reg_0121;
    84: op1_06_in07 = imem07_in[39:36];
    85: op1_06_in07 = reg_0689;
    86: op1_06_in07 = reg_0060;
    87: op1_06_in07 = reg_0605;
    88: op1_06_in07 = reg_0414;
    89: op1_06_in07 = imem07_in[31:28];
    90: op1_06_in07 = reg_0267;
    91: op1_06_in07 = reg_0443;
    94: op1_06_in07 = imem01_in[111:108];
    95: op1_06_in07 = imem02_in[103:100];
    96: op1_06_in07 = reg_0171;
    default: op1_06_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_06_inv07 = 1;
    10: op1_06_inv07 = 1;
    11: op1_06_inv07 = 1;
    15: op1_06_inv07 = 1;
    16: op1_06_inv07 = 1;
    18: op1_06_inv07 = 1;
    20: op1_06_inv07 = 1;
    21: op1_06_inv07 = 1;
    24: op1_06_inv07 = 1;
    25: op1_06_inv07 = 1;
    26: op1_06_inv07 = 1;
    28: op1_06_inv07 = 1;
    29: op1_06_inv07 = 1;
    30: op1_06_inv07 = 1;
    31: op1_06_inv07 = 1;
    32: op1_06_inv07 = 1;
    33: op1_06_inv07 = 1;
    34: op1_06_inv07 = 1;
    37: op1_06_inv07 = 1;
    39: op1_06_inv07 = 1;
    40: op1_06_inv07 = 1;
    41: op1_06_inv07 = 1;
    42: op1_06_inv07 = 1;
    47: op1_06_inv07 = 1;
    50: op1_06_inv07 = 1;
    52: op1_06_inv07 = 1;
    55: op1_06_inv07 = 1;
    57: op1_06_inv07 = 1;
    63: op1_06_inv07 = 1;
    65: op1_06_inv07 = 1;
    71: op1_06_inv07 = 1;
    77: op1_06_inv07 = 1;
    80: op1_06_inv07 = 1;
    81: op1_06_inv07 = 1;
    84: op1_06_inv07 = 1;
    86: op1_06_inv07 = 1;
    87: op1_06_inv07 = 1;
    88: op1_06_inv07 = 1;
    89: op1_06_inv07 = 1;
    90: op1_06_inv07 = 1;
    91: op1_06_inv07 = 1;
    92: op1_06_inv07 = 1;
    94: op1_06_inv07 = 1;
    96: op1_06_inv07 = 1;
    default: op1_06_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in08 = imem02_in[127:124];
    5: op1_06_in08 = reg_0454;
    6: op1_06_in08 = reg_0529;
    7: op1_06_in08 = imem07_in[15:12];
    8: op1_06_in08 = imem02_in[123:120];
    9: op1_06_in08 = reg_0457;
    10: op1_06_in08 = reg_0114;
    11: op1_06_in08 = reg_0453;
    3: op1_06_in08 = reg_0161;
    12: op1_06_in08 = reg_0067;
    13: op1_06_in08 = imem07_in[107:104];
    14: op1_06_in08 = reg_0691;
    15: op1_06_in08 = reg_0804;
    16: op1_06_in08 = imem05_in[103:100];
    17: op1_06_in08 = reg_0335;
    18: op1_06_in08 = reg_0607;
    2: op1_06_in08 = reg_0175;
    19: op1_06_in08 = reg_0659;
    71: op1_06_in08 = reg_0659;
    20: op1_06_in08 = reg_0130;
    63: op1_06_in08 = reg_0130;
    21: op1_06_in08 = imem02_in[15:12];
    22: op1_06_in08 = imem02_in[31:28];
    93: op1_06_in08 = imem02_in[31:28];
    23: op1_06_in08 = reg_0467;
    24: op1_06_in08 = reg_0396;
    25: op1_06_in08 = imem06_in[71:68];
    26: op1_06_in08 = reg_0803;
    27: op1_06_in08 = reg_0063;
    28: op1_06_in08 = imem02_in[91:88];
    29: op1_06_in08 = reg_0341;
    30: op1_06_in08 = reg_0492;
    31: op1_06_in08 = reg_0674;
    32: op1_06_in08 = reg_0248;
    33: op1_06_in08 = reg_0802;
    34: op1_06_in08 = imem00_in[99:96];
    36: op1_06_in08 = reg_0698;
    37: op1_06_in08 = reg_0676;
    38: op1_06_in08 = imem02_in[71:68];
    39: op1_06_in08 = imem04_in[91:88];
    40: op1_06_in08 = reg_0526;
    41: op1_06_in08 = reg_0752;
    42: op1_06_in08 = reg_0460;
    43: op1_06_in08 = reg_0357;
    44: op1_06_in08 = reg_0276;
    45: op1_06_in08 = reg_0051;
    46: op1_06_in08 = imem02_in[51:48];
    47: op1_06_in08 = reg_0513;
    49: op1_06_in08 = imem06_in[107:104];
    50: op1_06_in08 = reg_0501;
    51: op1_06_in08 = reg_0666;
    52: op1_06_in08 = reg_0560;
    53: op1_06_in08 = imem05_in[55:52];
    54: op1_06_in08 = reg_0025;
    55: op1_06_in08 = reg_0777;
    57: op1_06_in08 = reg_0681;
    58: op1_06_in08 = reg_0166;
    59: op1_06_in08 = reg_0419;
    60: op1_06_in08 = reg_0474;
    61: op1_06_in08 = imem02_in[7:4];
    62: op1_06_in08 = reg_0226;
    64: op1_06_in08 = reg_0159;
    65: op1_06_in08 = reg_0266;
    66: op1_06_in08 = reg_0334;
    67: op1_06_in08 = reg_0455;
    68: op1_06_in08 = imem04_in[67:64];
    69: op1_06_in08 = reg_0624;
    70: op1_06_in08 = reg_0696;
    72: op1_06_in08 = imem07_in[119:116];
    74: op1_06_in08 = reg_0464;
    80: op1_06_in08 = reg_0464;
    75: op1_06_in08 = reg_0414;
    76: op1_06_in08 = reg_0647;
    77: op1_06_in08 = reg_0028;
    78: op1_06_in08 = reg_0814;
    79: op1_06_in08 = reg_0180;
    82: op1_06_in08 = reg_0052;
    83: op1_06_in08 = reg_0678;
    84: op1_06_in08 = imem07_in[51:48];
    89: op1_06_in08 = imem07_in[51:48];
    85: op1_06_in08 = reg_0684;
    86: op1_06_in08 = reg_0558;
    87: op1_06_in08 = reg_0038;
    88: op1_06_in08 = imem03_in[43:40];
    90: op1_06_in08 = reg_0181;
    91: op1_06_in08 = reg_0448;
    92: op1_06_in08 = reg_0642;
    94: op1_06_in08 = reg_0125;
    95: op1_06_in08 = reg_0541;
    96: op1_06_in08 = reg_0477;
    default: op1_06_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv08 = 1;
    6: op1_06_inv08 = 1;
    9: op1_06_inv08 = 1;
    10: op1_06_inv08 = 1;
    14: op1_06_inv08 = 1;
    17: op1_06_inv08 = 1;
    20: op1_06_inv08 = 1;
    23: op1_06_inv08 = 1;
    26: op1_06_inv08 = 1;
    27: op1_06_inv08 = 1;
    31: op1_06_inv08 = 1;
    32: op1_06_inv08 = 1;
    33: op1_06_inv08 = 1;
    37: op1_06_inv08 = 1;
    38: op1_06_inv08 = 1;
    39: op1_06_inv08 = 1;
    40: op1_06_inv08 = 1;
    42: op1_06_inv08 = 1;
    44: op1_06_inv08 = 1;
    49: op1_06_inv08 = 1;
    51: op1_06_inv08 = 1;
    52: op1_06_inv08 = 1;
    53: op1_06_inv08 = 1;
    54: op1_06_inv08 = 1;
    55: op1_06_inv08 = 1;
    57: op1_06_inv08 = 1;
    58: op1_06_inv08 = 1;
    59: op1_06_inv08 = 1;
    61: op1_06_inv08 = 1;
    65: op1_06_inv08 = 1;
    68: op1_06_inv08 = 1;
    69: op1_06_inv08 = 1;
    71: op1_06_inv08 = 1;
    72: op1_06_inv08 = 1;
    76: op1_06_inv08 = 1;
    78: op1_06_inv08 = 1;
    79: op1_06_inv08 = 1;
    86: op1_06_inv08 = 1;
    87: op1_06_inv08 = 1;
    89: op1_06_inv08 = 1;
    90: op1_06_inv08 = 1;
    91: op1_06_inv08 = 1;
    96: op1_06_inv08 = 1;
    default: op1_06_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in09 = reg_0650;
    5: op1_06_in09 = reg_0451;
    6: op1_06_in09 = reg_0555;
    7: op1_06_in09 = imem07_in[63:60];
    8: op1_06_in09 = reg_0642;
    9: op1_06_in09 = reg_0469;
    10: op1_06_in09 = reg_0109;
    11: op1_06_in09 = reg_0464;
    3: op1_06_in09 = reg_0159;
    12: op1_06_in09 = reg_0068;
    13: op1_06_in09 = reg_0721;
    14: op1_06_in09 = reg_0692;
    15: op1_06_in09 = reg_0015;
    33: op1_06_in09 = reg_0015;
    16: op1_06_in09 = imem05_in[107:104];
    17: op1_06_in09 = imem03_in[7:4];
    18: op1_06_in09 = reg_0605;
    69: op1_06_in09 = reg_0605;
    2: op1_06_in09 = reg_0165;
    19: op1_06_in09 = reg_0325;
    20: op1_06_in09 = reg_0140;
    21: op1_06_in09 = imem02_in[31:28];
    22: op1_06_in09 = imem02_in[47:44];
    23: op1_06_in09 = reg_0468;
    24: op1_06_in09 = reg_0804;
    25: op1_06_in09 = imem06_in[75:72];
    26: op1_06_in09 = reg_0007;
    27: op1_06_in09 = imem05_in[3:0];
    28: op1_06_in09 = imem02_in[99:96];
    29: op1_06_in09 = reg_0351;
    30: op1_06_in09 = reg_0793;
    31: op1_06_in09 = reg_0678;
    32: op1_06_in09 = reg_0245;
    34: op1_06_in09 = imem00_in[103:100];
    36: op1_06_in09 = reg_0670;
    37: op1_06_in09 = reg_0674;
    38: op1_06_in09 = imem02_in[87:84];
    39: op1_06_in09 = imem04_in[115:112];
    40: op1_06_in09 = imem03_in[47:44];
    41: op1_06_in09 = reg_0367;
    42: op1_06_in09 = reg_0210;
    43: op1_06_in09 = reg_0358;
    44: op1_06_in09 = reg_0145;
    45: op1_06_in09 = reg_0635;
    65: op1_06_in09 = reg_0635;
    46: op1_06_in09 = imem02_in[95:92];
    47: op1_06_in09 = reg_0065;
    49: op1_06_in09 = reg_0628;
    50: op1_06_in09 = imem05_in[19:16];
    51: op1_06_in09 = reg_0637;
    52: op1_06_in09 = reg_0552;
    53: op1_06_in09 = reg_0791;
    54: op1_06_in09 = reg_0369;
    55: op1_06_in09 = reg_0238;
    57: op1_06_in09 = reg_0684;
    58: op1_06_in09 = reg_0184;
    59: op1_06_in09 = reg_0424;
    60: op1_06_in09 = reg_0452;
    61: op1_06_in09 = imem02_in[75:72];
    62: op1_06_in09 = reg_0133;
    63: op1_06_in09 = imem06_in[3:0];
    66: op1_06_in09 = reg_0441;
    67: op1_06_in09 = reg_0474;
    68: op1_06_in09 = reg_0545;
    70: op1_06_in09 = reg_0690;
    71: op1_06_in09 = reg_0593;
    72: op1_06_in09 = reg_0710;
    74: op1_06_in09 = reg_0477;
    80: op1_06_in09 = reg_0477;
    75: op1_06_in09 = reg_0527;
    76: op1_06_in09 = reg_0753;
    95: op1_06_in09 = reg_0753;
    77: op1_06_in09 = reg_0564;
    78: op1_06_in09 = reg_0404;
    79: op1_06_in09 = reg_0182;
    82: op1_06_in09 = reg_0616;
    83: op1_06_in09 = reg_0518;
    84: op1_06_in09 = imem07_in[83:80];
    85: op1_06_in09 = reg_0658;
    86: op1_06_in09 = reg_0551;
    87: op1_06_in09 = reg_0401;
    88: op1_06_in09 = imem03_in[55:52];
    89: op1_06_in09 = imem07_in[59:56];
    90: op1_06_in09 = reg_0099;
    91: op1_06_in09 = reg_0183;
    92: op1_06_in09 = reg_0533;
    93: op1_06_in09 = imem02_in[51:48];
    94: op1_06_in09 = reg_0120;
    96: op1_06_in09 = reg_0481;
    default: op1_06_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv09 = 1;
    7: op1_06_inv09 = 1;
    8: op1_06_inv09 = 1;
    9: op1_06_inv09 = 1;
    10: op1_06_inv09 = 1;
    3: op1_06_inv09 = 1;
    14: op1_06_inv09 = 1;
    17: op1_06_inv09 = 1;
    18: op1_06_inv09 = 1;
    2: op1_06_inv09 = 1;
    20: op1_06_inv09 = 1;
    21: op1_06_inv09 = 1;
    23: op1_06_inv09 = 1;
    27: op1_06_inv09 = 1;
    31: op1_06_inv09 = 1;
    36: op1_06_inv09 = 1;
    38: op1_06_inv09 = 1;
    39: op1_06_inv09 = 1;
    40: op1_06_inv09 = 1;
    41: op1_06_inv09 = 1;
    44: op1_06_inv09 = 1;
    45: op1_06_inv09 = 1;
    46: op1_06_inv09 = 1;
    47: op1_06_inv09 = 1;
    50: op1_06_inv09 = 1;
    53: op1_06_inv09 = 1;
    54: op1_06_inv09 = 1;
    55: op1_06_inv09 = 1;
    57: op1_06_inv09 = 1;
    58: op1_06_inv09 = 1;
    59: op1_06_inv09 = 1;
    60: op1_06_inv09 = 1;
    61: op1_06_inv09 = 1;
    62: op1_06_inv09 = 1;
    66: op1_06_inv09 = 1;
    68: op1_06_inv09 = 1;
    71: op1_06_inv09 = 1;
    72: op1_06_inv09 = 1;
    76: op1_06_inv09 = 1;
    78: op1_06_inv09 = 1;
    79: op1_06_inv09 = 1;
    80: op1_06_inv09 = 1;
    82: op1_06_inv09 = 1;
    83: op1_06_inv09 = 1;
    84: op1_06_inv09 = 1;
    87: op1_06_inv09 = 1;
    88: op1_06_inv09 = 1;
    93: op1_06_inv09 = 1;
    94: op1_06_inv09 = 1;
    default: op1_06_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in10 = reg_0637;
    5: op1_06_in10 = reg_0470;
    6: op1_06_in10 = reg_0556;
    7: op1_06_in10 = imem07_in[67:64];
    8: op1_06_in10 = reg_0646;
    9: op1_06_in10 = reg_0476;
    10: op1_06_in10 = reg_0110;
    11: op1_06_in10 = reg_0469;
    74: op1_06_in10 = reg_0469;
    3: op1_06_in10 = reg_0171;
    12: op1_06_in10 = reg_0048;
    13: op1_06_in10 = reg_0703;
    76: op1_06_in10 = reg_0703;
    14: op1_06_in10 = reg_0463;
    15: op1_06_in10 = reg_0016;
    16: op1_06_in10 = imem05_in[111:108];
    17: op1_06_in10 = imem03_in[31:28];
    18: op1_06_in10 = reg_0621;
    2: op1_06_in10 = reg_0185;
    79: op1_06_in10 = reg_0185;
    91: op1_06_in10 = reg_0185;
    19: op1_06_in10 = reg_0354;
    20: op1_06_in10 = imem06_in[3:0];
    21: op1_06_in10 = imem02_in[63:60];
    22: op1_06_in10 = imem02_in[51:48];
    23: op1_06_in10 = reg_0200;
    24: op1_06_in10 = reg_0805;
    25: op1_06_in10 = reg_0614;
    26: op1_06_in10 = reg_0014;
    27: op1_06_in10 = imem05_in[15:12];
    28: op1_06_in10 = imem02_in[107:104];
    29: op1_06_in10 = reg_0743;
    30: op1_06_in10 = reg_0786;
    31: op1_06_in10 = reg_0688;
    85: op1_06_in10 = reg_0688;
    32: op1_06_in10 = reg_0111;
    33: op1_06_in10 = reg_0799;
    34: op1_06_in10 = reg_0681;
    36: op1_06_in10 = reg_0690;
    37: op1_06_in10 = reg_0671;
    38: op1_06_in10 = reg_0642;
    39: op1_06_in10 = reg_0542;
    40: op1_06_in10 = imem03_in[83:80];
    41: op1_06_in10 = imem07_in[27:24];
    55: op1_06_in10 = imem07_in[27:24];
    42: op1_06_in10 = reg_0187;
    43: op1_06_in10 = reg_0360;
    44: op1_06_in10 = reg_0142;
    45: op1_06_in10 = reg_0434;
    65: op1_06_in10 = reg_0434;
    46: op1_06_in10 = imem02_in[115:112];
    47: op1_06_in10 = reg_0519;
    49: op1_06_in10 = reg_0624;
    50: op1_06_in10 = imem05_in[23:20];
    51: op1_06_in10 = imem02_in[3:0];
    52: op1_06_in10 = reg_0043;
    53: op1_06_in10 = reg_0798;
    54: op1_06_in10 = reg_0377;
    57: op1_06_in10 = reg_0691;
    59: op1_06_in10 = reg_0123;
    60: op1_06_in10 = reg_0478;
    61: op1_06_in10 = imem02_in[79:76];
    62: op1_06_in10 = reg_0138;
    63: op1_06_in10 = imem06_in[87:84];
    66: op1_06_in10 = reg_0436;
    67: op1_06_in10 = reg_0471;
    68: op1_06_in10 = reg_0316;
    69: op1_06_in10 = reg_0618;
    70: op1_06_in10 = reg_0758;
    71: op1_06_in10 = reg_0035;
    72: op1_06_in10 = reg_0726;
    75: op1_06_in10 = reg_0518;
    77: op1_06_in10 = reg_0368;
    78: op1_06_in10 = reg_0293;
    80: op1_06_in10 = reg_0460;
    82: op1_06_in10 = reg_0297;
    83: op1_06_in10 = reg_0055;
    84: op1_06_in10 = reg_0391;
    86: op1_06_in10 = reg_0331;
    87: op1_06_in10 = reg_0578;
    88: op1_06_in10 = imem03_in[123:120];
    89: op1_06_in10 = imem07_in[111:108];
    90: op1_06_in10 = reg_0228;
    92: op1_06_in10 = reg_0639;
    93: op1_06_in10 = imem02_in[75:72];
    94: op1_06_in10 = reg_0660;
    95: op1_06_in10 = reg_0075;
    96: op1_06_in10 = reg_0473;
    default: op1_06_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv10 = 1;
    5: op1_06_inv10 = 1;
    7: op1_06_inv10 = 1;
    10: op1_06_inv10 = 1;
    11: op1_06_inv10 = 1;
    3: op1_06_inv10 = 1;
    12: op1_06_inv10 = 1;
    13: op1_06_inv10 = 1;
    14: op1_06_inv10 = 1;
    15: op1_06_inv10 = 1;
    19: op1_06_inv10 = 1;
    20: op1_06_inv10 = 1;
    21: op1_06_inv10 = 1;
    27: op1_06_inv10 = 1;
    28: op1_06_inv10 = 1;
    29: op1_06_inv10 = 1;
    31: op1_06_inv10 = 1;
    32: op1_06_inv10 = 1;
    33: op1_06_inv10 = 1;
    37: op1_06_inv10 = 1;
    39: op1_06_inv10 = 1;
    41: op1_06_inv10 = 1;
    43: op1_06_inv10 = 1;
    45: op1_06_inv10 = 1;
    47: op1_06_inv10 = 1;
    53: op1_06_inv10 = 1;
    54: op1_06_inv10 = 1;
    55: op1_06_inv10 = 1;
    59: op1_06_inv10 = 1;
    61: op1_06_inv10 = 1;
    62: op1_06_inv10 = 1;
    68: op1_06_inv10 = 1;
    69: op1_06_inv10 = 1;
    71: op1_06_inv10 = 1;
    72: op1_06_inv10 = 1;
    74: op1_06_inv10 = 1;
    75: op1_06_inv10 = 1;
    83: op1_06_inv10 = 1;
    84: op1_06_inv10 = 1;
    89: op1_06_inv10 = 1;
    90: op1_06_inv10 = 1;
    91: op1_06_inv10 = 1;
    92: op1_06_inv10 = 1;
    93: op1_06_inv10 = 1;
    94: op1_06_inv10 = 1;
    95: op1_06_inv10 = 1;
    default: op1_06_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in11 = reg_0660;
    21: op1_06_in11 = reg_0660;
    5: op1_06_in11 = reg_0208;
    23: op1_06_in11 = reg_0208;
    6: op1_06_in11 = reg_0304;
    7: op1_06_in11 = imem07_in[75:72];
    8: op1_06_in11 = reg_0661;
    9: op1_06_in11 = reg_0198;
    10: op1_06_in11 = imem02_in[47:44];
    11: op1_06_in11 = reg_0460;
    12: op1_06_in11 = reg_0050;
    13: op1_06_in11 = reg_0712;
    72: op1_06_in11 = reg_0712;
    14: op1_06_in11 = reg_0477;
    15: op1_06_in11 = reg_0810;
    33: op1_06_in11 = reg_0810;
    16: op1_06_in11 = reg_0792;
    17: op1_06_in11 = imem03_in[39:36];
    18: op1_06_in11 = reg_0619;
    19: op1_06_in11 = reg_0345;
    95: op1_06_in11 = reg_0345;
    20: op1_06_in11 = imem06_in[15:12];
    22: op1_06_in11 = imem02_in[111:108];
    24: op1_06_in11 = reg_0015;
    25: op1_06_in11 = reg_0613;
    26: op1_06_in11 = reg_0805;
    27: op1_06_in11 = imem05_in[31:28];
    28: op1_06_in11 = reg_0658;
    29: op1_06_in11 = reg_0532;
    30: op1_06_in11 = reg_0737;
    31: op1_06_in11 = reg_0687;
    32: op1_06_in11 = reg_0116;
    34: op1_06_in11 = reg_0696;
    36: op1_06_in11 = reg_0699;
    37: op1_06_in11 = reg_0668;
    38: op1_06_in11 = reg_0645;
    39: op1_06_in11 = reg_0043;
    40: op1_06_in11 = imem03_in[99:96];
    41: op1_06_in11 = imem07_in[79:76];
    42: op1_06_in11 = reg_0211;
    43: op1_06_in11 = reg_0324;
    44: op1_06_in11 = reg_0143;
    45: op1_06_in11 = reg_0442;
    46: op1_06_in11 = reg_0639;
    47: op1_06_in11 = reg_0549;
    49: op1_06_in11 = reg_0606;
    50: op1_06_in11 = imem05_in[63:60];
    51: op1_06_in11 = imem02_in[35:32];
    52: op1_06_in11 = reg_0060;
    53: op1_06_in11 = reg_0488;
    54: op1_06_in11 = reg_0409;
    55: op1_06_in11 = imem07_in[51:48];
    57: op1_06_in11 = reg_0758;
    59: op1_06_in11 = reg_0104;
    60: op1_06_in11 = reg_0214;
    61: op1_06_in11 = imem02_in[115:112];
    62: op1_06_in11 = imem06_in[91:88];
    63: op1_06_in11 = reg_0299;
    65: op1_06_in11 = reg_0440;
    66: op1_06_in11 = reg_0636;
    67: op1_06_in11 = reg_0210;
    68: op1_06_in11 = reg_0087;
    69: op1_06_in11 = reg_0031;
    70: op1_06_in11 = reg_0688;
    71: op1_06_in11 = reg_0515;
    74: op1_06_in11 = reg_0468;
    75: op1_06_in11 = reg_0080;
    76: op1_06_in11 = reg_0138;
    77: op1_06_in11 = reg_0562;
    78: op1_06_in11 = reg_0401;
    80: op1_06_in11 = reg_0473;
    82: op1_06_in11 = reg_0627;
    83: op1_06_in11 = reg_0117;
    84: op1_06_in11 = reg_0167;
    85: op1_06_in11 = reg_0465;
    86: op1_06_in11 = reg_0516;
    87: op1_06_in11 = reg_0654;
    88: op1_06_in11 = imem03_in[127:124];
    89: op1_06_in11 = reg_0784;
    90: op1_06_in11 = reg_0141;
    92: op1_06_in11 = reg_0498;
    93: op1_06_in11 = imem02_in[79:76];
    94: op1_06_in11 = reg_0669;
    96: op1_06_in11 = reg_0474;
    default: op1_06_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv11 = 1;
    7: op1_06_inv11 = 1;
    8: op1_06_inv11 = 1;
    10: op1_06_inv11 = 1;
    14: op1_06_inv11 = 1;
    16: op1_06_inv11 = 1;
    18: op1_06_inv11 = 1;
    21: op1_06_inv11 = 1;
    22: op1_06_inv11 = 1;
    23: op1_06_inv11 = 1;
    25: op1_06_inv11 = 1;
    29: op1_06_inv11 = 1;
    32: op1_06_inv11 = 1;
    36: op1_06_inv11 = 1;
    38: op1_06_inv11 = 1;
    39: op1_06_inv11 = 1;
    40: op1_06_inv11 = 1;
    43: op1_06_inv11 = 1;
    47: op1_06_inv11 = 1;
    49: op1_06_inv11 = 1;
    50: op1_06_inv11 = 1;
    52: op1_06_inv11 = 1;
    54: op1_06_inv11 = 1;
    55: op1_06_inv11 = 1;
    57: op1_06_inv11 = 1;
    59: op1_06_inv11 = 1;
    60: op1_06_inv11 = 1;
    63: op1_06_inv11 = 1;
    65: op1_06_inv11 = 1;
    67: op1_06_inv11 = 1;
    69: op1_06_inv11 = 1;
    76: op1_06_inv11 = 1;
    80: op1_06_inv11 = 1;
    82: op1_06_inv11 = 1;
    88: op1_06_inv11 = 1;
    89: op1_06_inv11 = 1;
    92: op1_06_inv11 = 1;
    95: op1_06_inv11 = 1;
    default: op1_06_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in12 = reg_0661;
    5: op1_06_in12 = reg_0210;
    60: op1_06_in12 = reg_0210;
    6: op1_06_in12 = reg_0294;
    7: op1_06_in12 = imem07_in[91:88];
    8: op1_06_in12 = reg_0648;
    9: op1_06_in12 = reg_0738;
    10: op1_06_in12 = imem02_in[55:52];
    11: op1_06_in12 = reg_0481;
    12: op1_06_in12 = reg_0792;
    13: op1_06_in12 = reg_0715;
    14: op1_06_in12 = reg_0469;
    85: op1_06_in12 = reg_0469;
    15: op1_06_in12 = imem04_in[3:0];
    16: op1_06_in12 = reg_0483;
    17: op1_06_in12 = imem03_in[79:76];
    18: op1_06_in12 = reg_0615;
    19: op1_06_in12 = reg_0355;
    20: op1_06_in12 = imem06_in[35:32];
    21: op1_06_in12 = reg_0656;
    22: op1_06_in12 = imem02_in[115:112];
    23: op1_06_in12 = reg_0207;
    24: op1_06_in12 = reg_0016;
    25: op1_06_in12 = reg_0605;
    26: op1_06_in12 = reg_0799;
    27: op1_06_in12 = imem05_in[39:36];
    28: op1_06_in12 = reg_0664;
    29: op1_06_in12 = imem03_in[15:12];
    30: op1_06_in12 = reg_0276;
    31: op1_06_in12 = reg_0454;
    32: op1_06_in12 = reg_0114;
    33: op1_06_in12 = imem04_in[7:4];
    34: op1_06_in12 = reg_0677;
    36: op1_06_in12 = reg_0463;
    37: op1_06_in12 = reg_0669;
    38: op1_06_in12 = reg_0651;
    39: op1_06_in12 = reg_0536;
    40: op1_06_in12 = imem03_in[127:124];
    41: op1_06_in12 = imem07_in[115:112];
    42: op1_06_in12 = reg_0186;
    43: op1_06_in12 = reg_0353;
    76: op1_06_in12 = reg_0353;
    44: op1_06_in12 = reg_0140;
    45: op1_06_in12 = reg_0180;
    46: op1_06_in12 = reg_0665;
    47: op1_06_in12 = imem05_in[31:28];
    49: op1_06_in12 = reg_0622;
    50: op1_06_in12 = imem05_in[71:68];
    51: op1_06_in12 = imem02_in[79:76];
    52: op1_06_in12 = reg_0057;
    53: op1_06_in12 = reg_0788;
    54: op1_06_in12 = reg_0821;
    55: op1_06_in12 = imem07_in[59:56];
    57: op1_06_in12 = reg_0476;
    59: op1_06_in12 = reg_0120;
    61: op1_06_in12 = reg_0666;
    62: op1_06_in12 = imem06_in[123:120];
    63: op1_06_in12 = reg_0577;
    65: op1_06_in12 = reg_0448;
    66: op1_06_in12 = reg_0067;
    67: op1_06_in12 = reg_0194;
    68: op1_06_in12 = reg_0055;
    69: op1_06_in12 = reg_0580;
    70: op1_06_in12 = reg_0247;
    71: op1_06_in12 = reg_0039;
    72: op1_06_in12 = reg_0724;
    74: op1_06_in12 = reg_0479;
    80: op1_06_in12 = reg_0479;
    75: op1_06_in12 = reg_0096;
    77: op1_06_in12 = reg_0398;
    78: op1_06_in12 = reg_0031;
    82: op1_06_in12 = reg_0679;
    83: op1_06_in12 = imem02_in[19:16];
    84: op1_06_in12 = reg_0713;
    86: op1_06_in12 = reg_0556;
    87: op1_06_in12 = reg_0307;
    88: op1_06_in12 = reg_0010;
    89: op1_06_in12 = reg_0061;
    90: op1_06_in12 = reg_0325;
    92: op1_06_in12 = reg_0485;
    93: op1_06_in12 = imem02_in[103:100];
    94: op1_06_in12 = reg_0601;
    95: op1_06_in12 = reg_0361;
    96: op1_06_in12 = reg_0478;
    default: op1_06_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv12 = 1;
    6: op1_06_inv12 = 1;
    7: op1_06_inv12 = 1;
    8: op1_06_inv12 = 1;
    12: op1_06_inv12 = 1;
    16: op1_06_inv12 = 1;
    18: op1_06_inv12 = 1;
    22: op1_06_inv12 = 1;
    23: op1_06_inv12 = 1;
    24: op1_06_inv12 = 1;
    27: op1_06_inv12 = 1;
    28: op1_06_inv12 = 1;
    30: op1_06_inv12 = 1;
    34: op1_06_inv12 = 1;
    37: op1_06_inv12 = 1;
    39: op1_06_inv12 = 1;
    40: op1_06_inv12 = 1;
    42: op1_06_inv12 = 1;
    44: op1_06_inv12 = 1;
    53: op1_06_inv12 = 1;
    59: op1_06_inv12 = 1;
    62: op1_06_inv12 = 1;
    65: op1_06_inv12 = 1;
    66: op1_06_inv12 = 1;
    67: op1_06_inv12 = 1;
    72: op1_06_inv12 = 1;
    74: op1_06_inv12 = 1;
    80: op1_06_inv12 = 1;
    85: op1_06_inv12 = 1;
    89: op1_06_inv12 = 1;
    92: op1_06_inv12 = 1;
    94: op1_06_inv12 = 1;
    default: op1_06_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in13 = reg_0639;
    5: op1_06_in13 = reg_0204;
    6: op1_06_in13 = reg_0277;
    7: op1_06_in13 = imem07_in[95:92];
    8: op1_06_in13 = reg_0638;
    9: op1_06_in13 = reg_0497;
    10: op1_06_in13 = imem02_in[63:60];
    11: op1_06_in13 = reg_0473;
    12: op1_06_in13 = reg_0796;
    13: op1_06_in13 = reg_0701;
    14: op1_06_in13 = reg_0466;
    85: op1_06_in13 = reg_0466;
    15: op1_06_in13 = imem04_in[75:72];
    16: op1_06_in13 = reg_0785;
    17: op1_06_in13 = imem03_in[115:112];
    18: op1_06_in13 = reg_0601;
    19: op1_06_in13 = reg_0314;
    20: op1_06_in13 = imem06_in[39:36];
    21: op1_06_in13 = reg_0641;
    22: op1_06_in13 = imem02_in[123:120];
    23: op1_06_in13 = reg_0211;
    74: op1_06_in13 = reg_0211;
    24: op1_06_in13 = imem04_in[3:0];
    25: op1_06_in13 = reg_0616;
    26: op1_06_in13 = reg_0004;
    27: op1_06_in13 = imem05_in[63:60];
    28: op1_06_in13 = reg_0647;
    29: op1_06_in13 = imem03_in[43:40];
    30: op1_06_in13 = reg_0282;
    31: op1_06_in13 = reg_0469;
    32: op1_06_in13 = reg_0100;
    33: op1_06_in13 = imem04_in[11:8];
    34: op1_06_in13 = reg_0691;
    36: op1_06_in13 = reg_0450;
    37: op1_06_in13 = reg_0465;
    38: op1_06_in13 = reg_0358;
    39: op1_06_in13 = reg_0556;
    68: op1_06_in13 = reg_0556;
    40: op1_06_in13 = reg_0602;
    41: op1_06_in13 = reg_0722;
    42: op1_06_in13 = reg_0201;
    43: op1_06_in13 = reg_0541;
    44: op1_06_in13 = imem06_in[31:28];
    45: op1_06_in13 = reg_0167;
    46: op1_06_in13 = reg_0341;
    92: op1_06_in13 = reg_0341;
    47: op1_06_in13 = imem05_in[67:64];
    49: op1_06_in13 = reg_0369;
    50: op1_06_in13 = imem05_in[87:84];
    51: op1_06_in13 = imem02_in[91:88];
    52: op1_06_in13 = reg_0079;
    53: op1_06_in13 = reg_0789;
    54: op1_06_in13 = reg_0242;
    55: op1_06_in13 = imem07_in[99:96];
    57: op1_06_in13 = reg_0480;
    59: op1_06_in13 = reg_0672;
    60: op1_06_in13 = reg_0188;
    61: op1_06_in13 = reg_0637;
    62: op1_06_in13 = reg_0625;
    63: op1_06_in13 = reg_0624;
    65: op1_06_in13 = reg_0268;
    66: op1_06_in13 = reg_0444;
    67: op1_06_in13 = imem01_in[15:12];
    69: op1_06_in13 = reg_0700;
    70: op1_06_in13 = reg_0464;
    71: op1_06_in13 = reg_0787;
    72: op1_06_in13 = reg_0713;
    75: op1_06_in13 = reg_0539;
    76: op1_06_in13 = reg_0351;
    77: op1_06_in13 = reg_0496;
    78: op1_06_in13 = reg_0408;
    80: op1_06_in13 = reg_0186;
    82: op1_06_in13 = reg_0301;
    83: op1_06_in13 = imem02_in[35:32];
    84: op1_06_in13 = reg_0064;
    86: op1_06_in13 = reg_0174;
    87: op1_06_in13 = reg_0748;
    88: op1_06_in13 = reg_0507;
    89: op1_06_in13 = reg_0445;
    93: op1_06_in13 = imem02_in[111:108];
    94: op1_06_in13 = reg_0674;
    95: op1_06_in13 = reg_0353;
    96: op1_06_in13 = reg_0212;
    default: op1_06_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv13 = 1;
    5: op1_06_inv13 = 1;
    7: op1_06_inv13 = 1;
    10: op1_06_inv13 = 1;
    13: op1_06_inv13 = 1;
    18: op1_06_inv13 = 1;
    19: op1_06_inv13 = 1;
    20: op1_06_inv13 = 1;
    22: op1_06_inv13 = 1;
    23: op1_06_inv13 = 1;
    24: op1_06_inv13 = 1;
    28: op1_06_inv13 = 1;
    30: op1_06_inv13 = 1;
    34: op1_06_inv13 = 1;
    37: op1_06_inv13 = 1;
    38: op1_06_inv13 = 1;
    39: op1_06_inv13 = 1;
    40: op1_06_inv13 = 1;
    41: op1_06_inv13 = 1;
    46: op1_06_inv13 = 1;
    49: op1_06_inv13 = 1;
    51: op1_06_inv13 = 1;
    52: op1_06_inv13 = 1;
    54: op1_06_inv13 = 1;
    55: op1_06_inv13 = 1;
    57: op1_06_inv13 = 1;
    63: op1_06_inv13 = 1;
    65: op1_06_inv13 = 1;
    66: op1_06_inv13 = 1;
    68: op1_06_inv13 = 1;
    72: op1_06_inv13 = 1;
    74: op1_06_inv13 = 1;
    75: op1_06_inv13 = 1;
    76: op1_06_inv13 = 1;
    77: op1_06_inv13 = 1;
    82: op1_06_inv13 = 1;
    84: op1_06_inv13 = 1;
    85: op1_06_inv13 = 1;
    87: op1_06_inv13 = 1;
    89: op1_06_inv13 = 1;
    93: op1_06_inv13 = 1;
    94: op1_06_inv13 = 1;
    96: op1_06_inv13 = 1;
    default: op1_06_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in14 = reg_0640;
    5: op1_06_in14 = reg_0203;
    6: op1_06_in14 = reg_0059;
    7: op1_06_in14 = imem07_in[111:108];
    55: op1_06_in14 = imem07_in[111:108];
    8: op1_06_in14 = reg_0659;
    9: op1_06_in14 = reg_0499;
    10: op1_06_in14 = reg_0642;
    11: op1_06_in14 = reg_0467;
    12: op1_06_in14 = reg_0490;
    88: op1_06_in14 = reg_0490;
    13: op1_06_in14 = reg_0700;
    14: op1_06_in14 = reg_0468;
    15: op1_06_in14 = imem04_in[99:96];
    16: op1_06_in14 = reg_0495;
    17: op1_06_in14 = reg_0602;
    18: op1_06_in14 = reg_0402;
    19: op1_06_in14 = reg_0096;
    20: op1_06_in14 = reg_0628;
    21: op1_06_in14 = reg_0345;
    22: op1_06_in14 = reg_0666;
    23: op1_06_in14 = imem01_in[23:20];
    24: op1_06_in14 = imem04_in[15:12];
    25: op1_06_in14 = reg_0619;
    26: op1_06_in14 = imem04_in[71:68];
    27: op1_06_in14 = imem05_in[115:112];
    28: op1_06_in14 = reg_0667;
    29: op1_06_in14 = reg_0598;
    30: op1_06_in14 = reg_0269;
    31: op1_06_in14 = reg_0472;
    32: op1_06_in14 = imem02_in[11:8];
    33: op1_06_in14 = imem04_in[19:16];
    34: op1_06_in14 = reg_0688;
    36: op1_06_in14 = reg_0455;
    37: op1_06_in14 = reg_0450;
    38: op1_06_in14 = reg_0229;
    39: op1_06_in14 = reg_0301;
    40: op1_06_in14 = reg_0586;
    41: op1_06_in14 = reg_0719;
    42: op1_06_in14 = reg_0212;
    43: op1_06_in14 = reg_0080;
    44: op1_06_in14 = imem06_in[79:76];
    45: op1_06_in14 = reg_0160;
    46: op1_06_in14 = reg_0361;
    47: op1_06_in14 = imem05_in[71:68];
    49: op1_06_in14 = reg_0577;
    50: op1_06_in14 = imem05_in[111:108];
    51: op1_06_in14 = imem02_in[127:124];
    52: op1_06_in14 = reg_0076;
    53: op1_06_in14 = reg_0494;
    54: op1_06_in14 = reg_0812;
    57: op1_06_in14 = reg_0214;
    59: op1_06_in14 = reg_0675;
    60: op1_06_in14 = reg_0213;
    61: op1_06_in14 = reg_0661;
    62: op1_06_in14 = reg_0346;
    63: op1_06_in14 = reg_0298;
    65: op1_06_in14 = reg_0162;
    66: op1_06_in14 = reg_0442;
    67: op1_06_in14 = reg_0735;
    68: op1_06_in14 = reg_0305;
    69: op1_06_in14 = reg_0813;
    70: op1_06_in14 = reg_0461;
    71: op1_06_in14 = imem07_in[11:8];
    72: op1_06_in14 = reg_0636;
    74: op1_06_in14 = reg_0201;
    75: op1_06_in14 = reg_0757;
    76: op1_06_in14 = reg_0514;
    77: op1_06_in14 = reg_0637;
    78: op1_06_in14 = reg_0375;
    80: op1_06_in14 = reg_0198;
    82: op1_06_in14 = reg_0513;
    83: op1_06_in14 = imem02_in[39:36];
    84: op1_06_in14 = reg_0253;
    85: op1_06_in14 = reg_0475;
    86: op1_06_in14 = reg_0283;
    87: op1_06_in14 = reg_0763;
    89: op1_06_in14 = reg_0439;
    92: op1_06_in14 = reg_0359;
    93: op1_06_in14 = imem02_in[115:112];
    94: op1_06_in14 = reg_0678;
    95: op1_06_in14 = reg_0566;
    96: op1_06_in14 = imem01_in[11:8];
    default: op1_06_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv14 = 1;
    6: op1_06_inv14 = 1;
    10: op1_06_inv14 = 1;
    14: op1_06_inv14 = 1;
    15: op1_06_inv14 = 1;
    18: op1_06_inv14 = 1;
    21: op1_06_inv14 = 1;
    23: op1_06_inv14 = 1;
    25: op1_06_inv14 = 1;
    28: op1_06_inv14 = 1;
    31: op1_06_inv14 = 1;
    32: op1_06_inv14 = 1;
    34: op1_06_inv14 = 1;
    41: op1_06_inv14 = 1;
    42: op1_06_inv14 = 1;
    43: op1_06_inv14 = 1;
    44: op1_06_inv14 = 1;
    47: op1_06_inv14 = 1;
    51: op1_06_inv14 = 1;
    55: op1_06_inv14 = 1;
    59: op1_06_inv14 = 1;
    60: op1_06_inv14 = 1;
    61: op1_06_inv14 = 1;
    66: op1_06_inv14 = 1;
    74: op1_06_inv14 = 1;
    75: op1_06_inv14 = 1;
    77: op1_06_inv14 = 1;
    78: op1_06_inv14 = 1;
    80: op1_06_inv14 = 1;
    82: op1_06_inv14 = 1;
    83: op1_06_inv14 = 1;
    84: op1_06_inv14 = 1;
    86: op1_06_inv14 = 1;
    87: op1_06_inv14 = 1;
    88: op1_06_inv14 = 1;
    89: op1_06_inv14 = 1;
    93: op1_06_inv14 = 1;
    94: op1_06_inv14 = 1;
    95: op1_06_inv14 = 1;
    96: op1_06_inv14 = 1;
    default: op1_06_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in15 = reg_0641;
    5: op1_06_in15 = reg_0213;
    80: op1_06_in15 = reg_0213;
    6: op1_06_in15 = reg_0062;
    7: op1_06_in15 = reg_0723;
    8: op1_06_in15 = reg_0636;
    9: op1_06_in15 = reg_0230;
    10: op1_06_in15 = reg_0654;
    11: op1_06_in15 = reg_0474;
    12: op1_06_in15 = reg_0784;
    13: op1_06_in15 = reg_0441;
    14: op1_06_in15 = reg_0459;
    15: op1_06_in15 = reg_0544;
    16: op1_06_in15 = reg_0485;
    17: op1_06_in15 = reg_0591;
    18: op1_06_in15 = reg_0332;
    19: op1_06_in15 = reg_0097;
    20: op1_06_in15 = reg_0632;
    21: op1_06_in15 = reg_0318;
    22: op1_06_in15 = reg_0646;
    23: op1_06_in15 = imem01_in[107:104];
    24: op1_06_in15 = imem04_in[59:56];
    25: op1_06_in15 = reg_0601;
    26: op1_06_in15 = imem04_in[79:76];
    27: op1_06_in15 = reg_0798;
    28: op1_06_in15 = reg_0364;
    29: op1_06_in15 = reg_0582;
    30: op1_06_in15 = reg_0142;
    31: op1_06_in15 = reg_0189;
    32: op1_06_in15 = imem02_in[35:32];
    33: op1_06_in15 = imem04_in[23:20];
    34: op1_06_in15 = reg_0453;
    36: op1_06_in15 = reg_0466;
    37: op1_06_in15 = reg_0208;
    57: op1_06_in15 = reg_0208;
    38: op1_06_in15 = reg_0341;
    39: op1_06_in15 = reg_0273;
    40: op1_06_in15 = reg_0566;
    41: op1_06_in15 = reg_0710;
    42: op1_06_in15 = reg_0190;
    43: op1_06_in15 = reg_0095;
    92: op1_06_in15 = reg_0095;
    44: op1_06_in15 = imem06_in[87:84];
    45: op1_06_in15 = reg_0183;
    46: op1_06_in15 = reg_0351;
    47: op1_06_in15 = imem05_in[79:76];
    49: op1_06_in15 = reg_0405;
    50: op1_06_in15 = imem05_in[119:116];
    51: op1_06_in15 = reg_0518;
    52: op1_06_in15 = reg_0071;
    53: op1_06_in15 = reg_0787;
    54: op1_06_in15 = reg_0372;
    55: op1_06_in15 = imem07_in[123:120];
    59: op1_06_in15 = reg_0669;
    60: op1_06_in15 = reg_0205;
    61: op1_06_in15 = reg_0344;
    62: op1_06_in15 = reg_0609;
    63: op1_06_in15 = reg_0578;
    66: op1_06_in15 = reg_0267;
    67: op1_06_in15 = reg_0733;
    68: op1_06_in15 = reg_0280;
    86: op1_06_in15 = reg_0280;
    69: op1_06_in15 = reg_0752;
    70: op1_06_in15 = reg_0473;
    71: op1_06_in15 = imem07_in[27:24];
    72: op1_06_in15 = reg_0445;
    74: op1_06_in15 = imem01_in[39:36];
    75: op1_06_in15 = imem03_in[7:4];
    76: op1_06_in15 = reg_0323;
    77: op1_06_in15 = reg_0396;
    78: op1_06_in15 = reg_0764;
    82: op1_06_in15 = reg_0640;
    83: op1_06_in15 = imem02_in[71:68];
    84: op1_06_in15 = reg_0295;
    85: op1_06_in15 = reg_0472;
    87: op1_06_in15 = reg_0025;
    88: op1_06_in15 = reg_0549;
    89: op1_06_in15 = reg_0434;
    93: op1_06_in15 = reg_0642;
    94: op1_06_in15 = imem02_in[103:100];
    95: op1_06_in15 = reg_0514;
    96: op1_06_in15 = imem01_in[67:64];
    default: op1_06_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv15 = 1;
    8: op1_06_inv15 = 1;
    9: op1_06_inv15 = 1;
    11: op1_06_inv15 = 1;
    12: op1_06_inv15 = 1;
    14: op1_06_inv15 = 1;
    19: op1_06_inv15 = 1;
    20: op1_06_inv15 = 1;
    24: op1_06_inv15 = 1;
    25: op1_06_inv15 = 1;
    26: op1_06_inv15 = 1;
    27: op1_06_inv15 = 1;
    28: op1_06_inv15 = 1;
    31: op1_06_inv15 = 1;
    36: op1_06_inv15 = 1;
    37: op1_06_inv15 = 1;
    39: op1_06_inv15 = 1;
    40: op1_06_inv15 = 1;
    42: op1_06_inv15 = 1;
    43: op1_06_inv15 = 1;
    46: op1_06_inv15 = 1;
    47: op1_06_inv15 = 1;
    49: op1_06_inv15 = 1;
    50: op1_06_inv15 = 1;
    51: op1_06_inv15 = 1;
    52: op1_06_inv15 = 1;
    53: op1_06_inv15 = 1;
    55: op1_06_inv15 = 1;
    57: op1_06_inv15 = 1;
    59: op1_06_inv15 = 1;
    62: op1_06_inv15 = 1;
    70: op1_06_inv15 = 1;
    72: op1_06_inv15 = 1;
    75: op1_06_inv15 = 1;
    76: op1_06_inv15 = 1;
    77: op1_06_inv15 = 1;
    78: op1_06_inv15 = 1;
    80: op1_06_inv15 = 1;
    87: op1_06_inv15 = 1;
    88: op1_06_inv15 = 1;
    89: op1_06_inv15 = 1;
    94: op1_06_inv15 = 1;
    96: op1_06_inv15 = 1;
    default: op1_06_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in16 = reg_0333;
    5: op1_06_in16 = reg_0202;
    42: op1_06_in16 = reg_0202;
    6: op1_06_in16 = reg_0058;
    7: op1_06_in16 = reg_0430;
    8: op1_06_in16 = reg_0358;
    9: op1_06_in16 = reg_0736;
    12: op1_06_in16 = reg_0736;
    53: op1_06_in16 = reg_0736;
    10: op1_06_in16 = reg_0646;
    11: op1_06_in16 = reg_0471;
    13: op1_06_in16 = reg_0422;
    14: op1_06_in16 = reg_0204;
    15: op1_06_in16 = reg_0536;
    16: op1_06_in16 = reg_0787;
    17: op1_06_in16 = reg_0570;
    18: op1_06_in16 = reg_0372;
    19: op1_06_in16 = imem03_in[7:4];
    20: op1_06_in16 = reg_0402;
    21: op1_06_in16 = reg_0330;
    22: op1_06_in16 = reg_0648;
    23: op1_06_in16 = imem01_in[115:112];
    24: op1_06_in16 = imem04_in[67:64];
    25: op1_06_in16 = reg_0379;
    26: op1_06_in16 = imem04_in[111:108];
    27: op1_06_in16 = reg_0485;
    28: op1_06_in16 = reg_0359;
    29: op1_06_in16 = reg_0596;
    30: op1_06_in16 = reg_0139;
    31: op1_06_in16 = reg_0193;
    32: op1_06_in16 = imem02_in[43:40];
    33: op1_06_in16 = imem04_in[35:32];
    34: op1_06_in16 = reg_0451;
    36: op1_06_in16 = reg_0459;
    37: op1_06_in16 = reg_0203;
    38: op1_06_in16 = reg_0345;
    61: op1_06_in16 = reg_0345;
    39: op1_06_in16 = reg_0268;
    40: op1_06_in16 = reg_0594;
    41: op1_06_in16 = reg_0731;
    43: op1_06_in16 = reg_0096;
    51: op1_06_in16 = reg_0096;
    44: op1_06_in16 = imem06_in[107:104];
    45: op1_06_in16 = reg_0177;
    46: op1_06_in16 = reg_0347;
    47: op1_06_in16 = imem05_in[83:80];
    49: op1_06_in16 = reg_0775;
    50: op1_06_in16 = reg_0482;
    52: op1_06_in16 = reg_0292;
    54: op1_06_in16 = reg_0819;
    55: op1_06_in16 = reg_0720;
    57: op1_06_in16 = reg_0195;
    59: op1_06_in16 = reg_0678;
    60: op1_06_in16 = reg_0190;
    62: op1_06_in16 = reg_0401;
    63: op1_06_in16 = reg_0377;
    66: op1_06_in16 = reg_0448;
    67: op1_06_in16 = reg_0759;
    68: op1_06_in16 = reg_0076;
    69: op1_06_in16 = reg_0632;
    70: op1_06_in16 = reg_0470;
    71: op1_06_in16 = imem07_in[43:40];
    72: op1_06_in16 = reg_0181;
    74: op1_06_in16 = imem01_in[59:56];
    75: op1_06_in16 = imem03_in[39:36];
    76: op1_06_in16 = reg_0541;
    77: op1_06_in16 = reg_0006;
    78: op1_06_in16 = reg_0515;
    80: op1_06_in16 = reg_0196;
    82: op1_06_in16 = reg_0416;
    83: op1_06_in16 = imem02_in[111:108];
    94: op1_06_in16 = imem02_in[111:108];
    84: op1_06_in16 = reg_0436;
    85: op1_06_in16 = reg_0456;
    86: op1_06_in16 = reg_0074;
    87: op1_06_in16 = reg_0663;
    88: op1_06_in16 = reg_0496;
    89: op1_06_in16 = reg_0440;
    92: op1_06_in16 = reg_0255;
    93: op1_06_in16 = reg_0088;
    95: op1_06_in16 = reg_0109;
    96: op1_06_in16 = imem01_in[71:68];
    default: op1_06_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv16 = 1;
    6: op1_06_inv16 = 1;
    7: op1_06_inv16 = 1;
    10: op1_06_inv16 = 1;
    11: op1_06_inv16 = 1;
    13: op1_06_inv16 = 1;
    15: op1_06_inv16 = 1;
    21: op1_06_inv16 = 1;
    23: op1_06_inv16 = 1;
    24: op1_06_inv16 = 1;
    36: op1_06_inv16 = 1;
    37: op1_06_inv16 = 1;
    40: op1_06_inv16 = 1;
    42: op1_06_inv16 = 1;
    44: op1_06_inv16 = 1;
    45: op1_06_inv16 = 1;
    46: op1_06_inv16 = 1;
    51: op1_06_inv16 = 1;
    54: op1_06_inv16 = 1;
    55: op1_06_inv16 = 1;
    57: op1_06_inv16 = 1;
    59: op1_06_inv16 = 1;
    61: op1_06_inv16 = 1;
    70: op1_06_inv16 = 1;
    77: op1_06_inv16 = 1;
    78: op1_06_inv16 = 1;
    82: op1_06_inv16 = 1;
    83: op1_06_inv16 = 1;
    85: op1_06_inv16 = 1;
    92: op1_06_inv16 = 1;
    93: op1_06_inv16 = 1;
    96: op1_06_inv16 = 1;
    default: op1_06_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in17 = reg_0345;
    5: op1_06_in17 = imem01_in[35:32];
    6: op1_06_in17 = reg_0066;
    7: op1_06_in17 = reg_0445;
    8: op1_06_in17 = reg_0364;
    9: op1_06_in17 = reg_0224;
    10: op1_06_in17 = reg_0656;
    11: op1_06_in17 = reg_0468;
    12: op1_06_in17 = reg_0737;
    13: op1_06_in17 = reg_0447;
    14: op1_06_in17 = reg_0198;
    15: op1_06_in17 = reg_0542;
    16: op1_06_in17 = reg_0498;
    17: op1_06_in17 = reg_0590;
    18: op1_06_in17 = reg_0408;
    19: op1_06_in17 = imem03_in[11:8];
    20: op1_06_in17 = reg_0348;
    21: op1_06_in17 = reg_0541;
    22: op1_06_in17 = reg_0636;
    23: op1_06_in17 = reg_0497;
    24: op1_06_in17 = imem04_in[107:104];
    25: op1_06_in17 = reg_0381;
    26: op1_06_in17 = imem04_in[119:116];
    27: op1_06_in17 = reg_0090;
    28: op1_06_in17 = reg_0363;
    29: op1_06_in17 = reg_0599;
    30: op1_06_in17 = reg_0129;
    31: op1_06_in17 = reg_0194;
    32: op1_06_in17 = imem02_in[63:60];
    33: op1_06_in17 = imem04_in[43:40];
    34: op1_06_in17 = reg_0466;
    36: op1_06_in17 = reg_0452;
    37: op1_06_in17 = reg_0193;
    38: op1_06_in17 = reg_0347;
    39: op1_06_in17 = reg_0295;
    40: op1_06_in17 = reg_0588;
    41: op1_06_in17 = reg_0723;
    42: op1_06_in17 = reg_0195;
    43: op1_06_in17 = reg_0097;
    44: op1_06_in17 = imem06_in[115:112];
    45: op1_06_in17 = reg_0158;
    46: op1_06_in17 = reg_0092;
    47: op1_06_in17 = imem05_in[111:108];
    49: op1_06_in17 = reg_0404;
    50: op1_06_in17 = reg_0488;
    51: op1_06_in17 = reg_0094;
    52: op1_06_in17 = reg_0512;
    78: op1_06_in17 = reg_0512;
    53: op1_06_in17 = reg_0245;
    54: op1_06_in17 = reg_0752;
    55: op1_06_in17 = reg_0721;
    57: op1_06_in17 = reg_0192;
    80: op1_06_in17 = reg_0192;
    59: op1_06_in17 = imem02_in[7:4];
    60: op1_06_in17 = imem01_in[39:36];
    61: op1_06_in17 = reg_0343;
    62: op1_06_in17 = reg_0031;
    63: op1_06_in17 = reg_0773;
    66: op1_06_in17 = reg_0268;
    67: op1_06_in17 = reg_0306;
    68: op1_06_in17 = reg_0503;
    69: op1_06_in17 = imem07_in[95:92];
    70: op1_06_in17 = reg_0478;
    71: op1_06_in17 = imem07_in[55:52];
    72: op1_06_in17 = reg_0179;
    74: op1_06_in17 = reg_0653;
    75: op1_06_in17 = imem03_in[95:92];
    76: op1_06_in17 = reg_0535;
    77: op1_06_in17 = reg_0808;
    82: op1_06_in17 = imem05_in[107:104];
    83: op1_06_in17 = imem02_in[127:124];
    84: op1_06_in17 = reg_0089;
    85: op1_06_in17 = reg_0458;
    86: op1_06_in17 = reg_0610;
    87: op1_06_in17 = reg_0218;
    88: op1_06_in17 = reg_0623;
    89: op1_06_in17 = reg_0443;
    92: op1_06_in17 = reg_0757;
    93: op1_06_in17 = reg_0392;
    94: op1_06_in17 = imem02_in[119:116];
    95: op1_06_in17 = reg_0136;
    96: op1_06_in17 = imem01_in[107:104];
    default: op1_06_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv17 = 1;
    11: op1_06_inv17 = 1;
    14: op1_06_inv17 = 1;
    17: op1_06_inv17 = 1;
    18: op1_06_inv17 = 1;
    19: op1_06_inv17 = 1;
    23: op1_06_inv17 = 1;
    24: op1_06_inv17 = 1;
    25: op1_06_inv17 = 1;
    28: op1_06_inv17 = 1;
    30: op1_06_inv17 = 1;
    33: op1_06_inv17 = 1;
    37: op1_06_inv17 = 1;
    38: op1_06_inv17 = 1;
    39: op1_06_inv17 = 1;
    41: op1_06_inv17 = 1;
    42: op1_06_inv17 = 1;
    45: op1_06_inv17 = 1;
    47: op1_06_inv17 = 1;
    51: op1_06_inv17 = 1;
    52: op1_06_inv17 = 1;
    66: op1_06_inv17 = 1;
    67: op1_06_inv17 = 1;
    68: op1_06_inv17 = 1;
    71: op1_06_inv17 = 1;
    72: op1_06_inv17 = 1;
    74: op1_06_inv17 = 1;
    77: op1_06_inv17 = 1;
    78: op1_06_inv17 = 1;
    85: op1_06_inv17 = 1;
    87: op1_06_inv17 = 1;
    88: op1_06_inv17 = 1;
    89: op1_06_inv17 = 1;
    92: op1_06_inv17 = 1;
    96: op1_06_inv17 = 1;
    default: op1_06_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in18 = reg_0346;
    5: op1_06_in18 = imem01_in[103:100];
    6: op1_06_in18 = reg_0043;
    7: op1_06_in18 = reg_0167;
    8: op1_06_in18 = reg_0326;
    9: op1_06_in18 = reg_0734;
    10: op1_06_in18 = reg_0662;
    11: op1_06_in18 = reg_0478;
    12: op1_06_in18 = reg_0733;
    16: op1_06_in18 = reg_0733;
    13: op1_06_in18 = reg_0445;
    14: op1_06_in18 = reg_0212;
    15: op1_06_in18 = reg_0558;
    17: op1_06_in18 = reg_0395;
    18: op1_06_in18 = reg_0351;
    19: op1_06_in18 = imem03_in[31:28];
    20: op1_06_in18 = reg_0356;
    21: op1_06_in18 = reg_0769;
    43: op1_06_in18 = reg_0769;
    22: op1_06_in18 = reg_0663;
    23: op1_06_in18 = reg_0512;
    24: op1_06_in18 = imem04_in[127:124];
    26: op1_06_in18 = imem04_in[127:124];
    25: op1_06_in18 = reg_0392;
    27: op1_06_in18 = reg_0741;
    28: op1_06_in18 = reg_0355;
    29: op1_06_in18 = reg_0583;
    30: op1_06_in18 = reg_0141;
    31: op1_06_in18 = reg_0198;
    32: op1_06_in18 = imem02_in[95:92];
    33: op1_06_in18 = imem04_in[115:112];
    34: op1_06_in18 = reg_0472;
    36: op1_06_in18 = reg_0456;
    37: op1_06_in18 = reg_0194;
    70: op1_06_in18 = reg_0194;
    38: op1_06_in18 = reg_0743;
    39: op1_06_in18 = reg_0257;
    40: op1_06_in18 = reg_0573;
    78: op1_06_in18 = reg_0573;
    41: op1_06_in18 = reg_0725;
    42: op1_06_in18 = imem01_in[11:8];
    44: op1_06_in18 = reg_0020;
    46: op1_06_in18 = reg_0533;
    47: op1_06_in18 = imem05_in[123:120];
    49: op1_06_in18 = reg_0406;
    50: op1_06_in18 = reg_0793;
    51: op1_06_in18 = reg_0532;
    52: op1_06_in18 = reg_0065;
    53: op1_06_in18 = reg_0276;
    54: op1_06_in18 = imem07_in[3:0];
    55: op1_06_in18 = reg_0723;
    57: op1_06_in18 = imem01_in[19:16];
    59: op1_06_in18 = imem02_in[15:12];
    60: op1_06_in18 = imem01_in[43:40];
    61: op1_06_in18 = reg_0092;
    62: op1_06_in18 = reg_0369;
    63: op1_06_in18 = reg_0764;
    66: op1_06_in18 = reg_0174;
    67: op1_06_in18 = reg_0574;
    68: op1_06_in18 = reg_0617;
    69: op1_06_in18 = imem07_in[107:104];
    71: op1_06_in18 = imem07_in[71:68];
    72: op1_06_in18 = reg_0161;
    74: op1_06_in18 = reg_0772;
    75: op1_06_in18 = reg_0528;
    76: op1_06_in18 = imem03_in[39:36];
    77: op1_06_in18 = reg_0003;
    80: op1_06_in18 = imem01_in[3:0];
    82: op1_06_in18 = imem05_in[119:116];
    83: op1_06_in18 = reg_0344;
    84: op1_06_in18 = reg_0730;
    85: op1_06_in18 = reg_0214;
    86: op1_06_in18 = reg_0679;
    87: op1_06_in18 = reg_0657;
    88: op1_06_in18 = reg_0019;
    89: op1_06_in18 = reg_0438;
    92: op1_06_in18 = reg_0740;
    93: op1_06_in18 = reg_0639;
    94: op1_06_in18 = imem02_in[127:124];
    95: op1_06_in18 = reg_0703;
    96: op1_06_in18 = imem01_in[111:108];
    default: op1_06_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv18 = 1;
    5: op1_06_inv18 = 1;
    8: op1_06_inv18 = 1;
    10: op1_06_inv18 = 1;
    11: op1_06_inv18 = 1;
    13: op1_06_inv18 = 1;
    14: op1_06_inv18 = 1;
    15: op1_06_inv18 = 1;
    18: op1_06_inv18 = 1;
    19: op1_06_inv18 = 1;
    20: op1_06_inv18 = 1;
    23: op1_06_inv18 = 1;
    24: op1_06_inv18 = 1;
    25: op1_06_inv18 = 1;
    28: op1_06_inv18 = 1;
    29: op1_06_inv18 = 1;
    30: op1_06_inv18 = 1;
    32: op1_06_inv18 = 1;
    33: op1_06_inv18 = 1;
    34: op1_06_inv18 = 1;
    38: op1_06_inv18 = 1;
    40: op1_06_inv18 = 1;
    41: op1_06_inv18 = 1;
    42: op1_06_inv18 = 1;
    43: op1_06_inv18 = 1;
    50: op1_06_inv18 = 1;
    51: op1_06_inv18 = 1;
    55: op1_06_inv18 = 1;
    57: op1_06_inv18 = 1;
    59: op1_06_inv18 = 1;
    60: op1_06_inv18 = 1;
    61: op1_06_inv18 = 1;
    62: op1_06_inv18 = 1;
    66: op1_06_inv18 = 1;
    68: op1_06_inv18 = 1;
    71: op1_06_inv18 = 1;
    72: op1_06_inv18 = 1;
    74: op1_06_inv18 = 1;
    76: op1_06_inv18 = 1;
    80: op1_06_inv18 = 1;
    85: op1_06_inv18 = 1;
    87: op1_06_inv18 = 1;
    88: op1_06_inv18 = 1;
    89: op1_06_inv18 = 1;
    95: op1_06_inv18 = 1;
    default: op1_06_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in19 = reg_0347;
    5: op1_06_in19 = reg_0500;
    33: op1_06_in19 = reg_0500;
    6: op1_06_in19 = reg_0053;
    7: op1_06_in19 = reg_0169;
    8: op1_06_in19 = reg_0329;
    9: op1_06_in19 = reg_0735;
    27: op1_06_in19 = reg_0735;
    10: op1_06_in19 = reg_0358;
    11: op1_06_in19 = reg_0204;
    12: op1_06_in19 = reg_0260;
    16: op1_06_in19 = reg_0260;
    13: op1_06_in19 = reg_0428;
    14: op1_06_in19 = reg_0190;
    15: op1_06_in19 = reg_0533;
    17: op1_06_in19 = reg_0384;
    18: op1_06_in19 = reg_0405;
    19: op1_06_in19 = imem03_in[55:52];
    20: op1_06_in19 = reg_0382;
    21: op1_06_in19 = imem03_in[59:56];
    22: op1_06_in19 = reg_0352;
    23: op1_06_in19 = reg_0506;
    24: op1_06_in19 = reg_0560;
    25: op1_06_in19 = reg_0383;
    26: op1_06_in19 = reg_0262;
    28: op1_06_in19 = reg_0073;
    29: op1_06_in19 = reg_0592;
    30: op1_06_in19 = imem06_in[47:44];
    31: op1_06_in19 = imem01_in[31:28];
    42: op1_06_in19 = imem01_in[31:28];
    57: op1_06_in19 = imem01_in[31:28];
    32: op1_06_in19 = imem02_in[107:104];
    34: op1_06_in19 = reg_0470;
    36: op1_06_in19 = reg_0187;
    37: op1_06_in19 = reg_0201;
    38: op1_06_in19 = reg_0096;
    39: op1_06_in19 = reg_0281;
    40: op1_06_in19 = reg_0568;
    41: op1_06_in19 = reg_0703;
    43: op1_06_in19 = reg_0540;
    44: op1_06_in19 = reg_0298;
    46: op1_06_in19 = reg_0769;
    47: op1_06_in19 = reg_0792;
    49: op1_06_in19 = reg_0242;
    50: op1_06_in19 = reg_0495;
    51: op1_06_in19 = imem03_in[7:4];
    52: op1_06_in19 = reg_0598;
    53: op1_06_in19 = reg_0249;
    54: op1_06_in19 = imem07_in[19:16];
    55: op1_06_in19 = reg_0717;
    59: op1_06_in19 = imem02_in[27:24];
    60: op1_06_in19 = imem01_in[91:88];
    61: op1_06_in19 = reg_0081;
    62: op1_06_in19 = reg_0763;
    63: op1_06_in19 = reg_0512;
    66: op1_06_in19 = reg_0172;
    67: op1_06_in19 = reg_0674;
    68: op1_06_in19 = reg_0679;
    69: op1_06_in19 = imem07_in[111:108];
    70: op1_06_in19 = imem01_in[11:8];
    71: op1_06_in19 = imem07_in[123:120];
    72: op1_06_in19 = reg_0167;
    74: op1_06_in19 = reg_0737;
    75: op1_06_in19 = reg_0488;
    76: op1_06_in19 = imem03_in[71:68];
    77: op1_06_in19 = reg_0803;
    78: op1_06_in19 = reg_0777;
    80: op1_06_in19 = imem01_in[7:4];
    82: op1_06_in19 = reg_0791;
    83: op1_06_in19 = reg_0341;
    84: op1_06_in19 = reg_0185;
    85: op1_06_in19 = reg_0191;
    86: op1_06_in19 = reg_0069;
    87: op1_06_in19 = reg_0664;
    88: op1_06_in19 = reg_0808;
    89: op1_06_in19 = reg_0730;
    92: op1_06_in19 = imem03_in[31:28];
    93: op1_06_in19 = reg_0304;
    94: op1_06_in19 = reg_0086;
    95: op1_06_in19 = reg_0532;
    96: op1_06_in19 = reg_0513;
    default: op1_06_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv19 = 1;
    7: op1_06_inv19 = 1;
    8: op1_06_inv19 = 1;
    9: op1_06_inv19 = 1;
    11: op1_06_inv19 = 1;
    12: op1_06_inv19 = 1;
    14: op1_06_inv19 = 1;
    18: op1_06_inv19 = 1;
    19: op1_06_inv19 = 1;
    20: op1_06_inv19 = 1;
    23: op1_06_inv19 = 1;
    24: op1_06_inv19 = 1;
    25: op1_06_inv19 = 1;
    28: op1_06_inv19 = 1;
    36: op1_06_inv19 = 1;
    38: op1_06_inv19 = 1;
    39: op1_06_inv19 = 1;
    40: op1_06_inv19 = 1;
    43: op1_06_inv19 = 1;
    52: op1_06_inv19 = 1;
    53: op1_06_inv19 = 1;
    55: op1_06_inv19 = 1;
    59: op1_06_inv19 = 1;
    60: op1_06_inv19 = 1;
    61: op1_06_inv19 = 1;
    66: op1_06_inv19 = 1;
    70: op1_06_inv19 = 1;
    76: op1_06_inv19 = 1;
    78: op1_06_inv19 = 1;
    82: op1_06_inv19 = 1;
    83: op1_06_inv19 = 1;
    84: op1_06_inv19 = 1;
    85: op1_06_inv19 = 1;
    87: op1_06_inv19 = 1;
    93: op1_06_inv19 = 1;
    95: op1_06_inv19 = 1;
    96: op1_06_inv19 = 1;
    default: op1_06_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in20 = reg_0092;
    5: op1_06_in20 = reg_0519;
    6: op1_06_in20 = reg_0071;
    7: op1_06_in20 = reg_0160;
    8: op1_06_in20 = reg_0339;
    9: op1_06_in20 = reg_0225;
    10: op1_06_in20 = reg_0353;
    11: op1_06_in20 = reg_0198;
    12: op1_06_in20 = reg_0261;
    13: op1_06_in20 = reg_0444;
    14: op1_06_in20 = reg_0197;
    15: op1_06_in20 = reg_0531;
    16: op1_06_in20 = reg_0269;
    17: op1_06_in20 = reg_0360;
    18: op1_06_in20 = reg_0371;
    19: op1_06_in20 = imem03_in[103:100];
    20: op1_06_in20 = reg_0315;
    21: op1_06_in20 = imem03_in[91:88];
    22: op1_06_in20 = reg_0364;
    23: op1_06_in20 = reg_0122;
    24: op1_06_in20 = reg_0552;
    25: op1_06_in20 = reg_0404;
    26: op1_06_in20 = reg_0544;
    27: op1_06_in20 = reg_0275;
    28: op1_06_in20 = reg_0096;
    29: op1_06_in20 = reg_0591;
    30: op1_06_in20 = imem06_in[63:60];
    31: op1_06_in20 = imem01_in[35:32];
    57: op1_06_in20 = imem01_in[35:32];
    32: op1_06_in20 = reg_0661;
    87: op1_06_in20 = reg_0661;
    33: op1_06_in20 = reg_0054;
    34: op1_06_in20 = reg_0474;
    36: op1_06_in20 = reg_0203;
    37: op1_06_in20 = reg_0190;
    38: op1_06_in20 = reg_0097;
    39: op1_06_in20 = reg_0066;
    40: op1_06_in20 = reg_0571;
    75: op1_06_in20 = reg_0571;
    41: op1_06_in20 = reg_0729;
    42: op1_06_in20 = imem01_in[43:40];
    43: op1_06_in20 = imem03_in[11:8];
    44: op1_06_in20 = reg_0619;
    46: op1_06_in20 = reg_0535;
    47: op1_06_in20 = reg_0798;
    49: op1_06_in20 = reg_0372;
    50: op1_06_in20 = reg_0782;
    51: op1_06_in20 = imem03_in[75:72];
    52: op1_06_in20 = reg_0399;
    53: op1_06_in20 = reg_0307;
    54: op1_06_in20 = imem07_in[27:24];
    55: op1_06_in20 = reg_0725;
    59: op1_06_in20 = imem02_in[35:32];
    60: op1_06_in20 = imem01_in[123:120];
    61: op1_06_in20 = reg_0530;
    62: op1_06_in20 = reg_0035;
    63: op1_06_in20 = reg_0607;
    66: op1_06_in20 = reg_0179;
    67: op1_06_in20 = reg_0121;
    68: op1_06_in20 = reg_0068;
    69: op1_06_in20 = reg_0718;
    70: op1_06_in20 = imem01_in[67:64];
    71: op1_06_in20 = reg_0721;
    74: op1_06_in20 = reg_0507;
    76: op1_06_in20 = imem03_in[87:84];
    77: op1_06_in20 = imem04_in[75:72];
    78: op1_06_in20 = reg_0794;
    80: op1_06_in20 = imem01_in[31:28];
    82: op1_06_in20 = reg_0146;
    83: op1_06_in20 = reg_0361;
    85: op1_06_in20 = reg_0210;
    86: op1_06_in20 = reg_0774;
    88: op1_06_in20 = reg_0007;
    89: op1_06_in20 = reg_0099;
    92: op1_06_in20 = imem03_in[67:64];
    93: op1_06_in20 = reg_0274;
    94: op1_06_in20 = reg_0705;
    95: op1_06_in20 = imem03_in[31:28];
    96: op1_06_in20 = reg_0499;
    default: op1_06_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv20 = 1;
    7: op1_06_inv20 = 1;
    8: op1_06_inv20 = 1;
    9: op1_06_inv20 = 1;
    11: op1_06_inv20 = 1;
    12: op1_06_inv20 = 1;
    15: op1_06_inv20 = 1;
    17: op1_06_inv20 = 1;
    18: op1_06_inv20 = 1;
    20: op1_06_inv20 = 1;
    22: op1_06_inv20 = 1;
    24: op1_06_inv20 = 1;
    26: op1_06_inv20 = 1;
    29: op1_06_inv20 = 1;
    31: op1_06_inv20 = 1;
    32: op1_06_inv20 = 1;
    36: op1_06_inv20 = 1;
    37: op1_06_inv20 = 1;
    38: op1_06_inv20 = 1;
    40: op1_06_inv20 = 1;
    47: op1_06_inv20 = 1;
    51: op1_06_inv20 = 1;
    59: op1_06_inv20 = 1;
    71: op1_06_inv20 = 1;
    75: op1_06_inv20 = 1;
    76: op1_06_inv20 = 1;
    77: op1_06_inv20 = 1;
    80: op1_06_inv20 = 1;
    85: op1_06_inv20 = 1;
    86: op1_06_inv20 = 1;
    88: op1_06_inv20 = 1;
    89: op1_06_inv20 = 1;
    94: op1_06_inv20 = 1;
    96: op1_06_inv20 = 1;
    default: op1_06_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in21 = reg_0051;
    5: op1_06_in21 = reg_0499;
    6: op1_06_in21 = reg_0064;
    7: op1_06_in21 = reg_0166;
    8: op1_06_in21 = reg_0355;
    9: op1_06_in21 = reg_0522;
    10: op1_06_in21 = reg_0342;
    11: op1_06_in21 = reg_0205;
    12: op1_06_in21 = reg_0228;
    13: op1_06_in21 = reg_0442;
    14: op1_06_in21 = imem01_in[27:24];
    15: op1_06_in21 = reg_0305;
    16: op1_06_in21 = reg_0744;
    17: op1_06_in21 = reg_0370;
    18: op1_06_in21 = reg_0313;
    19: op1_06_in21 = imem03_in[127:124];
    20: op1_06_in21 = reg_0813;
    63: op1_06_in21 = reg_0813;
    21: op1_06_in21 = reg_0582;
    22: op1_06_in21 = reg_0339;
    23: op1_06_in21 = reg_0125;
    24: op1_06_in21 = reg_0542;
    25: op1_06_in21 = reg_0368;
    26: op1_06_in21 = reg_0315;
    27: op1_06_in21 = reg_0260;
    28: op1_06_in21 = reg_0094;
    29: op1_06_in21 = reg_0589;
    30: op1_06_in21 = imem06_in[115:112];
    31: op1_06_in21 = imem01_in[43:40];
    32: op1_06_in21 = reg_0639;
    33: op1_06_in21 = reg_0301;
    34: op1_06_in21 = reg_0459;
    36: op1_06_in21 = reg_0207;
    37: op1_06_in21 = imem01_in[11:8];
    38: op1_06_in21 = imem03_in[35:32];
    39: op1_06_in21 = reg_0067;
    40: op1_06_in21 = reg_0569;
    41: op1_06_in21 = reg_0718;
    42: op1_06_in21 = imem01_in[47:44];
    43: op1_06_in21 = imem03_in[27:24];
    44: op1_06_in21 = reg_0766;
    46: op1_06_in21 = reg_0531;
    47: op1_06_in21 = reg_0495;
    49: op1_06_in21 = reg_0620;
    50: op1_06_in21 = reg_0786;
    51: op1_06_in21 = imem03_in[87:84];
    92: op1_06_in21 = imem03_in[87:84];
    52: op1_06_in21 = reg_0068;
    53: op1_06_in21 = reg_0066;
    54: op1_06_in21 = imem07_in[43:40];
    55: op1_06_in21 = reg_0709;
    57: op1_06_in21 = imem01_in[39:36];
    59: op1_06_in21 = imem02_in[75:72];
    60: op1_06_in21 = reg_0772;
    61: op1_06_in21 = imem03_in[43:40];
    62: op1_06_in21 = reg_0667;
    66: op1_06_in21 = reg_0160;
    67: op1_06_in21 = reg_0678;
    68: op1_06_in21 = reg_0771;
    69: op1_06_in21 = reg_0253;
    70: op1_06_in21 = imem01_in[75:72];
    71: op1_06_in21 = reg_0717;
    74: op1_06_in21 = reg_0294;
    75: op1_06_in21 = reg_0398;
    76: op1_06_in21 = imem03_in[107:104];
    77: op1_06_in21 = imem04_in[83:80];
    78: op1_06_in21 = reg_0657;
    80: op1_06_in21 = imem01_in[55:52];
    82: op1_06_in21 = reg_0550;
    83: op1_06_in21 = reg_0356;
    85: op1_06_in21 = imem01_in[3:0];
    86: op1_06_in21 = reg_0010;
    87: op1_06_in21 = imem07_in[7:4];
    88: op1_06_in21 = reg_0809;
    89: op1_06_in21 = reg_0184;
    93: op1_06_in21 = reg_0344;
    94: op1_06_in21 = reg_0059;
    95: op1_06_in21 = imem03_in[63:60];
    96: op1_06_in21 = reg_0238;
    default: op1_06_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv21 = 1;
    7: op1_06_inv21 = 1;
    8: op1_06_inv21 = 1;
    9: op1_06_inv21 = 1;
    11: op1_06_inv21 = 1;
    12: op1_06_inv21 = 1;
    13: op1_06_inv21 = 1;
    14: op1_06_inv21 = 1;
    15: op1_06_inv21 = 1;
    16: op1_06_inv21 = 1;
    19: op1_06_inv21 = 1;
    21: op1_06_inv21 = 1;
    22: op1_06_inv21 = 1;
    24: op1_06_inv21 = 1;
    26: op1_06_inv21 = 1;
    27: op1_06_inv21 = 1;
    29: op1_06_inv21 = 1;
    33: op1_06_inv21 = 1;
    34: op1_06_inv21 = 1;
    36: op1_06_inv21 = 1;
    37: op1_06_inv21 = 1;
    39: op1_06_inv21 = 1;
    41: op1_06_inv21 = 1;
    42: op1_06_inv21 = 1;
    43: op1_06_inv21 = 1;
    46: op1_06_inv21 = 1;
    47: op1_06_inv21 = 1;
    49: op1_06_inv21 = 1;
    50: op1_06_inv21 = 1;
    53: op1_06_inv21 = 1;
    55: op1_06_inv21 = 1;
    61: op1_06_inv21 = 1;
    62: op1_06_inv21 = 1;
    67: op1_06_inv21 = 1;
    68: op1_06_inv21 = 1;
    71: op1_06_inv21 = 1;
    76: op1_06_inv21 = 1;
    82: op1_06_inv21 = 1;
    85: op1_06_inv21 = 1;
    95: op1_06_inv21 = 1;
    96: op1_06_inv21 = 1;
    default: op1_06_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in22 = reg_0084;
    5: op1_06_in22 = reg_0507;
    6: op1_06_in22 = reg_0050;
    7: op1_06_in22 = reg_0177;
    66: op1_06_in22 = reg_0177;
    8: op1_06_in22 = reg_0097;
    9: op1_06_in22 = reg_0520;
    10: op1_06_in22 = reg_0082;
    11: op1_06_in22 = reg_0202;
    12: op1_06_in22 = reg_0132;
    13: op1_06_in22 = reg_0175;
    14: op1_06_in22 = imem01_in[35:32];
    15: op1_06_in22 = reg_0290;
    16: op1_06_in22 = reg_0266;
    17: op1_06_in22 = reg_0312;
    18: op1_06_in22 = reg_0406;
    19: op1_06_in22 = reg_0586;
    20: op1_06_in22 = reg_0817;
    21: op1_06_in22 = reg_0599;
    22: op1_06_in22 = reg_0081;
    23: op1_06_in22 = reg_0108;
    24: op1_06_in22 = reg_0537;
    25: op1_06_in22 = reg_0033;
    26: op1_06_in22 = reg_0542;
    27: op1_06_in22 = reg_0307;
    28: op1_06_in22 = imem03_in[39:36];
    29: op1_06_in22 = reg_0593;
    30: op1_06_in22 = reg_0625;
    31: op1_06_in22 = imem01_in[111:108];
    32: op1_06_in22 = reg_0651;
    33: op1_06_in22 = reg_0268;
    34: op1_06_in22 = reg_0478;
    36: op1_06_in22 = reg_0211;
    37: op1_06_in22 = imem01_in[15:12];
    38: op1_06_in22 = imem03_in[63:60];
    61: op1_06_in22 = imem03_in[63:60];
    39: op1_06_in22 = reg_0075;
    40: op1_06_in22 = reg_0398;
    41: op1_06_in22 = reg_0449;
    42: op1_06_in22 = imem01_in[59:56];
    57: op1_06_in22 = imem01_in[59:56];
    43: op1_06_in22 = imem03_in[75:72];
    44: op1_06_in22 = reg_0612;
    46: op1_06_in22 = reg_0526;
    47: op1_06_in22 = reg_0790;
    49: op1_06_in22 = reg_0621;
    50: op1_06_in22 = reg_0787;
    51: op1_06_in22 = reg_0596;
    52: op1_06_in22 = reg_0549;
    53: op1_06_in22 = reg_0732;
    54: op1_06_in22 = imem07_in[51:48];
    55: op1_06_in22 = reg_0705;
    59: op1_06_in22 = imem02_in[83:80];
    60: op1_06_in22 = reg_0645;
    62: op1_06_in22 = reg_0534;
    63: op1_06_in22 = reg_0032;
    67: op1_06_in22 = imem02_in[3:0];
    68: op1_06_in22 = reg_0640;
    69: op1_06_in22 = reg_0446;
    70: op1_06_in22 = reg_0376;
    71: op1_06_in22 = reg_0729;
    74: op1_06_in22 = reg_0425;
    75: op1_06_in22 = reg_0623;
    76: op1_06_in22 = reg_0347;
    77: op1_06_in22 = imem04_in[87:84];
    78: op1_06_in22 = reg_0664;
    80: op1_06_in22 = imem01_in[63:60];
    82: op1_06_in22 = reg_0386;
    83: op1_06_in22 = reg_0353;
    85: op1_06_in22 = imem01_in[55:52];
    86: op1_06_in22 = reg_0278;
    87: op1_06_in22 = imem07_in[19:16];
    88: op1_06_in22 = imem04_in[3:0];
    92: op1_06_in22 = imem03_in[95:92];
    93: op1_06_in22 = reg_0341;
    94: op1_06_in22 = reg_0485;
    95: op1_06_in22 = reg_0602;
    96: op1_06_in22 = reg_0232;
    default: op1_06_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv22 = 1;
    9: op1_06_inv22 = 1;
    11: op1_06_inv22 = 1;
    13: op1_06_inv22 = 1;
    14: op1_06_inv22 = 1;
    19: op1_06_inv22 = 1;
    20: op1_06_inv22 = 1;
    24: op1_06_inv22 = 1;
    25: op1_06_inv22 = 1;
    30: op1_06_inv22 = 1;
    31: op1_06_inv22 = 1;
    32: op1_06_inv22 = 1;
    33: op1_06_inv22 = 1;
    38: op1_06_inv22 = 1;
    42: op1_06_inv22 = 1;
    46: op1_06_inv22 = 1;
    50: op1_06_inv22 = 1;
    51: op1_06_inv22 = 1;
    52: op1_06_inv22 = 1;
    57: op1_06_inv22 = 1;
    59: op1_06_inv22 = 1;
    60: op1_06_inv22 = 1;
    62: op1_06_inv22 = 1;
    63: op1_06_inv22 = 1;
    67: op1_06_inv22 = 1;
    71: op1_06_inv22 = 1;
    74: op1_06_inv22 = 1;
    75: op1_06_inv22 = 1;
    80: op1_06_inv22 = 1;
    82: op1_06_inv22 = 1;
    83: op1_06_inv22 = 1;
    86: op1_06_inv22 = 1;
    87: op1_06_inv22 = 1;
    88: op1_06_inv22 = 1;
    92: op1_06_inv22 = 1;
    95: op1_06_inv22 = 1;
    default: op1_06_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in23 = reg_0093;
    5: op1_06_in23 = reg_0235;
    6: op1_06_in23 = imem05_in[91:88];
    7: op1_06_in23 = reg_0185;
    8: op1_06_in23 = reg_0091;
    9: op1_06_in23 = reg_0514;
    10: op1_06_in23 = reg_0073;
    11: op1_06_in23 = reg_0195;
    12: op1_06_in23 = reg_0148;
    16: op1_06_in23 = reg_0148;
    13: op1_06_in23 = reg_0169;
    14: op1_06_in23 = imem01_in[39:36];
    15: op1_06_in23 = reg_0295;
    33: op1_06_in23 = reg_0295;
    17: op1_06_in23 = reg_0811;
    18: op1_06_in23 = reg_0028;
    19: op1_06_in23 = reg_0579;
    21: op1_06_in23 = reg_0579;
    20: op1_06_in23 = reg_0818;
    22: op1_06_in23 = imem03_in[7:4];
    23: op1_06_in23 = imem02_in[15:12];
    24: op1_06_in23 = reg_0083;
    25: op1_06_in23 = reg_0815;
    26: op1_06_in23 = reg_0556;
    27: op1_06_in23 = reg_0277;
    28: op1_06_in23 = imem03_in[63:60];
    29: op1_06_in23 = reg_0595;
    30: op1_06_in23 = reg_0604;
    31: op1_06_in23 = imem01_in[119:116];
    32: op1_06_in23 = reg_0647;
    34: op1_06_in23 = reg_0200;
    36: op1_06_in23 = reg_0194;
    37: op1_06_in23 = imem01_in[19:16];
    38: op1_06_in23 = reg_0565;
    39: op1_06_in23 = reg_0256;
    40: op1_06_in23 = reg_0397;
    41: op1_06_in23 = reg_0444;
    42: op1_06_in23 = imem01_in[103:100];
    43: op1_06_in23 = imem03_in[91:88];
    44: op1_06_in23 = reg_0318;
    46: op1_06_in23 = imem03_in[39:36];
    47: op1_06_in23 = reg_0309;
    49: op1_06_in23 = reg_0368;
    50: op1_06_in23 = reg_0489;
    51: op1_06_in23 = reg_0580;
    52: op1_06_in23 = reg_0350;
    53: op1_06_in23 = reg_0744;
    54: op1_06_in23 = imem07_in[55:52];
    55: op1_06_in23 = reg_0707;
    71: op1_06_in23 = reg_0707;
    57: op1_06_in23 = imem01_in[87:84];
    59: op1_06_in23 = reg_0642;
    60: op1_06_in23 = reg_0820;
    61: op1_06_in23 = imem03_in[95:92];
    62: op1_06_in23 = reg_0032;
    63: op1_06_in23 = reg_0777;
    66: op1_06_in23 = reg_0157;
    67: op1_06_in23 = imem02_in[19:16];
    68: op1_06_in23 = reg_0776;
    69: op1_06_in23 = reg_0442;
    70: op1_06_in23 = reg_0645;
    74: op1_06_in23 = reg_0419;
    75: op1_06_in23 = reg_0006;
    76: op1_06_in23 = reg_0493;
    77: op1_06_in23 = imem04_in[111:108];
    78: op1_06_in23 = reg_0730;
    80: op1_06_in23 = reg_0336;
    82: op1_06_in23 = reg_0491;
    83: op1_06_in23 = reg_0342;
    85: op1_06_in23 = imem01_in[83:80];
    86: op1_06_in23 = reg_0008;
    87: op1_06_in23 = imem07_in[31:28];
    88: op1_06_in23 = reg_0173;
    92: op1_06_in23 = imem03_in[107:104];
    93: op1_06_in23 = reg_0356;
    94: op1_06_in23 = reg_0358;
    95: op1_06_in23 = reg_0338;
    96: op1_06_in23 = reg_0111;
    default: op1_06_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv23 = 1;
    6: op1_06_inv23 = 1;
    7: op1_06_inv23 = 1;
    8: op1_06_inv23 = 1;
    9: op1_06_inv23 = 1;
    11: op1_06_inv23 = 1;
    13: op1_06_inv23 = 1;
    14: op1_06_inv23 = 1;
    15: op1_06_inv23 = 1;
    18: op1_06_inv23 = 1;
    19: op1_06_inv23 = 1;
    22: op1_06_inv23 = 1;
    23: op1_06_inv23 = 1;
    24: op1_06_inv23 = 1;
    27: op1_06_inv23 = 1;
    29: op1_06_inv23 = 1;
    31: op1_06_inv23 = 1;
    32: op1_06_inv23 = 1;
    34: op1_06_inv23 = 1;
    36: op1_06_inv23 = 1;
    37: op1_06_inv23 = 1;
    40: op1_06_inv23 = 1;
    41: op1_06_inv23 = 1;
    47: op1_06_inv23 = 1;
    50: op1_06_inv23 = 1;
    52: op1_06_inv23 = 1;
    53: op1_06_inv23 = 1;
    57: op1_06_inv23 = 1;
    59: op1_06_inv23 = 1;
    61: op1_06_inv23 = 1;
    63: op1_06_inv23 = 1;
    66: op1_06_inv23 = 1;
    67: op1_06_inv23 = 1;
    71: op1_06_inv23 = 1;
    74: op1_06_inv23 = 1;
    75: op1_06_inv23 = 1;
    77: op1_06_inv23 = 1;
    78: op1_06_inv23 = 1;
    83: op1_06_inv23 = 1;
    85: op1_06_inv23 = 1;
    86: op1_06_inv23 = 1;
    88: op1_06_inv23 = 1;
    92: op1_06_inv23 = 1;
    95: op1_06_inv23 = 1;
    96: op1_06_inv23 = 1;
    default: op1_06_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in24 = imem03_in[59:56];
    5: op1_06_in24 = reg_0222;
    6: op1_06_in24 = imem05_in[99:96];
    7: op1_06_in24 = reg_0168;
    8: op1_06_in24 = reg_0084;
    9: op1_06_in24 = reg_0521;
    10: op1_06_in24 = imem03_in[3:0];
    11: op1_06_in24 = reg_0199;
    12: op1_06_in24 = reg_0154;
    13: op1_06_in24 = reg_0163;
    14: op1_06_in24 = imem01_in[55:52];
    15: op1_06_in24 = reg_0059;
    16: op1_06_in24 = reg_0152;
    17: op1_06_in24 = reg_0008;
    18: op1_06_in24 = reg_0039;
    38: op1_06_in24 = reg_0039;
    19: op1_06_in24 = reg_0585;
    20: op1_06_in24 = reg_0038;
    21: op1_06_in24 = reg_0572;
    22: op1_06_in24 = imem03_in[43:40];
    23: op1_06_in24 = imem02_in[31:28];
    24: op1_06_in24 = reg_0555;
    25: op1_06_in24 = reg_0817;
    26: op1_06_in24 = reg_0547;
    27: op1_06_in24 = reg_0089;
    28: op1_06_in24 = imem03_in[87:84];
    29: op1_06_in24 = reg_0588;
    30: op1_06_in24 = reg_0605;
    31: op1_06_in24 = imem01_in[123:120];
    32: op1_06_in24 = reg_0638;
    33: op1_06_in24 = reg_0286;
    34: op1_06_in24 = reg_0193;
    36: op1_06_in24 = imem01_in[23:20];
    37: op1_06_in24 = imem01_in[43:40];
    39: op1_06_in24 = imem05_in[7:4];
    40: op1_06_in24 = reg_0803;
    41: op1_06_in24 = reg_0442;
    42: op1_06_in24 = imem01_in[127:124];
    43: op1_06_in24 = reg_0601;
    44: op1_06_in24 = reg_0369;
    46: op1_06_in24 = imem03_in[47:44];
    47: op1_06_in24 = reg_0260;
    49: op1_06_in24 = reg_0231;
    50: op1_06_in24 = reg_0304;
    51: op1_06_in24 = reg_0595;
    52: op1_06_in24 = reg_0519;
    53: op1_06_in24 = reg_0147;
    54: op1_06_in24 = imem07_in[83:80];
    55: op1_06_in24 = reg_0701;
    57: op1_06_in24 = imem01_in[95:92];
    59: op1_06_in24 = reg_0666;
    60: op1_06_in24 = reg_0761;
    61: op1_06_in24 = imem03_in[107:104];
    62: op1_06_in24 = reg_0620;
    63: op1_06_in24 = reg_0620;
    67: op1_06_in24 = imem02_in[79:76];
    68: op1_06_in24 = reg_0109;
    69: op1_06_in24 = reg_0172;
    70: op1_06_in24 = reg_0820;
    80: op1_06_in24 = reg_0820;
    71: op1_06_in24 = reg_0706;
    74: op1_06_in24 = reg_0424;
    75: op1_06_in24 = reg_0019;
    76: op1_06_in24 = reg_0319;
    77: op1_06_in24 = imem04_in[115:112];
    78: op1_06_in24 = reg_0718;
    82: op1_06_in24 = reg_0720;
    83: op1_06_in24 = reg_0590;
    85: op1_06_in24 = imem01_in[107:104];
    86: op1_06_in24 = reg_0146;
    87: op1_06_in24 = imem07_in[35:32];
    88: op1_06_in24 = reg_0553;
    92: op1_06_in24 = imem03_in[119:116];
    93: op1_06_in24 = reg_0353;
    94: op1_06_in24 = reg_0362;
    95: op1_06_in24 = reg_0494;
    96: op1_06_in24 = reg_0068;
    default: op1_06_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_06_inv24 = 1;
    6: op1_06_inv24 = 1;
    7: op1_06_inv24 = 1;
    8: op1_06_inv24 = 1;
    12: op1_06_inv24 = 1;
    17: op1_06_inv24 = 1;
    19: op1_06_inv24 = 1;
    20: op1_06_inv24 = 1;
    21: op1_06_inv24 = 1;
    22: op1_06_inv24 = 1;
    23: op1_06_inv24 = 1;
    25: op1_06_inv24 = 1;
    27: op1_06_inv24 = 1;
    28: op1_06_inv24 = 1;
    29: op1_06_inv24 = 1;
    30: op1_06_inv24 = 1;
    31: op1_06_inv24 = 1;
    32: op1_06_inv24 = 1;
    33: op1_06_inv24 = 1;
    39: op1_06_inv24 = 1;
    40: op1_06_inv24 = 1;
    41: op1_06_inv24 = 1;
    43: op1_06_inv24 = 1;
    46: op1_06_inv24 = 1;
    49: op1_06_inv24 = 1;
    51: op1_06_inv24 = 1;
    52: op1_06_inv24 = 1;
    53: op1_06_inv24 = 1;
    55: op1_06_inv24 = 1;
    57: op1_06_inv24 = 1;
    59: op1_06_inv24 = 1;
    60: op1_06_inv24 = 1;
    69: op1_06_inv24 = 1;
    74: op1_06_inv24 = 1;
    75: op1_06_inv24 = 1;
    76: op1_06_inv24 = 1;
    77: op1_06_inv24 = 1;
    78: op1_06_inv24 = 1;
    80: op1_06_inv24 = 1;
    82: op1_06_inv24 = 1;
    85: op1_06_inv24 = 1;
    86: op1_06_inv24 = 1;
    87: op1_06_inv24 = 1;
    88: op1_06_inv24 = 1;
    92: op1_06_inv24 = 1;
    93: op1_06_inv24 = 1;
    94: op1_06_inv24 = 1;
    95: op1_06_inv24 = 1;
    96: op1_06_inv24 = 1;
    default: op1_06_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in25 = imem03_in[95:92];
    22: op1_06_in25 = imem03_in[95:92];
    5: op1_06_in25 = reg_0240;
    6: op1_06_in25 = imem05_in[123:120];
    8: op1_06_in25 = reg_0055;
    9: op1_06_in25 = reg_0518;
    10: op1_06_in25 = imem03_in[115:112];
    11: op1_06_in25 = reg_0197;
    34: op1_06_in25 = reg_0197;
    12: op1_06_in25 = reg_0153;
    14: op1_06_in25 = imem01_in[59:56];
    15: op1_06_in25 = reg_0054;
    17: op1_06_in25 = reg_0054;
    16: op1_06_in25 = reg_0142;
    18: op1_06_in25 = reg_0813;
    19: op1_06_in25 = reg_0578;
    20: op1_06_in25 = imem07_in[11:8];
    49: op1_06_in25 = imem07_in[11:8];
    21: op1_06_in25 = reg_0593;
    23: op1_06_in25 = imem02_in[39:36];
    24: op1_06_in25 = reg_0523;
    25: op1_06_in25 = imem07_in[71:68];
    26: op1_06_in25 = reg_0534;
    27: op1_06_in25 = reg_0132;
    28: op1_06_in25 = imem03_in[123:120];
    29: op1_06_in25 = reg_0392;
    30: op1_06_in25 = reg_0616;
    31: op1_06_in25 = reg_0513;
    32: op1_06_in25 = reg_0636;
    33: op1_06_in25 = reg_0258;
    36: op1_06_in25 = imem01_in[115:112];
    85: op1_06_in25 = imem01_in[115:112];
    37: op1_06_in25 = imem01_in[63:60];
    38: op1_06_in25 = reg_0595;
    39: op1_06_in25 = imem05_in[35:32];
    40: op1_06_in25 = reg_0799;
    41: op1_06_in25 = reg_0443;
    42: op1_06_in25 = reg_0759;
    43: op1_06_in25 = reg_0599;
    44: op1_06_in25 = reg_0408;
    46: op1_06_in25 = imem03_in[59:56];
    47: op1_06_in25 = reg_0272;
    50: op1_06_in25 = reg_0102;
    70: op1_06_in25 = reg_0102;
    51: op1_06_in25 = reg_0755;
    52: op1_06_in25 = reg_0275;
    53: op1_06_in25 = reg_0129;
    54: op1_06_in25 = reg_0704;
    55: op1_06_in25 = reg_0700;
    57: op1_06_in25 = reg_0085;
    59: op1_06_in25 = reg_0647;
    60: op1_06_in25 = reg_0765;
    61: op1_06_in25 = imem03_in[111:108];
    62: op1_06_in25 = reg_0496;
    63: op1_06_in25 = reg_0819;
    67: op1_06_in25 = imem02_in[95:92];
    68: op1_06_in25 = imem05_in[23:20];
    69: op1_06_in25 = reg_0161;
    71: op1_06_in25 = reg_0051;
    74: op1_06_in25 = reg_0124;
    75: op1_06_in25 = reg_0007;
    76: op1_06_in25 = reg_0646;
    77: op1_06_in25 = reg_0057;
    78: op1_06_in25 = reg_0714;
    80: op1_06_in25 = reg_0224;
    82: op1_06_in25 = reg_0229;
    83: op1_06_in25 = reg_0098;
    86: op1_06_in25 = imem05_in[11:8];
    87: op1_06_in25 = reg_0162;
    88: op1_06_in25 = reg_0261;
    92: op1_06_in25 = reg_0602;
    93: op1_06_in25 = reg_0527;
    94: op1_06_in25 = reg_0092;
    95: op1_06_in25 = reg_0384;
    96: op1_06_in25 = reg_0520;
    default: op1_06_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv25 = 1;
    5: op1_06_inv25 = 1;
    6: op1_06_inv25 = 1;
    8: op1_06_inv25 = 1;
    14: op1_06_inv25 = 1;
    21: op1_06_inv25 = 1;
    22: op1_06_inv25 = 1;
    24: op1_06_inv25 = 1;
    28: op1_06_inv25 = 1;
    29: op1_06_inv25 = 1;
    30: op1_06_inv25 = 1;
    31: op1_06_inv25 = 1;
    32: op1_06_inv25 = 1;
    38: op1_06_inv25 = 1;
    39: op1_06_inv25 = 1;
    41: op1_06_inv25 = 1;
    42: op1_06_inv25 = 1;
    44: op1_06_inv25 = 1;
    47: op1_06_inv25 = 1;
    49: op1_06_inv25 = 1;
    51: op1_06_inv25 = 1;
    52: op1_06_inv25 = 1;
    53: op1_06_inv25 = 1;
    55: op1_06_inv25 = 1;
    61: op1_06_inv25 = 1;
    69: op1_06_inv25 = 1;
    70: op1_06_inv25 = 1;
    74: op1_06_inv25 = 1;
    75: op1_06_inv25 = 1;
    76: op1_06_inv25 = 1;
    78: op1_06_inv25 = 1;
    82: op1_06_inv25 = 1;
    88: op1_06_inv25 = 1;
    94: op1_06_inv25 = 1;
    default: op1_06_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in26 = reg_0563;
    5: op1_06_in26 = reg_0216;
    6: op1_06_in26 = reg_0788;
    8: op1_06_in26 = imem03_in[7:4];
    9: op1_06_in26 = reg_0515;
    42: op1_06_in26 = reg_0515;
    10: op1_06_in26 = reg_0582;
    11: op1_06_in26 = imem01_in[11:8];
    12: op1_06_in26 = reg_0131;
    70: op1_06_in26 = reg_0131;
    14: op1_06_in26 = reg_0822;
    15: op1_06_in26 = reg_0058;
    16: op1_06_in26 = reg_0138;
    17: op1_06_in26 = reg_0043;
    93: op1_06_in26 = reg_0043;
    18: op1_06_in26 = reg_0040;
    19: op1_06_in26 = reg_0360;
    20: op1_06_in26 = imem07_in[15:12];
    21: op1_06_in26 = reg_0394;
    22: op1_06_in26 = imem03_in[99:96];
    23: op1_06_in26 = imem02_in[43:40];
    24: op1_06_in26 = reg_0556;
    25: op1_06_in26 = imem07_in[99:96];
    26: op1_06_in26 = reg_0306;
    27: op1_06_in26 = reg_0149;
    28: op1_06_in26 = reg_0585;
    29: op1_06_in26 = imem04_in[35:32];
    30: op1_06_in26 = reg_0606;
    31: op1_06_in26 = reg_0520;
    32: op1_06_in26 = reg_0652;
    33: op1_06_in26 = reg_0068;
    34: op1_06_in26 = imem01_in[55:52];
    36: op1_06_in26 = reg_0336;
    37: op1_06_in26 = imem01_in[67:64];
    38: op1_06_in26 = reg_0751;
    39: op1_06_in26 = imem05_in[75:72];
    40: op1_06_in26 = reg_0809;
    41: op1_06_in26 = reg_0448;
    43: op1_06_in26 = reg_0589;
    44: op1_06_in26 = reg_0370;
    46: op1_06_in26 = imem03_in[67:64];
    47: op1_06_in26 = reg_0132;
    49: op1_06_in26 = imem07_in[23:20];
    50: op1_06_in26 = reg_0224;
    51: op1_06_in26 = reg_0373;
    52: op1_06_in26 = reg_0288;
    53: op1_06_in26 = reg_0144;
    54: op1_06_in26 = reg_0719;
    55: op1_06_in26 = reg_0334;
    57: op1_06_in26 = reg_0497;
    59: op1_06_in26 = reg_0355;
    60: op1_06_in26 = reg_0759;
    61: op1_06_in26 = imem03_in[119:116];
    62: op1_06_in26 = imem07_in[67:64];
    63: op1_06_in26 = reg_0642;
    67: op1_06_in26 = reg_0639;
    68: op1_06_in26 = imem05_in[51:48];
    69: op1_06_in26 = reg_0182;
    71: op1_06_in26 = reg_0439;
    74: op1_06_in26 = reg_0108;
    75: op1_06_in26 = reg_0800;
    76: op1_06_in26 = reg_0490;
    77: op1_06_in26 = reg_0516;
    78: op1_06_in26 = imem07_in[3:0];
    80: op1_06_in26 = reg_0760;
    82: op1_06_in26 = reg_0277;
    83: op1_06_in26 = reg_0757;
    85: op1_06_in26 = reg_0741;
    86: op1_06_in26 = imem05_in[15:12];
    87: op1_06_in26 = reg_0382;
    88: op1_06_in26 = reg_0429;
    92: op1_06_in26 = reg_0486;
    94: op1_06_in26 = reg_0055;
    95: op1_06_in26 = reg_0549;
    96: op1_06_in26 = reg_0101;
    default: op1_06_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv26 = 1;
    5: op1_06_inv26 = 1;
    8: op1_06_inv26 = 1;
    10: op1_06_inv26 = 1;
    11: op1_06_inv26 = 1;
    17: op1_06_inv26 = 1;
    18: op1_06_inv26 = 1;
    21: op1_06_inv26 = 1;
    23: op1_06_inv26 = 1;
    24: op1_06_inv26 = 1;
    26: op1_06_inv26 = 1;
    27: op1_06_inv26 = 1;
    33: op1_06_inv26 = 1;
    38: op1_06_inv26 = 1;
    43: op1_06_inv26 = 1;
    55: op1_06_inv26 = 1;
    62: op1_06_inv26 = 1;
    67: op1_06_inv26 = 1;
    68: op1_06_inv26 = 1;
    70: op1_06_inv26 = 1;
    74: op1_06_inv26 = 1;
    76: op1_06_inv26 = 1;
    82: op1_06_inv26 = 1;
    83: op1_06_inv26 = 1;
    85: op1_06_inv26 = 1;
    87: op1_06_inv26 = 1;
    88: op1_06_inv26 = 1;
    93: op1_06_inv26 = 1;
    95: op1_06_inv26 = 1;
    96: op1_06_inv26 = 1;
    default: op1_06_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in27 = reg_0322;
    5: op1_06_in27 = reg_0123;
    96: op1_06_in27 = reg_0123;
    6: op1_06_in27 = reg_0795;
    8: op1_06_in27 = imem03_in[11:8];
    9: op1_06_in27 = reg_0516;
    10: op1_06_in27 = reg_0573;
    11: op1_06_in27 = imem01_in[27:24];
    12: op1_06_in27 = imem06_in[47:44];
    14: op1_06_in27 = reg_0514;
    15: op1_06_in27 = reg_0076;
    16: op1_06_in27 = reg_0153;
    17: op1_06_in27 = reg_0055;
    18: op1_06_in27 = reg_0037;
    19: op1_06_in27 = reg_0311;
    20: op1_06_in27 = imem07_in[19:16];
    21: op1_06_in27 = reg_0395;
    22: op1_06_in27 = imem03_in[127:124];
    61: op1_06_in27 = imem03_in[127:124];
    23: op1_06_in27 = imem02_in[67:64];
    24: op1_06_in27 = reg_0308;
    25: op1_06_in27 = imem07_in[107:104];
    26: op1_06_in27 = reg_0297;
    27: op1_06_in27 = reg_0145;
    28: op1_06_in27 = reg_0578;
    29: op1_06_in27 = imem04_in[63:60];
    30: op1_06_in27 = reg_0627;
    31: op1_06_in27 = reg_0215;
    32: op1_06_in27 = reg_0663;
    33: op1_06_in27 = reg_0077;
    34: op1_06_in27 = imem01_in[59:56];
    36: op1_06_in27 = reg_0513;
    37: op1_06_in27 = imem01_in[87:84];
    38: op1_06_in27 = reg_0394;
    39: op1_06_in27 = imem05_in[83:80];
    40: op1_06_in27 = imem04_in[3:0];
    41: op1_06_in27 = reg_0160;
    42: op1_06_in27 = reg_0567;
    43: op1_06_in27 = reg_0590;
    44: op1_06_in27 = reg_0407;
    46: op1_06_in27 = imem03_in[83:80];
    47: op1_06_in27 = reg_0133;
    49: op1_06_in27 = imem07_in[35:32];
    50: op1_06_in27 = reg_0066;
    51: op1_06_in27 = reg_0012;
    52: op1_06_in27 = imem05_in[27:24];
    86: op1_06_in27 = imem05_in[27:24];
    53: op1_06_in27 = reg_0628;
    54: op1_06_in27 = reg_0721;
    55: op1_06_in27 = reg_0441;
    57: op1_06_in27 = reg_0653;
    59: op1_06_in27 = reg_0665;
    60: op1_06_in27 = reg_0235;
    62: op1_06_in27 = imem07_in[127:124];
    63: op1_06_in27 = reg_0029;
    67: op1_06_in27 = reg_0647;
    68: op1_06_in27 = imem05_in[71:68];
    70: op1_06_in27 = reg_0110;
    71: op1_06_in27 = reg_0444;
    74: op1_06_in27 = reg_0677;
    75: op1_06_in27 = reg_0802;
    76: op1_06_in27 = reg_0019;
    77: op1_06_in27 = reg_0500;
    78: op1_06_in27 = imem07_in[11:8];
    80: op1_06_in27 = reg_0423;
    82: op1_06_in27 = reg_0812;
    83: op1_06_in27 = reg_0093;
    93: op1_06_in27 = reg_0093;
    85: op1_06_in27 = reg_0224;
    87: op1_06_in27 = reg_0712;
    88: op1_06_in27 = reg_0079;
    92: op1_06_in27 = reg_0389;
    94: op1_06_in27 = imem03_in[3:0];
    95: op1_06_in27 = reg_0811;
    default: op1_06_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv27 = 1;
    5: op1_06_inv27 = 1;
    9: op1_06_inv27 = 1;
    10: op1_06_inv27 = 1;
    11: op1_06_inv27 = 1;
    12: op1_06_inv27 = 1;
    17: op1_06_inv27 = 1;
    18: op1_06_inv27 = 1;
    19: op1_06_inv27 = 1;
    22: op1_06_inv27 = 1;
    24: op1_06_inv27 = 1;
    25: op1_06_inv27 = 1;
    26: op1_06_inv27 = 1;
    28: op1_06_inv27 = 1;
    29: op1_06_inv27 = 1;
    30: op1_06_inv27 = 1;
    31: op1_06_inv27 = 1;
    33: op1_06_inv27 = 1;
    36: op1_06_inv27 = 1;
    46: op1_06_inv27 = 1;
    50: op1_06_inv27 = 1;
    52: op1_06_inv27 = 1;
    53: op1_06_inv27 = 1;
    54: op1_06_inv27 = 1;
    59: op1_06_inv27 = 1;
    62: op1_06_inv27 = 1;
    68: op1_06_inv27 = 1;
    70: op1_06_inv27 = 1;
    74: op1_06_inv27 = 1;
    75: op1_06_inv27 = 1;
    76: op1_06_inv27 = 1;
    82: op1_06_inv27 = 1;
    86: op1_06_inv27 = 1;
    88: op1_06_inv27 = 1;
    94: op1_06_inv27 = 1;
    95: op1_06_inv27 = 1;
    96: op1_06_inv27 = 1;
    default: op1_06_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in28 = reg_0323;
    5: op1_06_in28 = reg_0105;
    96: op1_06_in28 = reg_0105;
    6: op1_06_in28 = reg_0493;
    8: op1_06_in28 = imem03_in[43:40];
    9: op1_06_in28 = imem01_in[19:16];
    10: op1_06_in28 = reg_0578;
    11: op1_06_in28 = imem01_in[35:32];
    12: op1_06_in28 = imem06_in[71:68];
    14: op1_06_in28 = reg_0825;
    15: op1_06_in28 = imem05_in[3:0];
    33: op1_06_in28 = imem05_in[3:0];
    16: op1_06_in28 = imem06_in[43:40];
    17: op1_06_in28 = reg_0057;
    18: op1_06_in28 = reg_0751;
    19: op1_06_in28 = reg_0374;
    20: op1_06_in28 = imem07_in[51:48];
    21: op1_06_in28 = reg_0369;
    22: op1_06_in28 = reg_0592;
    23: op1_06_in28 = imem02_in[75:72];
    24: op1_06_in28 = reg_0301;
    25: op1_06_in28 = imem07_in[115:112];
    26: op1_06_in28 = reg_0286;
    27: op1_06_in28 = reg_0136;
    28: op1_06_in28 = reg_0568;
    29: op1_06_in28 = imem04_in[123:120];
    30: op1_06_in28 = reg_0615;
    31: op1_06_in28 = reg_0242;
    32: op1_06_in28 = reg_0229;
    34: op1_06_in28 = imem01_in[71:68];
    36: op1_06_in28 = reg_0337;
    37: op1_06_in28 = imem01_in[111:108];
    38: op1_06_in28 = reg_0387;
    43: op1_06_in28 = reg_0387;
    39: op1_06_in28 = imem05_in[87:84];
    40: op1_06_in28 = imem04_in[107:104];
    41: op1_06_in28 = reg_0183;
    42: op1_06_in28 = reg_0123;
    44: op1_06_in28 = reg_0406;
    46: op1_06_in28 = imem03_in[99:96];
    47: op1_06_in28 = reg_0144;
    49: op1_06_in28 = imem07_in[39:36];
    50: op1_06_in28 = reg_0101;
    51: op1_06_in28 = reg_0001;
    52: op1_06_in28 = imem05_in[31:28];
    53: op1_06_in28 = reg_0625;
    54: op1_06_in28 = reg_0726;
    55: op1_06_in28 = reg_0266;
    57: op1_06_in28 = reg_0772;
    59: op1_06_in28 = reg_0427;
    60: op1_06_in28 = reg_0421;
    61: op1_06_in28 = reg_0602;
    62: op1_06_in28 = reg_0728;
    63: op1_06_in28 = reg_0752;
    67: op1_06_in28 = reg_0655;
    68: op1_06_in28 = imem05_in[95:92];
    70: op1_06_in28 = reg_0760;
    71: op1_06_in28 = reg_0174;
    74: op1_06_in28 = reg_0601;
    75: op1_06_in28 = reg_0799;
    76: op1_06_in28 = reg_0803;
    77: op1_06_in28 = reg_0556;
    78: op1_06_in28 = imem07_in[47:44];
    80: op1_06_in28 = reg_0108;
    82: op1_06_in28 = reg_0148;
    83: op1_06_in28 = imem03_in[39:36];
    85: op1_06_in28 = reg_0388;
    86: op1_06_in28 = imem05_in[71:68];
    87: op1_06_in28 = reg_0157;
    88: op1_06_in28 = reg_0283;
    92: op1_06_in28 = reg_0395;
    93: op1_06_in28 = imem03_in[11:8];
    94: op1_06_in28 = imem03_in[55:52];
    95: op1_06_in28 = reg_0368;
    default: op1_06_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_06_inv28 = 1;
    10: op1_06_inv28 = 1;
    18: op1_06_inv28 = 1;
    21: op1_06_inv28 = 1;
    22: op1_06_inv28 = 1;
    23: op1_06_inv28 = 1;
    25: op1_06_inv28 = 1;
    26: op1_06_inv28 = 1;
    27: op1_06_inv28 = 1;
    29: op1_06_inv28 = 1;
    30: op1_06_inv28 = 1;
    32: op1_06_inv28 = 1;
    37: op1_06_inv28 = 1;
    39: op1_06_inv28 = 1;
    40: op1_06_inv28 = 1;
    41: op1_06_inv28 = 1;
    42: op1_06_inv28 = 1;
    46: op1_06_inv28 = 1;
    47: op1_06_inv28 = 1;
    49: op1_06_inv28 = 1;
    50: op1_06_inv28 = 1;
    51: op1_06_inv28 = 1;
    54: op1_06_inv28 = 1;
    55: op1_06_inv28 = 1;
    57: op1_06_inv28 = 1;
    60: op1_06_inv28 = 1;
    67: op1_06_inv28 = 1;
    68: op1_06_inv28 = 1;
    75: op1_06_inv28 = 1;
    82: op1_06_inv28 = 1;
    85: op1_06_inv28 = 1;
    87: op1_06_inv28 = 1;
    88: op1_06_inv28 = 1;
    93: op1_06_inv28 = 1;
    default: op1_06_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in29 = reg_0006;
    5: op1_06_in29 = reg_0124;
    42: op1_06_in29 = reg_0124;
    6: op1_06_in29 = reg_0794;
    8: op1_06_in29 = imem03_in[55:52];
    9: op1_06_in29 = imem01_in[75:72];
    10: op1_06_in29 = reg_0581;
    11: op1_06_in29 = imem01_in[127:124];
    12: op1_06_in29 = imem06_in[115:112];
    14: op1_06_in29 = reg_0507;
    15: op1_06_in29 = imem05_in[7:4];
    16: op1_06_in29 = imem06_in[67:64];
    17: op1_06_in29 = reg_0058;
    18: op1_06_in29 = imem07_in[3:0];
    19: op1_06_in29 = reg_0389;
    20: op1_06_in29 = imem07_in[63:60];
    78: op1_06_in29 = imem07_in[63:60];
    21: op1_06_in29 = reg_0000;
    22: op1_06_in29 = reg_0591;
    23: op1_06_in29 = imem02_in[79:76];
    24: op1_06_in29 = reg_0283;
    25: op1_06_in29 = reg_0716;
    62: op1_06_in29 = reg_0716;
    26: op1_06_in29 = reg_0079;
    27: op1_06_in29 = reg_0133;
    28: op1_06_in29 = reg_0373;
    29: op1_06_in29 = reg_0262;
    30: op1_06_in29 = reg_0025;
    31: op1_06_in29 = reg_0220;
    32: op1_06_in29 = reg_0353;
    33: op1_06_in29 = imem05_in[23:20];
    34: op1_06_in29 = imem01_in[87:84];
    36: op1_06_in29 = reg_0771;
    37: op1_06_in29 = imem01_in[115:112];
    38: op1_06_in29 = reg_0571;
    39: op1_06_in29 = reg_0788;
    40: op1_06_in29 = imem04_in[111:108];
    41: op1_06_in29 = reg_0164;
    43: op1_06_in29 = reg_0383;
    44: op1_06_in29 = reg_0812;
    46: op1_06_in29 = reg_0579;
    47: op1_06_in29 = imem06_in[43:40];
    49: op1_06_in29 = imem07_in[83:80];
    50: op1_06_in29 = reg_0086;
    51: op1_06_in29 = reg_0002;
    52: op1_06_in29 = imem05_in[39:36];
    53: op1_06_in29 = reg_0291;
    54: op1_06_in29 = reg_0717;
    55: op1_06_in29 = reg_0061;
    57: op1_06_in29 = reg_0663;
    59: op1_06_in29 = reg_0364;
    60: op1_06_in29 = reg_0511;
    61: op1_06_in29 = reg_0582;
    63: op1_06_in29 = imem07_in[7:4];
    67: op1_06_in29 = reg_0548;
    68: op1_06_in29 = imem05_in[99:96];
    70: op1_06_in29 = reg_0225;
    71: op1_06_in29 = reg_0181;
    74: op1_06_in29 = reg_0678;
    75: op1_06_in29 = imem04_in[7:4];
    76: op1_06_in29 = reg_0807;
    77: op1_06_in29 = reg_0611;
    80: op1_06_in29 = reg_0677;
    96: op1_06_in29 = reg_0677;
    82: op1_06_in29 = reg_0742;
    83: op1_06_in29 = imem03_in[43:40];
    85: op1_06_in29 = reg_0397;
    86: op1_06_in29 = imem05_in[87:84];
    87: op1_06_in29 = reg_0727;
    88: op1_06_in29 = reg_0617;
    92: op1_06_in29 = reg_0384;
    93: op1_06_in29 = imem03_in[123:120];
    94: op1_06_in29 = imem03_in[79:76];
    95: op1_06_in29 = reg_0800;
    default: op1_06_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv29 = 1;
    5: op1_06_inv29 = 1;
    6: op1_06_inv29 = 1;
    9: op1_06_inv29 = 1;
    10: op1_06_inv29 = 1;
    11: op1_06_inv29 = 1;
    12: op1_06_inv29 = 1;
    14: op1_06_inv29 = 1;
    16: op1_06_inv29 = 1;
    18: op1_06_inv29 = 1;
    20: op1_06_inv29 = 1;
    21: op1_06_inv29 = 1;
    22: op1_06_inv29 = 1;
    23: op1_06_inv29 = 1;
    28: op1_06_inv29 = 1;
    29: op1_06_inv29 = 1;
    30: op1_06_inv29 = 1;
    33: op1_06_inv29 = 1;
    37: op1_06_inv29 = 1;
    39: op1_06_inv29 = 1;
    41: op1_06_inv29 = 1;
    44: op1_06_inv29 = 1;
    46: op1_06_inv29 = 1;
    47: op1_06_inv29 = 1;
    51: op1_06_inv29 = 1;
    52: op1_06_inv29 = 1;
    53: op1_06_inv29 = 1;
    55: op1_06_inv29 = 1;
    57: op1_06_inv29 = 1;
    59: op1_06_inv29 = 1;
    60: op1_06_inv29 = 1;
    61: op1_06_inv29 = 1;
    63: op1_06_inv29 = 1;
    68: op1_06_inv29 = 1;
    70: op1_06_inv29 = 1;
    71: op1_06_inv29 = 1;
    75: op1_06_inv29 = 1;
    76: op1_06_inv29 = 1;
    77: op1_06_inv29 = 1;
    78: op1_06_inv29 = 1;
    80: op1_06_inv29 = 1;
    85: op1_06_inv29 = 1;
    86: op1_06_inv29 = 1;
    87: op1_06_inv29 = 1;
    88: op1_06_inv29 = 1;
    92: op1_06_inv29 = 1;
    94: op1_06_inv29 = 1;
    96: op1_06_inv29 = 1;
    default: op1_06_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_06_in30 = reg_0001;
    21: op1_06_in30 = reg_0001;
    5: op1_06_in30 = reg_0125;
    6: op1_06_in30 = reg_0790;
    8: op1_06_in30 = imem03_in[59:56];
    9: op1_06_in30 = imem01_in[79:76];
    10: op1_06_in30 = reg_0398;
    11: op1_06_in30 = reg_0500;
    12: op1_06_in30 = reg_0621;
    14: op1_06_in30 = reg_0821;
    15: op1_06_in30 = imem05_in[27:24];
    16: op1_06_in30 = imem06_in[95:92];
    47: op1_06_in30 = imem06_in[95:92];
    17: op1_06_in30 = reg_0552;
    18: op1_06_in30 = imem07_in[27:24];
    19: op1_06_in30 = reg_0808;
    20: op1_06_in30 = imem07_in[75:72];
    22: op1_06_in30 = reg_0593;
    23: op1_06_in30 = reg_0656;
    24: op1_06_in30 = reg_0534;
    25: op1_06_in30 = reg_0704;
    26: op1_06_in30 = reg_0074;
    27: op1_06_in30 = reg_0131;
    28: op1_06_in30 = reg_0571;
    29: op1_06_in30 = reg_0553;
    30: op1_06_in30 = reg_0369;
    31: op1_06_in30 = reg_0247;
    32: op1_06_in30 = reg_0351;
    33: op1_06_in30 = imem05_in[95:92];
    34: op1_06_in30 = reg_0758;
    36: op1_06_in30 = reg_0235;
    70: op1_06_in30 = reg_0235;
    37: op1_06_in30 = reg_0334;
    38: op1_06_in30 = reg_0397;
    39: op1_06_in30 = reg_0789;
    40: op1_06_in30 = imem04_in[115:112];
    42: op1_06_in30 = reg_0119;
    43: op1_06_in30 = reg_0385;
    44: op1_06_in30 = reg_0620;
    46: op1_06_in30 = reg_0587;
    49: op1_06_in30 = reg_0722;
    50: op1_06_in30 = reg_0137;
    51: op1_06_in30 = reg_0003;
    52: op1_06_in30 = imem05_in[75:72];
    53: op1_06_in30 = reg_0624;
    54: op1_06_in30 = reg_0702;
    55: op1_06_in30 = reg_0434;
    57: op1_06_in30 = reg_0649;
    59: op1_06_in30 = reg_0586;
    60: op1_06_in30 = reg_0422;
    61: op1_06_in30 = reg_0599;
    62: op1_06_in30 = reg_0710;
    63: op1_06_in30 = imem07_in[67:64];
    67: op1_06_in30 = reg_0114;
    68: op1_06_in30 = reg_0792;
    71: op1_06_in30 = reg_0160;
    74: op1_06_in30 = imem02_in[7:4];
    75: op1_06_in30 = imem04_in[11:8];
    76: op1_06_in30 = reg_0801;
    77: op1_06_in30 = reg_0430;
    78: op1_06_in30 = imem07_in[95:92];
    80: op1_06_in30 = imem02_in[23:20];
    82: op1_06_in30 = imem06_in[19:16];
    83: op1_06_in30 = imem03_in[99:96];
    85: op1_06_in30 = reg_0258;
    86: op1_06_in30 = imem05_in[115:112];
    87: op1_06_in30 = reg_0636;
    88: op1_06_in30 = reg_0513;
    92: op1_06_in30 = reg_0417;
    93: op1_06_in30 = reg_0383;
    94: op1_06_in30 = reg_0597;
    95: op1_06_in30 = reg_0306;
    96: op1_06_in30 = imem02_in[27:24];
    default: op1_06_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_06_inv30 = 1;
    5: op1_06_inv30 = 1;
    8: op1_06_inv30 = 1;
    10: op1_06_inv30 = 1;
    11: op1_06_inv30 = 1;
    12: op1_06_inv30 = 1;
    14: op1_06_inv30 = 1;
    16: op1_06_inv30 = 1;
    17: op1_06_inv30 = 1;
    19: op1_06_inv30 = 1;
    20: op1_06_inv30 = 1;
    23: op1_06_inv30 = 1;
    26: op1_06_inv30 = 1;
    29: op1_06_inv30 = 1;
    31: op1_06_inv30 = 1;
    32: op1_06_inv30 = 1;
    38: op1_06_inv30 = 1;
    39: op1_06_inv30 = 1;
    43: op1_06_inv30 = 1;
    44: op1_06_inv30 = 1;
    46: op1_06_inv30 = 1;
    49: op1_06_inv30 = 1;
    50: op1_06_inv30 = 1;
    51: op1_06_inv30 = 1;
    52: op1_06_inv30 = 1;
    54: op1_06_inv30 = 1;
    55: op1_06_inv30 = 1;
    57: op1_06_inv30 = 1;
    62: op1_06_inv30 = 1;
    67: op1_06_inv30 = 1;
    68: op1_06_inv30 = 1;
    75: op1_06_inv30 = 1;
    85: op1_06_inv30 = 1;
    88: op1_06_inv30 = 1;
    93: op1_06_inv30 = 1;
    94: op1_06_inv30 = 1;
    95: op1_06_inv30 = 1;
    default: op1_06_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_06_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_06_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in00 = reg_0007;
    5: op1_07_in00 = reg_0102;
    6: op1_07_in00 = reg_0784;
    7: op1_07_in00 = imem00_in[23:20];
    66: op1_07_in00 = imem00_in[23:20];
    84: op1_07_in00 = imem00_in[23:20];
    8: op1_07_in00 = imem03_in[83:80];
    9: op1_07_in00 = imem01_in[91:88];
    10: op1_07_in00 = reg_0397;
    43: op1_07_in00 = reg_0397;
    11: op1_07_in00 = reg_0824;
    12: op1_07_in00 = reg_0606;
    13: op1_07_in00 = imem00_in[11:8];
    45: op1_07_in00 = imem00_in[11:8];
    56: op1_07_in00 = imem00_in[11:8];
    3: op1_07_in00 = imem07_in[91:88];
    14: op1_07_in00 = reg_0220;
    15: op1_07_in00 = imem05_in[31:28];
    16: op1_07_in00 = imem06_in[123:120];
    17: op1_07_in00 = reg_0534;
    18: op1_07_in00 = imem07_in[35:32];
    19: op1_07_in00 = imem04_in[3:0];
    20: op1_07_in00 = imem07_in[87:84];
    2: op1_07_in00 = imem07_in[55:52];
    1: op1_07_in00 = imem07_in[55:52];
    21: op1_07_in00 = reg_0003;
    22: op1_07_in00 = reg_0580;
    23: op1_07_in00 = reg_0651;
    24: op1_07_in00 = reg_0306;
    25: op1_07_in00 = imem00_in[43:40];
    35: op1_07_in00 = imem00_in[43:40];
    26: op1_07_in00 = imem05_in[11:8];
    27: op1_07_in00 = imem06_in[43:40];
    82: op1_07_in00 = imem06_in[43:40];
    28: op1_07_in00 = reg_0392;
    29: op1_07_in00 = reg_0500;
    30: op1_07_in00 = reg_0408;
    31: op1_07_in00 = reg_0237;
    32: op1_07_in00 = reg_0342;
    33: op1_07_in00 = imem05_in[115:112];
    34: op1_07_in00 = reg_0501;
    36: op1_07_in00 = reg_0246;
    37: op1_07_in00 = reg_0549;
    38: op1_07_in00 = reg_0393;
    39: op1_07_in00 = reg_0493;
    40: op1_07_in00 = imem04_in[123:120];
    41: op1_07_in00 = imem00_in[99:96];
    91: op1_07_in00 = imem00_in[99:96];
    42: op1_07_in00 = reg_0100;
    44: op1_07_in00 = reg_0029;
    46: op1_07_in00 = reg_0592;
    47: op1_07_in00 = imem06_in[99:96];
    48: op1_07_in00 = imem00_in[7:4];
    69: op1_07_in00 = imem00_in[7:4];
    49: op1_07_in00 = reg_0717;
    50: op1_07_in00 = imem06_in[3:0];
    51: op1_07_in00 = reg_0810;
    52: op1_07_in00 = reg_0795;
    53: op1_07_in00 = reg_0416;
    54: op1_07_in00 = reg_0703;
    55: op1_07_in00 = reg_0437;
    57: op1_07_in00 = reg_0322;
    58: op1_07_in00 = imem00_in[31:28];
    72: op1_07_in00 = imem00_in[31:28];
    73: op1_07_in00 = imem00_in[31:28];
    59: op1_07_in00 = reg_0341;
    60: op1_07_in00 = reg_0217;
    61: op1_07_in00 = reg_0751;
    62: op1_07_in00 = reg_0726;
    63: op1_07_in00 = imem07_in[83:80];
    64: op1_07_in00 = imem00_in[27:24];
    65: op1_07_in00 = imem00_in[39:36];
    67: op1_07_in00 = reg_0372;
    68: op1_07_in00 = reg_0781;
    70: op1_07_in00 = reg_0418;
    71: op1_07_in00 = reg_0163;
    74: op1_07_in00 = imem02_in[15:12];
    75: op1_07_in00 = imem04_in[51:48];
    76: op1_07_in00 = reg_0800;
    77: op1_07_in00 = reg_0078;
    78: op1_07_in00 = imem07_in[103:100];
    79: op1_07_in00 = imem00_in[59:56];
    80: op1_07_in00 = imem02_in[31:28];
    81: op1_07_in00 = imem00_in[3:0];
    83: op1_07_in00 = imem03_in[107:104];
    85: op1_07_in00 = reg_0422;
    86: op1_07_in00 = reg_0742;
    87: op1_07_in00 = reg_0449;
    88: op1_07_in00 = reg_0771;
    89: op1_07_in00 = imem00_in[15:12];
    90: op1_07_in00 = reg_0019;
    92: op1_07_in00 = reg_0483;
    93: op1_07_in00 = reg_0599;
    94: op1_07_in00 = reg_0801;
    95: op1_07_in00 = reg_0802;
    96: op1_07_in00 = imem02_in[123:120];
    default: op1_07_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_07_inv00 = 1;
    8: op1_07_inv00 = 1;
    10: op1_07_inv00 = 1;
    11: op1_07_inv00 = 1;
    3: op1_07_inv00 = 1;
    15: op1_07_inv00 = 1;
    16: op1_07_inv00 = 1;
    18: op1_07_inv00 = 1;
    19: op1_07_inv00 = 1;
    20: op1_07_inv00 = 1;
    21: op1_07_inv00 = 1;
    23: op1_07_inv00 = 1;
    25: op1_07_inv00 = 1;
    30: op1_07_inv00 = 1;
    31: op1_07_inv00 = 1;
    33: op1_07_inv00 = 1;
    34: op1_07_inv00 = 1;
    36: op1_07_inv00 = 1;
    37: op1_07_inv00 = 1;
    39: op1_07_inv00 = 1;
    44: op1_07_inv00 = 1;
    47: op1_07_inv00 = 1;
    48: op1_07_inv00 = 1;
    49: op1_07_inv00 = 1;
    50: op1_07_inv00 = 1;
    52: op1_07_inv00 = 1;
    57: op1_07_inv00 = 1;
    61: op1_07_inv00 = 1;
    65: op1_07_inv00 = 1;
    70: op1_07_inv00 = 1;
    73: op1_07_inv00 = 1;
    74: op1_07_inv00 = 1;
    76: op1_07_inv00 = 1;
    77: op1_07_inv00 = 1;
    78: op1_07_inv00 = 1;
    79: op1_07_inv00 = 1;
    82: op1_07_inv00 = 1;
    90: op1_07_inv00 = 1;
    91: op1_07_inv00 = 1;
    92: op1_07_inv00 = 1;
    93: op1_07_inv00 = 1;
    95: op1_07_inv00 = 1;
    96: op1_07_inv00 = 1;
    default: op1_07_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in01 = reg_0008;
    94: op1_07_in01 = reg_0008;
    5: op1_07_in01 = reg_0115;
    90: op1_07_in01 = reg_0115;
    6: op1_07_in01 = reg_0259;
    7: op1_07_in01 = imem00_in[27:24];
    66: op1_07_in01 = imem00_in[27:24];
    8: op1_07_in01 = imem03_in[87:84];
    9: op1_07_in01 = imem01_in[111:108];
    10: op1_07_in01 = reg_0361;
    11: op1_07_in01 = reg_0778;
    12: op1_07_in01 = reg_0609;
    13: op1_07_in01 = imem00_in[15:12];
    48: op1_07_in01 = imem00_in[15:12];
    3: op1_07_in01 = reg_0443;
    14: op1_07_in01 = reg_0236;
    15: op1_07_in01 = imem05_in[63:60];
    16: op1_07_in01 = reg_0610;
    17: op1_07_in01 = reg_0535;
    32: op1_07_in01 = reg_0535;
    18: op1_07_in01 = imem07_in[63:60];
    1: op1_07_in01 = imem07_in[63:60];
    19: op1_07_in01 = imem04_in[47:44];
    20: op1_07_in01 = imem07_in[99:96];
    2: op1_07_in01 = imem07_in[103:100];
    21: op1_07_in01 = reg_0799;
    22: op1_07_in01 = reg_0384;
    23: op1_07_in01 = reg_0652;
    24: op1_07_in01 = reg_0293;
    25: op1_07_in01 = imem00_in[95:92];
    56: op1_07_in01 = imem00_in[95:92];
    26: op1_07_in01 = imem05_in[23:20];
    27: op1_07_in01 = imem06_in[71:68];
    28: op1_07_in01 = reg_0006;
    38: op1_07_in01 = reg_0006;
    29: op1_07_in01 = reg_0301;
    30: op1_07_in01 = reg_0776;
    31: op1_07_in01 = reg_0041;
    33: op1_07_in01 = imem05_in[123:120];
    34: op1_07_in01 = reg_0497;
    35: op1_07_in01 = imem00_in[63:60];
    36: op1_07_in01 = reg_0244;
    37: op1_07_in01 = reg_0563;
    39: op1_07_in01 = reg_0793;
    40: op1_07_in01 = reg_0544;
    41: op1_07_in01 = imem00_in[119:116];
    42: op1_07_in01 = reg_0107;
    43: op1_07_in01 = reg_0811;
    44: op1_07_in01 = imem07_in[11:8];
    45: op1_07_in01 = imem00_in[31:28];
    84: op1_07_in01 = imem00_in[31:28];
    46: op1_07_in01 = reg_0751;
    47: op1_07_in01 = imem06_in[119:116];
    49: op1_07_in01 = reg_0718;
    50: op1_07_in01 = imem06_in[15:12];
    51: op1_07_in01 = reg_0809;
    52: op1_07_in01 = reg_0494;
    53: op1_07_in01 = reg_0286;
    54: op1_07_in01 = reg_0724;
    55: op1_07_in01 = reg_0180;
    57: op1_07_in01 = reg_0100;
    58: op1_07_in01 = imem00_in[87:84];
    59: op1_07_in01 = reg_0360;
    60: op1_07_in01 = reg_0240;
    61: op1_07_in01 = reg_0394;
    62: op1_07_in01 = reg_0725;
    63: op1_07_in01 = imem07_in[123:120];
    64: op1_07_in01 = imem00_in[51:48];
    65: op1_07_in01 = imem00_in[43:40];
    72: op1_07_in01 = imem00_in[43:40];
    67: op1_07_in01 = reg_0237;
    68: op1_07_in01 = reg_0282;
    69: op1_07_in01 = imem00_in[107:104];
    70: op1_07_in01 = reg_0425;
    71: op1_07_in01 = reg_0166;
    73: op1_07_in01 = imem00_in[39:36];
    74: op1_07_in01 = imem02_in[19:16];
    75: op1_07_in01 = imem04_in[67:64];
    76: op1_07_in01 = reg_0014;
    77: op1_07_in01 = reg_0065;
    78: op1_07_in01 = imem07_in[107:104];
    79: op1_07_in01 = reg_0612;
    80: op1_07_in01 = imem02_in[63:60];
    81: op1_07_in01 = imem00_in[67:64];
    82: op1_07_in01 = imem06_in[51:48];
    83: op1_07_in01 = imem03_in[115:112];
    85: op1_07_in01 = reg_0217;
    86: op1_07_in01 = reg_0154;
    87: op1_07_in01 = reg_0440;
    88: op1_07_in01 = reg_0233;
    89: op1_07_in01 = imem00_in[75:72];
    91: op1_07_in01 = imem00_in[123:120];
    92: op1_07_in01 = reg_0372;
    93: op1_07_in01 = reg_0591;
    95: op1_07_in01 = imem04_in[15:12];
    96: op1_07_in01 = reg_0642;
    default: op1_07_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv01 = 1;
    5: op1_07_inv01 = 1;
    8: op1_07_inv01 = 1;
    11: op1_07_inv01 = 1;
    13: op1_07_inv01 = 1;
    3: op1_07_inv01 = 1;
    15: op1_07_inv01 = 1;
    17: op1_07_inv01 = 1;
    19: op1_07_inv01 = 1;
    22: op1_07_inv01 = 1;
    23: op1_07_inv01 = 1;
    1: op1_07_inv01 = 1;
    26: op1_07_inv01 = 1;
    33: op1_07_inv01 = 1;
    34: op1_07_inv01 = 1;
    35: op1_07_inv01 = 1;
    36: op1_07_inv01 = 1;
    38: op1_07_inv01 = 1;
    39: op1_07_inv01 = 1;
    40: op1_07_inv01 = 1;
    41: op1_07_inv01 = 1;
    43: op1_07_inv01 = 1;
    45: op1_07_inv01 = 1;
    47: op1_07_inv01 = 1;
    48: op1_07_inv01 = 1;
    49: op1_07_inv01 = 1;
    50: op1_07_inv01 = 1;
    51: op1_07_inv01 = 1;
    52: op1_07_inv01 = 1;
    54: op1_07_inv01 = 1;
    57: op1_07_inv01 = 1;
    60: op1_07_inv01 = 1;
    66: op1_07_inv01 = 1;
    67: op1_07_inv01 = 1;
    69: op1_07_inv01 = 1;
    72: op1_07_inv01 = 1;
    73: op1_07_inv01 = 1;
    74: op1_07_inv01 = 1;
    75: op1_07_inv01 = 1;
    76: op1_07_inv01 = 1;
    79: op1_07_inv01 = 1;
    80: op1_07_inv01 = 1;
    85: op1_07_inv01 = 1;
    86: op1_07_inv01 = 1;
    87: op1_07_inv01 = 1;
    91: op1_07_inv01 = 1;
    92: op1_07_inv01 = 1;
    93: op1_07_inv01 = 1;
    95: op1_07_inv01 = 1;
    default: op1_07_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in02 = reg_0009;
    21: op1_07_in02 = reg_0009;
    94: op1_07_in02 = reg_0009;
    5: op1_07_in02 = reg_0109;
    6: op1_07_in02 = reg_0241;
    7: op1_07_in02 = imem00_in[35:32];
    45: op1_07_in02 = imem00_in[35:32];
    66: op1_07_in02 = imem00_in[35:32];
    8: op1_07_in02 = imem03_in[107:104];
    9: op1_07_in02 = imem01_in[115:112];
    10: op1_07_in02 = reg_0002;
    43: op1_07_in02 = reg_0002;
    11: op1_07_in02 = reg_0518;
    12: op1_07_in02 = reg_0623;
    13: op1_07_in02 = imem00_in[55:52];
    3: op1_07_in02 = reg_0438;
    14: op1_07_in02 = reg_0248;
    15: op1_07_in02 = imem05_in[87:84];
    16: op1_07_in02 = reg_0604;
    17: op1_07_in02 = reg_0539;
    18: op1_07_in02 = imem07_in[75:72];
    19: op1_07_in02 = imem04_in[51:48];
    20: op1_07_in02 = imem07_in[119:116];
    78: op1_07_in02 = imem07_in[119:116];
    2: op1_07_in02 = imem07_in[111:108];
    22: op1_07_in02 = reg_0391;
    23: op1_07_in02 = reg_0352;
    24: op1_07_in02 = reg_0290;
    1: op1_07_in02 = imem07_in[83:80];
    25: op1_07_in02 = imem00_in[127:124];
    41: op1_07_in02 = imem00_in[127:124];
    26: op1_07_in02 = imem05_in[47:44];
    27: op1_07_in02 = imem06_in[103:100];
    28: op1_07_in02 = reg_0811;
    29: op1_07_in02 = reg_0273;
    30: op1_07_in02 = reg_0404;
    31: op1_07_in02 = reg_0105;
    32: op1_07_in02 = reg_0770;
    33: op1_07_in02 = reg_0488;
    34: op1_07_in02 = reg_0513;
    35: op1_07_in02 = imem00_in[107:104];
    36: op1_07_in02 = reg_0119;
    37: op1_07_in02 = reg_0771;
    38: op1_07_in02 = reg_0012;
    39: op1_07_in02 = reg_0794;
    40: op1_07_in02 = reg_0560;
    42: op1_07_in02 = imem02_in[3:0];
    44: op1_07_in02 = imem07_in[55:52];
    46: op1_07_in02 = reg_0575;
    47: op1_07_in02 = reg_0317;
    48: op1_07_in02 = imem00_in[71:68];
    49: op1_07_in02 = reg_0707;
    50: op1_07_in02 = imem06_in[23:20];
    51: op1_07_in02 = imem04_in[11:8];
    52: op1_07_in02 = reg_0495;
    53: op1_07_in02 = reg_0371;
    54: op1_07_in02 = reg_0715;
    55: op1_07_in02 = reg_0178;
    56: op1_07_in02 = imem00_in[119:116];
    57: op1_07_in02 = reg_0825;
    58: op1_07_in02 = reg_0683;
    59: op1_07_in02 = reg_0594;
    60: op1_07_in02 = reg_0294;
    61: op1_07_in02 = reg_0561;
    62: op1_07_in02 = reg_0705;
    63: op1_07_in02 = reg_0728;
    64: op1_07_in02 = imem00_in[59:56];
    65: op1_07_in02 = imem00_in[83:80];
    84: op1_07_in02 = imem00_in[83:80];
    67: op1_07_in02 = reg_0361;
    68: op1_07_in02 = reg_0374;
    69: op1_07_in02 = imem00_in[111:108];
    70: op1_07_in02 = reg_0603;
    72: op1_07_in02 = imem00_in[91:88];
    73: op1_07_in02 = imem00_in[51:48];
    74: op1_07_in02 = imem02_in[23:20];
    75: op1_07_in02 = imem04_in[91:88];
    76: op1_07_in02 = reg_0802;
    77: op1_07_in02 = reg_0774;
    79: op1_07_in02 = reg_0690;
    80: op1_07_in02 = reg_0045;
    81: op1_07_in02 = imem00_in[103:100];
    82: op1_07_in02 = imem06_in[115:112];
    83: op1_07_in02 = reg_0347;
    85: op1_07_in02 = reg_0502;
    86: op1_07_in02 = reg_0829;
    87: op1_07_in02 = reg_0442;
    88: op1_07_in02 = imem05_in[19:16];
    89: op1_07_in02 = imem00_in[95:92];
    90: op1_07_in02 = imem00_in[11:8];
    91: op1_07_in02 = reg_0697;
    92: op1_07_in02 = reg_0398;
    93: op1_07_in02 = reg_0318;
    95: op1_07_in02 = imem04_in[107:104];
    96: op1_07_in02 = reg_0081;
    default: op1_07_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_07_inv02 = 1;
    13: op1_07_inv02 = 1;
    15: op1_07_inv02 = 1;
    17: op1_07_inv02 = 1;
    18: op1_07_inv02 = 1;
    19: op1_07_inv02 = 1;
    20: op1_07_inv02 = 1;
    22: op1_07_inv02 = 1;
    23: op1_07_inv02 = 1;
    26: op1_07_inv02 = 1;
    27: op1_07_inv02 = 1;
    29: op1_07_inv02 = 1;
    33: op1_07_inv02 = 1;
    34: op1_07_inv02 = 1;
    37: op1_07_inv02 = 1;
    45: op1_07_inv02 = 1;
    51: op1_07_inv02 = 1;
    52: op1_07_inv02 = 1;
    54: op1_07_inv02 = 1;
    56: op1_07_inv02 = 1;
    57: op1_07_inv02 = 1;
    59: op1_07_inv02 = 1;
    62: op1_07_inv02 = 1;
    63: op1_07_inv02 = 1;
    64: op1_07_inv02 = 1;
    66: op1_07_inv02 = 1;
    68: op1_07_inv02 = 1;
    70: op1_07_inv02 = 1;
    73: op1_07_inv02 = 1;
    77: op1_07_inv02 = 1;
    81: op1_07_inv02 = 1;
    84: op1_07_inv02 = 1;
    92: op1_07_inv02 = 1;
    93: op1_07_inv02 = 1;
    94: op1_07_inv02 = 1;
    default: op1_07_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in03 = reg_0010;
    5: op1_07_in03 = imem02_in[67:64];
    6: op1_07_in03 = reg_0264;
    7: op1_07_in03 = imem00_in[95:92];
    13: op1_07_in03 = imem00_in[95:92];
    8: op1_07_in03 = reg_0579;
    9: op1_07_in03 = imem01_in[123:120];
    10: op1_07_in03 = reg_0800;
    11: op1_07_in03 = reg_0225;
    12: op1_07_in03 = reg_0612;
    3: op1_07_in03 = reg_0159;
    14: op1_07_in03 = reg_0238;
    15: op1_07_in03 = imem05_in[115:112];
    16: op1_07_in03 = reg_0605;
    17: op1_07_in03 = reg_0546;
    18: op1_07_in03 = imem07_in[115:112];
    19: op1_07_in03 = imem04_in[71:68];
    51: op1_07_in03 = imem04_in[71:68];
    20: op1_07_in03 = reg_0720;
    2: op1_07_in03 = reg_0179;
    21: op1_07_in03 = reg_0262;
    22: op1_07_in03 = reg_0343;
    23: op1_07_in03 = reg_0333;
    24: op1_07_in03 = reg_0292;
    1: op1_07_in03 = imem07_in[111:108];
    25: op1_07_in03 = reg_0679;
    26: op1_07_in03 = imem05_in[83:80];
    27: op1_07_in03 = imem06_in[111:108];
    28: op1_07_in03 = reg_0001;
    29: op1_07_in03 = reg_0534;
    30: op1_07_in03 = reg_0576;
    31: op1_07_in03 = reg_0114;
    32: op1_07_in03 = reg_0531;
    33: op1_07_in03 = reg_0789;
    34: op1_07_in03 = reg_0337;
    35: op1_07_in03 = imem00_in[115:112];
    36: op1_07_in03 = reg_0102;
    37: op1_07_in03 = reg_0515;
    38: op1_07_in03 = reg_0003;
    39: op1_07_in03 = reg_0485;
    40: op1_07_in03 = reg_0087;
    41: op1_07_in03 = reg_0695;
    42: op1_07_in03 = imem02_in[15:12];
    43: op1_07_in03 = reg_0805;
    44: op1_07_in03 = imem07_in[123:120];
    45: op1_07_in03 = imem00_in[59:56];
    46: op1_07_in03 = reg_0568;
    47: op1_07_in03 = reg_0331;
    48: op1_07_in03 = imem00_in[111:108];
    49: op1_07_in03 = reg_0727;
    50: op1_07_in03 = imem06_in[55:52];
    52: op1_07_in03 = reg_0790;
    53: op1_07_in03 = reg_0265;
    54: op1_07_in03 = reg_0706;
    55: op1_07_in03 = reg_0170;
    56: op1_07_in03 = reg_0696;
    57: op1_07_in03 = reg_0734;
    58: op1_07_in03 = reg_0694;
    59: op1_07_in03 = reg_0324;
    60: op1_07_in03 = reg_0122;
    61: op1_07_in03 = reg_0564;
    62: op1_07_in03 = reg_0447;
    63: op1_07_in03 = reg_0716;
    64: op1_07_in03 = imem00_in[107:104];
    65: op1_07_in03 = imem00_in[103:100];
    72: op1_07_in03 = imem00_in[103:100];
    84: op1_07_in03 = imem00_in[103:100];
    66: op1_07_in03 = imem00_in[39:36];
    90: op1_07_in03 = imem00_in[39:36];
    67: op1_07_in03 = reg_0406;
    68: op1_07_in03 = reg_0322;
    69: op1_07_in03 = reg_0749;
    70: op1_07_in03 = reg_0234;
    73: op1_07_in03 = imem00_in[99:96];
    74: op1_07_in03 = imem02_in[31:28];
    75: op1_07_in03 = imem04_in[95:92];
    76: op1_07_in03 = reg_0009;
    93: op1_07_in03 = reg_0009;
    77: op1_07_in03 = reg_0416;
    78: op1_07_in03 = reg_0441;
    79: op1_07_in03 = reg_0407;
    80: op1_07_in03 = reg_0141;
    81: op1_07_in03 = imem00_in[123:120];
    82: op1_07_in03 = imem06_in[127:124];
    83: op1_07_in03 = reg_0317;
    85: op1_07_in03 = reg_0216;
    86: op1_07_in03 = reg_0824;
    87: op1_07_in03 = reg_0084;
    88: op1_07_in03 = imem05_in[47:44];
    89: op1_07_in03 = reg_0685;
    91: op1_07_in03 = reg_0686;
    92: op1_07_in03 = reg_0186;
    94: op1_07_in03 = reg_0595;
    95: op1_07_in03 = imem04_in[123:120];
    96: op1_07_in03 = reg_0056;
    default: op1_07_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv03 = 1;
    7: op1_07_inv03 = 1;
    8: op1_07_inv03 = 1;
    10: op1_07_inv03 = 1;
    11: op1_07_inv03 = 1;
    12: op1_07_inv03 = 1;
    13: op1_07_inv03 = 1;
    3: op1_07_inv03 = 1;
    14: op1_07_inv03 = 1;
    15: op1_07_inv03 = 1;
    16: op1_07_inv03 = 1;
    17: op1_07_inv03 = 1;
    18: op1_07_inv03 = 1;
    19: op1_07_inv03 = 1;
    2: op1_07_inv03 = 1;
    22: op1_07_inv03 = 1;
    24: op1_07_inv03 = 1;
    1: op1_07_inv03 = 1;
    25: op1_07_inv03 = 1;
    27: op1_07_inv03 = 1;
    30: op1_07_inv03 = 1;
    33: op1_07_inv03 = 1;
    35: op1_07_inv03 = 1;
    36: op1_07_inv03 = 1;
    39: op1_07_inv03 = 1;
    40: op1_07_inv03 = 1;
    42: op1_07_inv03 = 1;
    47: op1_07_inv03 = 1;
    49: op1_07_inv03 = 1;
    50: op1_07_inv03 = 1;
    51: op1_07_inv03 = 1;
    54: op1_07_inv03 = 1;
    55: op1_07_inv03 = 1;
    59: op1_07_inv03 = 1;
    60: op1_07_inv03 = 1;
    61: op1_07_inv03 = 1;
    62: op1_07_inv03 = 1;
    63: op1_07_inv03 = 1;
    65: op1_07_inv03 = 1;
    66: op1_07_inv03 = 1;
    68: op1_07_inv03 = 1;
    69: op1_07_inv03 = 1;
    70: op1_07_inv03 = 1;
    75: op1_07_inv03 = 1;
    77: op1_07_inv03 = 1;
    79: op1_07_inv03 = 1;
    80: op1_07_inv03 = 1;
    81: op1_07_inv03 = 1;
    82: op1_07_inv03 = 1;
    83: op1_07_inv03 = 1;
    84: op1_07_inv03 = 1;
    85: op1_07_inv03 = 1;
    87: op1_07_inv03 = 1;
    89: op1_07_inv03 = 1;
    95: op1_07_inv03 = 1;
    default: op1_07_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in04 = reg_0004;
    5: op1_07_in04 = imem02_in[91:88];
    6: op1_07_in04 = reg_0251;
    7: op1_07_in04 = reg_0682;
    8: op1_07_in04 = reg_0572;
    9: op1_07_in04 = reg_0108;
    10: op1_07_in04 = reg_0799;
    11: op1_07_in04 = reg_0235;
    12: op1_07_in04 = reg_0344;
    13: op1_07_in04 = reg_0679;
    3: op1_07_in04 = reg_0173;
    14: op1_07_in04 = reg_0219;
    15: op1_07_in04 = imem05_in[119:116];
    26: op1_07_in04 = imem05_in[119:116];
    16: op1_07_in04 = reg_0621;
    17: op1_07_in04 = reg_0532;
    18: op1_07_in04 = imem07_in[123:120];
    19: op1_07_in04 = imem04_in[111:108];
    20: op1_07_in04 = reg_0701;
    2: op1_07_in04 = reg_0183;
    21: op1_07_in04 = reg_0536;
    22: op1_07_in04 = reg_0362;
    23: op1_07_in04 = reg_0359;
    24: op1_07_in04 = reg_0298;
    25: op1_07_in04 = reg_0668;
    27: op1_07_in04 = reg_0577;
    28: op1_07_in04 = reg_0801;
    29: op1_07_in04 = reg_0290;
    30: op1_07_in04 = reg_0817;
    31: op1_07_in04 = reg_0106;
    32: op1_07_in04 = imem03_in[3:0];
    33: op1_07_in04 = reg_0492;
    34: op1_07_in04 = reg_0514;
    35: op1_07_in04 = imem00_in[119:116];
    84: op1_07_in04 = imem00_in[119:116];
    36: op1_07_in04 = reg_0114;
    37: op1_07_in04 = reg_0557;
    38: op1_07_in04 = reg_0807;
    39: op1_07_in04 = reg_0271;
    40: op1_07_in04 = reg_0547;
    41: op1_07_in04 = reg_0670;
    42: op1_07_in04 = imem02_in[31:28];
    43: op1_07_in04 = reg_0015;
    44: op1_07_in04 = reg_0716;
    45: op1_07_in04 = imem00_in[63:60];
    46: op1_07_in04 = reg_0388;
    47: op1_07_in04 = reg_0407;
    48: op1_07_in04 = reg_0681;
    49: op1_07_in04 = reg_0636;
    50: op1_07_in04 = imem06_in[59:56];
    51: op1_07_in04 = imem04_in[107:104];
    52: op1_07_in04 = reg_0787;
    53: op1_07_in04 = reg_0318;
    54: op1_07_in04 = reg_0441;
    55: op1_07_in04 = reg_0176;
    56: op1_07_in04 = reg_0744;
    89: op1_07_in04 = reg_0744;
    57: op1_07_in04 = reg_0321;
    58: op1_07_in04 = reg_0634;
    59: op1_07_in04 = reg_0527;
    60: op1_07_in04 = reg_0118;
    61: op1_07_in04 = reg_0392;
    62: op1_07_in04 = reg_0445;
    63: op1_07_in04 = reg_0731;
    64: op1_07_in04 = reg_0693;
    65: op1_07_in04 = imem00_in[111:108];
    66: op1_07_in04 = imem00_in[51:48];
    67: op1_07_in04 = reg_0314;
    68: op1_07_in04 = reg_0386;
    69: op1_07_in04 = reg_0117;
    70: op1_07_in04 = reg_0506;
    72: op1_07_in04 = reg_0695;
    73: op1_07_in04 = imem00_in[123:120];
    74: op1_07_in04 = imem02_in[47:44];
    75: op1_07_in04 = imem04_in[103:100];
    76: op1_07_in04 = reg_0010;
    77: op1_07_in04 = imem05_in[91:88];
    78: op1_07_in04 = reg_0175;
    79: op1_07_in04 = reg_0699;
    80: op1_07_in04 = reg_0374;
    81: op1_07_in04 = reg_0694;
    82: op1_07_in04 = reg_0115;
    83: op1_07_in04 = reg_0599;
    85: op1_07_in04 = reg_0248;
    86: op1_07_in04 = imem06_in[55:52];
    87: op1_07_in04 = reg_0435;
    88: op1_07_in04 = reg_0792;
    90: op1_07_in04 = imem00_in[59:56];
    91: op1_07_in04 = reg_0691;
    92: op1_07_in04 = reg_0013;
    93: op1_07_in04 = reg_0507;
    94: op1_07_in04 = reg_0648;
    95: op1_07_in04 = reg_0058;
    96: op1_07_in04 = reg_0639;
    default: op1_07_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv04 = 1;
    5: op1_07_inv04 = 1;
    7: op1_07_inv04 = 1;
    11: op1_07_inv04 = 1;
    12: op1_07_inv04 = 1;
    3: op1_07_inv04 = 1;
    14: op1_07_inv04 = 1;
    15: op1_07_inv04 = 1;
    17: op1_07_inv04 = 1;
    19: op1_07_inv04 = 1;
    20: op1_07_inv04 = 1;
    2: op1_07_inv04 = 1;
    22: op1_07_inv04 = 1;
    24: op1_07_inv04 = 1;
    28: op1_07_inv04 = 1;
    29: op1_07_inv04 = 1;
    30: op1_07_inv04 = 1;
    32: op1_07_inv04 = 1;
    33: op1_07_inv04 = 1;
    36: op1_07_inv04 = 1;
    39: op1_07_inv04 = 1;
    41: op1_07_inv04 = 1;
    42: op1_07_inv04 = 1;
    44: op1_07_inv04 = 1;
    46: op1_07_inv04 = 1;
    47: op1_07_inv04 = 1;
    50: op1_07_inv04 = 1;
    56: op1_07_inv04 = 1;
    57: op1_07_inv04 = 1;
    58: op1_07_inv04 = 1;
    59: op1_07_inv04 = 1;
    61: op1_07_inv04 = 1;
    67: op1_07_inv04 = 1;
    69: op1_07_inv04 = 1;
    70: op1_07_inv04 = 1;
    72: op1_07_inv04 = 1;
    75: op1_07_inv04 = 1;
    78: op1_07_inv04 = 1;
    81: op1_07_inv04 = 1;
    84: op1_07_inv04 = 1;
    86: op1_07_inv04 = 1;
    92: op1_07_inv04 = 1;
    94: op1_07_inv04 = 1;
    default: op1_07_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in05 = imem04_in[11:8];
    5: op1_07_in05 = imem02_in[99:96];
    6: op1_07_in05 = reg_0254;
    7: op1_07_in05 = reg_0697;
    8: op1_07_in05 = reg_0569;
    9: op1_07_in05 = reg_0115;
    10: op1_07_in05 = imem04_in[43:40];
    11: op1_07_in05 = reg_0233;
    12: op1_07_in05 = reg_0392;
    46: op1_07_in05 = reg_0392;
    13: op1_07_in05 = reg_0463;
    79: op1_07_in05 = reg_0463;
    14: op1_07_in05 = reg_0123;
    15: op1_07_in05 = imem05_in[123:120];
    16: op1_07_in05 = reg_0616;
    17: op1_07_in05 = reg_0533;
    18: op1_07_in05 = reg_0722;
    19: op1_07_in05 = imem04_in[115:112];
    51: op1_07_in05 = imem04_in[115:112];
    20: op1_07_in05 = reg_0423;
    2: op1_07_in05 = reg_0178;
    21: op1_07_in05 = reg_0264;
    22: op1_07_in05 = reg_0385;
    23: op1_07_in05 = reg_0330;
    24: op1_07_in05 = reg_0284;
    25: op1_07_in05 = reg_0699;
    26: op1_07_in05 = reg_0484;
    27: op1_07_in05 = reg_0622;
    28: op1_07_in05 = reg_0008;
    29: op1_07_in05 = reg_0291;
    30: op1_07_in05 = reg_0819;
    31: op1_07_in05 = reg_0126;
    32: op1_07_in05 = imem03_in[7:4];
    33: op1_07_in05 = reg_0783;
    34: op1_07_in05 = reg_0820;
    35: op1_07_in05 = reg_0689;
    36: op1_07_in05 = reg_0107;
    37: op1_07_in05 = reg_0760;
    38: op1_07_in05 = reg_0801;
    39: op1_07_in05 = reg_0304;
    40: op1_07_in05 = reg_0283;
    41: op1_07_in05 = reg_0678;
    42: op1_07_in05 = reg_0655;
    43: op1_07_in05 = imem04_in[35:32];
    44: op1_07_in05 = reg_0731;
    45: op1_07_in05 = imem00_in[107:104];
    47: op1_07_in05 = reg_0607;
    48: op1_07_in05 = reg_0686;
    84: op1_07_in05 = reg_0686;
    49: op1_07_in05 = reg_0447;
    50: op1_07_in05 = imem06_in[71:68];
    52: op1_07_in05 = reg_0489;
    53: op1_07_in05 = reg_0369;
    54: op1_07_in05 = reg_0295;
    56: op1_07_in05 = reg_0690;
    57: op1_07_in05 = reg_0421;
    58: op1_07_in05 = reg_0476;
    59: op1_07_in05 = reg_0541;
    60: op1_07_in05 = reg_0592;
    61: op1_07_in05 = reg_0019;
    62: op1_07_in05 = reg_0449;
    63: op1_07_in05 = reg_0718;
    64: op1_07_in05 = reg_0612;
    65: op1_07_in05 = reg_0696;
    66: op1_07_in05 = imem00_in[67:64];
    67: op1_07_in05 = imem03_in[3:0];
    68: op1_07_in05 = reg_0326;
    69: op1_07_in05 = reg_0407;
    70: op1_07_in05 = reg_0419;
    72: op1_07_in05 = reg_0698;
    73: op1_07_in05 = reg_0685;
    74: op1_07_in05 = imem02_in[83:80];
    75: op1_07_in05 = reg_0545;
    76: op1_07_in05 = reg_0809;
    77: op1_07_in05 = imem05_in[99:96];
    78: op1_07_in05 = reg_0169;
    80: op1_07_in05 = reg_0485;
    81: op1_07_in05 = reg_0658;
    82: op1_07_in05 = reg_0404;
    83: op1_07_in05 = reg_0604;
    85: op1_07_in05 = reg_0424;
    86: op1_07_in05 = imem06_in[99:96];
    87: op1_07_in05 = reg_0139;
    88: op1_07_in05 = reg_0666;
    89: op1_07_in05 = reg_0691;
    90: op1_07_in05 = imem00_in[75:72];
    91: op1_07_in05 = reg_0145;
    92: op1_07_in05 = reg_0244;
    93: op1_07_in05 = reg_0028;
    94: op1_07_in05 = reg_0321;
    95: op1_07_in05 = reg_0555;
    96: op1_07_in05 = reg_0705;
    default: op1_07_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_07_inv05 = 1;
    10: op1_07_inv05 = 1;
    11: op1_07_inv05 = 1;
    14: op1_07_inv05 = 1;
    15: op1_07_inv05 = 1;
    16: op1_07_inv05 = 1;
    17: op1_07_inv05 = 1;
    18: op1_07_inv05 = 1;
    19: op1_07_inv05 = 1;
    21: op1_07_inv05 = 1;
    22: op1_07_inv05 = 1;
    23: op1_07_inv05 = 1;
    26: op1_07_inv05 = 1;
    27: op1_07_inv05 = 1;
    29: op1_07_inv05 = 1;
    30: op1_07_inv05 = 1;
    31: op1_07_inv05 = 1;
    33: op1_07_inv05 = 1;
    34: op1_07_inv05 = 1;
    35: op1_07_inv05 = 1;
    36: op1_07_inv05 = 1;
    37: op1_07_inv05 = 1;
    41: op1_07_inv05 = 1;
    42: op1_07_inv05 = 1;
    45: op1_07_inv05 = 1;
    49: op1_07_inv05 = 1;
    50: op1_07_inv05 = 1;
    51: op1_07_inv05 = 1;
    53: op1_07_inv05 = 1;
    58: op1_07_inv05 = 1;
    59: op1_07_inv05 = 1;
    63: op1_07_inv05 = 1;
    64: op1_07_inv05 = 1;
    65: op1_07_inv05 = 1;
    66: op1_07_inv05 = 1;
    69: op1_07_inv05 = 1;
    72: op1_07_inv05 = 1;
    75: op1_07_inv05 = 1;
    78: op1_07_inv05 = 1;
    79: op1_07_inv05 = 1;
    80: op1_07_inv05 = 1;
    81: op1_07_inv05 = 1;
    84: op1_07_inv05 = 1;
    89: op1_07_inv05 = 1;
    91: op1_07_inv05 = 1;
    92: op1_07_inv05 = 1;
    95: op1_07_inv05 = 1;
    96: op1_07_inv05 = 1;
    default: op1_07_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in06 = imem04_in[31:28];
    5: op1_07_in06 = imem02_in[119:116];
    6: op1_07_in06 = reg_0148;
    7: op1_07_in06 = reg_0681;
    8: op1_07_in06 = reg_0600;
    9: op1_07_in06 = reg_0109;
    10: op1_07_in06 = reg_0536;
    11: op1_07_in06 = reg_0506;
    12: op1_07_in06 = reg_0390;
    13: op1_07_in06 = reg_0461;
    14: op1_07_in06 = reg_0124;
    15: op1_07_in06 = reg_0797;
    16: op1_07_in06 = reg_0626;
    17: op1_07_in06 = reg_0531;
    18: op1_07_in06 = reg_0719;
    19: op1_07_in06 = reg_0545;
    20: op1_07_in06 = reg_0428;
    21: op1_07_in06 = reg_0542;
    22: op1_07_in06 = reg_0322;
    23: op1_07_in06 = reg_0346;
    24: op1_07_in06 = reg_0281;
    25: op1_07_in06 = reg_0455;
    26: op1_07_in06 = reg_0491;
    27: op1_07_in06 = reg_0601;
    28: op1_07_in06 = reg_0799;
    29: op1_07_in06 = reg_0298;
    30: op1_07_in06 = imem07_in[71:68];
    31: op1_07_in06 = imem02_in[75:72];
    32: op1_07_in06 = imem03_in[27:24];
    33: op1_07_in06 = reg_0784;
    34: op1_07_in06 = reg_0227;
    35: op1_07_in06 = reg_0684;
    73: op1_07_in06 = reg_0684;
    36: op1_07_in06 = reg_0121;
    37: op1_07_in06 = reg_0505;
    38: op1_07_in06 = imem04_in[19:16];
    39: op1_07_in06 = reg_0309;
    52: op1_07_in06 = reg_0309;
    40: op1_07_in06 = reg_0292;
    41: op1_07_in06 = reg_0688;
    84: op1_07_in06 = reg_0688;
    42: op1_07_in06 = reg_0653;
    43: op1_07_in06 = imem04_in[83:80];
    44: op1_07_in06 = reg_0714;
    45: op1_07_in06 = imem00_in[111:108];
    46: op1_07_in06 = reg_0499;
    47: op1_07_in06 = reg_0620;
    48: op1_07_in06 = reg_0677;
    49: op1_07_in06 = reg_0061;
    63: op1_07_in06 = reg_0061;
    50: op1_07_in06 = imem06_in[87:84];
    51: op1_07_in06 = reg_0316;
    53: op1_07_in06 = reg_0331;
    54: op1_07_in06 = reg_0439;
    56: op1_07_in06 = reg_0658;
    57: op1_07_in06 = reg_0418;
    58: op1_07_in06 = reg_0466;
    59: op1_07_in06 = reg_0314;
    60: op1_07_in06 = reg_0676;
    61: op1_07_in06 = reg_0002;
    62: op1_07_in06 = reg_0442;
    64: op1_07_in06 = reg_0633;
    65: op1_07_in06 = reg_0612;
    66: op1_07_in06 = imem00_in[83:80];
    67: op1_07_in06 = imem03_in[11:8];
    68: op1_07_in06 = reg_0246;
    69: op1_07_in06 = reg_0477;
    70: op1_07_in06 = reg_0105;
    72: op1_07_in06 = reg_0690;
    74: op1_07_in06 = imem02_in[127:124];
    75: op1_07_in06 = reg_0553;
    76: op1_07_in06 = imem04_in[67:64];
    77: op1_07_in06 = reg_0791;
    78: op1_07_in06 = reg_0177;
    79: op1_07_in06 = reg_0450;
    80: op1_07_in06 = reg_0320;
    81: op1_07_in06 = reg_0117;
    82: op1_07_in06 = reg_0659;
    83: op1_07_in06 = reg_0338;
    85: op1_07_in06 = reg_0119;
    86: op1_07_in06 = imem06_in[103:100];
    87: op1_07_in06 = reg_0089;
    88: op1_07_in06 = reg_0355;
    89: op1_07_in06 = reg_0451;
    90: op1_07_in06 = imem00_in[87:84];
    91: op1_07_in06 = reg_0460;
    92: op1_07_in06 = imem04_in[11:8];
    93: op1_07_in06 = reg_0321;
    94: op1_07_in06 = reg_0575;
    95: op1_07_in06 = reg_0174;
    96: op1_07_in06 = reg_0274;
    default: op1_07_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv06 = 1;
    5: op1_07_inv06 = 1;
    7: op1_07_inv06 = 1;
    8: op1_07_inv06 = 1;
    9: op1_07_inv06 = 1;
    11: op1_07_inv06 = 1;
    12: op1_07_inv06 = 1;
    13: op1_07_inv06 = 1;
    15: op1_07_inv06 = 1;
    16: op1_07_inv06 = 1;
    18: op1_07_inv06 = 1;
    19: op1_07_inv06 = 1;
    23: op1_07_inv06 = 1;
    24: op1_07_inv06 = 1;
    29: op1_07_inv06 = 1;
    30: op1_07_inv06 = 1;
    31: op1_07_inv06 = 1;
    32: op1_07_inv06 = 1;
    33: op1_07_inv06 = 1;
    35: op1_07_inv06 = 1;
    36: op1_07_inv06 = 1;
    37: op1_07_inv06 = 1;
    39: op1_07_inv06 = 1;
    41: op1_07_inv06 = 1;
    42: op1_07_inv06 = 1;
    44: op1_07_inv06 = 1;
    47: op1_07_inv06 = 1;
    50: op1_07_inv06 = 1;
    51: op1_07_inv06 = 1;
    52: op1_07_inv06 = 1;
    57: op1_07_inv06 = 1;
    58: op1_07_inv06 = 1;
    59: op1_07_inv06 = 1;
    60: op1_07_inv06 = 1;
    62: op1_07_inv06 = 1;
    65: op1_07_inv06 = 1;
    66: op1_07_inv06 = 1;
    67: op1_07_inv06 = 1;
    69: op1_07_inv06 = 1;
    72: op1_07_inv06 = 1;
    74: op1_07_inv06 = 1;
    80: op1_07_inv06 = 1;
    81: op1_07_inv06 = 1;
    82: op1_07_inv06 = 1;
    83: op1_07_inv06 = 1;
    84: op1_07_inv06 = 1;
    86: op1_07_inv06 = 1;
    87: op1_07_inv06 = 1;
    89: op1_07_inv06 = 1;
    90: op1_07_inv06 = 1;
    92: op1_07_inv06 = 1;
    93: op1_07_inv06 = 1;
    94: op1_07_inv06 = 1;
    96: op1_07_inv06 = 1;
    default: op1_07_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in07 = imem04_in[59:56];
    5: op1_07_in07 = reg_0658;
    65: op1_07_in07 = reg_0658;
    6: op1_07_in07 = reg_0145;
    7: op1_07_in07 = reg_0698;
    8: op1_07_in07 = reg_0581;
    9: op1_07_in07 = reg_0126;
    10: op1_07_in07 = reg_0553;
    11: op1_07_in07 = reg_0217;
    57: op1_07_in07 = reg_0217;
    12: op1_07_in07 = reg_0037;
    13: op1_07_in07 = reg_0466;
    14: op1_07_in07 = reg_0116;
    15: op1_07_in07 = reg_0781;
    16: op1_07_in07 = reg_0619;
    17: op1_07_in07 = reg_0556;
    18: op1_07_in07 = reg_0720;
    19: op1_07_in07 = reg_0542;
    20: op1_07_in07 = reg_0434;
    21: op1_07_in07 = imem04_in[19:16];
    92: op1_07_in07 = imem04_in[19:16];
    22: op1_07_in07 = reg_0323;
    23: op1_07_in07 = reg_0338;
    24: op1_07_in07 = reg_0079;
    25: op1_07_in07 = reg_0472;
    26: op1_07_in07 = reg_0492;
    27: op1_07_in07 = reg_0402;
    28: op1_07_in07 = reg_0004;
    29: op1_07_in07 = reg_0299;
    30: op1_07_in07 = imem07_in[91:88];
    31: op1_07_in07 = imem02_in[79:76];
    32: op1_07_in07 = imem03_in[35:32];
    33: op1_07_in07 = reg_0485;
    34: op1_07_in07 = reg_0549;
    35: op1_07_in07 = reg_0679;
    36: op1_07_in07 = imem02_in[39:36];
    37: op1_07_in07 = reg_0246;
    38: op1_07_in07 = imem04_in[27:24];
    39: op1_07_in07 = reg_0737;
    40: op1_07_in07 = reg_0256;
    41: op1_07_in07 = reg_0692;
    42: op1_07_in07 = reg_0661;
    43: op1_07_in07 = reg_0315;
    44: op1_07_in07 = reg_0724;
    45: op1_07_in07 = reg_0682;
    46: op1_07_in07 = reg_0396;
    47: op1_07_in07 = imem07_in[7:4];
    48: op1_07_in07 = reg_0671;
    49: op1_07_in07 = reg_0333;
    50: op1_07_in07 = reg_0604;
    51: op1_07_in07 = reg_0544;
    52: op1_07_in07 = reg_0245;
    53: op1_07_in07 = reg_0329;
    54: op1_07_in07 = reg_0443;
    56: op1_07_in07 = reg_0680;
    58: op1_07_in07 = reg_0467;
    59: op1_07_in07 = reg_0743;
    60: op1_07_in07 = imem02_in[19:16];
    61: op1_07_in07 = reg_0801;
    62: op1_07_in07 = reg_0180;
    63: op1_07_in07 = reg_0448;
    64: op1_07_in07 = reg_0455;
    66: op1_07_in07 = imem00_in[99:96];
    90: op1_07_in07 = imem00_in[99:96];
    67: op1_07_in07 = imem03_in[67:64];
    68: op1_07_in07 = reg_0491;
    69: op1_07_in07 = reg_0476;
    79: op1_07_in07 = reg_0476;
    70: op1_07_in07 = reg_0073;
    72: op1_07_in07 = reg_0477;
    73: op1_07_in07 = reg_0255;
    74: op1_07_in07 = reg_0392;
    75: op1_07_in07 = reg_0056;
    76: op1_07_in07 = imem04_in[83:80];
    77: op1_07_in07 = reg_0641;
    78: op1_07_in07 = reg_0168;
    80: op1_07_in07 = reg_0341;
    81: op1_07_in07 = reg_0247;
    82: op1_07_in07 = reg_0375;
    83: op1_07_in07 = reg_0319;
    84: op1_07_in07 = reg_0634;
    85: op1_07_in07 = reg_0669;
    86: op1_07_in07 = reg_0348;
    87: op1_07_in07 = reg_0236;
    88: op1_07_in07 = reg_0732;
    89: op1_07_in07 = reg_0470;
    91: op1_07_in07 = reg_0480;
    93: op1_07_in07 = reg_0186;
    94: op1_07_in07 = reg_0372;
    95: op1_07_in07 = reg_0615;
    96: op1_07_in07 = reg_0059;
    default: op1_07_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv07 = 1;
    11: op1_07_inv07 = 1;
    12: op1_07_inv07 = 1;
    15: op1_07_inv07 = 1;
    19: op1_07_inv07 = 1;
    22: op1_07_inv07 = 1;
    25: op1_07_inv07 = 1;
    27: op1_07_inv07 = 1;
    29: op1_07_inv07 = 1;
    31: op1_07_inv07 = 1;
    32: op1_07_inv07 = 1;
    34: op1_07_inv07 = 1;
    36: op1_07_inv07 = 1;
    40: op1_07_inv07 = 1;
    44: op1_07_inv07 = 1;
    45: op1_07_inv07 = 1;
    46: op1_07_inv07 = 1;
    48: op1_07_inv07 = 1;
    50: op1_07_inv07 = 1;
    53: op1_07_inv07 = 1;
    57: op1_07_inv07 = 1;
    61: op1_07_inv07 = 1;
    62: op1_07_inv07 = 1;
    67: op1_07_inv07 = 1;
    70: op1_07_inv07 = 1;
    72: op1_07_inv07 = 1;
    75: op1_07_inv07 = 1;
    78: op1_07_inv07 = 1;
    79: op1_07_inv07 = 1;
    80: op1_07_inv07 = 1;
    82: op1_07_inv07 = 1;
    84: op1_07_inv07 = 1;
    90: op1_07_inv07 = 1;
    92: op1_07_inv07 = 1;
    95: op1_07_inv07 = 1;
    default: op1_07_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in08 = imem04_in[67:64];
    5: op1_07_in08 = reg_0654;
    6: op1_07_in08 = reg_0143;
    7: op1_07_in08 = reg_0670;
    8: op1_07_in08 = reg_0595;
    9: op1_07_in08 = reg_0110;
    10: op1_07_in08 = reg_0550;
    11: op1_07_in08 = reg_0237;
    12: op1_07_in08 = reg_0029;
    13: op1_07_in08 = reg_0460;
    79: op1_07_in08 = reg_0460;
    14: op1_07_in08 = reg_0101;
    15: op1_07_in08 = reg_0489;
    16: op1_07_in08 = reg_0608;
    17: op1_07_in08 = reg_0303;
    18: op1_07_in08 = reg_0729;
    44: op1_07_in08 = reg_0729;
    19: op1_07_in08 = reg_0554;
    20: op1_07_in08 = reg_0444;
    21: op1_07_in08 = imem04_in[27:24];
    22: op1_07_in08 = reg_0019;
    23: op1_07_in08 = reg_0355;
    24: op1_07_in08 = reg_0067;
    25: op1_07_in08 = reg_0467;
    91: op1_07_in08 = reg_0467;
    26: op1_07_in08 = reg_0785;
    27: op1_07_in08 = reg_0404;
    28: op1_07_in08 = imem04_in[11:8];
    29: op1_07_in08 = reg_0064;
    30: op1_07_in08 = imem07_in[95:92];
    31: op1_07_in08 = imem02_in[91:88];
    32: op1_07_in08 = imem03_in[39:36];
    33: op1_07_in08 = reg_0090;
    34: op1_07_in08 = reg_0333;
    35: op1_07_in08 = reg_0463;
    56: op1_07_in08 = reg_0463;
    36: op1_07_in08 = imem02_in[47:44];
    37: op1_07_in08 = reg_0218;
    38: op1_07_in08 = imem04_in[55:52];
    39: op1_07_in08 = reg_0527;
    40: op1_07_in08 = imem05_in[55:52];
    41: op1_07_in08 = reg_0455;
    81: op1_07_in08 = reg_0455;
    42: op1_07_in08 = reg_0656;
    43: op1_07_in08 = reg_0328;
    45: op1_07_in08 = reg_0693;
    46: op1_07_in08 = reg_0570;
    47: op1_07_in08 = imem07_in[15:12];
    48: op1_07_in08 = reg_0454;
    49: op1_07_in08 = reg_0434;
    50: op1_07_in08 = reg_0291;
    86: op1_07_in08 = reg_0291;
    51: op1_07_in08 = reg_0315;
    52: op1_07_in08 = reg_0258;
    53: op1_07_in08 = reg_0028;
    54: op1_07_in08 = reg_0084;
    57: op1_07_in08 = reg_0567;
    58: op1_07_in08 = reg_0200;
    59: op1_07_in08 = reg_0080;
    60: op1_07_in08 = imem02_in[43:40];
    61: op1_07_in08 = reg_0805;
    62: op1_07_in08 = reg_0181;
    63: op1_07_in08 = reg_0180;
    64: op1_07_in08 = reg_0461;
    65: op1_07_in08 = reg_0255;
    66: op1_07_in08 = reg_0694;
    67: op1_07_in08 = imem03_in[91:88];
    68: op1_07_in08 = reg_0236;
    69: op1_07_in08 = reg_0475;
    70: op1_07_in08 = reg_0660;
    72: op1_07_in08 = reg_0452;
    73: op1_07_in08 = reg_0477;
    74: op1_07_in08 = reg_0139;
    75: op1_07_in08 = reg_0088;
    76: op1_07_in08 = imem04_in[99:96];
    77: op1_07_in08 = reg_0309;
    78: op1_07_in08 = reg_0170;
    80: op1_07_in08 = reg_0565;
    82: op1_07_in08 = reg_0583;
    83: op1_07_in08 = reg_0281;
    84: op1_07_in08 = reg_0457;
    85: op1_07_in08 = reg_0601;
    87: op1_07_in08 = reg_0182;
    88: op1_07_in08 = reg_0226;
    89: op1_07_in08 = reg_0189;
    90: op1_07_in08 = imem00_in[115:112];
    92: op1_07_in08 = imem04_in[51:48];
    93: op1_07_in08 = reg_0271;
    94: op1_07_in08 = reg_0569;
    95: op1_07_in08 = reg_0616;
    96: op1_07_in08 = reg_0251;
    default: op1_07_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv08 = 1;
    7: op1_07_inv08 = 1;
    11: op1_07_inv08 = 1;
    12: op1_07_inv08 = 1;
    13: op1_07_inv08 = 1;
    14: op1_07_inv08 = 1;
    15: op1_07_inv08 = 1;
    17: op1_07_inv08 = 1;
    20: op1_07_inv08 = 1;
    23: op1_07_inv08 = 1;
    24: op1_07_inv08 = 1;
    33: op1_07_inv08 = 1;
    35: op1_07_inv08 = 1;
    36: op1_07_inv08 = 1;
    37: op1_07_inv08 = 1;
    38: op1_07_inv08 = 1;
    39: op1_07_inv08 = 1;
    43: op1_07_inv08 = 1;
    44: op1_07_inv08 = 1;
    47: op1_07_inv08 = 1;
    49: op1_07_inv08 = 1;
    50: op1_07_inv08 = 1;
    51: op1_07_inv08 = 1;
    52: op1_07_inv08 = 1;
    56: op1_07_inv08 = 1;
    57: op1_07_inv08 = 1;
    58: op1_07_inv08 = 1;
    64: op1_07_inv08 = 1;
    65: op1_07_inv08 = 1;
    70: op1_07_inv08 = 1;
    73: op1_07_inv08 = 1;
    74: op1_07_inv08 = 1;
    75: op1_07_inv08 = 1;
    76: op1_07_inv08 = 1;
    79: op1_07_inv08 = 1;
    81: op1_07_inv08 = 1;
    84: op1_07_inv08 = 1;
    85: op1_07_inv08 = 1;
    87: op1_07_inv08 = 1;
    90: op1_07_inv08 = 1;
    93: op1_07_inv08 = 1;
    default: op1_07_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in09 = imem04_in[79:76];
    5: op1_07_in09 = reg_0637;
    6: op1_07_in09 = imem06_in[35:32];
    7: op1_07_in09 = reg_0677;
    8: op1_07_in09 = reg_0360;
    9: op1_07_in09 = imem02_in[3:0];
    10: op1_07_in09 = reg_0531;
    11: op1_07_in09 = reg_0245;
    12: op1_07_in09 = reg_0038;
    13: op1_07_in09 = reg_0481;
    69: op1_07_in09 = reg_0481;
    84: op1_07_in09 = reg_0481;
    14: op1_07_in09 = reg_0109;
    15: op1_07_in09 = reg_0267;
    16: op1_07_in09 = reg_0622;
    17: op1_07_in09 = reg_0305;
    18: op1_07_in09 = reg_0713;
    19: op1_07_in09 = reg_0551;
    20: op1_07_in09 = reg_0438;
    21: op1_07_in09 = imem04_in[51:48];
    22: op1_07_in09 = reg_0013;
    23: op1_07_in09 = reg_0347;
    24: op1_07_in09 = reg_0064;
    25: op1_07_in09 = reg_0479;
    26: op1_07_in09 = reg_0782;
    27: op1_07_in09 = reg_0401;
    28: op1_07_in09 = imem04_in[47:44];
    29: op1_07_in09 = imem05_in[103:100];
    30: op1_07_in09 = imem07_in[127:124];
    31: op1_07_in09 = imem02_in[127:124];
    32: op1_07_in09 = imem03_in[51:48];
    33: op1_07_in09 = reg_0225;
    34: op1_07_in09 = reg_0771;
    35: op1_07_in09 = reg_0464;
    36: op1_07_in09 = imem02_in[87:84];
    37: op1_07_in09 = reg_0239;
    38: op1_07_in09 = imem04_in[127:124];
    39: op1_07_in09 = reg_0085;
    40: op1_07_in09 = imem05_in[87:84];
    41: op1_07_in09 = reg_0466;
    42: op1_07_in09 = reg_0648;
    43: op1_07_in09 = reg_0087;
    44: op1_07_in09 = reg_0711;
    45: op1_07_in09 = reg_0683;
    46: op1_07_in09 = reg_0006;
    47: op1_07_in09 = imem07_in[31:28];
    48: op1_07_in09 = reg_0457;
    49: op1_07_in09 = reg_0444;
    50: op1_07_in09 = reg_0613;
    51: op1_07_in09 = reg_0552;
    52: op1_07_in09 = reg_0277;
    53: op1_07_in09 = reg_0753;
    54: op1_07_in09 = reg_0437;
    56: op1_07_in09 = reg_0450;
    57: op1_07_in09 = reg_0216;
    58: op1_07_in09 = reg_0210;
    59: op1_07_in09 = reg_0530;
    60: op1_07_in09 = imem02_in[51:48];
    61: op1_07_in09 = reg_0010;
    62: op1_07_in09 = reg_0179;
    63: op1_07_in09 = reg_0172;
    64: op1_07_in09 = reg_0469;
    81: op1_07_in09 = reg_0469;
    65: op1_07_in09 = reg_0494;
    66: op1_07_in09 = reg_0690;
    67: op1_07_in09 = imem03_in[95:92];
    68: op1_07_in09 = reg_0132;
    70: op1_07_in09 = reg_0675;
    72: op1_07_in09 = reg_0456;
    73: op1_07_in09 = reg_0473;
    74: op1_07_in09 = reg_0647;
    75: op1_07_in09 = reg_0083;
    76: op1_07_in09 = reg_0059;
    77: op1_07_in09 = reg_0789;
    78: op1_07_in09 = reg_0173;
    79: op1_07_in09 = reg_0208;
    80: op1_07_in09 = reg_0363;
    82: op1_07_in09 = reg_0573;
    83: op1_07_in09 = reg_0751;
    85: op1_07_in09 = reg_0671;
    86: op1_07_in09 = reg_0624;
    87: op1_07_in09 = reg_0427;
    88: op1_07_in09 = reg_0797;
    89: op1_07_in09 = reg_0204;
    90: op1_07_in09 = reg_0455;
    91: op1_07_in09 = reg_0474;
    92: op1_07_in09 = imem04_in[55:52];
    93: op1_07_in09 = reg_0811;
    94: op1_07_in09 = reg_0496;
    95: op1_07_in09 = reg_0629;
    96: op1_07_in09 = reg_0352;
    default: op1_07_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv09 = 1;
    13: op1_07_inv09 = 1;
    14: op1_07_inv09 = 1;
    17: op1_07_inv09 = 1;
    20: op1_07_inv09 = 1;
    22: op1_07_inv09 = 1;
    23: op1_07_inv09 = 1;
    24: op1_07_inv09 = 1;
    25: op1_07_inv09 = 1;
    26: op1_07_inv09 = 1;
    27: op1_07_inv09 = 1;
    30: op1_07_inv09 = 1;
    31: op1_07_inv09 = 1;
    34: op1_07_inv09 = 1;
    35: op1_07_inv09 = 1;
    36: op1_07_inv09 = 1;
    38: op1_07_inv09 = 1;
    40: op1_07_inv09 = 1;
    43: op1_07_inv09 = 1;
    44: op1_07_inv09 = 1;
    45: op1_07_inv09 = 1;
    46: op1_07_inv09 = 1;
    47: op1_07_inv09 = 1;
    48: op1_07_inv09 = 1;
    49: op1_07_inv09 = 1;
    50: op1_07_inv09 = 1;
    51: op1_07_inv09 = 1;
    52: op1_07_inv09 = 1;
    54: op1_07_inv09 = 1;
    57: op1_07_inv09 = 1;
    58: op1_07_inv09 = 1;
    63: op1_07_inv09 = 1;
    64: op1_07_inv09 = 1;
    66: op1_07_inv09 = 1;
    68: op1_07_inv09 = 1;
    69: op1_07_inv09 = 1;
    72: op1_07_inv09 = 1;
    77: op1_07_inv09 = 1;
    78: op1_07_inv09 = 1;
    79: op1_07_inv09 = 1;
    81: op1_07_inv09 = 1;
    82: op1_07_inv09 = 1;
    84: op1_07_inv09 = 1;
    89: op1_07_inv09 = 1;
    91: op1_07_inv09 = 1;
    92: op1_07_inv09 = 1;
    93: op1_07_inv09 = 1;
    95: op1_07_inv09 = 1;
    default: op1_07_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in10 = imem04_in[99:96];
    5: op1_07_in10 = reg_0649;
    42: op1_07_in10 = reg_0649;
    6: op1_07_in10 = imem06_in[67:64];
    7: op1_07_in10 = reg_0691;
    66: op1_07_in10 = reg_0691;
    8: op1_07_in10 = reg_0311;
    9: op1_07_in10 = imem02_in[67:64];
    10: op1_07_in10 = reg_0541;
    19: op1_07_in10 = reg_0541;
    11: op1_07_in10 = reg_0219;
    12: op1_07_in10 = imem07_in[7:4];
    13: op1_07_in10 = reg_0480;
    69: op1_07_in10 = reg_0480;
    14: op1_07_in10 = reg_0110;
    15: op1_07_in10 = reg_0498;
    16: op1_07_in10 = reg_0601;
    17: op1_07_in10 = imem04_in[31:28];
    18: op1_07_in10 = reg_0425;
    20: op1_07_in10 = reg_0448;
    21: op1_07_in10 = imem04_in[87:84];
    22: op1_07_in10 = reg_0807;
    23: op1_07_in10 = reg_0097;
    24: op1_07_in10 = imem05_in[23:20];
    25: op1_07_in10 = reg_0478;
    26: op1_07_in10 = reg_0783;
    27: op1_07_in10 = reg_0031;
    28: op1_07_in10 = imem04_in[103:100];
    29: op1_07_in10 = reg_0492;
    30: op1_07_in10 = reg_0704;
    31: op1_07_in10 = reg_0658;
    32: op1_07_in10 = imem03_in[59:56];
    33: op1_07_in10 = reg_0304;
    34: op1_07_in10 = reg_0515;
    35: op1_07_in10 = reg_0466;
    36: op1_07_in10 = imem02_in[111:108];
    37: op1_07_in10 = reg_0502;
    38: op1_07_in10 = reg_0315;
    39: op1_07_in10 = reg_0152;
    40: op1_07_in10 = imem05_in[115:112];
    41: op1_07_in10 = reg_0472;
    84: op1_07_in10 = reg_0472;
    43: op1_07_in10 = reg_0058;
    44: op1_07_in10 = reg_0727;
    45: op1_07_in10 = reg_0685;
    46: op1_07_in10 = reg_0802;
    47: op1_07_in10 = imem07_in[43:40];
    48: op1_07_in10 = reg_0470;
    64: op1_07_in10 = reg_0470;
    49: op1_07_in10 = reg_0084;
    50: op1_07_in10 = reg_0605;
    51: op1_07_in10 = reg_0055;
    52: op1_07_in10 = reg_0142;
    53: op1_07_in10 = reg_0819;
    54: op1_07_in10 = reg_0160;
    56: op1_07_in10 = reg_0474;
    57: op1_07_in10 = reg_0220;
    58: op1_07_in10 = reg_0203;
    59: op1_07_in10 = reg_0526;
    60: op1_07_in10 = imem02_in[99:96];
    61: op1_07_in10 = imem04_in[7:4];
    62: op1_07_in10 = reg_0169;
    63: op1_07_in10 = reg_0181;
    65: op1_07_in10 = reg_0464;
    67: op1_07_in10 = imem03_in[103:100];
    68: op1_07_in10 = reg_0136;
    70: op1_07_in10 = reg_0671;
    72: op1_07_in10 = reg_0201;
    73: op1_07_in10 = reg_0467;
    74: op1_07_in10 = reg_0138;
    75: op1_07_in10 = reg_0079;
    76: op1_07_in10 = reg_0316;
    77: op1_07_in10 = reg_0785;
    79: op1_07_in10 = reg_0194;
    80: op1_07_in10 = reg_0324;
    81: op1_07_in10 = reg_0475;
    82: op1_07_in10 = reg_0322;
    83: op1_07_in10 = reg_0384;
    85: op1_07_in10 = reg_0127;
    86: op1_07_in10 = reg_0815;
    88: op1_07_in10 = reg_0252;
    89: op1_07_in10 = reg_0198;
    90: op1_07_in10 = reg_0457;
    91: op1_07_in10 = reg_0471;
    92: op1_07_in10 = imem04_in[71:68];
    93: op1_07_in10 = reg_0319;
    94: op1_07_in10 = reg_0637;
    95: op1_07_in10 = reg_0679;
    96: op1_07_in10 = reg_0587;
    default: op1_07_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv10 = 1;
    10: op1_07_inv10 = 1;
    13: op1_07_inv10 = 1;
    14: op1_07_inv10 = 1;
    15: op1_07_inv10 = 1;
    16: op1_07_inv10 = 1;
    17: op1_07_inv10 = 1;
    19: op1_07_inv10 = 1;
    21: op1_07_inv10 = 1;
    22: op1_07_inv10 = 1;
    23: op1_07_inv10 = 1;
    24: op1_07_inv10 = 1;
    26: op1_07_inv10 = 1;
    27: op1_07_inv10 = 1;
    29: op1_07_inv10 = 1;
    30: op1_07_inv10 = 1;
    31: op1_07_inv10 = 1;
    34: op1_07_inv10 = 1;
    37: op1_07_inv10 = 1;
    40: op1_07_inv10 = 1;
    41: op1_07_inv10 = 1;
    42: op1_07_inv10 = 1;
    46: op1_07_inv10 = 1;
    47: op1_07_inv10 = 1;
    48: op1_07_inv10 = 1;
    49: op1_07_inv10 = 1;
    50: op1_07_inv10 = 1;
    56: op1_07_inv10 = 1;
    57: op1_07_inv10 = 1;
    62: op1_07_inv10 = 1;
    63: op1_07_inv10 = 1;
    64: op1_07_inv10 = 1;
    65: op1_07_inv10 = 1;
    66: op1_07_inv10 = 1;
    68: op1_07_inv10 = 1;
    76: op1_07_inv10 = 1;
    77: op1_07_inv10 = 1;
    79: op1_07_inv10 = 1;
    81: op1_07_inv10 = 1;
    84: op1_07_inv10 = 1;
    85: op1_07_inv10 = 1;
    86: op1_07_inv10 = 1;
    89: op1_07_inv10 = 1;
    90: op1_07_inv10 = 1;
    93: op1_07_inv10 = 1;
    96: op1_07_inv10 = 1;
    default: op1_07_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in11 = imem04_in[103:100];
    92: op1_07_in11 = imem04_in[103:100];
    5: op1_07_in11 = reg_0643;
    6: op1_07_in11 = imem06_in[75:72];
    7: op1_07_in11 = reg_0450;
    8: op1_07_in11 = reg_0385;
    9: op1_07_in11 = imem02_in[111:108];
    10: op1_07_in11 = reg_0301;
    11: op1_07_in11 = reg_0123;
    12: op1_07_in11 = imem07_in[27:24];
    13: op1_07_in11 = reg_0467;
    14: op1_07_in11 = imem02_in[31:28];
    15: op1_07_in11 = reg_0259;
    16: op1_07_in11 = reg_0379;
    17: op1_07_in11 = imem04_in[43:40];
    18: op1_07_in11 = reg_0429;
    19: op1_07_in11 = reg_0529;
    20: op1_07_in11 = reg_0166;
    21: op1_07_in11 = imem04_in[91:88];
    22: op1_07_in11 = imem04_in[51:48];
    23: op1_07_in11 = reg_0531;
    24: op1_07_in11 = reg_0484;
    25: op1_07_in11 = reg_0204;
    26: op1_07_in11 = reg_0787;
    27: op1_07_in11 = reg_0753;
    28: op1_07_in11 = reg_0316;
    29: op1_07_in11 = reg_0225;
    30: op1_07_in11 = reg_0714;
    31: op1_07_in11 = reg_0666;
    32: op1_07_in11 = imem03_in[103:100];
    33: op1_07_in11 = reg_0285;
    34: op1_07_in11 = reg_0550;
    35: op1_07_in11 = reg_0480;
    36: op1_07_in11 = imem02_in[115:112];
    37: op1_07_in11 = reg_0244;
    38: op1_07_in11 = reg_0043;
    39: op1_07_in11 = reg_0146;
    52: op1_07_in11 = reg_0146;
    40: op1_07_in11 = reg_0796;
    41: op1_07_in11 = reg_0459;
    48: op1_07_in11 = reg_0459;
    42: op1_07_in11 = reg_0662;
    43: op1_07_in11 = reg_0303;
    44: op1_07_in11 = reg_0253;
    45: op1_07_in11 = reg_0672;
    46: op1_07_in11 = reg_0799;
    47: op1_07_in11 = imem07_in[51:48];
    49: op1_07_in11 = reg_0161;
    63: op1_07_in11 = reg_0161;
    50: op1_07_in11 = reg_0025;
    51: op1_07_in11 = reg_0558;
    53: op1_07_in11 = reg_0338;
    54: op1_07_in11 = reg_0185;
    56: op1_07_in11 = reg_0479;
    84: op1_07_in11 = reg_0479;
    57: op1_07_in11 = reg_0290;
    58: op1_07_in11 = reg_0207;
    59: op1_07_in11 = imem03_in[31:28];
    60: op1_07_in11 = reg_0639;
    61: op1_07_in11 = imem04_in[39:36];
    62: op1_07_in11 = reg_0163;
    64: op1_07_in11 = reg_0474;
    65: op1_07_in11 = reg_0462;
    66: op1_07_in11 = reg_0117;
    67: op1_07_in11 = imem03_in[107:104];
    68: op1_07_in11 = reg_0140;
    69: op1_07_in11 = reg_0208;
    70: op1_07_in11 = reg_0676;
    72: op1_07_in11 = imem01_in[27:24];
    73: op1_07_in11 = reg_0470;
    74: op1_07_in11 = reg_0485;
    75: op1_07_in11 = reg_0280;
    76: op1_07_in11 = reg_0537;
    77: op1_07_in11 = reg_0825;
    79: op1_07_in11 = reg_0196;
    80: op1_07_in11 = reg_0406;
    81: op1_07_in11 = reg_0481;
    82: op1_07_in11 = reg_0777;
    83: op1_07_in11 = reg_0568;
    85: op1_07_in11 = reg_0121;
    86: op1_07_in11 = reg_0817;
    88: op1_07_in11 = reg_0580;
    89: op1_07_in11 = reg_0190;
    90: op1_07_in11 = reg_0461;
    91: op1_07_in11 = reg_0203;
    93: op1_07_in11 = reg_0278;
    94: op1_07_in11 = reg_0747;
    95: op1_07_in11 = reg_0687;
    96: op1_07_in11 = reg_0358;
    default: op1_07_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv11 = 1;
    8: op1_07_inv11 = 1;
    9: op1_07_inv11 = 1;
    12: op1_07_inv11 = 1;
    13: op1_07_inv11 = 1;
    16: op1_07_inv11 = 1;
    17: op1_07_inv11 = 1;
    18: op1_07_inv11 = 1;
    19: op1_07_inv11 = 1;
    21: op1_07_inv11 = 1;
    23: op1_07_inv11 = 1;
    25: op1_07_inv11 = 1;
    26: op1_07_inv11 = 1;
    28: op1_07_inv11 = 1;
    29: op1_07_inv11 = 1;
    30: op1_07_inv11 = 1;
    31: op1_07_inv11 = 1;
    34: op1_07_inv11 = 1;
    35: op1_07_inv11 = 1;
    37: op1_07_inv11 = 1;
    43: op1_07_inv11 = 1;
    45: op1_07_inv11 = 1;
    46: op1_07_inv11 = 1;
    47: op1_07_inv11 = 1;
    49: op1_07_inv11 = 1;
    57: op1_07_inv11 = 1;
    58: op1_07_inv11 = 1;
    59: op1_07_inv11 = 1;
    60: op1_07_inv11 = 1;
    62: op1_07_inv11 = 1;
    63: op1_07_inv11 = 1;
    66: op1_07_inv11 = 1;
    70: op1_07_inv11 = 1;
    74: op1_07_inv11 = 1;
    79: op1_07_inv11 = 1;
    80: op1_07_inv11 = 1;
    89: op1_07_inv11 = 1;
    92: op1_07_inv11 = 1;
    93: op1_07_inv11 = 1;
    95: op1_07_inv11 = 1;
    96: op1_07_inv11 = 1;
    default: op1_07_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in12 = imem04_in[127:124];
    21: op1_07_in12 = imem04_in[127:124];
    5: op1_07_in12 = reg_0357;
    6: op1_07_in12 = imem06_in[79:76];
    7: op1_07_in12 = reg_0461;
    8: op1_07_in12 = reg_0393;
    9: op1_07_in12 = imem02_in[119:116];
    36: op1_07_in12 = imem02_in[119:116];
    10: op1_07_in12 = reg_0285;
    11: op1_07_in12 = reg_0103;
    12: op1_07_in12 = imem07_in[51:48];
    13: op1_07_in12 = reg_0479;
    14: op1_07_in12 = imem02_in[47:44];
    15: op1_07_in12 = reg_0270;
    16: op1_07_in12 = reg_0375;
    17: op1_07_in12 = imem04_in[51:48];
    61: op1_07_in12 = imem04_in[51:48];
    18: op1_07_in12 = reg_0433;
    19: op1_07_in12 = reg_0258;
    20: op1_07_in12 = reg_0171;
    22: op1_07_in12 = imem04_in[99:96];
    23: op1_07_in12 = reg_0498;
    24: op1_07_in12 = reg_0492;
    25: op1_07_in12 = reg_0196;
    58: op1_07_in12 = reg_0196;
    69: op1_07_in12 = reg_0196;
    26: op1_07_in12 = reg_0486;
    27: op1_07_in12 = reg_0035;
    28: op1_07_in12 = reg_0328;
    29: op1_07_in12 = reg_0733;
    30: op1_07_in12 = reg_0712;
    31: op1_07_in12 = reg_0646;
    32: op1_07_in12 = imem03_in[111:108];
    33: op1_07_in12 = reg_0089;
    34: op1_07_in12 = reg_0235;
    35: op1_07_in12 = reg_0208;
    37: op1_07_in12 = reg_0247;
    38: op1_07_in12 = reg_0554;
    39: op1_07_in12 = reg_0140;
    40: op1_07_in12 = reg_0483;
    41: op1_07_in12 = reg_0211;
    42: op1_07_in12 = reg_0665;
    60: op1_07_in12 = reg_0665;
    43: op1_07_in12 = reg_0429;
    44: op1_07_in12 = reg_0061;
    45: op1_07_in12 = reg_0689;
    46: op1_07_in12 = reg_0806;
    47: op1_07_in12 = imem07_in[55:52];
    48: op1_07_in12 = reg_0452;
    84: op1_07_in12 = reg_0452;
    49: op1_07_in12 = reg_0162;
    50: op1_07_in12 = reg_0405;
    51: op1_07_in12 = reg_0305;
    52: op1_07_in12 = imem06_in[11:8];
    53: op1_07_in12 = reg_0368;
    54: op1_07_in12 = reg_0168;
    56: op1_07_in12 = reg_0459;
    57: op1_07_in12 = reg_0425;
    59: op1_07_in12 = imem03_in[43:40];
    62: op1_07_in12 = reg_0166;
    63: op1_07_in12 = reg_0166;
    64: op1_07_in12 = reg_0186;
    65: op1_07_in12 = reg_0480;
    90: op1_07_in12 = reg_0480;
    66: op1_07_in12 = reg_0210;
    67: op1_07_in12 = reg_0317;
    68: op1_07_in12 = imem06_in[27:24];
    70: op1_07_in12 = reg_0674;
    72: op1_07_in12 = imem01_in[51:48];
    73: op1_07_in12 = reg_0474;
    74: op1_07_in12 = reg_0359;
    75: op1_07_in12 = reg_0052;
    76: op1_07_in12 = reg_0057;
    77: op1_07_in12 = reg_0765;
    79: op1_07_in12 = reg_0205;
    80: op1_07_in12 = reg_0566;
    81: op1_07_in12 = reg_0473;
    82: op1_07_in12 = reg_0652;
    83: op1_07_in12 = reg_0570;
    85: op1_07_in12 = imem02_in[63:60];
    86: op1_07_in12 = reg_0370;
    88: op1_07_in12 = reg_0531;
    89: op1_07_in12 = reg_0202;
    91: op1_07_in12 = reg_0193;
    92: op1_07_in12 = imem04_in[107:104];
    93: op1_07_in12 = imem04_in[11:8];
    94: op1_07_in12 = reg_0396;
    95: op1_07_in12 = reg_0780;
    96: op1_07_in12 = reg_0586;
    default: op1_07_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv12 = 1;
    5: op1_07_inv12 = 1;
    6: op1_07_inv12 = 1;
    8: op1_07_inv12 = 1;
    9: op1_07_inv12 = 1;
    10: op1_07_inv12 = 1;
    12: op1_07_inv12 = 1;
    15: op1_07_inv12 = 1;
    16: op1_07_inv12 = 1;
    17: op1_07_inv12 = 1;
    18: op1_07_inv12 = 1;
    20: op1_07_inv12 = 1;
    28: op1_07_inv12 = 1;
    30: op1_07_inv12 = 1;
    32: op1_07_inv12 = 1;
    33: op1_07_inv12 = 1;
    34: op1_07_inv12 = 1;
    35: op1_07_inv12 = 1;
    37: op1_07_inv12 = 1;
    38: op1_07_inv12 = 1;
    40: op1_07_inv12 = 1;
    42: op1_07_inv12 = 1;
    47: op1_07_inv12 = 1;
    49: op1_07_inv12 = 1;
    51: op1_07_inv12 = 1;
    52: op1_07_inv12 = 1;
    53: op1_07_inv12 = 1;
    56: op1_07_inv12 = 1;
    57: op1_07_inv12 = 1;
    59: op1_07_inv12 = 1;
    60: op1_07_inv12 = 1;
    61: op1_07_inv12 = 1;
    62: op1_07_inv12 = 1;
    65: op1_07_inv12 = 1;
    68: op1_07_inv12 = 1;
    72: op1_07_inv12 = 1;
    73: op1_07_inv12 = 1;
    75: op1_07_inv12 = 1;
    76: op1_07_inv12 = 1;
    77: op1_07_inv12 = 1;
    81: op1_07_inv12 = 1;
    82: op1_07_inv12 = 1;
    88: op1_07_inv12 = 1;
    91: op1_07_inv12 = 1;
    92: op1_07_inv12 = 1;
    93: op1_07_inv12 = 1;
    94: op1_07_inv12 = 1;
    default: op1_07_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in13 = reg_0548;
    5: op1_07_in13 = reg_0358;
    6: op1_07_in13 = imem06_in[111:108];
    7: op1_07_in13 = reg_0477;
    8: op1_07_in13 = reg_0001;
    9: op1_07_in13 = reg_0642;
    36: op1_07_in13 = reg_0642;
    10: op1_07_in13 = reg_0059;
    11: op1_07_in13 = reg_0116;
    12: op1_07_in13 = imem07_in[63:60];
    13: op1_07_in13 = reg_0208;
    48: op1_07_in13 = reg_0208;
    14: op1_07_in13 = imem02_in[51:48];
    15: op1_07_in13 = reg_0735;
    16: op1_07_in13 = reg_0315;
    17: op1_07_in13 = imem04_in[59:56];
    18: op1_07_in13 = reg_0423;
    19: op1_07_in13 = reg_0079;
    21: op1_07_in13 = reg_0265;
    22: op1_07_in13 = imem04_in[119:116];
    23: op1_07_in13 = reg_0538;
    24: op1_07_in13 = reg_0793;
    25: op1_07_in13 = reg_0205;
    26: op1_07_in13 = reg_0527;
    27: op1_07_in13 = reg_0005;
    28: op1_07_in13 = reg_0542;
    29: op1_07_in13 = reg_0307;
    30: op1_07_in13 = reg_0707;
    31: op1_07_in13 = reg_0639;
    32: op1_07_in13 = imem03_in[127:124];
    33: op1_07_in13 = reg_0151;
    34: op1_07_in13 = reg_0511;
    35: op1_07_in13 = reg_0210;
    37: op1_07_in13 = reg_0504;
    38: op1_07_in13 = reg_0294;
    39: op1_07_in13 = imem06_in[51:48];
    40: op1_07_in13 = reg_0491;
    41: op1_07_in13 = reg_0201;
    42: op1_07_in13 = reg_0652;
    43: op1_07_in13 = reg_0302;
    44: op1_07_in13 = reg_0434;
    45: op1_07_in13 = reg_0670;
    46: op1_07_in13 = imem04_in[7:4];
    47: op1_07_in13 = imem07_in[59:56];
    49: op1_07_in13 = reg_0159;
    50: op1_07_in13 = reg_0329;
    51: op1_07_in13 = reg_0052;
    52: op1_07_in13 = imem06_in[23:20];
    53: op1_07_in13 = reg_0037;
    56: op1_07_in13 = reg_0214;
    57: op1_07_in13 = reg_0424;
    58: op1_07_in13 = imem01_in[47:44];
    59: op1_07_in13 = imem03_in[59:56];
    60: op1_07_in13 = reg_0352;
    61: op1_07_in13 = imem04_in[67:64];
    62: op1_07_in13 = reg_0185;
    63: op1_07_in13 = reg_0164;
    64: op1_07_in13 = reg_0213;
    65: op1_07_in13 = reg_0471;
    73: op1_07_in13 = reg_0471;
    66: op1_07_in13 = reg_0203;
    67: op1_07_in13 = reg_0579;
    68: op1_07_in13 = imem06_in[63:60];
    69: op1_07_in13 = reg_0195;
    84: op1_07_in13 = reg_0195;
    70: op1_07_in13 = imem02_in[55:52];
    72: op1_07_in13 = imem01_in[67:64];
    74: op1_07_in13 = reg_0360;
    75: op1_07_in13 = reg_0611;
    76: op1_07_in13 = reg_0536;
    77: op1_07_in13 = reg_0828;
    79: op1_07_in13 = reg_0192;
    80: op1_07_in13 = reg_0081;
    81: op1_07_in13 = reg_0187;
    82: op1_07_in13 = reg_0787;
    83: op1_07_in13 = reg_0000;
    85: op1_07_in13 = imem02_in[71:68];
    86: op1_07_in13 = reg_0409;
    88: op1_07_in13 = reg_0148;
    89: op1_07_in13 = reg_0206;
    90: op1_07_in13 = reg_0470;
    91: op1_07_in13 = reg_0198;
    92: op1_07_in13 = reg_0247;
    93: op1_07_in13 = imem04_in[19:16];
    94: op1_07_in13 = reg_0811;
    95: op1_07_in13 = reg_0774;
    96: op1_07_in13 = reg_0353;
    default: op1_07_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv13 = 1;
    5: op1_07_inv13 = 1;
    6: op1_07_inv13 = 1;
    7: op1_07_inv13 = 1;
    12: op1_07_inv13 = 1;
    13: op1_07_inv13 = 1;
    14: op1_07_inv13 = 1;
    16: op1_07_inv13 = 1;
    17: op1_07_inv13 = 1;
    19: op1_07_inv13 = 1;
    21: op1_07_inv13 = 1;
    23: op1_07_inv13 = 1;
    24: op1_07_inv13 = 1;
    26: op1_07_inv13 = 1;
    27: op1_07_inv13 = 1;
    30: op1_07_inv13 = 1;
    31: op1_07_inv13 = 1;
    33: op1_07_inv13 = 1;
    35: op1_07_inv13 = 1;
    37: op1_07_inv13 = 1;
    39: op1_07_inv13 = 1;
    40: op1_07_inv13 = 1;
    41: op1_07_inv13 = 1;
    42: op1_07_inv13 = 1;
    47: op1_07_inv13 = 1;
    48: op1_07_inv13 = 1;
    49: op1_07_inv13 = 1;
    50: op1_07_inv13 = 1;
    51: op1_07_inv13 = 1;
    58: op1_07_inv13 = 1;
    59: op1_07_inv13 = 1;
    62: op1_07_inv13 = 1;
    63: op1_07_inv13 = 1;
    64: op1_07_inv13 = 1;
    65: op1_07_inv13 = 1;
    66: op1_07_inv13 = 1;
    72: op1_07_inv13 = 1;
    75: op1_07_inv13 = 1;
    77: op1_07_inv13 = 1;
    79: op1_07_inv13 = 1;
    82: op1_07_inv13 = 1;
    83: op1_07_inv13 = 1;
    84: op1_07_inv13 = 1;
    85: op1_07_inv13 = 1;
    88: op1_07_inv13 = 1;
    89: op1_07_inv13 = 1;
    90: op1_07_inv13 = 1;
    91: op1_07_inv13 = 1;
    92: op1_07_inv13 = 1;
    96: op1_07_inv13 = 1;
    default: op1_07_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in14 = reg_0549;
    5: op1_07_in14 = reg_0318;
    6: op1_07_in14 = reg_0625;
    7: op1_07_in14 = reg_0460;
    8: op1_07_in14 = reg_0009;
    9: op1_07_in14 = reg_0637;
    10: op1_07_in14 = reg_0066;
    11: op1_07_in14 = reg_0108;
    12: op1_07_in14 = imem07_in[111:108];
    13: op1_07_in14 = reg_0196;
    41: op1_07_in14 = reg_0196;
    14: op1_07_in14 = imem02_in[67:64];
    15: op1_07_in14 = reg_0527;
    16: op1_07_in14 = reg_0367;
    17: op1_07_in14 = imem04_in[67:64];
    18: op1_07_in14 = reg_0175;
    19: op1_07_in14 = reg_0255;
    21: op1_07_in14 = reg_0051;
    22: op1_07_in14 = reg_0055;
    23: op1_07_in14 = imem03_in[7:4];
    24: op1_07_in14 = reg_0495;
    25: op1_07_in14 = imem01_in[15:12];
    26: op1_07_in14 = reg_0224;
    27: op1_07_in14 = reg_0751;
    28: op1_07_in14 = reg_0057;
    29: op1_07_in14 = reg_0744;
    30: op1_07_in14 = reg_0727;
    31: op1_07_in14 = reg_0651;
    32: op1_07_in14 = reg_0586;
    33: op1_07_in14 = reg_0142;
    34: op1_07_in14 = reg_0217;
    35: op1_07_in14 = reg_0194;
    36: op1_07_in14 = reg_0645;
    37: op1_07_in14 = reg_0245;
    38: op1_07_in14 = reg_0268;
    39: op1_07_in14 = imem06_in[91:88];
    40: op1_07_in14 = reg_0492;
    42: op1_07_in14 = reg_0358;
    43: op1_07_in14 = reg_0258;
    44: op1_07_in14 = reg_0443;
    45: op1_07_in14 = reg_0687;
    46: op1_07_in14 = imem04_in[55:52];
    47: op1_07_in14 = imem07_in[79:76];
    48: op1_07_in14 = reg_0191;
    49: op1_07_in14 = reg_0185;
    50: op1_07_in14 = reg_0319;
    67: op1_07_in14 = reg_0319;
    51: op1_07_in14 = reg_0611;
    52: op1_07_in14 = imem06_in[31:28];
    53: op1_07_in14 = reg_0818;
    56: op1_07_in14 = reg_0189;
    57: op1_07_in14 = reg_0420;
    58: op1_07_in14 = imem01_in[67:64];
    59: op1_07_in14 = imem03_in[63:60];
    60: op1_07_in14 = reg_0344;
    61: op1_07_in14 = imem04_in[71:68];
    62: op1_07_in14 = reg_0157;
    63: op1_07_in14 = reg_0157;
    64: op1_07_in14 = imem01_in[75:72];
    65: op1_07_in14 = reg_0200;
    90: op1_07_in14 = reg_0200;
    66: op1_07_in14 = reg_0207;
    68: op1_07_in14 = imem06_in[67:64];
    69: op1_07_in14 = imem01_in[23:20];
    70: op1_07_in14 = imem02_in[99:96];
    72: op1_07_in14 = imem01_in[91:88];
    73: op1_07_in14 = reg_0468;
    74: op1_07_in14 = reg_0590;
    96: op1_07_in14 = reg_0590;
    75: op1_07_in14 = reg_0508;
    76: op1_07_in14 = reg_0547;
    77: op1_07_in14 = imem06_in[43:40];
    79: op1_07_in14 = reg_0197;
    80: op1_07_in14 = reg_0096;
    81: op1_07_in14 = reg_0192;
    82: op1_07_in14 = reg_0767;
    83: op1_07_in14 = reg_0012;
    84: op1_07_in14 = imem01_in[31:28];
    85: op1_07_in14 = imem02_in[107:104];
    86: op1_07_in14 = reg_0814;
    88: op1_07_in14 = reg_0153;
    89: op1_07_in14 = imem01_in[43:40];
    91: op1_07_in14 = reg_0213;
    92: op1_07_in14 = reg_0553;
    93: op1_07_in14 = imem04_in[27:24];
    94: op1_07_in14 = reg_0607;
    95: op1_07_in14 = reg_0771;
    default: op1_07_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv14 = 1;
    6: op1_07_inv14 = 1;
    8: op1_07_inv14 = 1;
    12: op1_07_inv14 = 1;
    13: op1_07_inv14 = 1;
    14: op1_07_inv14 = 1;
    15: op1_07_inv14 = 1;
    17: op1_07_inv14 = 1;
    22: op1_07_inv14 = 1;
    23: op1_07_inv14 = 1;
    25: op1_07_inv14 = 1;
    27: op1_07_inv14 = 1;
    28: op1_07_inv14 = 1;
    30: op1_07_inv14 = 1;
    32: op1_07_inv14 = 1;
    33: op1_07_inv14 = 1;
    40: op1_07_inv14 = 1;
    41: op1_07_inv14 = 1;
    43: op1_07_inv14 = 1;
    46: op1_07_inv14 = 1;
    47: op1_07_inv14 = 1;
    51: op1_07_inv14 = 1;
    53: op1_07_inv14 = 1;
    56: op1_07_inv14 = 1;
    59: op1_07_inv14 = 1;
    61: op1_07_inv14 = 1;
    63: op1_07_inv14 = 1;
    65: op1_07_inv14 = 1;
    66: op1_07_inv14 = 1;
    67: op1_07_inv14 = 1;
    80: op1_07_inv14 = 1;
    83: op1_07_inv14 = 1;
    85: op1_07_inv14 = 1;
    86: op1_07_inv14 = 1;
    92: op1_07_inv14 = 1;
    93: op1_07_inv14 = 1;
    96: op1_07_inv14 = 1;
    default: op1_07_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in15 = reg_0546;
    5: op1_07_in15 = reg_0330;
    6: op1_07_in15 = reg_0626;
    7: op1_07_in15 = reg_0472;
    8: op1_07_in15 = imem04_in[27:24];
    9: op1_07_in15 = reg_0656;
    10: op1_07_in15 = reg_0076;
    11: op1_07_in15 = reg_0114;
    12: op1_07_in15 = reg_0722;
    13: op1_07_in15 = reg_0205;
    14: op1_07_in15 = imem02_in[71:68];
    15: op1_07_in15 = reg_0260;
    16: op1_07_in15 = reg_0337;
    17: op1_07_in15 = imem04_in[71:68];
    18: op1_07_in15 = reg_0165;
    19: op1_07_in15 = reg_0296;
    21: op1_07_in15 = reg_0078;
    22: op1_07_in15 = reg_0088;
    23: op1_07_in15 = imem03_in[11:8];
    24: op1_07_in15 = reg_0783;
    25: op1_07_in15 = imem01_in[19:16];
    26: op1_07_in15 = reg_0285;
    27: op1_07_in15 = imem07_in[23:20];
    28: op1_07_in15 = reg_0516;
    29: op1_07_in15 = reg_0086;
    30: op1_07_in15 = reg_0430;
    31: op1_07_in15 = reg_0641;
    32: op1_07_in15 = reg_0259;
    33: op1_07_in15 = reg_0138;
    34: op1_07_in15 = reg_0244;
    35: op1_07_in15 = reg_0213;
    36: op1_07_in15 = reg_0664;
    37: op1_07_in15 = reg_0111;
    38: op1_07_in15 = reg_0266;
    39: op1_07_in15 = imem06_in[123:120];
    40: op1_07_in15 = reg_0495;
    41: op1_07_in15 = reg_0212;
    42: op1_07_in15 = reg_0345;
    43: op1_07_in15 = reg_0255;
    44: op1_07_in15 = reg_0438;
    45: op1_07_in15 = reg_0475;
    46: op1_07_in15 = imem04_in[59:56];
    47: op1_07_in15 = imem07_in[83:80];
    48: op1_07_in15 = reg_0210;
    49: op1_07_in15 = reg_0176;
    63: op1_07_in15 = reg_0176;
    50: op1_07_in15 = reg_0406;
    51: op1_07_in15 = reg_0074;
    52: op1_07_in15 = imem06_in[47:44];
    53: op1_07_in15 = reg_0238;
    56: op1_07_in15 = reg_0190;
    91: op1_07_in15 = reg_0190;
    57: op1_07_in15 = reg_0123;
    58: op1_07_in15 = imem01_in[75:72];
    59: op1_07_in15 = imem03_in[75:72];
    60: op1_07_in15 = reg_0581;
    61: op1_07_in15 = imem04_in[95:92];
    64: op1_07_in15 = imem01_in[87:84];
    65: op1_07_in15 = reg_0208;
    66: op1_07_in15 = imem01_in[27:24];
    69: op1_07_in15 = imem01_in[27:24];
    67: op1_07_in15 = reg_0528;
    68: op1_07_in15 = imem06_in[71:68];
    77: op1_07_in15 = imem06_in[71:68];
    70: op1_07_in15 = imem02_in[119:116];
    72: op1_07_in15 = imem01_in[115:112];
    73: op1_07_in15 = reg_0452;
    74: op1_07_in15 = reg_0081;
    75: op1_07_in15 = reg_0050;
    76: op1_07_in15 = reg_0052;
    79: op1_07_in15 = imem01_in[55:52];
    80: op1_07_in15 = imem03_in[7:4];
    81: op1_07_in15 = reg_0197;
    82: op1_07_in15 = reg_0661;
    83: op1_07_in15 = reg_0803;
    84: op1_07_in15 = imem01_in[67:64];
    85: op1_07_in15 = reg_0530;
    86: op1_07_in15 = reg_0298;
    88: op1_07_in15 = reg_0155;
    89: op1_07_in15 = imem01_in[91:88];
    90: op1_07_in15 = reg_0204;
    92: op1_07_in15 = reg_0548;
    93: op1_07_in15 = imem04_in[31:28];
    94: op1_07_in15 = reg_0561;
    95: op1_07_in15 = reg_0640;
    96: op1_07_in15 = reg_0343;
    default: op1_07_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv15 = 1;
    7: op1_07_inv15 = 1;
    10: op1_07_inv15 = 1;
    11: op1_07_inv15 = 1;
    15: op1_07_inv15 = 1;
    17: op1_07_inv15 = 1;
    23: op1_07_inv15 = 1;
    25: op1_07_inv15 = 1;
    26: op1_07_inv15 = 1;
    29: op1_07_inv15 = 1;
    32: op1_07_inv15 = 1;
    36: op1_07_inv15 = 1;
    37: op1_07_inv15 = 1;
    42: op1_07_inv15 = 1;
    44: op1_07_inv15 = 1;
    45: op1_07_inv15 = 1;
    47: op1_07_inv15 = 1;
    48: op1_07_inv15 = 1;
    49: op1_07_inv15 = 1;
    50: op1_07_inv15 = 1;
    53: op1_07_inv15 = 1;
    56: op1_07_inv15 = 1;
    58: op1_07_inv15 = 1;
    63: op1_07_inv15 = 1;
    64: op1_07_inv15 = 1;
    65: op1_07_inv15 = 1;
    66: op1_07_inv15 = 1;
    68: op1_07_inv15 = 1;
    69: op1_07_inv15 = 1;
    70: op1_07_inv15 = 1;
    72: op1_07_inv15 = 1;
    73: op1_07_inv15 = 1;
    79: op1_07_inv15 = 1;
    82: op1_07_inv15 = 1;
    88: op1_07_inv15 = 1;
    89: op1_07_inv15 = 1;
    90: op1_07_inv15 = 1;
    93: op1_07_inv15 = 1;
    94: op1_07_inv15 = 1;
    96: op1_07_inv15 = 1;
    default: op1_07_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in16 = reg_0301;
    5: op1_07_in16 = reg_0310;
    6: op1_07_in16 = reg_0633;
    7: op1_07_in16 = reg_0208;
    8: op1_07_in16 = imem04_in[31:28];
    9: op1_07_in16 = reg_0641;
    10: op1_07_in16 = reg_0048;
    11: op1_07_in16 = reg_0101;
    12: op1_07_in16 = reg_0723;
    13: op1_07_in16 = reg_0195;
    56: op1_07_in16 = reg_0195;
    14: op1_07_in16 = imem02_in[79:76];
    15: op1_07_in16 = reg_0266;
    16: op1_07_in16 = reg_0034;
    17: op1_07_in16 = imem05_in[23:20];
    18: op1_07_in16 = reg_0181;
    19: op1_07_in16 = reg_0064;
    21: op1_07_in16 = reg_0062;
    22: op1_07_in16 = reg_0555;
    23: op1_07_in16 = imem03_in[19:16];
    24: op1_07_in16 = reg_0790;
    25: op1_07_in16 = imem01_in[31:28];
    26: op1_07_in16 = reg_0132;
    27: op1_07_in16 = imem07_in[47:44];
    28: op1_07_in16 = reg_0547;
    29: op1_07_in16 = reg_0145;
    30: op1_07_in16 = reg_0426;
    31: op1_07_in16 = reg_0361;
    32: op1_07_in16 = reg_0583;
    33: op1_07_in16 = reg_0130;
    34: op1_07_in16 = reg_0238;
    35: op1_07_in16 = imem01_in[39:36];
    81: op1_07_in16 = imem01_in[39:36];
    36: op1_07_in16 = reg_0661;
    37: op1_07_in16 = reg_0125;
    38: op1_07_in16 = reg_0050;
    51: op1_07_in16 = reg_0050;
    39: op1_07_in16 = reg_0289;
    40: op1_07_in16 = reg_0486;
    41: op1_07_in16 = reg_0197;
    42: op1_07_in16 = reg_0348;
    43: op1_07_in16 = imem05_in[3:0];
    95: op1_07_in16 = imem05_in[3:0];
    44: op1_07_in16 = reg_0175;
    45: op1_07_in16 = reg_0460;
    46: op1_07_in16 = imem04_in[71:68];
    47: op1_07_in16 = reg_0730;
    48: op1_07_in16 = reg_0204;
    65: op1_07_in16 = reg_0204;
    50: op1_07_in16 = reg_0038;
    52: op1_07_in16 = imem06_in[63:60];
    53: op1_07_in16 = reg_0029;
    57: op1_07_in16 = reg_0124;
    58: op1_07_in16 = reg_0663;
    59: op1_07_in16 = imem03_in[83:80];
    60: op1_07_in16 = reg_0345;
    61: op1_07_in16 = imem04_in[123:120];
    64: op1_07_in16 = imem01_in[95:92];
    66: op1_07_in16 = imem01_in[51:48];
    67: op1_07_in16 = reg_0281;
    68: op1_07_in16 = imem06_in[111:108];
    69: op1_07_in16 = imem01_in[35:32];
    70: op1_07_in16 = reg_0089;
    72: op1_07_in16 = imem01_in[119:116];
    73: op1_07_in16 = reg_0456;
    74: op1_07_in16 = reg_0531;
    75: op1_07_in16 = reg_0223;
    76: op1_07_in16 = reg_0611;
    77: op1_07_in16 = imem06_in[79:76];
    79: op1_07_in16 = imem01_in[99:96];
    80: op1_07_in16 = imem03_in[11:8];
    82: op1_07_in16 = imem07_in[31:28];
    83: op1_07_in16 = reg_0016;
    84: op1_07_in16 = imem01_in[79:76];
    85: op1_07_in16 = reg_0056;
    86: op1_07_in16 = reg_0404;
    88: op1_07_in16 = reg_0607;
    89: op1_07_in16 = reg_0376;
    90: op1_07_in16 = reg_0193;
    91: op1_07_in16 = reg_0199;
    92: op1_07_in16 = reg_0551;
    93: op1_07_in16 = imem04_in[39:36];
    94: op1_07_in16 = reg_0368;
    96: op1_07_in16 = reg_0323;
    default: op1_07_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_07_inv16 = 1;
    7: op1_07_inv16 = 1;
    9: op1_07_inv16 = 1;
    11: op1_07_inv16 = 1;
    13: op1_07_inv16 = 1;
    14: op1_07_inv16 = 1;
    17: op1_07_inv16 = 1;
    18: op1_07_inv16 = 1;
    22: op1_07_inv16 = 1;
    23: op1_07_inv16 = 1;
    24: op1_07_inv16 = 1;
    27: op1_07_inv16 = 1;
    28: op1_07_inv16 = 1;
    29: op1_07_inv16 = 1;
    30: op1_07_inv16 = 1;
    31: op1_07_inv16 = 1;
    34: op1_07_inv16 = 1;
    35: op1_07_inv16 = 1;
    36: op1_07_inv16 = 1;
    46: op1_07_inv16 = 1;
    48: op1_07_inv16 = 1;
    50: op1_07_inv16 = 1;
    51: op1_07_inv16 = 1;
    57: op1_07_inv16 = 1;
    61: op1_07_inv16 = 1;
    67: op1_07_inv16 = 1;
    68: op1_07_inv16 = 1;
    69: op1_07_inv16 = 1;
    70: op1_07_inv16 = 1;
    75: op1_07_inv16 = 1;
    77: op1_07_inv16 = 1;
    79: op1_07_inv16 = 1;
    80: op1_07_inv16 = 1;
    84: op1_07_inv16 = 1;
    86: op1_07_inv16 = 1;
    88: op1_07_inv16 = 1;
    90: op1_07_inv16 = 1;
    default: op1_07_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in17 = reg_0289;
    5: op1_07_in17 = reg_0336;
    6: op1_07_in17 = reg_0615;
    7: op1_07_in17 = reg_0210;
    8: op1_07_in17 = imem04_in[95:92];
    9: op1_07_in17 = reg_0662;
    10: op1_07_in17 = reg_0063;
    11: op1_07_in17 = reg_0126;
    12: op1_07_in17 = reg_0703;
    13: op1_07_in17 = imem01_in[27:24];
    14: op1_07_in17 = imem02_in[91:88];
    15: op1_07_in17 = reg_0228;
    16: op1_07_in17 = reg_0040;
    17: op1_07_in17 = imem05_in[63:60];
    18: op1_07_in17 = reg_0161;
    19: op1_07_in17 = reg_0270;
    21: op1_07_in17 = reg_0253;
    22: op1_07_in17 = reg_0554;
    23: op1_07_in17 = imem03_in[47:44];
    24: op1_07_in17 = reg_0225;
    40: op1_07_in17 = reg_0225;
    25: op1_07_in17 = imem01_in[47:44];
    26: op1_07_in17 = reg_0135;
    27: op1_07_in17 = imem07_in[111:108];
    28: op1_07_in17 = reg_0053;
    29: op1_07_in17 = reg_0151;
    30: op1_07_in17 = reg_0445;
    31: op1_07_in17 = reg_0360;
    32: op1_07_in17 = reg_0039;
    33: op1_07_in17 = reg_0140;
    34: op1_07_in17 = reg_0104;
    35: op1_07_in17 = imem01_in[79:76];
    36: op1_07_in17 = reg_0644;
    37: op1_07_in17 = reg_0112;
    38: op1_07_in17 = reg_0078;
    39: op1_07_in17 = reg_0291;
    41: op1_07_in17 = imem01_in[3:0];
    42: op1_07_in17 = reg_0342;
    43: op1_07_in17 = imem05_in[7:4];
    95: op1_07_in17 = imem05_in[7:4];
    44: op1_07_in17 = reg_0163;
    45: op1_07_in17 = reg_0473;
    46: op1_07_in17 = imem04_in[91:88];
    47: op1_07_in17 = reg_0731;
    48: op1_07_in17 = reg_0188;
    50: op1_07_in17 = reg_0614;
    51: op1_07_in17 = reg_0512;
    52: op1_07_in17 = imem06_in[115:112];
    53: op1_07_in17 = imem07_in[23:20];
    56: op1_07_in17 = imem01_in[11:8];
    57: op1_07_in17 = reg_0120;
    58: op1_07_in17 = reg_0820;
    64: op1_07_in17 = reg_0820;
    59: op1_07_in17 = imem03_in[95:92];
    60: op1_07_in17 = reg_0356;
    61: op1_07_in17 = reg_0542;
    65: op1_07_in17 = reg_0193;
    66: op1_07_in17 = imem01_in[59:56];
    67: op1_07_in17 = reg_0394;
    68: op1_07_in17 = imem06_in[127:124];
    69: op1_07_in17 = imem01_in[55:52];
    70: op1_07_in17 = reg_0739;
    72: op1_07_in17 = reg_0111;
    73: op1_07_in17 = reg_0208;
    74: op1_07_in17 = reg_0498;
    75: op1_07_in17 = reg_0643;
    76: op1_07_in17 = reg_0311;
    77: op1_07_in17 = imem06_in[107:104];
    79: op1_07_in17 = imem01_in[103:100];
    80: op1_07_in17 = imem03_in[27:24];
    81: op1_07_in17 = imem01_in[43:40];
    82: op1_07_in17 = imem07_in[67:64];
    83: op1_07_in17 = imem04_in[43:40];
    84: op1_07_in17 = imem01_in[99:96];
    85: op1_07_in17 = reg_0656;
    86: op1_07_in17 = reg_0618;
    88: op1_07_in17 = reg_0652;
    89: op1_07_in17 = reg_0085;
    90: op1_07_in17 = reg_0211;
    91: op1_07_in17 = imem01_in[67:64];
    92: op1_07_in17 = reg_0510;
    93: op1_07_in17 = imem04_in[67:64];
    94: op1_07_in17 = reg_0306;
    96: op1_07_in17 = reg_0540;
    default: op1_07_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv17 = 1;
    6: op1_07_inv17 = 1;
    7: op1_07_inv17 = 1;
    11: op1_07_inv17 = 1;
    12: op1_07_inv17 = 1;
    13: op1_07_inv17 = 1;
    14: op1_07_inv17 = 1;
    16: op1_07_inv17 = 1;
    18: op1_07_inv17 = 1;
    21: op1_07_inv17 = 1;
    24: op1_07_inv17 = 1;
    25: op1_07_inv17 = 1;
    33: op1_07_inv17 = 1;
    35: op1_07_inv17 = 1;
    36: op1_07_inv17 = 1;
    37: op1_07_inv17 = 1;
    38: op1_07_inv17 = 1;
    42: op1_07_inv17 = 1;
    43: op1_07_inv17 = 1;
    44: op1_07_inv17 = 1;
    45: op1_07_inv17 = 1;
    47: op1_07_inv17 = 1;
    48: op1_07_inv17 = 1;
    53: op1_07_inv17 = 1;
    58: op1_07_inv17 = 1;
    60: op1_07_inv17 = 1;
    65: op1_07_inv17 = 1;
    67: op1_07_inv17 = 1;
    74: op1_07_inv17 = 1;
    76: op1_07_inv17 = 1;
    79: op1_07_inv17 = 1;
    81: op1_07_inv17 = 1;
    83: op1_07_inv17 = 1;
    84: op1_07_inv17 = 1;
    86: op1_07_inv17 = 1;
    89: op1_07_inv17 = 1;
    90: op1_07_inv17 = 1;
    93: op1_07_inv17 = 1;
    95: op1_07_inv17 = 1;
    default: op1_07_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in18 = reg_0290;
    88: op1_07_in18 = reg_0290;
    5: op1_07_in18 = reg_0083;
    6: op1_07_in18 = reg_0348;
    7: op1_07_in18 = reg_0203;
    8: op1_07_in18 = imem04_in[107:104];
    9: op1_07_in18 = reg_0358;
    10: op1_07_in18 = reg_0075;
    11: op1_07_in18 = imem02_in[63:60];
    12: op1_07_in18 = reg_0705;
    13: op1_07_in18 = imem01_in[35:32];
    14: op1_07_in18 = reg_0657;
    15: op1_07_in18 = reg_0134;
    16: op1_07_in18 = reg_0817;
    17: op1_07_in18 = imem05_in[111:108];
    18: op1_07_in18 = reg_0167;
    19: op1_07_in18 = reg_0080;
    21: op1_07_in18 = reg_0299;
    22: op1_07_in18 = reg_0057;
    23: op1_07_in18 = reg_0596;
    24: op1_07_in18 = reg_0736;
    25: op1_07_in18 = imem01_in[91:88];
    26: op1_07_in18 = reg_0136;
    27: op1_07_in18 = imem07_in[127:124];
    28: op1_07_in18 = reg_0301;
    29: op1_07_in18 = reg_0155;
    30: op1_07_in18 = reg_0160;
    31: op1_07_in18 = reg_0353;
    32: op1_07_in18 = reg_0587;
    33: op1_07_in18 = imem06_in[39:36];
    34: op1_07_in18 = reg_0119;
    35: op1_07_in18 = imem01_in[83:80];
    36: op1_07_in18 = reg_0659;
    37: op1_07_in18 = reg_0100;
    38: op1_07_in18 = reg_0255;
    96: op1_07_in18 = reg_0255;
    39: op1_07_in18 = reg_0624;
    40: op1_07_in18 = reg_0309;
    41: op1_07_in18 = imem01_in[15:12];
    42: op1_07_in18 = reg_0343;
    43: op1_07_in18 = imem05_in[27:24];
    44: op1_07_in18 = reg_0184;
    45: op1_07_in18 = reg_0458;
    46: op1_07_in18 = imem04_in[127:124];
    47: op1_07_in18 = reg_0714;
    48: op1_07_in18 = reg_0196;
    65: op1_07_in18 = reg_0196;
    50: op1_07_in18 = reg_0028;
    51: op1_07_in18 = reg_0513;
    76: op1_07_in18 = reg_0513;
    52: op1_07_in18 = imem06_in[123:120];
    53: op1_07_in18 = imem07_in[39:36];
    56: op1_07_in18 = imem01_in[43:40];
    57: op1_07_in18 = reg_0672;
    58: op1_07_in18 = reg_0550;
    59: op1_07_in18 = reg_0559;
    60: op1_07_in18 = reg_0360;
    61: op1_07_in18 = reg_0088;
    64: op1_07_in18 = reg_0761;
    66: op1_07_in18 = imem01_in[111:108];
    84: op1_07_in18 = imem01_in[111:108];
    67: op1_07_in18 = reg_0384;
    68: op1_07_in18 = reg_0346;
    69: op1_07_in18 = imem01_in[95:92];
    70: op1_07_in18 = reg_0427;
    72: op1_07_in18 = reg_0520;
    73: op1_07_in18 = reg_0211;
    74: op1_07_in18 = reg_0538;
    75: op1_07_in18 = reg_0311;
    77: op1_07_in18 = imem06_in[111:108];
    79: op1_07_in18 = imem01_in[107:104];
    80: op1_07_in18 = imem03_in[39:36];
    81: op1_07_in18 = imem01_in[115:112];
    82: op1_07_in18 = imem07_in[71:68];
    83: op1_07_in18 = imem04_in[59:56];
    85: op1_07_in18 = reg_0639;
    86: op1_07_in18 = reg_0265;
    89: op1_07_in18 = reg_0772;
    90: op1_07_in18 = reg_0213;
    91: op1_07_in18 = reg_0085;
    92: op1_07_in18 = reg_0556;
    93: op1_07_in18 = imem04_in[87:84];
    94: op1_07_in18 = reg_0806;
    95: op1_07_in18 = imem05_in[55:52];
    default: op1_07_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_07_inv18 = 1;
    7: op1_07_inv18 = 1;
    9: op1_07_inv18 = 1;
    10: op1_07_inv18 = 1;
    12: op1_07_inv18 = 1;
    16: op1_07_inv18 = 1;
    17: op1_07_inv18 = 1;
    21: op1_07_inv18 = 1;
    23: op1_07_inv18 = 1;
    24: op1_07_inv18 = 1;
    26: op1_07_inv18 = 1;
    32: op1_07_inv18 = 1;
    34: op1_07_inv18 = 1;
    37: op1_07_inv18 = 1;
    39: op1_07_inv18 = 1;
    41: op1_07_inv18 = 1;
    42: op1_07_inv18 = 1;
    43: op1_07_inv18 = 1;
    44: op1_07_inv18 = 1;
    45: op1_07_inv18 = 1;
    46: op1_07_inv18 = 1;
    48: op1_07_inv18 = 1;
    51: op1_07_inv18 = 1;
    52: op1_07_inv18 = 1;
    57: op1_07_inv18 = 1;
    58: op1_07_inv18 = 1;
    60: op1_07_inv18 = 1;
    61: op1_07_inv18 = 1;
    64: op1_07_inv18 = 1;
    65: op1_07_inv18 = 1;
    67: op1_07_inv18 = 1;
    68: op1_07_inv18 = 1;
    74: op1_07_inv18 = 1;
    76: op1_07_inv18 = 1;
    77: op1_07_inv18 = 1;
    80: op1_07_inv18 = 1;
    82: op1_07_inv18 = 1;
    84: op1_07_inv18 = 1;
    86: op1_07_inv18 = 1;
    88: op1_07_inv18 = 1;
    90: op1_07_inv18 = 1;
    92: op1_07_inv18 = 1;
    93: op1_07_inv18 = 1;
    96: op1_07_inv18 = 1;
    default: op1_07_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in19 = reg_0291;
    77: op1_07_in19 = reg_0291;
    5: op1_07_in19 = reg_0092;
    6: op1_07_in19 = reg_0372;
    7: op1_07_in19 = reg_0207;
    8: op1_07_in19 = reg_0552;
    9: op1_07_in19 = reg_0359;
    10: op1_07_in19 = imem05_in[39:36];
    11: op1_07_in19 = imem02_in[75:72];
    12: op1_07_in19 = reg_0424;
    13: op1_07_in19 = imem01_in[47:44];
    14: op1_07_in19 = reg_0639;
    15: op1_07_in19 = imem06_in[15:12];
    16: op1_07_in19 = reg_0748;
    17: op1_07_in19 = imem05_in[115:112];
    18: op1_07_in19 = reg_0159;
    19: op1_07_in19 = reg_0526;
    21: op1_07_in19 = reg_0077;
    22: op1_07_in19 = reg_0551;
    23: op1_07_in19 = reg_0583;
    24: op1_07_in19 = reg_0735;
    25: op1_07_in19 = imem01_in[95:92];
    35: op1_07_in19 = imem01_in[95:92];
    26: op1_07_in19 = reg_0133;
    27: op1_07_in19 = reg_0724;
    28: op1_07_in19 = reg_0280;
    29: op1_07_in19 = imem06_in[35:32];
    30: op1_07_in19 = reg_0183;
    31: op1_07_in19 = reg_0365;
    32: op1_07_in19 = reg_0592;
    33: op1_07_in19 = imem06_in[43:40];
    34: op1_07_in19 = reg_0102;
    72: op1_07_in19 = reg_0102;
    81: op1_07_in19 = reg_0102;
    36: op1_07_in19 = reg_0663;
    37: op1_07_in19 = reg_0106;
    38: op1_07_in19 = reg_0256;
    39: op1_07_in19 = reg_0416;
    40: op1_07_in19 = reg_0272;
    41: op1_07_in19 = imem01_in[43:40];
    42: op1_07_in19 = reg_0347;
    43: op1_07_in19 = imem05_in[31:28];
    45: op1_07_in19 = reg_0187;
    46: op1_07_in19 = reg_0553;
    47: op1_07_in19 = reg_0713;
    48: op1_07_in19 = reg_0205;
    65: op1_07_in19 = reg_0205;
    50: op1_07_in19 = reg_0368;
    51: op1_07_in19 = reg_0644;
    52: op1_07_in19 = reg_0289;
    53: op1_07_in19 = imem07_in[59:56];
    56: op1_07_in19 = imem01_in[63:60];
    57: op1_07_in19 = reg_0108;
    58: op1_07_in19 = reg_0760;
    59: op1_07_in19 = reg_0281;
    60: op1_07_in19 = reg_0342;
    61: op1_07_in19 = reg_0055;
    64: op1_07_in19 = reg_0765;
    66: op1_07_in19 = reg_0322;
    67: op1_07_in19 = reg_0568;
    68: op1_07_in19 = reg_0115;
    69: op1_07_in19 = reg_0741;
    84: op1_07_in19 = reg_0741;
    70: op1_07_in19 = reg_0320;
    73: op1_07_in19 = reg_0212;
    74: op1_07_in19 = imem03_in[115:112];
    75: op1_07_in19 = imem05_in[15:12];
    76: op1_07_in19 = reg_0640;
    79: op1_07_in19 = reg_0645;
    80: op1_07_in19 = imem03_in[87:84];
    82: op1_07_in19 = reg_0716;
    83: op1_07_in19 = imem04_in[71:68];
    85: op1_07_in19 = reg_0351;
    86: op1_07_in19 = reg_0519;
    88: op1_07_in19 = reg_0011;
    89: op1_07_in19 = reg_0385;
    90: op1_07_in19 = reg_0199;
    91: op1_07_in19 = reg_0497;
    92: op1_07_in19 = reg_0631;
    93: op1_07_in19 = imem04_in[119:116];
    94: op1_07_in19 = imem04_in[47:44];
    95: op1_07_in19 = reg_0231;
    96: op1_07_in19 = reg_0756;
    default: op1_07_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_07_inv19 = 1;
    8: op1_07_inv19 = 1;
    9: op1_07_inv19 = 1;
    12: op1_07_inv19 = 1;
    14: op1_07_inv19 = 1;
    15: op1_07_inv19 = 1;
    16: op1_07_inv19 = 1;
    17: op1_07_inv19 = 1;
    21: op1_07_inv19 = 1;
    23: op1_07_inv19 = 1;
    24: op1_07_inv19 = 1;
    25: op1_07_inv19 = 1;
    26: op1_07_inv19 = 1;
    27: op1_07_inv19 = 1;
    28: op1_07_inv19 = 1;
    30: op1_07_inv19 = 1;
    34: op1_07_inv19 = 1;
    35: op1_07_inv19 = 1;
    37: op1_07_inv19 = 1;
    38: op1_07_inv19 = 1;
    39: op1_07_inv19 = 1;
    43: op1_07_inv19 = 1;
    47: op1_07_inv19 = 1;
    50: op1_07_inv19 = 1;
    51: op1_07_inv19 = 1;
    52: op1_07_inv19 = 1;
    53: op1_07_inv19 = 1;
    56: op1_07_inv19 = 1;
    58: op1_07_inv19 = 1;
    59: op1_07_inv19 = 1;
    60: op1_07_inv19 = 1;
    64: op1_07_inv19 = 1;
    68: op1_07_inv19 = 1;
    70: op1_07_inv19 = 1;
    72: op1_07_inv19 = 1;
    74: op1_07_inv19 = 1;
    75: op1_07_inv19 = 1;
    76: op1_07_inv19 = 1;
    82: op1_07_inv19 = 1;
    83: op1_07_inv19 = 1;
    84: op1_07_inv19 = 1;
    86: op1_07_inv19 = 1;
    90: op1_07_inv19 = 1;
    91: op1_07_inv19 = 1;
    92: op1_07_inv19 = 1;
    93: op1_07_inv19 = 1;
    default: op1_07_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in20 = reg_0292;
    5: op1_07_in20 = reg_0089;
    6: op1_07_in20 = reg_0349;
    68: op1_07_in20 = reg_0349;
    7: op1_07_in20 = reg_0198;
    8: op1_07_in20 = reg_0542;
    9: op1_07_in20 = reg_0330;
    10: op1_07_in20 = imem05_in[51:48];
    11: op1_07_in20 = imem02_in[87:84];
    12: op1_07_in20 = reg_0432;
    13: op1_07_in20 = imem01_in[87:84];
    14: op1_07_in20 = reg_0638;
    15: op1_07_in20 = imem06_in[35:32];
    16: op1_07_in20 = reg_0818;
    17: op1_07_in20 = reg_0792;
    18: op1_07_in20 = reg_0160;
    19: op1_07_in20 = reg_0081;
    21: op1_07_in20 = imem05_in[43:40];
    22: op1_07_in20 = reg_0058;
    23: op1_07_in20 = reg_0387;
    24: op1_07_in20 = reg_0282;
    25: op1_07_in20 = reg_0497;
    26: op1_07_in20 = reg_0151;
    27: op1_07_in20 = reg_0709;
    28: op1_07_in20 = reg_0306;
    29: op1_07_in20 = imem06_in[39:36];
    30: op1_07_in20 = reg_0178;
    31: op1_07_in20 = reg_0092;
    32: op1_07_in20 = reg_0589;
    33: op1_07_in20 = reg_0616;
    34: op1_07_in20 = reg_0127;
    35: op1_07_in20 = imem01_in[99:96];
    36: op1_07_in20 = reg_0354;
    37: op1_07_in20 = reg_0109;
    38: op1_07_in20 = reg_0288;
    39: op1_07_in20 = reg_0218;
    40: op1_07_in20 = reg_0136;
    41: op1_07_in20 = imem01_in[51:48];
    42: op1_07_in20 = reg_0314;
    85: op1_07_in20 = reg_0314;
    43: op1_07_in20 = imem05_in[83:80];
    45: op1_07_in20 = reg_0194;
    46: op1_07_in20 = reg_0555;
    47: op1_07_in20 = reg_0253;
    48: op1_07_in20 = reg_0190;
    50: op1_07_in20 = reg_0037;
    51: op1_07_in20 = imem05_in[15:12];
    52: op1_07_in20 = reg_0604;
    53: op1_07_in20 = imem07_in[67:64];
    56: op1_07_in20 = imem01_in[107:104];
    57: op1_07_in20 = reg_0675;
    58: op1_07_in20 = reg_0225;
    59: op1_07_in20 = reg_0388;
    67: op1_07_in20 = reg_0388;
    60: op1_07_in20 = reg_0406;
    61: op1_07_in20 = reg_0547;
    64: op1_07_in20 = reg_0649;
    65: op1_07_in20 = reg_0199;
    66: op1_07_in20 = reg_0734;
    69: op1_07_in20 = reg_0224;
    70: op1_07_in20 = reg_0581;
    72: op1_07_in20 = reg_0423;
    73: op1_07_in20 = imem01_in[3:0];
    74: op1_07_in20 = imem03_in[123:120];
    75: op1_07_in20 = imem05_in[39:36];
    76: op1_07_in20 = reg_0644;
    77: op1_07_in20 = reg_0624;
    79: op1_07_in20 = reg_0114;
    84: op1_07_in20 = reg_0114;
    80: op1_07_in20 = imem03_in[95:92];
    81: op1_07_in20 = reg_0235;
    82: op1_07_in20 = reg_0167;
    83: op1_07_in20 = imem04_in[87:84];
    86: op1_07_in20 = reg_0578;
    88: op1_07_in20 = reg_0390;
    89: op1_07_in20 = reg_0820;
    90: op1_07_in20 = reg_0192;
    91: op1_07_in20 = reg_0772;
    92: op1_07_in20 = reg_0302;
    93: op1_07_in20 = imem04_in[123:120];
    94: op1_07_in20 = imem04_in[63:60];
    95: op1_07_in20 = reg_0144;
    96: op1_07_in20 = imem03_in[59:56];
    default: op1_07_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv20 = 1;
    6: op1_07_inv20 = 1;
    7: op1_07_inv20 = 1;
    8: op1_07_inv20 = 1;
    10: op1_07_inv20 = 1;
    11: op1_07_inv20 = 1;
    15: op1_07_inv20 = 1;
    19: op1_07_inv20 = 1;
    21: op1_07_inv20 = 1;
    23: op1_07_inv20 = 1;
    29: op1_07_inv20 = 1;
    30: op1_07_inv20 = 1;
    31: op1_07_inv20 = 1;
    32: op1_07_inv20 = 1;
    34: op1_07_inv20 = 1;
    35: op1_07_inv20 = 1;
    36: op1_07_inv20 = 1;
    37: op1_07_inv20 = 1;
    40: op1_07_inv20 = 1;
    43: op1_07_inv20 = 1;
    45: op1_07_inv20 = 1;
    46: op1_07_inv20 = 1;
    47: op1_07_inv20 = 1;
    51: op1_07_inv20 = 1;
    53: op1_07_inv20 = 1;
    56: op1_07_inv20 = 1;
    58: op1_07_inv20 = 1;
    59: op1_07_inv20 = 1;
    64: op1_07_inv20 = 1;
    66: op1_07_inv20 = 1;
    68: op1_07_inv20 = 1;
    69: op1_07_inv20 = 1;
    70: op1_07_inv20 = 1;
    73: op1_07_inv20 = 1;
    79: op1_07_inv20 = 1;
    82: op1_07_inv20 = 1;
    84: op1_07_inv20 = 1;
    89: op1_07_inv20 = 1;
    92: op1_07_inv20 = 1;
    93: op1_07_inv20 = 1;
    default: op1_07_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in21 = reg_0288;
    5: op1_07_in21 = reg_0049;
    6: op1_07_in21 = reg_0404;
    7: op1_07_in21 = reg_0201;
    8: op1_07_in21 = reg_0555;
    9: op1_07_in21 = reg_0339;
    10: op1_07_in21 = imem05_in[63:60];
    11: op1_07_in21 = imem02_in[99:96];
    12: op1_07_in21 = reg_0422;
    13: op1_07_in21 = imem01_in[103:100];
    14: op1_07_in21 = reg_0644;
    15: op1_07_in21 = imem06_in[55:52];
    16: op1_07_in21 = reg_0751;
    17: op1_07_in21 = reg_0796;
    18: op1_07_in21 = reg_0183;
    19: op1_07_in21 = reg_0082;
    21: op1_07_in21 = imem05_in[55:52];
    75: op1_07_in21 = imem05_in[55:52];
    22: op1_07_in21 = reg_0053;
    47: op1_07_in21 = reg_0053;
    23: op1_07_in21 = reg_0007;
    24: op1_07_in21 = reg_0277;
    25: op1_07_in21 = reg_0496;
    26: op1_07_in21 = imem06_in[7:4];
    40: op1_07_in21 = imem06_in[7:4];
    27: op1_07_in21 = reg_0715;
    28: op1_07_in21 = reg_0291;
    29: op1_07_in21 = imem06_in[59:56];
    30: op1_07_in21 = reg_0157;
    31: op1_07_in21 = reg_0541;
    60: op1_07_in21 = reg_0541;
    32: op1_07_in21 = reg_0593;
    33: op1_07_in21 = reg_0631;
    34: op1_07_in21 = reg_0126;
    35: op1_07_in21 = imem01_in[107:104];
    36: op1_07_in21 = reg_0342;
    37: op1_07_in21 = reg_0107;
    38: op1_07_in21 = imem05_in[3:0];
    39: op1_07_in21 = reg_0817;
    41: op1_07_in21 = imem01_in[75:72];
    42: op1_07_in21 = reg_0095;
    43: op1_07_in21 = imem05_in[103:100];
    45: op1_07_in21 = reg_0192;
    46: op1_07_in21 = reg_0060;
    48: op1_07_in21 = reg_0206;
    50: op1_07_in21 = reg_0029;
    51: op1_07_in21 = imem05_in[23:20];
    52: op1_07_in21 = reg_0624;
    53: op1_07_in21 = imem07_in[103:100];
    56: op1_07_in21 = imem01_in[115:112];
    57: op1_07_in21 = reg_0127;
    58: op1_07_in21 = reg_0232;
    59: op1_07_in21 = reg_0383;
    61: op1_07_in21 = reg_0429;
    64: op1_07_in21 = reg_0322;
    65: op1_07_in21 = imem01_in[39:36];
    90: op1_07_in21 = imem01_in[39:36];
    66: op1_07_in21 = reg_0487;
    67: op1_07_in21 = reg_0398;
    68: op1_07_in21 = reg_0814;
    69: op1_07_in21 = reg_0102;
    89: op1_07_in21 = reg_0102;
    70: op1_07_in21 = reg_0356;
    72: op1_07_in21 = reg_0505;
    73: op1_07_in21 = imem01_in[7:4];
    74: op1_07_in21 = reg_0602;
    76: op1_07_in21 = reg_0109;
    77: op1_07_in21 = reg_0609;
    79: op1_07_in21 = reg_0101;
    80: op1_07_in21 = reg_0599;
    81: op1_07_in21 = reg_0306;
    82: op1_07_in21 = reg_0159;
    83: op1_07_in21 = reg_0247;
    84: op1_07_in21 = reg_0131;
    85: op1_07_in21 = reg_0097;
    86: op1_07_in21 = reg_0654;
    88: op1_07_in21 = reg_0625;
    91: op1_07_in21 = reg_0737;
    92: op1_07_in21 = reg_0616;
    93: op1_07_in21 = imem04_in[127:124];
    94: op1_07_in21 = imem04_in[79:76];
    95: op1_07_in21 = reg_0386;
    96: op1_07_in21 = imem03_in[83:80];
    default: op1_07_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv21 = 1;
    6: op1_07_inv21 = 1;
    10: op1_07_inv21 = 1;
    11: op1_07_inv21 = 1;
    12: op1_07_inv21 = 1;
    13: op1_07_inv21 = 1;
    14: op1_07_inv21 = 1;
    17: op1_07_inv21 = 1;
    18: op1_07_inv21 = 1;
    21: op1_07_inv21 = 1;
    22: op1_07_inv21 = 1;
    23: op1_07_inv21 = 1;
    24: op1_07_inv21 = 1;
    25: op1_07_inv21 = 1;
    26: op1_07_inv21 = 1;
    33: op1_07_inv21 = 1;
    34: op1_07_inv21 = 1;
    35: op1_07_inv21 = 1;
    36: op1_07_inv21 = 1;
    37: op1_07_inv21 = 1;
    38: op1_07_inv21 = 1;
    39: op1_07_inv21 = 1;
    40: op1_07_inv21 = 1;
    41: op1_07_inv21 = 1;
    42: op1_07_inv21 = 1;
    43: op1_07_inv21 = 1;
    46: op1_07_inv21 = 1;
    47: op1_07_inv21 = 1;
    48: op1_07_inv21 = 1;
    52: op1_07_inv21 = 1;
    53: op1_07_inv21 = 1;
    60: op1_07_inv21 = 1;
    64: op1_07_inv21 = 1;
    66: op1_07_inv21 = 1;
    68: op1_07_inv21 = 1;
    72: op1_07_inv21 = 1;
    73: op1_07_inv21 = 1;
    76: op1_07_inv21 = 1;
    77: op1_07_inv21 = 1;
    80: op1_07_inv21 = 1;
    81: op1_07_inv21 = 1;
    83: op1_07_inv21 = 1;
    85: op1_07_inv21 = 1;
    86: op1_07_inv21 = 1;
    91: op1_07_inv21 = 1;
    92: op1_07_inv21 = 1;
    93: op1_07_inv21 = 1;
    94: op1_07_inv21 = 1;
    95: op1_07_inv21 = 1;
    default: op1_07_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in22 = reg_0047;
    5: op1_07_in22 = reg_0732;
    6: op1_07_in22 = reg_0380;
    7: op1_07_in22 = reg_0212;
    8: op1_07_in22 = reg_0546;
    9: op1_07_in22 = reg_0353;
    10: op1_07_in22 = imem05_in[83:80];
    11: op1_07_in22 = imem02_in[119:116];
    12: op1_07_in22 = reg_0421;
    13: op1_07_in22 = imem01_in[111:108];
    35: op1_07_in22 = imem01_in[111:108];
    14: op1_07_in22 = reg_0329;
    15: op1_07_in22 = imem06_in[79:76];
    16: op1_07_in22 = imem07_in[23:20];
    17: op1_07_in22 = reg_0482;
    18: op1_07_in22 = reg_0184;
    19: op1_07_in22 = reg_0789;
    21: op1_07_in22 = imem05_in[107:104];
    22: op1_07_in22 = reg_0294;
    23: op1_07_in22 = reg_0805;
    24: op1_07_in22 = reg_0150;
    25: op1_07_in22 = reg_0520;
    26: op1_07_in22 = imem06_in[39:36];
    40: op1_07_in22 = imem06_in[39:36];
    27: op1_07_in22 = reg_0424;
    28: op1_07_in22 = reg_0268;
    29: op1_07_in22 = reg_0624;
    31: op1_07_in22 = reg_0096;
    32: op1_07_in22 = reg_0597;
    33: op1_07_in22 = reg_0633;
    34: op1_07_in22 = imem02_in[3:0];
    36: op1_07_in22 = reg_0322;
    37: op1_07_in22 = imem02_in[15:12];
    38: op1_07_in22 = imem05_in[35:32];
    39: op1_07_in22 = reg_0608;
    41: op1_07_in22 = imem01_in[127:124];
    42: op1_07_in22 = reg_0535;
    43: op1_07_in22 = imem05_in[119:116];
    75: op1_07_in22 = imem05_in[119:116];
    45: op1_07_in22 = imem01_in[87:84];
    46: op1_07_in22 = reg_0558;
    47: op1_07_in22 = reg_0051;
    48: op1_07_in22 = reg_0736;
    50: op1_07_in22 = reg_0236;
    51: op1_07_in22 = imem05_in[47:44];
    52: op1_07_in22 = reg_0613;
    53: op1_07_in22 = imem07_in[123:120];
    56: op1_07_in22 = reg_0646;
    57: op1_07_in22 = reg_0678;
    58: op1_07_in22 = reg_0567;
    59: op1_07_in22 = reg_0373;
    60: op1_07_in22 = reg_0082;
    61: op1_07_in22 = reg_0079;
    64: op1_07_in22 = reg_0100;
    65: op1_07_in22 = imem01_in[59:56];
    66: op1_07_in22 = reg_0574;
    67: op1_07_in22 = reg_0376;
    68: op1_07_in22 = reg_0293;
    69: op1_07_in22 = reg_0235;
    70: op1_07_in22 = reg_0518;
    72: op1_07_in22 = reg_0120;
    73: op1_07_in22 = imem01_in[75:72];
    74: op1_07_in22 = reg_0599;
    96: op1_07_in22 = reg_0599;
    76: op1_07_in22 = imem05_in[39:36];
    77: op1_07_in22 = reg_0238;
    79: op1_07_in22 = reg_0258;
    80: op1_07_in22 = reg_0559;
    81: op1_07_in22 = reg_0217;
    82: op1_07_in22 = reg_0731;
    83: op1_07_in22 = reg_0262;
    84: op1_07_in22 = reg_0225;
    85: op1_07_in22 = reg_0255;
    86: op1_07_in22 = reg_0405;
    88: op1_07_in22 = reg_0291;
    89: op1_07_in22 = reg_0114;
    90: op1_07_in22 = imem01_in[55:52];
    91: op1_07_in22 = reg_0502;
    92: op1_07_in22 = reg_0585;
    93: op1_07_in22 = reg_0553;
    94: op1_07_in22 = imem04_in[83:80];
    95: op1_07_in22 = reg_0326;
    default: op1_07_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_07_inv22 = 1;
    11: op1_07_inv22 = 1;
    12: op1_07_inv22 = 1;
    13: op1_07_inv22 = 1;
    14: op1_07_inv22 = 1;
    15: op1_07_inv22 = 1;
    18: op1_07_inv22 = 1;
    19: op1_07_inv22 = 1;
    21: op1_07_inv22 = 1;
    24: op1_07_inv22 = 1;
    26: op1_07_inv22 = 1;
    28: op1_07_inv22 = 1;
    31: op1_07_inv22 = 1;
    35: op1_07_inv22 = 1;
    36: op1_07_inv22 = 1;
    37: op1_07_inv22 = 1;
    38: op1_07_inv22 = 1;
    39: op1_07_inv22 = 1;
    40: op1_07_inv22 = 1;
    41: op1_07_inv22 = 1;
    43: op1_07_inv22 = 1;
    46: op1_07_inv22 = 1;
    47: op1_07_inv22 = 1;
    52: op1_07_inv22 = 1;
    56: op1_07_inv22 = 1;
    59: op1_07_inv22 = 1;
    60: op1_07_inv22 = 1;
    61: op1_07_inv22 = 1;
    64: op1_07_inv22 = 1;
    65: op1_07_inv22 = 1;
    66: op1_07_inv22 = 1;
    68: op1_07_inv22 = 1;
    69: op1_07_inv22 = 1;
    70: op1_07_inv22 = 1;
    74: op1_07_inv22 = 1;
    77: op1_07_inv22 = 1;
    80: op1_07_inv22 = 1;
    84: op1_07_inv22 = 1;
    85: op1_07_inv22 = 1;
    86: op1_07_inv22 = 1;
    88: op1_07_inv22 = 1;
    90: op1_07_inv22 = 1;
    92: op1_07_inv22 = 1;
    95: op1_07_inv22 = 1;
    96: op1_07_inv22 = 1;
    default: op1_07_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in23 = reg_0065;
    5: op1_07_in23 = reg_0745;
    6: op1_07_in23 = reg_0368;
    7: op1_07_in23 = reg_0205;
    8: op1_07_in23 = reg_0551;
    46: op1_07_in23 = reg_0551;
    9: op1_07_in23 = reg_0350;
    10: op1_07_in23 = imem05_in[87:84];
    11: op1_07_in23 = imem02_in[123:120];
    12: op1_07_in23 = reg_0426;
    13: op1_07_in23 = reg_0523;
    14: op1_07_in23 = reg_0086;
    15: op1_07_in23 = reg_0614;
    16: op1_07_in23 = imem07_in[55:52];
    17: op1_07_in23 = reg_0484;
    19: op1_07_in23 = reg_0783;
    21: op1_07_in23 = imem05_in[111:108];
    22: op1_07_in23 = reg_0293;
    23: op1_07_in23 = reg_0319;
    24: op1_07_in23 = reg_0152;
    25: op1_07_in23 = reg_0771;
    26: op1_07_in23 = imem06_in[51:48];
    27: op1_07_in23 = reg_0429;
    28: op1_07_in23 = reg_0281;
    29: op1_07_in23 = reg_0617;
    31: op1_07_in23 = reg_0540;
    32: op1_07_in23 = reg_0581;
    33: op1_07_in23 = reg_0369;
    34: op1_07_in23 = imem02_in[11:8];
    35: op1_07_in23 = reg_0758;
    36: op1_07_in23 = reg_0355;
    37: op1_07_in23 = imem02_in[43:40];
    38: op1_07_in23 = imem05_in[47:44];
    39: op1_07_in23 = reg_0618;
    77: op1_07_in23 = reg_0618;
    40: op1_07_in23 = imem06_in[91:88];
    41: op1_07_in23 = reg_0496;
    42: op1_07_in23 = reg_0498;
    43: op1_07_in23 = imem05_in[123:120];
    45: op1_07_in23 = imem01_in[111:108];
    47: op1_07_in23 = reg_0084;
    48: op1_07_in23 = reg_0514;
    50: op1_07_in23 = imem07_in[23:20];
    51: op1_07_in23 = imem05_in[95:92];
    52: op1_07_in23 = reg_0605;
    53: op1_07_in23 = reg_0704;
    56: op1_07_in23 = reg_0733;
    57: op1_07_in23 = imem02_in[27:24];
    58: op1_07_in23 = reg_0244;
    59: op1_07_in23 = reg_0499;
    60: op1_07_in23 = reg_0094;
    61: op1_07_in23 = reg_0631;
    64: op1_07_in23 = reg_0825;
    65: op1_07_in23 = imem01_in[83:80];
    66: op1_07_in23 = reg_0502;
    67: op1_07_in23 = reg_0397;
    68: op1_07_in23 = reg_0377;
    69: op1_07_in23 = reg_0421;
    70: op1_07_in23 = reg_0093;
    72: op1_07_in23 = imem02_in[15:12];
    73: op1_07_in23 = reg_0376;
    74: op1_07_in23 = reg_0591;
    75: op1_07_in23 = reg_0227;
    76: op1_07_in23 = imem05_in[43:40];
    79: op1_07_in23 = reg_0110;
    80: op1_07_in23 = reg_0596;
    81: op1_07_in23 = reg_0294;
    82: op1_07_in23 = reg_0727;
    83: op1_07_in23 = reg_0275;
    84: op1_07_in23 = reg_0423;
    85: op1_07_in23 = reg_0098;
    86: op1_07_in23 = reg_0638;
    88: op1_07_in23 = reg_0814;
    89: op1_07_in23 = reg_0388;
    90: op1_07_in23 = imem01_in[75:72];
    91: op1_07_in23 = reg_0220;
    92: op1_07_in23 = reg_0371;
    93: op1_07_in23 = reg_0548;
    94: op1_07_in23 = imem04_in[111:108];
    95: op1_07_in23 = reg_0552;
    96: op1_07_in23 = reg_0008;
    default: op1_07_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv23 = 1;
    5: op1_07_inv23 = 1;
    7: op1_07_inv23 = 1;
    8: op1_07_inv23 = 1;
    10: op1_07_inv23 = 1;
    12: op1_07_inv23 = 1;
    14: op1_07_inv23 = 1;
    15: op1_07_inv23 = 1;
    16: op1_07_inv23 = 1;
    17: op1_07_inv23 = 1;
    21: op1_07_inv23 = 1;
    22: op1_07_inv23 = 1;
    25: op1_07_inv23 = 1;
    26: op1_07_inv23 = 1;
    27: op1_07_inv23 = 1;
    29: op1_07_inv23 = 1;
    31: op1_07_inv23 = 1;
    37: op1_07_inv23 = 1;
    42: op1_07_inv23 = 1;
    43: op1_07_inv23 = 1;
    46: op1_07_inv23 = 1;
    50: op1_07_inv23 = 1;
    51: op1_07_inv23 = 1;
    52: op1_07_inv23 = 1;
    53: op1_07_inv23 = 1;
    58: op1_07_inv23 = 1;
    59: op1_07_inv23 = 1;
    60: op1_07_inv23 = 1;
    64: op1_07_inv23 = 1;
    66: op1_07_inv23 = 1;
    67: op1_07_inv23 = 1;
    68: op1_07_inv23 = 1;
    70: op1_07_inv23 = 1;
    72: op1_07_inv23 = 1;
    74: op1_07_inv23 = 1;
    75: op1_07_inv23 = 1;
    76: op1_07_inv23 = 1;
    80: op1_07_inv23 = 1;
    82: op1_07_inv23 = 1;
    83: op1_07_inv23 = 1;
    84: op1_07_inv23 = 1;
    88: op1_07_inv23 = 1;
    89: op1_07_inv23 = 1;
    91: op1_07_inv23 = 1;
    92: op1_07_inv23 = 1;
    95: op1_07_inv23 = 1;
    96: op1_07_inv23 = 1;
    default: op1_07_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in24 = reg_0066;
    5: op1_07_in24 = reg_0746;
    6: op1_07_in24 = reg_0027;
    7: op1_07_in24 = reg_0206;
    8: op1_07_in24 = reg_0277;
    9: op1_07_in24 = reg_0095;
    10: op1_07_in24 = imem05_in[103:100];
    11: op1_07_in24 = reg_0646;
    12: op1_07_in24 = reg_0165;
    13: op1_07_in24 = reg_0497;
    14: op1_07_in24 = reg_0087;
    15: op1_07_in24 = reg_0624;
    16: op1_07_in24 = imem07_in[59:56];
    17: op1_07_in24 = reg_0782;
    19: op1_07_in24 = reg_0787;
    21: op1_07_in24 = imem05_in[115:112];
    22: op1_07_in24 = reg_0062;
    23: op1_07_in24 = reg_0557;
    25: op1_07_in24 = reg_0557;
    41: op1_07_in24 = reg_0557;
    24: op1_07_in24 = reg_0153;
    26: op1_07_in24 = reg_0625;
    27: op1_07_in24 = reg_0419;
    28: op1_07_in24 = reg_0065;
    29: op1_07_in24 = reg_0331;
    31: op1_07_in24 = reg_0082;
    32: op1_07_in24 = reg_0394;
    33: op1_07_in24 = reg_0748;
    34: op1_07_in24 = imem02_in[19:16];
    35: op1_07_in24 = reg_0822;
    36: op1_07_in24 = reg_0321;
    37: op1_07_in24 = imem02_in[55:52];
    38: op1_07_in24 = imem05_in[59:56];
    39: op1_07_in24 = reg_0318;
    40: op1_07_in24 = imem06_in[107:104];
    42: op1_07_in24 = reg_0538;
    43: op1_07_in24 = reg_0792;
    45: op1_07_in24 = reg_0501;
    46: op1_07_in24 = reg_0303;
    47: op1_07_in24 = reg_0448;
    48: op1_07_in24 = reg_0086;
    50: op1_07_in24 = imem07_in[67:64];
    51: op1_07_in24 = imem05_in[111:108];
    52: op1_07_in24 = reg_0339;
    53: op1_07_in24 = reg_0719;
    56: op1_07_in24 = reg_0663;
    57: op1_07_in24 = imem02_in[123:120];
    58: op1_07_in24 = reg_0243;
    59: op1_07_in24 = reg_0397;
    60: op1_07_in24 = imem03_in[31:28];
    61: op1_07_in24 = reg_0508;
    64: op1_07_in24 = reg_0487;
    65: op1_07_in24 = imem01_in[99:96];
    66: op1_07_in24 = reg_0220;
    67: op1_07_in24 = reg_0570;
    68: op1_07_in24 = reg_0816;
    69: op1_07_in24 = reg_0418;
    84: op1_07_in24 = reg_0418;
    70: op1_07_in24 = imem03_in[19:16];
    72: op1_07_in24 = imem02_in[27:24];
    73: op1_07_in24 = reg_0645;
    74: op1_07_in24 = reg_0488;
    75: op1_07_in24 = reg_0641;
    76: op1_07_in24 = imem05_in[79:76];
    77: op1_07_in24 = reg_0405;
    79: op1_07_in24 = reg_0241;
    80: op1_07_in24 = reg_0319;
    81: op1_07_in24 = reg_0504;
    82: op1_07_in24 = reg_0334;
    83: op1_07_in24 = reg_0542;
    85: op1_07_in24 = reg_0093;
    86: op1_07_in24 = reg_0169;
    88: op1_07_in24 = reg_0354;
    89: op1_07_in24 = reg_0225;
    90: op1_07_in24 = imem01_in[91:88];
    91: op1_07_in24 = reg_0425;
    92: op1_07_in24 = reg_0640;
    93: op1_07_in24 = reg_0555;
    94: op1_07_in24 = imem04_in[119:116];
    95: op1_07_in24 = reg_0245;
    96: op1_07_in24 = reg_0799;
    default: op1_07_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv24 = 1;
    8: op1_07_inv24 = 1;
    9: op1_07_inv24 = 1;
    10: op1_07_inv24 = 1;
    11: op1_07_inv24 = 1;
    17: op1_07_inv24 = 1;
    19: op1_07_inv24 = 1;
    21: op1_07_inv24 = 1;
    23: op1_07_inv24 = 1;
    24: op1_07_inv24 = 1;
    26: op1_07_inv24 = 1;
    29: op1_07_inv24 = 1;
    39: op1_07_inv24 = 1;
    41: op1_07_inv24 = 1;
    42: op1_07_inv24 = 1;
    43: op1_07_inv24 = 1;
    48: op1_07_inv24 = 1;
    50: op1_07_inv24 = 1;
    52: op1_07_inv24 = 1;
    58: op1_07_inv24 = 1;
    59: op1_07_inv24 = 1;
    61: op1_07_inv24 = 1;
    64: op1_07_inv24 = 1;
    67: op1_07_inv24 = 1;
    69: op1_07_inv24 = 1;
    70: op1_07_inv24 = 1;
    72: op1_07_inv24 = 1;
    75: op1_07_inv24 = 1;
    80: op1_07_inv24 = 1;
    82: op1_07_inv24 = 1;
    88: op1_07_inv24 = 1;
    93: op1_07_inv24 = 1;
    default: op1_07_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in25 = reg_0067;
    5: op1_07_in25 = reg_0739;
    6: op1_07_in25 = reg_0026;
    7: op1_07_in25 = imem01_in[47:44];
    8: op1_07_in25 = reg_0285;
    9: op1_07_in25 = reg_0090;
    10: op1_07_in25 = imem05_in[111:108];
    11: op1_07_in25 = reg_0651;
    12: op1_07_in25 = reg_0161;
    13: op1_07_in25 = reg_0496;
    14: op1_07_in25 = imem03_in[19:16];
    15: op1_07_in25 = reg_0621;
    16: op1_07_in25 = imem07_in[103:100];
    17: op1_07_in25 = reg_0784;
    19: op1_07_in25 = reg_0489;
    21: op1_07_in25 = reg_0482;
    22: op1_07_in25 = reg_0299;
    23: op1_07_in25 = reg_0550;
    25: op1_07_in25 = reg_0550;
    24: op1_07_in25 = reg_0144;
    26: op1_07_in25 = reg_0624;
    27: op1_07_in25 = reg_0434;
    28: op1_07_in25 = reg_0254;
    29: op1_07_in25 = reg_0370;
    31: op1_07_in25 = reg_0093;
    42: op1_07_in25 = reg_0093;
    32: op1_07_in25 = reg_0573;
    86: op1_07_in25 = reg_0573;
    33: op1_07_in25 = reg_0776;
    34: op1_07_in25 = imem02_in[27:24];
    35: op1_07_in25 = reg_0511;
    69: op1_07_in25 = reg_0511;
    36: op1_07_in25 = reg_0081;
    37: op1_07_in25 = imem02_in[91:88];
    38: op1_07_in25 = imem05_in[75:72];
    39: op1_07_in25 = reg_0319;
    40: op1_07_in25 = reg_0605;
    41: op1_07_in25 = reg_0507;
    43: op1_07_in25 = reg_0483;
    45: op1_07_in25 = reg_0497;
    46: op1_07_in25 = reg_0308;
    47: op1_07_in25 = reg_0268;
    48: op1_07_in25 = imem01_in[63:60];
    50: op1_07_in25 = imem07_in[71:68];
    51: op1_07_in25 = reg_0494;
    52: op1_07_in25 = reg_0293;
    53: op1_07_in25 = reg_0723;
    56: op1_07_in25 = reg_0322;
    57: op1_07_in25 = reg_0664;
    58: op1_07_in25 = reg_0123;
    59: op1_07_in25 = reg_0747;
    60: op1_07_in25 = imem03_in[63:60];
    61: op1_07_in25 = reg_0617;
    64: op1_07_in25 = reg_0652;
    65: op1_07_in25 = imem01_in[103:100];
    66: op1_07_in25 = reg_0243;
    67: op1_07_in25 = reg_0000;
    68: op1_07_in25 = reg_0593;
    70: op1_07_in25 = imem03_in[35:32];
    72: op1_07_in25 = imem02_in[75:72];
    73: op1_07_in25 = reg_0258;
    74: op1_07_in25 = reg_0399;
    75: op1_07_in25 = reg_0027;
    76: op1_07_in25 = imem05_in[87:84];
    77: op1_07_in25 = reg_0375;
    79: op1_07_in25 = reg_0073;
    80: op1_07_in25 = reg_0591;
    81: op1_07_in25 = reg_0660;
    82: op1_07_in25 = reg_0449;
    83: op1_07_in25 = reg_0060;
    84: op1_07_in25 = reg_0306;
    85: op1_07_in25 = imem03_in[3:0];
    88: op1_07_in25 = reg_0618;
    89: op1_07_in25 = reg_0235;
    90: op1_07_in25 = imem01_in[119:116];
    91: op1_07_in25 = reg_0603;
    92: op1_07_in25 = reg_0644;
    93: op1_07_in25 = reg_0516;
    94: op1_07_in25 = reg_0544;
    95: op1_07_in25 = reg_0500;
    96: op1_07_in25 = reg_0589;
    default: op1_07_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_07_inv25 = 1;
    8: op1_07_inv25 = 1;
    10: op1_07_inv25 = 1;
    14: op1_07_inv25 = 1;
    17: op1_07_inv25 = 1;
    22: op1_07_inv25 = 1;
    23: op1_07_inv25 = 1;
    24: op1_07_inv25 = 1;
    25: op1_07_inv25 = 1;
    27: op1_07_inv25 = 1;
    28: op1_07_inv25 = 1;
    29: op1_07_inv25 = 1;
    31: op1_07_inv25 = 1;
    34: op1_07_inv25 = 1;
    36: op1_07_inv25 = 1;
    43: op1_07_inv25 = 1;
    45: op1_07_inv25 = 1;
    47: op1_07_inv25 = 1;
    48: op1_07_inv25 = 1;
    51: op1_07_inv25 = 1;
    52: op1_07_inv25 = 1;
    58: op1_07_inv25 = 1;
    60: op1_07_inv25 = 1;
    64: op1_07_inv25 = 1;
    65: op1_07_inv25 = 1;
    69: op1_07_inv25 = 1;
    70: op1_07_inv25 = 1;
    72: op1_07_inv25 = 1;
    79: op1_07_inv25 = 1;
    80: op1_07_inv25 = 1;
    83: op1_07_inv25 = 1;
    86: op1_07_inv25 = 1;
    88: op1_07_inv25 = 1;
    90: op1_07_inv25 = 1;
    91: op1_07_inv25 = 1;
    92: op1_07_inv25 = 1;
    93: op1_07_inv25 = 1;
    94: op1_07_inv25 = 1;
    95: op1_07_inv25 = 1;
    default: op1_07_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in26 = reg_0068;
    5: op1_07_in26 = reg_0569;
    6: op1_07_in26 = reg_0036;
    7: op1_07_in26 = imem01_in[51:48];
    8: op1_07_in26 = reg_0046;
    9: op1_07_in26 = reg_0093;
    10: op1_07_in26 = imem05_in[123:120];
    11: op1_07_in26 = reg_0652;
    12: op1_07_in26 = reg_0167;
    13: op1_07_in26 = reg_0820;
    14: op1_07_in26 = imem03_in[43:40];
    15: op1_07_in26 = reg_0609;
    16: op1_07_in26 = reg_0722;
    17: op1_07_in26 = reg_0267;
    19: op1_07_in26 = imem05_in[15:12];
    21: op1_07_in26 = reg_0789;
    22: op1_07_in26 = reg_0077;
    23: op1_07_in26 = reg_0270;
    24: op1_07_in26 = imem06_in[35:32];
    25: op1_07_in26 = reg_0760;
    26: op1_07_in26 = reg_0622;
    27: op1_07_in26 = reg_0446;
    28: op1_07_in26 = reg_0074;
    29: op1_07_in26 = reg_0401;
    31: op1_07_in26 = reg_0740;
    32: op1_07_in26 = reg_0398;
    33: op1_07_in26 = reg_0406;
    34: op1_07_in26 = imem02_in[43:40];
    35: op1_07_in26 = reg_0248;
    36: op1_07_in26 = reg_0082;
    37: op1_07_in26 = imem02_in[107:104];
    38: op1_07_in26 = imem05_in[79:76];
    39: op1_07_in26 = reg_0764;
    40: op1_07_in26 = reg_0020;
    41: op1_07_in26 = reg_0232;
    48: op1_07_in26 = reg_0232;
    42: op1_07_in26 = imem03_in[3:0];
    43: op1_07_in26 = reg_0484;
    45: op1_07_in26 = reg_0496;
    46: op1_07_in26 = reg_0302;
    47: op1_07_in26 = reg_0180;
    50: op1_07_in26 = imem07_in[79:76];
    51: op1_07_in26 = reg_0783;
    52: op1_07_in26 = reg_0318;
    53: op1_07_in26 = reg_0726;
    56: op1_07_in26 = reg_0563;
    57: op1_07_in26 = reg_0656;
    58: op1_07_in26 = reg_0073;
    59: op1_07_in26 = reg_0396;
    60: op1_07_in26 = imem03_in[83:80];
    61: op1_07_in26 = reg_0233;
    64: op1_07_in26 = reg_0567;
    65: op1_07_in26 = imem01_in[111:108];
    66: op1_07_in26 = reg_0670;
    79: op1_07_in26 = reg_0670;
    67: op1_07_in26 = reg_0010;
    68: op1_07_in26 = reg_0035;
    69: op1_07_in26 = reg_0425;
    70: op1_07_in26 = imem03_in[39:36];
    72: op1_07_in26 = imem02_in[123:120];
    73: op1_07_in26 = reg_0217;
    84: op1_07_in26 = reg_0217;
    89: op1_07_in26 = reg_0217;
    74: op1_07_in26 = reg_0588;
    75: op1_07_in26 = reg_0134;
    76: op1_07_in26 = reg_0133;
    77: op1_07_in26 = reg_0580;
    95: op1_07_in26 = reg_0580;
    80: op1_07_in26 = reg_0750;
    81: op1_07_in26 = reg_0677;
    82: op1_07_in26 = reg_0268;
    83: op1_07_in26 = reg_0516;
    85: op1_07_in26 = imem03_in[15:12];
    86: op1_07_in26 = reg_0700;
    88: op1_07_in26 = reg_0265;
    90: op1_07_in26 = imem01_in[123:120];
    91: op1_07_in26 = reg_0424;
    92: op1_07_in26 = imem05_in[11:8];
    93: op1_07_in26 = reg_0308;
    94: op1_07_in26 = reg_0058;
    96: op1_07_in26 = reg_0572;
    default: op1_07_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_07_inv26 = 1;
    11: op1_07_inv26 = 1;
    13: op1_07_inv26 = 1;
    14: op1_07_inv26 = 1;
    16: op1_07_inv26 = 1;
    21: op1_07_inv26 = 1;
    23: op1_07_inv26 = 1;
    24: op1_07_inv26 = 1;
    33: op1_07_inv26 = 1;
    34: op1_07_inv26 = 1;
    36: op1_07_inv26 = 1;
    40: op1_07_inv26 = 1;
    42: op1_07_inv26 = 1;
    45: op1_07_inv26 = 1;
    46: op1_07_inv26 = 1;
    47: op1_07_inv26 = 1;
    48: op1_07_inv26 = 1;
    50: op1_07_inv26 = 1;
    51: op1_07_inv26 = 1;
    56: op1_07_inv26 = 1;
    61: op1_07_inv26 = 1;
    64: op1_07_inv26 = 1;
    65: op1_07_inv26 = 1;
    68: op1_07_inv26 = 1;
    70: op1_07_inv26 = 1;
    73: op1_07_inv26 = 1;
    75: op1_07_inv26 = 1;
    76: op1_07_inv26 = 1;
    79: op1_07_inv26 = 1;
    81: op1_07_inv26 = 1;
    85: op1_07_inv26 = 1;
    86: op1_07_inv26 = 1;
    92: op1_07_inv26 = 1;
    93: op1_07_inv26 = 1;
    default: op1_07_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in27 = reg_0063;
    22: op1_07_in27 = reg_0063;
    5: op1_07_in27 = reg_0591;
    6: op1_07_in27 = reg_0030;
    7: op1_07_in27 = imem01_in[91:88];
    8: op1_07_in27 = reg_0054;
    9: op1_07_in27 = imem03_in[55:52];
    10: op1_07_in27 = reg_0791;
    11: op1_07_in27 = reg_0325;
    12: op1_07_in27 = reg_0169;
    13: op1_07_in27 = reg_0500;
    14: op1_07_in27 = imem03_in[51:48];
    15: op1_07_in27 = reg_0619;
    16: op1_07_in27 = reg_0704;
    17: op1_07_in27 = reg_0498;
    19: op1_07_in27 = imem05_in[35:32];
    21: op1_07_in27 = reg_0785;
    43: op1_07_in27 = reg_0785;
    23: op1_07_in27 = reg_0515;
    24: op1_07_in27 = imem06_in[43:40];
    25: op1_07_in27 = reg_0559;
    26: op1_07_in27 = reg_0379;
    27: op1_07_in27 = reg_0438;
    28: op1_07_in27 = reg_0256;
    29: op1_07_in27 = reg_0033;
    31: op1_07_in27 = imem03_in[87:84];
    60: op1_07_in27 = imem03_in[87:84];
    32: op1_07_in27 = reg_0499;
    33: op1_07_in27 = reg_0814;
    34: op1_07_in27 = imem02_in[51:48];
    35: op1_07_in27 = reg_0245;
    51: op1_07_in27 = reg_0245;
    36: op1_07_in27 = reg_0757;
    37: op1_07_in27 = imem02_in[111:108];
    38: op1_07_in27 = imem05_in[111:108];
    39: op1_07_in27 = reg_0242;
    40: op1_07_in27 = reg_0371;
    41: op1_07_in27 = reg_0235;
    42: op1_07_in27 = imem03_in[7:4];
    45: op1_07_in27 = reg_0563;
    46: op1_07_in27 = reg_0431;
    47: op1_07_in27 = reg_0161;
    48: op1_07_in27 = reg_0241;
    50: op1_07_in27 = imem07_in[115:112];
    52: op1_07_in27 = reg_0317;
    53: op1_07_in27 = reg_0724;
    56: op1_07_in27 = reg_0652;
    57: op1_07_in27 = reg_0301;
    58: op1_07_in27 = reg_0118;
    59: op1_07_in27 = reg_0374;
    61: op1_07_in27 = reg_0416;
    64: op1_07_in27 = reg_0244;
    65: op1_07_in27 = reg_0761;
    66: op1_07_in27 = reg_0108;
    67: op1_07_in27 = reg_0809;
    68: op1_07_in27 = reg_0812;
    69: op1_07_in27 = reg_0419;
    70: op1_07_in27 = imem03_in[75:72];
    72: op1_07_in27 = reg_0650;
    73: op1_07_in27 = reg_0502;
    74: op1_07_in27 = reg_0368;
    75: op1_07_in27 = reg_0386;
    76: op1_07_in27 = reg_0227;
    77: op1_07_in27 = reg_0029;
    79: op1_07_in27 = reg_0119;
    80: op1_07_in27 = reg_0350;
    81: op1_07_in27 = imem02_in[19:16];
    82: op1_07_in27 = reg_0185;
    83: op1_07_in27 = reg_0303;
    84: op1_07_in27 = reg_0425;
    85: op1_07_in27 = imem03_in[23:20];
    86: op1_07_in27 = reg_0813;
    88: op1_07_in27 = reg_0519;
    89: op1_07_in27 = reg_0567;
    90: op1_07_in27 = reg_0336;
    91: op1_07_in27 = reg_0219;
    92: op1_07_in27 = imem05_in[63:60];
    93: op1_07_in27 = reg_0508;
    94: op1_07_in27 = reg_0177;
    95: op1_07_in27 = reg_0547;
    96: op1_07_in27 = reg_0646;
    default: op1_07_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv27 = 1;
    7: op1_07_inv27 = 1;
    9: op1_07_inv27 = 1;
    11: op1_07_inv27 = 1;
    12: op1_07_inv27 = 1;
    13: op1_07_inv27 = 1;
    14: op1_07_inv27 = 1;
    16: op1_07_inv27 = 1;
    17: op1_07_inv27 = 1;
    21: op1_07_inv27 = 1;
    22: op1_07_inv27 = 1;
    24: op1_07_inv27 = 1;
    25: op1_07_inv27 = 1;
    27: op1_07_inv27 = 1;
    29: op1_07_inv27 = 1;
    33: op1_07_inv27 = 1;
    34: op1_07_inv27 = 1;
    35: op1_07_inv27 = 1;
    36: op1_07_inv27 = 1;
    39: op1_07_inv27 = 1;
    40: op1_07_inv27 = 1;
    43: op1_07_inv27 = 1;
    52: op1_07_inv27 = 1;
    53: op1_07_inv27 = 1;
    56: op1_07_inv27 = 1;
    59: op1_07_inv27 = 1;
    65: op1_07_inv27 = 1;
    66: op1_07_inv27 = 1;
    67: op1_07_inv27 = 1;
    69: op1_07_inv27 = 1;
    73: op1_07_inv27 = 1;
    74: op1_07_inv27 = 1;
    75: op1_07_inv27 = 1;
    76: op1_07_inv27 = 1;
    77: op1_07_inv27 = 1;
    81: op1_07_inv27 = 1;
    85: op1_07_inv27 = 1;
    88: op1_07_inv27 = 1;
    90: op1_07_inv27 = 1;
    91: op1_07_inv27 = 1;
    92: op1_07_inv27 = 1;
    93: op1_07_inv27 = 1;
    94: op1_07_inv27 = 1;
    default: op1_07_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in28 = reg_0069;
    5: op1_07_in28 = reg_0588;
    6: op1_07_in28 = imem07_in[11:8];
    7: op1_07_in28 = reg_0523;
    8: op1_07_in28 = reg_0078;
    9: op1_07_in28 = imem03_in[75:72];
    10: op1_07_in28 = reg_0495;
    11: op1_07_in28 = reg_0310;
    12: op1_07_in28 = reg_0164;
    13: op1_07_in28 = reg_0519;
    14: op1_07_in28 = imem03_in[67:64];
    15: op1_07_in28 = reg_0615;
    16: op1_07_in28 = reg_0720;
    17: op1_07_in28 = reg_0273;
    19: op1_07_in28 = reg_0130;
    21: op1_07_in28 = reg_0794;
    22: op1_07_in28 = reg_0075;
    23: op1_07_in28 = reg_0264;
    24: op1_07_in28 = imem06_in[47:44];
    25: op1_07_in28 = reg_0241;
    41: op1_07_in28 = reg_0241;
    26: op1_07_in28 = reg_0392;
    27: op1_07_in28 = reg_0174;
    28: op1_07_in28 = reg_0288;
    29: op1_07_in28 = reg_0813;
    68: op1_07_in28 = reg_0813;
    31: op1_07_in28 = imem03_in[95:92];
    85: op1_07_in28 = imem03_in[95:92];
    32: op1_07_in28 = reg_0396;
    33: op1_07_in28 = reg_0031;
    34: op1_07_in28 = imem02_in[63:60];
    35: op1_07_in28 = reg_0219;
    36: op1_07_in28 = imem03_in[79:76];
    37: op1_07_in28 = imem02_in[127:124];
    38: op1_07_in28 = reg_0798;
    39: op1_07_in28 = reg_0620;
    40: op1_07_in28 = reg_0608;
    42: op1_07_in28 = imem03_in[71:68];
    43: op1_07_in28 = reg_0736;
    45: op1_07_in28 = reg_0557;
    46: op1_07_in28 = reg_0066;
    47: op1_07_in28 = reg_0166;
    48: op1_07_in28 = reg_0421;
    50: op1_07_in28 = reg_0722;
    51: op1_07_in28 = reg_0256;
    52: op1_07_in28 = reg_0407;
    53: op1_07_in28 = reg_0718;
    56: op1_07_in28 = reg_0423;
    57: op1_07_in28 = reg_0352;
    58: op1_07_in28 = reg_0671;
    59: op1_07_in28 = reg_0801;
    60: op1_07_in28 = reg_0602;
    70: op1_07_in28 = reg_0602;
    61: op1_07_in28 = imem05_in[19:16];
    64: op1_07_in28 = reg_0234;
    65: op1_07_in28 = reg_0737;
    66: op1_07_in28 = reg_0677;
    67: op1_07_in28 = imem04_in[3:0];
    69: op1_07_in28 = reg_0073;
    72: op1_07_in28 = reg_0534;
    73: op1_07_in28 = reg_0244;
    74: op1_07_in28 = reg_0747;
    75: op1_07_in28 = reg_0040;
    76: op1_07_in28 = reg_0550;
    77: op1_07_in28 = reg_0039;
    79: op1_07_in28 = reg_0107;
    80: op1_07_in28 = reg_0600;
    81: op1_07_in28 = imem02_in[35:32];
    83: op1_07_in28 = reg_0631;
    84: op1_07_in28 = reg_0603;
    86: op1_07_in28 = reg_0777;
    88: op1_07_in28 = reg_0578;
    89: op1_07_in28 = reg_0425;
    90: op1_07_in28 = reg_0085;
    91: op1_07_in28 = reg_0123;
    92: op1_07_in28 = imem05_in[71:68];
    93: op1_07_in28 = reg_0617;
    94: op1_07_in28 = reg_0303;
    95: op1_07_in28 = reg_0560;
    96: op1_07_in28 = reg_0562;
    default: op1_07_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv28 = 1;
    8: op1_07_inv28 = 1;
    13: op1_07_inv28 = 1;
    15: op1_07_inv28 = 1;
    16: op1_07_inv28 = 1;
    22: op1_07_inv28 = 1;
    23: op1_07_inv28 = 1;
    26: op1_07_inv28 = 1;
    27: op1_07_inv28 = 1;
    28: op1_07_inv28 = 1;
    31: op1_07_inv28 = 1;
    32: op1_07_inv28 = 1;
    34: op1_07_inv28 = 1;
    42: op1_07_inv28 = 1;
    43: op1_07_inv28 = 1;
    45: op1_07_inv28 = 1;
    47: op1_07_inv28 = 1;
    50: op1_07_inv28 = 1;
    51: op1_07_inv28 = 1;
    60: op1_07_inv28 = 1;
    61: op1_07_inv28 = 1;
    64: op1_07_inv28 = 1;
    69: op1_07_inv28 = 1;
    73: op1_07_inv28 = 1;
    75: op1_07_inv28 = 1;
    80: op1_07_inv28 = 1;
    84: op1_07_inv28 = 1;
    91: op1_07_inv28 = 1;
    94: op1_07_inv28 = 1;
    95: op1_07_inv28 = 1;
    default: op1_07_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in29 = reg_0070;
    5: op1_07_in29 = reg_0384;
    6: op1_07_in29 = imem07_in[19:16];
    7: op1_07_in29 = reg_0522;
    8: op1_07_in29 = reg_0041;
    9: op1_07_in29 = imem03_in[103:100];
    42: op1_07_in29 = imem03_in[103:100];
    10: op1_07_in29 = reg_0486;
    11: op1_07_in29 = reg_0342;
    12: op1_07_in29 = reg_0185;
    13: op1_07_in29 = reg_0521;
    14: op1_07_in29 = imem03_in[71:68];
    15: op1_07_in29 = reg_0386;
    16: op1_07_in29 = reg_0726;
    17: op1_07_in29 = reg_0270;
    19: op1_07_in29 = reg_0134;
    21: op1_07_in29 = reg_0783;
    22: op1_07_in29 = reg_0256;
    23: op1_07_in29 = reg_0317;
    70: op1_07_in29 = reg_0317;
    24: op1_07_in29 = imem06_in[67:64];
    25: op1_07_in29 = reg_0244;
    26: op1_07_in29 = reg_0404;
    27: op1_07_in29 = reg_0179;
    28: op1_07_in29 = imem05_in[3:0];
    29: op1_07_in29 = reg_0032;
    31: op1_07_in29 = reg_0565;
    32: op1_07_in29 = reg_0000;
    33: op1_07_in29 = reg_0778;
    34: op1_07_in29 = imem02_in[123:120];
    35: op1_07_in29 = reg_0118;
    36: op1_07_in29 = imem03_in[99:96];
    85: op1_07_in29 = imem03_in[99:96];
    37: op1_07_in29 = reg_0658;
    38: op1_07_in29 = reg_0483;
    39: op1_07_in29 = reg_0040;
    40: op1_07_in29 = reg_0618;
    41: op1_07_in29 = reg_0240;
    43: op1_07_in29 = reg_0279;
    45: op1_07_in29 = reg_0761;
    46: op1_07_in29 = reg_0065;
    83: op1_07_in29 = reg_0065;
    48: op1_07_in29 = reg_0306;
    50: op1_07_in29 = reg_0704;
    51: op1_07_in29 = reg_0103;
    52: op1_07_in29 = reg_0607;
    53: op1_07_in29 = reg_0061;
    56: op1_07_in29 = reg_0574;
    57: op1_07_in29 = reg_0361;
    58: op1_07_in29 = reg_0676;
    59: op1_07_in29 = reg_0806;
    60: op1_07_in29 = reg_0591;
    61: op1_07_in29 = imem05_in[31:28];
    64: op1_07_in29 = reg_0506;
    65: op1_07_in29 = reg_0241;
    66: op1_07_in29 = reg_0675;
    69: op1_07_in29 = reg_0675;
    67: op1_07_in29 = imem04_in[111:108];
    68: op1_07_in29 = reg_0642;
    72: op1_07_in29 = reg_0639;
    73: op1_07_in29 = reg_0294;
    74: op1_07_in29 = reg_0396;
    75: op1_07_in29 = reg_0812;
    76: op1_07_in29 = reg_0090;
    77: op1_07_in29 = reg_0664;
    79: op1_07_in29 = imem02_in[75:72];
    80: op1_07_in29 = reg_0648;
    81: op1_07_in29 = imem02_in[51:48];
    84: op1_07_in29 = reg_0105;
    86: op1_07_in29 = reg_0794;
    88: op1_07_in29 = reg_0775;
    89: op1_07_in29 = reg_0419;
    90: op1_07_in29 = reg_0111;
    91: op1_07_in29 = reg_0673;
    92: op1_07_in29 = imem05_in[103:100];
    93: op1_07_in29 = reg_0614;
    94: op1_07_in29 = reg_0079;
    95: op1_07_in29 = reg_0781;
    96: op1_07_in29 = reg_0398;
    default: op1_07_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_07_inv29 = 1;
    7: op1_07_inv29 = 1;
    8: op1_07_inv29 = 1;
    11: op1_07_inv29 = 1;
    13: op1_07_inv29 = 1;
    16: op1_07_inv29 = 1;
    22: op1_07_inv29 = 1;
    24: op1_07_inv29 = 1;
    25: op1_07_inv29 = 1;
    26: op1_07_inv29 = 1;
    27: op1_07_inv29 = 1;
    29: op1_07_inv29 = 1;
    32: op1_07_inv29 = 1;
    33: op1_07_inv29 = 1;
    35: op1_07_inv29 = 1;
    37: op1_07_inv29 = 1;
    40: op1_07_inv29 = 1;
    41: op1_07_inv29 = 1;
    42: op1_07_inv29 = 1;
    45: op1_07_inv29 = 1;
    53: op1_07_inv29 = 1;
    59: op1_07_inv29 = 1;
    60: op1_07_inv29 = 1;
    61: op1_07_inv29 = 1;
    64: op1_07_inv29 = 1;
    65: op1_07_inv29 = 1;
    66: op1_07_inv29 = 1;
    67: op1_07_inv29 = 1;
    68: op1_07_inv29 = 1;
    73: op1_07_inv29 = 1;
    75: op1_07_inv29 = 1;
    79: op1_07_inv29 = 1;
    80: op1_07_inv29 = 1;
    86: op1_07_inv29 = 1;
    88: op1_07_inv29 = 1;
    91: op1_07_inv29 = 1;
    94: op1_07_inv29 = 1;
    default: op1_07_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_07_in30 = imem05_in[23:20];
    5: op1_07_in30 = reg_0387;
    6: op1_07_in30 = imem07_in[27:24];
    7: op1_07_in30 = reg_0511;
    8: op1_07_in30 = reg_0057;
    9: op1_07_in30 = imem03_in[111:108];
    10: op1_07_in30 = reg_0262;
    11: op1_07_in30 = reg_0045;
    12: op1_07_in30 = reg_0171;
    13: op1_07_in30 = reg_0515;
    14: op1_07_in30 = imem03_in[75:72];
    15: op1_07_in30 = reg_0409;
    16: op1_07_in30 = reg_0702;
    17: op1_07_in30 = reg_0269;
    19: op1_07_in30 = imem06_in[15:12];
    21: op1_07_in30 = reg_0486;
    22: op1_07_in30 = imem05_in[15:12];
    23: op1_07_in30 = reg_0311;
    24: op1_07_in30 = imem06_in[71:68];
    25: op1_07_in30 = reg_0238;
    26: op1_07_in30 = reg_0401;
    27: op1_07_in30 = reg_0161;
    28: op1_07_in30 = imem05_in[83:80];
    29: op1_07_in30 = reg_0815;
    31: op1_07_in30 = reg_0597;
    32: op1_07_in30 = reg_0006;
    33: op1_07_in30 = reg_0777;
    34: op1_07_in30 = reg_0666;
    37: op1_07_in30 = reg_0666;
    35: op1_07_in30 = reg_0120;
    36: op1_07_in30 = imem03_in[107:104];
    38: op1_07_in30 = reg_0788;
    39: op1_07_in30 = reg_0621;
    40: op1_07_in30 = reg_0293;
    41: op1_07_in30 = reg_0502;
    56: op1_07_in30 = reg_0502;
    42: op1_07_in30 = imem03_in[115:112];
    43: op1_07_in30 = reg_0742;
    45: op1_07_in30 = reg_0760;
    46: op1_07_in30 = reg_0519;
    48: op1_07_in30 = reg_0234;
    73: op1_07_in30 = reg_0234;
    50: op1_07_in30 = reg_0719;
    51: op1_07_in30 = reg_0150;
    52: op1_07_in30 = reg_0620;
    53: op1_07_in30 = reg_0029;
    57: op1_07_in30 = reg_0363;
    58: op1_07_in30 = reg_0678;
    59: op1_07_in30 = reg_0010;
    60: op1_07_in30 = reg_0528;
    61: op1_07_in30 = imem05_in[71:68];
    64: op1_07_in30 = reg_0506;
    65: op1_07_in30 = reg_0423;
    66: op1_07_in30 = reg_0106;
    67: op1_07_in30 = reg_0316;
    68: op1_07_in30 = reg_0752;
    69: op1_07_in30 = imem02_in[27:24];
    70: op1_07_in30 = reg_0329;
    72: op1_07_in30 = reg_0647;
    74: op1_07_in30 = reg_0570;
    75: op1_07_in30 = reg_0149;
    76: op1_07_in30 = reg_0665;
    77: op1_07_in30 = reg_0256;
    79: op1_07_in30 = imem02_in[91:88];
    80: op1_07_in30 = reg_0321;
    81: op1_07_in30 = imem02_in[67:64];
    83: op1_07_in30 = reg_0643;
    84: op1_07_in30 = reg_0108;
    91: op1_07_in30 = reg_0108;
    85: op1_07_in30 = imem03_in[103:100];
    86: op1_07_in30 = reg_0651;
    88: op1_07_in30 = reg_0246;
    89: op1_07_in30 = reg_0424;
    90: op1_07_in30 = reg_0385;
    92: op1_07_in30 = imem05_in[107:104];
    93: op1_07_in30 = reg_0779;
    94: op1_07_in30 = reg_0052;
    95: op1_07_in30 = reg_0828;
    96: op1_07_in30 = reg_0637;
    default: op1_07_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_07_inv30 = 1;
    8: op1_07_inv30 = 1;
    10: op1_07_inv30 = 1;
    11: op1_07_inv30 = 1;
    16: op1_07_inv30 = 1;
    17: op1_07_inv30 = 1;
    19: op1_07_inv30 = 1;
    24: op1_07_inv30 = 1;
    25: op1_07_inv30 = 1;
    26: op1_07_inv30 = 1;
    27: op1_07_inv30 = 1;
    28: op1_07_inv30 = 1;
    29: op1_07_inv30 = 1;
    31: op1_07_inv30 = 1;
    34: op1_07_inv30 = 1;
    35: op1_07_inv30 = 1;
    36: op1_07_inv30 = 1;
    37: op1_07_inv30 = 1;
    38: op1_07_inv30 = 1;
    40: op1_07_inv30 = 1;
    51: op1_07_inv30 = 1;
    56: op1_07_inv30 = 1;
    59: op1_07_inv30 = 1;
    64: op1_07_inv30 = 1;
    74: op1_07_inv30 = 1;
    76: op1_07_inv30 = 1;
    81: op1_07_inv30 = 1;
    83: op1_07_inv30 = 1;
    84: op1_07_inv30 = 1;
    86: op1_07_inv30 = 1;
    89: op1_07_inv30 = 1;
    90: op1_07_inv30 = 1;
    91: op1_07_inv30 = 1;
    92: op1_07_inv30 = 1;
    default: op1_07_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_07_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_07_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in00 = imem05_in[31:28];
    83: op1_08_in00 = imem05_in[31:28];
    5: op1_08_in00 = reg_0391;
    6: op1_08_in00 = imem07_in[47:44];
    2: op1_08_in00 = imem07_in[47:44];
    7: op1_08_in00 = reg_0503;
    8: op1_08_in00 = imem05_in[39:36];
    9: op1_08_in00 = reg_0586;
    10: op1_08_in00 = reg_0259;
    11: op1_08_in00 = reg_0052;
    12: op1_08_in00 = imem00_in[11:8];
    13: op1_08_in00 = reg_0755;
    14: op1_08_in00 = imem03_in[95:92];
    3: op1_08_in00 = imem07_in[15:12];
    15: op1_08_in00 = reg_0313;
    16: op1_08_in00 = imem00_in[59:56];
    63: op1_08_in00 = imem00_in[59:56];
    17: op1_08_in00 = reg_0732;
    18: op1_08_in00 = imem00_in[91:88];
    19: op1_08_in00 = imem06_in[43:40];
    20: op1_08_in00 = imem00_in[15:12];
    27: op1_08_in00 = imem00_in[15:12];
    82: op1_08_in00 = imem00_in[15:12];
    21: op1_08_in00 = reg_0279;
    22: op1_08_in00 = imem05_in[47:44];
    23: op1_08_in00 = reg_0529;
    24: op1_08_in00 = imem06_in[123:120];
    25: op1_08_in00 = reg_0123;
    26: op1_08_in00 = reg_0028;
    1: op1_08_in00 = imem07_in[95:92];
    28: op1_08_in00 = imem05_in[99:96];
    29: op1_08_in00 = reg_0816;
    30: op1_08_in00 = imem00_in[43:40];
    31: op1_08_in00 = reg_0595;
    32: op1_08_in00 = reg_0802;
    33: op1_08_in00 = reg_0368;
    39: op1_08_in00 = reg_0368;
    34: op1_08_in00 = reg_0647;
    35: op1_08_in00 = reg_0112;
    36: op1_08_in00 = reg_0039;
    37: op1_08_in00 = reg_0664;
    38: op1_08_in00 = reg_0495;
    40: op1_08_in00 = reg_0369;
    41: op1_08_in00 = reg_0244;
    42: op1_08_in00 = reg_0602;
    85: op1_08_in00 = reg_0602;
    43: op1_08_in00 = reg_0277;
    44: op1_08_in00 = imem00_in[71:68];
    55: op1_08_in00 = imem00_in[71:68];
    45: op1_08_in00 = reg_0241;
    46: op1_08_in00 = reg_0229;
    47: op1_08_in00 = imem00_in[31:28];
    78: op1_08_in00 = imem00_in[31:28];
    48: op1_08_in00 = reg_0120;
    49: op1_08_in00 = imem00_in[19:16];
    50: op1_08_in00 = reg_0717;
    51: op1_08_in00 = reg_0138;
    52: op1_08_in00 = reg_0815;
    53: op1_08_in00 = reg_0443;
    54: op1_08_in00 = reg_0113;
    56: op1_08_in00 = reg_0234;
    57: op1_08_in00 = reg_0324;
    58: op1_08_in00 = imem02_in[19:16];
    59: op1_08_in00 = imem04_in[59:56];
    60: op1_08_in00 = reg_0588;
    61: op1_08_in00 = imem05_in[87:84];
    62: op1_08_in00 = imem00_in[55:52];
    64: op1_08_in00 = reg_0419;
    65: op1_08_in00 = reg_0424;
    66: op1_08_in00 = reg_0601;
    67: op1_08_in00 = reg_0328;
    68: op1_08_in00 = imem07_in[11:8];
    69: op1_08_in00 = imem02_in[51:48];
    70: op1_08_in00 = reg_0600;
    71: op1_08_in00 = imem00_in[63:60];
    72: op1_08_in00 = reg_0607;
    73: op1_08_in00 = reg_0243;
    89: op1_08_in00 = reg_0243;
    74: op1_08_in00 = reg_0000;
    75: op1_08_in00 = reg_0827;
    76: op1_08_in00 = reg_0144;
    77: op1_08_in00 = imem07_in[67:64];
    79: op1_08_in00 = imem02_in[99:96];
    80: op1_08_in00 = reg_0575;
    81: op1_08_in00 = imem02_in[115:112];
    84: op1_08_in00 = reg_0127;
    86: op1_08_in00 = reg_0787;
    87: op1_08_in00 = imem00_in[7:4];
    88: op1_08_in00 = imem06_in[3:0];
    90: op1_08_in00 = reg_0102;
    91: op1_08_in00 = reg_0675;
    92: op1_08_in00 = reg_0135;
    93: op1_08_in00 = reg_0301;
    94: op1_08_in00 = reg_0433;
    95: op1_08_in00 = imem06_in[15:12];
    96: op1_08_in00 = reg_0649;
    default: op1_08_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv00 = 1;
    6: op1_08_inv00 = 1;
    9: op1_08_inv00 = 1;
    10: op1_08_inv00 = 1;
    11: op1_08_inv00 = 1;
    12: op1_08_inv00 = 1;
    3: op1_08_inv00 = 1;
    17: op1_08_inv00 = 1;
    19: op1_08_inv00 = 1;
    21: op1_08_inv00 = 1;
    25: op1_08_inv00 = 1;
    26: op1_08_inv00 = 1;
    31: op1_08_inv00 = 1;
    32: op1_08_inv00 = 1;
    38: op1_08_inv00 = 1;
    39: op1_08_inv00 = 1;
    40: op1_08_inv00 = 1;
    42: op1_08_inv00 = 1;
    44: op1_08_inv00 = 1;
    46: op1_08_inv00 = 1;
    47: op1_08_inv00 = 1;
    48: op1_08_inv00 = 1;
    53: op1_08_inv00 = 1;
    54: op1_08_inv00 = 1;
    59: op1_08_inv00 = 1;
    63: op1_08_inv00 = 1;
    69: op1_08_inv00 = 1;
    70: op1_08_inv00 = 1;
    75: op1_08_inv00 = 1;
    76: op1_08_inv00 = 1;
    78: op1_08_inv00 = 1;
    81: op1_08_inv00 = 1;
    82: op1_08_inv00 = 1;
    83: op1_08_inv00 = 1;
    85: op1_08_inv00 = 1;
    86: op1_08_inv00 = 1;
    90: op1_08_inv00 = 1;
    91: op1_08_inv00 = 1;
    93: op1_08_inv00 = 1;
    94: op1_08_inv00 = 1;
    95: op1_08_inv00 = 1;
    96: op1_08_inv00 = 1;
    default: op1_08_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in01 = imem05_in[35:32];
    5: op1_08_in01 = reg_0321;
    6: op1_08_in01 = imem07_in[59:56];
    7: op1_08_in01 = reg_0235;
    8: op1_08_in01 = imem05_in[55:52];
    9: op1_08_in01 = reg_0587;
    10: op1_08_in01 = reg_0260;
    11: op1_08_in01 = reg_0098;
    12: op1_08_in01 = imem00_in[15:12];
    13: op1_08_in01 = reg_0821;
    14: op1_08_in01 = reg_0582;
    3: op1_08_in01 = imem07_in[47:44];
    15: op1_08_in01 = reg_0383;
    16: op1_08_in01 = imem00_in[75:72];
    17: op1_08_in01 = reg_0139;
    18: op1_08_in01 = imem00_in[123:120];
    30: op1_08_in01 = imem00_in[123:120];
    19: op1_08_in01 = imem06_in[63:60];
    20: op1_08_in01 = imem00_in[27:24];
    2: op1_08_in01 = imem07_in[99:96];
    1: op1_08_in01 = imem07_in[99:96];
    21: op1_08_in01 = reg_0275;
    22: op1_08_in01 = imem05_in[67:64];
    23: op1_08_in01 = reg_0302;
    24: op1_08_in01 = reg_0610;
    25: op1_08_in01 = reg_0122;
    73: op1_08_in01 = reg_0122;
    26: op1_08_in01 = reg_0032;
    27: op1_08_in01 = imem00_in[59:56];
    28: op1_08_in01 = reg_0792;
    29: op1_08_in01 = reg_0037;
    52: op1_08_in01 = reg_0037;
    31: op1_08_in01 = reg_0588;
    32: op1_08_in01 = reg_0016;
    33: op1_08_in01 = reg_0380;
    34: op1_08_in01 = reg_0229;
    35: op1_08_in01 = reg_0102;
    48: op1_08_in01 = reg_0102;
    36: op1_08_in01 = reg_0387;
    37: op1_08_in01 = reg_0657;
    38: op1_08_in01 = reg_0790;
    39: op1_08_in01 = reg_0238;
    40: op1_08_in01 = reg_0577;
    41: op1_08_in01 = reg_0216;
    42: op1_08_in01 = reg_0586;
    43: op1_08_in01 = reg_0132;
    44: op1_08_in01 = reg_0682;
    45: op1_08_in01 = reg_0240;
    46: op1_08_in01 = reg_0256;
    47: op1_08_in01 = imem00_in[55:52];
    49: op1_08_in01 = imem00_in[55:52];
    50: op1_08_in01 = reg_0705;
    51: op1_08_in01 = reg_0129;
    53: op1_08_in01 = reg_0267;
    54: op1_08_in01 = reg_0112;
    55: op1_08_in01 = imem00_in[127:124];
    56: op1_08_in01 = reg_0123;
    57: op1_08_in01 = reg_0092;
    58: op1_08_in01 = imem02_in[31:28];
    59: op1_08_in01 = imem04_in[71:68];
    60: op1_08_in01 = reg_0395;
    61: op1_08_in01 = reg_0781;
    62: op1_08_in01 = imem00_in[67:64];
    63: op1_08_in01 = imem00_in[71:68];
    71: op1_08_in01 = imem00_in[71:68];
    64: op1_08_in01 = reg_0243;
    65: op1_08_in01 = reg_0505;
    66: op1_08_in01 = reg_0671;
    67: op1_08_in01 = reg_0056;
    68: op1_08_in01 = imem07_in[23:20];
    69: op1_08_in01 = imem02_in[99:96];
    70: op1_08_in01 = reg_0357;
    72: op1_08_in01 = reg_0140;
    74: op1_08_in01 = reg_0001;
    75: op1_08_in01 = reg_0765;
    76: op1_08_in01 = reg_0326;
    77: op1_08_in01 = imem07_in[91:88];
    78: op1_08_in01 = imem00_in[47:44];
    79: op1_08_in01 = imem02_in[119:116];
    80: op1_08_in01 = reg_0568;
    81: op1_08_in01 = reg_0642;
    82: op1_08_in01 = imem00_in[23:20];
    83: op1_08_in01 = imem05_in[51:48];
    84: op1_08_in01 = reg_0121;
    85: op1_08_in01 = reg_0579;
    86: op1_08_in01 = reg_0661;
    87: op1_08_in01 = imem00_in[11:8];
    88: op1_08_in01 = imem06_in[23:20];
    89: op1_08_in01 = reg_0420;
    90: op1_08_in01 = reg_0114;
    91: op1_08_in01 = reg_0669;
    92: op1_08_in01 = reg_0133;
    93: op1_08_in01 = reg_0062;
    94: op1_08_in01 = reg_0503;
    95: op1_08_in01 = imem06_in[39:36];
    96: op1_08_in01 = reg_0186;
    default: op1_08_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_08_inv01 = 1;
    8: op1_08_inv01 = 1;
    9: op1_08_inv01 = 1;
    12: op1_08_inv01 = 1;
    14: op1_08_inv01 = 1;
    15: op1_08_inv01 = 1;
    2: op1_08_inv01 = 1;
    21: op1_08_inv01 = 1;
    24: op1_08_inv01 = 1;
    25: op1_08_inv01 = 1;
    1: op1_08_inv01 = 1;
    27: op1_08_inv01 = 1;
    29: op1_08_inv01 = 1;
    31: op1_08_inv01 = 1;
    35: op1_08_inv01 = 1;
    37: op1_08_inv01 = 1;
    39: op1_08_inv01 = 1;
    41: op1_08_inv01 = 1;
    44: op1_08_inv01 = 1;
    45: op1_08_inv01 = 1;
    46: op1_08_inv01 = 1;
    47: op1_08_inv01 = 1;
    50: op1_08_inv01 = 1;
    52: op1_08_inv01 = 1;
    53: op1_08_inv01 = 1;
    54: op1_08_inv01 = 1;
    56: op1_08_inv01 = 1;
    58: op1_08_inv01 = 1;
    60: op1_08_inv01 = 1;
    64: op1_08_inv01 = 1;
    65: op1_08_inv01 = 1;
    66: op1_08_inv01 = 1;
    67: op1_08_inv01 = 1;
    68: op1_08_inv01 = 1;
    72: op1_08_inv01 = 1;
    74: op1_08_inv01 = 1;
    76: op1_08_inv01 = 1;
    78: op1_08_inv01 = 1;
    80: op1_08_inv01 = 1;
    81: op1_08_inv01 = 1;
    82: op1_08_inv01 = 1;
    83: op1_08_inv01 = 1;
    85: op1_08_inv01 = 1;
    86: op1_08_inv01 = 1;
    88: op1_08_inv01 = 1;
    90: op1_08_inv01 = 1;
    94: op1_08_inv01 = 1;
    95: op1_08_inv01 = 1;
    96: op1_08_inv01 = 1;
    default: op1_08_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in02 = imem05_in[39:36];
    5: op1_08_in02 = reg_0370;
    6: op1_08_in02 = imem07_in[67:64];
    7: op1_08_in02 = reg_0242;
    8: op1_08_in02 = imem05_in[63:60];
    9: op1_08_in02 = reg_0597;
    10: op1_08_in02 = reg_0266;
    11: op1_08_in02 = reg_0060;
    12: op1_08_in02 = imem00_in[39:36];
    20: op1_08_in02 = imem00_in[39:36];
    13: op1_08_in02 = reg_0225;
    14: op1_08_in02 = reg_0573;
    3: op1_08_in02 = imem07_in[55:52];
    15: op1_08_in02 = reg_0337;
    16: op1_08_in02 = imem00_in[83:80];
    17: op1_08_in02 = reg_0138;
    18: op1_08_in02 = imem00_in[127:124];
    19: op1_08_in02 = imem06_in[83:80];
    2: op1_08_in02 = imem07_in[107:104];
    21: op1_08_in02 = reg_0282;
    22: op1_08_in02 = imem05_in[71:68];
    83: op1_08_in02 = imem05_in[71:68];
    23: op1_08_in02 = reg_0293;
    24: op1_08_in02 = reg_0604;
    25: op1_08_in02 = reg_0103;
    26: op1_08_in02 = reg_0815;
    27: op1_08_in02 = imem00_in[71:68];
    28: op1_08_in02 = reg_0490;
    29: op1_08_in02 = reg_0005;
    30: op1_08_in02 = reg_0686;
    31: op1_08_in02 = reg_0749;
    32: op1_08_in02 = reg_0010;
    33: op1_08_in02 = imem07_in[27:24];
    34: op1_08_in02 = reg_0361;
    35: op1_08_in02 = reg_0126;
    84: op1_08_in02 = reg_0126;
    36: op1_08_in02 = reg_0391;
    37: op1_08_in02 = reg_0640;
    38: op1_08_in02 = reg_0090;
    39: op1_08_in02 = imem07_in[3:0];
    40: op1_08_in02 = reg_0748;
    41: op1_08_in02 = reg_0419;
    42: op1_08_in02 = reg_0589;
    43: op1_08_in02 = reg_0148;
    44: op1_08_in02 = reg_0670;
    45: op1_08_in02 = reg_0234;
    46: op1_08_in02 = imem05_in[31:28];
    47: op1_08_in02 = imem00_in[119:116];
    48: op1_08_in02 = reg_0101;
    49: op1_08_in02 = imem00_in[99:96];
    50: op1_08_in02 = reg_0715;
    51: op1_08_in02 = reg_0130;
    52: op1_08_in02 = imem07_in[47:44];
    53: op1_08_in02 = reg_0162;
    54: op1_08_in02 = reg_0114;
    55: op1_08_in02 = reg_0693;
    63: op1_08_in02 = reg_0693;
    56: op1_08_in02 = reg_0124;
    64: op1_08_in02 = reg_0124;
    57: op1_08_in02 = reg_0541;
    58: op1_08_in02 = imem02_in[75:72];
    59: op1_08_in02 = imem04_in[119:116];
    60: op1_08_in02 = reg_0387;
    61: op1_08_in02 = reg_0113;
    62: op1_08_in02 = imem00_in[87:84];
    65: op1_08_in02 = reg_0123;
    66: op1_08_in02 = reg_0678;
    67: op1_08_in02 = reg_0043;
    68: op1_08_in02 = imem07_in[51:48];
    69: op1_08_in02 = reg_0666;
    70: op1_08_in02 = reg_0384;
    71: op1_08_in02 = reg_0682;
    72: op1_08_in02 = reg_0702;
    73: op1_08_in02 = reg_0673;
    74: op1_08_in02 = reg_0007;
    75: op1_08_in02 = imem06_in[15:12];
    76: op1_08_in02 = reg_0797;
    77: op1_08_in02 = imem07_in[95:92];
    78: op1_08_in02 = imem00_in[63:60];
    79: op1_08_in02 = imem02_in[127:124];
    80: op1_08_in02 = reg_0572;
    81: op1_08_in02 = reg_0045;
    82: op1_08_in02 = imem00_in[35:32];
    85: op1_08_in02 = reg_0318;
    86: op1_08_in02 = reg_0752;
    87: op1_08_in02 = imem00_in[31:28];
    88: op1_08_in02 = imem06_in[39:36];
    89: op1_08_in02 = reg_0118;
    90: op1_08_in02 = reg_0760;
    91: op1_08_in02 = reg_0671;
    92: op1_08_in02 = reg_0788;
    93: op1_08_in02 = reg_0622;
    94: op1_08_in02 = reg_0508;
    95: op1_08_in02 = imem06_in[67:64];
    96: op1_08_in02 = reg_0607;
    default: op1_08_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_08_inv02 = 1;
    8: op1_08_inv02 = 1;
    10: op1_08_inv02 = 1;
    11: op1_08_inv02 = 1;
    13: op1_08_inv02 = 1;
    3: op1_08_inv02 = 1;
    16: op1_08_inv02 = 1;
    17: op1_08_inv02 = 1;
    18: op1_08_inv02 = 1;
    2: op1_08_inv02 = 1;
    21: op1_08_inv02 = 1;
    24: op1_08_inv02 = 1;
    25: op1_08_inv02 = 1;
    27: op1_08_inv02 = 1;
    28: op1_08_inv02 = 1;
    29: op1_08_inv02 = 1;
    30: op1_08_inv02 = 1;
    33: op1_08_inv02 = 1;
    35: op1_08_inv02 = 1;
    36: op1_08_inv02 = 1;
    37: op1_08_inv02 = 1;
    41: op1_08_inv02 = 1;
    44: op1_08_inv02 = 1;
    46: op1_08_inv02 = 1;
    50: op1_08_inv02 = 1;
    51: op1_08_inv02 = 1;
    55: op1_08_inv02 = 1;
    57: op1_08_inv02 = 1;
    62: op1_08_inv02 = 1;
    63: op1_08_inv02 = 1;
    66: op1_08_inv02 = 1;
    69: op1_08_inv02 = 1;
    71: op1_08_inv02 = 1;
    72: op1_08_inv02 = 1;
    73: op1_08_inv02 = 1;
    74: op1_08_inv02 = 1;
    76: op1_08_inv02 = 1;
    77: op1_08_inv02 = 1;
    78: op1_08_inv02 = 1;
    80: op1_08_inv02 = 1;
    82: op1_08_inv02 = 1;
    83: op1_08_inv02 = 1;
    84: op1_08_inv02 = 1;
    87: op1_08_inv02 = 1;
    89: op1_08_inv02 = 1;
    93: op1_08_inv02 = 1;
    94: op1_08_inv02 = 1;
    default: op1_08_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in03 = imem05_in[75:72];
    5: op1_08_in03 = reg_0322;
    6: op1_08_in03 = imem07_in[83:80];
    7: op1_08_in03 = reg_0228;
    8: op1_08_in03 = reg_0490;
    9: op1_08_in03 = reg_0595;
    10: op1_08_in03 = reg_0152;
    11: op1_08_in03 = reg_0073;
    12: op1_08_in03 = imem00_in[43:40];
    13: op1_08_in03 = reg_0235;
    14: op1_08_in03 = reg_0583;
    3: op1_08_in03 = imem07_in[87:84];
    15: op1_08_in03 = reg_0368;
    16: op1_08_in03 = imem00_in[111:108];
    17: op1_08_in03 = reg_0130;
    18: op1_08_in03 = reg_0682;
    19: op1_08_in03 = reg_0625;
    20: op1_08_in03 = imem00_in[75:72];
    2: op1_08_in03 = imem07_in[127:124];
    21: op1_08_in03 = reg_0277;
    22: op1_08_in03 = imem05_in[119:116];
    23: op1_08_in03 = reg_0268;
    24: op1_08_in03 = reg_0630;
    25: op1_08_in03 = reg_0120;
    26: op1_08_in03 = reg_0037;
    27: op1_08_in03 = imem00_in[103:100];
    62: op1_08_in03 = imem00_in[103:100];
    28: op1_08_in03 = reg_0495;
    29: op1_08_in03 = imem07_in[19:16];
    30: op1_08_in03 = reg_0674;
    31: op1_08_in03 = reg_0391;
    32: op1_08_in03 = reg_0004;
    33: op1_08_in03 = imem07_in[35:32];
    34: op1_08_in03 = reg_0343;
    35: op1_08_in03 = imem02_in[3:0];
    36: op1_08_in03 = reg_0568;
    37: op1_08_in03 = reg_0648;
    38: op1_08_in03 = reg_0736;
    39: op1_08_in03 = imem07_in[23:20];
    40: op1_08_in03 = reg_0329;
    41: op1_08_in03 = reg_0219;
    42: op1_08_in03 = reg_0384;
    43: op1_08_in03 = reg_0142;
    44: op1_08_in03 = reg_0690;
    45: op1_08_in03 = reg_0419;
    46: op1_08_in03 = imem05_in[51:48];
    47: op1_08_in03 = reg_0685;
    55: op1_08_in03 = reg_0685;
    48: op1_08_in03 = reg_0115;
    49: op1_08_in03 = reg_0697;
    50: op1_08_in03 = reg_0707;
    51: op1_08_in03 = reg_0140;
    52: op1_08_in03 = imem07_in[107:104];
    53: op1_08_in03 = reg_0167;
    54: op1_08_in03 = reg_0679;
    94: op1_08_in03 = reg_0679;
    56: op1_08_in03 = reg_0118;
    57: op1_08_in03 = reg_0530;
    58: op1_08_in03 = imem02_in[111:108];
    59: op1_08_in03 = reg_0545;
    60: op1_08_in03 = reg_0571;
    70: op1_08_in03 = reg_0571;
    85: op1_08_in03 = reg_0571;
    61: op1_08_in03 = reg_0288;
    63: op1_08_in03 = reg_0696;
    64: op1_08_in03 = reg_0119;
    65: op1_08_in03 = reg_0105;
    66: op1_08_in03 = imem02_in[11:8];
    67: op1_08_in03 = reg_0303;
    68: op1_08_in03 = imem07_in[67:64];
    69: op1_08_in03 = reg_0651;
    71: op1_08_in03 = reg_0693;
    72: op1_08_in03 = reg_0581;
    73: op1_08_in03 = reg_0660;
    74: op1_08_in03 = imem04_in[51:48];
    75: op1_08_in03 = imem06_in[27:24];
    76: op1_08_in03 = reg_0245;
    77: op1_08_in03 = reg_0728;
    78: op1_08_in03 = imem00_in[91:88];
    79: op1_08_in03 = reg_0642;
    80: op1_08_in03 = reg_0569;
    81: op1_08_in03 = reg_0621;
    82: op1_08_in03 = imem00_in[55:52];
    83: op1_08_in03 = reg_0791;
    84: op1_08_in03 = reg_0678;
    86: op1_08_in03 = imem07_in[3:0];
    87: op1_08_in03 = imem00_in[123:120];
    88: op1_08_in03 = imem06_in[51:48];
    89: op1_08_in03 = reg_0670;
    90: op1_08_in03 = reg_0241;
    91: op1_08_in03 = imem02_in[31:28];
    92: op1_08_in03 = reg_0146;
    93: op1_08_in03 = reg_0771;
    95: op1_08_in03 = imem06_in[83:80];
    96: op1_08_in03 = reg_0001;
    default: op1_08_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv03 = 1;
    9: op1_08_inv03 = 1;
    10: op1_08_inv03 = 1;
    13: op1_08_inv03 = 1;
    14: op1_08_inv03 = 1;
    16: op1_08_inv03 = 1;
    20: op1_08_inv03 = 1;
    21: op1_08_inv03 = 1;
    22: op1_08_inv03 = 1;
    23: op1_08_inv03 = 1;
    24: op1_08_inv03 = 1;
    26: op1_08_inv03 = 1;
    27: op1_08_inv03 = 1;
    30: op1_08_inv03 = 1;
    31: op1_08_inv03 = 1;
    32: op1_08_inv03 = 1;
    36: op1_08_inv03 = 1;
    37: op1_08_inv03 = 1;
    38: op1_08_inv03 = 1;
    39: op1_08_inv03 = 1;
    41: op1_08_inv03 = 1;
    42: op1_08_inv03 = 1;
    43: op1_08_inv03 = 1;
    45: op1_08_inv03 = 1;
    48: op1_08_inv03 = 1;
    51: op1_08_inv03 = 1;
    52: op1_08_inv03 = 1;
    53: op1_08_inv03 = 1;
    54: op1_08_inv03 = 1;
    55: op1_08_inv03 = 1;
    57: op1_08_inv03 = 1;
    62: op1_08_inv03 = 1;
    65: op1_08_inv03 = 1;
    67: op1_08_inv03 = 1;
    69: op1_08_inv03 = 1;
    70: op1_08_inv03 = 1;
    75: op1_08_inv03 = 1;
    76: op1_08_inv03 = 1;
    77: op1_08_inv03 = 1;
    79: op1_08_inv03 = 1;
    82: op1_08_inv03 = 1;
    85: op1_08_inv03 = 1;
    86: op1_08_inv03 = 1;
    88: op1_08_inv03 = 1;
    90: op1_08_inv03 = 1;
    92: op1_08_inv03 = 1;
    93: op1_08_inv03 = 1;
    94: op1_08_inv03 = 1;
    95: op1_08_inv03 = 1;
    default: op1_08_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in04 = imem05_in[91:88];
    5: op1_08_in04 = imem03_in[95:92];
    6: op1_08_in04 = imem07_in[119:116];
    7: op1_08_in04 = reg_0102;
    8: op1_08_in04 = reg_0789;
    9: op1_08_in04 = reg_0388;
    31: op1_08_in04 = reg_0388;
    10: op1_08_in04 = reg_0153;
    11: op1_08_in04 = imem03_in[59:56];
    12: op1_08_in04 = imem00_in[71:68];
    13: op1_08_in04 = reg_0246;
    14: op1_08_in04 = reg_0592;
    3: op1_08_in04 = imem07_in[127:124];
    15: op1_08_in04 = reg_0033;
    16: op1_08_in04 = reg_0697;
    17: op1_08_in04 = imem06_in[7:4];
    18: op1_08_in04 = reg_0696;
    19: op1_08_in04 = reg_0626;
    20: op1_08_in04 = imem00_in[99:96];
    2: op1_08_in04 = reg_0174;
    21: op1_08_in04 = reg_0744;
    22: op1_08_in04 = reg_0791;
    23: op1_08_in04 = reg_0298;
    24: op1_08_in04 = reg_0618;
    25: op1_08_in04 = reg_0112;
    26: op1_08_in04 = reg_0818;
    27: op1_08_in04 = reg_0686;
    63: op1_08_in04 = reg_0686;
    28: op1_08_in04 = reg_0783;
    29: op1_08_in04 = imem07_in[27:24];
    30: op1_08_in04 = reg_0678;
    32: op1_08_in04 = imem04_in[15:12];
    33: op1_08_in04 = imem07_in[39:36];
    34: op1_08_in04 = reg_0347;
    35: op1_08_in04 = imem02_in[55:52];
    36: op1_08_in04 = reg_0392;
    37: op1_08_in04 = reg_0638;
    38: op1_08_in04 = reg_0741;
    39: op1_08_in04 = imem07_in[107:104];
    40: op1_08_in04 = reg_0614;
    41: op1_08_in04 = reg_0106;
    42: op1_08_in04 = reg_0391;
    43: op1_08_in04 = reg_0134;
    44: op1_08_in04 = reg_0688;
    45: op1_08_in04 = imem02_in[35:32];
    46: op1_08_in04 = imem05_in[79:76];
    47: op1_08_in04 = reg_0676;
    49: op1_08_in04 = reg_0676;
    48: op1_08_in04 = reg_0127;
    50: op1_08_in04 = reg_0706;
    51: op1_08_in04 = imem06_in[63:60];
    52: op1_08_in04 = reg_0716;
    53: op1_08_in04 = reg_0166;
    54: op1_08_in04 = reg_0110;
    55: op1_08_in04 = reg_0698;
    56: op1_08_in04 = reg_0670;
    57: op1_08_in04 = reg_0535;
    58: op1_08_in04 = imem02_in[115:112];
    59: op1_08_in04 = reg_0056;
    60: op1_08_in04 = reg_0562;
    80: op1_08_in04 = reg_0562;
    61: op1_08_in04 = reg_0736;
    62: op1_08_in04 = reg_0682;
    64: op1_08_in04 = reg_0120;
    65: op1_08_in04 = reg_0672;
    66: op1_08_in04 = imem02_in[15:12];
    67: op1_08_in04 = reg_0280;
    68: op1_08_in04 = imem07_in[87:84];
    69: op1_08_in04 = reg_0484;
    70: op1_08_in04 = reg_0368;
    71: op1_08_in04 = reg_0492;
    78: op1_08_in04 = reg_0492;
    72: op1_08_in04 = reg_0356;
    73: op1_08_in04 = reg_0601;
    74: op1_08_in04 = imem04_in[71:68];
    75: op1_08_in04 = imem06_in[55:52];
    76: op1_08_in04 = reg_0383;
    77: op1_08_in04 = reg_0731;
    79: op1_08_in04 = reg_0703;
    81: op1_08_in04 = reg_0320;
    82: op1_08_in04 = imem00_in[83:80];
    83: op1_08_in04 = reg_0145;
    84: op1_08_in04 = reg_0607;
    85: op1_08_in04 = reg_0564;
    86: op1_08_in04 = imem07_in[15:12];
    87: op1_08_in04 = reg_0683;
    88: op1_08_in04 = imem06_in[115:112];
    89: op1_08_in04 = reg_0669;
    90: op1_08_in04 = reg_0423;
    91: op1_08_in04 = imem02_in[39:36];
    92: op1_08_in04 = reg_0782;
    93: op1_08_in04 = reg_0233;
    94: op1_08_in04 = reg_0065;
    95: op1_08_in04 = imem06_in[103:100];
    96: op1_08_in04 = reg_0800;
    default: op1_08_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv04 = 1;
    5: op1_08_inv04 = 1;
    6: op1_08_inv04 = 1;
    8: op1_08_inv04 = 1;
    9: op1_08_inv04 = 1;
    10: op1_08_inv04 = 1;
    14: op1_08_inv04 = 1;
    3: op1_08_inv04 = 1;
    18: op1_08_inv04 = 1;
    20: op1_08_inv04 = 1;
    23: op1_08_inv04 = 1;
    25: op1_08_inv04 = 1;
    27: op1_08_inv04 = 1;
    28: op1_08_inv04 = 1;
    32: op1_08_inv04 = 1;
    33: op1_08_inv04 = 1;
    35: op1_08_inv04 = 1;
    41: op1_08_inv04 = 1;
    44: op1_08_inv04 = 1;
    46: op1_08_inv04 = 1;
    48: op1_08_inv04 = 1;
    52: op1_08_inv04 = 1;
    54: op1_08_inv04 = 1;
    55: op1_08_inv04 = 1;
    56: op1_08_inv04 = 1;
    59: op1_08_inv04 = 1;
    62: op1_08_inv04 = 1;
    65: op1_08_inv04 = 1;
    68: op1_08_inv04 = 1;
    72: op1_08_inv04 = 1;
    76: op1_08_inv04 = 1;
    82: op1_08_inv04 = 1;
    83: op1_08_inv04 = 1;
    84: op1_08_inv04 = 1;
    87: op1_08_inv04 = 1;
    88: op1_08_inv04 = 1;
    89: op1_08_inv04 = 1;
    90: op1_08_inv04 = 1;
    91: op1_08_inv04 = 1;
    94: op1_08_inv04 = 1;
    default: op1_08_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in05 = imem05_in[95:92];
    5: op1_08_in05 = imem04_in[23:20];
    6: op1_08_in05 = reg_0717;
    7: op1_08_in05 = reg_0107;
    8: op1_08_in05 = reg_0793;
    9: op1_08_in05 = reg_0377;
    10: op1_08_in05 = reg_0140;
    11: op1_08_in05 = imem03_in[63:60];
    12: op1_08_in05 = reg_0698;
    18: op1_08_in05 = reg_0698;
    62: op1_08_in05 = reg_0698;
    13: op1_08_in05 = reg_0242;
    40: op1_08_in05 = reg_0242;
    14: op1_08_in05 = reg_0600;
    3: op1_08_in05 = reg_0446;
    15: op1_08_in05 = reg_0753;
    16: op1_08_in05 = reg_0694;
    17: op1_08_in05 = imem06_in[27:24];
    19: op1_08_in05 = reg_0611;
    20: op1_08_in05 = reg_0695;
    2: op1_08_in05 = reg_0167;
    21: op1_08_in05 = reg_0734;
    22: op1_08_in05 = reg_0788;
    23: op1_08_in05 = reg_0065;
    24: op1_08_in05 = reg_0612;
    25: op1_08_in05 = reg_0317;
    26: op1_08_in05 = imem07_in[11:8];
    27: op1_08_in05 = reg_0688;
    28: op1_08_in05 = reg_0279;
    38: op1_08_in05 = reg_0279;
    29: op1_08_in05 = imem07_in[31:28];
    86: op1_08_in05 = imem07_in[31:28];
    30: op1_08_in05 = reg_0668;
    31: op1_08_in05 = reg_0385;
    32: op1_08_in05 = imem04_in[43:40];
    96: op1_08_in05 = imem04_in[43:40];
    33: op1_08_in05 = imem07_in[87:84];
    34: op1_08_in05 = reg_0769;
    35: op1_08_in05 = imem02_in[119:116];
    36: op1_08_in05 = reg_0398;
    37: op1_08_in05 = reg_0636;
    39: op1_08_in05 = reg_0722;
    41: op1_08_in05 = imem02_in[43:40];
    42: op1_08_in05 = reg_0575;
    43: op1_08_in05 = imem06_in[15:12];
    44: op1_08_in05 = reg_0687;
    47: op1_08_in05 = reg_0687;
    45: op1_08_in05 = imem02_in[111:108];
    46: op1_08_in05 = imem05_in[103:100];
    48: op1_08_in05 = reg_0110;
    49: op1_08_in05 = reg_0689;
    50: op1_08_in05 = reg_0053;
    51: op1_08_in05 = reg_0624;
    52: op1_08_in05 = reg_0704;
    54: op1_08_in05 = reg_0111;
    55: op1_08_in05 = reg_0749;
    63: op1_08_in05 = reg_0749;
    56: op1_08_in05 = reg_0671;
    57: op1_08_in05 = reg_0531;
    58: op1_08_in05 = reg_0657;
    59: op1_08_in05 = reg_0083;
    60: op1_08_in05 = reg_0747;
    61: op1_08_in05 = reg_0309;
    64: op1_08_in05 = reg_0675;
    65: op1_08_in05 = reg_0675;
    66: op1_08_in05 = imem02_in[87:84];
    67: op1_08_in05 = reg_0292;
    68: op1_08_in05 = imem07_in[99:96];
    69: op1_08_in05 = reg_0641;
    70: op1_08_in05 = reg_0403;
    71: op1_08_in05 = reg_0686;
    72: op1_08_in05 = reg_0414;
    73: op1_08_in05 = imem02_in[63:60];
    74: op1_08_in05 = imem04_in[79:76];
    75: op1_08_in05 = imem06_in[83:80];
    76: op1_08_in05 = reg_0812;
    77: op1_08_in05 = reg_0239;
    78: op1_08_in05 = reg_0744;
    87: op1_08_in05 = reg_0744;
    79: op1_08_in05 = reg_0427;
    80: op1_08_in05 = reg_0496;
    81: op1_08_in05 = reg_0586;
    82: op1_08_in05 = imem00_in[87:84];
    83: op1_08_in05 = reg_0795;
    84: op1_08_in05 = reg_0541;
    85: op1_08_in05 = reg_0013;
    88: op1_08_in05 = reg_0715;
    89: op1_08_in05 = reg_0674;
    90: op1_08_in05 = reg_0421;
    91: op1_08_in05 = imem02_in[67:64];
    92: op1_08_in05 = reg_0732;
    93: op1_08_in05 = imem05_in[11:8];
    94: op1_08_in05 = reg_0643;
    95: op1_08_in05 = reg_0289;
    default: op1_08_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv05 = 1;
    8: op1_08_inv05 = 1;
    10: op1_08_inv05 = 1;
    12: op1_08_inv05 = 1;
    13: op1_08_inv05 = 1;
    3: op1_08_inv05 = 1;
    16: op1_08_inv05 = 1;
    18: op1_08_inv05 = 1;
    21: op1_08_inv05 = 1;
    22: op1_08_inv05 = 1;
    24: op1_08_inv05 = 1;
    26: op1_08_inv05 = 1;
    27: op1_08_inv05 = 1;
    28: op1_08_inv05 = 1;
    31: op1_08_inv05 = 1;
    32: op1_08_inv05 = 1;
    34: op1_08_inv05 = 1;
    35: op1_08_inv05 = 1;
    37: op1_08_inv05 = 1;
    38: op1_08_inv05 = 1;
    42: op1_08_inv05 = 1;
    44: op1_08_inv05 = 1;
    45: op1_08_inv05 = 1;
    46: op1_08_inv05 = 1;
    48: op1_08_inv05 = 1;
    50: op1_08_inv05 = 1;
    51: op1_08_inv05 = 1;
    52: op1_08_inv05 = 1;
    54: op1_08_inv05 = 1;
    58: op1_08_inv05 = 1;
    59: op1_08_inv05 = 1;
    60: op1_08_inv05 = 1;
    67: op1_08_inv05 = 1;
    70: op1_08_inv05 = 1;
    74: op1_08_inv05 = 1;
    75: op1_08_inv05 = 1;
    76: op1_08_inv05 = 1;
    79: op1_08_inv05 = 1;
    80: op1_08_inv05 = 1;
    84: op1_08_inv05 = 1;
    85: op1_08_inv05 = 1;
    87: op1_08_inv05 = 1;
    91: op1_08_inv05 = 1;
    92: op1_08_inv05 = 1;
    93: op1_08_inv05 = 1;
    94: op1_08_inv05 = 1;
    95: op1_08_inv05 = 1;
    default: op1_08_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in06 = imem05_in[115:112];
    5: op1_08_in06 = imem04_in[27:24];
    6: op1_08_in06 = reg_0724;
    7: op1_08_in06 = imem02_in[11:8];
    8: op1_08_in06 = reg_0780;
    9: op1_08_in06 = reg_0322;
    10: op1_08_in06 = imem06_in[51:48];
    11: op1_08_in06 = imem03_in[79:76];
    12: op1_08_in06 = reg_0691;
    13: op1_08_in06 = reg_0237;
    14: op1_08_in06 = reg_0578;
    3: op1_08_in06 = reg_0161;
    15: op1_08_in06 = reg_0816;
    16: op1_08_in06 = reg_0698;
    17: op1_08_in06 = imem06_in[71:68];
    18: op1_08_in06 = reg_0688;
    19: op1_08_in06 = reg_0618;
    20: op1_08_in06 = reg_0696;
    2: op1_08_in06 = reg_0164;
    21: op1_08_in06 = reg_0285;
    22: op1_08_in06 = reg_0493;
    23: op1_08_in06 = reg_0075;
    24: op1_08_in06 = reg_0356;
    25: op1_08_in06 = reg_0264;
    26: op1_08_in06 = imem07_in[27:24];
    27: op1_08_in06 = reg_0457;
    28: op1_08_in06 = reg_0139;
    29: op1_08_in06 = imem07_in[51:48];
    30: op1_08_in06 = reg_0675;
    31: op1_08_in06 = reg_0572;
    32: op1_08_in06 = imem04_in[99:96];
    33: op1_08_in06 = reg_0731;
    88: op1_08_in06 = reg_0731;
    34: op1_08_in06 = reg_0531;
    35: op1_08_in06 = reg_0655;
    36: op1_08_in06 = reg_0000;
    37: op1_08_in06 = reg_0320;
    38: op1_08_in06 = reg_0742;
    39: op1_08_in06 = reg_0721;
    40: op1_08_in06 = reg_0620;
    41: op1_08_in06 = imem02_in[63:60];
    42: op1_08_in06 = reg_0569;
    43: op1_08_in06 = imem06_in[43:40];
    44: op1_08_in06 = reg_0692;
    45: op1_08_in06 = imem02_in[115:112];
    46: op1_08_in06 = imem05_in[123:120];
    47: op1_08_in06 = reg_0463;
    48: op1_08_in06 = imem02_in[35:32];
    49: op1_08_in06 = reg_0690;
    78: op1_08_in06 = reg_0690;
    50: op1_08_in06 = reg_0267;
    51: op1_08_in06 = reg_0416;
    52: op1_08_in06 = reg_0719;
    54: op1_08_in06 = imem00_in[15:12];
    55: op1_08_in06 = reg_0658;
    63: op1_08_in06 = reg_0658;
    56: op1_08_in06 = reg_0674;
    57: op1_08_in06 = reg_0526;
    58: op1_08_in06 = reg_0661;
    59: op1_08_in06 = reg_0555;
    60: op1_08_in06 = reg_0396;
    61: op1_08_in06 = reg_0245;
    62: op1_08_in06 = reg_0686;
    64: op1_08_in06 = reg_0669;
    65: op1_08_in06 = reg_0106;
    66: op1_08_in06 = imem02_in[103:100];
    67: op1_08_in06 = reg_0610;
    68: op1_08_in06 = imem07_in[103:100];
    69: op1_08_in06 = reg_0426;
    70: op1_08_in06 = reg_0387;
    80: op1_08_in06 = reg_0387;
    71: op1_08_in06 = reg_0749;
    87: op1_08_in06 = reg_0749;
    72: op1_08_in06 = reg_0527;
    73: op1_08_in06 = imem02_in[79:76];
    74: op1_08_in06 = imem04_in[87:84];
    75: op1_08_in06 = reg_0115;
    76: op1_08_in06 = reg_0147;
    77: op1_08_in06 = reg_0434;
    79: op1_08_in06 = reg_0581;
    81: op1_08_in06 = reg_0359;
    82: op1_08_in06 = reg_0695;
    83: op1_08_in06 = reg_0315;
    84: op1_08_in06 = reg_0081;
    85: op1_08_in06 = reg_0007;
    86: op1_08_in06 = imem07_in[39:36];
    89: op1_08_in06 = reg_0678;
    90: op1_08_in06 = reg_0054;
    91: op1_08_in06 = imem02_in[107:104];
    92: op1_08_in06 = reg_0492;
    93: op1_08_in06 = imem05_in[23:20];
    94: op1_08_in06 = reg_0233;
    95: op1_08_in06 = reg_0817;
    96: op1_08_in06 = imem04_in[47:44];
    default: op1_08_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv06 = 1;
    6: op1_08_inv06 = 1;
    7: op1_08_inv06 = 1;
    10: op1_08_inv06 = 1;
    11: op1_08_inv06 = 1;
    15: op1_08_inv06 = 1;
    19: op1_08_inv06 = 1;
    20: op1_08_inv06 = 1;
    2: op1_08_inv06 = 1;
    21: op1_08_inv06 = 1;
    24: op1_08_inv06 = 1;
    25: op1_08_inv06 = 1;
    26: op1_08_inv06 = 1;
    27: op1_08_inv06 = 1;
    28: op1_08_inv06 = 1;
    29: op1_08_inv06 = 1;
    31: op1_08_inv06 = 1;
    35: op1_08_inv06 = 1;
    38: op1_08_inv06 = 1;
    41: op1_08_inv06 = 1;
    45: op1_08_inv06 = 1;
    47: op1_08_inv06 = 1;
    48: op1_08_inv06 = 1;
    49: op1_08_inv06 = 1;
    50: op1_08_inv06 = 1;
    54: op1_08_inv06 = 1;
    57: op1_08_inv06 = 1;
    59: op1_08_inv06 = 1;
    60: op1_08_inv06 = 1;
    62: op1_08_inv06 = 1;
    63: op1_08_inv06 = 1;
    65: op1_08_inv06 = 1;
    66: op1_08_inv06 = 1;
    67: op1_08_inv06 = 1;
    70: op1_08_inv06 = 1;
    71: op1_08_inv06 = 1;
    72: op1_08_inv06 = 1;
    74: op1_08_inv06 = 1;
    75: op1_08_inv06 = 1;
    77: op1_08_inv06 = 1;
    78: op1_08_inv06 = 1;
    80: op1_08_inv06 = 1;
    82: op1_08_inv06 = 1;
    84: op1_08_inv06 = 1;
    85: op1_08_inv06 = 1;
    86: op1_08_inv06 = 1;
    88: op1_08_inv06 = 1;
    89: op1_08_inv06 = 1;
    90: op1_08_inv06 = 1;
    91: op1_08_inv06 = 1;
    92: op1_08_inv06 = 1;
    94: op1_08_inv06 = 1;
    95: op1_08_inv06 = 1;
    default: op1_08_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in07 = reg_0488;
    5: op1_08_in07 = imem04_in[43:40];
    6: op1_08_in07 = reg_0711;
    7: op1_08_in07 = imem02_in[83:80];
    8: op1_08_in07 = reg_0787;
    9: op1_08_in07 = reg_0309;
    10: op1_08_in07 = imem06_in[59:56];
    11: op1_08_in07 = imem03_in[99:96];
    12: op1_08_in07 = reg_0675;
    13: op1_08_in07 = reg_0245;
    14: op1_08_in07 = reg_0590;
    72: op1_08_in07 = reg_0590;
    3: op1_08_in07 = reg_0162;
    15: op1_08_in07 = reg_0029;
    40: op1_08_in07 = reg_0029;
    16: op1_08_in07 = reg_0677;
    17: op1_08_in07 = imem06_in[79:76];
    18: op1_08_in07 = reg_0451;
    19: op1_08_in07 = reg_0615;
    20: op1_08_in07 = reg_0686;
    2: op1_08_in07 = reg_0185;
    21: op1_08_in07 = reg_0086;
    22: op1_08_in07 = reg_0794;
    23: op1_08_in07 = reg_0256;
    61: op1_08_in07 = reg_0256;
    24: op1_08_in07 = reg_0405;
    25: op1_08_in07 = reg_0259;
    26: op1_08_in07 = imem07_in[39:36];
    27: op1_08_in07 = reg_0469;
    28: op1_08_in07 = reg_0141;
    29: op1_08_in07 = imem07_in[111:108];
    30: op1_08_in07 = reg_0476;
    31: op1_08_in07 = reg_0398;
    32: op1_08_in07 = imem04_in[123:120];
    33: op1_08_in07 = reg_0726;
    34: op1_08_in07 = reg_0094;
    35: op1_08_in07 = reg_0638;
    36: op1_08_in07 = reg_0006;
    37: op1_08_in07 = reg_0356;
    38: op1_08_in07 = reg_0272;
    39: op1_08_in07 = reg_0725;
    41: op1_08_in07 = reg_0654;
    42: op1_08_in07 = reg_0562;
    43: op1_08_in07 = reg_0289;
    44: op1_08_in07 = reg_0464;
    45: op1_08_in07 = reg_0337;
    46: op1_08_in07 = reg_0792;
    47: op1_08_in07 = reg_0465;
    48: op1_08_in07 = imem02_in[43:40];
    49: op1_08_in07 = reg_0688;
    50: op1_08_in07 = reg_0448;
    51: op1_08_in07 = reg_0371;
    52: op1_08_in07 = reg_0720;
    54: op1_08_in07 = imem00_in[79:76];
    55: op1_08_in07 = reg_0758;
    56: op1_08_in07 = reg_0121;
    57: op1_08_in07 = reg_0093;
    58: op1_08_in07 = reg_0667;
    59: op1_08_in07 = reg_0060;
    60: op1_08_in07 = reg_0374;
    62: op1_08_in07 = reg_0247;
    63: op1_08_in07 = reg_0494;
    64: op1_08_in07 = reg_0671;
    65: op1_08_in07 = reg_0127;
    66: op1_08_in07 = imem02_in[127:124];
    67: op1_08_in07 = reg_0513;
    68: op1_08_in07 = imem07_in[119:116];
    69: op1_08_in07 = reg_0364;
    70: op1_08_in07 = reg_0000;
    71: op1_08_in07 = reg_0658;
    73: op1_08_in07 = imem02_in[111:108];
    74: op1_08_in07 = reg_0552;
    75: op1_08_in07 = reg_0762;
    76: op1_08_in07 = reg_0827;
    77: op1_08_in07 = reg_0446;
    78: op1_08_in07 = reg_0691;
    87: op1_08_in07 = reg_0691;
    79: op1_08_in07 = reg_0363;
    80: op1_08_in07 = reg_0623;
    81: op1_08_in07 = reg_0345;
    82: op1_08_in07 = reg_0492;
    83: op1_08_in07 = reg_0486;
    84: op1_08_in07 = reg_0392;
    85: op1_08_in07 = imem04_in[71:68];
    86: op1_08_in07 = imem07_in[83:80];
    88: op1_08_in07 = reg_0295;
    89: op1_08_in07 = imem02_in[3:0];
    90: op1_08_in07 = reg_0567;
    91: op1_08_in07 = reg_0533;
    92: op1_08_in07 = reg_0580;
    93: op1_08_in07 = imem05_in[43:40];
    94: op1_08_in07 = reg_0416;
    95: op1_08_in07 = reg_0814;
    96: op1_08_in07 = imem04_in[67:64];
    default: op1_08_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv07 = 1;
    6: op1_08_inv07 = 1;
    11: op1_08_inv07 = 1;
    12: op1_08_inv07 = 1;
    13: op1_08_inv07 = 1;
    14: op1_08_inv07 = 1;
    3: op1_08_inv07 = 1;
    16: op1_08_inv07 = 1;
    18: op1_08_inv07 = 1;
    21: op1_08_inv07 = 1;
    22: op1_08_inv07 = 1;
    25: op1_08_inv07 = 1;
    30: op1_08_inv07 = 1;
    31: op1_08_inv07 = 1;
    34: op1_08_inv07 = 1;
    35: op1_08_inv07 = 1;
    36: op1_08_inv07 = 1;
    37: op1_08_inv07 = 1;
    38: op1_08_inv07 = 1;
    39: op1_08_inv07 = 1;
    42: op1_08_inv07 = 1;
    43: op1_08_inv07 = 1;
    48: op1_08_inv07 = 1;
    49: op1_08_inv07 = 1;
    50: op1_08_inv07 = 1;
    51: op1_08_inv07 = 1;
    52: op1_08_inv07 = 1;
    54: op1_08_inv07 = 1;
    58: op1_08_inv07 = 1;
    60: op1_08_inv07 = 1;
    61: op1_08_inv07 = 1;
    63: op1_08_inv07 = 1;
    64: op1_08_inv07 = 1;
    65: op1_08_inv07 = 1;
    66: op1_08_inv07 = 1;
    68: op1_08_inv07 = 1;
    69: op1_08_inv07 = 1;
    72: op1_08_inv07 = 1;
    73: op1_08_inv07 = 1;
    79: op1_08_inv07 = 1;
    80: op1_08_inv07 = 1;
    82: op1_08_inv07 = 1;
    83: op1_08_inv07 = 1;
    84: op1_08_inv07 = 1;
    85: op1_08_inv07 = 1;
    90: op1_08_inv07 = 1;
    91: op1_08_inv07 = 1;
    95: op1_08_inv07 = 1;
    96: op1_08_inv07 = 1;
    default: op1_08_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in08 = reg_0489;
    5: op1_08_in08 = imem04_in[79:76];
    6: op1_08_in08 = reg_0707;
    7: op1_08_in08 = imem02_in[91:88];
    8: op1_08_in08 = reg_0268;
    9: op1_08_in08 = reg_0807;
    10: op1_08_in08 = imem06_in[67:64];
    11: op1_08_in08 = reg_0586;
    58: op1_08_in08 = reg_0586;
    12: op1_08_in08 = reg_0680;
    63: op1_08_in08 = reg_0680;
    13: op1_08_in08 = reg_0243;
    14: op1_08_in08 = reg_0576;
    3: op1_08_in08 = reg_0163;
    15: op1_08_in08 = imem07_in[31:28];
    16: op1_08_in08 = reg_0678;
    17: op1_08_in08 = imem06_in[83:80];
    18: op1_08_in08 = reg_0472;
    19: op1_08_in08 = reg_0612;
    20: op1_08_in08 = reg_0679;
    2: op1_08_in08 = reg_0170;
    21: op1_08_in08 = reg_0089;
    22: op1_08_in08 = reg_0783;
    23: op1_08_in08 = imem05_in[15:12];
    24: op1_08_in08 = reg_0383;
    25: op1_08_in08 = reg_0311;
    26: op1_08_in08 = imem07_in[47:44];
    27: op1_08_in08 = reg_0481;
    28: op1_08_in08 = reg_0372;
    29: op1_08_in08 = reg_0725;
    30: op1_08_in08 = reg_0458;
    31: op1_08_in08 = reg_0396;
    32: op1_08_in08 = reg_0544;
    33: op1_08_in08 = reg_0703;
    34: op1_08_in08 = imem03_in[55:52];
    35: op1_08_in08 = reg_0348;
    36: op1_08_in08 = reg_0013;
    37: op1_08_in08 = reg_0073;
    38: op1_08_in08 = reg_0732;
    39: op1_08_in08 = reg_0724;
    40: op1_08_in08 = imem07_in[15:12];
    41: op1_08_in08 = reg_0656;
    42: op1_08_in08 = reg_0012;
    43: op1_08_in08 = reg_0628;
    44: op1_08_in08 = reg_0187;
    45: op1_08_in08 = reg_0254;
    46: op1_08_in08 = reg_0488;
    47: op1_08_in08 = reg_0464;
    48: op1_08_in08 = imem02_in[71:68];
    49: op1_08_in08 = reg_0669;
    50: op1_08_in08 = reg_0435;
    51: op1_08_in08 = reg_0298;
    52: op1_08_in08 = reg_0726;
    54: op1_08_in08 = imem00_in[99:96];
    55: op1_08_in08 = reg_0699;
    56: op1_08_in08 = imem02_in[15:12];
    57: op1_08_in08 = imem03_in[3:0];
    59: op1_08_in08 = reg_0523;
    60: op1_08_in08 = reg_0019;
    61: op1_08_in08 = reg_0103;
    62: op1_08_in08 = reg_0465;
    64: op1_08_in08 = imem02_in[35:32];
    65: op1_08_in08 = imem02_in[11:8];
    89: op1_08_in08 = imem02_in[11:8];
    66: op1_08_in08 = reg_0785;
    67: op1_08_in08 = reg_0296;
    68: op1_08_in08 = reg_0716;
    69: op1_08_in08 = reg_0359;
    84: op1_08_in08 = reg_0359;
    70: op1_08_in08 = reg_0003;
    71: op1_08_in08 = reg_0691;
    72: op1_08_in08 = reg_0343;
    73: op1_08_in08 = reg_0142;
    74: op1_08_in08 = reg_0510;
    75: op1_08_in08 = reg_0401;
    76: op1_08_in08 = reg_0734;
    77: op1_08_in08 = reg_0175;
    78: op1_08_in08 = reg_0758;
    79: op1_08_in08 = reg_0365;
    80: op1_08_in08 = imem04_in[3:0];
    81: op1_08_in08 = reg_0324;
    82: op1_08_in08 = reg_0689;
    83: op1_08_in08 = reg_0735;
    85: op1_08_in08 = imem04_in[87:84];
    86: op1_08_in08 = imem07_in[95:92];
    87: op1_08_in08 = reg_0450;
    88: op1_08_in08 = reg_0636;
    90: op1_08_in08 = reg_0220;
    91: op1_08_in08 = reg_0639;
    92: op1_08_in08 = reg_0751;
    93: op1_08_in08 = imem05_in[55:52];
    94: op1_08_in08 = imem05_in[7:4];
    95: op1_08_in08 = reg_0619;
    96: op1_08_in08 = imem04_in[111:108];
    default: op1_08_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv08 = 1;
    5: op1_08_inv08 = 1;
    6: op1_08_inv08 = 1;
    8: op1_08_inv08 = 1;
    10: op1_08_inv08 = 1;
    11: op1_08_inv08 = 1;
    14: op1_08_inv08 = 1;
    15: op1_08_inv08 = 1;
    16: op1_08_inv08 = 1;
    17: op1_08_inv08 = 1;
    18: op1_08_inv08 = 1;
    20: op1_08_inv08 = 1;
    2: op1_08_inv08 = 1;
    21: op1_08_inv08 = 1;
    25: op1_08_inv08 = 1;
    27: op1_08_inv08 = 1;
    28: op1_08_inv08 = 1;
    33: op1_08_inv08 = 1;
    35: op1_08_inv08 = 1;
    36: op1_08_inv08 = 1;
    37: op1_08_inv08 = 1;
    38: op1_08_inv08 = 1;
    39: op1_08_inv08 = 1;
    41: op1_08_inv08 = 1;
    42: op1_08_inv08 = 1;
    44: op1_08_inv08 = 1;
    45: op1_08_inv08 = 1;
    46: op1_08_inv08 = 1;
    48: op1_08_inv08 = 1;
    49: op1_08_inv08 = 1;
    50: op1_08_inv08 = 1;
    52: op1_08_inv08 = 1;
    54: op1_08_inv08 = 1;
    57: op1_08_inv08 = 1;
    59: op1_08_inv08 = 1;
    62: op1_08_inv08 = 1;
    65: op1_08_inv08 = 1;
    68: op1_08_inv08 = 1;
    70: op1_08_inv08 = 1;
    71: op1_08_inv08 = 1;
    73: op1_08_inv08 = 1;
    74: op1_08_inv08 = 1;
    75: op1_08_inv08 = 1;
    76: op1_08_inv08 = 1;
    79: op1_08_inv08 = 1;
    80: op1_08_inv08 = 1;
    82: op1_08_inv08 = 1;
    86: op1_08_inv08 = 1;
    90: op1_08_inv08 = 1;
    93: op1_08_inv08 = 1;
    94: op1_08_inv08 = 1;
    96: op1_08_inv08 = 1;
    default: op1_08_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in09 = reg_0215;
    5: op1_08_in09 = imem04_in[107:104];
    6: op1_08_in09 = reg_0700;
    7: op1_08_in09 = imem02_in[115:112];
    8: op1_08_in09 = reg_0269;
    9: op1_08_in09 = reg_0804;
    10: op1_08_in09 = imem06_in[107:104];
    17: op1_08_in09 = imem06_in[107:104];
    11: op1_08_in09 = reg_0572;
    12: op1_08_in09 = reg_0455;
    13: op1_08_in09 = reg_0105;
    14: op1_08_in09 = reg_0360;
    69: op1_08_in09 = reg_0360;
    15: op1_08_in09 = reg_0722;
    16: op1_08_in09 = reg_0699;
    18: op1_08_in09 = reg_0480;
    27: op1_08_in09 = reg_0480;
    19: op1_08_in09 = reg_0349;
    20: op1_08_in09 = reg_0675;
    2: op1_08_in09 = reg_0173;
    21: op1_08_in09 = reg_0136;
    22: op1_08_in09 = reg_0787;
    23: op1_08_in09 = imem05_in[67:64];
    24: op1_08_in09 = reg_0404;
    25: op1_08_in09 = reg_0657;
    66: op1_08_in09 = reg_0657;
    26: op1_08_in09 = imem07_in[71:68];
    28: op1_08_in09 = reg_0338;
    29: op1_08_in09 = reg_0701;
    30: op1_08_in09 = reg_0187;
    31: op1_08_in09 = reg_0374;
    32: op1_08_in09 = reg_0328;
    33: op1_08_in09 = reg_0712;
    34: op1_08_in09 = imem03_in[107:104];
    35: op1_08_in09 = reg_0363;
    36: op1_08_in09 = imem04_in[63:60];
    37: op1_08_in09 = reg_0518;
    38: op1_08_in09 = reg_0086;
    39: op1_08_in09 = reg_0708;
    40: op1_08_in09 = imem07_in[43:40];
    41: op1_08_in09 = reg_0643;
    42: op1_08_in09 = reg_0808;
    43: op1_08_in09 = reg_0604;
    44: op1_08_in09 = reg_0194;
    45: op1_08_in09 = reg_0664;
    46: op1_08_in09 = reg_0793;
    47: op1_08_in09 = reg_0473;
    48: op1_08_in09 = imem02_in[107:104];
    49: op1_08_in09 = reg_0450;
    62: op1_08_in09 = reg_0450;
    50: op1_08_in09 = reg_0180;
    51: op1_08_in09 = reg_0766;
    52: op1_08_in09 = reg_0714;
    54: op1_08_in09 = reg_0457;
    55: op1_08_in09 = reg_0469;
    56: op1_08_in09 = imem02_in[47:44];
    57: op1_08_in09 = imem03_in[51:48];
    58: op1_08_in09 = reg_0581;
    59: op1_08_in09 = reg_0516;
    60: op1_08_in09 = reg_0008;
    61: op1_08_in09 = reg_0226;
    63: op1_08_in09 = reg_0247;
    96: op1_08_in09 = reg_0247;
    64: op1_08_in09 = imem02_in[59:56];
    65: op1_08_in09 = imem02_in[99:96];
    67: op1_08_in09 = reg_0336;
    68: op1_08_in09 = reg_0717;
    70: op1_08_in09 = reg_0803;
    71: op1_08_in09 = reg_0688;
    72: op1_08_in09 = reg_0323;
    73: op1_08_in09 = reg_0138;
    92: op1_08_in09 = reg_0138;
    74: op1_08_in09 = reg_0547;
    75: op1_08_in09 = reg_0242;
    76: op1_08_in09 = imem06_in[47:44];
    77: op1_08_in09 = reg_0167;
    78: op1_08_in09 = reg_0407;
    79: op1_08_in09 = reg_0514;
    80: op1_08_in09 = imem04_in[47:44];
    81: op1_08_in09 = reg_0527;
    82: op1_08_in09 = reg_0691;
    83: op1_08_in09 = reg_0383;
    84: op1_08_in09 = reg_0345;
    85: op1_08_in09 = imem04_in[119:116];
    86: op1_08_in09 = imem07_in[111:108];
    87: op1_08_in09 = reg_0461;
    88: op1_08_in09 = reg_0061;
    89: op1_08_in09 = imem02_in[35:32];
    90: op1_08_in09 = reg_0425;
    91: op1_08_in09 = reg_0342;
    93: op1_08_in09 = imem05_in[83:80];
    94: op1_08_in09 = imem05_in[51:48];
    95: op1_08_in09 = reg_0354;
    default: op1_08_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_08_inv09 = 1;
    8: op1_08_inv09 = 1;
    9: op1_08_inv09 = 1;
    12: op1_08_inv09 = 1;
    13: op1_08_inv09 = 1;
    14: op1_08_inv09 = 1;
    16: op1_08_inv09 = 1;
    17: op1_08_inv09 = 1;
    18: op1_08_inv09 = 1;
    2: op1_08_inv09 = 1;
    22: op1_08_inv09 = 1;
    23: op1_08_inv09 = 1;
    24: op1_08_inv09 = 1;
    25: op1_08_inv09 = 1;
    28: op1_08_inv09 = 1;
    30: op1_08_inv09 = 1;
    32: op1_08_inv09 = 1;
    35: op1_08_inv09 = 1;
    36: op1_08_inv09 = 1;
    38: op1_08_inv09 = 1;
    39: op1_08_inv09 = 1;
    41: op1_08_inv09 = 1;
    42: op1_08_inv09 = 1;
    43: op1_08_inv09 = 1;
    44: op1_08_inv09 = 1;
    45: op1_08_inv09 = 1;
    47: op1_08_inv09 = 1;
    52: op1_08_inv09 = 1;
    56: op1_08_inv09 = 1;
    59: op1_08_inv09 = 1;
    60: op1_08_inv09 = 1;
    61: op1_08_inv09 = 1;
    65: op1_08_inv09 = 1;
    67: op1_08_inv09 = 1;
    68: op1_08_inv09 = 1;
    73: op1_08_inv09 = 1;
    74: op1_08_inv09 = 1;
    75: op1_08_inv09 = 1;
    76: op1_08_inv09 = 1;
    81: op1_08_inv09 = 1;
    82: op1_08_inv09 = 1;
    84: op1_08_inv09 = 1;
    87: op1_08_inv09 = 1;
    89: op1_08_inv09 = 1;
    90: op1_08_inv09 = 1;
    91: op1_08_inv09 = 1;
    96: op1_08_inv09 = 1;
    default: op1_08_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in10 = reg_0261;
    5: op1_08_in10 = imem04_in[127:124];
    6: op1_08_in10 = reg_0429;
    7: op1_08_in10 = reg_0642;
    8: op1_08_in10 = reg_0244;
    9: op1_08_in10 = reg_0801;
    10: op1_08_in10 = reg_0614;
    11: op1_08_in10 = reg_0594;
    12: op1_08_in10 = reg_0470;
    18: op1_08_in10 = reg_0470;
    13: op1_08_in10 = reg_0111;
    14: op1_08_in10 = reg_0362;
    15: op1_08_in10 = reg_0730;
    16: op1_08_in10 = reg_0463;
    17: op1_08_in10 = reg_0619;
    19: op1_08_in10 = reg_0392;
    20: op1_08_in10 = reg_0680;
    78: op1_08_in10 = reg_0680;
    21: op1_08_in10 = reg_0151;
    22: op1_08_in10 = reg_0741;
    23: op1_08_in10 = imem05_in[71:68];
    24: op1_08_in10 = reg_0812;
    25: op1_08_in10 = reg_0651;
    26: op1_08_in10 = imem07_in[115:112];
    27: op1_08_in10 = reg_0214;
    54: op1_08_in10 = reg_0214;
    28: op1_08_in10 = reg_0371;
    29: op1_08_in10 = reg_0424;
    30: op1_08_in10 = reg_0212;
    31: op1_08_in10 = reg_0389;
    32: op1_08_in10 = reg_0087;
    33: op1_08_in10 = reg_0709;
    34: op1_08_in10 = imem03_in[119:116];
    35: op1_08_in10 = reg_0541;
    36: op1_08_in10 = reg_0545;
    85: op1_08_in10 = reg_0545;
    96: op1_08_in10 = reg_0545;
    37: op1_08_in10 = reg_0080;
    38: op1_08_in10 = reg_0145;
    39: op1_08_in10 = reg_0425;
    40: op1_08_in10 = imem07_in[79:76];
    41: op1_08_in10 = reg_0354;
    42: op1_08_in10 = reg_0007;
    43: op1_08_in10 = reg_0020;
    44: op1_08_in10 = reg_0213;
    45: op1_08_in10 = reg_0657;
    46: op1_08_in10 = reg_0304;
    47: op1_08_in10 = reg_0458;
    48: op1_08_in10 = imem02_in[111:108];
    49: op1_08_in10 = reg_0451;
    50: op1_08_in10 = reg_0172;
    51: op1_08_in10 = reg_0612;
    52: op1_08_in10 = reg_0708;
    55: op1_08_in10 = reg_0475;
    56: op1_08_in10 = imem02_in[63:60];
    57: op1_08_in10 = imem03_in[59:56];
    58: op1_08_in10 = reg_0341;
    59: op1_08_in10 = reg_0556;
    60: op1_08_in10 = imem04_in[87:84];
    61: op1_08_in10 = reg_0101;
    62: op1_08_in10 = reg_0481;
    63: op1_08_in10 = reg_0692;
    64: op1_08_in10 = imem02_in[103:100];
    65: op1_08_in10 = reg_0650;
    66: op1_08_in10 = reg_0483;
    67: op1_08_in10 = reg_0225;
    68: op1_08_in10 = reg_0724;
    69: op1_08_in10 = reg_0590;
    81: op1_08_in10 = reg_0590;
    70: op1_08_in10 = imem04_in[31:28];
    71: op1_08_in10 = reg_0247;
    72: op1_08_in10 = reg_0518;
    73: op1_08_in10 = reg_0344;
    74: op1_08_in10 = reg_0280;
    75: op1_08_in10 = reg_0583;
    76: op1_08_in10 = imem06_in[79:76];
    77: op1_08_in10 = reg_0183;
    79: op1_08_in10 = reg_0081;
    80: op1_08_in10 = imem04_in[59:56];
    82: op1_08_in10 = reg_0758;
    83: op1_08_in10 = reg_0156;
    84: op1_08_in10 = reg_0351;
    86: op1_08_in10 = imem07_in[123:120];
    87: op1_08_in10 = reg_0469;
    88: op1_08_in10 = reg_0439;
    89: op1_08_in10 = imem02_in[39:36];
    90: op1_08_in10 = reg_0603;
    91: op1_08_in10 = reg_0092;
    92: op1_08_in10 = reg_0149;
    93: op1_08_in10 = imem05_in[103:100];
    94: op1_08_in10 = imem05_in[55:52];
    95: op1_08_in10 = reg_0293;
    default: op1_08_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_08_inv10 = 1;
    12: op1_08_inv10 = 1;
    13: op1_08_inv10 = 1;
    14: op1_08_inv10 = 1;
    16: op1_08_inv10 = 1;
    17: op1_08_inv10 = 1;
    19: op1_08_inv10 = 1;
    20: op1_08_inv10 = 1;
    21: op1_08_inv10 = 1;
    24: op1_08_inv10 = 1;
    25: op1_08_inv10 = 1;
    27: op1_08_inv10 = 1;
    28: op1_08_inv10 = 1;
    30: op1_08_inv10 = 1;
    31: op1_08_inv10 = 1;
    32: op1_08_inv10 = 1;
    33: op1_08_inv10 = 1;
    35: op1_08_inv10 = 1;
    36: op1_08_inv10 = 1;
    38: op1_08_inv10 = 1;
    40: op1_08_inv10 = 1;
    41: op1_08_inv10 = 1;
    42: op1_08_inv10 = 1;
    44: op1_08_inv10 = 1;
    46: op1_08_inv10 = 1;
    52: op1_08_inv10 = 1;
    54: op1_08_inv10 = 1;
    55: op1_08_inv10 = 1;
    59: op1_08_inv10 = 1;
    65: op1_08_inv10 = 1;
    66: op1_08_inv10 = 1;
    69: op1_08_inv10 = 1;
    70: op1_08_inv10 = 1;
    71: op1_08_inv10 = 1;
    73: op1_08_inv10 = 1;
    77: op1_08_inv10 = 1;
    79: op1_08_inv10 = 1;
    82: op1_08_inv10 = 1;
    85: op1_08_inv10 = 1;
    86: op1_08_inv10 = 1;
    89: op1_08_inv10 = 1;
    92: op1_08_inv10 = 1;
    95: op1_08_inv10 = 1;
    96: op1_08_inv10 = 1;
    default: op1_08_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in11 = reg_0147;
    5: op1_08_in11 = reg_0545;
    6: op1_08_in11 = reg_0426;
    7: op1_08_in11 = reg_0645;
    8: op1_08_in11 = reg_0272;
    9: op1_08_in11 = reg_0800;
    10: op1_08_in11 = reg_0624;
    11: op1_08_in11 = reg_0593;
    12: op1_08_in11 = reg_0474;
    13: op1_08_in11 = reg_0118;
    14: op1_08_in11 = reg_0373;
    15: op1_08_in11 = reg_0705;
    16: op1_08_in11 = reg_0455;
    49: op1_08_in11 = reg_0455;
    17: op1_08_in11 = reg_0633;
    18: op1_08_in11 = reg_0471;
    19: op1_08_in11 = reg_0405;
    20: op1_08_in11 = reg_0687;
    21: op1_08_in11 = reg_0154;
    22: op1_08_in11 = reg_0309;
    23: op1_08_in11 = reg_0781;
    24: op1_08_in11 = reg_0813;
    25: op1_08_in11 = reg_0643;
    26: op1_08_in11 = reg_0716;
    86: op1_08_in11 = reg_0716;
    27: op1_08_in11 = imem01_in[3:0];
    28: op1_08_in11 = reg_0367;
    29: op1_08_in11 = reg_0447;
    30: op1_08_in11 = imem01_in[15:12];
    31: op1_08_in11 = reg_0570;
    32: op1_08_in11 = reg_0043;
    33: op1_08_in11 = reg_0715;
    34: op1_08_in11 = imem03_in[123:120];
    35: op1_08_in11 = reg_0081;
    72: op1_08_in11 = reg_0081;
    36: op1_08_in11 = reg_0315;
    37: op1_08_in11 = reg_0740;
    38: op1_08_in11 = reg_0136;
    39: op1_08_in11 = reg_0424;
    40: op1_08_in11 = imem07_in[123:120];
    41: op1_08_in11 = reg_0341;
    42: op1_08_in11 = reg_0014;
    43: op1_08_in11 = reg_0622;
    44: op1_08_in11 = reg_0202;
    55: op1_08_in11 = reg_0202;
    45: op1_08_in11 = reg_0639;
    66: op1_08_in11 = reg_0639;
    46: op1_08_in11 = reg_0279;
    47: op1_08_in11 = reg_0191;
    48: op1_08_in11 = reg_0658;
    50: op1_08_in11 = reg_0159;
    51: op1_08_in11 = reg_0402;
    52: op1_08_in11 = reg_0707;
    54: op1_08_in11 = reg_0209;
    56: op1_08_in11 = imem02_in[67:64];
    57: op1_08_in11 = imem03_in[103:100];
    58: op1_08_in11 = reg_0363;
    59: op1_08_in11 = reg_0283;
    60: op1_08_in11 = reg_0056;
    61: op1_08_in11 = reg_0285;
    62: op1_08_in11 = reg_0470;
    63: op1_08_in11 = reg_0472;
    64: op1_08_in11 = reg_0563;
    65: op1_08_in11 = reg_0045;
    67: op1_08_in11 = reg_0258;
    68: op1_08_in11 = reg_0709;
    69: op1_08_in11 = reg_0314;
    91: op1_08_in11 = reg_0314;
    70: op1_08_in11 = imem04_in[39:36];
    71: op1_08_in11 = reg_0692;
    78: op1_08_in11 = reg_0692;
    73: op1_08_in11 = reg_0356;
    74: op1_08_in11 = reg_0076;
    75: op1_08_in11 = reg_0025;
    76: op1_08_in11 = imem06_in[115:112];
    77: op1_08_in11 = reg_0168;
    79: op1_08_in11 = reg_0535;
    80: op1_08_in11 = imem04_in[111:108];
    81: op1_08_in11 = reg_0538;
    82: op1_08_in11 = reg_0688;
    83: op1_08_in11 = reg_0257;
    84: op1_08_in11 = reg_0365;
    85: op1_08_in11 = reg_0544;
    87: op1_08_in11 = reg_0475;
    88: op1_08_in11 = reg_0181;
    89: op1_08_in11 = reg_0533;
    90: op1_08_in11 = reg_0420;
    92: op1_08_in11 = reg_0785;
    93: op1_08_in11 = imem05_in[107:104];
    94: op1_08_in11 = reg_0736;
    95: op1_08_in11 = reg_0401;
    96: op1_08_in11 = reg_0060;
    default: op1_08_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv11 = 1;
    9: op1_08_inv11 = 1;
    10: op1_08_inv11 = 1;
    11: op1_08_inv11 = 1;
    12: op1_08_inv11 = 1;
    13: op1_08_inv11 = 1;
    14: op1_08_inv11 = 1;
    15: op1_08_inv11 = 1;
    16: op1_08_inv11 = 1;
    19: op1_08_inv11 = 1;
    20: op1_08_inv11 = 1;
    21: op1_08_inv11 = 1;
    22: op1_08_inv11 = 1;
    23: op1_08_inv11 = 1;
    24: op1_08_inv11 = 1;
    27: op1_08_inv11 = 1;
    29: op1_08_inv11 = 1;
    30: op1_08_inv11 = 1;
    33: op1_08_inv11 = 1;
    35: op1_08_inv11 = 1;
    37: op1_08_inv11 = 1;
    44: op1_08_inv11 = 1;
    46: op1_08_inv11 = 1;
    47: op1_08_inv11 = 1;
    50: op1_08_inv11 = 1;
    51: op1_08_inv11 = 1;
    52: op1_08_inv11 = 1;
    54: op1_08_inv11 = 1;
    58: op1_08_inv11 = 1;
    60: op1_08_inv11 = 1;
    63: op1_08_inv11 = 1;
    65: op1_08_inv11 = 1;
    66: op1_08_inv11 = 1;
    69: op1_08_inv11 = 1;
    76: op1_08_inv11 = 1;
    78: op1_08_inv11 = 1;
    79: op1_08_inv11 = 1;
    80: op1_08_inv11 = 1;
    81: op1_08_inv11 = 1;
    82: op1_08_inv11 = 1;
    83: op1_08_inv11 = 1;
    84: op1_08_inv11 = 1;
    85: op1_08_inv11 = 1;
    89: op1_08_inv11 = 1;
    91: op1_08_inv11 = 1;
    94: op1_08_inv11 = 1;
    95: op1_08_inv11 = 1;
    96: op1_08_inv11 = 1;
    default: op1_08_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in12 = reg_0148;
    5: op1_08_in12 = reg_0536;
    6: op1_08_in12 = reg_0172;
    7: op1_08_in12 = reg_0665;
    8: op1_08_in12 = reg_0261;
    9: op1_08_in12 = reg_0802;
    42: op1_08_in12 = reg_0802;
    10: op1_08_in12 = reg_0577;
    11: op1_08_in12 = reg_0311;
    12: op1_08_in12 = reg_0187;
    13: op1_08_in12 = reg_0112;
    14: op1_08_in12 = reg_0396;
    15: op1_08_in12 = reg_0701;
    52: op1_08_in12 = reg_0701;
    16: op1_08_in12 = reg_0461;
    49: op1_08_in12 = reg_0461;
    17: op1_08_in12 = reg_0623;
    18: op1_08_in12 = reg_0191;
    19: op1_08_in12 = reg_0386;
    20: op1_08_in12 = reg_0454;
    21: op1_08_in12 = imem06_in[3:0];
    22: op1_08_in12 = reg_0279;
    23: op1_08_in12 = reg_0488;
    24: op1_08_in12 = reg_0032;
    25: op1_08_in12 = reg_0652;
    26: op1_08_in12 = reg_0710;
    86: op1_08_in12 = reg_0710;
    27: op1_08_in12 = imem01_in[27:24];
    28: op1_08_in12 = reg_0610;
    29: op1_08_in12 = reg_0434;
    30: op1_08_in12 = imem01_in[23:20];
    31: op1_08_in12 = reg_0013;
    32: op1_08_in12 = reg_0088;
    33: op1_08_in12 = reg_0436;
    34: op1_08_in12 = reg_0582;
    35: op1_08_in12 = imem03_in[23:20];
    36: op1_08_in12 = reg_0558;
    37: op1_08_in12 = reg_0532;
    38: op1_08_in12 = reg_0128;
    39: op1_08_in12 = reg_0445;
    40: op1_08_in12 = reg_0704;
    41: op1_08_in12 = reg_0363;
    73: op1_08_in12 = reg_0363;
    43: op1_08_in12 = reg_0369;
    44: op1_08_in12 = imem01_in[15:12];
    45: op1_08_in12 = reg_0427;
    46: op1_08_in12 = reg_0224;
    47: op1_08_in12 = reg_0210;
    48: op1_08_in12 = reg_0666;
    51: op1_08_in12 = reg_0318;
    54: op1_08_in12 = reg_0186;
    55: op1_08_in12 = imem01_in[19:16];
    56: op1_08_in12 = imem02_in[87:84];
    57: op1_08_in12 = reg_0063;
    58: op1_08_in12 = reg_0342;
    59: op1_08_in12 = reg_0305;
    60: op1_08_in12 = reg_0555;
    61: op1_08_in12 = reg_0089;
    62: op1_08_in12 = reg_0474;
    63: op1_08_in12 = reg_0480;
    64: op1_08_in12 = reg_0483;
    65: op1_08_in12 = reg_0657;
    66: op1_08_in12 = reg_0355;
    67: op1_08_in12 = imem05_in[7:4];
    68: op1_08_in12 = reg_0706;
    69: op1_08_in12 = reg_0095;
    70: op1_08_in12 = imem04_in[59:56];
    71: op1_08_in12 = reg_0451;
    72: op1_08_in12 = reg_0538;
    74: op1_08_in12 = reg_0631;
    75: op1_08_in12 = reg_0700;
    76: op1_08_in12 = reg_0115;
    77: op1_08_in12 = reg_0184;
    78: op1_08_in12 = reg_0453;
    82: op1_08_in12 = reg_0453;
    79: op1_08_in12 = reg_0098;
    80: op1_08_in12 = reg_0545;
    81: op1_08_in12 = reg_0094;
    83: op1_08_in12 = reg_0765;
    84: op1_08_in12 = reg_0323;
    85: op1_08_in12 = reg_0173;
    87: op1_08_in12 = reg_0207;
    88: op1_08_in12 = reg_0142;
    89: op1_08_in12 = reg_0322;
    90: op1_08_in12 = reg_0105;
    91: op1_08_in12 = reg_0526;
    92: op1_08_in12 = reg_0156;
    93: op1_08_in12 = reg_0499;
    94: op1_08_in12 = reg_0133;
    95: op1_08_in12 = reg_0408;
    96: op1_08_in12 = reg_0554;
    default: op1_08_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv12 = 1;
    5: op1_08_inv12 = 1;
    6: op1_08_inv12 = 1;
    7: op1_08_inv12 = 1;
    8: op1_08_inv12 = 1;
    9: op1_08_inv12 = 1;
    10: op1_08_inv12 = 1;
    11: op1_08_inv12 = 1;
    13: op1_08_inv12 = 1;
    15: op1_08_inv12 = 1;
    18: op1_08_inv12 = 1;
    19: op1_08_inv12 = 1;
    27: op1_08_inv12 = 1;
    28: op1_08_inv12 = 1;
    30: op1_08_inv12 = 1;
    31: op1_08_inv12 = 1;
    32: op1_08_inv12 = 1;
    33: op1_08_inv12 = 1;
    34: op1_08_inv12 = 1;
    36: op1_08_inv12 = 1;
    46: op1_08_inv12 = 1;
    47: op1_08_inv12 = 1;
    49: op1_08_inv12 = 1;
    51: op1_08_inv12 = 1;
    52: op1_08_inv12 = 1;
    55: op1_08_inv12 = 1;
    56: op1_08_inv12 = 1;
    58: op1_08_inv12 = 1;
    60: op1_08_inv12 = 1;
    65: op1_08_inv12 = 1;
    67: op1_08_inv12 = 1;
    68: op1_08_inv12 = 1;
    71: op1_08_inv12 = 1;
    72: op1_08_inv12 = 1;
    75: op1_08_inv12 = 1;
    77: op1_08_inv12 = 1;
    78: op1_08_inv12 = 1;
    79: op1_08_inv12 = 1;
    80: op1_08_inv12 = 1;
    81: op1_08_inv12 = 1;
    83: op1_08_inv12 = 1;
    84: op1_08_inv12 = 1;
    85: op1_08_inv12 = 1;
    86: op1_08_inv12 = 1;
    88: op1_08_inv12 = 1;
    89: op1_08_inv12 = 1;
    94: op1_08_inv12 = 1;
    95: op1_08_inv12 = 1;
    default: op1_08_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in13 = reg_0149;
    5: op1_08_in13 = reg_0553;
    80: op1_08_in13 = reg_0553;
    6: op1_08_in13 = reg_0170;
    7: op1_08_in13 = reg_0659;
    8: op1_08_in13 = reg_0266;
    9: op1_08_in13 = reg_0010;
    10: op1_08_in13 = reg_0618;
    11: op1_08_in13 = reg_0319;
    12: op1_08_in13 = reg_0209;
    13: op1_08_in13 = reg_0121;
    14: op1_08_in13 = reg_0000;
    15: op1_08_in13 = reg_0700;
    16: op1_08_in13 = reg_0466;
    17: op1_08_in13 = reg_0612;
    18: op1_08_in13 = reg_0187;
    19: op1_08_in13 = reg_0390;
    20: op1_08_in13 = reg_0451;
    21: op1_08_in13 = imem06_in[27:24];
    22: op1_08_in13 = reg_0742;
    23: op1_08_in13 = reg_0780;
    24: op1_08_in13 = reg_0816;
    25: op1_08_in13 = imem02_in[3:0];
    84: op1_08_in13 = imem02_in[3:0];
    26: op1_08_in13 = reg_0723;
    27: op1_08_in13 = imem01_in[31:28];
    28: op1_08_in13 = reg_0611;
    74: op1_08_in13 = reg_0611;
    29: op1_08_in13 = reg_0444;
    30: op1_08_in13 = imem01_in[27:24];
    31: op1_08_in13 = reg_0804;
    32: op1_08_in13 = reg_0060;
    60: op1_08_in13 = reg_0060;
    33: op1_08_in13 = reg_0433;
    34: op1_08_in13 = reg_0591;
    35: op1_08_in13 = reg_0602;
    36: op1_08_in13 = reg_0551;
    37: op1_08_in13 = imem03_in[31:28];
    38: op1_08_in13 = reg_0156;
    39: op1_08_in13 = reg_0434;
    40: op1_08_in13 = reg_0726;
    41: op1_08_in13 = reg_0351;
    42: op1_08_in13 = imem04_in[27:24];
    43: op1_08_in13 = reg_0821;
    44: op1_08_in13 = imem01_in[35:32];
    45: op1_08_in13 = reg_0345;
    46: op1_08_in13 = reg_0307;
    47: op1_08_in13 = reg_0203;
    48: op1_08_in13 = reg_0637;
    49: op1_08_in13 = reg_0473;
    51: op1_08_in13 = reg_0404;
    52: op1_08_in13 = reg_0334;
    54: op1_08_in13 = imem01_in[15:12];
    55: op1_08_in13 = imem01_in[23:20];
    56: op1_08_in13 = imem02_in[119:116];
    57: op1_08_in13 = reg_0597;
    58: op1_08_in13 = reg_0527;
    59: op1_08_in13 = reg_0280;
    61: op1_08_in13 = reg_0132;
    62: op1_08_in13 = reg_0471;
    63: op1_08_in13 = reg_0467;
    64: op1_08_in13 = reg_0484;
    65: op1_08_in13 = reg_0237;
    66: op1_08_in13 = reg_0343;
    67: op1_08_in13 = imem05_in[51:48];
    68: op1_08_in13 = reg_0067;
    69: op1_08_in13 = reg_0097;
    70: op1_08_in13 = imem04_in[67:64];
    71: op1_08_in13 = reg_0457;
    72: op1_08_in13 = reg_0093;
    81: op1_08_in13 = reg_0093;
    73: op1_08_in13 = reg_0324;
    75: op1_08_in13 = reg_0767;
    76: op1_08_in13 = reg_0349;
    78: op1_08_in13 = reg_0477;
    79: op1_08_in13 = reg_0757;
    82: op1_08_in13 = reg_0462;
    83: op1_08_in13 = imem06_in[59:56];
    85: op1_08_in13 = reg_0534;
    86: op1_08_in13 = reg_0159;
    87: op1_08_in13 = reg_0211;
    88: op1_08_in13 = reg_0426;
    89: op1_08_in13 = reg_0359;
    90: op1_08_in13 = reg_0670;
    91: op1_08_in13 = imem03_in[15:12];
    92: op1_08_in13 = reg_0153;
    93: op1_08_in13 = reg_0134;
    94: op1_08_in13 = reg_0227;
    95: op1_08_in13 = reg_0246;
    96: op1_08_in13 = reg_0261;
    default: op1_08_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv13 = 1;
    5: op1_08_inv13 = 1;
    6: op1_08_inv13 = 1;
    8: op1_08_inv13 = 1;
    10: op1_08_inv13 = 1;
    11: op1_08_inv13 = 1;
    12: op1_08_inv13 = 1;
    13: op1_08_inv13 = 1;
    16: op1_08_inv13 = 1;
    17: op1_08_inv13 = 1;
    18: op1_08_inv13 = 1;
    20: op1_08_inv13 = 1;
    22: op1_08_inv13 = 1;
    23: op1_08_inv13 = 1;
    24: op1_08_inv13 = 1;
    28: op1_08_inv13 = 1;
    30: op1_08_inv13 = 1;
    32: op1_08_inv13 = 1;
    34: op1_08_inv13 = 1;
    35: op1_08_inv13 = 1;
    41: op1_08_inv13 = 1;
    43: op1_08_inv13 = 1;
    44: op1_08_inv13 = 1;
    47: op1_08_inv13 = 1;
    54: op1_08_inv13 = 1;
    59: op1_08_inv13 = 1;
    60: op1_08_inv13 = 1;
    64: op1_08_inv13 = 1;
    65: op1_08_inv13 = 1;
    66: op1_08_inv13 = 1;
    68: op1_08_inv13 = 1;
    70: op1_08_inv13 = 1;
    72: op1_08_inv13 = 1;
    74: op1_08_inv13 = 1;
    75: op1_08_inv13 = 1;
    78: op1_08_inv13 = 1;
    80: op1_08_inv13 = 1;
    82: op1_08_inv13 = 1;
    84: op1_08_inv13 = 1;
    86: op1_08_inv13 = 1;
    87: op1_08_inv13 = 1;
    88: op1_08_inv13 = 1;
    90: op1_08_inv13 = 1;
    92: op1_08_inv13 = 1;
    93: op1_08_inv13 = 1;
    94: op1_08_inv13 = 1;
    default: op1_08_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in14 = reg_0150;
    5: op1_08_in14 = reg_0303;
    7: op1_08_in14 = reg_0325;
    88: op1_08_in14 = reg_0325;
    8: op1_08_in14 = reg_0136;
    9: op1_08_in14 = reg_0004;
    10: op1_08_in14 = reg_0627;
    11: op1_08_in14 = reg_0369;
    12: op1_08_in14 = reg_0199;
    13: op1_08_in14 = imem02_in[23:20];
    14: op1_08_in14 = reg_0019;
    15: op1_08_in14 = reg_0424;
    16: op1_08_in14 = reg_0456;
    17: op1_08_in14 = reg_0402;
    18: op1_08_in14 = reg_0213;
    19: op1_08_in14 = reg_0401;
    20: op1_08_in14 = reg_0200;
    49: op1_08_in14 = reg_0200;
    21: op1_08_in14 = imem06_in[55:52];
    22: op1_08_in14 = reg_0276;
    23: op1_08_in14 = reg_0489;
    24: op1_08_in14 = reg_0750;
    25: op1_08_in14 = imem02_in[55:52];
    26: op1_08_in14 = reg_0717;
    40: op1_08_in14 = reg_0717;
    27: op1_08_in14 = imem01_in[119:116];
    28: op1_08_in14 = reg_0623;
    29: op1_08_in14 = reg_0420;
    30: op1_08_in14 = imem01_in[55:52];
    31: op1_08_in14 = reg_0801;
    32: op1_08_in14 = reg_0554;
    33: op1_08_in14 = reg_0428;
    34: op1_08_in14 = reg_0594;
    35: op1_08_in14 = reg_0596;
    36: op1_08_in14 = reg_0510;
    60: op1_08_in14 = reg_0510;
    37: op1_08_in14 = imem03_in[59:56];
    38: op1_08_in14 = reg_0130;
    39: op1_08_in14 = reg_0443;
    41: op1_08_in14 = reg_0322;
    42: op1_08_in14 = imem04_in[35:32];
    43: op1_08_in14 = reg_0270;
    44: op1_08_in14 = imem01_in[115:112];
    45: op1_08_in14 = reg_0365;
    46: op1_08_in14 = reg_0147;
    47: op1_08_in14 = reg_0196;
    48: op1_08_in14 = reg_0656;
    51: op1_08_in14 = reg_0329;
    52: op1_08_in14 = reg_0253;
    54: op1_08_in14 = imem01_in[35:32];
    55: op1_08_in14 = imem01_in[39:36];
    56: op1_08_in14 = imem02_in[127:124];
    57: op1_08_in14 = reg_0599;
    58: op1_08_in14 = reg_0095;
    59: op1_08_in14 = reg_0611;
    61: op1_08_in14 = reg_0135;
    62: op1_08_in14 = reg_0479;
    63: op1_08_in14 = reg_0471;
    64: op1_08_in14 = reg_0641;
    65: op1_08_in14 = reg_0358;
    66: op1_08_in14 = reg_0514;
    67: op1_08_in14 = imem05_in[79:76];
    68: op1_08_in14 = reg_0061;
    69: op1_08_in14 = reg_0082;
    70: op1_08_in14 = reg_0059;
    71: op1_08_in14 = reg_0476;
    72: op1_08_in14 = reg_0740;
    73: op1_08_in14 = reg_0406;
    74: op1_08_in14 = reg_0302;
    75: op1_08_in14 = reg_0752;
    76: op1_08_in14 = reg_0619;
    78: op1_08_in14 = reg_0473;
    79: op1_08_in14 = imem03_in[3:0];
    81: op1_08_in14 = imem03_in[3:0];
    80: op1_08_in14 = reg_0087;
    82: op1_08_in14 = reg_0191;
    83: op1_08_in14 = imem06_in[91:88];
    84: op1_08_in14 = imem02_in[11:8];
    85: op1_08_in14 = reg_0179;
    86: op1_08_in14 = reg_0726;
    87: op1_08_in14 = reg_0205;
    89: op1_08_in14 = reg_0565;
    90: op1_08_in14 = reg_0119;
    91: op1_08_in14 = imem03_in[47:44];
    92: op1_08_in14 = imem06_in[23:20];
    93: op1_08_in14 = reg_0517;
    94: op1_08_in14 = reg_0788;
    95: op1_08_in14 = reg_0215;
    96: op1_08_in14 = reg_0308;
    default: op1_08_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv14 = 1;
    5: op1_08_inv14 = 1;
    8: op1_08_inv14 = 1;
    10: op1_08_inv14 = 1;
    11: op1_08_inv14 = 1;
    13: op1_08_inv14 = 1;
    15: op1_08_inv14 = 1;
    17: op1_08_inv14 = 1;
    22: op1_08_inv14 = 1;
    23: op1_08_inv14 = 1;
    25: op1_08_inv14 = 1;
    26: op1_08_inv14 = 1;
    32: op1_08_inv14 = 1;
    35: op1_08_inv14 = 1;
    36: op1_08_inv14 = 1;
    37: op1_08_inv14 = 1;
    38: op1_08_inv14 = 1;
    41: op1_08_inv14 = 1;
    43: op1_08_inv14 = 1;
    45: op1_08_inv14 = 1;
    49: op1_08_inv14 = 1;
    52: op1_08_inv14 = 1;
    55: op1_08_inv14 = 1;
    58: op1_08_inv14 = 1;
    60: op1_08_inv14 = 1;
    62: op1_08_inv14 = 1;
    64: op1_08_inv14 = 1;
    70: op1_08_inv14 = 1;
    72: op1_08_inv14 = 1;
    76: op1_08_inv14 = 1;
    79: op1_08_inv14 = 1;
    81: op1_08_inv14 = 1;
    82: op1_08_inv14 = 1;
    83: op1_08_inv14 = 1;
    85: op1_08_inv14 = 1;
    86: op1_08_inv14 = 1;
    91: op1_08_inv14 = 1;
    default: op1_08_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in15 = reg_0129;
    5: op1_08_in15 = reg_0289;
    7: op1_08_in15 = reg_0324;
    8: op1_08_in15 = reg_0142;
    9: op1_08_in15 = imem04_in[11:8];
    10: op1_08_in15 = reg_0622;
    11: op1_08_in15 = reg_0309;
    12: op1_08_in15 = imem01_in[7:4];
    13: op1_08_in15 = imem02_in[39:36];
    14: op1_08_in15 = reg_0808;
    15: op1_08_in15 = reg_0434;
    16: op1_08_in15 = reg_0207;
    82: op1_08_in15 = reg_0207;
    17: op1_08_in15 = reg_0344;
    18: op1_08_in15 = reg_0212;
    19: op1_08_in15 = reg_0747;
    20: op1_08_in15 = reg_0203;
    21: op1_08_in15 = imem06_in[59:56];
    22: op1_08_in15 = reg_0148;
    23: op1_08_in15 = reg_0279;
    24: op1_08_in15 = imem07_in[11:8];
    25: op1_08_in15 = imem02_in[63:60];
    26: op1_08_in15 = reg_0724;
    27: op1_08_in15 = imem01_in[123:120];
    28: op1_08_in15 = imem06_in[31:28];
    29: op1_08_in15 = reg_0180;
    30: op1_08_in15 = reg_0501;
    31: op1_08_in15 = reg_0800;
    32: op1_08_in15 = reg_0057;
    33: op1_08_in15 = reg_0438;
    34: op1_08_in15 = reg_0585;
    35: op1_08_in15 = reg_0591;
    36: op1_08_in15 = reg_0053;
    37: op1_08_in15 = imem03_in[63:60];
    38: op1_08_in15 = reg_0051;
    39: op1_08_in15 = reg_0437;
    40: op1_08_in15 = reg_0714;
    41: op1_08_in15 = reg_0343;
    42: op1_08_in15 = imem04_in[67:64];
    43: op1_08_in15 = reg_0815;
    44: op1_08_in15 = imem01_in[127:124];
    45: op1_08_in15 = reg_0342;
    46: op1_08_in15 = reg_0133;
    47: op1_08_in15 = reg_0068;
    48: op1_08_in15 = reg_0639;
    49: op1_08_in15 = imem01_in[43:40];
    51: op1_08_in15 = reg_0401;
    52: op1_08_in15 = reg_0061;
    54: op1_08_in15 = imem01_in[47:44];
    55: op1_08_in15 = imem01_in[47:44];
    56: op1_08_in15 = reg_0655;
    57: op1_08_in15 = reg_0319;
    58: op1_08_in15 = reg_0540;
    59: op1_08_in15 = reg_0687;
    60: op1_08_in15 = reg_0280;
    61: op1_08_in15 = reg_0139;
    62: op1_08_in15 = reg_0208;
    63: op1_08_in15 = reg_0479;
    64: op1_08_in15 = reg_0372;
    65: op1_08_in15 = reg_0362;
    66: op1_08_in15 = reg_0092;
    67: op1_08_in15 = imem05_in[119:116];
    68: op1_08_in15 = reg_0439;
    69: op1_08_in15 = reg_0573;
    70: op1_08_in15 = reg_0560;
    71: op1_08_in15 = reg_0462;
    72: op1_08_in15 = imem03_in[7:4];
    73: op1_08_in15 = reg_0518;
    74: op1_08_in15 = reg_0616;
    75: op1_08_in15 = reg_0011;
    76: op1_08_in15 = reg_0638;
    78: op1_08_in15 = reg_0456;
    79: op1_08_in15 = imem03_in[99:96];
    80: op1_08_in15 = reg_0056;
    81: op1_08_in15 = imem03_in[15:12];
    83: op1_08_in15 = imem06_in[103:100];
    84: op1_08_in15 = imem02_in[19:16];
    85: op1_08_in15 = reg_0537;
    86: op1_08_in15 = reg_0158;
    87: op1_08_in15 = reg_0192;
    88: op1_08_in15 = reg_0091;
    89: op1_08_in15 = reg_0360;
    90: op1_08_in15 = reg_0601;
    91: op1_08_in15 = imem03_in[59:56];
    92: op1_08_in15 = imem06_in[55:52];
    93: op1_08_in15 = reg_0563;
    94: op1_08_in15 = reg_0550;
    95: op1_08_in15 = reg_0576;
    96: op1_08_in15 = reg_0631;
    default: op1_08_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv15 = 1;
    5: op1_08_inv15 = 1;
    9: op1_08_inv15 = 1;
    11: op1_08_inv15 = 1;
    14: op1_08_inv15 = 1;
    15: op1_08_inv15 = 1;
    16: op1_08_inv15 = 1;
    17: op1_08_inv15 = 1;
    21: op1_08_inv15 = 1;
    22: op1_08_inv15 = 1;
    27: op1_08_inv15 = 1;
    28: op1_08_inv15 = 1;
    34: op1_08_inv15 = 1;
    36: op1_08_inv15 = 1;
    38: op1_08_inv15 = 1;
    45: op1_08_inv15 = 1;
    47: op1_08_inv15 = 1;
    54: op1_08_inv15 = 1;
    55: op1_08_inv15 = 1;
    58: op1_08_inv15 = 1;
    63: op1_08_inv15 = 1;
    66: op1_08_inv15 = 1;
    69: op1_08_inv15 = 1;
    70: op1_08_inv15 = 1;
    72: op1_08_inv15 = 1;
    73: op1_08_inv15 = 1;
    74: op1_08_inv15 = 1;
    75: op1_08_inv15 = 1;
    79: op1_08_inv15 = 1;
    80: op1_08_inv15 = 1;
    82: op1_08_inv15 = 1;
    83: op1_08_inv15 = 1;
    84: op1_08_inv15 = 1;
    85: op1_08_inv15 = 1;
    86: op1_08_inv15 = 1;
    87: op1_08_inv15 = 1;
    88: op1_08_inv15 = 1;
    89: op1_08_inv15 = 1;
    92: op1_08_inv15 = 1;
    93: op1_08_inv15 = 1;
    default: op1_08_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in16 = imem06_in[11:8];
    61: op1_08_in16 = imem06_in[11:8];
    5: op1_08_in16 = reg_0054;
    7: op1_08_in16 = reg_0353;
    8: op1_08_in16 = reg_0143;
    9: op1_08_in16 = imem04_in[15:12];
    10: op1_08_in16 = reg_0381;
    11: op1_08_in16 = reg_0006;
    12: op1_08_in16 = imem01_in[15:12];
    13: op1_08_in16 = imem02_in[103:100];
    14: op1_08_in16 = reg_0013;
    15: op1_08_in16 = reg_0440;
    16: op1_08_in16 = reg_0186;
    17: op1_08_in16 = reg_0372;
    18: op1_08_in16 = reg_0199;
    19: op1_08_in16 = imem07_in[23:20];
    20: op1_08_in16 = reg_0194;
    21: op1_08_in16 = imem06_in[83:80];
    22: op1_08_in16 = reg_0133;
    23: op1_08_in16 = reg_0085;
    55: op1_08_in16 = reg_0085;
    24: op1_08_in16 = imem07_in[19:16];
    25: op1_08_in16 = imem02_in[119:116];
    26: op1_08_in16 = reg_0705;
    27: op1_08_in16 = reg_0520;
    28: op1_08_in16 = imem06_in[47:44];
    29: op1_08_in16 = reg_0165;
    39: op1_08_in16 = reg_0165;
    30: op1_08_in16 = reg_0824;
    31: op1_08_in16 = reg_0809;
    32: op1_08_in16 = reg_0283;
    33: op1_08_in16 = reg_0180;
    34: op1_08_in16 = reg_0595;
    35: op1_08_in16 = reg_0750;
    36: op1_08_in16 = reg_0265;
    37: op1_08_in16 = imem03_in[71:68];
    38: op1_08_in16 = reg_0629;
    40: op1_08_in16 = reg_0703;
    41: op1_08_in16 = reg_0321;
    45: op1_08_in16 = reg_0321;
    42: op1_08_in16 = imem04_in[79:76];
    43: op1_08_in16 = reg_0231;
    44: op1_08_in16 = reg_0758;
    46: op1_08_in16 = reg_0156;
    47: op1_08_in16 = reg_0069;
    59: op1_08_in16 = reg_0069;
    48: op1_08_in16 = reg_0349;
    49: op1_08_in16 = imem01_in[47:44];
    51: op1_08_in16 = reg_0812;
    52: op1_08_in16 = reg_0333;
    54: op1_08_in16 = imem01_in[119:116];
    56: op1_08_in16 = reg_0661;
    57: op1_08_in16 = reg_0561;
    58: op1_08_in16 = imem03_in[7:4];
    60: op1_08_in16 = reg_0611;
    62: op1_08_in16 = reg_0191;
    63: op1_08_in16 = reg_0209;
    64: op1_08_in16 = reg_0344;
    65: op1_08_in16 = reg_0363;
    66: op1_08_in16 = reg_0540;
    67: op1_08_in16 = imem05_in[127:124];
    68: op1_08_in16 = reg_0435;
    69: op1_08_in16 = reg_0735;
    70: op1_08_in16 = reg_0055;
    71: op1_08_in16 = reg_0471;
    72: op1_08_in16 = imem03_in[11:8];
    73: op1_08_in16 = reg_0095;
    74: op1_08_in16 = reg_0626;
    75: op1_08_in16 = imem07_in[79:76];
    76: op1_08_in16 = reg_0218;
    78: op1_08_in16 = reg_0478;
    79: op1_08_in16 = reg_0596;
    80: op1_08_in16 = reg_0523;
    81: op1_08_in16 = imem03_in[27:24];
    82: op1_08_in16 = reg_0198;
    83: op1_08_in16 = imem06_in[115:112];
    84: op1_08_in16 = imem02_in[27:24];
    85: op1_08_in16 = reg_0554;
    86: op1_08_in16 = reg_0334;
    87: op1_08_in16 = imem01_in[11:8];
    88: op1_08_in16 = reg_0184;
    89: op1_08_in16 = reg_0324;
    90: op1_08_in16 = reg_0107;
    91: op1_08_in16 = imem03_in[119:116];
    92: op1_08_in16 = imem06_in[91:88];
    93: op1_08_in16 = reg_0245;
    94: op1_08_in16 = reg_0793;
    95: op1_08_in16 = reg_0657;
    96: op1_08_in16 = reg_0301;
    default: op1_08_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv16 = 1;
    7: op1_08_inv16 = 1;
    8: op1_08_inv16 = 1;
    9: op1_08_inv16 = 1;
    10: op1_08_inv16 = 1;
    14: op1_08_inv16 = 1;
    17: op1_08_inv16 = 1;
    18: op1_08_inv16 = 1;
    19: op1_08_inv16 = 1;
    21: op1_08_inv16 = 1;
    24: op1_08_inv16 = 1;
    28: op1_08_inv16 = 1;
    29: op1_08_inv16 = 1;
    30: op1_08_inv16 = 1;
    31: op1_08_inv16 = 1;
    33: op1_08_inv16 = 1;
    34: op1_08_inv16 = 1;
    35: op1_08_inv16 = 1;
    37: op1_08_inv16 = 1;
    40: op1_08_inv16 = 1;
    44: op1_08_inv16 = 1;
    45: op1_08_inv16 = 1;
    46: op1_08_inv16 = 1;
    49: op1_08_inv16 = 1;
    51: op1_08_inv16 = 1;
    55: op1_08_inv16 = 1;
    56: op1_08_inv16 = 1;
    57: op1_08_inv16 = 1;
    59: op1_08_inv16 = 1;
    60: op1_08_inv16 = 1;
    61: op1_08_inv16 = 1;
    62: op1_08_inv16 = 1;
    65: op1_08_inv16 = 1;
    66: op1_08_inv16 = 1;
    67: op1_08_inv16 = 1;
    68: op1_08_inv16 = 1;
    70: op1_08_inv16 = 1;
    74: op1_08_inv16 = 1;
    78: op1_08_inv16 = 1;
    79: op1_08_inv16 = 1;
    82: op1_08_inv16 = 1;
    86: op1_08_inv16 = 1;
    87: op1_08_inv16 = 1;
    88: op1_08_inv16 = 1;
    89: op1_08_inv16 = 1;
    90: op1_08_inv16 = 1;
    91: op1_08_inv16 = 1;
    92: op1_08_inv16 = 1;
    94: op1_08_inv16 = 1;
    default: op1_08_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in17 = reg_0607;
    5: op1_08_in17 = reg_0043;
    7: op1_08_in17 = reg_0310;
    8: op1_08_in17 = reg_0130;
    9: op1_08_in17 = imem04_in[71:68];
    10: op1_08_in17 = reg_0367;
    11: op1_08_in17 = reg_0803;
    12: op1_08_in17 = imem01_in[55:52];
    13: op1_08_in17 = imem02_in[107:104];
    14: op1_08_in17 = reg_0007;
    15: op1_08_in17 = reg_0427;
    16: op1_08_in17 = reg_0198;
    17: op1_08_in17 = reg_0407;
    18: op1_08_in17 = imem01_in[7:4];
    19: op1_08_in17 = imem07_in[75:72];
    20: op1_08_in17 = imem01_in[11:8];
    21: op1_08_in17 = imem06_in[95:92];
    22: op1_08_in17 = reg_0150;
    23: op1_08_in17 = reg_0307;
    24: op1_08_in17 = imem07_in[43:40];
    43: op1_08_in17 = imem07_in[43:40];
    25: op1_08_in17 = reg_0314;
    26: op1_08_in17 = reg_0711;
    27: op1_08_in17 = reg_0514;
    28: op1_08_in17 = imem06_in[51:48];
    29: op1_08_in17 = reg_0177;
    39: op1_08_in17 = reg_0177;
    30: op1_08_in17 = reg_0227;
    31: op1_08_in17 = imem04_in[31:28];
    32: op1_08_in17 = reg_0529;
    33: op1_08_in17 = reg_0172;
    34: op1_08_in17 = reg_0394;
    35: op1_08_in17 = reg_0584;
    36: op1_08_in17 = reg_0291;
    37: op1_08_in17 = imem03_in[87:84];
    38: op1_08_in17 = reg_0617;
    40: op1_08_in17 = reg_0708;
    41: op1_08_in17 = reg_0323;
    42: op1_08_in17 = imem04_in[127:124];
    44: op1_08_in17 = reg_0501;
    45: op1_08_in17 = reg_0541;
    46: op1_08_in17 = reg_0143;
    47: op1_08_in17 = reg_0075;
    48: op1_08_in17 = reg_0345;
    49: op1_08_in17 = imem01_in[51:48];
    51: op1_08_in17 = reg_0621;
    52: op1_08_in17 = reg_0180;
    54: op1_08_in17 = reg_0085;
    55: op1_08_in17 = reg_0322;
    56: op1_08_in17 = reg_0638;
    57: op1_08_in17 = reg_0562;
    58: op1_08_in17 = imem03_in[39:36];
    59: op1_08_in17 = reg_0640;
    60: op1_08_in17 = reg_0077;
    61: op1_08_in17 = reg_0817;
    62: op1_08_in17 = reg_0207;
    63: op1_08_in17 = reg_0190;
    64: op1_08_in17 = reg_0341;
    65: op1_08_in17 = reg_0533;
    66: op1_08_in17 = reg_0526;
    67: op1_08_in17 = reg_0246;
    68: op1_08_in17 = reg_0174;
    69: op1_08_in17 = reg_0039;
    70: op1_08_in17 = reg_0554;
    71: op1_08_in17 = reg_0479;
    72: op1_08_in17 = imem03_in[27:24];
    73: op1_08_in17 = reg_0769;
    74: op1_08_in17 = reg_0301;
    75: op1_08_in17 = imem07_in[91:88];
    76: op1_08_in17 = imem07_in[31:28];
    78: op1_08_in17 = reg_0458;
    79: op1_08_in17 = reg_0751;
    80: op1_08_in17 = reg_0305;
    81: op1_08_in17 = imem03_in[31:28];
    82: op1_08_in17 = reg_0201;
    83: op1_08_in17 = reg_0299;
    84: op1_08_in17 = imem02_in[103:100];
    85: op1_08_in17 = reg_0536;
    86: op1_08_in17 = reg_0266;
    87: op1_08_in17 = imem01_in[87:84];
    89: op1_08_in17 = reg_0406;
    90: op1_08_in17 = imem02_in[55:52];
    91: op1_08_in17 = imem03_in[123:120];
    92: op1_08_in17 = reg_0348;
    93: op1_08_in17 = reg_0531;
    94: op1_08_in17 = reg_0231;
    95: op1_08_in17 = imem07_in[51:48];
    96: op1_08_in17 = reg_0780;
    default: op1_08_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_08_inv17 = 1;
    9: op1_08_inv17 = 1;
    12: op1_08_inv17 = 1;
    14: op1_08_inv17 = 1;
    16: op1_08_inv17 = 1;
    18: op1_08_inv17 = 1;
    19: op1_08_inv17 = 1;
    20: op1_08_inv17 = 1;
    22: op1_08_inv17 = 1;
    23: op1_08_inv17 = 1;
    25: op1_08_inv17 = 1;
    28: op1_08_inv17 = 1;
    29: op1_08_inv17 = 1;
    31: op1_08_inv17 = 1;
    32: op1_08_inv17 = 1;
    34: op1_08_inv17 = 1;
    35: op1_08_inv17 = 1;
    37: op1_08_inv17 = 1;
    38: op1_08_inv17 = 1;
    40: op1_08_inv17 = 1;
    44: op1_08_inv17 = 1;
    45: op1_08_inv17 = 1;
    46: op1_08_inv17 = 1;
    47: op1_08_inv17 = 1;
    52: op1_08_inv17 = 1;
    54: op1_08_inv17 = 1;
    56: op1_08_inv17 = 1;
    58: op1_08_inv17 = 1;
    61: op1_08_inv17 = 1;
    62: op1_08_inv17 = 1;
    64: op1_08_inv17 = 1;
    69: op1_08_inv17 = 1;
    72: op1_08_inv17 = 1;
    73: op1_08_inv17 = 1;
    74: op1_08_inv17 = 1;
    79: op1_08_inv17 = 1;
    80: op1_08_inv17 = 1;
    84: op1_08_inv17 = 1;
    86: op1_08_inv17 = 1;
    87: op1_08_inv17 = 1;
    92: op1_08_inv17 = 1;
    93: op1_08_inv17 = 1;
    94: op1_08_inv17 = 1;
    default: op1_08_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in18 = reg_0616;
    38: op1_08_in18 = reg_0616;
    5: op1_08_in18 = reg_0063;
    69: op1_08_in18 = reg_0063;
    7: op1_08_in18 = reg_0350;
    8: op1_08_in18 = reg_0155;
    9: op1_08_in18 = imem04_in[79:76];
    31: op1_08_in18 = imem04_in[79:76];
    10: op1_08_in18 = reg_0337;
    11: op1_08_in18 = reg_0007;
    12: op1_08_in18 = imem01_in[87:84];
    13: op1_08_in18 = imem02_in[123:120];
    14: op1_08_in18 = reg_0015;
    15: op1_08_in18 = reg_0435;
    16: op1_08_in18 = reg_0213;
    17: op1_08_in18 = reg_0383;
    34: op1_08_in18 = reg_0383;
    18: op1_08_in18 = imem01_in[11:8];
    62: op1_08_in18 = imem01_in[11:8];
    19: op1_08_in18 = reg_0719;
    20: op1_08_in18 = imem01_in[43:40];
    21: op1_08_in18 = imem06_in[103:100];
    22: op1_08_in18 = reg_0144;
    23: op1_08_in18 = reg_0089;
    24: op1_08_in18 = imem07_in[51:48];
    43: op1_08_in18 = imem07_in[51:48];
    25: op1_08_in18 = reg_0082;
    26: op1_08_in18 = reg_0433;
    27: op1_08_in18 = reg_0227;
    28: op1_08_in18 = imem06_in[67:64];
    30: op1_08_in18 = reg_0232;
    32: op1_08_in18 = reg_0268;
    36: op1_08_in18 = reg_0268;
    33: op1_08_in18 = reg_0177;
    35: op1_08_in18 = reg_0578;
    37: op1_08_in18 = imem03_in[91:88];
    39: op1_08_in18 = reg_0184;
    40: op1_08_in18 = reg_0727;
    41: op1_08_in18 = reg_0080;
    42: op1_08_in18 = reg_0328;
    44: op1_08_in18 = reg_0496;
    45: op1_08_in18 = reg_0533;
    90: op1_08_in18 = reg_0533;
    46: op1_08_in18 = reg_0139;
    47: op1_08_in18 = imem01_in[27:24];
    48: op1_08_in18 = reg_0365;
    49: op1_08_in18 = imem01_in[91:88];
    51: op1_08_in18 = imem07_in[19:16];
    52: op1_08_in18 = reg_0181;
    54: op1_08_in18 = reg_0100;
    55: op1_08_in18 = reg_0054;
    56: op1_08_in18 = reg_0362;
    57: op1_08_in18 = reg_0376;
    58: op1_08_in18 = imem03_in[55:52];
    72: op1_08_in18 = imem03_in[55:52];
    59: op1_08_in18 = reg_0109;
    60: op1_08_in18 = reg_0626;
    61: op1_08_in18 = reg_0618;
    63: op1_08_in18 = reg_0199;
    64: op1_08_in18 = reg_0565;
    65: op1_08_in18 = reg_0535;
    66: op1_08_in18 = imem03_in[43:40];
    67: op1_08_in18 = reg_0491;
    68: op1_08_in18 = reg_0162;
    70: op1_08_in18 = reg_0510;
    71: op1_08_in18 = reg_0191;
    73: op1_08_in18 = reg_0770;
    74: op1_08_in18 = reg_0311;
    75: op1_08_in18 = imem07_in[95:92];
    76: op1_08_in18 = imem07_in[47:44];
    78: op1_08_in18 = reg_0189;
    79: op1_08_in18 = reg_0509;
    80: op1_08_in18 = reg_0631;
    81: op1_08_in18 = imem03_in[51:48];
    82: op1_08_in18 = reg_0212;
    83: op1_08_in18 = reg_0625;
    84: op1_08_in18 = imem02_in[111:108];
    85: op1_08_in18 = reg_0308;
    86: op1_08_in18 = reg_0333;
    87: op1_08_in18 = reg_0653;
    89: op1_08_in18 = reg_0092;
    91: op1_08_in18 = reg_0604;
    92: op1_08_in18 = reg_0346;
    93: op1_08_in18 = reg_0785;
    94: op1_08_in18 = reg_0355;
    95: op1_08_in18 = imem07_in[67:64];
    96: op1_08_in18 = reg_0643;
    default: op1_08_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv18 = 1;
    11: op1_08_inv18 = 1;
    15: op1_08_inv18 = 1;
    18: op1_08_inv18 = 1;
    23: op1_08_inv18 = 1;
    25: op1_08_inv18 = 1;
    26: op1_08_inv18 = 1;
    28: op1_08_inv18 = 1;
    30: op1_08_inv18 = 1;
    31: op1_08_inv18 = 1;
    33: op1_08_inv18 = 1;
    35: op1_08_inv18 = 1;
    42: op1_08_inv18 = 1;
    43: op1_08_inv18 = 1;
    49: op1_08_inv18 = 1;
    52: op1_08_inv18 = 1;
    54: op1_08_inv18 = 1;
    55: op1_08_inv18 = 1;
    57: op1_08_inv18 = 1;
    59: op1_08_inv18 = 1;
    60: op1_08_inv18 = 1;
    61: op1_08_inv18 = 1;
    63: op1_08_inv18 = 1;
    64: op1_08_inv18 = 1;
    66: op1_08_inv18 = 1;
    78: op1_08_inv18 = 1;
    80: op1_08_inv18 = 1;
    82: op1_08_inv18 = 1;
    83: op1_08_inv18 = 1;
    84: op1_08_inv18 = 1;
    85: op1_08_inv18 = 1;
    89: op1_08_inv18 = 1;
    91: op1_08_inv18 = 1;
    92: op1_08_inv18 = 1;
    93: op1_08_inv18 = 1;
    94: op1_08_inv18 = 1;
    default: op1_08_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in19 = reg_0609;
    5: op1_08_in19 = reg_0072;
    7: op1_08_in19 = reg_0080;
    8: op1_08_in19 = reg_0137;
    9: op1_08_in19 = imem04_in[87:84];
    10: op1_08_in19 = reg_0815;
    11: op1_08_in19 = reg_0800;
    12: op1_08_in19 = imem01_in[91:88];
    13: op1_08_in19 = reg_0666;
    14: op1_08_in19 = reg_0809;
    15: op1_08_in19 = reg_0159;
    16: op1_08_in19 = reg_0205;
    17: op1_08_in19 = reg_0033;
    18: op1_08_in19 = imem01_in[15:12];
    63: op1_08_in19 = imem01_in[15:12];
    19: op1_08_in19 = reg_0723;
    20: op1_08_in19 = imem01_in[51:48];
    21: op1_08_in19 = reg_0630;
    22: op1_08_in19 = imem06_in[19:16];
    23: op1_08_in19 = reg_0135;
    24: op1_08_in19 = imem07_in[63:60];
    43: op1_08_in19 = imem07_in[63:60];
    25: op1_08_in19 = reg_0757;
    26: op1_08_in19 = reg_0442;
    27: op1_08_in19 = reg_0333;
    28: op1_08_in19 = imem06_in[83:80];
    30: op1_08_in19 = reg_0505;
    31: op1_08_in19 = imem04_in[99:96];
    32: op1_08_in19 = reg_0050;
    33: op1_08_in19 = reg_0164;
    34: op1_08_in19 = reg_0569;
    35: op1_08_in19 = reg_0395;
    36: op1_08_in19 = reg_0297;
    37: op1_08_in19 = reg_0587;
    38: op1_08_in19 = reg_0041;
    40: op1_08_in19 = reg_0430;
    41: op1_08_in19 = reg_0096;
    42: op1_08_in19 = reg_0058;
    44: op1_08_in19 = reg_0513;
    45: op1_08_in19 = reg_0538;
    46: op1_08_in19 = reg_0140;
    47: op1_08_in19 = imem01_in[47:44];
    48: op1_08_in19 = reg_0518;
    49: op1_08_in19 = imem01_in[99:96];
    51: op1_08_in19 = imem07_in[47:44];
    52: op1_08_in19 = reg_0179;
    54: op1_08_in19 = reg_0778;
    55: op1_08_in19 = reg_0217;
    56: op1_08_in19 = reg_0324;
    57: op1_08_in19 = reg_0393;
    58: op1_08_in19 = imem03_in[79:76];
    59: op1_08_in19 = imem05_in[11:8];
    60: op1_08_in19 = reg_0301;
    61: op1_08_in19 = reg_0519;
    62: op1_08_in19 = imem01_in[19:16];
    64: op1_08_in19 = reg_0351;
    65: op1_08_in19 = reg_0539;
    66: op1_08_in19 = imem03_in[71:68];
    67: op1_08_in19 = reg_0040;
    68: op1_08_in19 = reg_0160;
    69: op1_08_in19 = reg_0347;
    70: op1_08_in19 = reg_0516;
    71: op1_08_in19 = reg_0189;
    72: op1_08_in19 = imem03_in[107:104];
    73: op1_08_in19 = reg_0531;
    74: op1_08_in19 = reg_0371;
    75: op1_08_in19 = reg_0719;
    76: op1_08_in19 = imem07_in[55:52];
    78: op1_08_in19 = reg_0188;
    79: op1_08_in19 = reg_0648;
    80: op1_08_in19 = reg_0077;
    81: op1_08_in19 = imem03_in[55:52];
    82: op1_08_in19 = imem01_in[7:4];
    83: op1_08_in19 = reg_0346;
    84: op1_08_in19 = imem03_in[3:0];
    85: op1_08_in19 = reg_0429;
    86: op1_08_in19 = reg_0438;
    87: op1_08_in19 = reg_0385;
    89: op1_08_in19 = reg_0109;
    90: op1_08_in19 = reg_0081;
    91: op1_08_in19 = reg_0494;
    92: op1_08_in19 = reg_0349;
    93: op1_08_in19 = reg_0154;
    94: op1_08_in19 = reg_0489;
    95: op1_08_in19 = reg_0391;
    96: op1_08_in19 = imem05_in[19:16];
    default: op1_08_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv19 = 1;
    7: op1_08_inv19 = 1;
    8: op1_08_inv19 = 1;
    12: op1_08_inv19 = 1;
    13: op1_08_inv19 = 1;
    14: op1_08_inv19 = 1;
    16: op1_08_inv19 = 1;
    19: op1_08_inv19 = 1;
    21: op1_08_inv19 = 1;
    22: op1_08_inv19 = 1;
    24: op1_08_inv19 = 1;
    25: op1_08_inv19 = 1;
    26: op1_08_inv19 = 1;
    30: op1_08_inv19 = 1;
    31: op1_08_inv19 = 1;
    32: op1_08_inv19 = 1;
    34: op1_08_inv19 = 1;
    35: op1_08_inv19 = 1;
    37: op1_08_inv19 = 1;
    38: op1_08_inv19 = 1;
    40: op1_08_inv19 = 1;
    41: op1_08_inv19 = 1;
    42: op1_08_inv19 = 1;
    43: op1_08_inv19 = 1;
    45: op1_08_inv19 = 1;
    46: op1_08_inv19 = 1;
    51: op1_08_inv19 = 1;
    52: op1_08_inv19 = 1;
    58: op1_08_inv19 = 1;
    59: op1_08_inv19 = 1;
    60: op1_08_inv19 = 1;
    62: op1_08_inv19 = 1;
    63: op1_08_inv19 = 1;
    66: op1_08_inv19 = 1;
    67: op1_08_inv19 = 1;
    68: op1_08_inv19 = 1;
    69: op1_08_inv19 = 1;
    70: op1_08_inv19 = 1;
    72: op1_08_inv19 = 1;
    73: op1_08_inv19 = 1;
    74: op1_08_inv19 = 1;
    75: op1_08_inv19 = 1;
    76: op1_08_inv19 = 1;
    78: op1_08_inv19 = 1;
    81: op1_08_inv19 = 1;
    82: op1_08_inv19 = 1;
    87: op1_08_inv19 = 1;
    89: op1_08_inv19 = 1;
    90: op1_08_inv19 = 1;
    91: op1_08_inv19 = 1;
    92: op1_08_inv19 = 1;
    93: op1_08_inv19 = 1;
    95: op1_08_inv19 = 1;
    default: op1_08_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in20 = reg_0402;
    5: op1_08_in20 = reg_0742;
    7: op1_08_in20 = reg_0090;
    8: op1_08_in20 = reg_0131;
    9: op1_08_in20 = imem04_in[91:88];
    10: op1_08_in20 = reg_0819;
    11: op1_08_in20 = reg_0004;
    12: op1_08_in20 = reg_0512;
    13: op1_08_in20 = reg_0639;
    14: op1_08_in20 = imem04_in[35:32];
    15: op1_08_in20 = reg_0182;
    16: op1_08_in20 = reg_0197;
    17: op1_08_in20 = reg_0812;
    18: op1_08_in20 = imem01_in[23:20];
    19: op1_08_in20 = reg_0712;
    20: op1_08_in20 = imem01_in[55:52];
    47: op1_08_in20 = imem01_in[55:52];
    21: op1_08_in20 = reg_0605;
    22: op1_08_in20 = imem06_in[31:28];
    38: op1_08_in20 = imem06_in[31:28];
    23: op1_08_in20 = reg_0152;
    24: op1_08_in20 = imem07_in[67:64];
    76: op1_08_in20 = imem07_in[67:64];
    25: op1_08_in20 = imem03_in[15:12];
    26: op1_08_in20 = reg_0443;
    27: op1_08_in20 = reg_0515;
    28: op1_08_in20 = imem06_in[87:84];
    30: op1_08_in20 = reg_0246;
    31: op1_08_in20 = imem04_in[111:108];
    32: op1_08_in20 = reg_0257;
    33: op1_08_in20 = reg_0171;
    34: op1_08_in20 = reg_0398;
    35: op1_08_in20 = reg_0575;
    36: op1_08_in20 = reg_0295;
    37: op1_08_in20 = reg_0750;
    40: op1_08_in20 = reg_0433;
    85: op1_08_in20 = reg_0433;
    41: op1_08_in20 = reg_0540;
    89: op1_08_in20 = reg_0540;
    42: op1_08_in20 = reg_0547;
    43: op1_08_in20 = imem07_in[87:84];
    44: op1_08_in20 = reg_0822;
    45: op1_08_in20 = imem03_in[63:60];
    46: op1_08_in20 = imem06_in[19:16];
    48: op1_08_in20 = reg_0541;
    49: op1_08_in20 = imem01_in[103:100];
    51: op1_08_in20 = imem07_in[51:48];
    52: op1_08_in20 = reg_0177;
    54: op1_08_in20 = reg_0321;
    55: op1_08_in20 = reg_0502;
    56: op1_08_in20 = reg_0365;
    57: op1_08_in20 = reg_0389;
    58: op1_08_in20 = imem03_in[91:88];
    59: op1_08_in20 = imem05_in[55:52];
    60: op1_08_in20 = reg_0078;
    61: op1_08_in20 = reg_0630;
    62: op1_08_in20 = imem01_in[39:36];
    63: op1_08_in20 = imem01_in[27:24];
    64: op1_08_in20 = reg_0590;
    65: op1_08_in20 = reg_0757;
    66: op1_08_in20 = imem03_in[87:84];
    67: op1_08_in20 = reg_0288;
    68: op1_08_in20 = reg_0166;
    69: op1_08_in20 = reg_0493;
    70: op1_08_in20 = reg_0432;
    71: op1_08_in20 = reg_0187;
    72: op1_08_in20 = imem03_in[119:116];
    73: op1_08_in20 = imem03_in[27:24];
    74: op1_08_in20 = imem05_in[15:12];
    75: op1_08_in20 = reg_0723;
    78: op1_08_in20 = imem01_in[15:12];
    79: op1_08_in20 = reg_0384;
    80: op1_08_in20 = reg_0065;
    81: op1_08_in20 = imem03_in[71:68];
    82: op1_08_in20 = imem01_in[87:84];
    83: op1_08_in20 = reg_0291;
    84: op1_08_in20 = imem03_in[7:4];
    86: op1_08_in20 = reg_0236;
    87: op1_08_in20 = reg_0101;
    90: op1_08_in20 = reg_0080;
    91: op1_08_in20 = reg_0318;
    92: op1_08_in20 = reg_0339;
    93: op1_08_in20 = reg_0137;
    94: op1_08_in20 = reg_0386;
    95: op1_08_in20 = reg_0725;
    96: op1_08_in20 = imem05_in[39:36];
    default: op1_08_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_08_inv20 = 1;
    11: op1_08_inv20 = 1;
    12: op1_08_inv20 = 1;
    14: op1_08_inv20 = 1;
    17: op1_08_inv20 = 1;
    18: op1_08_inv20 = 1;
    24: op1_08_inv20 = 1;
    26: op1_08_inv20 = 1;
    27: op1_08_inv20 = 1;
    30: op1_08_inv20 = 1;
    31: op1_08_inv20 = 1;
    32: op1_08_inv20 = 1;
    33: op1_08_inv20 = 1;
    34: op1_08_inv20 = 1;
    37: op1_08_inv20 = 1;
    40: op1_08_inv20 = 1;
    42: op1_08_inv20 = 1;
    43: op1_08_inv20 = 1;
    44: op1_08_inv20 = 1;
    45: op1_08_inv20 = 1;
    49: op1_08_inv20 = 1;
    52: op1_08_inv20 = 1;
    54: op1_08_inv20 = 1;
    56: op1_08_inv20 = 1;
    57: op1_08_inv20 = 1;
    58: op1_08_inv20 = 1;
    59: op1_08_inv20 = 1;
    60: op1_08_inv20 = 1;
    61: op1_08_inv20 = 1;
    63: op1_08_inv20 = 1;
    64: op1_08_inv20 = 1;
    66: op1_08_inv20 = 1;
    70: op1_08_inv20 = 1;
    74: op1_08_inv20 = 1;
    76: op1_08_inv20 = 1;
    79: op1_08_inv20 = 1;
    80: op1_08_inv20 = 1;
    85: op1_08_inv20 = 1;
    86: op1_08_inv20 = 1;
    89: op1_08_inv20 = 1;
    90: op1_08_inv20 = 1;
    91: op1_08_inv20 = 1;
    92: op1_08_inv20 = 1;
    93: op1_08_inv20 = 1;
    94: op1_08_inv20 = 1;
    95: op1_08_inv20 = 1;
    96: op1_08_inv20 = 1;
    default: op1_08_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in21 = reg_0348;
    5: op1_08_in21 = reg_0737;
    7: op1_08_in21 = reg_0055;
    8: op1_08_in21 = reg_0134;
    9: op1_08_in21 = imem04_in[107:104];
    10: op1_08_in21 = reg_0818;
    11: op1_08_in21 = imem04_in[7:4];
    12: op1_08_in21 = reg_0514;
    13: op1_08_in21 = reg_0649;
    14: op1_08_in21 = imem04_in[55:52];
    15: op1_08_in21 = reg_0177;
    16: op1_08_in21 = imem01_in[83:80];
    62: op1_08_in21 = imem01_in[83:80];
    78: op1_08_in21 = imem01_in[83:80];
    17: op1_08_in21 = reg_0815;
    18: op1_08_in21 = imem01_in[31:28];
    19: op1_08_in21 = reg_0709;
    20: op1_08_in21 = imem01_in[67:64];
    21: op1_08_in21 = reg_0626;
    22: op1_08_in21 = imem06_in[35:32];
    93: op1_08_in21 = imem06_in[35:32];
    23: op1_08_in21 = reg_0156;
    24: op1_08_in21 = imem07_in[91:88];
    43: op1_08_in21 = imem07_in[91:88];
    25: op1_08_in21 = imem03_in[39:36];
    73: op1_08_in21 = imem03_in[39:36];
    26: op1_08_in21 = reg_0431;
    27: op1_08_in21 = reg_0760;
    28: op1_08_in21 = reg_0028;
    30: op1_08_in21 = reg_0503;
    31: op1_08_in21 = reg_0059;
    32: op1_08_in21 = reg_0079;
    34: op1_08_in21 = reg_0397;
    35: op1_08_in21 = reg_0373;
    36: op1_08_in21 = reg_0298;
    37: op1_08_in21 = reg_0600;
    38: op1_08_in21 = imem06_in[39:36];
    40: op1_08_in21 = reg_0426;
    41: op1_08_in21 = reg_0756;
    42: op1_08_in21 = reg_0615;
    44: op1_08_in21 = reg_0824;
    45: op1_08_in21 = imem03_in[71:68];
    46: op1_08_in21 = imem06_in[83:80];
    47: op1_08_in21 = imem01_in[99:96];
    48: op1_08_in21 = reg_0095;
    49: op1_08_in21 = imem01_in[111:108];
    51: op1_08_in21 = imem07_in[63:60];
    52: op1_08_in21 = reg_0178;
    54: op1_08_in21 = reg_0294;
    55: op1_08_in21 = reg_0290;
    56: op1_08_in21 = reg_0342;
    57: op1_08_in21 = reg_0000;
    58: op1_08_in21 = imem03_in[95:92];
    59: op1_08_in21 = imem05_in[59:56];
    74: op1_08_in21 = imem05_in[59:56];
    60: op1_08_in21 = reg_0311;
    61: op1_08_in21 = reg_0816;
    63: op1_08_in21 = imem01_in[39:36];
    64: op1_08_in21 = reg_0743;
    65: op1_08_in21 = imem03_in[127:124];
    66: op1_08_in21 = imem03_in[127:124];
    67: op1_08_in21 = reg_0066;
    68: op1_08_in21 = reg_0168;
    69: op1_08_in21 = reg_0488;
    70: op1_08_in21 = reg_0280;
    71: op1_08_in21 = reg_0202;
    72: op1_08_in21 = reg_0317;
    75: op1_08_in21 = reg_0103;
    76: op1_08_in21 = imem07_in[111:108];
    79: op1_08_in21 = reg_0568;
    80: op1_08_in21 = reg_0771;
    81: op1_08_in21 = imem03_in[75:72];
    82: op1_08_in21 = reg_0388;
    83: op1_08_in21 = reg_0605;
    84: op1_08_in21 = imem03_in[11:8];
    85: op1_08_in21 = reg_0679;
    86: op1_08_in21 = reg_0183;
    87: op1_08_in21 = reg_0306;
    89: op1_08_in21 = reg_0526;
    90: op1_08_in21 = reg_0392;
    91: op1_08_in21 = reg_0009;
    92: op1_08_in21 = reg_0265;
    94: op1_08_in21 = reg_0245;
    95: op1_08_in21 = reg_0253;
    96: op1_08_in21 = imem05_in[67:64];
    default: op1_08_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv21 = 1;
    7: op1_08_inv21 = 1;
    8: op1_08_inv21 = 1;
    10: op1_08_inv21 = 1;
    11: op1_08_inv21 = 1;
    12: op1_08_inv21 = 1;
    15: op1_08_inv21 = 1;
    16: op1_08_inv21 = 1;
    20: op1_08_inv21 = 1;
    21: op1_08_inv21 = 1;
    23: op1_08_inv21 = 1;
    24: op1_08_inv21 = 1;
    26: op1_08_inv21 = 1;
    27: op1_08_inv21 = 1;
    28: op1_08_inv21 = 1;
    30: op1_08_inv21 = 1;
    32: op1_08_inv21 = 1;
    34: op1_08_inv21 = 1;
    35: op1_08_inv21 = 1;
    36: op1_08_inv21 = 1;
    38: op1_08_inv21 = 1;
    43: op1_08_inv21 = 1;
    44: op1_08_inv21 = 1;
    46: op1_08_inv21 = 1;
    47: op1_08_inv21 = 1;
    48: op1_08_inv21 = 1;
    49: op1_08_inv21 = 1;
    51: op1_08_inv21 = 1;
    54: op1_08_inv21 = 1;
    56: op1_08_inv21 = 1;
    57: op1_08_inv21 = 1;
    59: op1_08_inv21 = 1;
    61: op1_08_inv21 = 1;
    62: op1_08_inv21 = 1;
    64: op1_08_inv21 = 1;
    65: op1_08_inv21 = 1;
    67: op1_08_inv21 = 1;
    68: op1_08_inv21 = 1;
    71: op1_08_inv21 = 1;
    76: op1_08_inv21 = 1;
    79: op1_08_inv21 = 1;
    80: op1_08_inv21 = 1;
    82: op1_08_inv21 = 1;
    86: op1_08_inv21 = 1;
    87: op1_08_inv21 = 1;
    92: op1_08_inv21 = 1;
    94: op1_08_inv21 = 1;
    default: op1_08_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in22 = reg_0379;
    5: op1_08_in22 = reg_0743;
    7: op1_08_in22 = reg_0060;
    8: op1_08_in22 = reg_0026;
    9: op1_08_in22 = reg_0536;
    10: op1_08_in22 = reg_0750;
    17: op1_08_in22 = reg_0750;
    11: op1_08_in22 = imem04_in[27:24];
    12: op1_08_in22 = reg_0778;
    13: op1_08_in22 = reg_0663;
    14: op1_08_in22 = imem04_in[59:56];
    15: op1_08_in22 = reg_0164;
    16: op1_08_in22 = imem01_in[87:84];
    18: op1_08_in22 = imem01_in[59:56];
    19: op1_08_in22 = reg_0706;
    20: op1_08_in22 = imem01_in[123:120];
    21: op1_08_in22 = reg_0611;
    22: op1_08_in22 = imem06_in[103:100];
    23: op1_08_in22 = reg_0143;
    24: op1_08_in22 = imem07_in[95:92];
    25: op1_08_in22 = imem03_in[99:96];
    45: op1_08_in22 = imem03_in[99:96];
    26: op1_08_in22 = reg_0172;
    27: op1_08_in22 = reg_0233;
    85: op1_08_in22 = reg_0233;
    28: op1_08_in22 = reg_0749;
    30: op1_08_in22 = reg_0504;
    31: op1_08_in22 = reg_0328;
    32: op1_08_in22 = reg_0065;
    34: op1_08_in22 = reg_0396;
    35: op1_08_in22 = reg_0001;
    36: op1_08_in22 = reg_0258;
    37: op1_08_in22 = reg_0595;
    38: op1_08_in22 = imem06_in[55:52];
    40: op1_08_in22 = reg_0434;
    41: op1_08_in22 = imem03_in[71:68];
    42: op1_08_in22 = reg_0302;
    43: op1_08_in22 = reg_0728;
    44: op1_08_in22 = reg_0825;
    46: op1_08_in22 = imem06_in[95:92];
    47: op1_08_in22 = reg_0235;
    48: op1_08_in22 = reg_0538;
    49: op1_08_in22 = reg_0646;
    51: op1_08_in22 = imem07_in[79:76];
    54: op1_08_in22 = reg_0248;
    55: op1_08_in22 = reg_0234;
    56: op1_08_in22 = reg_0414;
    57: op1_08_in22 = reg_0019;
    58: op1_08_in22 = reg_0063;
    59: op1_08_in22 = imem05_in[63:60];
    60: op1_08_in22 = reg_0640;
    61: op1_08_in22 = reg_0035;
    62: op1_08_in22 = imem01_in[107:104];
    63: op1_08_in22 = imem01_in[43:40];
    64: op1_08_in22 = reg_0097;
    65: op1_08_in22 = reg_0317;
    66: op1_08_in22 = reg_0317;
    67: op1_08_in22 = reg_0145;
    69: op1_08_in22 = reg_0331;
    70: op1_08_in22 = reg_0629;
    71: op1_08_in22 = imem01_in[79:76];
    72: op1_08_in22 = reg_0591;
    73: op1_08_in22 = imem03_in[91:88];
    81: op1_08_in22 = imem03_in[91:88];
    74: op1_08_in22 = imem05_in[103:100];
    75: op1_08_in22 = reg_0334;
    76: op1_08_in22 = imem07_in[123:120];
    78: op1_08_in22 = imem01_in[103:100];
    79: op1_08_in22 = reg_0368;
    80: op1_08_in22 = imem05_in[3:0];
    82: op1_08_in22 = reg_0306;
    83: op1_08_in22 = reg_0814;
    84: op1_08_in22 = imem03_in[35:32];
    86: op1_08_in22 = reg_0325;
    87: op1_08_in22 = reg_0105;
    89: op1_08_in22 = reg_0740;
    90: op1_08_in22 = reg_0056;
    91: op1_08_in22 = reg_0648;
    92: op1_08_in22 = reg_0032;
    93: op1_08_in22 = imem06_in[43:40];
    94: op1_08_in22 = reg_0583;
    95: op1_08_in22 = reg_0447;
    96: op1_08_in22 = imem05_in[79:76];
    default: op1_08_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv22 = 1;
    7: op1_08_inv22 = 1;
    8: op1_08_inv22 = 1;
    10: op1_08_inv22 = 1;
    11: op1_08_inv22 = 1;
    13: op1_08_inv22 = 1;
    14: op1_08_inv22 = 1;
    16: op1_08_inv22 = 1;
    17: op1_08_inv22 = 1;
    19: op1_08_inv22 = 1;
    21: op1_08_inv22 = 1;
    23: op1_08_inv22 = 1;
    27: op1_08_inv22 = 1;
    30: op1_08_inv22 = 1;
    38: op1_08_inv22 = 1;
    40: op1_08_inv22 = 1;
    42: op1_08_inv22 = 1;
    46: op1_08_inv22 = 1;
    57: op1_08_inv22 = 1;
    58: op1_08_inv22 = 1;
    59: op1_08_inv22 = 1;
    62: op1_08_inv22 = 1;
    63: op1_08_inv22 = 1;
    65: op1_08_inv22 = 1;
    67: op1_08_inv22 = 1;
    70: op1_08_inv22 = 1;
    79: op1_08_inv22 = 1;
    80: op1_08_inv22 = 1;
    85: op1_08_inv22 = 1;
    87: op1_08_inv22 = 1;
    89: op1_08_inv22 = 1;
    92: op1_08_inv22 = 1;
    93: op1_08_inv22 = 1;
    95: op1_08_inv22 = 1;
    default: op1_08_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in23 = reg_0349;
    5: op1_08_in23 = reg_0734;
    7: op1_08_in23 = imem03_in[19:16];
    8: op1_08_in23 = reg_0216;
    9: op1_08_in23 = reg_0557;
    10: op1_08_in23 = imem07_in[55:52];
    11: op1_08_in23 = imem04_in[75:72];
    12: op1_08_in23 = reg_0510;
    13: op1_08_in23 = reg_0325;
    14: op1_08_in23 = reg_0544;
    15: op1_08_in23 = reg_0185;
    16: op1_08_in23 = imem01_in[119:116];
    17: op1_08_in23 = reg_0749;
    18: op1_08_in23 = imem01_in[63:60];
    19: op1_08_in23 = reg_0441;
    20: op1_08_in23 = reg_0229;
    94: op1_08_in23 = reg_0229;
    21: op1_08_in23 = reg_0622;
    22: op1_08_in23 = imem06_in[127:124];
    23: op1_08_in23 = reg_0139;
    24: op1_08_in23 = imem07_in[103:100];
    25: op1_08_in23 = reg_0597;
    26: op1_08_in23 = reg_0166;
    27: op1_08_in23 = reg_0511;
    82: op1_08_in23 = reg_0511;
    28: op1_08_in23 = imem07_in[19:16];
    30: op1_08_in23 = reg_0243;
    31: op1_08_in23 = reg_0552;
    32: op1_08_in23 = imem05_in[59:56];
    34: op1_08_in23 = reg_0801;
    57: op1_08_in23 = reg_0801;
    35: op1_08_in23 = reg_0014;
    36: op1_08_in23 = reg_0074;
    70: op1_08_in23 = reg_0074;
    37: op1_08_in23 = reg_0751;
    38: op1_08_in23 = imem06_in[91:88];
    40: op1_08_in23 = reg_0427;
    41: op1_08_in23 = imem03_in[119:116];
    42: op1_08_in23 = reg_0430;
    43: op1_08_in23 = reg_0719;
    44: op1_08_in23 = reg_0759;
    45: op1_08_in23 = imem03_in[115:112];
    46: op1_08_in23 = imem06_in[99:96];
    47: op1_08_in23 = reg_0423;
    48: op1_08_in23 = reg_0093;
    49: op1_08_in23 = reg_0668;
    51: op1_08_in23 = imem07_in[83:80];
    54: op1_08_in23 = reg_0219;
    55: op1_08_in23 = reg_0424;
    56: op1_08_in23 = reg_0590;
    58: op1_08_in23 = reg_0604;
    59: op1_08_in23 = imem05_in[87:84];
    96: op1_08_in23 = imem05_in[87:84];
    60: op1_08_in23 = reg_0296;
    61: op1_08_in23 = reg_0620;
    62: op1_08_in23 = imem01_in[111:108];
    63: op1_08_in23 = imem01_in[67:64];
    64: op1_08_in23 = reg_0769;
    65: op1_08_in23 = reg_0579;
    66: op1_08_in23 = reg_0599;
    67: op1_08_in23 = reg_0142;
    69: op1_08_in23 = imem03_in[111:108];
    71: op1_08_in23 = imem01_in[83:80];
    72: op1_08_in23 = reg_0509;
    73: op1_08_in23 = imem03_in[103:100];
    74: op1_08_in23 = imem05_in[127:124];
    75: op1_08_in23 = reg_0436;
    76: op1_08_in23 = reg_0278;
    78: op1_08_in23 = imem01_in[115:112];
    79: op1_08_in23 = reg_0490;
    80: op1_08_in23 = imem05_in[7:4];
    81: op1_08_in23 = reg_0063;
    83: op1_08_in23 = reg_0298;
    84: op1_08_in23 = imem03_in[87:84];
    85: op1_08_in23 = imem05_in[19:16];
    86: op1_08_in23 = reg_0170;
    87: op1_08_in23 = reg_0670;
    89: op1_08_in23 = reg_0000;
    90: op1_08_in23 = reg_0304;
    91: op1_08_in23 = reg_0575;
    92: op1_08_in23 = reg_0654;
    93: op1_08_in23 = imem06_in[47:44];
    95: op1_08_in23 = reg_0440;
    default: op1_08_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_08_inv23 = 1;
    11: op1_08_inv23 = 1;
    12: op1_08_inv23 = 1;
    15: op1_08_inv23 = 1;
    18: op1_08_inv23 = 1;
    19: op1_08_inv23 = 1;
    24: op1_08_inv23 = 1;
    26: op1_08_inv23 = 1;
    28: op1_08_inv23 = 1;
    32: op1_08_inv23 = 1;
    35: op1_08_inv23 = 1;
    37: op1_08_inv23 = 1;
    40: op1_08_inv23 = 1;
    41: op1_08_inv23 = 1;
    43: op1_08_inv23 = 1;
    51: op1_08_inv23 = 1;
    57: op1_08_inv23 = 1;
    58: op1_08_inv23 = 1;
    59: op1_08_inv23 = 1;
    61: op1_08_inv23 = 1;
    65: op1_08_inv23 = 1;
    66: op1_08_inv23 = 1;
    70: op1_08_inv23 = 1;
    71: op1_08_inv23 = 1;
    73: op1_08_inv23 = 1;
    75: op1_08_inv23 = 1;
    76: op1_08_inv23 = 1;
    78: op1_08_inv23 = 1;
    79: op1_08_inv23 = 1;
    80: op1_08_inv23 = 1;
    83: op1_08_inv23 = 1;
    84: op1_08_inv23 = 1;
    87: op1_08_inv23 = 1;
    90: op1_08_inv23 = 1;
    93: op1_08_inv23 = 1;
    95: op1_08_inv23 = 1;
    default: op1_08_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in24 = reg_0403;
    5: op1_08_in24 = reg_0747;
    7: op1_08_in24 = imem03_in[23:20];
    8: op1_08_in24 = reg_0020;
    9: op1_08_in24 = reg_0534;
    10: op1_08_in24 = imem07_in[95:92];
    11: op1_08_in24 = imem04_in[87:84];
    12: op1_08_in24 = reg_0225;
    13: op1_08_in24 = reg_0326;
    14: op1_08_in24 = reg_0530;
    15: op1_08_in24 = reg_0158;
    16: op1_08_in24 = reg_0500;
    17: op1_08_in24 = imem07_in[19:16];
    18: op1_08_in24 = reg_0501;
    19: op1_08_in24 = reg_0429;
    20: op1_08_in24 = reg_0755;
    21: op1_08_in24 = reg_0402;
    22: op1_08_in24 = reg_0629;
    23: op1_08_in24 = reg_0129;
    24: op1_08_in24 = reg_0727;
    25: op1_08_in24 = reg_0581;
    26: op1_08_in24 = reg_0184;
    27: op1_08_in24 = reg_0242;
    28: op1_08_in24 = imem07_in[67:64];
    30: op1_08_in24 = reg_0111;
    31: op1_08_in24 = reg_0537;
    32: op1_08_in24 = imem05_in[115:112];
    34: op1_08_in24 = imem04_in[35:32];
    35: op1_08_in24 = reg_0008;
    36: op1_08_in24 = reg_0288;
    37: op1_08_in24 = reg_0395;
    38: op1_08_in24 = imem06_in[107:104];
    40: op1_08_in24 = reg_0437;
    41: op1_08_in24 = reg_0596;
    65: op1_08_in24 = reg_0596;
    89: op1_08_in24 = reg_0596;
    42: op1_08_in24 = reg_0071;
    43: op1_08_in24 = reg_0710;
    44: op1_08_in24 = reg_0771;
    45: op1_08_in24 = reg_0582;
    46: op1_08_in24 = reg_0247;
    47: op1_08_in24 = reg_0306;
    48: op1_08_in24 = imem03_in[7:4];
    49: op1_08_in24 = reg_0645;
    51: op1_08_in24 = imem07_in[99:96];
    54: op1_08_in24 = reg_0123;
    55: op1_08_in24 = reg_0073;
    56: op1_08_in24 = reg_0323;
    57: op1_08_in24 = reg_0800;
    58: op1_08_in24 = reg_0357;
    59: op1_08_in24 = reg_0791;
    60: op1_08_in24 = reg_0275;
    61: op1_08_in24 = reg_0819;
    62: op1_08_in24 = reg_0085;
    78: op1_08_in24 = reg_0085;
    63: op1_08_in24 = imem01_in[115:112];
    64: op1_08_in24 = reg_0756;
    66: op1_08_in24 = reg_0579;
    67: op1_08_in24 = reg_0134;
    69: op1_08_in24 = imem03_in[115:112];
    84: op1_08_in24 = imem03_in[115:112];
    70: op1_08_in24 = reg_0301;
    71: op1_08_in24 = reg_0497;
    72: op1_08_in24 = reg_0331;
    73: op1_08_in24 = reg_0589;
    74: op1_08_in24 = reg_0070;
    75: op1_08_in24 = reg_0333;
    76: op1_08_in24 = reg_0157;
    79: op1_08_in24 = reg_0569;
    80: op1_08_in24 = imem05_in[11:8];
    81: op1_08_in24 = reg_0347;
    82: op1_08_in24 = reg_0216;
    83: op1_08_in24 = reg_0238;
    85: op1_08_in24 = imem05_in[27:24];
    86: op1_08_in24 = reg_0427;
    87: op1_08_in24 = reg_0119;
    90: op1_08_in24 = reg_0256;
    91: op1_08_in24 = reg_0372;
    92: op1_08_in24 = reg_0307;
    93: op1_08_in24 = imem06_in[55:52];
    94: op1_08_in24 = reg_0827;
    95: op1_08_in24 = reg_0435;
    96: op1_08_in24 = imem05_in[107:104];
    default: op1_08_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv24 = 1;
    8: op1_08_inv24 = 1;
    10: op1_08_inv24 = 1;
    11: op1_08_inv24 = 1;
    14: op1_08_inv24 = 1;
    15: op1_08_inv24 = 1;
    17: op1_08_inv24 = 1;
    22: op1_08_inv24 = 1;
    26: op1_08_inv24 = 1;
    28: op1_08_inv24 = 1;
    34: op1_08_inv24 = 1;
    36: op1_08_inv24 = 1;
    37: op1_08_inv24 = 1;
    38: op1_08_inv24 = 1;
    41: op1_08_inv24 = 1;
    46: op1_08_inv24 = 1;
    47: op1_08_inv24 = 1;
    48: op1_08_inv24 = 1;
    49: op1_08_inv24 = 1;
    51: op1_08_inv24 = 1;
    56: op1_08_inv24 = 1;
    58: op1_08_inv24 = 1;
    59: op1_08_inv24 = 1;
    60: op1_08_inv24 = 1;
    61: op1_08_inv24 = 1;
    62: op1_08_inv24 = 1;
    64: op1_08_inv24 = 1;
    65: op1_08_inv24 = 1;
    69: op1_08_inv24 = 1;
    70: op1_08_inv24 = 1;
    72: op1_08_inv24 = 1;
    75: op1_08_inv24 = 1;
    80: op1_08_inv24 = 1;
    81: op1_08_inv24 = 1;
    83: op1_08_inv24 = 1;
    84: op1_08_inv24 = 1;
    86: op1_08_inv24 = 1;
    87: op1_08_inv24 = 1;
    90: op1_08_inv24 = 1;
    91: op1_08_inv24 = 1;
    93: op1_08_inv24 = 1;
    default: op1_08_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in25 = reg_0367;
    5: op1_08_in25 = imem05_in[19:16];
    7: op1_08_in25 = imem03_in[51:48];
    8: op1_08_in25 = reg_0220;
    9: op1_08_in25 = reg_0555;
    10: op1_08_in25 = imem07_in[103:100];
    28: op1_08_in25 = imem07_in[103:100];
    11: op1_08_in25 = imem04_in[127:124];
    12: op1_08_in25 = reg_0232;
    13: op1_08_in25 = reg_0359;
    14: op1_08_in25 = reg_0553;
    16: op1_08_in25 = reg_0225;
    17: op1_08_in25 = imem07_in[23:20];
    18: op1_08_in25 = reg_0509;
    19: op1_08_in25 = reg_0428;
    20: op1_08_in25 = reg_0241;
    21: op1_08_in25 = reg_0379;
    22: op1_08_in25 = reg_0616;
    23: op1_08_in25 = reg_0141;
    24: op1_08_in25 = reg_0175;
    25: op1_08_in25 = reg_0590;
    27: op1_08_in25 = reg_0216;
    30: op1_08_in25 = reg_0116;
    31: op1_08_in25 = reg_0056;
    32: op1_08_in25 = reg_0798;
    59: op1_08_in25 = reg_0798;
    34: op1_08_in25 = imem04_in[43:40];
    35: op1_08_in25 = reg_0015;
    36: op1_08_in25 = imem05_in[3:0];
    37: op1_08_in25 = reg_0387;
    38: op1_08_in25 = imem06_in[127:124];
    40: op1_08_in25 = reg_0438;
    41: op1_08_in25 = reg_0592;
    55: op1_08_in25 = reg_0592;
    42: op1_08_in25 = reg_0627;
    43: op1_08_in25 = reg_0731;
    44: op1_08_in25 = reg_0761;
    45: op1_08_in25 = reg_0601;
    46: op1_08_in25 = reg_0609;
    47: op1_08_in25 = reg_0294;
    82: op1_08_in25 = reg_0294;
    48: op1_08_in25 = imem03_in[47:44];
    49: op1_08_in25 = reg_0825;
    51: op1_08_in25 = imem07_in[107:104];
    54: op1_08_in25 = reg_0671;
    56: op1_08_in25 = reg_0541;
    57: op1_08_in25 = reg_0014;
    58: op1_08_in25 = reg_0573;
    60: op1_08_in25 = reg_0483;
    61: op1_08_in25 = reg_0368;
    62: op1_08_in25 = reg_0497;
    63: op1_08_in25 = reg_0668;
    64: op1_08_in25 = reg_0098;
    65: op1_08_in25 = reg_0591;
    66: op1_08_in25 = reg_0488;
    67: op1_08_in25 = imem06_in[11:8];
    69: op1_08_in25 = reg_0012;
    70: op1_08_in25 = reg_0640;
    71: op1_08_in25 = reg_0772;
    72: op1_08_in25 = reg_0568;
    73: op1_08_in25 = reg_0596;
    74: op1_08_in25 = reg_0146;
    75: op1_08_in25 = reg_0439;
    76: op1_08_in25 = reg_0727;
    78: op1_08_in25 = reg_0520;
    79: op1_08_in25 = reg_0398;
    80: op1_08_in25 = imem05_in[51:48];
    81: op1_08_in25 = reg_0589;
    83: op1_08_in25 = reg_0293;
    84: op1_08_in25 = reg_0317;
    85: op1_08_in25 = imem05_in[35:32];
    86: op1_08_in25 = reg_0184;
    87: op1_08_in25 = reg_0677;
    89: op1_08_in25 = reg_0803;
    90: op1_08_in25 = reg_0251;
    91: op1_08_in25 = reg_0490;
    92: op1_08_in25 = reg_0750;
    93: op1_08_in25 = imem06_in[83:80];
    94: op1_08_in25 = reg_0742;
    95: op1_08_in25 = reg_0228;
    96: op1_08_in25 = imem05_in[123:120];
    default: op1_08_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv25 = 1;
    7: op1_08_inv25 = 1;
    8: op1_08_inv25 = 1;
    10: op1_08_inv25 = 1;
    11: op1_08_inv25 = 1;
    12: op1_08_inv25 = 1;
    13: op1_08_inv25 = 1;
    16: op1_08_inv25 = 1;
    18: op1_08_inv25 = 1;
    20: op1_08_inv25 = 1;
    22: op1_08_inv25 = 1;
    24: op1_08_inv25 = 1;
    28: op1_08_inv25 = 1;
    31: op1_08_inv25 = 1;
    36: op1_08_inv25 = 1;
    37: op1_08_inv25 = 1;
    38: op1_08_inv25 = 1;
    40: op1_08_inv25 = 1;
    43: op1_08_inv25 = 1;
    46: op1_08_inv25 = 1;
    54: op1_08_inv25 = 1;
    55: op1_08_inv25 = 1;
    56: op1_08_inv25 = 1;
    58: op1_08_inv25 = 1;
    59: op1_08_inv25 = 1;
    62: op1_08_inv25 = 1;
    66: op1_08_inv25 = 1;
    67: op1_08_inv25 = 1;
    71: op1_08_inv25 = 1;
    72: op1_08_inv25 = 1;
    73: op1_08_inv25 = 1;
    74: op1_08_inv25 = 1;
    78: op1_08_inv25 = 1;
    79: op1_08_inv25 = 1;
    83: op1_08_inv25 = 1;
    84: op1_08_inv25 = 1;
    85: op1_08_inv25 = 1;
    89: op1_08_inv25 = 1;
    93: op1_08_inv25 = 1;
    94: op1_08_inv25 = 1;
    95: op1_08_inv25 = 1;
    96: op1_08_inv25 = 1;
    default: op1_08_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in26 = reg_0380;
    5: op1_08_in26 = imem05_in[67:64];
    7: op1_08_in26 = imem03_in[63:60];
    8: op1_08_in26 = reg_0630;
    9: op1_08_in26 = reg_0558;
    10: op1_08_in26 = imem07_in[107:104];
    11: op1_08_in26 = reg_0540;
    12: op1_08_in26 = reg_0506;
    13: op1_08_in26 = reg_0339;
    14: op1_08_in26 = reg_0529;
    16: op1_08_in26 = reg_0505;
    20: op1_08_in26 = reg_0505;
    17: op1_08_in26 = imem07_in[27:24];
    18: op1_08_in26 = reg_0520;
    19: op1_08_in26 = reg_0446;
    21: op1_08_in26 = reg_0372;
    22: op1_08_in26 = reg_0618;
    23: op1_08_in26 = imem06_in[63:60];
    24: op1_08_in26 = reg_0165;
    25: op1_08_in26 = reg_0370;
    27: op1_08_in26 = reg_0245;
    28: op1_08_in26 = imem07_in[119:116];
    30: op1_08_in26 = imem02_in[79:76];
    31: op1_08_in26 = reg_0055;
    32: op1_08_in26 = reg_0788;
    34: op1_08_in26 = imem04_in[59:56];
    35: op1_08_in26 = reg_0799;
    36: op1_08_in26 = imem05_in[7:4];
    37: op1_08_in26 = reg_0755;
    38: op1_08_in26 = reg_0025;
    40: op1_08_in26 = reg_0435;
    41: op1_08_in26 = reg_0590;
    42: op1_08_in26 = reg_0281;
    66: op1_08_in26 = reg_0281;
    43: op1_08_in26 = reg_0723;
    44: op1_08_in26 = reg_0422;
    45: op1_08_in26 = reg_0579;
    46: op1_08_in26 = reg_0633;
    47: op1_08_in26 = reg_0234;
    48: op1_08_in26 = imem03_in[51:48];
    49: op1_08_in26 = reg_0237;
    51: op1_08_in26 = reg_0728;
    54: op1_08_in26 = imem02_in[15:12];
    55: op1_08_in26 = imem02_in[3:0];
    56: op1_08_in26 = reg_0530;
    57: op1_08_in26 = reg_0016;
    58: op1_08_in26 = reg_0572;
    59: op1_08_in26 = reg_0796;
    60: op1_08_in26 = reg_0336;
    61: op1_08_in26 = reg_0787;
    62: op1_08_in26 = reg_0668;
    63: op1_08_in26 = reg_0759;
    64: op1_08_in26 = reg_0498;
    65: op1_08_in26 = reg_0528;
    67: op1_08_in26 = imem06_in[15:12];
    69: op1_08_in26 = reg_0803;
    70: op1_08_in26 = reg_0296;
    71: op1_08_in26 = reg_0110;
    72: op1_08_in26 = reg_0483;
    73: op1_08_in26 = reg_0318;
    74: op1_08_in26 = reg_0782;
    75: op1_08_in26 = reg_0267;
    76: op1_08_in26 = reg_0295;
    78: op1_08_in26 = reg_0645;
    79: op1_08_in26 = reg_0802;
    80: op1_08_in26 = imem05_in[63:60];
    81: op1_08_in26 = reg_0599;
    82: op1_08_in26 = reg_0425;
    83: op1_08_in26 = reg_0401;
    84: op1_08_in26 = reg_0493;
    85: op1_08_in26 = imem05_in[87:84];
    87: op1_08_in26 = reg_0127;
    89: op1_08_in26 = reg_0329;
    90: op1_08_in26 = reg_0364;
    91: op1_08_in26 = reg_0396;
    92: op1_08_in26 = reg_0576;
    93: op1_08_in26 = imem06_in[103:100];
    94: op1_08_in26 = reg_0830;
    96: op1_08_in26 = reg_0791;
    default: op1_08_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv26 = 1;
    5: op1_08_inv26 = 1;
    7: op1_08_inv26 = 1;
    8: op1_08_inv26 = 1;
    9: op1_08_inv26 = 1;
    11: op1_08_inv26 = 1;
    14: op1_08_inv26 = 1;
    17: op1_08_inv26 = 1;
    18: op1_08_inv26 = 1;
    22: op1_08_inv26 = 1;
    23: op1_08_inv26 = 1;
    30: op1_08_inv26 = 1;
    31: op1_08_inv26 = 1;
    34: op1_08_inv26 = 1;
    36: op1_08_inv26 = 1;
    38: op1_08_inv26 = 1;
    40: op1_08_inv26 = 1;
    41: op1_08_inv26 = 1;
    45: op1_08_inv26 = 1;
    47: op1_08_inv26 = 1;
    49: op1_08_inv26 = 1;
    51: op1_08_inv26 = 1;
    54: op1_08_inv26 = 1;
    55: op1_08_inv26 = 1;
    61: op1_08_inv26 = 1;
    64: op1_08_inv26 = 1;
    65: op1_08_inv26 = 1;
    66: op1_08_inv26 = 1;
    67: op1_08_inv26 = 1;
    69: op1_08_inv26 = 1;
    71: op1_08_inv26 = 1;
    73: op1_08_inv26 = 1;
    76: op1_08_inv26 = 1;
    78: op1_08_inv26 = 1;
    81: op1_08_inv26 = 1;
    87: op1_08_inv26 = 1;
    89: op1_08_inv26 = 1;
    93: op1_08_inv26 = 1;
    94: op1_08_inv26 = 1;
    96: op1_08_inv26 = 1;
    default: op1_08_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in27 = reg_0026;
    5: op1_08_in27 = imem05_in[75:72];
    7: op1_08_in27 = reg_0579;
    8: op1_08_in27 = reg_0624;
    9: op1_08_in27 = reg_0559;
    10: op1_08_in27 = imem07_in[115:112];
    11: op1_08_in27 = reg_0304;
    12: op1_08_in27 = reg_0217;
    13: op1_08_in27 = reg_0346;
    14: op1_08_in27 = reg_0537;
    16: op1_08_in27 = reg_0503;
    17: op1_08_in27 = imem07_in[31:28];
    18: op1_08_in27 = reg_0519;
    19: op1_08_in27 = reg_0175;
    20: op1_08_in27 = reg_0506;
    82: op1_08_in27 = reg_0506;
    21: op1_08_in27 = reg_0407;
    22: op1_08_in27 = reg_0402;
    23: op1_08_in27 = imem06_in[95:92];
    24: op1_08_in27 = reg_0179;
    25: op1_08_in27 = reg_0369;
    27: op1_08_in27 = reg_0238;
    28: op1_08_in27 = reg_0714;
    30: op1_08_in27 = imem02_in[83:80];
    31: op1_08_in27 = reg_0083;
    32: op1_08_in27 = reg_0493;
    81: op1_08_in27 = reg_0493;
    34: op1_08_in27 = imem04_in[63:60];
    35: op1_08_in27 = imem04_in[43:40];
    36: op1_08_in27 = imem05_in[39:36];
    37: op1_08_in27 = reg_0562;
    38: op1_08_in27 = reg_0317;
    40: op1_08_in27 = reg_0431;
    41: op1_08_in27 = reg_0385;
    42: op1_08_in27 = reg_0065;
    43: op1_08_in27 = reg_0700;
    44: op1_08_in27 = reg_0425;
    45: op1_08_in27 = reg_0597;
    46: op1_08_in27 = reg_0618;
    47: op1_08_in27 = reg_0505;
    48: op1_08_in27 = imem03_in[67:64];
    49: op1_08_in27 = reg_0737;
    51: op1_08_in27 = reg_0720;
    54: op1_08_in27 = imem02_in[31:28];
    55: op1_08_in27 = imem02_in[7:4];
    56: op1_08_in27 = reg_0540;
    57: op1_08_in27 = reg_0806;
    58: op1_08_in27 = reg_0386;
    59: op1_08_in27 = reg_0490;
    60: op1_08_in27 = reg_0788;
    61: op1_08_in27 = reg_0495;
    62: op1_08_in27 = reg_0663;
    63: op1_08_in27 = reg_0557;
    64: op1_08_in27 = reg_0094;
    65: op1_08_in27 = reg_0329;
    66: op1_08_in27 = reg_0575;
    67: op1_08_in27 = imem06_in[39:36];
    69: op1_08_in27 = reg_0807;
    70: op1_08_in27 = reg_0233;
    71: op1_08_in27 = reg_0507;
    72: op1_08_in27 = reg_0012;
    73: op1_08_in27 = reg_0528;
    74: op1_08_in27 = reg_0245;
    75: op1_08_in27 = reg_0448;
    76: op1_08_in27 = reg_0447;
    78: op1_08_in27 = reg_0114;
    79: op1_08_in27 = reg_0015;
    80: op1_08_in27 = imem05_in[83:80];
    83: op1_08_in27 = reg_0578;
    84: op1_08_in27 = reg_0600;
    85: op1_08_in27 = reg_0792;
    87: op1_08_in27 = reg_0126;
    89: op1_08_in27 = reg_0145;
    90: op1_08_in27 = reg_0586;
    91: op1_08_in27 = reg_0623;
    92: op1_08_in27 = reg_0335;
    93: op1_08_in27 = imem06_in[115:112];
    94: op1_08_in27 = reg_0155;
    96: op1_08_in27 = reg_0667;
    default: op1_08_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv27 = 1;
    5: op1_08_inv27 = 1;
    7: op1_08_inv27 = 1;
    8: op1_08_inv27 = 1;
    10: op1_08_inv27 = 1;
    11: op1_08_inv27 = 1;
    12: op1_08_inv27 = 1;
    13: op1_08_inv27 = 1;
    14: op1_08_inv27 = 1;
    17: op1_08_inv27 = 1;
    18: op1_08_inv27 = 1;
    19: op1_08_inv27 = 1;
    20: op1_08_inv27 = 1;
    21: op1_08_inv27 = 1;
    22: op1_08_inv27 = 1;
    24: op1_08_inv27 = 1;
    25: op1_08_inv27 = 1;
    27: op1_08_inv27 = 1;
    31: op1_08_inv27 = 1;
    36: op1_08_inv27 = 1;
    41: op1_08_inv27 = 1;
    43: op1_08_inv27 = 1;
    45: op1_08_inv27 = 1;
    46: op1_08_inv27 = 1;
    48: op1_08_inv27 = 1;
    49: op1_08_inv27 = 1;
    54: op1_08_inv27 = 1;
    58: op1_08_inv27 = 1;
    59: op1_08_inv27 = 1;
    61: op1_08_inv27 = 1;
    63: op1_08_inv27 = 1;
    66: op1_08_inv27 = 1;
    67: op1_08_inv27 = 1;
    69: op1_08_inv27 = 1;
    71: op1_08_inv27 = 1;
    73: op1_08_inv27 = 1;
    75: op1_08_inv27 = 1;
    76: op1_08_inv27 = 1;
    78: op1_08_inv27 = 1;
    83: op1_08_inv27 = 1;
    85: op1_08_inv27 = 1;
    87: op1_08_inv27 = 1;
    91: op1_08_inv27 = 1;
    96: op1_08_inv27 = 1;
    default: op1_08_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in28 = reg_0020;
    5: op1_08_in28 = imem05_in[103:100];
    7: op1_08_in28 = reg_0569;
    8: op1_08_in28 = reg_0633;
    9: op1_08_in28 = reg_0531;
    56: op1_08_in28 = reg_0531;
    10: op1_08_in28 = imem07_in[127:124];
    11: op1_08_in28 = reg_0279;
    12: op1_08_in28 = reg_0242;
    13: op1_08_in28 = reg_0353;
    14: op1_08_in28 = reg_0549;
    16: op1_08_in28 = reg_0248;
    17: op1_08_in28 = imem07_in[67:64];
    18: op1_08_in28 = reg_0521;
    19: op1_08_in28 = reg_0180;
    20: op1_08_in28 = reg_0216;
    21: op1_08_in28 = reg_0403;
    22: op1_08_in28 = reg_0344;
    23: op1_08_in28 = imem06_in[127:124];
    24: op1_08_in28 = reg_0161;
    25: op1_08_in28 = reg_0377;
    89: op1_08_in28 = reg_0377;
    27: op1_08_in28 = reg_0243;
    28: op1_08_in28 = reg_0711;
    30: op1_08_in28 = imem02_in[87:84];
    31: op1_08_in28 = reg_0054;
    32: op1_08_in28 = reg_0494;
    34: op1_08_in28 = imem04_in[71:68];
    35: op1_08_in28 = imem04_in[55:52];
    36: op1_08_in28 = imem05_in[63:60];
    37: op1_08_in28 = reg_0747;
    38: op1_08_in28 = reg_0331;
    40: op1_08_in28 = reg_0166;
    41: op1_08_in28 = reg_0562;
    66: op1_08_in28 = reg_0562;
    42: op1_08_in28 = reg_0063;
    43: op1_08_in28 = reg_0727;
    44: op1_08_in28 = reg_0504;
    45: op1_08_in28 = reg_0595;
    46: op1_08_in28 = reg_0317;
    47: op1_08_in28 = reg_0123;
    48: op1_08_in28 = imem03_in[71:68];
    49: op1_08_in28 = reg_0550;
    51: op1_08_in28 = reg_0721;
    54: op1_08_in28 = imem02_in[79:76];
    55: op1_08_in28 = imem02_in[67:64];
    57: op1_08_in28 = reg_0809;
    58: op1_08_in28 = reg_0001;
    59: op1_08_in28 = reg_0795;
    60: op1_08_in28 = reg_0785;
    61: op1_08_in28 = imem07_in[3:0];
    62: op1_08_in28 = reg_0322;
    63: op1_08_in28 = reg_0421;
    64: op1_08_in28 = reg_0532;
    65: op1_08_in28 = reg_0281;
    67: op1_08_in28 = imem06_in[103:100];
    69: op1_08_in28 = reg_0014;
    70: op1_08_in28 = reg_0644;
    71: op1_08_in28 = reg_0306;
    72: op1_08_in28 = reg_0801;
    73: op1_08_in28 = reg_0350;
    74: op1_08_in28 = reg_0040;
    75: op1_08_in28 = reg_0162;
    76: op1_08_in28 = reg_0175;
    78: op1_08_in28 = reg_0131;
    79: op1_08_in28 = imem04_in[31:28];
    80: op1_08_in28 = imem05_in[127:124];
    81: op1_08_in28 = reg_0591;
    82: op1_08_in28 = reg_0219;
    83: op1_08_in28 = reg_0659;
    84: op1_08_in28 = reg_0588;
    85: op1_08_in28 = reg_0736;
    87: op1_08_in28 = imem02_in[19:16];
    90: op1_08_in28 = reg_0341;
    91: op1_08_in28 = reg_0649;
    92: op1_08_in28 = reg_0664;
    93: op1_08_in28 = reg_0289;
    94: op1_08_in28 = reg_0824;
    96: op1_08_in28 = reg_0788;
    default: op1_08_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv28 = 1;
    7: op1_08_inv28 = 1;
    12: op1_08_inv28 = 1;
    13: op1_08_inv28 = 1;
    17: op1_08_inv28 = 1;
    19: op1_08_inv28 = 1;
    20: op1_08_inv28 = 1;
    22: op1_08_inv28 = 1;
    25: op1_08_inv28 = 1;
    40: op1_08_inv28 = 1;
    44: op1_08_inv28 = 1;
    45: op1_08_inv28 = 1;
    46: op1_08_inv28 = 1;
    48: op1_08_inv28 = 1;
    51: op1_08_inv28 = 1;
    54: op1_08_inv28 = 1;
    55: op1_08_inv28 = 1;
    59: op1_08_inv28 = 1;
    61: op1_08_inv28 = 1;
    63: op1_08_inv28 = 1;
    64: op1_08_inv28 = 1;
    67: op1_08_inv28 = 1;
    69: op1_08_inv28 = 1;
    70: op1_08_inv28 = 1;
    71: op1_08_inv28 = 1;
    72: op1_08_inv28 = 1;
    74: op1_08_inv28 = 1;
    78: op1_08_inv28 = 1;
    81: op1_08_inv28 = 1;
    82: op1_08_inv28 = 1;
    83: op1_08_inv28 = 1;
    84: op1_08_inv28 = 1;
    87: op1_08_inv28 = 1;
    89: op1_08_inv28 = 1;
    90: op1_08_inv28 = 1;
    94: op1_08_inv28 = 1;
    96: op1_08_inv28 = 1;
    default: op1_08_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in29 = reg_0030;
    5: op1_08_in29 = imem05_in[107:104];
    7: op1_08_in29 = reg_0595;
    73: op1_08_in29 = reg_0595;
    81: op1_08_in29 = reg_0595;
    8: op1_08_in29 = reg_0608;
    9: op1_08_in29 = reg_0281;
    10: op1_08_in29 = reg_0719;
    11: op1_08_in29 = reg_0306;
    12: op1_08_in29 = reg_0216;
    13: op1_08_in29 = reg_0089;
    14: op1_08_in29 = reg_0558;
    16: op1_08_in29 = reg_0504;
    17: op1_08_in29 = imem07_in[79:76];
    18: op1_08_in29 = reg_0778;
    19: op1_08_in29 = reg_0159;
    20: op1_08_in29 = reg_0248;
    21: op1_08_in29 = reg_0390;
    22: op1_08_in29 = reg_0405;
    23: op1_08_in29 = reg_0628;
    24: op1_08_in29 = reg_0169;
    25: op1_08_in29 = reg_0398;
    27: op1_08_in29 = reg_0108;
    28: op1_08_in29 = reg_0706;
    30: op1_08_in29 = imem02_in[91:88];
    31: op1_08_in29 = reg_0301;
    32: op1_08_in29 = reg_0304;
    34: op1_08_in29 = imem04_in[83:80];
    35: op1_08_in29 = imem04_in[63:60];
    36: op1_08_in29 = imem05_in[91:88];
    37: op1_08_in29 = reg_0570;
    38: op1_08_in29 = reg_0577;
    46: op1_08_in29 = reg_0577;
    40: op1_08_in29 = reg_0157;
    41: op1_08_in29 = reg_0000;
    42: op1_08_in29 = reg_0069;
    43: op1_08_in29 = reg_0253;
    44: op1_08_in29 = reg_0424;
    45: op1_08_in29 = reg_0387;
    47: op1_08_in29 = reg_0122;
    48: op1_08_in29 = imem03_in[111:108];
    49: op1_08_in29 = reg_0235;
    51: op1_08_in29 = reg_0709;
    54: op1_08_in29 = imem02_in[123:120];
    55: op1_08_in29 = imem02_in[71:68];
    56: op1_08_in29 = reg_0094;
    57: op1_08_in29 = imem04_in[11:8];
    58: op1_08_in29 = reg_0800;
    59: op1_08_in29 = reg_0288;
    60: op1_08_in29 = reg_0269;
    61: op1_08_in29 = imem07_in[19:16];
    62: op1_08_in29 = reg_0100;
    63: op1_08_in29 = reg_0567;
    64: op1_08_in29 = imem03_in[43:40];
    65: op1_08_in29 = reg_0357;
    66: op1_08_in29 = reg_0572;
    67: op1_08_in29 = imem06_in[107:104];
    69: op1_08_in29 = reg_0802;
    70: op1_08_in29 = imem05_in[51:48];
    71: op1_08_in29 = reg_0217;
    72: op1_08_in29 = reg_0015;
    74: op1_08_in29 = reg_0812;
    75: op1_08_in29 = reg_0160;
    76: op1_08_in29 = reg_0172;
    78: op1_08_in29 = reg_0110;
    79: op1_08_in29 = imem04_in[35:32];
    80: op1_08_in29 = reg_0667;
    82: op1_08_in29 = reg_0420;
    83: op1_08_in29 = reg_0654;
    84: op1_08_in29 = reg_0648;
    85: op1_08_in29 = reg_0145;
    87: op1_08_in29 = imem02_in[51:48];
    89: op1_08_in29 = reg_0016;
    90: op1_08_in29 = reg_0359;
    91: op1_08_in29 = reg_0561;
    92: op1_08_in29 = reg_0037;
    93: op1_08_in29 = reg_0348;
    94: op1_08_in29 = reg_0734;
    96: op1_08_in29 = reg_0641;
    default: op1_08_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_08_inv29 = 1;
    5: op1_08_inv29 = 1;
    9: op1_08_inv29 = 1;
    11: op1_08_inv29 = 1;
    12: op1_08_inv29 = 1;
    14: op1_08_inv29 = 1;
    16: op1_08_inv29 = 1;
    17: op1_08_inv29 = 1;
    19: op1_08_inv29 = 1;
    21: op1_08_inv29 = 1;
    24: op1_08_inv29 = 1;
    25: op1_08_inv29 = 1;
    27: op1_08_inv29 = 1;
    28: op1_08_inv29 = 1;
    32: op1_08_inv29 = 1;
    38: op1_08_inv29 = 1;
    40: op1_08_inv29 = 1;
    41: op1_08_inv29 = 1;
    43: op1_08_inv29 = 1;
    44: op1_08_inv29 = 1;
    56: op1_08_inv29 = 1;
    60: op1_08_inv29 = 1;
    61: op1_08_inv29 = 1;
    65: op1_08_inv29 = 1;
    66: op1_08_inv29 = 1;
    67: op1_08_inv29 = 1;
    70: op1_08_inv29 = 1;
    71: op1_08_inv29 = 1;
    72: op1_08_inv29 = 1;
    79: op1_08_inv29 = 1;
    80: op1_08_inv29 = 1;
    81: op1_08_inv29 = 1;
    82: op1_08_inv29 = 1;
    84: op1_08_inv29 = 1;
    85: op1_08_inv29 = 1;
    90: op1_08_inv29 = 1;
    93: op1_08_inv29 = 1;
    94: op1_08_inv29 = 1;
    96: op1_08_inv29 = 1;
    default: op1_08_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_08_in30 = reg_0011;
    5: op1_08_in30 = imem05_in[119:116];
    7: op1_08_in30 = reg_0588;
    81: op1_08_in30 = reg_0588;
    8: op1_08_in30 = reg_0632;
    9: op1_08_in30 = reg_0279;
    10: op1_08_in30 = reg_0731;
    11: op1_08_in30 = reg_0291;
    12: op1_08_in30 = reg_0248;
    13: op1_08_in30 = reg_0095;
    14: op1_08_in30 = reg_0282;
    16: op1_08_in30 = reg_0245;
    17: op1_08_in30 = imem07_in[99:96];
    18: op1_08_in30 = reg_0232;
    19: op1_08_in30 = reg_0182;
    20: op1_08_in30 = reg_0504;
    21: op1_08_in30 = reg_0380;
    22: op1_08_in30 = reg_0812;
    23: op1_08_in30 = reg_0620;
    24: op1_08_in30 = reg_0183;
    25: op1_08_in30 = reg_0376;
    27: op1_08_in30 = reg_0114;
    28: op1_08_in30 = reg_0430;
    30: op1_08_in30 = imem02_in[111:108];
    31: op1_08_in30 = reg_0305;
    32: op1_08_in30 = reg_0085;
    34: op1_08_in30 = imem04_in[95:92];
    35: op1_08_in30 = imem04_in[83:80];
    36: op1_08_in30 = reg_0796;
    37: op1_08_in30 = reg_0002;
    38: op1_08_in30 = reg_0370;
    41: op1_08_in30 = reg_0006;
    42: op1_08_in30 = imem05_in[27:24];
    43: op1_08_in30 = reg_0053;
    44: op1_08_in30 = reg_0111;
    45: op1_08_in30 = reg_0573;
    46: op1_08_in30 = reg_0775;
    47: op1_08_in30 = reg_0119;
    48: op1_08_in30 = imem03_in[119:116];
    49: op1_08_in30 = reg_0306;
    51: op1_08_in30 = reg_0715;
    54: op1_08_in30 = reg_0662;
    55: op1_08_in30 = imem02_in[75:72];
    56: op1_08_in30 = reg_0093;
    57: op1_08_in30 = imem04_in[19:16];
    58: op1_08_in30 = reg_0484;
    59: op1_08_in30 = reg_0793;
    80: op1_08_in30 = reg_0793;
    60: op1_08_in30 = reg_0403;
    61: op1_08_in30 = imem07_in[23:20];
    62: op1_08_in30 = reg_0737;
    63: op1_08_in30 = reg_0240;
    64: op1_08_in30 = imem03_in[51:48];
    65: op1_08_in30 = reg_0755;
    66: op1_08_in30 = reg_0747;
    67: op1_08_in30 = imem06_in[119:116];
    69: op1_08_in30 = imem04_in[79:76];
    70: op1_08_in30 = imem05_in[87:84];
    71: op1_08_in30 = reg_0567;
    72: op1_08_in30 = reg_0806;
    73: op1_08_in30 = reg_0751;
    74: op1_08_in30 = reg_0147;
    75: op1_08_in30 = reg_0163;
    78: op1_08_in30 = reg_0574;
    79: op1_08_in30 = imem04_in[67:64];
    82: op1_08_in30 = reg_0104;
    83: op1_08_in30 = reg_0405;
    84: op1_08_in30 = reg_0564;
    85: op1_08_in30 = reg_0666;
    87: op1_08_in30 = imem02_in[79:76];
    89: op1_08_in30 = reg_0375;
    90: op1_08_in30 = reg_0361;
    91: op1_08_in30 = reg_0216;
    92: op1_08_in30 = imem07_in[27:24];
    93: op1_08_in30 = reg_0349;
    94: op1_08_in30 = imem06_in[27:24];
    96: op1_08_in30 = reg_0113;
    default: op1_08_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_08_inv30 = 1;
    10: op1_08_inv30 = 1;
    11: op1_08_inv30 = 1;
    12: op1_08_inv30 = 1;
    13: op1_08_inv30 = 1;
    14: op1_08_inv30 = 1;
    17: op1_08_inv30 = 1;
    18: op1_08_inv30 = 1;
    19: op1_08_inv30 = 1;
    20: op1_08_inv30 = 1;
    21: op1_08_inv30 = 1;
    23: op1_08_inv30 = 1;
    25: op1_08_inv30 = 1;
    27: op1_08_inv30 = 1;
    28: op1_08_inv30 = 1;
    32: op1_08_inv30 = 1;
    34: op1_08_inv30 = 1;
    36: op1_08_inv30 = 1;
    38: op1_08_inv30 = 1;
    46: op1_08_inv30 = 1;
    47: op1_08_inv30 = 1;
    49: op1_08_inv30 = 1;
    51: op1_08_inv30 = 1;
    54: op1_08_inv30 = 1;
    55: op1_08_inv30 = 1;
    57: op1_08_inv30 = 1;
    59: op1_08_inv30 = 1;
    63: op1_08_inv30 = 1;
    65: op1_08_inv30 = 1;
    69: op1_08_inv30 = 1;
    70: op1_08_inv30 = 1;
    71: op1_08_inv30 = 1;
    72: op1_08_inv30 = 1;
    73: op1_08_inv30 = 1;
    74: op1_08_inv30 = 1;
    78: op1_08_inv30 = 1;
    80: op1_08_inv30 = 1;
    82: op1_08_inv30 = 1;
    83: op1_08_inv30 = 1;
    87: op1_08_inv30 = 1;
    89: op1_08_inv30 = 1;
    93: op1_08_inv30 = 1;
    96: op1_08_inv30 = 1;
    default: op1_08_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_08_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_08_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in00 = imem07_in[43:40];
    5: op1_09_in00 = reg_0217;
    6: op1_09_in00 = imem00_in[79:76];
    7: op1_09_in00 = reg_0570;
    8: op1_09_in00 = reg_0623;
    9: op1_09_in00 = reg_0297;
    10: op1_09_in00 = imem00_in[35:32];
    53: op1_09_in00 = imem00_in[35:32];
    11: op1_09_in00 = reg_0292;
    12: op1_09_in00 = reg_0237;
    13: op1_09_in00 = reg_0085;
    14: op1_09_in00 = reg_0078;
    15: op1_09_in00 = imem00_in[31:28];
    40: op1_09_in00 = imem00_in[31:28];
    3: op1_09_in00 = imem07_in[79:76];
    16: op1_09_in00 = reg_0243;
    17: op1_09_in00 = imem00_in[15:12];
    86: op1_09_in00 = imem00_in[15:12];
    88: op1_09_in00 = imem00_in[15:12];
    18: op1_09_in00 = reg_0235;
    19: op1_09_in00 = imem00_in[19:16];
    20: op1_09_in00 = reg_0238;
    21: op1_09_in00 = reg_0028;
    22: op1_09_in00 = reg_0747;
    23: op1_09_in00 = reg_0631;
    2: op1_09_in00 = imem07_in[123:120];
    24: op1_09_in00 = imem00_in[39:36];
    25: op1_09_in00 = reg_0019;
    26: op1_09_in00 = imem00_in[59:56];
    27: op1_09_in00 = reg_0106;
    1: op1_09_in00 = imem07_in[51:48];
    28: op1_09_in00 = imem00_in[7:4];
    68: op1_09_in00 = imem00_in[7:4];
    95: op1_09_in00 = imem00_in[7:4];
    29: op1_09_in00 = imem00_in[75:72];
    30: op1_09_in00 = reg_0642;
    31: op1_09_in00 = reg_0302;
    32: op1_09_in00 = reg_0744;
    33: op1_09_in00 = imem00_in[11:8];
    52: op1_09_in00 = imem00_in[11:8];
    34: op1_09_in00 = imem04_in[119:116];
    35: op1_09_in00 = imem04_in[87:84];
    36: op1_09_in00 = reg_0789;
    37: op1_09_in00 = reg_0003;
    38: op1_09_in00 = reg_0329;
    39: op1_09_in00 = imem00_in[47:44];
    77: op1_09_in00 = imem00_in[47:44];
    41: op1_09_in00 = reg_0806;
    42: op1_09_in00 = imem05_in[39:36];
    43: op1_09_in00 = reg_0635;
    44: op1_09_in00 = reg_0104;
    45: op1_09_in00 = reg_0564;
    46: op1_09_in00 = reg_0406;
    47: op1_09_in00 = reg_0102;
    48: op1_09_in00 = imem03_in[127:124];
    49: op1_09_in00 = reg_0422;
    50: op1_09_in00 = imem00_in[3:0];
    76: op1_09_in00 = imem00_in[3:0];
    51: op1_09_in00 = reg_0440;
    54: op1_09_in00 = reg_0548;
    55: op1_09_in00 = reg_0637;
    56: op1_09_in00 = imem03_in[11:8];
    57: op1_09_in00 = imem04_in[35:32];
    58: op1_09_in00 = reg_0489;
    59: op1_09_in00 = reg_0278;
    60: op1_09_in00 = imem05_in[31:28];
    61: op1_09_in00 = imem07_in[27:24];
    62: op1_09_in00 = reg_0511;
    63: op1_09_in00 = reg_0216;
    64: op1_09_in00 = imem03_in[59:56];
    65: op1_09_in00 = reg_0392;
    66: op1_09_in00 = reg_0396;
    67: op1_09_in00 = imem06_in[127:124];
    69: op1_09_in00 = reg_0087;
    70: op1_09_in00 = imem05_in[115:112];
    71: op1_09_in00 = reg_0603;
    72: op1_09_in00 = imem04_in[15:12];
    91: op1_09_in00 = imem04_in[15:12];
    73: op1_09_in00 = reg_0395;
    74: op1_09_in00 = reg_0150;
    75: op1_09_in00 = reg_0164;
    78: op1_09_in00 = reg_0567;
    79: op1_09_in00 = reg_0544;
    80: op1_09_in00 = reg_0113;
    81: op1_09_in00 = reg_0331;
    82: op1_09_in00 = reg_0119;
    83: op1_09_in00 = reg_0763;
    84: op1_09_in00 = reg_0403;
    85: op1_09_in00 = reg_0128;
    87: op1_09_in00 = imem02_in[87:84];
    89: op1_09_in00 = reg_0588;
    90: op1_09_in00 = reg_0356;
    92: op1_09_in00 = imem07_in[31:28];
    93: op1_09_in00 = reg_0370;
    94: op1_09_in00 = imem06_in[91:88];
    96: op1_09_in00 = reg_0782;
    default: op1_09_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_09_inv00 = 1;
    6: op1_09_inv00 = 1;
    11: op1_09_inv00 = 1;
    13: op1_09_inv00 = 1;
    15: op1_09_inv00 = 1;
    18: op1_09_inv00 = 1;
    19: op1_09_inv00 = 1;
    24: op1_09_inv00 = 1;
    28: op1_09_inv00 = 1;
    30: op1_09_inv00 = 1;
    35: op1_09_inv00 = 1;
    37: op1_09_inv00 = 1;
    38: op1_09_inv00 = 1;
    40: op1_09_inv00 = 1;
    41: op1_09_inv00 = 1;
    42: op1_09_inv00 = 1;
    44: op1_09_inv00 = 1;
    49: op1_09_inv00 = 1;
    50: op1_09_inv00 = 1;
    51: op1_09_inv00 = 1;
    54: op1_09_inv00 = 1;
    55: op1_09_inv00 = 1;
    56: op1_09_inv00 = 1;
    58: op1_09_inv00 = 1;
    59: op1_09_inv00 = 1;
    61: op1_09_inv00 = 1;
    62: op1_09_inv00 = 1;
    63: op1_09_inv00 = 1;
    65: op1_09_inv00 = 1;
    73: op1_09_inv00 = 1;
    74: op1_09_inv00 = 1;
    75: op1_09_inv00 = 1;
    76: op1_09_inv00 = 1;
    78: op1_09_inv00 = 1;
    79: op1_09_inv00 = 1;
    80: op1_09_inv00 = 1;
    82: op1_09_inv00 = 1;
    85: op1_09_inv00 = 1;
    91: op1_09_inv00 = 1;
    93: op1_09_inv00 = 1;
    94: op1_09_inv00 = 1;
    95: op1_09_inv00 = 1;
    96: op1_09_inv00 = 1;
    default: op1_09_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in01 = imem07_in[115:112];
    5: op1_09_in01 = reg_0269;
    6: op1_09_in01 = imem00_in[87:84];
    7: op1_09_in01 = reg_0311;
    8: op1_09_in01 = reg_0348;
    9: op1_09_in01 = reg_0275;
    11: op1_09_in01 = reg_0275;
    58: op1_09_in01 = reg_0275;
    10: op1_09_in01 = imem00_in[75:72];
    26: op1_09_in01 = imem00_in[75:72];
    12: op1_09_in01 = reg_0238;
    13: op1_09_in01 = reg_0096;
    14: op1_09_in01 = reg_0065;
    15: op1_09_in01 = imem00_in[39:36];
    17: op1_09_in01 = imem00_in[39:36];
    19: op1_09_in01 = imem00_in[39:36];
    53: op1_09_in01 = imem00_in[39:36];
    88: op1_09_in01 = imem00_in[39:36];
    3: op1_09_in01 = imem07_in[91:88];
    16: op1_09_in01 = reg_0122;
    18: op1_09_in01 = reg_0246;
    20: op1_09_in01 = reg_0114;
    21: op1_09_in01 = reg_0815;
    22: op1_09_in01 = reg_0813;
    23: op1_09_in01 = reg_0608;
    2: op1_09_in01 = reg_0174;
    24: op1_09_in01 = imem00_in[71:68];
    25: op1_09_in01 = reg_0804;
    27: op1_09_in01 = reg_0110;
    1: op1_09_in01 = imem07_in[99:96];
    28: op1_09_in01 = imem00_in[27:24];
    76: op1_09_in01 = imem00_in[27:24];
    29: op1_09_in01 = imem00_in[99:96];
    30: op1_09_in01 = reg_0661;
    31: op1_09_in01 = reg_0290;
    78: op1_09_in01 = reg_0290;
    32: op1_09_in01 = reg_0135;
    33: op1_09_in01 = reg_0693;
    34: op1_09_in01 = reg_0542;
    35: op1_09_in01 = imem04_in[107:104];
    36: op1_09_in01 = reg_0491;
    37: op1_09_in01 = reg_0800;
    38: op1_09_in01 = reg_0028;
    73: op1_09_in01 = reg_0028;
    39: op1_09_in01 = imem00_in[51:48];
    40: op1_09_in01 = imem00_in[47:44];
    41: op1_09_in01 = reg_0239;
    42: op1_09_in01 = imem05_in[51:48];
    43: op1_09_in01 = reg_0446;
    44: op1_09_in01 = reg_0119;
    45: op1_09_in01 = reg_0000;
    46: op1_09_in01 = reg_0038;
    47: op1_09_in01 = reg_0107;
    48: op1_09_in01 = reg_0588;
    49: op1_09_in01 = reg_0574;
    50: op1_09_in01 = imem00_in[11:8];
    51: op1_09_in01 = reg_0438;
    52: op1_09_in01 = imem00_in[31:28];
    54: op1_09_in01 = reg_0665;
    96: op1_09_in01 = reg_0665;
    55: op1_09_in01 = reg_0426;
    56: op1_09_in01 = imem03_in[23:20];
    57: op1_09_in01 = imem04_in[43:40];
    59: op1_09_in01 = reg_0752;
    60: op1_09_in01 = imem05_in[115:112];
    61: op1_09_in01 = imem07_in[39:36];
    62: op1_09_in01 = reg_0054;
    63: op1_09_in01 = reg_0234;
    64: op1_09_in01 = imem03_in[83:80];
    65: op1_09_in01 = reg_0802;
    66: op1_09_in01 = reg_0570;
    67: op1_09_in01 = reg_0354;
    68: op1_09_in01 = imem00_in[35:32];
    69: op1_09_in01 = reg_0537;
    70: op1_09_in01 = reg_0793;
    71: op1_09_in01 = reg_0506;
    72: op1_09_in01 = imem04_in[23:20];
    74: op1_09_in01 = reg_0152;
    75: op1_09_in01 = reg_0185;
    77: op1_09_in01 = imem00_in[67:64];
    79: op1_09_in01 = reg_0560;
    80: op1_09_in01 = reg_0732;
    81: op1_09_in01 = reg_0321;
    82: op1_09_in01 = reg_0672;
    83: op1_09_in01 = reg_0270;
    84: op1_09_in01 = reg_0490;
    85: op1_09_in01 = reg_0489;
    86: op1_09_in01 = imem00_in[43:40];
    87: op1_09_in01 = imem02_in[123:120];
    89: op1_09_in01 = reg_0006;
    90: op1_09_in01 = reg_0342;
    91: op1_09_in01 = imem04_in[35:32];
    92: op1_09_in01 = imem07_in[51:48];
    93: op1_09_in01 = reg_0409;
    94: op1_09_in01 = imem06_in[107:104];
    95: op1_09_in01 = imem00_in[19:16];
    default: op1_09_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_09_inv01 = 1;
    5: op1_09_inv01 = 1;
    7: op1_09_inv01 = 1;
    14: op1_09_inv01 = 1;
    3: op1_09_inv01 = 1;
    16: op1_09_inv01 = 1;
    17: op1_09_inv01 = 1;
    19: op1_09_inv01 = 1;
    2: op1_09_inv01 = 1;
    24: op1_09_inv01 = 1;
    26: op1_09_inv01 = 1;
    27: op1_09_inv01 = 1;
    29: op1_09_inv01 = 1;
    32: op1_09_inv01 = 1;
    34: op1_09_inv01 = 1;
    36: op1_09_inv01 = 1;
    37: op1_09_inv01 = 1;
    39: op1_09_inv01 = 1;
    40: op1_09_inv01 = 1;
    41: op1_09_inv01 = 1;
    43: op1_09_inv01 = 1;
    44: op1_09_inv01 = 1;
    47: op1_09_inv01 = 1;
    48: op1_09_inv01 = 1;
    49: op1_09_inv01 = 1;
    51: op1_09_inv01 = 1;
    52: op1_09_inv01 = 1;
    53: op1_09_inv01 = 1;
    55: op1_09_inv01 = 1;
    56: op1_09_inv01 = 1;
    57: op1_09_inv01 = 1;
    58: op1_09_inv01 = 1;
    60: op1_09_inv01 = 1;
    61: op1_09_inv01 = 1;
    62: op1_09_inv01 = 1;
    64: op1_09_inv01 = 1;
    68: op1_09_inv01 = 1;
    69: op1_09_inv01 = 1;
    70: op1_09_inv01 = 1;
    71: op1_09_inv01 = 1;
    72: op1_09_inv01 = 1;
    74: op1_09_inv01 = 1;
    75: op1_09_inv01 = 1;
    80: op1_09_inv01 = 1;
    84: op1_09_inv01 = 1;
    86: op1_09_inv01 = 1;
    87: op1_09_inv01 = 1;
    90: op1_09_inv01 = 1;
    91: op1_09_inv01 = 1;
    93: op1_09_inv01 = 1;
    94: op1_09_inv01 = 1;
    96: op1_09_inv01 = 1;
    default: op1_09_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in02 = imem07_in[127:124];
    5: op1_09_in02 = reg_0263;
    6: op1_09_in02 = imem00_in[91:88];
    7: op1_09_in02 = reg_0376;
    8: op1_09_in02 = reg_0313;
    9: op1_09_in02 = reg_0065;
    10: op1_09_in02 = imem00_in[83:80];
    11: op1_09_in02 = reg_0054;
    12: op1_09_in02 = reg_0111;
    13: op1_09_in02 = reg_0097;
    14: op1_09_in02 = reg_0048;
    15: op1_09_in02 = imem00_in[47:44];
    17: op1_09_in02 = imem00_in[47:44];
    86: op1_09_in02 = imem00_in[47:44];
    3: op1_09_in02 = imem07_in[99:96];
    16: op1_09_in02 = reg_0116;
    18: op1_09_in02 = reg_0217;
    19: op1_09_in02 = imem00_in[55:52];
    40: op1_09_in02 = imem00_in[55:52];
    53: op1_09_in02 = imem00_in[55:52];
    20: op1_09_in02 = reg_0109;
    21: op1_09_in02 = reg_0040;
    22: op1_09_in02 = reg_0035;
    23: op1_09_in02 = reg_0632;
    2: op1_09_in02 = reg_0161;
    24: op1_09_in02 = imem00_in[99:96];
    25: op1_09_in02 = reg_0801;
    26: op1_09_in02 = imem00_in[115:112];
    27: op1_09_in02 = imem02_in[19:16];
    28: op1_09_in02 = imem00_in[35:32];
    95: op1_09_in02 = imem00_in[35:32];
    29: op1_09_in02 = reg_0682;
    30: op1_09_in02 = reg_0656;
    31: op1_09_in02 = reg_0267;
    32: op1_09_in02 = reg_0139;
    33: op1_09_in02 = reg_0694;
    34: op1_09_in02 = reg_0055;
    35: op1_09_in02 = reg_0328;
    36: op1_09_in02 = reg_0780;
    37: op1_09_in02 = reg_0806;
    38: op1_09_in02 = reg_0031;
    39: op1_09_in02 = imem00_in[71:68];
    41: op1_09_in02 = reg_0049;
    42: op1_09_in02 = imem05_in[71:68];
    43: op1_09_in02 = reg_0440;
    44: op1_09_in02 = reg_0100;
    45: op1_09_in02 = reg_0012;
    46: op1_09_in02 = reg_0028;
    47: op1_09_in02 = imem02_in[43:40];
    48: op1_09_in02 = reg_0749;
    49: op1_09_in02 = reg_0567;
    50: op1_09_in02 = imem00_in[19:16];
    51: op1_09_in02 = reg_0268;
    52: op1_09_in02 = imem00_in[59:56];
    54: op1_09_in02 = reg_0659;
    55: op1_09_in02 = reg_0362;
    56: op1_09_in02 = imem03_in[51:48];
    57: op1_09_in02 = imem04_in[59:56];
    58: op1_09_in02 = reg_0491;
    59: op1_09_in02 = reg_0114;
    60: op1_09_in02 = imem05_in[127:124];
    61: op1_09_in02 = imem07_in[107:104];
    62: op1_09_in02 = reg_0504;
    63: op1_09_in02 = reg_0105;
    64: op1_09_in02 = reg_0602;
    65: op1_09_in02 = reg_0009;
    66: op1_09_in02 = reg_0013;
    67: op1_09_in02 = reg_0402;
    68: op1_09_in02 = imem00_in[51:48];
    69: op1_09_in02 = reg_0056;
    70: op1_09_in02 = reg_0499;
    71: op1_09_in02 = reg_0424;
    72: op1_09_in02 = imem04_in[27:24];
    73: op1_09_in02 = reg_0575;
    74: op1_09_in02 = reg_0156;
    76: op1_09_in02 = imem00_in[43:40];
    77: op1_09_in02 = imem00_in[119:116];
    88: op1_09_in02 = imem00_in[119:116];
    78: op1_09_in02 = reg_0670;
    79: op1_09_in02 = reg_0542;
    80: op1_09_in02 = reg_0489;
    81: op1_09_in02 = reg_0755;
    82: op1_09_in02 = reg_0675;
    83: op1_09_in02 = reg_0638;
    84: op1_09_in02 = reg_0387;
    85: op1_09_in02 = reg_0517;
    87: op1_09_in02 = reg_0264;
    89: op1_09_in02 = reg_0509;
    90: op1_09_in02 = reg_0406;
    91: op1_09_in02 = imem04_in[55:52];
    92: op1_09_in02 = imem07_in[63:60];
    93: op1_09_in02 = reg_0519;
    94: op1_09_in02 = reg_0289;
    96: op1_09_in02 = reg_0134;
    default: op1_09_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_09_inv02 = 1;
    10: op1_09_inv02 = 1;
    11: op1_09_inv02 = 1;
    12: op1_09_inv02 = 1;
    3: op1_09_inv02 = 1;
    16: op1_09_inv02 = 1;
    23: op1_09_inv02 = 1;
    2: op1_09_inv02 = 1;
    25: op1_09_inv02 = 1;
    27: op1_09_inv02 = 1;
    29: op1_09_inv02 = 1;
    31: op1_09_inv02 = 1;
    34: op1_09_inv02 = 1;
    35: op1_09_inv02 = 1;
    39: op1_09_inv02 = 1;
    40: op1_09_inv02 = 1;
    41: op1_09_inv02 = 1;
    42: op1_09_inv02 = 1;
    44: op1_09_inv02 = 1;
    46: op1_09_inv02 = 1;
    50: op1_09_inv02 = 1;
    52: op1_09_inv02 = 1;
    54: op1_09_inv02 = 1;
    55: op1_09_inv02 = 1;
    56: op1_09_inv02 = 1;
    58: op1_09_inv02 = 1;
    59: op1_09_inv02 = 1;
    60: op1_09_inv02 = 1;
    65: op1_09_inv02 = 1;
    67: op1_09_inv02 = 1;
    70: op1_09_inv02 = 1;
    72: op1_09_inv02 = 1;
    73: op1_09_inv02 = 1;
    74: op1_09_inv02 = 1;
    79: op1_09_inv02 = 1;
    80: op1_09_inv02 = 1;
    81: op1_09_inv02 = 1;
    82: op1_09_inv02 = 1;
    86: op1_09_inv02 = 1;
    87: op1_09_inv02 = 1;
    93: op1_09_inv02 = 1;
    94: op1_09_inv02 = 1;
    default: op1_09_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in03 = reg_0719;
    5: op1_09_in03 = reg_0149;
    6: op1_09_in03 = imem00_in[103:100];
    7: op1_09_in03 = reg_0013;
    8: op1_09_in03 = imem06_in[27:24];
    9: op1_09_in03 = reg_0058;
    20: op1_09_in03 = reg_0058;
    10: op1_09_in03 = imem00_in[111:108];
    68: op1_09_in03 = imem00_in[111:108];
    11: op1_09_in03 = reg_0065;
    12: op1_09_in03 = reg_0116;
    13: op1_09_in03 = reg_0087;
    14: op1_09_in03 = reg_0050;
    15: op1_09_in03 = imem00_in[79:76];
    17: op1_09_in03 = imem00_in[79:76];
    3: op1_09_in03 = imem07_in[115:112];
    16: op1_09_in03 = reg_0120;
    63: op1_09_in03 = reg_0120;
    18: op1_09_in03 = reg_0244;
    19: op1_09_in03 = imem00_in[91:88];
    21: op1_09_in03 = imem07_in[19:16];
    22: op1_09_in03 = reg_0040;
    23: op1_09_in03 = reg_0332;
    2: op1_09_in03 = reg_0162;
    24: op1_09_in03 = imem00_in[123:120];
    25: op1_09_in03 = reg_0799;
    26: op1_09_in03 = imem00_in[127:124];
    39: op1_09_in03 = imem00_in[127:124];
    27: op1_09_in03 = imem02_in[47:44];
    47: op1_09_in03 = imem02_in[47:44];
    28: op1_09_in03 = imem00_in[67:64];
    53: op1_09_in03 = imem00_in[67:64];
    29: op1_09_in03 = reg_0693;
    30: op1_09_in03 = reg_0641;
    31: op1_09_in03 = reg_0286;
    32: op1_09_in03 = imem06_in[3:0];
    33: op1_09_in03 = reg_0689;
    34: op1_09_in03 = reg_0083;
    35: op1_09_in03 = reg_0555;
    36: op1_09_in03 = reg_0790;
    37: op1_09_in03 = reg_0010;
    38: op1_09_in03 = reg_0815;
    40: op1_09_in03 = imem00_in[83:80];
    52: op1_09_in03 = imem00_in[83:80];
    41: op1_09_in03 = reg_0084;
    42: op1_09_in03 = imem05_in[79:76];
    43: op1_09_in03 = reg_0442;
    44: op1_09_in03 = reg_0113;
    45: op1_09_in03 = reg_0007;
    46: op1_09_in03 = reg_0753;
    48: op1_09_in03 = reg_0373;
    49: op1_09_in03 = reg_0240;
    50: op1_09_in03 = imem00_in[35:32];
    51: op1_09_in03 = reg_0174;
    54: op1_09_in03 = reg_0427;
    55: op1_09_in03 = reg_0320;
    56: op1_09_in03 = imem03_in[71:68];
    57: op1_09_in03 = imem04_in[79:76];
    58: op1_09_in03 = reg_0088;
    79: op1_09_in03 = reg_0088;
    59: op1_09_in03 = reg_0090;
    60: op1_09_in03 = reg_0090;
    61: op1_09_in03 = reg_0726;
    62: op1_09_in03 = reg_0670;
    64: op1_09_in03 = reg_0604;
    89: op1_09_in03 = reg_0604;
    65: op1_09_in03 = reg_0004;
    66: op1_09_in03 = reg_0807;
    67: op1_09_in03 = reg_0654;
    69: op1_09_in03 = reg_0558;
    70: op1_09_in03 = reg_0389;
    71: op1_09_in03 = reg_0420;
    72: op1_09_in03 = imem04_in[59:56];
    73: op1_09_in03 = reg_0387;
    74: op1_09_in03 = reg_0143;
    76: op1_09_in03 = imem00_in[87:84];
    77: op1_09_in03 = reg_0696;
    78: op1_09_in03 = reg_0119;
    80: op1_09_in03 = reg_0315;
    81: op1_09_in03 = reg_0368;
    82: op1_09_in03 = reg_0669;
    83: op1_09_in03 = reg_0039;
    84: op1_09_in03 = reg_0623;
    85: op1_09_in03 = reg_0252;
    86: op1_09_in03 = imem00_in[99:96];
    87: op1_09_in03 = reg_0647;
    88: op1_09_in03 = reg_0697;
    90: op1_09_in03 = reg_0092;
    91: op1_09_in03 = imem04_in[63:60];
    92: op1_09_in03 = imem07_in[71:68];
    93: op1_09_in03 = reg_0578;
    94: op1_09_in03 = reg_0370;
    95: op1_09_in03 = imem00_in[43:40];
    96: op1_09_in03 = reg_0517;
    default: op1_09_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv03 = 1;
    6: op1_09_inv03 = 1;
    8: op1_09_inv03 = 1;
    10: op1_09_inv03 = 1;
    12: op1_09_inv03 = 1;
    13: op1_09_inv03 = 1;
    14: op1_09_inv03 = 1;
    15: op1_09_inv03 = 1;
    21: op1_09_inv03 = 1;
    2: op1_09_inv03 = 1;
    24: op1_09_inv03 = 1;
    28: op1_09_inv03 = 1;
    31: op1_09_inv03 = 1;
    33: op1_09_inv03 = 1;
    34: op1_09_inv03 = 1;
    37: op1_09_inv03 = 1;
    38: op1_09_inv03 = 1;
    39: op1_09_inv03 = 1;
    41: op1_09_inv03 = 1;
    42: op1_09_inv03 = 1;
    43: op1_09_inv03 = 1;
    45: op1_09_inv03 = 1;
    46: op1_09_inv03 = 1;
    48: op1_09_inv03 = 1;
    49: op1_09_inv03 = 1;
    50: op1_09_inv03 = 1;
    53: op1_09_inv03 = 1;
    54: op1_09_inv03 = 1;
    57: op1_09_inv03 = 1;
    58: op1_09_inv03 = 1;
    59: op1_09_inv03 = 1;
    61: op1_09_inv03 = 1;
    62: op1_09_inv03 = 1;
    63: op1_09_inv03 = 1;
    70: op1_09_inv03 = 1;
    73: op1_09_inv03 = 1;
    77: op1_09_inv03 = 1;
    78: op1_09_inv03 = 1;
    82: op1_09_inv03 = 1;
    84: op1_09_inv03 = 1;
    86: op1_09_inv03 = 1;
    87: op1_09_inv03 = 1;
    89: op1_09_inv03 = 1;
    91: op1_09_inv03 = 1;
    92: op1_09_inv03 = 1;
    93: op1_09_inv03 = 1;
    96: op1_09_inv03 = 1;
    default: op1_09_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in04 = reg_0720;
    80: op1_09_in04 = reg_0720;
    5: op1_09_in04 = reg_0150;
    6: op1_09_in04 = reg_0682;
    86: op1_09_in04 = reg_0682;
    7: op1_09_in04 = reg_0800;
    8: op1_09_in04 = imem07_in[39:36];
    9: op1_09_in04 = reg_0068;
    10: op1_09_in04 = reg_0685;
    11: op1_09_in04 = reg_0048;
    12: op1_09_in04 = reg_0113;
    13: op1_09_in04 = reg_0094;
    14: op1_09_in04 = imem05_in[39:36];
    15: op1_09_in04 = imem00_in[87:84];
    3: op1_09_in04 = reg_0422;
    16: op1_09_in04 = reg_0114;
    17: op1_09_in04 = imem00_in[95:92];
    40: op1_09_in04 = imem00_in[95:92];
    18: op1_09_in04 = reg_0041;
    19: op1_09_in04 = imem00_in[99:96];
    52: op1_09_in04 = imem00_in[99:96];
    20: op1_09_in04 = reg_0059;
    21: op1_09_in04 = imem07_in[59:56];
    22: op1_09_in04 = reg_0819;
    23: op1_09_in04 = reg_0381;
    2: op1_09_in04 = reg_0184;
    24: op1_09_in04 = reg_0693;
    25: op1_09_in04 = reg_0016;
    45: op1_09_in04 = reg_0016;
    26: op1_09_in04 = reg_0672;
    27: op1_09_in04 = imem02_in[51:48];
    28: op1_09_in04 = imem00_in[75:72];
    29: op1_09_in04 = reg_0697;
    39: op1_09_in04 = reg_0697;
    30: op1_09_in04 = reg_0636;
    31: op1_09_in04 = reg_0051;
    32: op1_09_in04 = imem06_in[87:84];
    33: op1_09_in04 = reg_0677;
    34: op1_09_in04 = reg_0057;
    58: op1_09_in04 = reg_0057;
    35: op1_09_in04 = reg_0551;
    36: op1_09_in04 = reg_0737;
    37: op1_09_in04 = imem04_in[11:8];
    38: op1_09_in04 = reg_0375;
    41: op1_09_in04 = reg_0328;
    42: op1_09_in04 = imem05_in[87:84];
    43: op1_09_in04 = reg_0437;
    44: op1_09_in04 = reg_0645;
    46: op1_09_in04 = reg_0620;
    47: op1_09_in04 = imem02_in[55:52];
    48: op1_09_in04 = reg_0572;
    49: op1_09_in04 = reg_0220;
    50: op1_09_in04 = imem00_in[43:40];
    51: op1_09_in04 = reg_0175;
    53: op1_09_in04 = imem00_in[83:80];
    54: op1_09_in04 = reg_0586;
    55: op1_09_in04 = reg_0586;
    56: op1_09_in04 = imem03_in[95:92];
    57: op1_09_in04 = imem04_in[91:88];
    59: op1_09_in04 = reg_0099;
    60: op1_09_in04 = reg_0276;
    61: op1_09_in04 = reg_0725;
    62: op1_09_in04 = reg_0592;
    63: op1_09_in04 = reg_0126;
    64: op1_09_in04 = reg_0596;
    65: op1_09_in04 = imem04_in[7:4];
    66: op1_09_in04 = reg_0801;
    67: op1_09_in04 = reg_0377;
    68: op1_09_in04 = reg_0689;
    69: op1_09_in04 = reg_0556;
    70: op1_09_in04 = reg_0215;
    71: op1_09_in04 = reg_0105;
    72: op1_09_in04 = imem04_in[95:92];
    73: op1_09_in04 = reg_0747;
    74: op1_09_in04 = reg_0828;
    76: op1_09_in04 = imem00_in[127:124];
    77: op1_09_in04 = reg_0686;
    78: op1_09_in04 = reg_0120;
    79: op1_09_in04 = reg_0283;
    81: op1_09_in04 = reg_0646;
    82: op1_09_in04 = reg_0601;
    83: op1_09_in04 = reg_0652;
    84: op1_09_in04 = reg_0649;
    85: op1_09_in04 = reg_0491;
    87: op1_09_in04 = reg_0485;
    88: op1_09_in04 = reg_0696;
    89: op1_09_in04 = reg_0559;
    90: op1_09_in04 = reg_0043;
    91: op1_09_in04 = reg_0553;
    92: op1_09_in04 = imem07_in[83:80];
    93: op1_09_in04 = reg_0408;
    94: op1_09_in04 = reg_0339;
    95: op1_09_in04 = imem00_in[47:44];
    96: op1_09_in04 = reg_0309;
    default: op1_09_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv04 = 1;
    11: op1_09_inv04 = 1;
    15: op1_09_inv04 = 1;
    16: op1_09_inv04 = 1;
    19: op1_09_inv04 = 1;
    23: op1_09_inv04 = 1;
    2: op1_09_inv04 = 1;
    24: op1_09_inv04 = 1;
    27: op1_09_inv04 = 1;
    30: op1_09_inv04 = 1;
    33: op1_09_inv04 = 1;
    34: op1_09_inv04 = 1;
    35: op1_09_inv04 = 1;
    38: op1_09_inv04 = 1;
    39: op1_09_inv04 = 1;
    41: op1_09_inv04 = 1;
    42: op1_09_inv04 = 1;
    46: op1_09_inv04 = 1;
    50: op1_09_inv04 = 1;
    51: op1_09_inv04 = 1;
    52: op1_09_inv04 = 1;
    53: op1_09_inv04 = 1;
    54: op1_09_inv04 = 1;
    55: op1_09_inv04 = 1;
    56: op1_09_inv04 = 1;
    59: op1_09_inv04 = 1;
    64: op1_09_inv04 = 1;
    67: op1_09_inv04 = 1;
    68: op1_09_inv04 = 1;
    69: op1_09_inv04 = 1;
    70: op1_09_inv04 = 1;
    71: op1_09_inv04 = 1;
    72: op1_09_inv04 = 1;
    73: op1_09_inv04 = 1;
    76: op1_09_inv04 = 1;
    77: op1_09_inv04 = 1;
    78: op1_09_inv04 = 1;
    80: op1_09_inv04 = 1;
    83: op1_09_inv04 = 1;
    84: op1_09_inv04 = 1;
    87: op1_09_inv04 = 1;
    90: op1_09_inv04 = 1;
    91: op1_09_inv04 = 1;
    93: op1_09_inv04 = 1;
    95: op1_09_inv04 = 1;
    default: op1_09_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in05 = reg_0721;
    5: op1_09_in05 = reg_0152;
    6: op1_09_in05 = reg_0684;
    88: op1_09_in05 = reg_0684;
    7: op1_09_in05 = reg_0805;
    8: op1_09_in05 = imem07_in[123:120];
    9: op1_09_in05 = reg_0048;
    10: op1_09_in05 = reg_0688;
    11: op1_09_in05 = reg_0254;
    12: op1_09_in05 = imem02_in[3:0];
    13: op1_09_in05 = imem03_in[7:4];
    14: op1_09_in05 = imem05_in[75:72];
    15: op1_09_in05 = imem00_in[107:104];
    3: op1_09_in05 = reg_0423;
    16: op1_09_in05 = reg_0127;
    17: op1_09_in05 = reg_0693;
    19: op1_09_in05 = reg_0693;
    18: op1_09_in05 = reg_0238;
    20: op1_09_in05 = reg_0666;
    21: op1_09_in05 = imem07_in[67:64];
    22: op1_09_in05 = reg_0816;
    23: op1_09_in05 = reg_0390;
    24: op1_09_in05 = reg_0689;
    25: op1_09_in05 = reg_0806;
    26: op1_09_in05 = reg_0670;
    27: op1_09_in05 = imem02_in[55:52];
    28: op1_09_in05 = imem00_in[99:96];
    50: op1_09_in05 = imem00_in[99:96];
    53: op1_09_in05 = imem00_in[99:96];
    29: op1_09_in05 = reg_0683;
    39: op1_09_in05 = reg_0683;
    30: op1_09_in05 = reg_0341;
    31: op1_09_in05 = reg_0257;
    32: op1_09_in05 = imem06_in[95:92];
    33: op1_09_in05 = reg_0678;
    82: op1_09_in05 = reg_0678;
    34: op1_09_in05 = reg_0295;
    35: op1_09_in05 = reg_0052;
    36: op1_09_in05 = reg_0149;
    37: op1_09_in05 = imem04_in[15:12];
    38: op1_09_in05 = reg_0752;
    40: op1_09_in05 = reg_0697;
    41: op1_09_in05 = imem04_in[7:4];
    42: op1_09_in05 = reg_0792;
    43: op1_09_in05 = reg_0438;
    44: op1_09_in05 = imem02_in[11:8];
    45: op1_09_in05 = reg_0245;
    46: op1_09_in05 = reg_0338;
    47: op1_09_in05 = reg_0650;
    48: op1_09_in05 = reg_0811;
    49: op1_09_in05 = reg_0603;
    51: op1_09_in05 = reg_0165;
    52: op1_09_in05 = reg_0695;
    54: op1_09_in05 = reg_0351;
    55: op1_09_in05 = reg_0594;
    56: op1_09_in05 = imem03_in[111:108];
    57: op1_09_in05 = imem04_in[127:124];
    58: op1_09_in05 = reg_0058;
    59: op1_09_in05 = reg_0309;
    60: op1_09_in05 = reg_0101;
    61: op1_09_in05 = reg_0729;
    62: op1_09_in05 = reg_0675;
    63: op1_09_in05 = imem02_in[27:24];
    64: op1_09_in05 = reg_0350;
    65: op1_09_in05 = imem04_in[43:40];
    66: op1_09_in05 = reg_0014;
    73: op1_09_in05 = reg_0014;
    67: op1_09_in05 = reg_0580;
    68: op1_09_in05 = reg_0691;
    69: op1_09_in05 = reg_0432;
    70: op1_09_in05 = reg_0797;
    71: op1_09_in05 = reg_0124;
    72: op1_09_in05 = reg_0560;
    74: op1_09_in05 = imem06_in[63:60];
    76: op1_09_in05 = reg_0696;
    77: op1_09_in05 = reg_0451;
    78: op1_09_in05 = reg_0671;
    79: op1_09_in05 = reg_0050;
    80: op1_09_in05 = reg_0393;
    81: op1_09_in05 = reg_0496;
    83: op1_09_in05 = reg_0787;
    84: op1_09_in05 = reg_0012;
    85: op1_09_in05 = reg_0277;
    86: op1_09_in05 = reg_0681;
    87: op1_09_in05 = reg_0359;
    89: op1_09_in05 = reg_0801;
    90: op1_09_in05 = reg_0109;
    91: op1_09_in05 = reg_0177;
    92: op1_09_in05 = imem07_in[95:92];
    93: op1_09_in05 = reg_0613;
    94: op1_09_in05 = reg_0293;
    95: op1_09_in05 = imem00_in[63:60];
    96: op1_09_in05 = reg_0830;
    default: op1_09_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv05 = 1;
    6: op1_09_inv05 = 1;
    8: op1_09_inv05 = 1;
    9: op1_09_inv05 = 1;
    11: op1_09_inv05 = 1;
    12: op1_09_inv05 = 1;
    13: op1_09_inv05 = 1;
    15: op1_09_inv05 = 1;
    16: op1_09_inv05 = 1;
    17: op1_09_inv05 = 1;
    19: op1_09_inv05 = 1;
    20: op1_09_inv05 = 1;
    21: op1_09_inv05 = 1;
    22: op1_09_inv05 = 1;
    23: op1_09_inv05 = 1;
    24: op1_09_inv05 = 1;
    25: op1_09_inv05 = 1;
    26: op1_09_inv05 = 1;
    28: op1_09_inv05 = 1;
    30: op1_09_inv05 = 1;
    32: op1_09_inv05 = 1;
    34: op1_09_inv05 = 1;
    36: op1_09_inv05 = 1;
    39: op1_09_inv05 = 1;
    42: op1_09_inv05 = 1;
    46: op1_09_inv05 = 1;
    49: op1_09_inv05 = 1;
    51: op1_09_inv05 = 1;
    54: op1_09_inv05 = 1;
    55: op1_09_inv05 = 1;
    57: op1_09_inv05 = 1;
    58: op1_09_inv05 = 1;
    59: op1_09_inv05 = 1;
    60: op1_09_inv05 = 1;
    63: op1_09_inv05 = 1;
    64: op1_09_inv05 = 1;
    65: op1_09_inv05 = 1;
    68: op1_09_inv05 = 1;
    69: op1_09_inv05 = 1;
    71: op1_09_inv05 = 1;
    73: op1_09_inv05 = 1;
    76: op1_09_inv05 = 1;
    77: op1_09_inv05 = 1;
    78: op1_09_inv05 = 1;
    80: op1_09_inv05 = 1;
    82: op1_09_inv05 = 1;
    83: op1_09_inv05 = 1;
    84: op1_09_inv05 = 1;
    88: op1_09_inv05 = 1;
    89: op1_09_inv05 = 1;
    92: op1_09_inv05 = 1;
    93: op1_09_inv05 = 1;
    96: op1_09_inv05 = 1;
    default: op1_09_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in06 = reg_0702;
    5: op1_09_in06 = reg_0141;
    6: op1_09_in06 = reg_0450;
    7: op1_09_in06 = reg_0008;
    8: op1_09_in06 = reg_0710;
    9: op1_09_in06 = imem05_in[55:52];
    10: op1_09_in06 = reg_0463;
    11: op1_09_in06 = reg_0253;
    12: op1_09_in06 = imem02_in[43:40];
    13: op1_09_in06 = imem03_in[11:8];
    14: op1_09_in06 = imem05_in[87:84];
    15: op1_09_in06 = reg_0685;
    76: op1_09_in06 = reg_0685;
    3: op1_09_in06 = reg_0445;
    16: op1_09_in06 = reg_0113;
    17: op1_09_in06 = reg_0697;
    18: op1_09_in06 = reg_0508;
    19: op1_09_in06 = reg_0694;
    20: op1_09_in06 = reg_0639;
    21: op1_09_in06 = imem07_in[111:108];
    22: op1_09_in06 = reg_0036;
    23: op1_09_in06 = reg_0032;
    24: op1_09_in06 = reg_0686;
    29: op1_09_in06 = reg_0686;
    25: op1_09_in06 = reg_0004;
    26: op1_09_in06 = reg_0688;
    27: op1_09_in06 = imem02_in[59:56];
    28: op1_09_in06 = imem00_in[115:112];
    30: op1_09_in06 = reg_0345;
    31: op1_09_in06 = reg_0078;
    32: op1_09_in06 = reg_0614;
    33: op1_09_in06 = reg_0687;
    34: op1_09_in06 = reg_0061;
    35: op1_09_in06 = reg_0291;
    36: op1_09_in06 = reg_0145;
    37: op1_09_in06 = imem04_in[27:24];
    38: op1_09_in06 = imem07_in[31:28];
    39: op1_09_in06 = reg_0696;
    40: op1_09_in06 = reg_0672;
    41: op1_09_in06 = imem04_in[11:8];
    81: op1_09_in06 = imem04_in[11:8];
    42: op1_09_in06 = reg_0797;
    43: op1_09_in06 = reg_0435;
    44: op1_09_in06 = imem02_in[35:32];
    45: op1_09_in06 = reg_0062;
    46: op1_09_in06 = reg_0029;
    47: op1_09_in06 = reg_0666;
    48: op1_09_in06 = reg_0007;
    49: op1_09_in06 = reg_0504;
    50: op1_09_in06 = imem00_in[127:124];
    51: op1_09_in06 = reg_0161;
    52: op1_09_in06 = reg_0683;
    53: op1_09_in06 = imem00_in[107:104];
    54: op1_09_in06 = reg_0365;
    55: op1_09_in06 = reg_0518;
    56: op1_09_in06 = reg_0317;
    57: op1_09_in06 = reg_0328;
    72: op1_09_in06 = reg_0328;
    58: op1_09_in06 = reg_0547;
    59: op1_09_in06 = reg_0103;
    60: op1_09_in06 = reg_0136;
    61: op1_09_in06 = reg_0708;
    62: op1_09_in06 = reg_0676;
    63: op1_09_in06 = imem02_in[39:36];
    64: op1_09_in06 = reg_0488;
    65: op1_09_in06 = imem04_in[87:84];
    66: op1_09_in06 = reg_0806;
    67: op1_09_in06 = reg_0035;
    68: op1_09_in06 = reg_0472;
    69: op1_09_in06 = reg_0305;
    70: op1_09_in06 = reg_0783;
    71: op1_09_in06 = reg_0106;
    73: op1_09_in06 = reg_0016;
    74: op1_09_in06 = imem06_in[67:64];
    77: op1_09_in06 = reg_0457;
    78: op1_09_in06 = reg_0127;
    79: op1_09_in06 = reg_0617;
    80: op1_09_in06 = reg_0383;
    82: op1_09_in06 = imem02_in[11:8];
    83: op1_09_in06 = imem07_in[19:16];
    84: op1_09_in06 = reg_0001;
    85: op1_09_in06 = reg_0149;
    86: op1_09_in06 = reg_0658;
    87: op1_09_in06 = reg_0324;
    88: op1_09_in06 = reg_0749;
    89: op1_09_in06 = reg_0318;
    90: op1_09_in06 = reg_0540;
    91: op1_09_in06 = reg_0539;
    92: op1_09_in06 = imem07_in[103:100];
    93: op1_09_in06 = reg_0763;
    94: op1_09_in06 = reg_0402;
    95: op1_09_in06 = imem00_in[95:92];
    96: op1_09_in06 = reg_0156;
    default: op1_09_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_09_inv06 = 1;
    6: op1_09_inv06 = 1;
    7: op1_09_inv06 = 1;
    8: op1_09_inv06 = 1;
    9: op1_09_inv06 = 1;
    10: op1_09_inv06 = 1;
    12: op1_09_inv06 = 1;
    3: op1_09_inv06 = 1;
    17: op1_09_inv06 = 1;
    18: op1_09_inv06 = 1;
    20: op1_09_inv06 = 1;
    22: op1_09_inv06 = 1;
    23: op1_09_inv06 = 1;
    24: op1_09_inv06 = 1;
    25: op1_09_inv06 = 1;
    27: op1_09_inv06 = 1;
    28: op1_09_inv06 = 1;
    32: op1_09_inv06 = 1;
    36: op1_09_inv06 = 1;
    39: op1_09_inv06 = 1;
    41: op1_09_inv06 = 1;
    44: op1_09_inv06 = 1;
    46: op1_09_inv06 = 1;
    49: op1_09_inv06 = 1;
    51: op1_09_inv06 = 1;
    57: op1_09_inv06 = 1;
    59: op1_09_inv06 = 1;
    61: op1_09_inv06 = 1;
    62: op1_09_inv06 = 1;
    63: op1_09_inv06 = 1;
    64: op1_09_inv06 = 1;
    66: op1_09_inv06 = 1;
    67: op1_09_inv06 = 1;
    68: op1_09_inv06 = 1;
    70: op1_09_inv06 = 1;
    71: op1_09_inv06 = 1;
    76: op1_09_inv06 = 1;
    77: op1_09_inv06 = 1;
    78: op1_09_inv06 = 1;
    79: op1_09_inv06 = 1;
    81: op1_09_inv06 = 1;
    84: op1_09_inv06 = 1;
    85: op1_09_inv06 = 1;
    86: op1_09_inv06 = 1;
    87: op1_09_inv06 = 1;
    88: op1_09_inv06 = 1;
    91: op1_09_inv06 = 1;
    93: op1_09_inv06 = 1;
    94: op1_09_inv06 = 1;
    95: op1_09_inv06 = 1;
    default: op1_09_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in07 = reg_0426;
    5: op1_09_in07 = reg_0130;
    6: op1_09_in07 = reg_0457;
    7: op1_09_in07 = reg_0015;
    8: op1_09_in07 = reg_0725;
    9: op1_09_in07 = imem05_in[75:72];
    10: op1_09_in07 = reg_0451;
    11: op1_09_in07 = reg_0255;
    31: op1_09_in07 = reg_0255;
    12: op1_09_in07 = imem02_in[91:88];
    13: op1_09_in07 = imem03_in[39:36];
    14: op1_09_in07 = reg_0781;
    85: op1_09_in07 = reg_0781;
    15: op1_09_in07 = reg_0680;
    3: op1_09_in07 = reg_0434;
    16: op1_09_in07 = imem02_in[35:32];
    17: op1_09_in07 = reg_0676;
    18: op1_09_in07 = reg_0111;
    19: op1_09_in07 = reg_0686;
    20: op1_09_in07 = reg_0643;
    21: op1_09_in07 = reg_0702;
    22: op1_09_in07 = reg_0030;
    23: op1_09_in07 = reg_0034;
    24: op1_09_in07 = reg_0691;
    88: op1_09_in07 = reg_0691;
    25: op1_09_in07 = imem04_in[27:24];
    41: op1_09_in07 = imem04_in[27:24];
    26: op1_09_in07 = reg_0455;
    27: op1_09_in07 = reg_0658;
    28: op1_09_in07 = reg_0682;
    29: op1_09_in07 = reg_0679;
    30: op1_09_in07 = reg_0365;
    32: op1_09_in07 = reg_0611;
    33: op1_09_in07 = reg_0453;
    34: op1_09_in07 = reg_0258;
    35: op1_09_in07 = reg_0292;
    36: op1_09_in07 = reg_0152;
    37: op1_09_in07 = imem04_in[39:36];
    38: op1_09_in07 = imem07_in[39:36];
    39: op1_09_in07 = reg_0672;
    40: op1_09_in07 = reg_0694;
    42: op1_09_in07 = reg_0793;
    43: op1_09_in07 = reg_0175;
    44: op1_09_in07 = imem02_in[63:60];
    45: op1_09_in07 = reg_0068;
    46: op1_09_in07 = imem07_in[19:16];
    47: op1_09_in07 = reg_0254;
    48: op1_09_in07 = reg_0800;
    49: op1_09_in07 = reg_0243;
    50: op1_09_in07 = reg_0693;
    51: op1_09_in07 = reg_0169;
    52: op1_09_in07 = reg_0685;
    53: op1_09_in07 = imem00_in[115:112];
    54: op1_09_in07 = reg_0527;
    55: op1_09_in07 = reg_0097;
    56: op1_09_in07 = reg_0589;
    57: op1_09_in07 = reg_0043;
    58: op1_09_in07 = reg_0305;
    59: op1_09_in07 = reg_0070;
    60: op1_09_in07 = reg_0133;
    61: op1_09_in07 = reg_0713;
    62: op1_09_in07 = reg_0645;
    63: op1_09_in07 = imem02_in[47:44];
    82: op1_09_in07 = imem02_in[47:44];
    64: op1_09_in07 = reg_0357;
    65: op1_09_in07 = reg_0262;
    66: op1_09_in07 = reg_0010;
    67: op1_09_in07 = reg_0520;
    68: op1_09_in07 = reg_0480;
    69: op1_09_in07 = reg_0052;
    70: op1_09_in07 = reg_0790;
    71: op1_09_in07 = reg_0107;
    72: op1_09_in07 = reg_0552;
    73: op1_09_in07 = imem04_in[3:0];
    74: op1_09_in07 = reg_0291;
    76: op1_09_in07 = reg_0744;
    77: op1_09_in07 = reg_0464;
    78: op1_09_in07 = reg_0678;
    79: op1_09_in07 = reg_0078;
    80: op1_09_in07 = reg_0149;
    81: op1_09_in07 = imem04_in[15:12];
    83: op1_09_in07 = imem07_in[23:20];
    84: op1_09_in07 = reg_0003;
    86: op1_09_in07 = reg_0758;
    87: op1_09_in07 = reg_0566;
    89: op1_09_in07 = reg_0009;
    90: op1_09_in07 = reg_0740;
    91: op1_09_in07 = reg_0516;
    92: op1_09_in07 = reg_0716;
    93: op1_09_in07 = reg_0215;
    94: op1_09_in07 = reg_0613;
    95: op1_09_in07 = reg_0695;
    96: op1_09_in07 = reg_0143;
    default: op1_09_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_09_inv07 = 1;
    5: op1_09_inv07 = 1;
    6: op1_09_inv07 = 1;
    7: op1_09_inv07 = 1;
    8: op1_09_inv07 = 1;
    10: op1_09_inv07 = 1;
    11: op1_09_inv07 = 1;
    12: op1_09_inv07 = 1;
    14: op1_09_inv07 = 1;
    18: op1_09_inv07 = 1;
    19: op1_09_inv07 = 1;
    23: op1_09_inv07 = 1;
    24: op1_09_inv07 = 1;
    25: op1_09_inv07 = 1;
    27: op1_09_inv07 = 1;
    31: op1_09_inv07 = 1;
    34: op1_09_inv07 = 1;
    36: op1_09_inv07 = 1;
    39: op1_09_inv07 = 1;
    43: op1_09_inv07 = 1;
    44: op1_09_inv07 = 1;
    45: op1_09_inv07 = 1;
    50: op1_09_inv07 = 1;
    58: op1_09_inv07 = 1;
    60: op1_09_inv07 = 1;
    61: op1_09_inv07 = 1;
    62: op1_09_inv07 = 1;
    63: op1_09_inv07 = 1;
    65: op1_09_inv07 = 1;
    66: op1_09_inv07 = 1;
    67: op1_09_inv07 = 1;
    71: op1_09_inv07 = 1;
    74: op1_09_inv07 = 1;
    77: op1_09_inv07 = 1;
    79: op1_09_inv07 = 1;
    80: op1_09_inv07 = 1;
    81: op1_09_inv07 = 1;
    84: op1_09_inv07 = 1;
    85: op1_09_inv07 = 1;
    86: op1_09_inv07 = 1;
    87: op1_09_inv07 = 1;
    88: op1_09_inv07 = 1;
    89: op1_09_inv07 = 1;
    90: op1_09_inv07 = 1;
    91: op1_09_inv07 = 1;
    92: op1_09_inv07 = 1;
    default: op1_09_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in08 = reg_0181;
    5: op1_09_in08 = imem06_in[3:0];
    96: op1_09_in08 = imem06_in[3:0];
    6: op1_09_in08 = reg_0469;
    10: op1_09_in08 = reg_0469;
    7: op1_09_in08 = reg_0009;
    8: op1_09_in08 = reg_0714;
    9: op1_09_in08 = imem05_in[99:96];
    11: op1_09_in08 = reg_0257;
    12: op1_09_in08 = imem02_in[95:92];
    13: op1_09_in08 = imem03_in[63:60];
    14: op1_09_in08 = reg_0490;
    15: op1_09_in08 = reg_0688;
    39: op1_09_in08 = reg_0688;
    3: op1_09_in08 = reg_0427;
    16: op1_09_in08 = imem02_in[59:56];
    17: op1_09_in08 = reg_0674;
    24: op1_09_in08 = reg_0674;
    18: op1_09_in08 = reg_0118;
    19: op1_09_in08 = reg_0690;
    20: op1_09_in08 = reg_0328;
    93: op1_09_in08 = reg_0328;
    21: op1_09_in08 = reg_0708;
    22: op1_09_in08 = reg_0038;
    23: op1_09_in08 = reg_0819;
    25: op1_09_in08 = reg_0544;
    65: op1_09_in08 = reg_0544;
    26: op1_09_in08 = reg_0457;
    27: op1_09_in08 = reg_0653;
    28: op1_09_in08 = reg_0681;
    29: op1_09_in08 = reg_0677;
    30: op1_09_in08 = reg_0322;
    31: op1_09_in08 = reg_0072;
    32: op1_09_in08 = reg_0618;
    33: op1_09_in08 = reg_0481;
    34: op1_09_in08 = reg_0062;
    35: op1_09_in08 = reg_0266;
    36: op1_09_in08 = reg_0143;
    85: op1_09_in08 = reg_0143;
    37: op1_09_in08 = imem04_in[79:76];
    38: op1_09_in08 = imem07_in[59:56];
    40: op1_09_in08 = reg_0689;
    41: op1_09_in08 = imem04_in[71:68];
    42: op1_09_in08 = reg_0787;
    43: op1_09_in08 = reg_0180;
    44: op1_09_in08 = reg_0357;
    45: op1_09_in08 = reg_0246;
    46: op1_09_in08 = imem07_in[35:32];
    47: op1_09_in08 = reg_0651;
    48: op1_09_in08 = reg_0805;
    49: op1_09_in08 = reg_0105;
    50: op1_09_in08 = reg_0676;
    51: op1_09_in08 = reg_0160;
    52: op1_09_in08 = reg_0698;
    53: op1_09_in08 = imem00_in[119:116];
    54: op1_09_in08 = reg_0530;
    55: op1_09_in08 = reg_0770;
    56: op1_09_in08 = reg_0750;
    57: op1_09_in08 = reg_0055;
    58: op1_09_in08 = reg_0433;
    59: op1_09_in08 = reg_0249;
    60: op1_09_in08 = reg_0134;
    61: op1_09_in08 = reg_0707;
    62: op1_09_in08 = reg_0227;
    63: op1_09_in08 = imem02_in[67:64];
    64: op1_09_in08 = reg_0394;
    66: op1_09_in08 = imem04_in[7:4];
    67: op1_09_in08 = reg_0777;
    68: op1_09_in08 = reg_0452;
    69: op1_09_in08 = reg_0076;
    70: op1_09_in08 = reg_0136;
    71: op1_09_in08 = reg_0126;
    72: op1_09_in08 = reg_0516;
    73: op1_09_in08 = imem04_in[39:36];
    74: op1_09_in08 = reg_0577;
    76: op1_09_in08 = reg_0407;
    77: op1_09_in08 = reg_0477;
    78: op1_09_in08 = imem02_in[19:16];
    79: op1_09_in08 = reg_0069;
    80: op1_09_in08 = reg_0785;
    81: op1_09_in08 = imem04_in[27:24];
    82: op1_09_in08 = imem02_in[55:52];
    83: op1_09_in08 = imem07_in[83:80];
    84: op1_09_in08 = reg_0015;
    86: op1_09_in08 = reg_0494;
    87: op1_09_in08 = reg_0540;
    88: op1_09_in08 = reg_0758;
    89: op1_09_in08 = reg_0648;
    90: op1_09_in08 = imem03_in[23:20];
    91: op1_09_in08 = reg_0052;
    92: op1_09_in08 = reg_0161;
    94: op1_09_in08 = reg_0659;
    95: op1_09_in08 = reg_0685;
    default: op1_09_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv08 = 1;
    11: op1_09_inv08 = 1;
    14: op1_09_inv08 = 1;
    15: op1_09_inv08 = 1;
    16: op1_09_inv08 = 1;
    18: op1_09_inv08 = 1;
    19: op1_09_inv08 = 1;
    21: op1_09_inv08 = 1;
    23: op1_09_inv08 = 1;
    28: op1_09_inv08 = 1;
    32: op1_09_inv08 = 1;
    35: op1_09_inv08 = 1;
    38: op1_09_inv08 = 1;
    39: op1_09_inv08 = 1;
    40: op1_09_inv08 = 1;
    44: op1_09_inv08 = 1;
    46: op1_09_inv08 = 1;
    50: op1_09_inv08 = 1;
    52: op1_09_inv08 = 1;
    53: op1_09_inv08 = 1;
    59: op1_09_inv08 = 1;
    62: op1_09_inv08 = 1;
    63: op1_09_inv08 = 1;
    66: op1_09_inv08 = 1;
    68: op1_09_inv08 = 1;
    69: op1_09_inv08 = 1;
    72: op1_09_inv08 = 1;
    73: op1_09_inv08 = 1;
    76: op1_09_inv08 = 1;
    79: op1_09_inv08 = 1;
    80: op1_09_inv08 = 1;
    81: op1_09_inv08 = 1;
    83: op1_09_inv08 = 1;
    89: op1_09_inv08 = 1;
    92: op1_09_inv08 = 1;
    94: op1_09_inv08 = 1;
    96: op1_09_inv08 = 1;
    default: op1_09_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in09 = reg_0182;
    5: op1_09_in09 = imem06_in[19:16];
    6: op1_09_in09 = reg_0471;
    7: op1_09_in09 = reg_0004;
    8: op1_09_in09 = reg_0712;
    9: op1_09_in09 = imem05_in[111:108];
    10: op1_09_in09 = reg_0474;
    11: op1_09_in09 = reg_0482;
    12: op1_09_in09 = imem02_in[107:104];
    13: op1_09_in09 = imem03_in[95:92];
    14: op1_09_in09 = reg_0788;
    15: op1_09_in09 = reg_0673;
    3: op1_09_in09 = reg_0435;
    16: op1_09_in09 = imem02_in[91:88];
    17: op1_09_in09 = reg_0671;
    18: op1_09_in09 = reg_0099;
    19: op1_09_in09 = reg_0691;
    29: op1_09_in09 = reg_0691;
    20: op1_09_in09 = imem02_in[7:4];
    21: op1_09_in09 = reg_0709;
    22: op1_09_in09 = reg_0749;
    23: op1_09_in09 = reg_0814;
    24: op1_09_in09 = reg_0675;
    25: op1_09_in09 = reg_0315;
    26: op1_09_in09 = reg_0452;
    27: op1_09_in09 = reg_0664;
    62: op1_09_in09 = reg_0664;
    28: op1_09_in09 = reg_0685;
    30: op1_09_in09 = reg_0323;
    31: op1_09_in09 = imem05_in[15:12];
    32: op1_09_in09 = reg_0622;
    33: op1_09_in09 = reg_0473;
    34: op1_09_in09 = reg_0067;
    35: op1_09_in09 = reg_0051;
    36: op1_09_in09 = reg_0138;
    37: op1_09_in09 = imem04_in[103:100];
    38: op1_09_in09 = imem07_in[67:64];
    39: op1_09_in09 = reg_0469;
    40: op1_09_in09 = reg_0668;
    41: op1_09_in09 = imem04_in[83:80];
    42: op1_09_in09 = reg_0741;
    43: op1_09_in09 = reg_0162;
    44: op1_09_in09 = reg_0362;
    45: op1_09_in09 = reg_0288;
    46: op1_09_in09 = imem07_in[47:44];
    47: op1_09_in09 = reg_0426;
    48: op1_09_in09 = reg_0809;
    49: op1_09_in09 = reg_0111;
    50: op1_09_in09 = reg_0677;
    51: op1_09_in09 = reg_0163;
    52: op1_09_in09 = reg_0686;
    53: op1_09_in09 = reg_0693;
    54: op1_09_in09 = reg_0097;
    55: op1_09_in09 = reg_0498;
    56: op1_09_in09 = reg_0116;
    57: op1_09_in09 = reg_0057;
    58: op1_09_in09 = reg_0529;
    59: op1_09_in09 = reg_0101;
    60: op1_09_in09 = reg_0075;
    61: op1_09_in09 = reg_0727;
    63: op1_09_in09 = imem02_in[123:120];
    64: op1_09_in09 = reg_0392;
    65: op1_09_in09 = reg_0328;
    66: op1_09_in09 = imem04_in[51:48];
    73: op1_09_in09 = imem04_in[51:48];
    67: op1_09_in09 = reg_0218;
    68: op1_09_in09 = reg_0189;
    77: op1_09_in09 = reg_0189;
    69: op1_09_in09 = reg_0430;
    70: op1_09_in09 = reg_0156;
    71: op1_09_in09 = reg_0678;
    72: op1_09_in09 = reg_0547;
    74: op1_09_in09 = reg_0762;
    76: op1_09_in09 = reg_0461;
    78: op1_09_in09 = imem02_in[55:52];
    79: op1_09_in09 = imem05_in[19:16];
    80: op1_09_in09 = reg_0152;
    81: op1_09_in09 = imem04_in[43:40];
    82: op1_09_in09 = imem02_in[63:60];
    83: op1_09_in09 = imem07_in[91:88];
    84: op1_09_in09 = reg_0806;
    85: op1_09_in09 = reg_0369;
    86: op1_09_in09 = reg_0634;
    87: op1_09_in09 = reg_0770;
    88: op1_09_in09 = reg_0453;
    89: op1_09_in09 = reg_0395;
    90: op1_09_in09 = imem03_in[67:64];
    91: op1_09_in09 = reg_0614;
    92: op1_09_in09 = reg_0167;
    93: op1_09_in09 = reg_0651;
    94: op1_09_in09 = reg_0242;
    95: op1_09_in09 = reg_0698;
    96: op1_09_in09 = imem06_in[7:4];
    default: op1_09_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv09 = 1;
    8: op1_09_inv09 = 1;
    9: op1_09_inv09 = 1;
    10: op1_09_inv09 = 1;
    12: op1_09_inv09 = 1;
    13: op1_09_inv09 = 1;
    14: op1_09_inv09 = 1;
    15: op1_09_inv09 = 1;
    3: op1_09_inv09 = 1;
    16: op1_09_inv09 = 1;
    17: op1_09_inv09 = 1;
    18: op1_09_inv09 = 1;
    20: op1_09_inv09 = 1;
    21: op1_09_inv09 = 1;
    22: op1_09_inv09 = 1;
    23: op1_09_inv09 = 1;
    28: op1_09_inv09 = 1;
    31: op1_09_inv09 = 1;
    34: op1_09_inv09 = 1;
    35: op1_09_inv09 = 1;
    41: op1_09_inv09 = 1;
    42: op1_09_inv09 = 1;
    44: op1_09_inv09 = 1;
    45: op1_09_inv09 = 1;
    46: op1_09_inv09 = 1;
    48: op1_09_inv09 = 1;
    50: op1_09_inv09 = 1;
    54: op1_09_inv09 = 1;
    55: op1_09_inv09 = 1;
    56: op1_09_inv09 = 1;
    59: op1_09_inv09 = 1;
    60: op1_09_inv09 = 1;
    63: op1_09_inv09 = 1;
    65: op1_09_inv09 = 1;
    66: op1_09_inv09 = 1;
    67: op1_09_inv09 = 1;
    69: op1_09_inv09 = 1;
    72: op1_09_inv09 = 1;
    78: op1_09_inv09 = 1;
    79: op1_09_inv09 = 1;
    80: op1_09_inv09 = 1;
    81: op1_09_inv09 = 1;
    82: op1_09_inv09 = 1;
    85: op1_09_inv09 = 1;
    86: op1_09_inv09 = 1;
    89: op1_09_inv09 = 1;
    92: op1_09_inv09 = 1;
    93: op1_09_inv09 = 1;
    94: op1_09_inv09 = 1;
    96: op1_09_inv09 = 1;
    default: op1_09_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_09_in10 = reg_0166;
    5: op1_09_in10 = imem06_in[67:64];
    6: op1_09_in10 = reg_0191;
    7: op1_09_in10 = imem04_in[11:8];
    8: op1_09_in10 = reg_0709;
    9: op1_09_in10 = reg_0271;
    42: op1_09_in10 = reg_0271;
    10: op1_09_in10 = reg_0193;
    68: op1_09_in10 = reg_0193;
    77: op1_09_in10 = reg_0193;
    11: op1_09_in10 = reg_0490;
    12: op1_09_in10 = imem02_in[127:124];
    13: op1_09_in10 = reg_0599;
    14: op1_09_in10 = reg_0793;
    15: op1_09_in10 = reg_0455;
    3: op1_09_in10 = reg_0183;
    16: op1_09_in10 = imem02_in[115:112];
    17: op1_09_in10 = reg_0465;
    40: op1_09_in10 = reg_0465;
    18: op1_09_in10 = reg_0114;
    19: op1_09_in10 = reg_0680;
    20: op1_09_in10 = imem02_in[31:28];
    21: op1_09_in10 = reg_0713;
    22: op1_09_in10 = imem07_in[7:4];
    23: op1_09_in10 = reg_0748;
    24: op1_09_in10 = reg_0463;
    25: op1_09_in10 = reg_0088;
    26: op1_09_in10 = reg_0458;
    27: op1_09_in10 = reg_0656;
    67: op1_09_in10 = reg_0656;
    28: op1_09_in10 = reg_0684;
    29: op1_09_in10 = reg_0453;
    30: op1_09_in10 = reg_0314;
    31: op1_09_in10 = imem05_in[35:32];
    32: op1_09_in10 = reg_0317;
    33: op1_09_in10 = reg_0214;
    34: op1_09_in10 = reg_0063;
    35: op1_09_in10 = reg_0281;
    36: op1_09_in10 = reg_0141;
    37: op1_09_in10 = imem04_in[115:112];
    38: op1_09_in10 = imem07_in[83:80];
    39: op1_09_in10 = reg_0460;
    41: op1_09_in10 = reg_0061;
    43: op1_09_in10 = reg_0170;
    44: op1_09_in10 = reg_0345;
    45: op1_09_in10 = reg_0249;
    46: op1_09_in10 = reg_0704;
    47: op1_09_in10 = reg_0344;
    48: op1_09_in10 = reg_0070;
    49: op1_09_in10 = reg_0104;
    50: op1_09_in10 = reg_0674;
    52: op1_09_in10 = reg_0688;
    53: op1_09_in10 = reg_0696;
    54: op1_09_in10 = reg_0348;
    55: op1_09_in10 = imem03_in[31:28];
    56: op1_09_in10 = reg_0588;
    57: op1_09_in10 = reg_0536;
    58: op1_09_in10 = reg_0071;
    69: op1_09_in10 = reg_0071;
    59: op1_09_in10 = reg_0285;
    60: op1_09_in10 = reg_0372;
    61: op1_09_in10 = reg_0436;
    62: op1_09_in10 = reg_0112;
    63: op1_09_in10 = reg_0501;
    64: op1_09_in10 = reg_0376;
    65: op1_09_in10 = reg_0552;
    66: op1_09_in10 = imem04_in[67:64];
    70: op1_09_in10 = reg_0138;
    71: op1_09_in10 = reg_0666;
    72: op1_09_in10 = reg_0433;
    73: op1_09_in10 = imem04_in[63:60];
    74: op1_09_in10 = reg_0370;
    76: op1_09_in10 = reg_0211;
    78: op1_09_in10 = imem02_in[63:60];
    79: op1_09_in10 = imem05_in[43:40];
    80: op1_09_in10 = reg_0796;
    81: op1_09_in10 = imem04_in[79:76];
    82: op1_09_in10 = imem02_in[107:104];
    83: op1_09_in10 = imem07_in[103:100];
    84: op1_09_in10 = imem04_in[23:20];
    85: op1_09_in10 = reg_0816;
    86: op1_09_in10 = reg_0461;
    87: op1_09_in10 = reg_0756;
    88: op1_09_in10 = reg_0207;
    89: op1_09_in10 = reg_0575;
    90: op1_09_in10 = imem03_in[87:84];
    91: op1_09_in10 = reg_0774;
    92: op1_09_in10 = reg_0164;
    93: op1_09_in10 = reg_0813;
    94: op1_09_in10 = reg_0576;
    95: op1_09_in10 = reg_0749;
    96: op1_09_in10 = imem06_in[31:28];
    default: op1_09_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_09_inv10 = 1;
    5: op1_09_inv10 = 1;
    7: op1_09_inv10 = 1;
    8: op1_09_inv10 = 1;
    9: op1_09_inv10 = 1;
    10: op1_09_inv10 = 1;
    11: op1_09_inv10 = 1;
    12: op1_09_inv10 = 1;
    14: op1_09_inv10 = 1;
    3: op1_09_inv10 = 1;
    16: op1_09_inv10 = 1;
    17: op1_09_inv10 = 1;
    19: op1_09_inv10 = 1;
    20: op1_09_inv10 = 1;
    22: op1_09_inv10 = 1;
    23: op1_09_inv10 = 1;
    25: op1_09_inv10 = 1;
    26: op1_09_inv10 = 1;
    27: op1_09_inv10 = 1;
    28: op1_09_inv10 = 1;
    29: op1_09_inv10 = 1;
    31: op1_09_inv10 = 1;
    32: op1_09_inv10 = 1;
    39: op1_09_inv10 = 1;
    43: op1_09_inv10 = 1;
    45: op1_09_inv10 = 1;
    46: op1_09_inv10 = 1;
    48: op1_09_inv10 = 1;
    49: op1_09_inv10 = 1;
    55: op1_09_inv10 = 1;
    57: op1_09_inv10 = 1;
    59: op1_09_inv10 = 1;
    60: op1_09_inv10 = 1;
    62: op1_09_inv10 = 1;
    64: op1_09_inv10 = 1;
    65: op1_09_inv10 = 1;
    67: op1_09_inv10 = 1;
    69: op1_09_inv10 = 1;
    73: op1_09_inv10 = 1;
    76: op1_09_inv10 = 1;
    77: op1_09_inv10 = 1;
    78: op1_09_inv10 = 1;
    79: op1_09_inv10 = 1;
    81: op1_09_inv10 = 1;
    86: op1_09_inv10 = 1;
    88: op1_09_inv10 = 1;
    89: op1_09_inv10 = 1;
    91: op1_09_inv10 = 1;
    93: op1_09_inv10 = 1;
    default: op1_09_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の11番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in11 = reg_0628;
    6: op1_09_in11 = reg_0212;
    10: op1_09_in11 = reg_0212;
    7: op1_09_in11 = imem04_in[15:12];
    8: op1_09_in11 = reg_0701;
    9: op1_09_in11 = reg_0259;
    11: op1_09_in11 = reg_0789;
    12: op1_09_in11 = reg_0648;
    13: op1_09_in11 = reg_0583;
    14: op1_09_in11 = reg_0785;
    15: op1_09_in11 = reg_0476;
    86: op1_09_in11 = reg_0476;
    3: op1_09_in11 = reg_0168;
    16: op1_09_in11 = reg_0647;
    17: op1_09_in11 = reg_0469;
    18: op1_09_in11 = reg_0113;
    19: op1_09_in11 = reg_0459;
    20: op1_09_in11 = imem03_in[7:4];
    21: op1_09_in11 = reg_0441;
    22: op1_09_in11 = imem07_in[23:20];
    23: op1_09_in11 = reg_0750;
    24: op1_09_in11 = reg_0457;
    25: op1_09_in11 = reg_0057;
    26: op1_09_in11 = reg_0188;
    27: op1_09_in11 = reg_0644;
    28: op1_09_in11 = reg_0690;
    29: op1_09_in11 = reg_0481;
    30: op1_09_in11 = reg_0082;
    31: op1_09_in11 = imem05_in[55:52];
    32: op1_09_in11 = reg_0408;
    33: op1_09_in11 = reg_0208;
    34: op1_09_in11 = reg_0064;
    35: op1_09_in11 = reg_0062;
    36: op1_09_in11 = reg_0130;
    37: op1_09_in11 = reg_0262;
    81: op1_09_in11 = reg_0262;
    38: op1_09_in11 = imem07_in[99:96];
    39: op1_09_in11 = reg_0473;
    40: op1_09_in11 = reg_0450;
    41: op1_09_in11 = reg_0066;
    42: op1_09_in11 = reg_0260;
    44: op1_09_in11 = reg_0363;
    45: op1_09_in11 = reg_0544;
    46: op1_09_in11 = reg_0719;
    47: op1_09_in11 = reg_0365;
    48: op1_09_in11 = reg_0229;
    49: op1_09_in11 = reg_0112;
    50: op1_09_in11 = reg_0678;
    52: op1_09_in11 = reg_0464;
    53: op1_09_in11 = reg_0698;
    54: op1_09_in11 = reg_0270;
    55: op1_09_in11 = imem03_in[43:40];
    56: op1_09_in11 = reg_0398;
    57: op1_09_in11 = reg_0280;
    58: op1_09_in11 = reg_0616;
    59: op1_09_in11 = reg_0089;
    60: op1_09_in11 = reg_0621;
    61: op1_09_in11 = reg_0051;
    62: op1_09_in11 = reg_0665;
    63: op1_09_in11 = reg_0045;
    64: op1_09_in11 = reg_0499;
    65: op1_09_in11 = reg_0542;
    66: op1_09_in11 = imem04_in[71:68];
    67: op1_09_in11 = reg_0507;
    68: op1_09_in11 = reg_0207;
    69: op1_09_in11 = reg_0297;
    72: op1_09_in11 = reg_0297;
    70: op1_09_in11 = reg_0607;
    71: op1_09_in11 = reg_0128;
    73: op1_09_in11 = imem04_in[75:72];
    74: op1_09_in11 = reg_0238;
    76: op1_09_in11 = imem01_in[67:64];
    77: op1_09_in11 = reg_0198;
    78: op1_09_in11 = imem02_in[107:104];
    79: op1_09_in11 = imem05_in[47:44];
    91: op1_09_in11 = imem05_in[47:44];
    80: op1_09_in11 = reg_0783;
    82: op1_09_in11 = imem02_in[123:120];
    83: op1_09_in11 = imem07_in[115:112];
    84: op1_09_in11 = imem04_in[43:40];
    85: op1_09_in11 = reg_0375;
    87: op1_09_in11 = reg_0094;
    88: op1_09_in11 = reg_0206;
    89: op1_09_in11 = reg_0755;
    90: op1_09_in11 = reg_0604;
    92: op1_09_in11 = reg_0708;
    93: op1_09_in11 = reg_0620;
    94: op1_09_in11 = reg_0681;
    95: op1_09_in11 = reg_0691;
    96: op1_09_in11 = imem06_in[47:44];
    default: op1_09_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv11 = 1;
    9: op1_09_inv11 = 1;
    10: op1_09_inv11 = 1;
    14: op1_09_inv11 = 1;
    18: op1_09_inv11 = 1;
    19: op1_09_inv11 = 1;
    20: op1_09_inv11 = 1;
    22: op1_09_inv11 = 1;
    23: op1_09_inv11 = 1;
    24: op1_09_inv11 = 1;
    25: op1_09_inv11 = 1;
    27: op1_09_inv11 = 1;
    28: op1_09_inv11 = 1;
    29: op1_09_inv11 = 1;
    36: op1_09_inv11 = 1;
    41: op1_09_inv11 = 1;
    42: op1_09_inv11 = 1;
    44: op1_09_inv11 = 1;
    46: op1_09_inv11 = 1;
    47: op1_09_inv11 = 1;
    48: op1_09_inv11 = 1;
    50: op1_09_inv11 = 1;
    52: op1_09_inv11 = 1;
    54: op1_09_inv11 = 1;
    55: op1_09_inv11 = 1;
    60: op1_09_inv11 = 1;
    61: op1_09_inv11 = 1;
    62: op1_09_inv11 = 1;
    63: op1_09_inv11 = 1;
    68: op1_09_inv11 = 1;
    71: op1_09_inv11 = 1;
    73: op1_09_inv11 = 1;
    74: op1_09_inv11 = 1;
    76: op1_09_inv11 = 1;
    79: op1_09_inv11 = 1;
    80: op1_09_inv11 = 1;
    81: op1_09_inv11 = 1;
    89: op1_09_inv11 = 1;
    93: op1_09_inv11 = 1;
    94: op1_09_inv11 = 1;
    default: op1_09_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の12番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in12 = reg_0610;
    6: op1_09_in12 = imem01_in[23:20];
    7: op1_09_in12 = imem04_in[23:20];
    8: op1_09_in12 = reg_0700;
    9: op1_09_in12 = reg_0252;
    10: op1_09_in12 = reg_0190;
    11: op1_09_in12 = reg_0494;
    12: op1_09_in12 = reg_0652;
    13: op1_09_in12 = reg_0591;
    14: op1_09_in12 = reg_0794;
    15: op1_09_in12 = reg_0479;
    16: op1_09_in12 = reg_0640;
    17: op1_09_in12 = reg_0476;
    18: op1_09_in12 = imem02_in[51:48];
    19: op1_09_in12 = reg_0191;
    20: op1_09_in12 = imem03_in[23:20];
    21: op1_09_in12 = reg_0430;
    22: op1_09_in12 = imem07_in[103:100];
    38: op1_09_in12 = imem07_in[103:100];
    23: op1_09_in12 = reg_0029;
    24: op1_09_in12 = reg_0475;
    25: op1_09_in12 = reg_0551;
    26: op1_09_in12 = reg_0203;
    27: op1_09_in12 = reg_0636;
    28: op1_09_in12 = reg_0668;
    29: op1_09_in12 = reg_0472;
    30: op1_09_in12 = reg_0756;
    31: op1_09_in12 = imem05_in[71:68];
    32: op1_09_in12 = reg_0329;
    33: op1_09_in12 = reg_0207;
    34: op1_09_in12 = reg_0256;
    35: op1_09_in12 = reg_0289;
    36: op1_09_in12 = reg_0144;
    37: op1_09_in12 = reg_0087;
    39: op1_09_in12 = reg_0470;
    40: op1_09_in12 = reg_0469;
    41: op1_09_in12 = reg_0068;
    42: op1_09_in12 = reg_0307;
    44: op1_09_in12 = reg_0347;
    45: op1_09_in12 = reg_0315;
    46: op1_09_in12 = reg_0710;
    83: op1_09_in12 = reg_0710;
    47: op1_09_in12 = reg_0342;
    48: op1_09_in12 = reg_0544;
    49: op1_09_in12 = reg_0106;
    50: op1_09_in12 = reg_0675;
    52: op1_09_in12 = reg_0478;
    53: op1_09_in12 = reg_0689;
    54: op1_09_in12 = reg_0401;
    55: op1_09_in12 = imem03_in[95:92];
    56: op1_09_in12 = reg_0386;
    64: op1_09_in12 = reg_0386;
    57: op1_09_in12 = reg_0077;
    58: op1_09_in12 = imem04_in[31:28];
    59: op1_09_in12 = reg_0147;
    60: op1_09_in12 = reg_0110;
    61: op1_09_in12 = reg_0442;
    62: op1_09_in12 = imem02_in[31:28];
    63: op1_09_in12 = reg_0666;
    65: op1_09_in12 = reg_0056;
    66: op1_09_in12 = imem04_in[87:84];
    67: op1_09_in12 = reg_0642;
    68: op1_09_in12 = reg_0194;
    69: op1_09_in12 = reg_0508;
    70: op1_09_in12 = reg_0034;
    71: op1_09_in12 = imem02_in[23:20];
    72: op1_09_in12 = reg_0780;
    73: op1_09_in12 = imem04_in[79:76];
    74: op1_09_in12 = reg_0293;
    76: op1_09_in12 = imem01_in[83:80];
    77: op1_09_in12 = reg_0199;
    78: op1_09_in12 = imem02_in[115:112];
    79: op1_09_in12 = imem05_in[55:52];
    80: op1_09_in12 = reg_0155;
    81: op1_09_in12 = reg_0537;
    82: op1_09_in12 = reg_0739;
    84: op1_09_in12 = imem04_in[103:100];
    85: op1_09_in12 = reg_0580;
    86: op1_09_in12 = reg_0471;
    87: op1_09_in12 = reg_0093;
    88: op1_09_in12 = reg_0197;
    89: op1_09_in12 = reg_0564;
    90: op1_09_in12 = reg_0338;
    91: op1_09_in12 = imem05_in[59:56];
    92: op1_09_in12 = reg_0789;
    93: op1_09_in12 = reg_0351;
    94: op1_09_in12 = reg_0650;
    95: op1_09_in12 = reg_0063;
    96: op1_09_in12 = reg_0577;
    default: op1_09_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv12 = 1;
    8: op1_09_inv12 = 1;
    11: op1_09_inv12 = 1;
    15: op1_09_inv12 = 1;
    16: op1_09_inv12 = 1;
    17: op1_09_inv12 = 1;
    18: op1_09_inv12 = 1;
    21: op1_09_inv12 = 1;
    23: op1_09_inv12 = 1;
    24: op1_09_inv12 = 1;
    26: op1_09_inv12 = 1;
    30: op1_09_inv12 = 1;
    33: op1_09_inv12 = 1;
    40: op1_09_inv12 = 1;
    41: op1_09_inv12 = 1;
    42: op1_09_inv12 = 1;
    44: op1_09_inv12 = 1;
    47: op1_09_inv12 = 1;
    50: op1_09_inv12 = 1;
    52: op1_09_inv12 = 1;
    55: op1_09_inv12 = 1;
    58: op1_09_inv12 = 1;
    59: op1_09_inv12 = 1;
    60: op1_09_inv12 = 1;
    61: op1_09_inv12 = 1;
    63: op1_09_inv12 = 1;
    64: op1_09_inv12 = 1;
    66: op1_09_inv12 = 1;
    68: op1_09_inv12 = 1;
    71: op1_09_inv12 = 1;
    74: op1_09_inv12 = 1;
    77: op1_09_inv12 = 1;
    78: op1_09_inv12 = 1;
    80: op1_09_inv12 = 1;
    81: op1_09_inv12 = 1;
    83: op1_09_inv12 = 1;
    86: op1_09_inv12 = 1;
    87: op1_09_inv12 = 1;
    89: op1_09_inv12 = 1;
    90: op1_09_inv12 = 1;
    default: op1_09_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の13番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in13 = reg_0629;
    6: op1_09_in13 = imem01_in[27:24];
    7: op1_09_in13 = imem04_in[55:52];
    8: op1_09_in13 = reg_0421;
    9: op1_09_in13 = reg_0258;
    10: op1_09_in13 = reg_0202;
    11: op1_09_in13 = reg_0783;
    12: op1_09_in13 = reg_0352;
    13: op1_09_in13 = reg_0563;
    14: op1_09_in13 = reg_0784;
    83: op1_09_in13 = reg_0784;
    15: op1_09_in13 = reg_0214;
    16: op1_09_in13 = reg_0648;
    17: op1_09_in13 = reg_0481;
    18: op1_09_in13 = imem02_in[63:60];
    19: op1_09_in13 = reg_0209;
    20: op1_09_in13 = reg_0584;
    82: op1_09_in13 = reg_0584;
    21: op1_09_in13 = reg_0447;
    22: op1_09_in13 = reg_0704;
    23: op1_09_in13 = imem07_in[23:20];
    24: op1_09_in13 = reg_0480;
    50: op1_09_in13 = reg_0480;
    25: op1_09_in13 = reg_0303;
    26: op1_09_in13 = imem01_in[3:0];
    77: op1_09_in13 = imem01_in[3:0];
    27: op1_09_in13 = reg_0344;
    28: op1_09_in13 = reg_0675;
    29: op1_09_in13 = reg_0470;
    30: op1_09_in13 = reg_0531;
    31: op1_09_in13 = reg_0791;
    32: op1_09_in13 = reg_0038;
    33: op1_09_in13 = reg_0213;
    34: op1_09_in13 = imem05_in[3:0];
    35: op1_09_in13 = reg_0254;
    36: op1_09_in13 = reg_0286;
    37: op1_09_in13 = reg_0542;
    38: op1_09_in13 = reg_0716;
    39: op1_09_in13 = reg_0193;
    40: op1_09_in13 = reg_0476;
    41: op1_09_in13 = reg_0063;
    42: op1_09_in13 = reg_0734;
    44: op1_09_in13 = reg_0080;
    45: op1_09_in13 = reg_0088;
    46: op1_09_in13 = reg_0723;
    47: op1_09_in13 = reg_0347;
    48: op1_09_in13 = reg_0055;
    65: op1_09_in13 = reg_0055;
    81: op1_09_in13 = reg_0055;
    49: op1_09_in13 = reg_0115;
    52: op1_09_in13 = reg_0208;
    53: op1_09_in13 = reg_0690;
    54: op1_09_in13 = imem03_in[15:12];
    55: op1_09_in13 = imem03_in[115:112];
    56: op1_09_in13 = reg_0002;
    57: op1_09_in13 = reg_0585;
    58: op1_09_in13 = imem04_in[47:44];
    59: op1_09_in13 = reg_0128;
    60: op1_09_in13 = reg_0037;
    61: op1_09_in13 = reg_0443;
    62: op1_09_in13 = imem02_in[55:52];
    63: op1_09_in13 = reg_0739;
    64: op1_09_in13 = reg_0374;
    66: op1_09_in13 = imem04_in[95:92];
    67: op1_09_in13 = reg_0368;
    68: op1_09_in13 = reg_0196;
    69: op1_09_in13 = reg_0626;
    70: op1_09_in13 = reg_0642;
    71: op1_09_in13 = imem02_in[51:48];
    72: op1_09_in13 = reg_0100;
    73: op1_09_in13 = imem04_in[119:116];
    74: op1_09_in13 = reg_0519;
    76: op1_09_in13 = imem01_in[87:84];
    78: op1_09_in13 = imem02_in[123:120];
    79: op1_09_in13 = imem05_in[71:68];
    80: op1_09_in13 = reg_0137;
    84: op1_09_in13 = reg_0262;
    85: op1_09_in13 = reg_0764;
    86: op1_09_in13 = reg_0468;
    87: op1_09_in13 = reg_0740;
    88: op1_09_in13 = imem01_in[19:16];
    89: op1_09_in13 = reg_0549;
    90: op1_09_in13 = reg_0599;
    91: op1_09_in13 = imem05_in[95:92];
    92: op1_09_in13 = reg_0334;
    93: op1_09_in13 = reg_0633;
    94: op1_09_in13 = imem07_in[15:12];
    95: op1_09_in13 = reg_0688;
    96: op1_09_in13 = reg_0605;
    default: op1_09_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv13 = 1;
    7: op1_09_inv13 = 1;
    10: op1_09_inv13 = 1;
    11: op1_09_inv13 = 1;
    13: op1_09_inv13 = 1;
    14: op1_09_inv13 = 1;
    17: op1_09_inv13 = 1;
    18: op1_09_inv13 = 1;
    20: op1_09_inv13 = 1;
    21: op1_09_inv13 = 1;
    22: op1_09_inv13 = 1;
    23: op1_09_inv13 = 1;
    29: op1_09_inv13 = 1;
    31: op1_09_inv13 = 1;
    33: op1_09_inv13 = 1;
    35: op1_09_inv13 = 1;
    38: op1_09_inv13 = 1;
    40: op1_09_inv13 = 1;
    41: op1_09_inv13 = 1;
    42: op1_09_inv13 = 1;
    44: op1_09_inv13 = 1;
    45: op1_09_inv13 = 1;
    46: op1_09_inv13 = 1;
    47: op1_09_inv13 = 1;
    52: op1_09_inv13 = 1;
    53: op1_09_inv13 = 1;
    54: op1_09_inv13 = 1;
    56: op1_09_inv13 = 1;
    57: op1_09_inv13 = 1;
    59: op1_09_inv13 = 1;
    60: op1_09_inv13 = 1;
    61: op1_09_inv13 = 1;
    66: op1_09_inv13 = 1;
    67: op1_09_inv13 = 1;
    68: op1_09_inv13 = 1;
    69: op1_09_inv13 = 1;
    70: op1_09_inv13 = 1;
    71: op1_09_inv13 = 1;
    72: op1_09_inv13 = 1;
    74: op1_09_inv13 = 1;
    76: op1_09_inv13 = 1;
    79: op1_09_inv13 = 1;
    81: op1_09_inv13 = 1;
    83: op1_09_inv13 = 1;
    86: op1_09_inv13 = 1;
    90: op1_09_inv13 = 1;
    93: op1_09_inv13 = 1;
    96: op1_09_inv13 = 1;
    default: op1_09_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の14番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in14 = reg_0630;
    6: op1_09_in14 = imem01_in[87:84];
    7: op1_09_in14 = imem04_in[95:92];
    8: op1_09_in14 = reg_0447;
    92: op1_09_in14 = reg_0447;
    9: op1_09_in14 = reg_0265;
    10: op1_09_in14 = reg_0738;
    11: op1_09_in14 = reg_0787;
    67: op1_09_in14 = reg_0787;
    12: op1_09_in14 = reg_0333;
    16: op1_09_in14 = reg_0333;
    13: op1_09_in14 = reg_0594;
    14: op1_09_in14 = reg_0486;
    15: op1_09_in14 = reg_0200;
    17: op1_09_in14 = reg_0470;
    18: op1_09_in14 = imem02_in[99:96];
    19: op1_09_in14 = reg_0207;
    20: op1_09_in14 = reg_0585;
    21: op1_09_in14 = reg_0418;
    22: op1_09_in14 = reg_0720;
    23: op1_09_in14 = imem07_in[55:52];
    24: op1_09_in14 = reg_0473;
    50: op1_09_in14 = reg_0473;
    25: op1_09_in14 = reg_0054;
    26: op1_09_in14 = imem01_in[67:64];
    27: op1_09_in14 = reg_0357;
    28: op1_09_in14 = reg_0673;
    29: op1_09_in14 = reg_0198;
    39: op1_09_in14 = reg_0198;
    30: op1_09_in14 = reg_0526;
    31: op1_09_in14 = reg_0798;
    32: op1_09_in14 = reg_0576;
    33: op1_09_in14 = reg_0195;
    34: op1_09_in14 = imem05_in[7:4];
    35: op1_09_in14 = reg_0256;
    36: op1_09_in14 = reg_0610;
    37: op1_09_in14 = reg_0536;
    38: op1_09_in14 = reg_0726;
    46: op1_09_in14 = reg_0726;
    40: op1_09_in14 = reg_0456;
    41: op1_09_in14 = imem05_in[11:8];
    42: op1_09_in14 = reg_0086;
    44: op1_09_in14 = imem03_in[7:4];
    45: op1_09_in14 = reg_0083;
    47: op1_09_in14 = reg_0314;
    48: op1_09_in14 = reg_0057;
    49: op1_09_in14 = reg_0127;
    52: op1_09_in14 = reg_0204;
    53: op1_09_in14 = reg_0688;
    54: op1_09_in14 = imem03_in[87:84];
    55: op1_09_in14 = imem03_in[119:116];
    56: op1_09_in14 = reg_0806;
    57: op1_09_in14 = reg_0065;
    58: op1_09_in14 = imem04_in[63:60];
    59: op1_09_in14 = reg_0142;
    60: op1_09_in14 = reg_0818;
    61: op1_09_in14 = reg_0448;
    62: op1_09_in14 = imem02_in[71:68];
    63: op1_09_in14 = reg_0039;
    64: op1_09_in14 = reg_0003;
    65: op1_09_in14 = reg_0516;
    66: op1_09_in14 = imem04_in[99:96];
    68: op1_09_in14 = reg_0663;
    69: op1_09_in14 = reg_0643;
    70: op1_09_in14 = reg_0132;
    71: op1_09_in14 = imem02_in[63:60];
    72: op1_09_in14 = imem05_in[67:64];
    73: op1_09_in14 = reg_0552;
    74: op1_09_in14 = reg_0816;
    76: op1_09_in14 = reg_0741;
    77: op1_09_in14 = imem01_in[11:8];
    78: op1_09_in14 = reg_0325;
    79: op1_09_in14 = imem05_in[83:80];
    80: op1_09_in14 = imem06_in[7:4];
    81: op1_09_in14 = reg_0551;
    82: op1_09_in14 = reg_0639;
    83: op1_09_in14 = reg_0725;
    84: op1_09_in14 = reg_0545;
    85: op1_09_in14 = reg_0348;
    86: op1_09_in14 = reg_0479;
    87: op1_09_in14 = reg_0377;
    88: op1_09_in14 = imem01_in[47:44];
    89: op1_09_in14 = reg_0398;
    90: op1_09_in14 = reg_0801;
    91: op1_09_in14 = reg_0146;
    93: op1_09_in14 = reg_0632;
    94: op1_09_in14 = imem07_in[23:20];
    95: op1_09_in14 = reg_0469;
    96: op1_09_in14 = reg_0370;
    default: op1_09_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_09_inv14 = 1;
    16: op1_09_inv14 = 1;
    18: op1_09_inv14 = 1;
    20: op1_09_inv14 = 1;
    23: op1_09_inv14 = 1;
    31: op1_09_inv14 = 1;
    32: op1_09_inv14 = 1;
    34: op1_09_inv14 = 1;
    37: op1_09_inv14 = 1;
    38: op1_09_inv14 = 1;
    39: op1_09_inv14 = 1;
    40: op1_09_inv14 = 1;
    42: op1_09_inv14 = 1;
    46: op1_09_inv14 = 1;
    49: op1_09_inv14 = 1;
    53: op1_09_inv14 = 1;
    54: op1_09_inv14 = 1;
    56: op1_09_inv14 = 1;
    59: op1_09_inv14 = 1;
    61: op1_09_inv14 = 1;
    66: op1_09_inv14 = 1;
    84: op1_09_inv14 = 1;
    85: op1_09_inv14 = 1;
    86: op1_09_inv14 = 1;
    88: op1_09_inv14 = 1;
    89: op1_09_inv14 = 1;
    95: op1_09_inv14 = 1;
    96: op1_09_inv14 = 1;
    default: op1_09_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の15番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in15 = reg_0631;
    6: op1_09_in15 = imem01_in[111:108];
    7: op1_09_in15 = imem04_in[119:116];
    8: op1_09_in15 = reg_0419;
    9: op1_09_in15 = reg_0272;
    10: op1_09_in15 = reg_0226;
    11: op1_09_in15 = imem05_in[63:60];
    35: op1_09_in15 = imem05_in[63:60];
    12: op1_09_in15 = reg_0320;
    13: op1_09_in15 = reg_0395;
    14: op1_09_in15 = reg_0736;
    15: op1_09_in15 = reg_0186;
    19: op1_09_in15 = reg_0186;
    16: op1_09_in15 = reg_0329;
    17: op1_09_in15 = reg_0456;
    18: op1_09_in15 = imem02_in[103:100];
    20: op1_09_in15 = reg_0578;
    21: op1_09_in15 = reg_0434;
    22: op1_09_in15 = reg_0721;
    23: op1_09_in15 = imem07_in[71:68];
    24: op1_09_in15 = reg_0452;
    86: op1_09_in15 = reg_0452;
    25: op1_09_in15 = reg_0301;
    26: op1_09_in15 = imem01_in[123:120];
    27: op1_09_in15 = reg_0364;
    28: op1_09_in15 = reg_0692;
    53: op1_09_in15 = reg_0692;
    29: op1_09_in15 = reg_0212;
    30: op1_09_in15 = reg_0538;
    31: op1_09_in15 = reg_0483;
    32: op1_09_in15 = reg_0040;
    33: op1_09_in15 = reg_0199;
    34: op1_09_in15 = imem05_in[23:20];
    36: op1_09_in15 = reg_0604;
    37: op1_09_in15 = reg_0058;
    38: op1_09_in15 = reg_0717;
    39: op1_09_in15 = reg_0197;
    40: op1_09_in15 = reg_0188;
    41: op1_09_in15 = imem05_in[55:52];
    42: op1_09_in15 = reg_0128;
    44: op1_09_in15 = imem03_in[15:12];
    45: op1_09_in15 = reg_0079;
    81: op1_09_in15 = reg_0079;
    46: op1_09_in15 = reg_0441;
    47: op1_09_in15 = reg_0095;
    48: op1_09_in15 = reg_0551;
    49: op1_09_in15 = reg_0110;
    50: op1_09_in15 = reg_0470;
    52: op1_09_in15 = reg_0194;
    54: op1_09_in15 = imem03_in[111:108];
    55: op1_09_in15 = reg_0317;
    56: op1_09_in15 = imem04_in[11:8];
    57: op1_09_in15 = reg_0640;
    58: op1_09_in15 = imem04_in[75:72];
    59: op1_09_in15 = reg_0146;
    60: op1_09_in15 = reg_0112;
    61: op1_09_in15 = reg_0161;
    62: op1_09_in15 = imem02_in[87:84];
    63: op1_09_in15 = reg_0548;
    64: op1_09_in15 = reg_0801;
    65: op1_09_in15 = reg_0556;
    66: op1_09_in15 = imem04_in[103:100];
    67: op1_09_in15 = reg_0029;
    68: op1_09_in15 = reg_0100;
    69: op1_09_in15 = reg_0311;
    70: op1_09_in15 = reg_0577;
    71: op1_09_in15 = imem02_in[71:68];
    72: op1_09_in15 = imem05_in[103:100];
    73: op1_09_in15 = reg_0537;
    74: op1_09_in15 = reg_0700;
    76: op1_09_in15 = reg_0131;
    77: op1_09_in15 = imem01_in[79:76];
    78: op1_09_in15 = reg_0392;
    79: op1_09_in15 = imem05_in[95:92];
    80: op1_09_in15 = imem06_in[15:12];
    82: op1_09_in15 = reg_0704;
    83: op1_09_in15 = reg_0446;
    84: op1_09_in15 = reg_0535;
    85: op1_09_in15 = reg_0762;
    87: op1_09_in15 = reg_0375;
    88: op1_09_in15 = reg_0085;
    89: op1_09_in15 = reg_0747;
    90: op1_09_in15 = reg_0403;
    91: op1_09_in15 = reg_0355;
    92: op1_09_in15 = reg_0061;
    93: op1_09_in15 = reg_0650;
    94: op1_09_in15 = imem07_in[31:28];
    95: op1_09_in15 = reg_0472;
    96: op1_09_in15 = reg_0814;
    default: op1_09_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv15 = 1;
    8: op1_09_inv15 = 1;
    12: op1_09_inv15 = 1;
    13: op1_09_inv15 = 1;
    14: op1_09_inv15 = 1;
    17: op1_09_inv15 = 1;
    19: op1_09_inv15 = 1;
    20: op1_09_inv15 = 1;
    22: op1_09_inv15 = 1;
    24: op1_09_inv15 = 1;
    25: op1_09_inv15 = 1;
    28: op1_09_inv15 = 1;
    32: op1_09_inv15 = 1;
    34: op1_09_inv15 = 1;
    35: op1_09_inv15 = 1;
    38: op1_09_inv15 = 1;
    40: op1_09_inv15 = 1;
    41: op1_09_inv15 = 1;
    42: op1_09_inv15 = 1;
    46: op1_09_inv15 = 1;
    47: op1_09_inv15 = 1;
    48: op1_09_inv15 = 1;
    49: op1_09_inv15 = 1;
    56: op1_09_inv15 = 1;
    58: op1_09_inv15 = 1;
    59: op1_09_inv15 = 1;
    60: op1_09_inv15 = 1;
    62: op1_09_inv15 = 1;
    63: op1_09_inv15 = 1;
    64: op1_09_inv15 = 1;
    69: op1_09_inv15 = 1;
    71: op1_09_inv15 = 1;
    72: op1_09_inv15 = 1;
    73: op1_09_inv15 = 1;
    74: op1_09_inv15 = 1;
    76: op1_09_inv15 = 1;
    77: op1_09_inv15 = 1;
    78: op1_09_inv15 = 1;
    79: op1_09_inv15 = 1;
    80: op1_09_inv15 = 1;
    84: op1_09_inv15 = 1;
    86: op1_09_inv15 = 1;
    87: op1_09_inv15 = 1;
    88: op1_09_inv15 = 1;
    89: op1_09_inv15 = 1;
    94: op1_09_inv15 = 1;
    96: op1_09_inv15 = 1;
    default: op1_09_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の16番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in16 = reg_0626;
    6: op1_09_in16 = imem01_in[127:124];
    7: op1_09_in16 = reg_0548;
    8: op1_09_in16 = reg_0434;
    9: op1_09_in16 = reg_0254;
    10: op1_09_in16 = reg_0736;
    11: op1_09_in16 = imem05_in[71:68];
    12: op1_09_in16 = reg_0359;
    13: op1_09_in16 = reg_0360;
    14: op1_09_in16 = reg_0259;
    15: op1_09_in16 = reg_0194;
    19: op1_09_in16 = reg_0194;
    16: op1_09_in16 = reg_0346;
    17: op1_09_in16 = reg_0196;
    52: op1_09_in16 = reg_0196;
    18: op1_09_in16 = imem02_in[115:112];
    20: op1_09_in16 = reg_0597;
    21: op1_09_in16 = reg_0443;
    22: op1_09_in16 = reg_0725;
    23: op1_09_in16 = imem07_in[79:76];
    24: op1_09_in16 = reg_0188;
    25: op1_09_in16 = reg_0284;
    26: op1_09_in16 = reg_0822;
    27: op1_09_in16 = reg_0342;
    28: op1_09_in16 = reg_0463;
    29: op1_09_in16 = imem01_in[47:44];
    30: op1_09_in16 = reg_0028;
    31: op1_09_in16 = reg_0488;
    32: op1_09_in16 = reg_0779;
    33: op1_09_in16 = imem01_in[51:48];
    34: op1_09_in16 = imem05_in[31:28];
    35: op1_09_in16 = imem05_in[87:84];
    36: op1_09_in16 = reg_0622;
    37: op1_09_in16 = reg_0295;
    38: op1_09_in16 = reg_0703;
    39: op1_09_in16 = reg_0217;
    40: op1_09_in16 = reg_0190;
    41: op1_09_in16 = imem05_in[63:60];
    42: op1_09_in16 = reg_0139;
    83: op1_09_in16 = reg_0139;
    44: op1_09_in16 = imem03_in[27:24];
    45: op1_09_in16 = reg_0283;
    46: op1_09_in16 = reg_0061;
    47: op1_09_in16 = reg_0498;
    48: op1_09_in16 = reg_0615;
    49: op1_09_in16 = imem02_in[3:0];
    50: op1_09_in16 = reg_0456;
    53: op1_09_in16 = reg_0454;
    54: op1_09_in16 = imem03_in[119:116];
    55: op1_09_in16 = reg_0596;
    56: op1_09_in16 = imem04_in[23:20];
    57: op1_09_in16 = imem05_in[3:0];
    58: op1_09_in16 = imem05_in[59:56];
    59: op1_09_in16 = reg_0153;
    60: op1_09_in16 = reg_0289;
    61: op1_09_in16 = reg_0185;
    62: op1_09_in16 = imem02_in[91:88];
    63: op1_09_in16 = reg_0320;
    64: op1_09_in16 = reg_0010;
    65: op1_09_in16 = reg_0303;
    66: op1_09_in16 = reg_0059;
    67: op1_09_in16 = imem07_in[23:20];
    68: op1_09_in16 = reg_0271;
    69: op1_09_in16 = reg_0371;
    70: op1_09_in16 = reg_0814;
    71: op1_09_in16 = imem02_in[79:76];
    72: op1_09_in16 = imem05_in[123:120];
    73: op1_09_in16 = reg_0631;
    74: op1_09_in16 = reg_0819;
    76: op1_09_in16 = reg_0394;
    77: op1_09_in16 = imem01_in[99:96];
    78: op1_09_in16 = reg_0487;
    79: op1_09_in16 = imem05_in[115:112];
    80: op1_09_in16 = imem06_in[71:68];
    81: op1_09_in16 = reg_0305;
    82: op1_09_in16 = reg_0753;
    84: op1_09_in16 = reg_0510;
    85: op1_09_in16 = reg_0409;
    86: op1_09_in16 = reg_0204;
    87: op1_09_in16 = reg_0588;
    88: op1_09_in16 = reg_0520;
    89: op1_09_in16 = reg_0396;
    90: op1_09_in16 = reg_0549;
    91: op1_09_in16 = reg_0552;
    92: op1_09_in16 = reg_0239;
    93: op1_09_in16 = imem07_in[43:40];
    94: op1_09_in16 = imem07_in[83:80];
    95: op1_09_in16 = reg_0480;
    96: op1_09_in16 = reg_0750;
    default: op1_09_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_09_inv16 = 1;
    9: op1_09_inv16 = 1;
    10: op1_09_inv16 = 1;
    11: op1_09_inv16 = 1;
    12: op1_09_inv16 = 1;
    15: op1_09_inv16 = 1;
    20: op1_09_inv16 = 1;
    22: op1_09_inv16 = 1;
    24: op1_09_inv16 = 1;
    25: op1_09_inv16 = 1;
    28: op1_09_inv16 = 1;
    30: op1_09_inv16 = 1;
    32: op1_09_inv16 = 1;
    34: op1_09_inv16 = 1;
    35: op1_09_inv16 = 1;
    36: op1_09_inv16 = 1;
    38: op1_09_inv16 = 1;
    39: op1_09_inv16 = 1;
    40: op1_09_inv16 = 1;
    52: op1_09_inv16 = 1;
    53: op1_09_inv16 = 1;
    54: op1_09_inv16 = 1;
    57: op1_09_inv16 = 1;
    59: op1_09_inv16 = 1;
    60: op1_09_inv16 = 1;
    61: op1_09_inv16 = 1;
    63: op1_09_inv16 = 1;
    67: op1_09_inv16 = 1;
    69: op1_09_inv16 = 1;
    70: op1_09_inv16 = 1;
    72: op1_09_inv16 = 1;
    73: op1_09_inv16 = 1;
    74: op1_09_inv16 = 1;
    78: op1_09_inv16 = 1;
    79: op1_09_inv16 = 1;
    80: op1_09_inv16 = 1;
    82: op1_09_inv16 = 1;
    83: op1_09_inv16 = 1;
    85: op1_09_inv16 = 1;
    90: op1_09_inv16 = 1;
    91: op1_09_inv16 = 1;
    95: op1_09_inv16 = 1;
    default: op1_09_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の17番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in17 = reg_0379;
    6: op1_09_in17 = reg_0509;
    7: op1_09_in17 = reg_0537;
    8: op1_09_in17 = reg_0444;
    9: op1_09_in17 = reg_0255;
    10: op1_09_in17 = reg_0224;
    11: op1_09_in17 = imem05_in[79:76];
    12: op1_09_in17 = reg_0355;
    27: op1_09_in17 = reg_0355;
    13: op1_09_in17 = reg_0343;
    14: op1_09_in17 = reg_0526;
    15: op1_09_in17 = reg_0198;
    16: op1_09_in17 = reg_0097;
    17: op1_09_in17 = reg_0202;
    18: op1_09_in17 = reg_0650;
    19: op1_09_in17 = imem01_in[27:24];
    20: op1_09_in17 = reg_0588;
    21: op1_09_in17 = reg_0172;
    22: op1_09_in17 = reg_0707;
    23: op1_09_in17 = imem07_in[111:108];
    24: op1_09_in17 = reg_0205;
    25: op1_09_in17 = reg_0068;
    26: op1_09_in17 = reg_0215;
    72: op1_09_in17 = reg_0215;
    28: op1_09_in17 = reg_0450;
    29: op1_09_in17 = imem01_in[75:72];
    30: op1_09_in17 = reg_0367;
    31: op1_09_in17 = reg_0484;
    32: op1_09_in17 = imem07_in[23:20];
    33: op1_09_in17 = imem01_in[67:64];
    34: op1_09_in17 = imem05_in[87:84];
    35: op1_09_in17 = imem05_in[95:92];
    36: op1_09_in17 = reg_0612;
    37: op1_09_in17 = reg_0298;
    38: op1_09_in17 = reg_0709;
    39: op1_09_in17 = reg_0502;
    40: op1_09_in17 = reg_0246;
    41: op1_09_in17 = imem05_in[115:112];
    42: op1_09_in17 = imem06_in[15:12];
    44: op1_09_in17 = imem03_in[67:64];
    45: op1_09_in17 = reg_0280;
    46: op1_09_in17 = reg_0439;
    47: op1_09_in17 = reg_0538;
    48: op1_09_in17 = reg_0611;
    81: op1_09_in17 = reg_0611;
    49: op1_09_in17 = imem02_in[23:20];
    50: op1_09_in17 = reg_0209;
    52: op1_09_in17 = reg_0212;
    53: op1_09_in17 = reg_0451;
    54: op1_09_in17 = imem03_in[123:120];
    55: op1_09_in17 = reg_0751;
    56: op1_09_in17 = imem04_in[75:72];
    57: op1_09_in17 = imem05_in[27:24];
    58: op1_09_in17 = imem05_in[91:88];
    59: op1_09_in17 = reg_0134;
    60: op1_09_in17 = reg_0625;
    61: op1_09_in17 = reg_0157;
    62: op1_09_in17 = imem02_in[115:112];
    63: op1_09_in17 = reg_0324;
    64: op1_09_in17 = imem04_in[7:4];
    65: op1_09_in17 = reg_0079;
    66: op1_09_in17 = reg_0552;
    67: op1_09_in17 = imem07_in[71:68];
    68: op1_09_in17 = reg_0734;
    69: op1_09_in17 = reg_0259;
    70: op1_09_in17 = reg_0238;
    71: op1_09_in17 = imem02_in[99:96];
    73: op1_09_in17 = reg_0529;
    74: op1_09_in17 = reg_0652;
    76: op1_09_in17 = reg_0759;
    77: op1_09_in17 = reg_0085;
    78: op1_09_in17 = reg_0548;
    79: op1_09_in17 = reg_0337;
    80: op1_09_in17 = imem06_in[83:80];
    82: op1_09_in17 = reg_0703;
    83: op1_09_in17 = reg_0175;
    84: op1_09_in17 = reg_0174;
    85: op1_09_in17 = reg_0618;
    86: op1_09_in17 = reg_0186;
    87: op1_09_in17 = imem03_in[7:4];
    88: op1_09_in17 = reg_0112;
    89: op1_09_in17 = imem03_in[51:48];
    90: op1_09_in17 = reg_0387;
    91: op1_09_in17 = reg_0500;
    92: op1_09_in17 = reg_0440;
    93: op1_09_in17 = imem07_in[47:44];
    94: op1_09_in17 = reg_0161;
    95: op1_09_in17 = reg_0473;
    96: op1_09_in17 = reg_0813;
    default: op1_09_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv17 = 1;
    7: op1_09_inv17 = 1;
    8: op1_09_inv17 = 1;
    11: op1_09_inv17 = 1;
    12: op1_09_inv17 = 1;
    14: op1_09_inv17 = 1;
    15: op1_09_inv17 = 1;
    16: op1_09_inv17 = 1;
    17: op1_09_inv17 = 1;
    18: op1_09_inv17 = 1;
    19: op1_09_inv17 = 1;
    20: op1_09_inv17 = 1;
    22: op1_09_inv17 = 1;
    23: op1_09_inv17 = 1;
    24: op1_09_inv17 = 1;
    25: op1_09_inv17 = 1;
    26: op1_09_inv17 = 1;
    27: op1_09_inv17 = 1;
    28: op1_09_inv17 = 1;
    34: op1_09_inv17 = 1;
    35: op1_09_inv17 = 1;
    37: op1_09_inv17 = 1;
    40: op1_09_inv17 = 1;
    42: op1_09_inv17 = 1;
    45: op1_09_inv17 = 1;
    46: op1_09_inv17 = 1;
    47: op1_09_inv17 = 1;
    49: op1_09_inv17 = 1;
    52: op1_09_inv17 = 1;
    54: op1_09_inv17 = 1;
    55: op1_09_inv17 = 1;
    56: op1_09_inv17 = 1;
    57: op1_09_inv17 = 1;
    59: op1_09_inv17 = 1;
    61: op1_09_inv17 = 1;
    65: op1_09_inv17 = 1;
    67: op1_09_inv17 = 1;
    70: op1_09_inv17 = 1;
    71: op1_09_inv17 = 1;
    72: op1_09_inv17 = 1;
    76: op1_09_inv17 = 1;
    77: op1_09_inv17 = 1;
    78: op1_09_inv17 = 1;
    81: op1_09_inv17 = 1;
    87: op1_09_inv17 = 1;
    89: op1_09_inv17 = 1;
    92: op1_09_inv17 = 1;
    93: op1_09_inv17 = 1;
    95: op1_09_inv17 = 1;
    96: op1_09_inv17 = 1;
    default: op1_09_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の18番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in18 = reg_0381;
    6: op1_09_in18 = reg_0503;
    7: op1_09_in18 = reg_0555;
    8: op1_09_in18 = reg_0442;
    9: op1_09_in18 = reg_0142;
    10: op1_09_in18 = reg_0744;
    11: op1_09_in18 = imem05_in[87:84];
    12: op1_09_in18 = reg_0350;
    13: op1_09_in18 = reg_0396;
    14: op1_09_in18 = reg_0230;
    15: op1_09_in18 = imem01_in[7:4];
    16: op1_09_in18 = reg_0082;
    17: op1_09_in18 = imem01_in[67:64];
    18: op1_09_in18 = reg_0658;
    19: op1_09_in18 = imem01_in[47:44];
    20: op1_09_in18 = reg_0388;
    21: op1_09_in18 = reg_0179;
    22: op1_09_in18 = reg_0426;
    23: op1_09_in18 = reg_0720;
    24: op1_09_in18 = reg_0199;
    25: op1_09_in18 = reg_0072;
    26: op1_09_in18 = reg_0246;
    72: op1_09_in18 = reg_0246;
    27: op1_09_in18 = reg_0539;
    28: op1_09_in18 = reg_0464;
    29: op1_09_in18 = imem01_in[87:84];
    30: op1_09_in18 = reg_0339;
    85: op1_09_in18 = reg_0339;
    31: op1_09_in18 = reg_0788;
    32: op1_09_in18 = imem07_in[39:36];
    33: op1_09_in18 = imem01_in[79:76];
    34: op1_09_in18 = imem05_in[99:96];
    35: op1_09_in18 = reg_0483;
    36: op1_09_in18 = reg_0402;
    37: op1_09_in18 = reg_0266;
    38: op1_09_in18 = reg_0701;
    39: op1_09_in18 = reg_0513;
    40: op1_09_in18 = reg_0245;
    41: op1_09_in18 = reg_0482;
    42: op1_09_in18 = imem06_in[19:16];
    44: op1_09_in18 = imem03_in[79:76];
    45: op1_09_in18 = reg_0076;
    46: op1_09_in18 = reg_0449;
    47: op1_09_in18 = reg_0093;
    48: op1_09_in18 = reg_0077;
    49: op1_09_in18 = imem02_in[95:92];
    50: op1_09_in18 = reg_0188;
    52: op1_09_in18 = reg_0197;
    53: op1_09_in18 = reg_0469;
    54: op1_09_in18 = imem03_in[127:124];
    55: op1_09_in18 = reg_0331;
    56: op1_09_in18 = imem04_in[79:76];
    57: op1_09_in18 = imem05_in[47:44];
    58: op1_09_in18 = imem05_in[111:108];
    59: op1_09_in18 = reg_0144;
    60: op1_09_in18 = reg_0618;
    62: op1_09_in18 = imem02_in[127:124];
    63: op1_09_in18 = reg_0514;
    64: op1_09_in18 = imem04_in[43:40];
    65: op1_09_in18 = reg_0283;
    66: op1_09_in18 = reg_0055;
    67: op1_09_in18 = imem07_in[87:84];
    68: op1_09_in18 = reg_0557;
    69: op1_09_in18 = reg_0233;
    70: op1_09_in18 = reg_0659;
    71: op1_09_in18 = reg_0362;
    73: op1_09_in18 = reg_0616;
    74: op1_09_in18 = reg_0787;
    76: op1_09_in18 = reg_0778;
    77: op1_09_in18 = reg_0111;
    78: op1_09_in18 = reg_0427;
    79: op1_09_in18 = reg_0145;
    80: op1_09_in18 = imem06_in[87:84];
    81: op1_09_in18 = reg_0508;
    82: op1_09_in18 = reg_0485;
    83: op1_09_in18 = reg_0236;
    84: op1_09_in18 = reg_0079;
    86: op1_09_in18 = reg_0198;
    87: op1_09_in18 = reg_0384;
    88: op1_09_in18 = reg_0114;
    89: op1_09_in18 = imem03_in[59:56];
    90: op1_09_in18 = reg_0747;
    91: op1_09_in18 = reg_0252;
    92: op1_09_in18 = reg_0267;
    93: op1_09_in18 = imem07_in[51:48];
    94: op1_09_in18 = reg_0725;
    95: op1_09_in18 = reg_0470;
    96: op1_09_in18 = reg_0664;
    default: op1_09_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_09_inv18 = 1;
    8: op1_09_inv18 = 1;
    12: op1_09_inv18 = 1;
    13: op1_09_inv18 = 1;
    16: op1_09_inv18 = 1;
    17: op1_09_inv18 = 1;
    23: op1_09_inv18 = 1;
    24: op1_09_inv18 = 1;
    26: op1_09_inv18 = 1;
    27: op1_09_inv18 = 1;
    28: op1_09_inv18 = 1;
    29: op1_09_inv18 = 1;
    30: op1_09_inv18 = 1;
    31: op1_09_inv18 = 1;
    35: op1_09_inv18 = 1;
    36: op1_09_inv18 = 1;
    37: op1_09_inv18 = 1;
    38: op1_09_inv18 = 1;
    39: op1_09_inv18 = 1;
    42: op1_09_inv18 = 1;
    44: op1_09_inv18 = 1;
    47: op1_09_inv18 = 1;
    48: op1_09_inv18 = 1;
    52: op1_09_inv18 = 1;
    53: op1_09_inv18 = 1;
    54: op1_09_inv18 = 1;
    56: op1_09_inv18 = 1;
    57: op1_09_inv18 = 1;
    58: op1_09_inv18 = 1;
    59: op1_09_inv18 = 1;
    60: op1_09_inv18 = 1;
    63: op1_09_inv18 = 1;
    64: op1_09_inv18 = 1;
    66: op1_09_inv18 = 1;
    69: op1_09_inv18 = 1;
    71: op1_09_inv18 = 1;
    72: op1_09_inv18 = 1;
    73: op1_09_inv18 = 1;
    77: op1_09_inv18 = 1;
    80: op1_09_inv18 = 1;
    83: op1_09_inv18 = 1;
    85: op1_09_inv18 = 1;
    87: op1_09_inv18 = 1;
    90: op1_09_inv18 = 1;
    92: op1_09_inv18 = 1;
    95: op1_09_inv18 = 1;
    96: op1_09_inv18 = 1;
    default: op1_09_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の19番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in19 = reg_0392;
    6: op1_09_in19 = reg_0506;
    7: op1_09_in19 = reg_0540;
    8: op1_09_in19 = reg_0443;
    9: op1_09_in19 = reg_0143;
    10: op1_09_in19 = reg_0228;
    11: op1_09_in19 = imem05_in[107:104];
    12: op1_09_in19 = reg_0347;
    13: op1_09_in19 = reg_0000;
    14: op1_09_in19 = reg_0732;
    15: op1_09_in19 = imem01_in[11:8];
    16: op1_09_in19 = reg_0084;
    46: op1_09_in19 = reg_0084;
    17: op1_09_in19 = imem01_in[71:68];
    19: op1_09_in19 = imem01_in[71:68];
    18: op1_09_in19 = reg_0653;
    20: op1_09_in19 = reg_0369;
    21: op1_09_in19 = reg_0161;
    22: op1_09_in19 = reg_0419;
    23: op1_09_in19 = reg_0710;
    24: op1_09_in19 = reg_0197;
    25: op1_09_in19 = reg_0256;
    26: op1_09_in19 = reg_0105;
    27: op1_09_in19 = reg_0756;
    28: op1_09_in19 = reg_0480;
    29: op1_09_in19 = imem01_in[91:88];
    30: op1_09_in19 = reg_0375;
    31: op1_09_in19 = reg_0790;
    32: op1_09_in19 = imem07_in[75:72];
    33: op1_09_in19 = reg_0549;
    34: op1_09_in19 = imem05_in[123:120];
    35: op1_09_in19 = reg_0788;
    36: op1_09_in19 = reg_0407;
    37: op1_09_in19 = reg_0278;
    38: op1_09_in19 = reg_0727;
    39: op1_09_in19 = reg_0772;
    40: op1_09_in19 = reg_0249;
    41: op1_09_in19 = reg_0797;
    42: op1_09_in19 = imem06_in[39:36];
    44: op1_09_in19 = imem03_in[91:88];
    45: op1_09_in19 = reg_0631;
    47: op1_09_in19 = imem03_in[19:16];
    48: op1_09_in19 = reg_0626;
    65: op1_09_in19 = reg_0626;
    49: op1_09_in19 = imem02_in[123:120];
    50: op1_09_in19 = reg_0193;
    52: op1_09_in19 = reg_0111;
    53: op1_09_in19 = reg_0472;
    54: op1_09_in19 = reg_0394;
    55: op1_09_in19 = reg_0568;
    56: op1_09_in19 = imem04_in[91:88];
    57: op1_09_in19 = imem05_in[67:64];
    58: op1_09_in19 = reg_0781;
    59: op1_09_in19 = imem06_in[7:4];
    60: op1_09_in19 = reg_0031;
    62: op1_09_in19 = reg_0587;
    63: op1_09_in19 = reg_0541;
    64: op1_09_in19 = imem04_in[51:48];
    66: op1_09_in19 = reg_0060;
    67: op1_09_in19 = imem07_in[107:104];
    68: op1_09_in19 = reg_0652;
    69: op1_09_in19 = reg_0416;
    70: op1_09_in19 = reg_0654;
    71: op1_09_in19 = reg_0514;
    72: op1_09_in19 = reg_0279;
    73: op1_09_in19 = reg_0292;
    74: op1_09_in19 = reg_0716;
    76: op1_09_in19 = reg_0237;
    77: op1_09_in19 = reg_0112;
    78: op1_09_in19 = reg_0352;
    79: op1_09_in19 = reg_0135;
    80: op1_09_in19 = imem06_in[107:104];
    81: op1_09_in19 = reg_0617;
    82: op1_09_in19 = reg_0320;
    83: op1_09_in19 = reg_0066;
    84: op1_09_in19 = reg_0433;
    85: op1_09_in19 = reg_0265;
    86: op1_09_in19 = reg_0212;
    87: op1_09_in19 = reg_0028;
    88: op1_09_in19 = reg_0759;
    89: op1_09_in19 = imem03_in[75:72];
    90: op1_09_in19 = reg_0319;
    91: op1_09_in19 = reg_0491;
    92: op1_09_in19 = reg_0438;
    93: op1_09_in19 = imem07_in[111:108];
    94: op1_09_in19 = reg_0713;
    95: op1_09_in19 = reg_0471;
    96: op1_09_in19 = reg_0661;
    default: op1_09_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv19 = 1;
    9: op1_09_inv19 = 1;
    10: op1_09_inv19 = 1;
    11: op1_09_inv19 = 1;
    12: op1_09_inv19 = 1;
    13: op1_09_inv19 = 1;
    14: op1_09_inv19 = 1;
    18: op1_09_inv19 = 1;
    20: op1_09_inv19 = 1;
    21: op1_09_inv19 = 1;
    25: op1_09_inv19 = 1;
    26: op1_09_inv19 = 1;
    27: op1_09_inv19 = 1;
    28: op1_09_inv19 = 1;
    29: op1_09_inv19 = 1;
    30: op1_09_inv19 = 1;
    31: op1_09_inv19 = 1;
    32: op1_09_inv19 = 1;
    34: op1_09_inv19 = 1;
    35: op1_09_inv19 = 1;
    38: op1_09_inv19 = 1;
    39: op1_09_inv19 = 1;
    40: op1_09_inv19 = 1;
    41: op1_09_inv19 = 1;
    44: op1_09_inv19 = 1;
    45: op1_09_inv19 = 1;
    46: op1_09_inv19 = 1;
    48: op1_09_inv19 = 1;
    53: op1_09_inv19 = 1;
    55: op1_09_inv19 = 1;
    58: op1_09_inv19 = 1;
    59: op1_09_inv19 = 1;
    60: op1_09_inv19 = 1;
    62: op1_09_inv19 = 1;
    63: op1_09_inv19 = 1;
    69: op1_09_inv19 = 1;
    71: op1_09_inv19 = 1;
    76: op1_09_inv19 = 1;
    77: op1_09_inv19 = 1;
    78: op1_09_inv19 = 1;
    79: op1_09_inv19 = 1;
    80: op1_09_inv19 = 1;
    85: op1_09_inv19 = 1;
    86: op1_09_inv19 = 1;
    87: op1_09_inv19 = 1;
    92: op1_09_inv19 = 1;
    94: op1_09_inv19 = 1;
    default: op1_09_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の20番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in20 = reg_0371;
    6: op1_09_in20 = reg_0233;
    7: op1_09_in20 = reg_0532;
    8: op1_09_in20 = reg_0435;
    9: op1_09_in20 = reg_0134;
    10: op1_09_in20 = reg_0737;
    11: op1_09_in20 = reg_0147;
    12: op1_09_in20 = reg_0083;
    13: op1_09_in20 = reg_0801;
    14: op1_09_in20 = reg_0744;
    15: op1_09_in20 = imem01_in[39:36];
    16: op1_09_in20 = reg_0079;
    17: op1_09_in20 = imem01_in[87:84];
    18: op1_09_in20 = reg_0637;
    19: op1_09_in20 = imem01_in[107:104];
    20: op1_09_in20 = reg_0377;
    21: op1_09_in20 = reg_0182;
    22: op1_09_in20 = reg_0439;
    23: op1_09_in20 = reg_0706;
    24: op1_09_in20 = reg_0229;
    25: op1_09_in20 = imem05_in[59:56];
    26: op1_09_in20 = reg_0107;
    27: op1_09_in20 = reg_0526;
    28: op1_09_in20 = reg_0470;
    29: op1_09_in20 = imem01_in[111:108];
    30: op1_09_in20 = imem03_in[3:0];
    63: op1_09_in20 = imem03_in[3:0];
    31: op1_09_in20 = reg_0271;
    32: op1_09_in20 = imem07_in[87:84];
    33: op1_09_in20 = reg_0515;
    34: op1_09_in20 = reg_0490;
    58: op1_09_in20 = reg_0490;
    35: op1_09_in20 = reg_0785;
    36: op1_09_in20 = reg_0270;
    37: op1_09_in20 = reg_0063;
    38: op1_09_in20 = reg_0441;
    39: op1_09_in20 = reg_0514;
    40: op1_09_in20 = reg_0758;
    41: op1_09_in20 = reg_0488;
    42: op1_09_in20 = imem06_in[43:40];
    44: op1_09_in20 = imem03_in[123:120];
    45: op1_09_in20 = reg_0071;
    46: op1_09_in20 = reg_0175;
    47: op1_09_in20 = imem03_in[67:64];
    48: op1_09_in20 = imem04_in[3:0];
    49: op1_09_in20 = reg_0656;
    50: op1_09_in20 = reg_0207;
    52: op1_09_in20 = reg_0509;
    53: op1_09_in20 = reg_0480;
    54: op1_09_in20 = reg_0384;
    55: op1_09_in20 = reg_0386;
    56: op1_09_in20 = imem04_in[111:108];
    57: op1_09_in20 = imem05_in[83:80];
    59: op1_09_in20 = imem06_in[31:28];
    60: op1_09_in20 = reg_0580;
    62: op1_09_in20 = reg_0358;
    78: op1_09_in20 = reg_0358;
    64: op1_09_in20 = imem04_in[55:52];
    65: op1_09_in20 = reg_0614;
    81: op1_09_in20 = reg_0614;
    66: op1_09_in20 = reg_0057;
    67: op1_09_in20 = reg_0719;
    68: op1_09_in20 = imem01_in[15:12];
    69: op1_09_in20 = imem05_in[7:4];
    70: op1_09_in20 = reg_0375;
    71: op1_09_in20 = reg_0533;
    72: op1_09_in20 = reg_0040;
    73: op1_09_in20 = reg_0508;
    74: op1_09_in20 = reg_0089;
    76: op1_09_in20 = reg_0388;
    77: op1_09_in20 = reg_0397;
    79: op1_09_in20 = reg_0090;
    80: op1_09_in20 = imem06_in[115:112];
    82: op1_09_in20 = reg_0581;
    83: op1_09_in20 = reg_0183;
    84: op1_09_in20 = reg_0616;
    85: op1_09_in20 = reg_0401;
    86: op1_09_in20 = imem01_in[47:44];
    87: op1_09_in20 = reg_0570;
    88: op1_09_in20 = reg_0778;
    89: op1_09_in20 = imem03_in[99:96];
    90: op1_09_in20 = reg_0800;
    91: op1_09_in20 = reg_0531;
    92: op1_09_in20 = reg_0116;
    93: op1_09_in20 = imem07_in[119:116];
    94: op1_09_in20 = reg_0724;
    95: op1_09_in20 = reg_0208;
    96: op1_09_in20 = imem07_in[43:40];
    default: op1_09_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv20 = 1;
    8: op1_09_inv20 = 1;
    11: op1_09_inv20 = 1;
    12: op1_09_inv20 = 1;
    13: op1_09_inv20 = 1;
    14: op1_09_inv20 = 1;
    15: op1_09_inv20 = 1;
    16: op1_09_inv20 = 1;
    18: op1_09_inv20 = 1;
    19: op1_09_inv20 = 1;
    20: op1_09_inv20 = 1;
    24: op1_09_inv20 = 1;
    26: op1_09_inv20 = 1;
    28: op1_09_inv20 = 1;
    33: op1_09_inv20 = 1;
    35: op1_09_inv20 = 1;
    38: op1_09_inv20 = 1;
    45: op1_09_inv20 = 1;
    48: op1_09_inv20 = 1;
    49: op1_09_inv20 = 1;
    50: op1_09_inv20 = 1;
    52: op1_09_inv20 = 1;
    56: op1_09_inv20 = 1;
    57: op1_09_inv20 = 1;
    62: op1_09_inv20 = 1;
    63: op1_09_inv20 = 1;
    64: op1_09_inv20 = 1;
    65: op1_09_inv20 = 1;
    66: op1_09_inv20 = 1;
    69: op1_09_inv20 = 1;
    71: op1_09_inv20 = 1;
    72: op1_09_inv20 = 1;
    77: op1_09_inv20 = 1;
    81: op1_09_inv20 = 1;
    82: op1_09_inv20 = 1;
    83: op1_09_inv20 = 1;
    85: op1_09_inv20 = 1;
    86: op1_09_inv20 = 1;
    89: op1_09_inv20 = 1;
    92: op1_09_inv20 = 1;
    93: op1_09_inv20 = 1;
    94: op1_09_inv20 = 1;
    default: op1_09_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の21番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in21 = reg_0390;
    6: op1_09_in21 = reg_0218;
    7: op1_09_in21 = reg_0301;
    8: op1_09_in21 = reg_0181;
    92: op1_09_in21 = reg_0181;
    9: op1_09_in21 = imem06_in[7:4];
    10: op1_09_in21 = reg_0498;
    11: op1_09_in21 = reg_0151;
    91: op1_09_in21 = reg_0151;
    12: op1_09_in21 = reg_0092;
    13: op1_09_in21 = imem04_in[95:92];
    14: op1_09_in21 = reg_0734;
    15: op1_09_in21 = imem01_in[47:44];
    68: op1_09_in21 = imem01_in[47:44];
    16: op1_09_in21 = imem03_in[39:36];
    17: op1_09_in21 = imem01_in[95:92];
    18: op1_09_in21 = reg_0648;
    19: op1_09_in21 = reg_0523;
    20: op1_09_in21 = reg_0803;
    21: op1_09_in21 = reg_0163;
    22: op1_09_in21 = reg_0428;
    23: op1_09_in21 = reg_0429;
    24: op1_09_in21 = reg_0322;
    25: op1_09_in21 = reg_0484;
    26: op1_09_in21 = reg_0113;
    27: op1_09_in21 = reg_0740;
    28: op1_09_in21 = reg_0459;
    29: op1_09_in21 = reg_0497;
    30: op1_09_in21 = imem03_in[47:44];
    31: op1_09_in21 = reg_0304;
    32: op1_09_in21 = imem07_in[111:108];
    33: op1_09_in21 = reg_0548;
    34: op1_09_in21 = reg_0492;
    35: op1_09_in21 = reg_0784;
    36: op1_09_in21 = reg_0776;
    37: op1_09_in21 = imem05_in[11:8];
    38: op1_09_in21 = reg_0445;
    39: op1_09_in21 = reg_0334;
    40: op1_09_in21 = reg_0514;
    41: op1_09_in21 = reg_0491;
    42: op1_09_in21 = imem06_in[67:64];
    44: op1_09_in21 = reg_0599;
    45: op1_09_in21 = reg_0292;
    84: op1_09_in21 = reg_0292;
    46: op1_09_in21 = reg_0179;
    47: op1_09_in21 = imem03_in[87:84];
    48: op1_09_in21 = imem04_in[11:8];
    49: op1_09_in21 = reg_0346;
    50: op1_09_in21 = reg_0196;
    52: op1_09_in21 = reg_0771;
    53: op1_09_in21 = reg_0471;
    54: op1_09_in21 = reg_0755;
    55: op1_09_in21 = reg_0019;
    56: op1_09_in21 = reg_0544;
    57: op1_09_in21 = imem05_in[103:100];
    58: op1_09_in21 = reg_0110;
    59: op1_09_in21 = imem06_in[59:56];
    60: op1_09_in21 = imem06_in[3:0];
    62: op1_09_in21 = reg_0353;
    63: op1_09_in21 = imem03_in[19:16];
    64: op1_09_in21 = imem04_in[87:84];
    65: op1_09_in21 = reg_0679;
    66: op1_09_in21 = reg_0536;
    67: op1_09_in21 = reg_0726;
    69: op1_09_in21 = imem05_in[91:88];
    70: op1_09_in21 = imem06_in[19:16];
    71: op1_09_in21 = reg_0540;
    72: op1_09_in21 = reg_0276;
    73: op1_09_in21 = reg_0614;
    74: op1_09_in21 = reg_0710;
    76: op1_09_in21 = reg_0225;
    77: op1_09_in21 = reg_0423;
    78: op1_09_in21 = reg_0320;
    79: op1_09_in21 = reg_0732;
    80: op1_09_in21 = reg_0348;
    81: op1_09_in21 = reg_0598;
    82: op1_09_in21 = reg_0341;
    83: op1_09_in21 = reg_0100;
    85: op1_09_in21 = imem06_in[23:20];
    86: op1_09_in21 = imem01_in[91:88];
    87: op1_09_in21 = reg_0006;
    88: op1_09_in21 = reg_0388;
    89: op1_09_in21 = imem04_in[3:0];
    90: op1_09_in21 = reg_0809;
    93: op1_09_in21 = reg_0716;
    94: op1_09_in21 = reg_0253;
    95: op1_09_in21 = reg_0204;
    96: op1_09_in21 = imem07_in[87:84];
    default: op1_09_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_09_inv21 = 1;
    14: op1_09_inv21 = 1;
    16: op1_09_inv21 = 1;
    20: op1_09_inv21 = 1;
    21: op1_09_inv21 = 1;
    24: op1_09_inv21 = 1;
    25: op1_09_inv21 = 1;
    32: op1_09_inv21 = 1;
    34: op1_09_inv21 = 1;
    35: op1_09_inv21 = 1;
    38: op1_09_inv21 = 1;
    39: op1_09_inv21 = 1;
    40: op1_09_inv21 = 1;
    41: op1_09_inv21 = 1;
    44: op1_09_inv21 = 1;
    45: op1_09_inv21 = 1;
    46: op1_09_inv21 = 1;
    47: op1_09_inv21 = 1;
    49: op1_09_inv21 = 1;
    57: op1_09_inv21 = 1;
    58: op1_09_inv21 = 1;
    59: op1_09_inv21 = 1;
    60: op1_09_inv21 = 1;
    62: op1_09_inv21 = 1;
    65: op1_09_inv21 = 1;
    66: op1_09_inv21 = 1;
    67: op1_09_inv21 = 1;
    68: op1_09_inv21 = 1;
    69: op1_09_inv21 = 1;
    70: op1_09_inv21 = 1;
    72: op1_09_inv21 = 1;
    73: op1_09_inv21 = 1;
    77: op1_09_inv21 = 1;
    79: op1_09_inv21 = 1;
    80: op1_09_inv21 = 1;
    86: op1_09_inv21 = 1;
    88: op1_09_inv21 = 1;
    89: op1_09_inv21 = 1;
    90: op1_09_inv21 = 1;
    92: op1_09_inv21 = 1;
    94: op1_09_inv21 = 1;
    95: op1_09_inv21 = 1;
    96: op1_09_inv21 = 1;
    default: op1_09_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の22番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in22 = reg_0367;
    6: op1_09_in22 = reg_0245;
    7: op1_09_in22 = reg_0279;
    83: op1_09_in22 = reg_0279;
    8: op1_09_in22 = reg_0162;
    9: op1_09_in22 = imem06_in[23:20];
    10: op1_09_in22 = reg_0740;
    11: op1_09_in22 = reg_0153;
    12: op1_09_in22 = reg_0049;
    13: op1_09_in22 = imem04_in[107:104];
    14: op1_09_in22 = reg_0148;
    15: op1_09_in22 = imem01_in[51:48];
    68: op1_09_in22 = imem01_in[51:48];
    16: op1_09_in22 = imem03_in[63:60];
    17: op1_09_in22 = imem01_in[99:96];
    18: op1_09_in22 = reg_0638;
    19: op1_09_in22 = reg_0513;
    20: op1_09_in22 = reg_0008;
    21: op1_09_in22 = reg_0178;
    22: op1_09_in22 = reg_0431;
    45: op1_09_in22 = reg_0431;
    23: op1_09_in22 = reg_0418;
    77: op1_09_in22 = reg_0418;
    24: op1_09_in22 = reg_0323;
    25: op1_09_in22 = reg_0789;
    26: op1_09_in22 = imem02_in[31:28];
    27: op1_09_in22 = reg_0317;
    28: op1_09_in22 = reg_0208;
    29: op1_09_in22 = reg_0822;
    30: op1_09_in22 = imem03_in[55:52];
    31: op1_09_in22 = reg_0309;
    32: op1_09_in22 = imem07_in[119:116];
    33: op1_09_in22 = reg_0550;
    34: op1_09_in22 = reg_0793;
    35: op1_09_in22 = reg_0485;
    36: op1_09_in22 = reg_0319;
    37: op1_09_in22 = imem05_in[15:12];
    38: op1_09_in22 = reg_0438;
    39: op1_09_in22 = reg_0515;
    40: op1_09_in22 = reg_0824;
    41: op1_09_in22 = reg_0492;
    42: op1_09_in22 = imem06_in[103:100];
    44: op1_09_in22 = reg_0583;
    46: op1_09_in22 = reg_0168;
    47: op1_09_in22 = imem03_in[115:112];
    48: op1_09_in22 = imem04_in[27:24];
    49: op1_09_in22 = reg_0355;
    50: op1_09_in22 = imem01_in[27:24];
    52: op1_09_in22 = reg_0113;
    53: op1_09_in22 = reg_0209;
    54: op1_09_in22 = reg_0376;
    55: op1_09_in22 = reg_0012;
    56: op1_09_in22 = reg_0553;
    57: op1_09_in22 = imem05_in[107:104];
    69: op1_09_in22 = imem05_in[107:104];
    58: op1_09_in22 = reg_0099;
    59: op1_09_in22 = imem06_in[71:68];
    60: op1_09_in22 = imem06_in[19:16];
    62: op1_09_in22 = reg_0365;
    63: op1_09_in22 = imem03_in[39:36];
    64: op1_09_in22 = imem04_in[103:100];
    65: op1_09_in22 = reg_0301;
    66: op1_09_in22 = reg_0516;
    67: op1_09_in22 = reg_0727;
    70: op1_09_in22 = imem06_in[27:24];
    71: op1_09_in22 = reg_0770;
    72: op1_09_in22 = reg_0786;
    73: op1_09_in22 = reg_0598;
    74: op1_09_in22 = reg_0712;
    76: op1_09_in22 = reg_0240;
    78: op1_09_in22 = reg_0360;
    79: op1_09_in22 = reg_0226;
    80: op1_09_in22 = reg_0349;
    81: op1_09_in22 = reg_0643;
    82: op1_09_in22 = reg_0353;
    84: op1_09_in22 = reg_0627;
    85: op1_09_in22 = imem06_in[43:40];
    86: op1_09_in22 = reg_0772;
    87: op1_09_in22 = reg_0805;
    88: op1_09_in22 = reg_0258;
    89: op1_09_in22 = imem04_in[31:28];
    90: op1_09_in22 = imem04_in[3:0];
    91: op1_09_in22 = reg_0830;
    92: op1_09_in22 = reg_0183;
    93: op1_09_in22 = reg_0711;
    94: op1_09_in22 = reg_0067;
    95: op1_09_in22 = reg_0203;
    96: op1_09_in22 = imem07_in[99:96];
    default: op1_09_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv22 = 1;
    8: op1_09_inv22 = 1;
    10: op1_09_inv22 = 1;
    12: op1_09_inv22 = 1;
    15: op1_09_inv22 = 1;
    16: op1_09_inv22 = 1;
    18: op1_09_inv22 = 1;
    24: op1_09_inv22 = 1;
    26: op1_09_inv22 = 1;
    28: op1_09_inv22 = 1;
    30: op1_09_inv22 = 1;
    31: op1_09_inv22 = 1;
    33: op1_09_inv22 = 1;
    34: op1_09_inv22 = 1;
    35: op1_09_inv22 = 1;
    38: op1_09_inv22 = 1;
    39: op1_09_inv22 = 1;
    40: op1_09_inv22 = 1;
    41: op1_09_inv22 = 1;
    44: op1_09_inv22 = 1;
    47: op1_09_inv22 = 1;
    48: op1_09_inv22 = 1;
    55: op1_09_inv22 = 1;
    56: op1_09_inv22 = 1;
    58: op1_09_inv22 = 1;
    59: op1_09_inv22 = 1;
    60: op1_09_inv22 = 1;
    62: op1_09_inv22 = 1;
    63: op1_09_inv22 = 1;
    64: op1_09_inv22 = 1;
    66: op1_09_inv22 = 1;
    68: op1_09_inv22 = 1;
    69: op1_09_inv22 = 1;
    72: op1_09_inv22 = 1;
    84: op1_09_inv22 = 1;
    85: op1_09_inv22 = 1;
    86: op1_09_inv22 = 1;
    89: op1_09_inv22 = 1;
    91: op1_09_inv22 = 1;
    93: op1_09_inv22 = 1;
    96: op1_09_inv22 = 1;
    default: op1_09_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の23番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in23 = reg_0035;
    6: op1_09_in23 = reg_0219;
    7: op1_09_in23 = reg_0293;
    8: op1_09_in23 = reg_0182;
    9: op1_09_in23 = imem06_in[55:52];
    10: op1_09_in23 = reg_0505;
    11: op1_09_in23 = imem06_in[43:40];
    12: op1_09_in23 = reg_0087;
    13: op1_09_in23 = reg_0560;
    14: op1_09_in23 = reg_0128;
    15: op1_09_in23 = imem01_in[63:60];
    16: op1_09_in23 = imem03_in[79:76];
    17: op1_09_in23 = imem01_in[111:108];
    18: op1_09_in23 = reg_0659;
    19: op1_09_in23 = reg_0820;
    20: op1_09_in23 = reg_0806;
    21: op1_09_in23 = reg_0157;
    22: op1_09_in23 = reg_0165;
    23: op1_09_in23 = reg_0442;
    24: op1_09_in23 = imem01_in[35:32];
    25: op1_09_in23 = reg_0780;
    41: op1_09_in23 = reg_0780;
    26: op1_09_in23 = imem02_in[107:104];
    27: op1_09_in23 = reg_0259;
    28: op1_09_in23 = reg_0201;
    29: op1_09_in23 = reg_0514;
    30: op1_09_in23 = imem03_in[99:96];
    31: op1_09_in23 = reg_0282;
    32: op1_09_in23 = imem07_in[123:120];
    33: op1_09_in23 = reg_0235;
    34: op1_09_in23 = reg_0494;
    35: op1_09_in23 = reg_0486;
    36: op1_09_in23 = reg_0764;
    37: op1_09_in23 = imem05_in[19:16];
    38: op1_09_in23 = reg_0175;
    39: op1_09_in23 = imem01_in[75:72];
    40: op1_09_in23 = reg_0519;
    42: op1_09_in23 = imem06_in[119:116];
    44: op1_09_in23 = reg_0592;
    45: op1_09_in23 = imem04_in[7:4];
    46: op1_09_in23 = reg_0170;
    92: op1_09_in23 = reg_0170;
    47: op1_09_in23 = reg_0598;
    48: op1_09_in23 = imem04_in[67:64];
    49: op1_09_in23 = reg_0665;
    50: op1_09_in23 = imem01_in[79:76];
    52: op1_09_in23 = reg_0117;
    53: op1_09_in23 = reg_0196;
    54: op1_09_in23 = reg_0747;
    55: op1_09_in23 = reg_0015;
    56: op1_09_in23 = reg_0542;
    57: op1_09_in23 = reg_0798;
    58: op1_09_in23 = reg_0269;
    59: op1_09_in23 = imem06_in[83:80];
    60: op1_09_in23 = imem06_in[47:44];
    62: op1_09_in23 = reg_0406;
    63: op1_09_in23 = imem03_in[95:92];
    64: op1_09_in23 = reg_0545;
    65: op1_09_in23 = reg_0622;
    66: op1_09_in23 = reg_0556;
    67: op1_09_in23 = reg_0266;
    68: op1_09_in23 = imem01_in[95:92];
    69: op1_09_in23 = imem05_in[119:116];
    70: op1_09_in23 = imem06_in[31:28];
    71: op1_09_in23 = reg_0539;
    72: op1_09_in23 = reg_0156;
    73: op1_09_in23 = reg_0068;
    74: op1_09_in23 = reg_0713;
    76: op1_09_in23 = reg_0502;
    77: op1_09_in23 = reg_0511;
    78: op1_09_in23 = reg_0527;
    79: op1_09_in23 = reg_0326;
    80: op1_09_in23 = reg_0609;
    81: op1_09_in23 = reg_0774;
    82: op1_09_in23 = reg_0365;
    84: op1_09_in23 = reg_0301;
    85: op1_09_in23 = imem06_in[95:92];
    86: op1_09_in23 = reg_0385;
    87: op1_09_in23 = imem04_in[15:12];
    88: op1_09_in23 = reg_0418;
    89: op1_09_in23 = imem04_in[43:40];
    90: op1_09_in23 = imem04_in[55:52];
    91: op1_09_in23 = reg_0153;
    93: op1_09_in23 = reg_0443;
    94: op1_09_in23 = reg_0635;
    95: op1_09_in23 = reg_0205;
    96: op1_09_in23 = imem07_in[103:100];
    default: op1_09_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv23 = 1;
    7: op1_09_inv23 = 1;
    10: op1_09_inv23 = 1;
    11: op1_09_inv23 = 1;
    14: op1_09_inv23 = 1;
    15: op1_09_inv23 = 1;
    16: op1_09_inv23 = 1;
    17: op1_09_inv23 = 1;
    18: op1_09_inv23 = 1;
    19: op1_09_inv23 = 1;
    21: op1_09_inv23 = 1;
    22: op1_09_inv23 = 1;
    23: op1_09_inv23 = 1;
    26: op1_09_inv23 = 1;
    29: op1_09_inv23 = 1;
    30: op1_09_inv23 = 1;
    31: op1_09_inv23 = 1;
    32: op1_09_inv23 = 1;
    37: op1_09_inv23 = 1;
    38: op1_09_inv23 = 1;
    40: op1_09_inv23 = 1;
    42: op1_09_inv23 = 1;
    44: op1_09_inv23 = 1;
    45: op1_09_inv23 = 1;
    46: op1_09_inv23 = 1;
    49: op1_09_inv23 = 1;
    53: op1_09_inv23 = 1;
    55: op1_09_inv23 = 1;
    58: op1_09_inv23 = 1;
    60: op1_09_inv23 = 1;
    64: op1_09_inv23 = 1;
    65: op1_09_inv23 = 1;
    66: op1_09_inv23 = 1;
    67: op1_09_inv23 = 1;
    68: op1_09_inv23 = 1;
    71: op1_09_inv23 = 1;
    76: op1_09_inv23 = 1;
    78: op1_09_inv23 = 1;
    79: op1_09_inv23 = 1;
    81: op1_09_inv23 = 1;
    90: op1_09_inv23 = 1;
    95: op1_09_inv23 = 1;
    default: op1_09_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の24番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in24 = reg_0020;
    6: op1_09_in24 = reg_0118;
    7: op1_09_in24 = reg_0307;
    8: op1_09_in24 = reg_0183;
    9: op1_09_in24 = imem06_in[75:72];
    10: op1_09_in24 = reg_0215;
    11: op1_09_in24 = imem06_in[51:48];
    12: op1_09_in24 = reg_0073;
    13: op1_09_in24 = reg_0554;
    14: op1_09_in24 = reg_0139;
    15: op1_09_in24 = reg_0522;
    16: op1_09_in24 = reg_0602;
    17: op1_09_in24 = reg_0514;
    78: op1_09_in24 = reg_0514;
    82: op1_09_in24 = reg_0514;
    18: op1_09_in24 = reg_0329;
    19: op1_09_in24 = reg_0824;
    29: op1_09_in24 = reg_0824;
    20: op1_09_in24 = imem04_in[23:20];
    22: op1_09_in24 = reg_0168;
    23: op1_09_in24 = reg_0165;
    24: op1_09_in24 = imem01_in[95:92];
    25: op1_09_in24 = reg_0785;
    26: op1_09_in24 = imem02_in[119:116];
    27: op1_09_in24 = reg_0319;
    28: op1_09_in24 = reg_0212;
    30: op1_09_in24 = imem03_in[115:112];
    31: op1_09_in24 = reg_0277;
    32: op1_09_in24 = imem07_in[127:124];
    33: op1_09_in24 = reg_0241;
    34: op1_09_in24 = reg_0780;
    73: op1_09_in24 = reg_0780;
    35: op1_09_in24 = reg_0225;
    36: op1_09_in24 = imem06_in[67:64];
    37: op1_09_in24 = imem05_in[27:24];
    38: op1_09_in24 = reg_0166;
    39: op1_09_in24 = imem01_in[83:80];
    40: op1_09_in24 = reg_0333;
    41: op1_09_in24 = reg_0091;
    42: op1_09_in24 = reg_0604;
    44: op1_09_in24 = reg_0578;
    45: op1_09_in24 = imem04_in[19:16];
    47: op1_09_in24 = reg_0587;
    48: op1_09_in24 = imem04_in[83:80];
    49: op1_09_in24 = reg_0344;
    50: op1_09_in24 = imem01_in[91:88];
    52: op1_09_in24 = reg_0559;
    53: op1_09_in24 = reg_0205;
    54: op1_09_in24 = reg_0386;
    55: op1_09_in24 = reg_0009;
    56: op1_09_in24 = reg_0056;
    57: op1_09_in24 = reg_0796;
    58: op1_09_in24 = reg_0089;
    59: op1_09_in24 = imem06_in[99:96];
    60: op1_09_in24 = imem06_in[91:88];
    62: op1_09_in24 = reg_0323;
    63: op1_09_in24 = reg_0589;
    64: op1_09_in24 = reg_0315;
    65: op1_09_in24 = reg_0643;
    66: op1_09_in24 = reg_0547;
    67: op1_09_in24 = reg_0436;
    68: op1_09_in24 = imem01_in[99:96];
    69: op1_09_in24 = reg_0788;
    70: op1_09_in24 = imem06_in[43:40];
    71: op1_09_in24 = reg_0538;
    72: op1_09_in24 = reg_0155;
    74: op1_09_in24 = reg_0708;
    76: op1_09_in24 = reg_0505;
    77: op1_09_in24 = reg_0220;
    79: op1_09_in24 = reg_0309;
    80: op1_09_in24 = reg_0606;
    81: op1_09_in24 = reg_0640;
    84: op1_09_in24 = reg_0687;
    85: op1_09_in24 = imem06_in[127:124];
    86: op1_09_in24 = reg_0224;
    87: op1_09_in24 = imem04_in[47:44];
    88: op1_09_in24 = reg_0567;
    89: op1_09_in24 = imem04_in[79:76];
    90: op1_09_in24 = imem04_in[59:56];
    91: op1_09_in24 = reg_0765;
    93: op1_09_in24 = reg_0084;
    94: op1_09_in24 = reg_0445;
    95: op1_09_in24 = reg_0202;
    96: op1_09_in24 = reg_0162;
    default: op1_09_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv24 = 1;
    6: op1_09_inv24 = 1;
    7: op1_09_inv24 = 1;
    8: op1_09_inv24 = 1;
    9: op1_09_inv24 = 1;
    10: op1_09_inv24 = 1;
    11: op1_09_inv24 = 1;
    12: op1_09_inv24 = 1;
    13: op1_09_inv24 = 1;
    14: op1_09_inv24 = 1;
    16: op1_09_inv24 = 1;
    18: op1_09_inv24 = 1;
    19: op1_09_inv24 = 1;
    20: op1_09_inv24 = 1;
    22: op1_09_inv24 = 1;
    24: op1_09_inv24 = 1;
    25: op1_09_inv24 = 1;
    26: op1_09_inv24 = 1;
    27: op1_09_inv24 = 1;
    28: op1_09_inv24 = 1;
    29: op1_09_inv24 = 1;
    30: op1_09_inv24 = 1;
    32: op1_09_inv24 = 1;
    37: op1_09_inv24 = 1;
    38: op1_09_inv24 = 1;
    40: op1_09_inv24 = 1;
    41: op1_09_inv24 = 1;
    42: op1_09_inv24 = 1;
    47: op1_09_inv24 = 1;
    49: op1_09_inv24 = 1;
    50: op1_09_inv24 = 1;
    52: op1_09_inv24 = 1;
    53: op1_09_inv24 = 1;
    54: op1_09_inv24 = 1;
    55: op1_09_inv24 = 1;
    57: op1_09_inv24 = 1;
    59: op1_09_inv24 = 1;
    62: op1_09_inv24 = 1;
    65: op1_09_inv24 = 1;
    66: op1_09_inv24 = 1;
    67: op1_09_inv24 = 1;
    69: op1_09_inv24 = 1;
    72: op1_09_inv24 = 1;
    76: op1_09_inv24 = 1;
    77: op1_09_inv24 = 1;
    78: op1_09_inv24 = 1;
    79: op1_09_inv24 = 1;
    81: op1_09_inv24 = 1;
    84: op1_09_inv24 = 1;
    85: op1_09_inv24 = 1;
    86: op1_09_inv24 = 1;
    87: op1_09_inv24 = 1;
    89: op1_09_inv24 = 1;
    93: op1_09_inv24 = 1;
    95: op1_09_inv24 = 1;
    default: op1_09_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の25番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in25 = reg_0023;
    6: op1_09_in25 = reg_0125;
    7: op1_09_in25 = reg_0059;
    8: op1_09_in25 = reg_0166;
    9: op1_09_in25 = imem06_in[95:92];
    60: op1_09_in25 = imem06_in[95:92];
    10: op1_09_in25 = reg_0504;
    11: op1_09_in25 = imem06_in[63:60];
    12: op1_09_in25 = imem03_in[43:40];
    13: op1_09_in25 = reg_0558;
    14: op1_09_in25 = reg_0140;
    15: op1_09_in25 = reg_0512;
    16: op1_09_in25 = reg_0579;
    17: op1_09_in25 = reg_0227;
    29: op1_09_in25 = reg_0227;
    18: op1_09_in25 = reg_0365;
    19: op1_09_in25 = reg_0521;
    20: op1_09_in25 = imem04_in[75:72];
    22: op1_09_in25 = reg_0170;
    23: op1_09_in25 = reg_0179;
    24: op1_09_in25 = imem01_in[103:100];
    25: op1_09_in25 = reg_0782;
    26: op1_09_in25 = reg_0655;
    27: op1_09_in25 = reg_0318;
    28: op1_09_in25 = imem01_in[11:8];
    30: op1_09_in25 = reg_0391;
    31: op1_09_in25 = reg_0149;
    32: op1_09_in25 = reg_0722;
    33: op1_09_in25 = reg_0218;
    85: op1_09_in25 = reg_0218;
    34: op1_09_in25 = reg_0226;
    35: op1_09_in25 = reg_0271;
    36: op1_09_in25 = imem06_in[87:84];
    37: op1_09_in25 = reg_0788;
    38: op1_09_in25 = reg_0177;
    39: op1_09_in25 = imem01_in[91:88];
    40: op1_09_in25 = imem01_in[15:12];
    41: op1_09_in25 = reg_0086;
    42: op1_09_in25 = reg_0613;
    44: op1_09_in25 = reg_0588;
    45: op1_09_in25 = imem04_in[47:44];
    47: op1_09_in25 = reg_0750;
    48: op1_09_in25 = imem04_in[111:108];
    49: op1_09_in25 = reg_0362;
    50: op1_09_in25 = imem01_in[95:92];
    52: op1_09_in25 = reg_0646;
    53: op1_09_in25 = reg_0190;
    54: op1_09_in25 = reg_0811;
    55: op1_09_in25 = imem04_in[15:12];
    56: op1_09_in25 = reg_0555;
    57: op1_09_in25 = reg_0259;
    58: op1_09_in25 = reg_0132;
    59: op1_09_in25 = imem06_in[103:100];
    62: op1_09_in25 = reg_0530;
    63: op1_09_in25 = reg_0599;
    64: op1_09_in25 = reg_0560;
    65: op1_09_in25 = reg_0311;
    66: op1_09_in25 = reg_0429;
    67: op1_09_in25 = reg_0067;
    68: op1_09_in25 = imem01_in[115:112];
    69: op1_09_in25 = reg_0793;
    70: op1_09_in25 = imem06_in[51:48];
    71: op1_09_in25 = imem03_in[59:56];
    72: op1_09_in25 = imem06_in[3:0];
    73: op1_09_in25 = reg_0109;
    74: op1_09_in25 = reg_0714;
    76: op1_09_in25 = reg_0105;
    77: op1_09_in25 = reg_0290;
    78: op1_09_in25 = reg_0756;
    79: op1_09_in25 = reg_0245;
    80: op1_09_in25 = reg_0659;
    81: op1_09_in25 = imem05_in[47:44];
    82: op1_09_in25 = reg_0323;
    84: op1_09_in25 = reg_0640;
    86: op1_09_in25 = reg_0418;
    87: op1_09_in25 = imem04_in[79:76];
    88: op1_09_in25 = reg_0216;
    89: op1_09_in25 = imem04_in[83:80];
    90: op1_09_in25 = imem04_in[83:80];
    91: op1_09_in25 = imem06_in[23:20];
    93: op1_09_in25 = reg_0116;
    94: op1_09_in25 = reg_0099;
    95: op1_09_in25 = reg_0241;
    96: op1_09_in25 = reg_0726;
    default: op1_09_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv25 = 1;
    7: op1_09_inv25 = 1;
    9: op1_09_inv25 = 1;
    10: op1_09_inv25 = 1;
    15: op1_09_inv25 = 1;
    16: op1_09_inv25 = 1;
    19: op1_09_inv25 = 1;
    20: op1_09_inv25 = 1;
    26: op1_09_inv25 = 1;
    27: op1_09_inv25 = 1;
    28: op1_09_inv25 = 1;
    29: op1_09_inv25 = 1;
    32: op1_09_inv25 = 1;
    35: op1_09_inv25 = 1;
    36: op1_09_inv25 = 1;
    38: op1_09_inv25 = 1;
    39: op1_09_inv25 = 1;
    40: op1_09_inv25 = 1;
    41: op1_09_inv25 = 1;
    45: op1_09_inv25 = 1;
    56: op1_09_inv25 = 1;
    58: op1_09_inv25 = 1;
    60: op1_09_inv25 = 1;
    64: op1_09_inv25 = 1;
    65: op1_09_inv25 = 1;
    68: op1_09_inv25 = 1;
    69: op1_09_inv25 = 1;
    76: op1_09_inv25 = 1;
    78: op1_09_inv25 = 1;
    80: op1_09_inv25 = 1;
    82: op1_09_inv25 = 1;
    84: op1_09_inv25 = 1;
    85: op1_09_inv25 = 1;
    89: op1_09_inv25 = 1;
    90: op1_09_inv25 = 1;
    91: op1_09_inv25 = 1;
    93: op1_09_inv25 = 1;
    94: op1_09_inv25 = 1;
    96: op1_09_inv25 = 1;
    default: op1_09_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の26番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in26 = imem07_in[15:12];
    6: op1_09_in26 = reg_0107;
    7: op1_09_in26 = reg_0076;
    8: op1_09_in26 = reg_0178;
    9: op1_09_in26 = imem06_in[99:96];
    10: op1_09_in26 = reg_0109;
    11: op1_09_in26 = reg_0610;
    12: op1_09_in26 = imem03_in[59:56];
    13: op1_09_in26 = reg_0531;
    14: op1_09_in26 = imem06_in[3:0];
    15: op1_09_in26 = reg_0820;
    16: op1_09_in26 = reg_0572;
    17: op1_09_in26 = reg_0515;
    18: op1_09_in26 = reg_0342;
    19: op1_09_in26 = reg_0518;
    20: op1_09_in26 = imem04_in[103:100];
    23: op1_09_in26 = reg_0162;
    24: op1_09_in26 = reg_0241;
    25: op1_09_in26 = reg_0086;
    26: op1_09_in26 = reg_0640;
    27: op1_09_in26 = reg_0377;
    28: op1_09_in26 = imem01_in[35:32];
    29: op1_09_in26 = reg_0759;
    30: op1_09_in26 = reg_0398;
    31: op1_09_in26 = reg_0133;
    32: op1_09_in26 = reg_0710;
    33: op1_09_in26 = reg_0240;
    34: op1_09_in26 = reg_0224;
    35: op1_09_in26 = reg_0742;
    36: op1_09_in26 = imem06_in[107:104];
    59: op1_09_in26 = imem06_in[107:104];
    37: op1_09_in26 = reg_0783;
    38: op1_09_in26 = reg_0158;
    39: op1_09_in26 = imem01_in[95:92];
    40: op1_09_in26 = imem01_in[107:104];
    50: op1_09_in26 = imem01_in[107:104];
    41: op1_09_in26 = reg_0132;
    42: op1_09_in26 = reg_0817;
    44: op1_09_in26 = reg_0575;
    45: op1_09_in26 = imem04_in[51:48];
    47: op1_09_in26 = reg_0589;
    48: op1_09_in26 = imem05_in[19:16];
    49: op1_09_in26 = reg_0364;
    52: op1_09_in26 = reg_0497;
    53: op1_09_in26 = imem01_in[11:8];
    54: op1_09_in26 = reg_0008;
    55: op1_09_in26 = imem04_in[27:24];
    56: op1_09_in26 = reg_0060;
    57: op1_09_in26 = reg_0490;
    58: op1_09_in26 = reg_0135;
    60: op1_09_in26 = imem07_in[51:48];
    62: op1_09_in26 = reg_0756;
    63: op1_09_in26 = reg_0604;
    64: op1_09_in26 = reg_0553;
    65: op1_09_in26 = reg_0771;
    66: op1_09_in26 = reg_0079;
    67: op1_09_in26 = reg_0438;
    68: op1_09_in26 = reg_0423;
    69: op1_09_in26 = reg_0227;
    70: op1_09_in26 = imem06_in[95:92];
    71: op1_09_in26 = imem03_in[75:72];
    72: op1_09_in26 = imem06_in[47:44];
    73: op1_09_in26 = reg_0136;
    74: op1_09_in26 = imem07_in[11:8];
    76: op1_09_in26 = reg_0073;
    77: op1_09_in26 = reg_0248;
    78: op1_09_in26 = imem03_in[11:8];
    79: op1_09_in26 = reg_0328;
    80: op1_09_in26 = reg_0593;
    81: op1_09_in26 = imem05_in[107:104];
    82: op1_09_in26 = reg_0092;
    84: op1_09_in26 = reg_0776;
    85: op1_09_in26 = reg_0752;
    86: op1_09_in26 = reg_0306;
    87: op1_09_in26 = imem04_in[95:92];
    88: op1_09_in26 = reg_0425;
    89: op1_09_in26 = reg_0545;
    90: op1_09_in26 = imem04_in[107:104];
    91: op1_09_in26 = imem06_in[43:40];
    93: op1_09_in26 = reg_0099;
    94: op1_09_in26 = reg_0141;
    95: op1_09_in26 = reg_0258;
    96: op1_09_in26 = reg_0789;
    default: op1_09_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv26 = 1;
    7: op1_09_inv26 = 1;
    10: op1_09_inv26 = 1;
    12: op1_09_inv26 = 1;
    13: op1_09_inv26 = 1;
    14: op1_09_inv26 = 1;
    17: op1_09_inv26 = 1;
    19: op1_09_inv26 = 1;
    23: op1_09_inv26 = 1;
    24: op1_09_inv26 = 1;
    25: op1_09_inv26 = 1;
    29: op1_09_inv26 = 1;
    30: op1_09_inv26 = 1;
    33: op1_09_inv26 = 1;
    36: op1_09_inv26 = 1;
    39: op1_09_inv26 = 1;
    41: op1_09_inv26 = 1;
    42: op1_09_inv26 = 1;
    44: op1_09_inv26 = 1;
    45: op1_09_inv26 = 1;
    47: op1_09_inv26 = 1;
    48: op1_09_inv26 = 1;
    49: op1_09_inv26 = 1;
    53: op1_09_inv26 = 1;
    56: op1_09_inv26 = 1;
    59: op1_09_inv26 = 1;
    60: op1_09_inv26 = 1;
    64: op1_09_inv26 = 1;
    70: op1_09_inv26 = 1;
    71: op1_09_inv26 = 1;
    72: op1_09_inv26 = 1;
    73: op1_09_inv26 = 1;
    74: op1_09_inv26 = 1;
    78: op1_09_inv26 = 1;
    79: op1_09_inv26 = 1;
    82: op1_09_inv26 = 1;
    87: op1_09_inv26 = 1;
    91: op1_09_inv26 = 1;
    94: op1_09_inv26 = 1;
    95: op1_09_inv26 = 1;
    96: op1_09_inv26 = 1;
    default: op1_09_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の27番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in27 = imem07_in[51:48];
    74: op1_09_in27 = imem07_in[51:48];
    6: op1_09_in27 = imem02_in[31:28];
    7: op1_09_in27 = reg_0048;
    8: op1_09_in27 = reg_0157;
    9: op1_09_in27 = reg_0625;
    10: op1_09_in27 = reg_0107;
    11: op1_09_in27 = reg_0626;
    12: op1_09_in27 = imem03_in[67:64];
    13: op1_09_in27 = reg_0541;
    82: op1_09_in27 = reg_0541;
    14: op1_09_in27 = imem06_in[39:36];
    15: op1_09_in27 = reg_0825;
    16: op1_09_in27 = reg_0576;
    17: op1_09_in27 = reg_0225;
    18: op1_09_in27 = reg_0314;
    19: op1_09_in27 = reg_0525;
    20: op1_09_in27 = reg_0543;
    23: op1_09_in27 = reg_0166;
    24: op1_09_in27 = reg_0233;
    25: op1_09_in27 = reg_0089;
    26: op1_09_in27 = reg_0362;
    27: op1_09_in27 = reg_0589;
    28: op1_09_in27 = imem01_in[39:36];
    29: op1_09_in27 = reg_0771;
    30: op1_09_in27 = reg_0570;
    31: op1_09_in27 = reg_0151;
    32: op1_09_in27 = reg_0717;
    33: op1_09_in27 = reg_0234;
    34: op1_09_in27 = reg_0734;
    35: op1_09_in27 = reg_0733;
    36: op1_09_in27 = imem07_in[19:16];
    37: op1_09_in27 = reg_0090;
    65: op1_09_in27 = reg_0090;
    39: op1_09_in27 = imem01_in[103:100];
    40: op1_09_in27 = imem01_in[111:108];
    41: op1_09_in27 = reg_0145;
    42: op1_09_in27 = reg_0286;
    44: op1_09_in27 = reg_0568;
    45: op1_09_in27 = imem04_in[111:108];
    47: op1_09_in27 = reg_0597;
    48: op1_09_in27 = imem05_in[35:32];
    49: op1_09_in27 = reg_0348;
    50: op1_09_in27 = reg_0646;
    52: op1_09_in27 = reg_0653;
    53: op1_09_in27 = imem01_in[31:28];
    54: op1_09_in27 = reg_0806;
    55: op1_09_in27 = reg_0262;
    56: op1_09_in27 = reg_0057;
    57: op1_09_in27 = reg_0793;
    58: op1_09_in27 = reg_0133;
    59: op1_09_in27 = imem06_in[111:108];
    60: op1_09_in27 = imem07_in[63:60];
    62: op1_09_in27 = reg_0098;
    63: op1_09_in27 = reg_0319;
    64: op1_09_in27 = reg_0537;
    66: op1_09_in27 = reg_0430;
    67: op1_09_in27 = reg_0176;
    68: op1_09_in27 = reg_0217;
    69: op1_09_in27 = reg_0322;
    70: op1_09_in27 = imem06_in[99:96];
    71: op1_09_in27 = imem03_in[79:76];
    72: op1_09_in27 = imem06_in[71:68];
    91: op1_09_in27 = imem06_in[71:68];
    73: op1_09_in27 = reg_0735;
    79: op1_09_in27 = reg_0735;
    76: op1_09_in27 = reg_0104;
    77: op1_09_in27 = reg_0505;
    78: op1_09_in27 = imem03_in[15:12];
    80: op1_09_in27 = reg_0764;
    81: op1_09_in27 = reg_0792;
    84: op1_09_in27 = imem05_in[39:36];
    85: op1_09_in27 = imem07_in[43:40];
    86: op1_09_in27 = reg_0216;
    87: op1_09_in27 = imem04_in[127:124];
    88: op1_09_in27 = reg_0506;
    89: op1_09_in27 = reg_0171;
    90: op1_09_in27 = reg_0545;
    93: op1_09_in27 = reg_0141;
    94: op1_09_in27 = reg_0325;
    95: op1_09_in27 = reg_0741;
    96: op1_09_in27 = reg_0715;
    default: op1_09_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_09_inv27 = 1;
    9: op1_09_inv27 = 1;
    11: op1_09_inv27 = 1;
    12: op1_09_inv27 = 1;
    13: op1_09_inv27 = 1;
    14: op1_09_inv27 = 1;
    15: op1_09_inv27 = 1;
    16: op1_09_inv27 = 1;
    18: op1_09_inv27 = 1;
    23: op1_09_inv27 = 1;
    24: op1_09_inv27 = 1;
    25: op1_09_inv27 = 1;
    26: op1_09_inv27 = 1;
    30: op1_09_inv27 = 1;
    32: op1_09_inv27 = 1;
    34: op1_09_inv27 = 1;
    35: op1_09_inv27 = 1;
    37: op1_09_inv27 = 1;
    41: op1_09_inv27 = 1;
    42: op1_09_inv27 = 1;
    44: op1_09_inv27 = 1;
    45: op1_09_inv27 = 1;
    49: op1_09_inv27 = 1;
    50: op1_09_inv27 = 1;
    53: op1_09_inv27 = 1;
    54: op1_09_inv27 = 1;
    60: op1_09_inv27 = 1;
    62: op1_09_inv27 = 1;
    66: op1_09_inv27 = 1;
    69: op1_09_inv27 = 1;
    76: op1_09_inv27 = 1;
    77: op1_09_inv27 = 1;
    78: op1_09_inv27 = 1;
    79: op1_09_inv27 = 1;
    81: op1_09_inv27 = 1;
    82: op1_09_inv27 = 1;
    84: op1_09_inv27 = 1;
    89: op1_09_inv27 = 1;
    90: op1_09_inv27 = 1;
    91: op1_09_inv27 = 1;
    93: op1_09_inv27 = 1;
    94: op1_09_inv27 = 1;
    default: op1_09_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の28番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in28 = imem07_in[115:112];
    6: op1_09_in28 = imem02_in[123:120];
    7: op1_09_in28 = imem05_in[7:4];
    9: op1_09_in28 = reg_0607;
    10: op1_09_in28 = reg_0117;
    11: op1_09_in28 = reg_0608;
    12: op1_09_in28 = reg_0596;
    13: op1_09_in28 = reg_0547;
    14: op1_09_in28 = imem06_in[43:40];
    15: op1_09_in28 = reg_0232;
    16: op1_09_in28 = reg_0394;
    17: op1_09_in28 = reg_0247;
    87: op1_09_in28 = reg_0247;
    18: op1_09_in28 = reg_0092;
    19: op1_09_in28 = reg_0241;
    20: op1_09_in28 = reg_0557;
    23: op1_09_in28 = reg_0176;
    93: op1_09_in28 = reg_0176;
    24: op1_09_in28 = reg_0217;
    25: op1_09_in28 = reg_0147;
    26: op1_09_in28 = reg_0320;
    27: op1_09_in28 = reg_0585;
    28: op1_09_in28 = imem01_in[51:48];
    29: op1_09_in28 = reg_0550;
    30: op1_09_in28 = reg_0811;
    31: op1_09_in28 = reg_0134;
    32: op1_09_in28 = reg_0708;
    33: op1_09_in28 = reg_0104;
    34: op1_09_in28 = reg_0086;
    35: op1_09_in28 = reg_0086;
    36: op1_09_in28 = imem07_in[31:28];
    37: op1_09_in28 = reg_0735;
    50: op1_09_in28 = reg_0735;
    39: op1_09_in28 = imem01_in[111:108];
    40: op1_09_in28 = imem01_in[115:112];
    41: op1_09_in28 = reg_0133;
    42: op1_09_in28 = reg_0339;
    44: op1_09_in28 = reg_0517;
    45: op1_09_in28 = imem05_in[3:0];
    47: op1_09_in28 = reg_0588;
    48: op1_09_in28 = imem05_in[39:36];
    49: op1_09_in28 = reg_0530;
    52: op1_09_in28 = reg_0645;
    53: op1_09_in28 = imem01_in[79:76];
    54: op1_09_in28 = imem04_in[35:32];
    55: op1_09_in28 = reg_0043;
    56: op1_09_in28 = reg_0500;
    57: op1_09_in28 = reg_0782;
    58: op1_09_in28 = reg_0151;
    59: op1_09_in28 = imem06_in[119:116];
    60: op1_09_in28 = imem07_in[95:92];
    62: op1_09_in28 = reg_0498;
    63: op1_09_in28 = reg_0116;
    64: op1_09_in28 = reg_0055;
    65: op1_09_in28 = reg_0224;
    66: op1_09_in28 = reg_0503;
    68: op1_09_in28 = reg_0567;
    69: op1_09_in28 = reg_0245;
    70: op1_09_in28 = imem07_in[15:12];
    71: op1_09_in28 = imem03_in[119:116];
    72: op1_09_in28 = imem06_in[95:92];
    73: op1_09_in28 = reg_0282;
    74: op1_09_in28 = imem07_in[59:56];
    76: op1_09_in28 = reg_0660;
    77: op1_09_in28 = reg_0123;
    78: op1_09_in28 = imem03_in[31:28];
    79: op1_09_in28 = reg_0393;
    80: op1_09_in28 = reg_0515;
    81: op1_09_in28 = reg_0128;
    82: op1_09_in28 = reg_0081;
    84: op1_09_in28 = imem05_in[63:60];
    85: op1_09_in28 = imem07_in[91:88];
    86: op1_09_in28 = reg_0118;
    88: op1_09_in28 = reg_0673;
    89: op1_09_in28 = reg_0553;
    90: op1_09_in28 = reg_0537;
    91: op1_09_in28 = imem06_in[111:108];
    94: op1_09_in28 = reg_0279;
    95: op1_09_in28 = reg_0165;
    96: op1_09_in28 = reg_0635;
    default: op1_09_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_09_inv28 = 1;
    10: op1_09_inv28 = 1;
    11: op1_09_inv28 = 1;
    14: op1_09_inv28 = 1;
    18: op1_09_inv28 = 1;
    19: op1_09_inv28 = 1;
    20: op1_09_inv28 = 1;
    23: op1_09_inv28 = 1;
    25: op1_09_inv28 = 1;
    26: op1_09_inv28 = 1;
    28: op1_09_inv28 = 1;
    34: op1_09_inv28 = 1;
    35: op1_09_inv28 = 1;
    37: op1_09_inv28 = 1;
    39: op1_09_inv28 = 1;
    40: op1_09_inv28 = 1;
    44: op1_09_inv28 = 1;
    47: op1_09_inv28 = 1;
    49: op1_09_inv28 = 1;
    54: op1_09_inv28 = 1;
    55: op1_09_inv28 = 1;
    58: op1_09_inv28 = 1;
    60: op1_09_inv28 = 1;
    62: op1_09_inv28 = 1;
    63: op1_09_inv28 = 1;
    65: op1_09_inv28 = 1;
    66: op1_09_inv28 = 1;
    69: op1_09_inv28 = 1;
    74: op1_09_inv28 = 1;
    76: op1_09_inv28 = 1;
    78: op1_09_inv28 = 1;
    81: op1_09_inv28 = 1;
    82: op1_09_inv28 = 1;
    85: op1_09_inv28 = 1;
    86: op1_09_inv28 = 1;
    87: op1_09_inv28 = 1;
    91: op1_09_inv28 = 1;
    93: op1_09_inv28 = 1;
    94: op1_09_inv28 = 1;
    default: op1_09_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の29番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in29 = reg_0728;
    6: op1_09_in29 = reg_0642;
    7: op1_09_in29 = imem05_in[39:36];
    9: op1_09_in29 = reg_0631;
    10: op1_09_in29 = imem02_in[3:0];
    11: op1_09_in29 = reg_0349;
    12: op1_09_in29 = reg_0587;
    13: op1_09_in29 = reg_0301;
    14: op1_09_in29 = imem06_in[47:44];
    15: op1_09_in29 = reg_0235;
    16: op1_09_in29 = reg_0373;
    17: op1_09_in29 = reg_0503;
    18: op1_09_in29 = reg_0085;
    19: op1_09_in29 = reg_0233;
    20: op1_09_in29 = reg_0552;
    24: op1_09_in29 = reg_0245;
    25: op1_09_in29 = reg_0145;
    26: op1_09_in29 = reg_0229;
    27: op1_09_in29 = reg_0588;
    63: op1_09_in29 = reg_0588;
    28: op1_09_in29 = imem01_in[67:64];
    29: op1_09_in29 = reg_0760;
    30: op1_09_in29 = reg_0808;
    31: op1_09_in29 = reg_0032;
    32: op1_09_in29 = reg_0713;
    33: op1_09_in29 = reg_0108;
    34: op1_09_in29 = reg_0132;
    35: op1_09_in29 = reg_0132;
    36: op1_09_in29 = imem07_in[63:60];
    37: op1_09_in29 = reg_0282;
    39: op1_09_in29 = imem01_in[119:116];
    40: op1_09_in29 = reg_0111;
    41: op1_09_in29 = reg_0129;
    42: op1_09_in29 = reg_0370;
    44: op1_09_in29 = reg_0571;
    45: op1_09_in29 = imem05_in[7:4];
    47: op1_09_in29 = reg_0755;
    48: op1_09_in29 = imem05_in[43:40];
    49: op1_09_in29 = reg_0097;
    50: op1_09_in29 = reg_0653;
    52: op1_09_in29 = reg_0322;
    53: op1_09_in29 = imem01_in[99:96];
    54: op1_09_in29 = imem04_in[63:60];
    55: op1_09_in29 = reg_0308;
    56: op1_09_in29 = reg_0052;
    57: op1_09_in29 = reg_0309;
    58: op1_09_in29 = reg_0152;
    59: op1_09_in29 = reg_0348;
    60: op1_09_in29 = imem07_in[115:112];
    62: op1_09_in29 = reg_0740;
    64: op1_09_in29 = reg_0523;
    65: op1_09_in29 = reg_0225;
    66: op1_09_in29 = reg_0627;
    68: op1_09_in29 = reg_0506;
    69: op1_09_in29 = reg_0128;
    70: op1_09_in29 = imem07_in[31:28];
    71: op1_09_in29 = reg_0319;
    72: op1_09_in29 = imem06_in[119:116];
    91: op1_09_in29 = imem06_in[119:116];
    73: op1_09_in29 = reg_0393;
    74: op1_09_in29 = imem07_in[75:72];
    76: op1_09_in29 = reg_0677;
    77: op1_09_in29 = reg_0677;
    88: op1_09_in29 = reg_0677;
    78: op1_09_in29 = imem03_in[39:36];
    79: op1_09_in29 = reg_0277;
    80: op1_09_in29 = reg_0620;
    81: op1_09_in29 = reg_0146;
    82: op1_09_in29 = reg_0095;
    84: op1_09_in29 = imem05_in[83:80];
    85: op1_09_in29 = imem07_in[95:92];
    86: op1_09_in29 = reg_0104;
    87: op1_09_in29 = reg_0177;
    89: op1_09_in29 = reg_0275;
    90: op1_09_in29 = reg_0060;
    95: op1_09_in29 = reg_0107;
    96: op1_09_in29 = reg_0442;
    default: op1_09_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv29 = 1;
    6: op1_09_inv29 = 1;
    7: op1_09_inv29 = 1;
    9: op1_09_inv29 = 1;
    11: op1_09_inv29 = 1;
    12: op1_09_inv29 = 1;
    13: op1_09_inv29 = 1;
    14: op1_09_inv29 = 1;
    17: op1_09_inv29 = 1;
    18: op1_09_inv29 = 1;
    19: op1_09_inv29 = 1;
    20: op1_09_inv29 = 1;
    25: op1_09_inv29 = 1;
    27: op1_09_inv29 = 1;
    29: op1_09_inv29 = 1;
    30: op1_09_inv29 = 1;
    31: op1_09_inv29 = 1;
    32: op1_09_inv29 = 1;
    33: op1_09_inv29 = 1;
    34: op1_09_inv29 = 1;
    39: op1_09_inv29 = 1;
    40: op1_09_inv29 = 1;
    41: op1_09_inv29 = 1;
    42: op1_09_inv29 = 1;
    45: op1_09_inv29 = 1;
    50: op1_09_inv29 = 1;
    52: op1_09_inv29 = 1;
    56: op1_09_inv29 = 1;
    62: op1_09_inv29 = 1;
    70: op1_09_inv29 = 1;
    73: op1_09_inv29 = 1;
    80: op1_09_inv29 = 1;
    81: op1_09_inv29 = 1;
    82: op1_09_inv29 = 1;
    84: op1_09_inv29 = 1;
    85: op1_09_inv29 = 1;
    86: op1_09_inv29 = 1;
    87: op1_09_inv29 = 1;
    88: op1_09_inv29 = 1;
    90: op1_09_inv29 = 1;
    default: op1_09_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の30番目の入力
  always @ ( * ) begin
    case ( state )
    5: op1_09_in30 = reg_0702;
    6: op1_09_in30 = reg_0646;
    7: op1_09_in30 = imem05_in[79:76];
    9: op1_09_in30 = reg_0626;
    10: op1_09_in30 = imem02_in[31:28];
    11: op1_09_in30 = reg_0404;
    12: op1_09_in30 = reg_0592;
    13: op1_09_in30 = reg_0306;
    14: op1_09_in30 = reg_0259;
    15: op1_09_in30 = reg_0505;
    16: op1_09_in30 = reg_0322;
    17: op1_09_in30 = reg_0236;
    18: op1_09_in30 = imem03_in[59:56];
    19: op1_09_in30 = reg_0215;
    20: op1_09_in30 = reg_0555;
    24: op1_09_in30 = reg_0238;
    25: op1_09_in30 = reg_0128;
    26: op1_09_in30 = reg_0324;
    27: op1_09_in30 = imem03_in[3:0];
    28: op1_09_in30 = imem01_in[79:76];
    29: op1_09_in30 = reg_0559;
    30: op1_09_in30 = reg_0803;
    31: op1_09_in30 = reg_0753;
    32: op1_09_in30 = reg_0701;
    33: op1_09_in30 = reg_0114;
    34: op1_09_in30 = reg_0135;
    35: op1_09_in30 = reg_0135;
    36: op1_09_in30 = imem07_in[75:72];
    37: op1_09_in30 = reg_0272;
    39: op1_09_in30 = reg_0123;
    40: op1_09_in30 = reg_0100;
    52: op1_09_in30 = reg_0100;
    41: op1_09_in30 = reg_0140;
    42: op1_09_in30 = reg_0748;
    44: op1_09_in30 = reg_0562;
    45: op1_09_in30 = imem05_in[123:120];
    47: op1_09_in30 = reg_0373;
    48: op1_09_in30 = imem05_in[91:88];
    49: op1_09_in30 = reg_0769;
    50: op1_09_in30 = reg_0663;
    53: op1_09_in30 = imem01_in[123:120];
    54: op1_09_in30 = imem04_in[103:100];
    55: op1_09_in30 = reg_0432;
    56: op1_09_in30 = reg_0076;
    57: op1_09_in30 = reg_0742;
    58: op1_09_in30 = reg_0154;
    59: op1_09_in30 = reg_0625;
    60: op1_09_in30 = reg_0722;
    62: op1_09_in30 = reg_0532;
    63: op1_09_in30 = reg_0388;
    64: op1_09_in30 = reg_0058;
    65: op1_09_in30 = reg_0490;
    66: op1_09_in30 = reg_0614;
    68: op1_09_in30 = reg_0424;
    69: op1_09_in30 = reg_0066;
    70: op1_09_in30 = imem07_in[59:56];
    71: op1_09_in30 = reg_0329;
    72: op1_09_in30 = reg_0817;
    73: op1_09_in30 = reg_0784;
    74: op1_09_in30 = imem07_in[83:80];
    76: op1_09_in30 = reg_0675;
    77: op1_09_in30 = reg_0675;
    78: op1_09_in30 = imem03_in[47:44];
    79: op1_09_in30 = reg_0827;
    80: op1_09_in30 = reg_0651;
    81: op1_09_in30 = reg_0782;
    82: op1_09_in30 = reg_0540;
    84: op1_09_in30 = imem05_in[87:84];
    85: op1_09_in30 = reg_0163;
    86: op1_09_in30 = reg_0119;
    87: op1_09_in30 = reg_0611;
    88: op1_09_in30 = reg_0671;
    89: op1_09_in30 = reg_0249;
    90: op1_09_in30 = reg_0551;
    91: op1_09_in30 = reg_0619;
    95: op1_09_in30 = reg_0234;
    96: op1_09_in30 = reg_0438;
    default: op1_09_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_09_inv30 = 1;
    6: op1_09_inv30 = 1;
    9: op1_09_inv30 = 1;
    10: op1_09_inv30 = 1;
    13: op1_09_inv30 = 1;
    16: op1_09_inv30 = 1;
    24: op1_09_inv30 = 1;
    25: op1_09_inv30 = 1;
    26: op1_09_inv30 = 1;
    27: op1_09_inv30 = 1;
    28: op1_09_inv30 = 1;
    30: op1_09_inv30 = 1;
    31: op1_09_inv30 = 1;
    33: op1_09_inv30 = 1;
    36: op1_09_inv30 = 1;
    37: op1_09_inv30 = 1;
    39: op1_09_inv30 = 1;
    41: op1_09_inv30 = 1;
    45: op1_09_inv30 = 1;
    48: op1_09_inv30 = 1;
    52: op1_09_inv30 = 1;
    62: op1_09_inv30 = 1;
    63: op1_09_inv30 = 1;
    64: op1_09_inv30 = 1;
    68: op1_09_inv30 = 1;
    79: op1_09_inv30 = 1;
    80: op1_09_inv30 = 1;
    82: op1_09_inv30 = 1;
    95: op1_09_inv30 = 1;
    96: op1_09_inv30 = 1;
    default: op1_09_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_09_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_09_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in00 = imem00_in[103:100];
    5: op1_10_in00 = imem00_in[31:28];
    92: op1_10_in00 = imem00_in[31:28];
    6: op1_10_in00 = reg_0664;
    80: op1_10_in00 = reg_0664;
    7: op1_10_in00 = imem05_in[107:104];
    8: op1_10_in00 = imem00_in[47:44];
    9: op1_10_in00 = reg_0601;
    76: op1_10_in00 = reg_0601;
    10: op1_10_in00 = imem02_in[83:80];
    11: op1_10_in00 = reg_0367;
    12: op1_10_in00 = reg_0589;
    13: op1_10_in00 = reg_0302;
    56: op1_10_in00 = reg_0302;
    14: op1_10_in00 = imem06_in[59:56];
    15: op1_10_in00 = reg_0218;
    16: op1_10_in00 = reg_0331;
    3: op1_10_in00 = imem07_in[31:28];
    17: op1_10_in00 = reg_0249;
    18: op1_10_in00 = imem03_in[79:76];
    19: op1_10_in00 = reg_0220;
    20: op1_10_in00 = reg_0551;
    21: op1_10_in00 = reg_0685;
    22: op1_10_in00 = imem00_in[59:56];
    23: op1_10_in00 = imem00_in[3:0];
    46: op1_10_in00 = imem00_in[3:0];
    24: op1_10_in00 = reg_0105;
    2: op1_10_in00 = imem07_in[107:104];
    70: op1_10_in00 = imem07_in[107:104];
    25: op1_10_in00 = reg_0156;
    26: op1_10_in00 = reg_0518;
    27: op1_10_in00 = imem03_in[27:24];
    28: op1_10_in00 = imem01_in[95:92];
    29: op1_10_in00 = reg_0505;
    30: op1_10_in00 = reg_0806;
    1: op1_10_in00 = imem07_in[67:64];
    31: op1_10_in00 = reg_0037;
    32: op1_10_in00 = reg_0706;
    33: op1_10_in00 = reg_0100;
    34: op1_10_in00 = reg_0150;
    35: op1_10_in00 = reg_0154;
    36: op1_10_in00 = imem07_in[79:76];
    37: op1_10_in00 = reg_0732;
    81: op1_10_in00 = reg_0732;
    38: op1_10_in00 = imem00_in[15:12];
    67: op1_10_in00 = imem00_in[15:12];
    75: op1_10_in00 = imem00_in[15:12];
    93: op1_10_in00 = imem00_in[15:12];
    39: op1_10_in00 = reg_0111;
    40: op1_10_in00 = reg_0106;
    41: op1_10_in00 = reg_0131;
    42: op1_10_in00 = reg_0270;
    43: op1_10_in00 = imem00_in[19:16];
    44: op1_10_in00 = reg_0376;
    45: op1_10_in00 = reg_0482;
    47: op1_10_in00 = reg_0392;
    48: op1_10_in00 = reg_0791;
    49: op1_10_in00 = reg_0770;
    50: op1_10_in00 = reg_0557;
    51: op1_10_in00 = imem00_in[7:4];
    83: op1_10_in00 = imem00_in[7:4];
    52: op1_10_in00 = reg_0563;
    53: op1_10_in00 = reg_0322;
    54: op1_10_in00 = imem04_in[111:108];
    55: op1_10_in00 = reg_0430;
    57: op1_10_in00 = reg_0229;
    58: op1_10_in00 = reg_0129;
    59: op1_10_in00 = reg_0346;
    60: op1_10_in00 = reg_0704;
    61: op1_10_in00 = imem00_in[67:64];
    62: op1_10_in00 = imem03_in[11:8];
    63: op1_10_in00 = reg_0385;
    64: op1_10_in00 = reg_0510;
    65: op1_10_in00 = reg_0085;
    66: op1_10_in00 = reg_0065;
    68: op1_10_in00 = reg_0219;
    69: op1_10_in00 = reg_0086;
    71: op1_10_in00 = reg_0399;
    72: op1_10_in00 = reg_0298;
    73: op1_10_in00 = reg_0389;
    74: op1_10_in00 = imem07_in[87:84];
    77: op1_10_in00 = reg_0674;
    78: op1_10_in00 = imem03_in[71:68];
    79: op1_10_in00 = reg_0785;
    82: op1_10_in00 = imem03_in[7:4];
    84: op1_10_in00 = imem05_in[111:108];
    85: op1_10_in00 = reg_0103;
    86: op1_10_in00 = reg_0660;
    87: op1_10_in00 = reg_0508;
    88: op1_10_in00 = imem02_in[39:36];
    89: op1_10_in00 = reg_0556;
    90: op1_10_in00 = reg_0556;
    91: op1_10_in00 = reg_0260;
    94: op1_10_in00 = imem00_in[71:68];
    95: op1_10_in00 = imem01_in[11:8];
    96: op1_10_in00 = reg_0448;
    default: op1_10_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv00 = 1;
    5: op1_10_inv00 = 1;
    10: op1_10_inv00 = 1;
    12: op1_10_inv00 = 1;
    13: op1_10_inv00 = 1;
    14: op1_10_inv00 = 1;
    16: op1_10_inv00 = 1;
    17: op1_10_inv00 = 1;
    18: op1_10_inv00 = 1;
    19: op1_10_inv00 = 1;
    20: op1_10_inv00 = 1;
    21: op1_10_inv00 = 1;
    23: op1_10_inv00 = 1;
    2: op1_10_inv00 = 1;
    26: op1_10_inv00 = 1;
    27: op1_10_inv00 = 1;
    28: op1_10_inv00 = 1;
    1: op1_10_inv00 = 1;
    32: op1_10_inv00 = 1;
    35: op1_10_inv00 = 1;
    36: op1_10_inv00 = 1;
    37: op1_10_inv00 = 1;
    40: op1_10_inv00 = 1;
    42: op1_10_inv00 = 1;
    44: op1_10_inv00 = 1;
    45: op1_10_inv00 = 1;
    46: op1_10_inv00 = 1;
    51: op1_10_inv00 = 1;
    56: op1_10_inv00 = 1;
    57: op1_10_inv00 = 1;
    59: op1_10_inv00 = 1;
    61: op1_10_inv00 = 1;
    62: op1_10_inv00 = 1;
    66: op1_10_inv00 = 1;
    68: op1_10_inv00 = 1;
    69: op1_10_inv00 = 1;
    70: op1_10_inv00 = 1;
    71: op1_10_inv00 = 1;
    75: op1_10_inv00 = 1;
    77: op1_10_inv00 = 1;
    82: op1_10_inv00 = 1;
    86: op1_10_inv00 = 1;
    87: op1_10_inv00 = 1;
    88: op1_10_inv00 = 1;
    89: op1_10_inv00 = 1;
    92: op1_10_inv00 = 1;
    93: op1_10_inv00 = 1;
    default: op1_10_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in01 = imem00_in[115:112];
    5: op1_10_in01 = imem00_in[35:32];
    6: op1_10_in01 = reg_0663;
    7: op1_10_in01 = reg_0796;
    8: op1_10_in01 = imem00_in[51:48];
    43: op1_10_in01 = imem00_in[51:48];
    9: op1_10_in01 = reg_0356;
    10: op1_10_in01 = reg_0650;
    11: op1_10_in01 = reg_0034;
    12: op1_10_in01 = reg_0580;
    13: op1_10_in01 = reg_0293;
    14: op1_10_in01 = reg_0614;
    15: op1_10_in01 = reg_0239;
    16: op1_10_in01 = reg_0002;
    3: op1_10_in01 = imem07_in[39:36];
    17: op1_10_in01 = reg_0118;
    18: op1_10_in01 = imem03_in[91:88];
    19: op1_10_in01 = reg_0111;
    20: op1_10_in01 = reg_0308;
    21: op1_10_in01 = reg_0686;
    22: op1_10_in01 = imem00_in[103:100];
    23: op1_10_in01 = imem00_in[11:8];
    83: op1_10_in01 = imem00_in[11:8];
    24: op1_10_in01 = reg_0122;
    2: op1_10_in01 = imem07_in[111:108];
    74: op1_10_in01 = imem07_in[111:108];
    25: op1_10_in01 = reg_0154;
    26: op1_10_in01 = reg_0540;
    27: op1_10_in01 = imem03_in[31:28];
    82: op1_10_in01 = imem03_in[31:28];
    28: op1_10_in01 = reg_0772;
    29: op1_10_in01 = reg_0511;
    30: op1_10_in01 = reg_0810;
    1: op1_10_in01 = imem07_in[103:100];
    31: op1_10_in01 = reg_0752;
    32: op1_10_in01 = reg_0436;
    33: op1_10_in01 = reg_0127;
    34: op1_10_in01 = reg_0156;
    35: op1_10_in01 = reg_0129;
    36: op1_10_in01 = imem07_in[91:88];
    37: op1_10_in01 = reg_0128;
    38: op1_10_in01 = imem00_in[47:44];
    39: op1_10_in01 = reg_0116;
    40: op1_10_in01 = reg_0115;
    41: op1_10_in01 = imem06_in[11:8];
    42: op1_10_in01 = reg_0764;
    44: op1_10_in01 = reg_0396;
    45: op1_10_in01 = reg_0797;
    46: op1_10_in01 = imem00_in[31:28];
    47: op1_10_in01 = reg_0570;
    48: op1_10_in01 = reg_0792;
    49: op1_10_in01 = reg_0539;
    50: op1_10_in01 = reg_0294;
    51: op1_10_in01 = imem00_in[15:12];
    52: op1_10_in01 = reg_0759;
    53: op1_10_in01 = reg_0550;
    54: op1_10_in01 = reg_0083;
    55: op1_10_in01 = reg_0508;
    56: op1_10_in01 = reg_0629;
    57: op1_10_in01 = reg_0224;
    58: op1_10_in01 = imem06_in[35:32];
    59: op1_10_in01 = reg_0409;
    60: op1_10_in01 = reg_0712;
    61: op1_10_in01 = imem00_in[83:80];
    62: op1_10_in01 = imem03_in[63:60];
    63: op1_10_in01 = reg_0572;
    64: op1_10_in01 = reg_0305;
    65: op1_10_in01 = reg_0039;
    66: op1_10_in01 = reg_0513;
    67: op1_10_in01 = imem00_in[59:56];
    68: op1_10_in01 = reg_0124;
    69: op1_10_in01 = reg_0136;
    70: op1_10_in01 = reg_0719;
    71: op1_10_in01 = reg_0568;
    72: op1_10_in01 = reg_0354;
    73: op1_10_in01 = reg_0736;
    75: op1_10_in01 = imem00_in[23:20];
    76: op1_10_in01 = reg_0674;
    77: op1_10_in01 = imem02_in[15:12];
    78: op1_10_in01 = imem03_in[107:104];
    79: op1_10_in01 = reg_0830;
    80: op1_10_in01 = reg_0652;
    81: op1_10_in01 = reg_0665;
    84: op1_10_in01 = reg_0791;
    85: op1_10_in01 = reg_0442;
    86: op1_10_in01 = imem02_in[35:32];
    87: op1_10_in01 = reg_0223;
    88: op1_10_in01 = imem02_in[47:44];
    89: op1_10_in01 = reg_0079;
    90: op1_10_in01 = reg_0174;
    91: op1_10_in01 = reg_0402;
    92: op1_10_in01 = imem00_in[55:52];
    93: op1_10_in01 = imem00_in[19:16];
    94: op1_10_in01 = reg_0698;
    95: op1_10_in01 = imem01_in[27:24];
    96: op1_10_in01 = reg_0180;
    default: op1_10_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv01 = 1;
    6: op1_10_inv01 = 1;
    7: op1_10_inv01 = 1;
    9: op1_10_inv01 = 1;
    15: op1_10_inv01 = 1;
    16: op1_10_inv01 = 1;
    17: op1_10_inv01 = 1;
    19: op1_10_inv01 = 1;
    20: op1_10_inv01 = 1;
    21: op1_10_inv01 = 1;
    23: op1_10_inv01 = 1;
    2: op1_10_inv01 = 1;
    25: op1_10_inv01 = 1;
    27: op1_10_inv01 = 1;
    28: op1_10_inv01 = 1;
    29: op1_10_inv01 = 1;
    30: op1_10_inv01 = 1;
    33: op1_10_inv01 = 1;
    34: op1_10_inv01 = 1;
    36: op1_10_inv01 = 1;
    37: op1_10_inv01 = 1;
    40: op1_10_inv01 = 1;
    41: op1_10_inv01 = 1;
    42: op1_10_inv01 = 1;
    47: op1_10_inv01 = 1;
    48: op1_10_inv01 = 1;
    51: op1_10_inv01 = 1;
    52: op1_10_inv01 = 1;
    53: op1_10_inv01 = 1;
    55: op1_10_inv01 = 1;
    57: op1_10_inv01 = 1;
    58: op1_10_inv01 = 1;
    61: op1_10_inv01 = 1;
    62: op1_10_inv01 = 1;
    63: op1_10_inv01 = 1;
    64: op1_10_inv01 = 1;
    65: op1_10_inv01 = 1;
    67: op1_10_inv01 = 1;
    70: op1_10_inv01 = 1;
    73: op1_10_inv01 = 1;
    74: op1_10_inv01 = 1;
    75: op1_10_inv01 = 1;
    76: op1_10_inv01 = 1;
    77: op1_10_inv01 = 1;
    80: op1_10_inv01 = 1;
    86: op1_10_inv01 = 1;
    91: op1_10_inv01 = 1;
    92: op1_10_inv01 = 1;
    96: op1_10_inv01 = 1;
    default: op1_10_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in02 = reg_0685;
    5: op1_10_in02 = imem00_in[47:44];
    6: op1_10_in02 = reg_0358;
    7: op1_10_in02 = reg_0483;
    8: op1_10_in02 = imem00_in[71:68];
    9: op1_10_in02 = reg_0344;
    10: op1_10_in02 = reg_0647;
    11: op1_10_in02 = reg_0815;
    12: op1_10_in02 = reg_0588;
    13: op1_10_in02 = reg_0048;
    14: op1_10_in02 = reg_0625;
    15: op1_10_in02 = reg_0217;
    53: op1_10_in02 = reg_0217;
    16: op1_10_in02 = reg_0015;
    3: op1_10_in02 = imem07_in[71:68];
    17: op1_10_in02 = reg_0116;
    18: op1_10_in02 = imem03_in[107:104];
    62: op1_10_in02 = imem03_in[107:104];
    19: op1_10_in02 = reg_0125;
    20: op1_10_in02 = reg_0534;
    21: op1_10_in02 = reg_0679;
    22: op1_10_in02 = reg_0679;
    23: op1_10_in02 = imem00_in[35:32];
    24: op1_10_in02 = reg_0104;
    2: op1_10_in02 = reg_0175;
    25: op1_10_in02 = imem06_in[115:112];
    26: op1_10_in02 = reg_0535;
    27: op1_10_in02 = imem03_in[79:76];
    28: op1_10_in02 = reg_0514;
    29: op1_10_in02 = reg_0242;
    30: op1_10_in02 = reg_0809;
    1: op1_10_in02 = imem07_in[111:108];
    31: op1_10_in02 = reg_0614;
    32: op1_10_in02 = reg_0434;
    33: op1_10_in02 = imem02_in[7:4];
    76: op1_10_in02 = imem02_in[7:4];
    34: op1_10_in02 = reg_0130;
    35: op1_10_in02 = reg_0141;
    36: op1_10_in02 = imem07_in[119:116];
    37: op1_10_in02 = reg_0154;
    69: op1_10_in02 = reg_0154;
    38: op1_10_in02 = imem00_in[59:56];
    39: op1_10_in02 = reg_0108;
    40: op1_10_in02 = reg_0126;
    41: op1_10_in02 = imem06_in[31:28];
    42: op1_10_in02 = reg_0778;
    43: op1_10_in02 = imem00_in[83:80];
    44: op1_10_in02 = reg_0001;
    45: op1_10_in02 = reg_0491;
    46: op1_10_in02 = imem00_in[39:36];
    75: op1_10_in02 = imem00_in[39:36];
    47: op1_10_in02 = reg_0019;
    48: op1_10_in02 = reg_0493;
    49: op1_10_in02 = reg_0756;
    50: op1_10_in02 = reg_0506;
    51: op1_10_in02 = imem00_in[51:48];
    52: op1_10_in02 = reg_0422;
    54: op1_10_in02 = reg_0523;
    55: op1_10_in02 = reg_0050;
    56: op1_10_in02 = reg_0078;
    57: op1_10_in02 = reg_0258;
    65: op1_10_in02 = reg_0258;
    58: op1_10_in02 = imem06_in[111:108];
    59: op1_10_in02 = reg_0298;
    60: op1_10_in02 = reg_0709;
    61: op1_10_in02 = imem00_in[115:112];
    92: op1_10_in02 = imem00_in[115:112];
    63: op1_10_in02 = reg_0374;
    64: op1_10_in02 = reg_0077;
    66: op1_10_in02 = reg_0109;
    67: op1_10_in02 = imem00_in[67:64];
    68: op1_10_in02 = reg_0073;
    70: op1_10_in02 = reg_0721;
    71: op1_10_in02 = reg_0623;
    72: op1_10_in02 = reg_0618;
    73: op1_10_in02 = reg_0227;
    84: op1_10_in02 = reg_0227;
    74: op1_10_in02 = reg_0064;
    77: op1_10_in02 = imem02_in[31:28];
    78: op1_10_in02 = imem03_in[115:112];
    79: op1_10_in02 = imem06_in[19:16];
    80: op1_10_in02 = reg_0767;
    81: op1_10_in02 = reg_0134;
    82: op1_10_in02 = imem03_in[39:36];
    83: op1_10_in02 = imem00_in[27:24];
    85: op1_10_in02 = reg_0279;
    86: op1_10_in02 = imem02_in[43:40];
    87: op1_10_in02 = imem05_in[47:44];
    88: op1_10_in02 = imem02_in[59:56];
    89: op1_10_in02 = reg_0433;
    90: op1_10_in02 = reg_0432;
    91: op1_10_in02 = reg_0039;
    93: op1_10_in02 = imem00_in[79:76];
    94: op1_10_in02 = reg_0690;
    95: op1_10_in02 = imem01_in[31:28];
    96: op1_10_in02 = reg_0236;
    default: op1_10_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv02 = 1;
    8: op1_10_inv02 = 1;
    10: op1_10_inv02 = 1;
    11: op1_10_inv02 = 1;
    13: op1_10_inv02 = 1;
    15: op1_10_inv02 = 1;
    3: op1_10_inv02 = 1;
    19: op1_10_inv02 = 1;
    20: op1_10_inv02 = 1;
    21: op1_10_inv02 = 1;
    22: op1_10_inv02 = 1;
    23: op1_10_inv02 = 1;
    2: op1_10_inv02 = 1;
    27: op1_10_inv02 = 1;
    28: op1_10_inv02 = 1;
    29: op1_10_inv02 = 1;
    30: op1_10_inv02 = 1;
    32: op1_10_inv02 = 1;
    33: op1_10_inv02 = 1;
    36: op1_10_inv02 = 1;
    38: op1_10_inv02 = 1;
    39: op1_10_inv02 = 1;
    41: op1_10_inv02 = 1;
    42: op1_10_inv02 = 1;
    44: op1_10_inv02 = 1;
    45: op1_10_inv02 = 1;
    46: op1_10_inv02 = 1;
    54: op1_10_inv02 = 1;
    55: op1_10_inv02 = 1;
    56: op1_10_inv02 = 1;
    57: op1_10_inv02 = 1;
    59: op1_10_inv02 = 1;
    61: op1_10_inv02 = 1;
    62: op1_10_inv02 = 1;
    63: op1_10_inv02 = 1;
    65: op1_10_inv02 = 1;
    67: op1_10_inv02 = 1;
    69: op1_10_inv02 = 1;
    70: op1_10_inv02 = 1;
    72: op1_10_inv02 = 1;
    73: op1_10_inv02 = 1;
    77: op1_10_inv02 = 1;
    79: op1_10_inv02 = 1;
    82: op1_10_inv02 = 1;
    83: op1_10_inv02 = 1;
    84: op1_10_inv02 = 1;
    85: op1_10_inv02 = 1;
    86: op1_10_inv02 = 1;
    87: op1_10_inv02 = 1;
    88: op1_10_inv02 = 1;
    90: op1_10_inv02 = 1;
    91: op1_10_inv02 = 1;
    92: op1_10_inv02 = 1;
    93: op1_10_inv02 = 1;
    95: op1_10_inv02 = 1;
    default: op1_10_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in03 = reg_0689;
    5: op1_10_in03 = imem00_in[51:48];
    46: op1_10_in03 = imem00_in[51:48];
    6: op1_10_in03 = reg_0325;
    7: op1_10_in03 = reg_0489;
    8: op1_10_in03 = imem00_in[75:72];
    9: op1_10_in03 = reg_0381;
    10: op1_10_in03 = reg_0648;
    11: op1_10_in03 = reg_0037;
    12: op1_10_in03 = reg_0590;
    13: op1_10_in03 = imem05_in[11:8];
    14: op1_10_in03 = reg_0630;
    15: op1_10_in03 = reg_0238;
    16: op1_10_in03 = reg_0810;
    3: op1_10_in03 = imem07_in[75:72];
    17: op1_10_in03 = reg_0119;
    18: op1_10_in03 = reg_0569;
    19: op1_10_in03 = reg_0106;
    20: op1_10_in03 = reg_0529;
    21: op1_10_in03 = reg_0691;
    22: op1_10_in03 = reg_0690;
    23: op1_10_in03 = imem00_in[43:40];
    24: op1_10_in03 = reg_0120;
    2: op1_10_in03 = reg_0181;
    25: op1_10_in03 = reg_0614;
    26: op1_10_in03 = imem03_in[47:44];
    27: op1_10_in03 = imem03_in[111:108];
    28: op1_10_in03 = reg_0824;
    29: op1_10_in03 = reg_0240;
    30: op1_10_in03 = imem04_in[15:12];
    31: op1_10_in03 = reg_0607;
    32: op1_10_in03 = reg_0446;
    33: op1_10_in03 = imem02_in[27:24];
    34: op1_10_in03 = imem06_in[11:8];
    35: op1_10_in03 = reg_0137;
    36: op1_10_in03 = reg_0713;
    37: op1_10_in03 = reg_0134;
    38: op1_10_in03 = imem00_in[83:80];
    39: op1_10_in03 = reg_0100;
    40: op1_10_in03 = imem02_in[7:4];
    41: op1_10_in03 = reg_0299;
    42: op1_10_in03 = reg_0375;
    43: op1_10_in03 = imem00_in[103:100];
    44: op1_10_in03 = reg_0800;
    45: op1_10_in03 = reg_0492;
    47: op1_10_in03 = reg_0803;
    48: op1_10_in03 = reg_0793;
    49: op1_10_in03 = reg_0526;
    50: op1_10_in03 = reg_0219;
    51: op1_10_in03 = reg_0695;
    52: op1_10_in03 = reg_0574;
    53: op1_10_in03 = reg_0567;
    54: op1_10_in03 = reg_0058;
    55: op1_10_in03 = reg_0520;
    56: op1_10_in03 = reg_0075;
    57: op1_10_in03 = reg_0249;
    58: op1_10_in03 = reg_0289;
    59: op1_10_in03 = reg_0293;
    60: op1_10_in03 = reg_0718;
    61: op1_10_in03 = imem00_in[119:116];
    62: op1_10_in03 = reg_0597;
    63: op1_10_in03 = reg_0389;
    64: op1_10_in03 = reg_0074;
    65: op1_10_in03 = reg_0277;
    66: op1_10_in03 = imem05_in[31:28];
    67: op1_10_in03 = imem00_in[95:92];
    93: op1_10_in03 = imem00_in[95:92];
    68: op1_10_in03 = reg_0125;
    69: op1_10_in03 = imem06_in[47:44];
    70: op1_10_in03 = reg_0723;
    71: op1_10_in03 = reg_0570;
    72: op1_10_in03 = reg_0260;
    73: op1_10_in03 = reg_0666;
    74: op1_10_in03 = reg_0266;
    75: op1_10_in03 = reg_0696;
    76: op1_10_in03 = imem02_in[15:12];
    77: op1_10_in03 = imem02_in[35:32];
    78: op1_10_in03 = reg_0347;
    79: op1_10_in03 = imem06_in[39:36];
    80: op1_10_in03 = reg_0256;
    81: op1_10_in03 = reg_0328;
    82: op1_10_in03 = imem03_in[75:72];
    83: op1_10_in03 = imem00_in[35:32];
    84: op1_10_in03 = reg_0499;
    86: op1_10_in03 = imem02_in[75:72];
    87: op1_10_in03 = imem05_in[51:48];
    88: op1_10_in03 = imem02_in[71:68];
    89: op1_10_in03 = reg_0076;
    90: op1_10_in03 = reg_0430;
    91: op1_10_in03 = reg_0519;
    92: op1_10_in03 = reg_0683;
    94: op1_10_in03 = reg_0758;
    95: op1_10_in03 = imem01_in[35:32];
    96: op1_10_in03 = reg_0426;
    default: op1_10_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv03 = 1;
    8: op1_10_inv03 = 1;
    9: op1_10_inv03 = 1;
    11: op1_10_inv03 = 1;
    14: op1_10_inv03 = 1;
    16: op1_10_inv03 = 1;
    3: op1_10_inv03 = 1;
    17: op1_10_inv03 = 1;
    18: op1_10_inv03 = 1;
    19: op1_10_inv03 = 1;
    21: op1_10_inv03 = 1;
    23: op1_10_inv03 = 1;
    24: op1_10_inv03 = 1;
    25: op1_10_inv03 = 1;
    26: op1_10_inv03 = 1;
    28: op1_10_inv03 = 1;
    31: op1_10_inv03 = 1;
    36: op1_10_inv03 = 1;
    38: op1_10_inv03 = 1;
    39: op1_10_inv03 = 1;
    40: op1_10_inv03 = 1;
    43: op1_10_inv03 = 1;
    45: op1_10_inv03 = 1;
    47: op1_10_inv03 = 1;
    48: op1_10_inv03 = 1;
    50: op1_10_inv03 = 1;
    52: op1_10_inv03 = 1;
    54: op1_10_inv03 = 1;
    56: op1_10_inv03 = 1;
    65: op1_10_inv03 = 1;
    66: op1_10_inv03 = 1;
    67: op1_10_inv03 = 1;
    70: op1_10_inv03 = 1;
    71: op1_10_inv03 = 1;
    72: op1_10_inv03 = 1;
    73: op1_10_inv03 = 1;
    74: op1_10_inv03 = 1;
    75: op1_10_inv03 = 1;
    76: op1_10_inv03 = 1;
    77: op1_10_inv03 = 1;
    78: op1_10_inv03 = 1;
    79: op1_10_inv03 = 1;
    80: op1_10_inv03 = 1;
    81: op1_10_inv03 = 1;
    86: op1_10_inv03 = 1;
    89: op1_10_inv03 = 1;
    91: op1_10_inv03 = 1;
    95: op1_10_inv03 = 1;
    96: op1_10_inv03 = 1;
    default: op1_10_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in04 = reg_0679;
    5: op1_10_in04 = imem00_in[99:96];
    6: op1_10_in04 = reg_0341;
    7: op1_10_in04 = reg_0486;
    8: op1_10_in04 = imem00_in[123:120];
    9: op1_10_in04 = reg_0372;
    10: op1_10_in04 = reg_0665;
    11: op1_10_in04 = reg_0030;
    12: op1_10_in04 = reg_0391;
    13: op1_10_in04 = imem05_in[15:12];
    14: op1_10_in04 = reg_0618;
    15: op1_10_in04 = reg_0122;
    16: op1_10_in04 = reg_0004;
    3: op1_10_in04 = imem07_in[111:108];
    17: op1_10_in04 = reg_0114;
    18: op1_10_in04 = reg_0369;
    19: op1_10_in04 = reg_0109;
    20: op1_10_in04 = reg_0267;
    21: op1_10_in04 = reg_0680;
    22: op1_10_in04 = reg_0677;
    23: op1_10_in04 = imem00_in[47:44];
    83: op1_10_in04 = imem00_in[47:44];
    24: op1_10_in04 = reg_0106;
    39: op1_10_in04 = reg_0106;
    2: op1_10_in04 = reg_0162;
    25: op1_10_in04 = reg_0625;
    58: op1_10_in04 = reg_0625;
    26: op1_10_in04 = imem03_in[103:100];
    27: op1_10_in04 = imem03_in[123:120];
    28: op1_10_in04 = reg_0227;
    29: op1_10_in04 = reg_0216;
    30: op1_10_in04 = imem04_in[23:20];
    31: op1_10_in04 = reg_0620;
    32: op1_10_in04 = reg_0449;
    33: op1_10_in04 = imem02_in[63:60];
    34: op1_10_in04 = imem06_in[15:12];
    35: op1_10_in04 = reg_0144;
    37: op1_10_in04 = reg_0144;
    36: op1_10_in04 = reg_0711;
    38: op1_10_in04 = imem00_in[87:84];
    40: op1_10_in04 = imem02_in[11:8];
    41: op1_10_in04 = reg_0624;
    42: op1_10_in04 = reg_0818;
    43: op1_10_in04 = imem00_in[127:124];
    44: op1_10_in04 = imem04_in[39:36];
    45: op1_10_in04 = reg_0793;
    46: op1_10_in04 = imem00_in[75:72];
    47: op1_10_in04 = imem04_in[15:12];
    48: op1_10_in04 = reg_0785;
    49: op1_10_in04 = imem03_in[43:40];
    50: op1_10_in04 = reg_0113;
    51: op1_10_in04 = reg_0681;
    52: op1_10_in04 = reg_0244;
    53: op1_10_in04 = reg_0244;
    54: op1_10_in04 = reg_0500;
    55: op1_10_in04 = reg_0078;
    56: op1_10_in04 = reg_0507;
    57: op1_10_in04 = reg_0257;
    59: op1_10_in04 = reg_0260;
    60: op1_10_in04 = reg_0441;
    61: op1_10_in04 = reg_0693;
    62: op1_10_in04 = reg_0493;
    63: op1_10_in04 = reg_0803;
    64: op1_10_in04 = reg_0617;
    65: op1_10_in04 = imem05_in[23:20];
    66: op1_10_in04 = imem05_in[51:48];
    67: op1_10_in04 = reg_0697;
    68: op1_10_in04 = reg_0592;
    69: op1_10_in04 = imem06_in[95:92];
    70: op1_10_in04 = reg_0715;
    71: op1_10_in04 = reg_0019;
    72: op1_10_in04 = reg_0578;
    73: op1_10_in04 = reg_0070;
    74: op1_10_in04 = reg_0061;
    75: op1_10_in04 = reg_0698;
    76: op1_10_in04 = imem02_in[19:16];
    77: op1_10_in04 = imem02_in[87:84];
    78: op1_10_in04 = reg_0028;
    79: op1_10_in04 = imem06_in[51:48];
    80: op1_10_in04 = reg_0175;
    81: op1_10_in04 = reg_0389;
    82: op1_10_in04 = imem03_in[91:88];
    84: op1_10_in04 = reg_0134;
    86: op1_10_in04 = imem02_in[83:80];
    88: op1_10_in04 = imem02_in[83:80];
    87: op1_10_in04 = imem05_in[67:64];
    89: op1_10_in04 = reg_0529;
    90: op1_10_in04 = reg_0503;
    91: op1_10_in04 = reg_0307;
    92: op1_10_in04 = reg_0689;
    93: op1_10_in04 = reg_0000;
    94: op1_10_in04 = reg_0130;
    95: op1_10_in04 = imem01_in[63:60];
    96: op1_10_in04 = reg_0182;
    default: op1_10_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv04 = 1;
    7: op1_10_inv04 = 1;
    8: op1_10_inv04 = 1;
    10: op1_10_inv04 = 1;
    15: op1_10_inv04 = 1;
    16: op1_10_inv04 = 1;
    19: op1_10_inv04 = 1;
    21: op1_10_inv04 = 1;
    22: op1_10_inv04 = 1;
    27: op1_10_inv04 = 1;
    28: op1_10_inv04 = 1;
    29: op1_10_inv04 = 1;
    30: op1_10_inv04 = 1;
    32: op1_10_inv04 = 1;
    35: op1_10_inv04 = 1;
    36: op1_10_inv04 = 1;
    37: op1_10_inv04 = 1;
    40: op1_10_inv04 = 1;
    41: op1_10_inv04 = 1;
    42: op1_10_inv04 = 1;
    43: op1_10_inv04 = 1;
    44: op1_10_inv04 = 1;
    45: op1_10_inv04 = 1;
    49: op1_10_inv04 = 1;
    51: op1_10_inv04 = 1;
    52: op1_10_inv04 = 1;
    54: op1_10_inv04 = 1;
    56: op1_10_inv04 = 1;
    58: op1_10_inv04 = 1;
    59: op1_10_inv04 = 1;
    61: op1_10_inv04 = 1;
    63: op1_10_inv04 = 1;
    67: op1_10_inv04 = 1;
    70: op1_10_inv04 = 1;
    71: op1_10_inv04 = 1;
    72: op1_10_inv04 = 1;
    74: op1_10_inv04 = 1;
    75: op1_10_inv04 = 1;
    76: op1_10_inv04 = 1;
    78: op1_10_inv04 = 1;
    79: op1_10_inv04 = 1;
    80: op1_10_inv04 = 1;
    83: op1_10_inv04 = 1;
    84: op1_10_inv04 = 1;
    87: op1_10_inv04 = 1;
    88: op1_10_inv04 = 1;
    89: op1_10_inv04 = 1;
    90: op1_10_inv04 = 1;
    92: op1_10_inv04 = 1;
    93: op1_10_inv04 = 1;
    95: op1_10_inv04 = 1;
    96: op1_10_inv04 = 1;
    default: op1_10_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in05 = reg_0690;
    51: op1_10_in05 = reg_0690;
    5: op1_10_in05 = reg_0693;
    6: op1_10_in05 = reg_0346;
    7: op1_10_in05 = reg_0256;
    8: op1_10_in05 = reg_0688;
    9: op1_10_in05 = reg_0408;
    10: op1_10_in05 = reg_0341;
    11: op1_10_in05 = imem07_in[15:12];
    12: op1_10_in05 = reg_0360;
    13: op1_10_in05 = imem05_in[51:48];
    14: op1_10_in05 = reg_0632;
    15: op1_10_in05 = reg_0124;
    16: op1_10_in05 = imem04_in[115:112];
    3: op1_10_in05 = imem07_in[119:116];
    17: op1_10_in05 = reg_0106;
    18: op1_10_in05 = reg_0396;
    19: op1_10_in05 = reg_0107;
    24: op1_10_in05 = reg_0107;
    20: op1_10_in05 = reg_0268;
    21: op1_10_in05 = reg_0687;
    22: op1_10_in05 = reg_0675;
    23: op1_10_in05 = imem00_in[71:68];
    2: op1_10_in05 = reg_0183;
    25: op1_10_in05 = reg_0613;
    72: op1_10_in05 = reg_0613;
    26: op1_10_in05 = imem03_in[107:104];
    82: op1_10_in05 = imem03_in[107:104];
    27: op1_10_in05 = reg_0803;
    28: op1_10_in05 = reg_0519;
    29: op1_10_in05 = reg_0245;
    30: op1_10_in05 = imem04_in[51:48];
    44: op1_10_in05 = imem04_in[51:48];
    31: op1_10_in05 = reg_0608;
    32: op1_10_in05 = reg_0442;
    33: op1_10_in05 = imem02_in[87:84];
    34: op1_10_in05 = imem06_in[19:16];
    35: op1_10_in05 = reg_0753;
    36: op1_10_in05 = reg_0707;
    37: op1_10_in05 = imem06_in[15:12];
    38: op1_10_in05 = reg_0695;
    46: op1_10_in05 = reg_0695;
    39: op1_10_in05 = reg_0115;
    40: op1_10_in05 = imem02_in[63:60];
    41: op1_10_in05 = reg_0298;
    42: op1_10_in05 = reg_0231;
    43: op1_10_in05 = reg_0682;
    45: op1_10_in05 = reg_0782;
    47: op1_10_in05 = imem04_in[31:28];
    48: op1_10_in05 = reg_0790;
    49: op1_10_in05 = imem03_in[87:84];
    50: op1_10_in05 = reg_0126;
    52: op1_10_in05 = imem01_in[15:12];
    53: op1_10_in05 = reg_0248;
    54: op1_10_in05 = reg_0077;
    55: op1_10_in05 = reg_0789;
    56: op1_10_in05 = reg_0515;
    57: op1_10_in05 = reg_0277;
    58: op1_10_in05 = reg_0609;
    59: op1_10_in05 = reg_0405;
    60: op1_10_in05 = reg_0253;
    61: op1_10_in05 = reg_0696;
    62: op1_10_in05 = reg_0573;
    63: op1_10_in05 = reg_0807;
    64: op1_10_in05 = reg_0065;
    65: op1_10_in05 = imem05_in[43:40];
    66: op1_10_in05 = imem05_in[59:56];
    67: op1_10_in05 = reg_0683;
    68: op1_10_in05 = reg_0119;
    69: op1_10_in05 = reg_0762;
    70: op1_10_in05 = reg_0718;
    71: op1_10_in05 = reg_0001;
    73: op1_10_in05 = reg_0027;
    74: op1_10_in05 = reg_0444;
    75: op1_10_in05 = reg_0684;
    76: op1_10_in05 = imem02_in[79:76];
    77: op1_10_in05 = imem02_in[103:100];
    86: op1_10_in05 = imem02_in[103:100];
    78: op1_10_in05 = reg_0575;
    79: op1_10_in05 = imem06_in[75:72];
    80: op1_10_in05 = reg_0179;
    81: op1_10_in05 = reg_0058;
    83: op1_10_in05 = imem00_in[55:52];
    84: op1_10_in05 = reg_0486;
    87: op1_10_in05 = imem05_in[99:96];
    88: op1_10_in05 = imem02_in[111:108];
    89: op1_10_in05 = reg_0430;
    90: op1_10_in05 = reg_0629;
    91: op1_10_in05 = reg_0748;
    92: op1_10_in05 = reg_0658;
    93: op1_10_in05 = reg_0691;
    94: op1_10_in05 = reg_0016;
    95: op1_10_in05 = imem01_in[67:64];
    96: op1_10_in05 = reg_0100;
    default: op1_10_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv05 = 1;
    8: op1_10_inv05 = 1;
    9: op1_10_inv05 = 1;
    13: op1_10_inv05 = 1;
    16: op1_10_inv05 = 1;
    18: op1_10_inv05 = 1;
    21: op1_10_inv05 = 1;
    22: op1_10_inv05 = 1;
    24: op1_10_inv05 = 1;
    25: op1_10_inv05 = 1;
    26: op1_10_inv05 = 1;
    27: op1_10_inv05 = 1;
    28: op1_10_inv05 = 1;
    29: op1_10_inv05 = 1;
    30: op1_10_inv05 = 1;
    31: op1_10_inv05 = 1;
    32: op1_10_inv05 = 1;
    33: op1_10_inv05 = 1;
    34: op1_10_inv05 = 1;
    36: op1_10_inv05 = 1;
    38: op1_10_inv05 = 1;
    40: op1_10_inv05 = 1;
    48: op1_10_inv05 = 1;
    49: op1_10_inv05 = 1;
    50: op1_10_inv05 = 1;
    52: op1_10_inv05 = 1;
    53: op1_10_inv05 = 1;
    54: op1_10_inv05 = 1;
    57: op1_10_inv05 = 1;
    61: op1_10_inv05 = 1;
    68: op1_10_inv05 = 1;
    69: op1_10_inv05 = 1;
    70: op1_10_inv05 = 1;
    72: op1_10_inv05 = 1;
    73: op1_10_inv05 = 1;
    75: op1_10_inv05 = 1;
    76: op1_10_inv05 = 1;
    77: op1_10_inv05 = 1;
    82: op1_10_inv05 = 1;
    89: op1_10_inv05 = 1;
    94: op1_10_inv05 = 1;
    95: op1_10_inv05 = 1;
    96: op1_10_inv05 = 1;
    default: op1_10_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in06 = reg_0691;
    51: op1_10_in06 = reg_0691;
    75: op1_10_in06 = reg_0691;
    92: op1_10_in06 = reg_0691;
    5: op1_10_in06 = reg_0694;
    6: op1_10_in06 = reg_0324;
    7: op1_10_in06 = reg_0252;
    8: op1_10_in06 = reg_0465;
    22: op1_10_in06 = reg_0465;
    9: op1_10_in06 = reg_0313;
    10: op1_10_in06 = reg_0353;
    11: op1_10_in06 = imem07_in[19:16];
    12: op1_10_in06 = reg_0317;
    13: op1_10_in06 = imem05_in[55:52];
    14: op1_10_in06 = reg_0623;
    15: op1_10_in06 = reg_0125;
    16: op1_10_in06 = imem04_in[119:116];
    3: op1_10_in06 = reg_0447;
    17: op1_10_in06 = reg_0110;
    18: op1_10_in06 = reg_0331;
    19: op1_10_in06 = reg_0127;
    20: op1_10_in06 = reg_0297;
    21: op1_10_in06 = reg_0699;
    23: op1_10_in06 = imem00_in[87:84];
    24: op1_10_in06 = imem02_in[19:16];
    2: op1_10_in06 = reg_0166;
    25: op1_10_in06 = reg_0606;
    26: op1_10_in06 = imem03_in[111:108];
    27: op1_10_in06 = reg_0807;
    28: op1_10_in06 = reg_0771;
    29: op1_10_in06 = reg_0119;
    30: op1_10_in06 = imem04_in[59:56];
    31: op1_10_in06 = reg_0622;
    32: op1_10_in06 = reg_0443;
    33: op1_10_in06 = imem02_in[103:100];
    34: op1_10_in06 = imem06_in[87:84];
    35: op1_10_in06 = reg_0812;
    81: op1_10_in06 = reg_0812;
    36: op1_10_in06 = reg_0701;
    37: op1_10_in06 = imem06_in[27:24];
    38: op1_10_in06 = reg_0670;
    39: op1_10_in06 = reg_0107;
    40: op1_10_in06 = imem02_in[107:104];
    86: op1_10_in06 = imem02_in[107:104];
    41: op1_10_in06 = reg_0265;
    42: op1_10_in06 = reg_0238;
    43: op1_10_in06 = reg_0457;
    44: op1_10_in06 = imem04_in[91:88];
    45: op1_10_in06 = reg_0737;
    46: op1_10_in06 = reg_0683;
    47: op1_10_in06 = imem04_in[63:60];
    48: op1_10_in06 = reg_0485;
    49: op1_10_in06 = imem03_in[95:92];
    50: op1_10_in06 = imem02_in[7:4];
    52: op1_10_in06 = imem01_in[27:24];
    53: op1_10_in06 = reg_0234;
    54: op1_10_in06 = reg_0071;
    55: op1_10_in06 = reg_0780;
    56: op1_10_in06 = reg_0227;
    57: op1_10_in06 = reg_0285;
    58: op1_10_in06 = reg_0618;
    59: op1_10_in06 = reg_0821;
    60: op1_10_in06 = reg_0266;
    61: op1_10_in06 = reg_0612;
    62: op1_10_in06 = reg_0755;
    63: op1_10_in06 = reg_0802;
    64: op1_10_in06 = reg_0259;
    65: op1_10_in06 = imem05_in[59:56];
    66: op1_10_in06 = reg_0791;
    67: op1_10_in06 = reg_0407;
    68: op1_10_in06 = reg_0120;
    69: op1_10_in06 = reg_0619;
    70: op1_10_in06 = reg_0334;
    71: op1_10_in06 = reg_0801;
    72: op1_10_in06 = reg_0377;
    73: op1_10_in06 = reg_0517;
    74: op1_10_in06 = reg_0438;
    76: op1_10_in06 = imem02_in[87:84];
    77: op1_10_in06 = reg_0142;
    78: op1_10_in06 = reg_0001;
    79: op1_10_in06 = reg_0348;
    80: op1_10_in06 = reg_0249;
    82: op1_10_in06 = reg_0602;
    83: op1_10_in06 = imem00_in[63:60];
    84: op1_10_in06 = reg_0328;
    87: op1_10_in06 = imem05_in[107:104];
    88: op1_10_in06 = reg_0533;
    89: op1_10_in06 = reg_0077;
    90: op1_10_in06 = reg_0508;
    91: op1_10_in06 = reg_0638;
    93: op1_10_in06 = reg_0688;
    94: op1_10_in06 = reg_0029;
    95: op1_10_in06 = imem01_in[91:88];
    96: op1_10_in06 = reg_0091;
    default: op1_10_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv06 = 1;
    8: op1_10_inv06 = 1;
    11: op1_10_inv06 = 1;
    12: op1_10_inv06 = 1;
    13: op1_10_inv06 = 1;
    15: op1_10_inv06 = 1;
    17: op1_10_inv06 = 1;
    20: op1_10_inv06 = 1;
    21: op1_10_inv06 = 1;
    23: op1_10_inv06 = 1;
    24: op1_10_inv06 = 1;
    25: op1_10_inv06 = 1;
    26: op1_10_inv06 = 1;
    28: op1_10_inv06 = 1;
    30: op1_10_inv06 = 1;
    31: op1_10_inv06 = 1;
    32: op1_10_inv06 = 1;
    33: op1_10_inv06 = 1;
    35: op1_10_inv06 = 1;
    36: op1_10_inv06 = 1;
    43: op1_10_inv06 = 1;
    44: op1_10_inv06 = 1;
    45: op1_10_inv06 = 1;
    47: op1_10_inv06 = 1;
    48: op1_10_inv06 = 1;
    49: op1_10_inv06 = 1;
    52: op1_10_inv06 = 1;
    55: op1_10_inv06 = 1;
    59: op1_10_inv06 = 1;
    60: op1_10_inv06 = 1;
    62: op1_10_inv06 = 1;
    63: op1_10_inv06 = 1;
    65: op1_10_inv06 = 1;
    66: op1_10_inv06 = 1;
    67: op1_10_inv06 = 1;
    68: op1_10_inv06 = 1;
    71: op1_10_inv06 = 1;
    72: op1_10_inv06 = 1;
    73: op1_10_inv06 = 1;
    74: op1_10_inv06 = 1;
    77: op1_10_inv06 = 1;
    79: op1_10_inv06 = 1;
    81: op1_10_inv06 = 1;
    82: op1_10_inv06 = 1;
    84: op1_10_inv06 = 1;
    88: op1_10_inv06 = 1;
    90: op1_10_inv06 = 1;
    91: op1_10_inv06 = 1;
    default: op1_10_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in07 = reg_0675;
    5: op1_10_in07 = reg_0676;
    6: op1_10_in07 = reg_0335;
    10: op1_10_in07 = reg_0335;
    7: op1_10_in07 = reg_0254;
    8: op1_10_in07 = reg_0453;
    21: op1_10_in07 = reg_0453;
    22: op1_10_in07 = reg_0453;
    9: op1_10_in07 = reg_0375;
    11: op1_10_in07 = imem07_in[31:28];
    12: op1_10_in07 = reg_0361;
    13: op1_10_in07 = imem05_in[59:56];
    14: op1_10_in07 = reg_0615;
    15: op1_10_in07 = reg_0114;
    16: op1_10_in07 = reg_0530;
    3: op1_10_in07 = reg_0419;
    17: op1_10_in07 = imem02_in[51:48];
    18: op1_10_in07 = reg_0013;
    19: op1_10_in07 = imem02_in[23:20];
    24: op1_10_in07 = imem02_in[23:20];
    20: op1_10_in07 = reg_0286;
    23: op1_10_in07 = imem00_in[103:100];
    25: op1_10_in07 = reg_0609;
    26: op1_10_in07 = imem03_in[123:120];
    27: op1_10_in07 = reg_0802;
    28: op1_10_in07 = reg_0515;
    29: op1_10_in07 = reg_0112;
    30: op1_10_in07 = imem04_in[75:72];
    31: op1_10_in07 = reg_0762;
    32: op1_10_in07 = reg_0169;
    33: op1_10_in07 = imem02_in[123:120];
    34: op1_10_in07 = reg_0625;
    35: op1_10_in07 = reg_0040;
    36: op1_10_in07 = reg_0425;
    37: op1_10_in07 = imem06_in[47:44];
    38: op1_10_in07 = reg_0687;
    39: op1_10_in07 = imem02_in[19:16];
    40: op1_10_in07 = imem02_in[127:124];
    41: op1_10_in07 = reg_0369;
    42: op1_10_in07 = reg_0632;
    43: op1_10_in07 = reg_0466;
    44: op1_10_in07 = reg_0542;
    45: op1_10_in07 = reg_0742;
    46: op1_10_in07 = reg_0696;
    47: op1_10_in07 = imem04_in[71:68];
    48: op1_10_in07 = reg_0279;
    49: op1_10_in07 = imem03_in[103:100];
    50: op1_10_in07 = imem02_in[99:96];
    51: op1_10_in07 = reg_0680;
    52: op1_10_in07 = imem01_in[83:80];
    53: op1_10_in07 = reg_0122;
    54: op1_10_in07 = reg_0431;
    55: op1_10_in07 = imem05_in[15:12];
    56: op1_10_in07 = reg_0519;
    57: op1_10_in07 = reg_0086;
    58: op1_10_in07 = reg_0593;
    59: op1_10_in07 = reg_0608;
    60: op1_10_in07 = reg_0439;
    61: op1_10_in07 = reg_0698;
    62: op1_10_in07 = reg_0568;
    63: op1_10_in07 = imem04_in[7:4];
    64: op1_10_in07 = reg_0090;
    65: op1_10_in07 = imem05_in[87:84];
    66: op1_10_in07 = reg_0792;
    67: op1_10_in07 = reg_0454;
    68: op1_10_in07 = reg_0106;
    69: op1_10_in07 = reg_0766;
    70: op1_10_in07 = reg_0441;
    71: op1_10_in07 = reg_0008;
    72: op1_10_in07 = reg_0405;
    73: op1_10_in07 = reg_0386;
    74: op1_10_in07 = reg_0435;
    75: op1_10_in07 = reg_0469;
    76: op1_10_in07 = imem02_in[119:116];
    77: op1_10_in07 = reg_0392;
    78: op1_10_in07 = reg_0806;
    79: op1_10_in07 = reg_0409;
    80: op1_10_in07 = reg_0100;
    81: op1_10_in07 = reg_0149;
    82: op1_10_in07 = reg_0317;
    83: op1_10_in07 = imem00_in[119:116];
    84: op1_10_in07 = reg_0500;
    86: op1_10_in07 = imem02_in[111:108];
    87: op1_10_in07 = imem05_in[123:120];
    88: op1_10_in07 = reg_0656;
    89: op1_10_in07 = reg_0629;
    90: op1_10_in07 = reg_0062;
    91: op1_10_in07 = reg_0328;
    92: op1_10_in07 = reg_0063;
    93: op1_10_in07 = reg_0029;
    94: op1_10_in07 = reg_0699;
    95: op1_10_in07 = imem01_in[95:92];
    default: op1_10_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv07 = 1;
    5: op1_10_inv07 = 1;
    9: op1_10_inv07 = 1;
    11: op1_10_inv07 = 1;
    12: op1_10_inv07 = 1;
    13: op1_10_inv07 = 1;
    15: op1_10_inv07 = 1;
    16: op1_10_inv07 = 1;
    3: op1_10_inv07 = 1;
    17: op1_10_inv07 = 1;
    19: op1_10_inv07 = 1;
    20: op1_10_inv07 = 1;
    25: op1_10_inv07 = 1;
    26: op1_10_inv07 = 1;
    29: op1_10_inv07 = 1;
    30: op1_10_inv07 = 1;
    31: op1_10_inv07 = 1;
    33: op1_10_inv07 = 1;
    35: op1_10_inv07 = 1;
    37: op1_10_inv07 = 1;
    39: op1_10_inv07 = 1;
    40: op1_10_inv07 = 1;
    44: op1_10_inv07 = 1;
    45: op1_10_inv07 = 1;
    47: op1_10_inv07 = 1;
    49: op1_10_inv07 = 1;
    50: op1_10_inv07 = 1;
    51: op1_10_inv07 = 1;
    52: op1_10_inv07 = 1;
    53: op1_10_inv07 = 1;
    54: op1_10_inv07 = 1;
    58: op1_10_inv07 = 1;
    59: op1_10_inv07 = 1;
    60: op1_10_inv07 = 1;
    61: op1_10_inv07 = 1;
    63: op1_10_inv07 = 1;
    67: op1_10_inv07 = 1;
    70: op1_10_inv07 = 1;
    73: op1_10_inv07 = 1;
    75: op1_10_inv07 = 1;
    76: op1_10_inv07 = 1;
    77: op1_10_inv07 = 1;
    79: op1_10_inv07 = 1;
    81: op1_10_inv07 = 1;
    83: op1_10_inv07 = 1;
    84: op1_10_inv07 = 1;
    87: op1_10_inv07 = 1;
    88: op1_10_inv07 = 1;
    89: op1_10_inv07 = 1;
    90: op1_10_inv07 = 1;
    91: op1_10_inv07 = 1;
    92: op1_10_inv07 = 1;
    default: op1_10_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in08 = reg_0680;
    5: op1_10_in08 = reg_0671;
    6: op1_10_in08 = reg_0347;
    7: op1_10_in08 = reg_0255;
    8: op1_10_in08 = reg_0460;
    9: op1_10_in08 = reg_0382;
    10: op1_10_in08 = reg_0328;
    11: op1_10_in08 = imem07_in[43:40];
    12: op1_10_in08 = reg_0396;
    13: op1_10_in08 = imem05_in[103:100];
    14: op1_10_in08 = reg_0405;
    15: op1_10_in08 = imem02_in[15:12];
    16: op1_10_in08 = reg_0534;
    3: op1_10_in08 = reg_0443;
    17: op1_10_in08 = imem02_in[71:68];
    18: op1_10_in08 = reg_0800;
    19: op1_10_in08 = imem02_in[47:44];
    20: op1_10_in08 = reg_0278;
    21: op1_10_in08 = reg_0454;
    22: op1_10_in08 = reg_0457;
    93: op1_10_in08 = reg_0457;
    23: op1_10_in08 = reg_0672;
    24: op1_10_in08 = imem02_in[115:112];
    25: op1_10_in08 = reg_0611;
    26: op1_10_in08 = reg_0572;
    27: op1_10_in08 = reg_0015;
    28: op1_10_in08 = reg_0232;
    29: op1_10_in08 = reg_0106;
    30: op1_10_in08 = reg_0316;
    31: op1_10_in08 = reg_0319;
    32: op1_10_in08 = reg_0177;
    33: op1_10_in08 = reg_0645;
    34: op1_10_in08 = reg_0629;
    35: op1_10_in08 = reg_0616;
    36: op1_10_in08 = reg_0433;
    37: op1_10_in08 = imem06_in[67:64];
    38: op1_10_in08 = reg_0450;
    67: op1_10_in08 = reg_0450;
    39: op1_10_in08 = imem02_in[51:48];
    40: op1_10_in08 = reg_0664;
    41: op1_10_in08 = reg_0762;
    42: op1_10_in08 = reg_0288;
    84: op1_10_in08 = reg_0288;
    43: op1_10_in08 = reg_0472;
    44: op1_10_in08 = reg_0060;
    45: op1_10_in08 = reg_0732;
    46: op1_10_in08 = reg_0676;
    47: op1_10_in08 = imem04_in[79:76];
    48: op1_10_in08 = reg_0269;
    49: op1_10_in08 = imem03_in[111:108];
    50: op1_10_in08 = reg_0642;
    51: op1_10_in08 = reg_0453;
    92: op1_10_in08 = reg_0453;
    52: op1_10_in08 = imem02_in[19:16];
    53: op1_10_in08 = reg_0670;
    54: op1_10_in08 = reg_0626;
    55: op1_10_in08 = imem05_in[31:28];
    56: op1_10_in08 = reg_0644;
    57: op1_10_in08 = reg_0089;
    58: op1_10_in08 = reg_0035;
    59: op1_10_in08 = reg_0764;
    60: op1_10_in08 = reg_0437;
    61: op1_10_in08 = reg_0684;
    62: op1_10_in08 = reg_0373;
    63: op1_10_in08 = imem04_in[11:8];
    64: op1_10_in08 = reg_0797;
    65: op1_10_in08 = reg_0132;
    66: op1_10_in08 = reg_0231;
    68: op1_10_in08 = reg_0601;
    69: op1_10_in08 = reg_0265;
    70: op1_10_in08 = reg_0636;
    71: op1_10_in08 = reg_0016;
    72: op1_10_in08 = reg_0515;
    73: op1_10_in08 = reg_0279;
    74: op1_10_in08 = reg_0174;
    75: op1_10_in08 = reg_0481;
    76: op1_10_in08 = imem02_in[123:120];
    86: op1_10_in08 = imem02_in[123:120];
    77: op1_10_in08 = reg_0426;
    78: op1_10_in08 = imem04_in[23:20];
    79: op1_10_in08 = reg_0609;
    80: op1_10_in08 = reg_0171;
    81: op1_10_in08 = reg_0827;
    82: op1_10_in08 = reg_0604;
    83: op1_10_in08 = reg_0682;
    87: op1_10_in08 = reg_0667;
    88: op1_10_in08 = reg_0647;
    89: op1_10_in08 = reg_0617;
    90: op1_10_in08 = reg_0065;
    91: op1_10_in08 = reg_0335;
    94: op1_10_in08 = reg_0464;
    95: op1_10_in08 = imem01_in[111:108];
    default: op1_10_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv08 = 1;
    8: op1_10_inv08 = 1;
    9: op1_10_inv08 = 1;
    11: op1_10_inv08 = 1;
    12: op1_10_inv08 = 1;
    13: op1_10_inv08 = 1;
    16: op1_10_inv08 = 1;
    3: op1_10_inv08 = 1;
    18: op1_10_inv08 = 1;
    21: op1_10_inv08 = 1;
    23: op1_10_inv08 = 1;
    29: op1_10_inv08 = 1;
    30: op1_10_inv08 = 1;
    31: op1_10_inv08 = 1;
    34: op1_10_inv08 = 1;
    36: op1_10_inv08 = 1;
    39: op1_10_inv08 = 1;
    41: op1_10_inv08 = 1;
    44: op1_10_inv08 = 1;
    47: op1_10_inv08 = 1;
    48: op1_10_inv08 = 1;
    49: op1_10_inv08 = 1;
    56: op1_10_inv08 = 1;
    58: op1_10_inv08 = 1;
    59: op1_10_inv08 = 1;
    60: op1_10_inv08 = 1;
    61: op1_10_inv08 = 1;
    63: op1_10_inv08 = 1;
    64: op1_10_inv08 = 1;
    69: op1_10_inv08 = 1;
    70: op1_10_inv08 = 1;
    72: op1_10_inv08 = 1;
    77: op1_10_inv08 = 1;
    78: op1_10_inv08 = 1;
    79: op1_10_inv08 = 1;
    81: op1_10_inv08 = 1;
    82: op1_10_inv08 = 1;
    84: op1_10_inv08 = 1;
    87: op1_10_inv08 = 1;
    88: op1_10_inv08 = 1;
    89: op1_10_inv08 = 1;
    92: op1_10_inv08 = 1;
    94: op1_10_inv08 = 1;
    default: op1_10_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in09 = reg_0451;
    5: op1_10_in09 = reg_0465;
    6: op1_10_in09 = imem03_in[35:32];
    7: op1_10_in09 = reg_0263;
    8: op1_10_in09 = reg_0480;
    9: op1_10_in09 = reg_0404;
    10: op1_10_in09 = reg_0097;
    11: op1_10_in09 = imem07_in[91:88];
    12: op1_10_in09 = reg_0000;
    13: op1_10_in09 = imem05_in[107:104];
    14: op1_10_in09 = reg_0029;
    15: op1_10_in09 = imem02_in[87:84];
    16: op1_10_in09 = reg_0537;
    3: op1_10_in09 = reg_0437;
    17: op1_10_in09 = imem02_in[115:112];
    19: op1_10_in09 = imem02_in[115:112];
    18: op1_10_in09 = reg_0014;
    20: op1_10_in09 = reg_0257;
    21: op1_10_in09 = reg_0469;
    22: op1_10_in09 = reg_0476;
    23: op1_10_in09 = reg_0670;
    24: op1_10_in09 = reg_0664;
    25: op1_10_in09 = reg_0577;
    26: op1_10_in09 = reg_0594;
    27: op1_10_in09 = reg_0009;
    28: op1_10_in09 = reg_0241;
    29: op1_10_in09 = reg_0115;
    30: op1_10_in09 = reg_0544;
    31: op1_10_in09 = imem06_in[27:24];
    32: op1_10_in09 = reg_0157;
    33: op1_10_in09 = reg_0654;
    34: op1_10_in09 = reg_0624;
    35: op1_10_in09 = reg_0286;
    36: op1_10_in09 = reg_0439;
    37: op1_10_in09 = imem06_in[87:84];
    38: op1_10_in09 = reg_0455;
    67: op1_10_in09 = reg_0455;
    39: op1_10_in09 = imem02_in[63:60];
    40: op1_10_in09 = reg_0661;
    41: op1_10_in09 = reg_0270;
    42: op1_10_in09 = reg_0245;
    43: op1_10_in09 = reg_0468;
    44: op1_10_in09 = reg_0510;
    45: op1_10_in09 = reg_0285;
    46: op1_10_in09 = reg_0688;
    47: op1_10_in09 = imem04_in[83:80];
    48: op1_10_in09 = reg_0732;
    49: op1_10_in09 = imem03_in[127:124];
    50: op1_10_in09 = reg_0355;
    51: op1_10_in09 = reg_0470;
    52: op1_10_in09 = imem02_in[55:52];
    53: op1_10_in09 = imem02_in[3:0];
    54: op1_10_in09 = reg_0501;
    55: op1_10_in09 = imem05_in[123:120];
    56: op1_10_in09 = reg_0275;
    77: op1_10_in09 = reg_0275;
    57: op1_10_in09 = reg_0148;
    65: op1_10_in09 = reg_0148;
    58: op1_10_in09 = reg_0372;
    59: op1_10_in09 = reg_0607;
    60: op1_10_in09 = reg_0268;
    61: op1_10_in09 = reg_0255;
    62: op1_10_in09 = reg_0385;
    63: op1_10_in09 = imem04_in[15:12];
    64: op1_10_in09 = reg_0112;
    66: op1_10_in09 = reg_0304;
    68: op1_10_in09 = reg_0678;
    69: op1_10_in09 = reg_0408;
    70: op1_10_in09 = reg_0061;
    71: op1_10_in09 = imem04_in[3:0];
    72: op1_10_in09 = reg_0813;
    73: op1_10_in09 = reg_0103;
    74: op1_10_in09 = reg_0182;
    75: op1_10_in09 = reg_0473;
    76: op1_10_in09 = reg_0642;
    78: op1_10_in09 = imem04_in[67:64];
    79: op1_10_in09 = reg_0238;
    80: op1_10_in09 = reg_0086;
    81: op1_10_in09 = reg_0742;
    82: op1_10_in09 = reg_0281;
    83: op1_10_in09 = reg_0744;
    84: op1_10_in09 = reg_0393;
    86: op1_10_in09 = reg_0057;
    87: op1_10_in09 = reg_0666;
    88: op1_10_in09 = reg_0256;
    89: op1_10_in09 = reg_0069;
    90: op1_10_in09 = reg_0069;
    91: op1_10_in09 = reg_0621;
    92: op1_10_in09 = reg_0454;
    93: op1_10_in09 = reg_0466;
    94: op1_10_in09 = reg_0461;
    95: op1_10_in09 = imem01_in[119:116];
    default: op1_10_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv09 = 1;
    12: op1_10_inv09 = 1;
    15: op1_10_inv09 = 1;
    17: op1_10_inv09 = 1;
    20: op1_10_inv09 = 1;
    24: op1_10_inv09 = 1;
    26: op1_10_inv09 = 1;
    27: op1_10_inv09 = 1;
    28: op1_10_inv09 = 1;
    29: op1_10_inv09 = 1;
    30: op1_10_inv09 = 1;
    32: op1_10_inv09 = 1;
    33: op1_10_inv09 = 1;
    34: op1_10_inv09 = 1;
    35: op1_10_inv09 = 1;
    38: op1_10_inv09 = 1;
    39: op1_10_inv09 = 1;
    42: op1_10_inv09 = 1;
    43: op1_10_inv09 = 1;
    44: op1_10_inv09 = 1;
    46: op1_10_inv09 = 1;
    47: op1_10_inv09 = 1;
    48: op1_10_inv09 = 1;
    49: op1_10_inv09 = 1;
    52: op1_10_inv09 = 1;
    53: op1_10_inv09 = 1;
    55: op1_10_inv09 = 1;
    56: op1_10_inv09 = 1;
    57: op1_10_inv09 = 1;
    58: op1_10_inv09 = 1;
    59: op1_10_inv09 = 1;
    61: op1_10_inv09 = 1;
    62: op1_10_inv09 = 1;
    65: op1_10_inv09 = 1;
    66: op1_10_inv09 = 1;
    67: op1_10_inv09 = 1;
    68: op1_10_inv09 = 1;
    69: op1_10_inv09 = 1;
    72: op1_10_inv09 = 1;
    75: op1_10_inv09 = 1;
    76: op1_10_inv09 = 1;
    80: op1_10_inv09 = 1;
    82: op1_10_inv09 = 1;
    84: op1_10_inv09 = 1;
    87: op1_10_inv09 = 1;
    89: op1_10_inv09 = 1;
    91: op1_10_inv09 = 1;
    92: op1_10_inv09 = 1;
    93: op1_10_inv09 = 1;
    95: op1_10_inv09 = 1;
    default: op1_10_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in10 = reg_0473;
    5: op1_10_in10 = reg_0457;
    6: op1_10_in10 = imem03_in[47:44];
    7: op1_10_in10 = reg_0154;
    8: op1_10_in10 = reg_0456;
    51: op1_10_in10 = reg_0456;
    9: op1_10_in10 = reg_0406;
    10: op1_10_in10 = reg_0051;
    11: op1_10_in10 = imem07_in[95:92];
    12: op1_10_in10 = reg_0808;
    13: op1_10_in10 = imem05_in[123:120];
    14: op1_10_in10 = imem07_in[3:0];
    15: op1_10_in10 = reg_0642;
    16: op1_10_in10 = reg_0541;
    3: op1_10_in10 = reg_0435;
    17: op1_10_in10 = imem02_in[127:124];
    19: op1_10_in10 = imem02_in[127:124];
    18: op1_10_in10 = reg_0008;
    20: op1_10_in10 = reg_0061;
    21: op1_10_in10 = reg_0480;
    22: op1_10_in10 = reg_0466;
    23: op1_10_in10 = reg_0679;
    24: op1_10_in10 = reg_0647;
    25: op1_10_in10 = reg_0618;
    26: op1_10_in10 = reg_0578;
    27: op1_10_in10 = reg_0809;
    28: op1_10_in10 = reg_0511;
    29: op1_10_in10 = reg_0110;
    30: op1_10_in10 = reg_0056;
    31: op1_10_in10 = imem06_in[35:32];
    32: op1_10_in10 = reg_0158;
    33: op1_10_in10 = reg_0660;
    34: op1_10_in10 = reg_0620;
    58: op1_10_in10 = reg_0620;
    35: op1_10_in10 = reg_0609;
    36: op1_10_in10 = reg_0449;
    37: op1_10_in10 = imem06_in[107:104];
    38: op1_10_in10 = reg_0469;
    39: op1_10_in10 = imem02_in[79:76];
    40: op1_10_in10 = reg_0639;
    41: op1_10_in10 = reg_0776;
    42: op1_10_in10 = reg_0301;
    43: op1_10_in10 = reg_0214;
    44: op1_10_in10 = reg_0516;
    45: op1_10_in10 = reg_0086;
    46: op1_10_in10 = reg_0673;
    47: op1_10_in10 = imem04_in[107:104];
    48: op1_10_in10 = reg_0285;
    49: op1_10_in10 = reg_0582;
    50: op1_10_in10 = reg_0426;
    52: op1_10_in10 = imem02_in[67:64];
    53: op1_10_in10 = imem02_in[111:108];
    54: op1_10_in10 = reg_0519;
    55: op1_10_in10 = reg_0309;
    56: op1_10_in10 = imem05_in[31:28];
    57: op1_10_in10 = reg_0149;
    59: op1_10_in10 = reg_0819;
    60: op1_10_in10 = reg_0159;
    61: op1_10_in10 = reg_0117;
    62: op1_10_in10 = reg_0569;
    63: op1_10_in10 = imem04_in[23:20];
    64: op1_10_in10 = reg_0486;
    65: op1_10_in10 = reg_0133;
    66: op1_10_in10 = reg_0742;
    67: op1_10_in10 = reg_0467;
    68: op1_10_in10 = imem02_in[43:40];
    69: op1_10_in10 = reg_0654;
    70: op1_10_in10 = reg_0434;
    71: op1_10_in10 = imem04_in[7:4];
    72: op1_10_in10 = reg_0794;
    73: op1_10_in10 = reg_0278;
    74: op1_10_in10 = reg_0177;
    75: op1_10_in10 = reg_0471;
    76: op1_10_in10 = reg_0142;
    77: op1_10_in10 = reg_0358;
    78: op1_10_in10 = imem04_in[71:68];
    79: op1_10_in10 = reg_0404;
    80: op1_10_in10 = reg_0728;
    81: op1_10_in10 = imem06_in[55:52];
    82: op1_10_in10 = reg_0357;
    83: op1_10_in10 = reg_0658;
    84: op1_10_in10 = reg_0383;
    86: op1_10_in10 = reg_0392;
    87: op1_10_in10 = reg_0795;
    88: op1_10_in10 = reg_0356;
    89: op1_10_in10 = reg_0780;
    90: op1_10_in10 = reg_0513;
    91: op1_10_in10 = imem07_in[75:72];
    92: op1_10_in10 = reg_0461;
    93: op1_10_in10 = reg_0472;
    94: op1_10_in10 = reg_0460;
    95: op1_10_in10 = reg_0062;
    default: op1_10_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_10_inv10 = 1;
    12: op1_10_inv10 = 1;
    16: op1_10_inv10 = 1;
    3: op1_10_inv10 = 1;
    20: op1_10_inv10 = 1;
    23: op1_10_inv10 = 1;
    25: op1_10_inv10 = 1;
    27: op1_10_inv10 = 1;
    31: op1_10_inv10 = 1;
    32: op1_10_inv10 = 1;
    34: op1_10_inv10 = 1;
    36: op1_10_inv10 = 1;
    43: op1_10_inv10 = 1;
    44: op1_10_inv10 = 1;
    45: op1_10_inv10 = 1;
    49: op1_10_inv10 = 1;
    50: op1_10_inv10 = 1;
    52: op1_10_inv10 = 1;
    53: op1_10_inv10 = 1;
    54: op1_10_inv10 = 1;
    55: op1_10_inv10 = 1;
    57: op1_10_inv10 = 1;
    58: op1_10_inv10 = 1;
    60: op1_10_inv10 = 1;
    64: op1_10_inv10 = 1;
    67: op1_10_inv10 = 1;
    68: op1_10_inv10 = 1;
    69: op1_10_inv10 = 1;
    73: op1_10_inv10 = 1;
    74: op1_10_inv10 = 1;
    78: op1_10_inv10 = 1;
    79: op1_10_inv10 = 1;
    80: op1_10_inv10 = 1;
    81: op1_10_inv10 = 1;
    82: op1_10_inv10 = 1;
    89: op1_10_inv10 = 1;
    92: op1_10_inv10 = 1;
    93: op1_10_inv10 = 1;
    94: op1_10_inv10 = 1;
    default: op1_10_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in11 = reg_0459;
    75: op1_10_in11 = reg_0459;
    5: op1_10_in11 = reg_0469;
    6: op1_10_in11 = imem03_in[79:76];
    7: op1_10_in11 = reg_0140;
    8: op1_10_in11 = reg_0209;
    9: op1_10_in11 = reg_0367;
    10: op1_10_in11 = reg_0094;
    11: op1_10_in11 = imem07_in[103:100];
    12: op1_10_in11 = reg_0013;
    13: op1_10_in11 = reg_0788;
    66: op1_10_in11 = reg_0788;
    14: op1_10_in11 = imem07_in[7:4];
    15: op1_10_in11 = reg_0650;
    16: op1_10_in11 = reg_0300;
    3: op1_10_in11 = reg_0174;
    17: op1_10_in11 = reg_0658;
    18: op1_10_in11 = reg_0809;
    19: op1_10_in11 = reg_0645;
    20: op1_10_in11 = reg_0281;
    21: op1_10_in11 = reg_0473;
    38: op1_10_in11 = reg_0473;
    94: op1_10_in11 = reg_0473;
    22: op1_10_in11 = reg_0187;
    23: op1_10_in11 = reg_0673;
    24: op1_10_in11 = reg_0352;
    25: op1_10_in11 = reg_0408;
    26: op1_10_in11 = reg_0393;
    27: op1_10_in11 = imem04_in[87:84];
    28: op1_10_in11 = reg_0217;
    29: op1_10_in11 = imem02_in[3:0];
    30: op1_10_in11 = reg_0554;
    31: op1_10_in11 = imem06_in[67:64];
    33: op1_10_in11 = reg_0640;
    34: op1_10_in11 = reg_0632;
    35: op1_10_in11 = reg_0608;
    36: op1_10_in11 = reg_0427;
    37: op1_10_in11 = reg_0630;
    39: op1_10_in11 = imem02_in[111:108];
    40: op1_10_in11 = reg_0649;
    41: op1_10_in11 = reg_0038;
    42: op1_10_in11 = reg_0355;
    43: op1_10_in11 = reg_0198;
    44: op1_10_in11 = reg_0280;
    45: op1_10_in11 = reg_0089;
    46: op1_10_in11 = reg_0699;
    47: op1_10_in11 = imem04_in[111:108];
    48: op1_10_in11 = reg_0148;
    84: op1_10_in11 = reg_0148;
    49: op1_10_in11 = reg_0591;
    50: op1_10_in11 = reg_0362;
    51: op1_10_in11 = reg_0478;
    52: op1_10_in11 = imem02_in[71:68];
    53: op1_10_in11 = reg_0642;
    54: op1_10_in11 = reg_0275;
    55: op1_10_in11 = reg_0256;
    56: op1_10_in11 = imem05_in[83:80];
    57: op1_10_in11 = reg_0135;
    58: op1_10_in11 = reg_0819;
    59: op1_10_in11 = reg_0368;
    61: op1_10_in11 = reg_0247;
    62: op1_10_in11 = reg_0000;
    63: op1_10_in11 = imem04_in[39:36];
    64: op1_10_in11 = imem05_in[15:12];
    65: op1_10_in11 = reg_0142;
    67: op1_10_in11 = reg_0468;
    93: op1_10_in11 = reg_0468;
    68: op1_10_in11 = imem02_in[47:44];
    69: op1_10_in11 = reg_0375;
    70: op1_10_in11 = reg_0449;
    71: op1_10_in11 = imem04_in[23:20];
    72: op1_10_in11 = reg_0818;
    73: op1_10_in11 = reg_0383;
    74: op1_10_in11 = reg_0173;
    76: op1_10_in11 = reg_0325;
    77: op1_10_in11 = reg_0565;
    78: op1_10_in11 = imem04_in[103:100];
    79: op1_10_in11 = reg_0613;
    80: op1_10_in11 = reg_0160;
    81: op1_10_in11 = imem06_in[59:56];
    82: op1_10_in11 = reg_0733;
    83: op1_10_in11 = reg_0691;
    86: op1_10_in11 = reg_0075;
    87: op1_10_in11 = reg_0782;
    88: op1_10_in11 = reg_0353;
    89: op1_10_in11 = reg_0513;
    90: op1_10_in11 = imem05_in[19:16];
    91: op1_10_in11 = imem07_in[87:84];
    92: op1_10_in11 = reg_0477;
    95: op1_10_in11 = reg_0111;
    default: op1_10_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv11 = 1;
    7: op1_10_inv11 = 1;
    12: op1_10_inv11 = 1;
    14: op1_10_inv11 = 1;
    15: op1_10_inv11 = 1;
    16: op1_10_inv11 = 1;
    3: op1_10_inv11 = 1;
    17: op1_10_inv11 = 1;
    19: op1_10_inv11 = 1;
    25: op1_10_inv11 = 1;
    26: op1_10_inv11 = 1;
    27: op1_10_inv11 = 1;
    28: op1_10_inv11 = 1;
    29: op1_10_inv11 = 1;
    30: op1_10_inv11 = 1;
    31: op1_10_inv11 = 1;
    34: op1_10_inv11 = 1;
    36: op1_10_inv11 = 1;
    37: op1_10_inv11 = 1;
    38: op1_10_inv11 = 1;
    44: op1_10_inv11 = 1;
    45: op1_10_inv11 = 1;
    46: op1_10_inv11 = 1;
    49: op1_10_inv11 = 1;
    50: op1_10_inv11 = 1;
    55: op1_10_inv11 = 1;
    59: op1_10_inv11 = 1;
    61: op1_10_inv11 = 1;
    63: op1_10_inv11 = 1;
    64: op1_10_inv11 = 1;
    66: op1_10_inv11 = 1;
    67: op1_10_inv11 = 1;
    70: op1_10_inv11 = 1;
    74: op1_10_inv11 = 1;
    75: op1_10_inv11 = 1;
    76: op1_10_inv11 = 1;
    77: op1_10_inv11 = 1;
    80: op1_10_inv11 = 1;
    82: op1_10_inv11 = 1;
    84: op1_10_inv11 = 1;
    87: op1_10_inv11 = 1;
    88: op1_10_inv11 = 1;
    92: op1_10_inv11 = 1;
    94: op1_10_inv11 = 1;
    default: op1_10_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in12 = reg_0452;
    5: op1_10_in12 = reg_0476;
    6: op1_10_in12 = reg_0572;
    7: op1_10_in12 = reg_0134;
    8: op1_10_in12 = reg_0205;
    9: op1_10_in12 = reg_0380;
    10: op1_10_in12 = reg_0093;
    11: op1_10_in12 = imem07_in[123:120];
    12: op1_10_in12 = reg_0807;
    13: op1_10_in12 = reg_0784;
    14: op1_10_in12 = imem07_in[15:12];
    15: op1_10_in12 = reg_0643;
    16: op1_10_in12 = reg_0299;
    3: op1_10_in12 = reg_0179;
    17: op1_10_in12 = reg_0653;
    18: op1_10_in12 = reg_0004;
    19: op1_10_in12 = reg_0661;
    20: op1_10_in12 = reg_0062;
    21: op1_10_in12 = reg_0470;
    22: op1_10_in12 = reg_0194;
    23: op1_10_in12 = reg_0669;
    24: op1_10_in12 = reg_0341;
    25: op1_10_in12 = reg_0386;
    26: op1_10_in12 = imem04_in[3:0];
    27: op1_10_in12 = imem04_in[103:100];
    28: op1_10_in12 = reg_0242;
    29: op1_10_in12 = imem02_in[23:20];
    30: op1_10_in12 = reg_0556;
    31: op1_10_in12 = imem06_in[71:68];
    33: op1_10_in12 = reg_0638;
    34: op1_10_in12 = reg_0627;
    35: op1_10_in12 = reg_0236;
    36: op1_10_in12 = reg_0438;
    37: op1_10_in12 = reg_0371;
    38: op1_10_in12 = reg_0474;
    94: op1_10_in12 = reg_0474;
    39: op1_10_in12 = imem02_in[119:116];
    40: op1_10_in12 = reg_0357;
    41: op1_10_in12 = reg_0576;
    42: op1_10_in12 = reg_0709;
    43: op1_10_in12 = reg_0197;
    44: op1_10_in12 = reg_0631;
    45: op1_10_in12 = reg_0136;
    46: op1_10_in12 = reg_0475;
    47: op1_10_in12 = reg_0544;
    48: op1_10_in12 = reg_0145;
    49: op1_10_in12 = reg_0594;
    50: op1_10_in12 = reg_0361;
    77: op1_10_in12 = reg_0361;
    51: op1_10_in12 = reg_0208;
    52: op1_10_in12 = imem02_in[91:88];
    53: op1_10_in12 = reg_0650;
    54: op1_10_in12 = imem05_in[3:0];
    55: op1_10_in12 = reg_0279;
    56: op1_10_in12 = imem05_in[115:112];
    57: op1_10_in12 = reg_0152;
    58: op1_10_in12 = reg_0231;
    59: op1_10_in12 = reg_0029;
    61: op1_10_in12 = reg_0692;
    62: op1_10_in12 = reg_0809;
    63: op1_10_in12 = imem04_in[71:68];
    64: op1_10_in12 = imem05_in[39:36];
    65: op1_10_in12 = imem06_in[3:0];
    66: op1_10_in12 = reg_0795;
    67: op1_10_in12 = reg_0210;
    75: op1_10_in12 = reg_0210;
    68: op1_10_in12 = imem02_in[79:76];
    69: op1_10_in12 = reg_0583;
    70: op1_10_in12 = reg_0444;
    71: op1_10_in12 = imem04_in[31:28];
    72: op1_10_in12 = reg_0787;
    73: op1_10_in12 = imem05_in[19:16];
    76: op1_10_in12 = reg_0141;
    78: op1_10_in12 = imem04_in[107:104];
    79: op1_10_in12 = reg_0405;
    80: op1_10_in12 = reg_0725;
    81: op1_10_in12 = imem06_in[83:80];
    82: op1_10_in12 = reg_0396;
    83: op1_10_in12 = reg_0407;
    84: op1_10_in12 = reg_0781;
    86: op1_10_in12 = reg_0304;
    87: op1_10_in12 = reg_0245;
    88: op1_10_in12 = reg_0406;
    89: op1_10_in12 = reg_0259;
    90: op1_10_in12 = imem05_in[35:32];
    91: op1_10_in12 = imem07_in[115:112];
    92: op1_10_in12 = reg_0462;
    93: op1_10_in12 = reg_0479;
    95: op1_10_in12 = reg_0567;
    default: op1_10_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv12 = 1;
    6: op1_10_inv12 = 1;
    7: op1_10_inv12 = 1;
    11: op1_10_inv12 = 1;
    12: op1_10_inv12 = 1;
    14: op1_10_inv12 = 1;
    15: op1_10_inv12 = 1;
    20: op1_10_inv12 = 1;
    22: op1_10_inv12 = 1;
    25: op1_10_inv12 = 1;
    26: op1_10_inv12 = 1;
    28: op1_10_inv12 = 1;
    31: op1_10_inv12 = 1;
    36: op1_10_inv12 = 1;
    40: op1_10_inv12 = 1;
    41: op1_10_inv12 = 1;
    42: op1_10_inv12 = 1;
    43: op1_10_inv12 = 1;
    50: op1_10_inv12 = 1;
    53: op1_10_inv12 = 1;
    57: op1_10_inv12 = 1;
    64: op1_10_inv12 = 1;
    66: op1_10_inv12 = 1;
    68: op1_10_inv12 = 1;
    71: op1_10_inv12 = 1;
    73: op1_10_inv12 = 1;
    77: op1_10_inv12 = 1;
    80: op1_10_inv12 = 1;
    84: op1_10_inv12 = 1;
    87: op1_10_inv12 = 1;
    89: op1_10_inv12 = 1;
    93: op1_10_inv12 = 1;
    95: op1_10_inv12 = 1;
    default: op1_10_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in13 = reg_0456;
    93: op1_10_in13 = reg_0456;
    5: op1_10_in13 = reg_0466;
    6: op1_10_in13 = reg_0593;
    7: op1_10_in13 = imem06_in[3:0];
    8: op1_10_in13 = reg_0195;
    9: op1_10_in13 = reg_0039;
    10: op1_10_in13 = imem03_in[15:12];
    11: op1_10_in13 = imem07_in[127:124];
    12: op1_10_in13 = reg_0010;
    13: op1_10_in13 = reg_0736;
    14: op1_10_in13 = imem07_in[39:36];
    15: op1_10_in13 = reg_0659;
    16: op1_10_in13 = reg_0289;
    3: op1_10_in13 = reg_0170;
    17: op1_10_in13 = reg_0661;
    52: op1_10_in13 = reg_0661;
    18: op1_10_in13 = reg_0277;
    19: op1_10_in13 = reg_0647;
    20: op1_10_in13 = reg_0074;
    21: op1_10_in13 = reg_0459;
    22: op1_10_in13 = imem01_in[15:12];
    23: op1_10_in13 = reg_0453;
    24: op1_10_in13 = reg_0359;
    40: op1_10_in13 = reg_0359;
    25: op1_10_in13 = reg_0375;
    26: op1_10_in13 = imem04_in[19:16];
    27: op1_10_in13 = imem04_in[107:104];
    28: op1_10_in13 = reg_0244;
    29: op1_10_in13 = imem02_in[27:24];
    30: op1_10_in13 = reg_0529;
    31: op1_10_in13 = imem06_in[79:76];
    33: op1_10_in13 = reg_0665;
    34: op1_10_in13 = reg_0622;
    35: op1_10_in13 = imem06_in[35:32];
    36: op1_10_in13 = reg_0167;
    37: op1_10_in13 = reg_0606;
    38: op1_10_in13 = reg_0478;
    39: op1_10_in13 = imem02_in[123:120];
    41: op1_10_in13 = reg_0753;
    42: op1_10_in13 = imem07_in[71:68];
    43: op1_10_in13 = imem01_in[19:16];
    44: op1_10_in13 = reg_0626;
    45: op1_10_in13 = reg_0152;
    46: op1_10_in13 = reg_0452;
    47: op1_10_in13 = reg_0055;
    48: op1_10_in13 = reg_0128;
    49: op1_10_in13 = reg_0387;
    50: op1_10_in13 = reg_0363;
    77: op1_10_in13 = reg_0363;
    51: op1_10_in13 = reg_0191;
    53: op1_10_in13 = reg_0655;
    54: op1_10_in13 = imem05_in[55:52];
    55: op1_10_in13 = reg_0224;
    56: op1_10_in13 = reg_0792;
    57: op1_10_in13 = reg_0142;
    58: op1_10_in13 = reg_0632;
    59: op1_10_in13 = reg_0632;
    61: op1_10_in13 = reg_0634;
    62: op1_10_in13 = imem04_in[15:12];
    63: op1_10_in13 = reg_0059;
    64: op1_10_in13 = imem05_in[63:60];
    65: op1_10_in13 = imem06_in[31:28];
    66: op1_10_in13 = reg_0793;
    67: op1_10_in13 = reg_0209;
    68: op1_10_in13 = imem02_in[87:84];
    69: op1_10_in13 = reg_0819;
    70: op1_10_in13 = reg_0435;
    71: op1_10_in13 = imem04_in[43:40];
    72: op1_10_in13 = imem07_in[3:0];
    73: op1_10_in13 = imem06_in[11:8];
    75: op1_10_in13 = reg_0186;
    76: op1_10_in13 = reg_0427;
    78: op1_10_in13 = imem04_in[123:120];
    79: op1_10_in13 = reg_0763;
    80: op1_10_in13 = reg_0158;
    81: op1_10_in13 = imem06_in[95:92];
    82: op1_10_in13 = reg_0003;
    83: op1_10_in13 = reg_0680;
    84: op1_10_in13 = reg_0151;
    86: op1_10_in13 = reg_0345;
    87: op1_10_in13 = reg_0488;
    88: op1_10_in13 = reg_0590;
    89: op1_10_in13 = reg_0776;
    90: op1_10_in13 = imem05_in[59:56];
    91: op1_10_in13 = reg_0716;
    92: op1_10_in13 = reg_0205;
    94: op1_10_in13 = reg_0471;
    95: op1_10_in13 = reg_0051;
    default: op1_10_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv13 = 1;
    5: op1_10_inv13 = 1;
    6: op1_10_inv13 = 1;
    10: op1_10_inv13 = 1;
    16: op1_10_inv13 = 1;
    18: op1_10_inv13 = 1;
    19: op1_10_inv13 = 1;
    20: op1_10_inv13 = 1;
    21: op1_10_inv13 = 1;
    22: op1_10_inv13 = 1;
    27: op1_10_inv13 = 1;
    34: op1_10_inv13 = 1;
    35: op1_10_inv13 = 1;
    36: op1_10_inv13 = 1;
    37: op1_10_inv13 = 1;
    40: op1_10_inv13 = 1;
    42: op1_10_inv13 = 1;
    45: op1_10_inv13 = 1;
    46: op1_10_inv13 = 1;
    48: op1_10_inv13 = 1;
    51: op1_10_inv13 = 1;
    53: op1_10_inv13 = 1;
    54: op1_10_inv13 = 1;
    56: op1_10_inv13 = 1;
    58: op1_10_inv13 = 1;
    59: op1_10_inv13 = 1;
    61: op1_10_inv13 = 1;
    62: op1_10_inv13 = 1;
    65: op1_10_inv13 = 1;
    66: op1_10_inv13 = 1;
    67: op1_10_inv13 = 1;
    70: op1_10_inv13 = 1;
    71: op1_10_inv13 = 1;
    73: op1_10_inv13 = 1;
    76: op1_10_inv13 = 1;
    77: op1_10_inv13 = 1;
    80: op1_10_inv13 = 1;
    82: op1_10_inv13 = 1;
    84: op1_10_inv13 = 1;
    86: op1_10_inv13 = 1;
    88: op1_10_inv13 = 1;
    90: op1_10_inv13 = 1;
    91: op1_10_inv13 = 1;
    95: op1_10_inv13 = 1;
    default: op1_10_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in14 = reg_0191;
    5: op1_10_in14 = reg_0470;
    6: op1_10_in14 = reg_0395;
    7: op1_10_in14 = imem06_in[15:12];
    8: op1_10_in14 = imem01_in[35:32];
    75: op1_10_in14 = imem01_in[35:32];
    9: op1_10_in14 = reg_0814;
    10: op1_10_in14 = imem03_in[19:16];
    11: op1_10_in14 = reg_0731;
    12: op1_10_in14 = imem04_in[11:8];
    13: op1_10_in14 = reg_0733;
    14: op1_10_in14 = imem07_in[95:92];
    15: op1_10_in14 = reg_0352;
    16: op1_10_in14 = reg_0306;
    3: op1_10_in14 = reg_0176;
    17: op1_10_in14 = reg_0641;
    18: op1_10_in14 = reg_0276;
    19: op1_10_in14 = reg_0640;
    20: op1_10_in14 = reg_0072;
    21: op1_10_in14 = reg_0209;
    22: op1_10_in14 = imem01_in[59:56];
    23: op1_10_in14 = reg_0450;
    24: op1_10_in14 = reg_0345;
    25: op1_10_in14 = reg_0404;
    26: op1_10_in14 = imem04_in[27:24];
    27: op1_10_in14 = reg_0059;
    78: op1_10_in14 = reg_0059;
    28: op1_10_in14 = reg_0503;
    29: op1_10_in14 = imem02_in[47:44];
    30: op1_10_in14 = reg_0290;
    31: op1_10_in14 = imem06_in[103:100];
    33: op1_10_in14 = reg_0652;
    34: op1_10_in14 = reg_0402;
    35: op1_10_in14 = imem06_in[51:48];
    36: op1_10_in14 = reg_0169;
    37: op1_10_in14 = reg_0618;
    38: op1_10_in14 = reg_0198;
    39: op1_10_in14 = imem02_in[127:124];
    40: op1_10_in14 = reg_0348;
    41: op1_10_in14 = reg_0620;
    42: op1_10_in14 = imem07_in[107:104];
    43: op1_10_in14 = imem01_in[23:20];
    44: op1_10_in14 = reg_0258;
    45: op1_10_in14 = reg_0130;
    46: op1_10_in14 = reg_0456;
    47: op1_10_in14 = reg_0303;
    48: op1_10_in14 = reg_0154;
    49: op1_10_in14 = reg_0561;
    50: op1_10_in14 = reg_0324;
    51: op1_10_in14 = reg_0186;
    52: op1_10_in14 = reg_0651;
    53: op1_10_in14 = reg_0659;
    54: op1_10_in14 = imem05_in[79:76];
    55: op1_10_in14 = reg_0132;
    56: op1_10_in14 = reg_0797;
    57: op1_10_in14 = reg_0137;
    58: op1_10_in14 = reg_0236;
    59: op1_10_in14 = imem07_in[39:36];
    61: op1_10_in14 = reg_0473;
    62: op1_10_in14 = imem04_in[51:48];
    63: op1_10_in14 = reg_0055;
    64: op1_10_in14 = imem05_in[67:64];
    65: op1_10_in14 = imem06_in[43:40];
    66: op1_10_in14 = reg_0227;
    67: op1_10_in14 = imem01_in[7:4];
    68: op1_10_in14 = imem02_in[103:100];
    69: op1_10_in14 = reg_0787;
    70: op1_10_in14 = reg_0161;
    91: op1_10_in14 = reg_0161;
    71: op1_10_in14 = imem04_in[47:44];
    72: op1_10_in14 = imem07_in[7:4];
    73: op1_10_in14 = imem06_in[63:60];
    76: op1_10_in14 = reg_0587;
    77: op1_10_in14 = reg_0594;
    79: op1_10_in14 = reg_0593;
    80: op1_10_in14 = reg_0253;
    81: op1_10_in14 = imem06_in[99:96];
    82: op1_10_in14 = reg_0801;
    83: op1_10_in14 = reg_0454;
    84: op1_10_in14 = reg_0830;
    86: op1_10_in14 = reg_0363;
    87: op1_10_in14 = reg_0583;
    88: op1_10_in14 = reg_0514;
    89: op1_10_in14 = imem05_in[27:24];
    90: op1_10_in14 = imem05_in[71:68];
    92: op1_10_in14 = reg_0522;
    93: op1_10_in14 = reg_0458;
    94: op1_10_in14 = reg_0200;
    95: op1_10_in14 = reg_0260;
    default: op1_10_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv14 = 1;
    5: op1_10_inv14 = 1;
    7: op1_10_inv14 = 1;
    8: op1_10_inv14 = 1;
    11: op1_10_inv14 = 1;
    12: op1_10_inv14 = 1;
    13: op1_10_inv14 = 1;
    14: op1_10_inv14 = 1;
    16: op1_10_inv14 = 1;
    23: op1_10_inv14 = 1;
    24: op1_10_inv14 = 1;
    26: op1_10_inv14 = 1;
    28: op1_10_inv14 = 1;
    29: op1_10_inv14 = 1;
    36: op1_10_inv14 = 1;
    39: op1_10_inv14 = 1;
    40: op1_10_inv14 = 1;
    41: op1_10_inv14 = 1;
    43: op1_10_inv14 = 1;
    44: op1_10_inv14 = 1;
    45: op1_10_inv14 = 1;
    46: op1_10_inv14 = 1;
    48: op1_10_inv14 = 1;
    52: op1_10_inv14 = 1;
    53: op1_10_inv14 = 1;
    54: op1_10_inv14 = 1;
    55: op1_10_inv14 = 1;
    61: op1_10_inv14 = 1;
    64: op1_10_inv14 = 1;
    66: op1_10_inv14 = 1;
    67: op1_10_inv14 = 1;
    70: op1_10_inv14 = 1;
    71: op1_10_inv14 = 1;
    72: op1_10_inv14 = 1;
    73: op1_10_inv14 = 1;
    77: op1_10_inv14 = 1;
    78: op1_10_inv14 = 1;
    81: op1_10_inv14 = 1;
    83: op1_10_inv14 = 1;
    84: op1_10_inv14 = 1;
    87: op1_10_inv14 = 1;
    90: op1_10_inv14 = 1;
    91: op1_10_inv14 = 1;
    92: op1_10_inv14 = 1;
    93: op1_10_inv14 = 1;
    94: op1_10_inv14 = 1;
    default: op1_10_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in15 = reg_0210;
    5: op1_10_in15 = reg_0203;
    21: op1_10_in15 = reg_0203;
    94: op1_10_in15 = reg_0203;
    6: op1_10_in15 = reg_0391;
    7: op1_10_in15 = imem06_in[47:44];
    8: op1_10_in15 = imem01_in[55:52];
    67: op1_10_in15 = imem01_in[55:52];
    9: op1_10_in15 = reg_0036;
    10: op1_10_in15 = imem03_in[47:44];
    11: op1_10_in15 = reg_0702;
    12: op1_10_in15 = imem04_in[59:56];
    13: op1_10_in15 = reg_0264;
    14: op1_10_in15 = imem07_in[103:100];
    15: op1_10_in15 = reg_0364;
    16: op1_10_in15 = reg_0302;
    3: op1_10_in15 = reg_0158;
    17: op1_10_in15 = reg_0325;
    18: op1_10_in15 = reg_0226;
    19: op1_10_in15 = reg_0649;
    20: op1_10_in15 = imem05_in[11:8];
    22: op1_10_in15 = imem01_in[79:76];
    23: op1_10_in15 = reg_0464;
    24: op1_10_in15 = reg_0363;
    25: op1_10_in15 = reg_0753;
    26: op1_10_in15 = imem04_in[43:40];
    27: op1_10_in15 = reg_0262;
    28: op1_10_in15 = reg_0237;
    29: op1_10_in15 = imem02_in[123:120];
    30: op1_10_in15 = reg_0291;
    31: op1_10_in15 = imem07_in[3:0];
    33: op1_10_in15 = reg_0359;
    34: op1_10_in15 = reg_0317;
    35: op1_10_in15 = imem06_in[71:68];
    36: op1_10_in15 = reg_0170;
    37: op1_10_in15 = reg_0627;
    38: op1_10_in15 = reg_0196;
    39: op1_10_in15 = reg_0666;
    40: op1_10_in15 = reg_0353;
    77: op1_10_in15 = reg_0353;
    41: op1_10_in15 = reg_0819;
    42: op1_10_in15 = imem07_in[115:112];
    43: op1_10_in15 = imem01_in[27:24];
    44: op1_10_in15 = reg_0070;
    45: op1_10_in15 = reg_0155;
    46: op1_10_in15 = reg_0209;
    47: op1_10_in15 = reg_0611;
    48: op1_10_in15 = reg_0139;
    49: op1_10_in15 = reg_0386;
    50: op1_10_in15 = reg_0541;
    51: op1_10_in15 = reg_0194;
    93: op1_10_in15 = reg_0194;
    52: op1_10_in15 = reg_0662;
    53: op1_10_in15 = reg_0341;
    54: op1_10_in15 = imem05_in[103:100];
    55: op1_10_in15 = reg_0154;
    56: op1_10_in15 = reg_0091;
    57: op1_10_in15 = reg_0109;
    58: op1_10_in15 = reg_0623;
    59: op1_10_in15 = imem07_in[67:64];
    61: op1_10_in15 = reg_0467;
    62: op1_10_in15 = imem04_in[67:64];
    63: op1_10_in15 = reg_0057;
    64: op1_10_in15 = imem05_in[87:84];
    65: op1_10_in15 = imem06_in[55:52];
    66: op1_10_in15 = reg_0039;
    68: op1_10_in15 = imem02_in[107:104];
    69: op1_10_in15 = reg_0767;
    70: op1_10_in15 = reg_0169;
    71: op1_10_in15 = imem04_in[75:72];
    72: op1_10_in15 = imem07_in[35:32];
    73: op1_10_in15 = imem06_in[91:88];
    75: op1_10_in15 = imem01_in[63:60];
    76: op1_10_in15 = reg_0358;
    78: op1_10_in15 = reg_0560;
    79: op1_10_in15 = reg_0663;
    80: op1_10_in15 = reg_0636;
    81: op1_10_in15 = imem06_in[111:108];
    82: op1_10_in15 = reg_0015;
    83: op1_10_in15 = reg_0450;
    84: op1_10_in15 = reg_0156;
    86: op1_10_in15 = reg_0590;
    87: op1_10_in15 = reg_0252;
    88: op1_10_in15 = reg_0093;
    89: op1_10_in15 = reg_0135;
    90: op1_10_in15 = imem05_in[91:88];
    91: op1_10_in15 = reg_0167;
    92: op1_10_in15 = reg_0421;
    95: op1_10_in15 = reg_0425;
    default: op1_10_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv15 = 1;
    7: op1_10_inv15 = 1;
    14: op1_10_inv15 = 1;
    15: op1_10_inv15 = 1;
    16: op1_10_inv15 = 1;
    3: op1_10_inv15 = 1;
    17: op1_10_inv15 = 1;
    19: op1_10_inv15 = 1;
    20: op1_10_inv15 = 1;
    21: op1_10_inv15 = 1;
    24: op1_10_inv15 = 1;
    25: op1_10_inv15 = 1;
    26: op1_10_inv15 = 1;
    27: op1_10_inv15 = 1;
    28: op1_10_inv15 = 1;
    29: op1_10_inv15 = 1;
    33: op1_10_inv15 = 1;
    34: op1_10_inv15 = 1;
    36: op1_10_inv15 = 1;
    38: op1_10_inv15 = 1;
    39: op1_10_inv15 = 1;
    41: op1_10_inv15 = 1;
    43: op1_10_inv15 = 1;
    44: op1_10_inv15 = 1;
    47: op1_10_inv15 = 1;
    50: op1_10_inv15 = 1;
    51: op1_10_inv15 = 1;
    54: op1_10_inv15 = 1;
    55: op1_10_inv15 = 1;
    56: op1_10_inv15 = 1;
    58: op1_10_inv15 = 1;
    59: op1_10_inv15 = 1;
    61: op1_10_inv15 = 1;
    63: op1_10_inv15 = 1;
    66: op1_10_inv15 = 1;
    70: op1_10_inv15 = 1;
    71: op1_10_inv15 = 1;
    73: op1_10_inv15 = 1;
    75: op1_10_inv15 = 1;
    80: op1_10_inv15 = 1;
    81: op1_10_inv15 = 1;
    83: op1_10_inv15 = 1;
    87: op1_10_inv15 = 1;
    88: op1_10_inv15 = 1;
    91: op1_10_inv15 = 1;
    93: op1_10_inv15 = 1;
    94: op1_10_inv15 = 1;
    95: op1_10_inv15 = 1;
    default: op1_10_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in16 = reg_0204;
    5: op1_10_in16 = reg_0193;
    6: op1_10_in16 = reg_0362;
    7: op1_10_in16 = imem06_in[71:68];
    8: op1_10_in16 = imem01_in[111:108];
    9: op1_10_in16 = reg_0037;
    10: op1_10_in16 = imem03_in[55:52];
    11: op1_10_in16 = reg_0718;
    12: op1_10_in16 = imem04_in[87:84];
    13: op1_10_in16 = reg_0230;
    14: op1_10_in16 = imem07_in[107:104];
    15: op1_10_in16 = reg_0310;
    16: op1_10_in16 = reg_0291;
    3: op1_10_in16 = reg_0171;
    17: op1_10_in16 = reg_0359;
    18: op1_10_in16 = reg_0057;
    19: op1_10_in16 = reg_0644;
    20: op1_10_in16 = imem05_in[55:52];
    21: op1_10_in16 = reg_0207;
    22: op1_10_in16 = reg_0523;
    63: op1_10_in16 = reg_0523;
    23: op1_10_in16 = reg_0459;
    24: op1_10_in16 = reg_0365;
    25: op1_10_in16 = reg_0032;
    26: op1_10_in16 = imem04_in[103:100];
    27: op1_10_in16 = reg_0545;
    28: op1_10_in16 = reg_0234;
    29: op1_10_in16 = reg_0658;
    30: op1_10_in16 = reg_0266;
    31: op1_10_in16 = imem07_in[15:12];
    33: op1_10_in16 = reg_0322;
    34: op1_10_in16 = reg_0577;
    73: op1_10_in16 = reg_0577;
    35: op1_10_in16 = imem06_in[95:92];
    36: op1_10_in16 = reg_0184;
    37: op1_10_in16 = reg_0612;
    38: op1_10_in16 = reg_0206;
    39: op1_10_in16 = reg_0637;
    40: op1_10_in16 = reg_0321;
    41: op1_10_in16 = reg_0338;
    42: op1_10_in16 = imem07_in[123:120];
    43: op1_10_in16 = imem01_in[35:32];
    44: op1_10_in16 = reg_0796;
    45: op1_10_in16 = reg_0131;
    46: op1_10_in16 = reg_0186;
    47: op1_10_in16 = reg_0503;
    48: op1_10_in16 = reg_0130;
    49: op1_10_in16 = reg_0006;
    50: op1_10_in16 = reg_0096;
    51: op1_10_in16 = reg_0190;
    52: op1_10_in16 = reg_0548;
    53: op1_10_in16 = reg_0356;
    54: op1_10_in16 = imem05_in[111:108];
    55: op1_10_in16 = reg_0139;
    56: op1_10_in16 = reg_0215;
    57: op1_10_in16 = reg_0020;
    58: op1_10_in16 = imem07_in[31:28];
    59: op1_10_in16 = imem07_in[87:84];
    61: op1_10_in16 = reg_0470;
    62: op1_10_in16 = imem04_in[95:92];
    64: op1_10_in16 = imem05_in[91:88];
    65: op1_10_in16 = imem06_in[87:84];
    66: op1_10_in16 = reg_0277;
    67: op1_10_in16 = imem01_in[71:68];
    68: op1_10_in16 = reg_0403;
    69: op1_10_in16 = reg_0632;
    70: op1_10_in16 = reg_0182;
    71: op1_10_in16 = imem04_in[107:104];
    72: op1_10_in16 = imem07_in[43:40];
    75: op1_10_in16 = imem01_in[99:96];
    76: op1_10_in16 = reg_0320;
    77: op1_10_in16 = reg_0414;
    78: op1_10_in16 = reg_0552;
    79: op1_10_in16 = reg_0651;
    80: op1_10_in16 = reg_0053;
    81: op1_10_in16 = imem06_in[115:112];
    82: op1_10_in16 = reg_0806;
    83: op1_10_in16 = reg_0464;
    84: op1_10_in16 = reg_0143;
    86: op1_10_in16 = reg_0743;
    87: op1_10_in16 = reg_0288;
    88: op1_10_in16 = imem03_in[39:36];
    89: op1_10_in16 = reg_0355;
    90: op1_10_in16 = reg_0666;
    91: op1_10_in16 = reg_0157;
    92: op1_10_in16 = reg_0098;
    93: op1_10_in16 = reg_0198;
    94: op1_10_in16 = reg_0152;
    95: op1_10_in16 = reg_0304;
    default: op1_10_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv16 = 1;
    8: op1_10_inv16 = 1;
    9: op1_10_inv16 = 1;
    15: op1_10_inv16 = 1;
    16: op1_10_inv16 = 1;
    21: op1_10_inv16 = 1;
    22: op1_10_inv16 = 1;
    25: op1_10_inv16 = 1;
    26: op1_10_inv16 = 1;
    28: op1_10_inv16 = 1;
    29: op1_10_inv16 = 1;
    33: op1_10_inv16 = 1;
    34: op1_10_inv16 = 1;
    35: op1_10_inv16 = 1;
    36: op1_10_inv16 = 1;
    37: op1_10_inv16 = 1;
    38: op1_10_inv16 = 1;
    39: op1_10_inv16 = 1;
    40: op1_10_inv16 = 1;
    42: op1_10_inv16 = 1;
    44: op1_10_inv16 = 1;
    47: op1_10_inv16 = 1;
    48: op1_10_inv16 = 1;
    50: op1_10_inv16 = 1;
    54: op1_10_inv16 = 1;
    56: op1_10_inv16 = 1;
    58: op1_10_inv16 = 1;
    59: op1_10_inv16 = 1;
    61: op1_10_inv16 = 1;
    64: op1_10_inv16 = 1;
    66: op1_10_inv16 = 1;
    68: op1_10_inv16 = 1;
    78: op1_10_inv16 = 1;
    82: op1_10_inv16 = 1;
    84: op1_10_inv16 = 1;
    88: op1_10_inv16 = 1;
    89: op1_10_inv16 = 1;
    90: op1_10_inv16 = 1;
    91: op1_10_inv16 = 1;
    93: op1_10_inv16 = 1;
    94: op1_10_inv16 = 1;
    default: op1_10_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in17 = reg_0211;
    5: op1_10_in17 = reg_0207;
    6: op1_10_in17 = reg_0373;
    7: op1_10_in17 = imem06_in[111:108];
    8: op1_10_in17 = reg_0514;
    9: op1_10_in17 = reg_0029;
    41: op1_10_in17 = reg_0029;
    10: op1_10_in17 = imem03_in[95:92];
    11: op1_10_in17 = reg_0711;
    12: op1_10_in17 = reg_0549;
    13: op1_10_in17 = reg_0132;
    14: op1_10_in17 = reg_0722;
    15: op1_10_in17 = reg_0365;
    16: op1_10_in17 = reg_0297;
    17: op1_10_in17 = reg_0083;
    18: op1_10_in17 = reg_0224;
    19: op1_10_in17 = reg_0663;
    20: op1_10_in17 = reg_0490;
    21: op1_10_in17 = reg_0206;
    22: op1_10_in17 = reg_0820;
    92: op1_10_in17 = reg_0820;
    23: op1_10_in17 = reg_0214;
    24: op1_10_in17 = reg_0342;
    25: op1_10_in17 = imem07_in[35:32];
    26: op1_10_in17 = reg_0551;
    27: op1_10_in17 = reg_0544;
    28: op1_10_in17 = reg_0245;
    29: op1_10_in17 = reg_0656;
    30: op1_10_in17 = reg_0050;
    31: op1_10_in17 = imem07_in[39:36];
    33: op1_10_in17 = reg_0092;
    34: op1_10_in17 = reg_0408;
    35: op1_10_in17 = imem06_in[115:112];
    65: op1_10_in17 = imem06_in[115:112];
    37: op1_10_in17 = reg_0370;
    38: op1_10_in17 = imem01_in[7:4];
    51: op1_10_in17 = imem01_in[7:4];
    39: op1_10_in17 = reg_0640;
    40: op1_10_in17 = reg_0347;
    42: op1_10_in17 = reg_0181;
    43: op1_10_in17 = imem01_in[43:40];
    44: op1_10_in17 = reg_0795;
    45: op1_10_in17 = imem06_in[27:24];
    46: op1_10_in17 = imem01_in[3:0];
    47: op1_10_in17 = reg_0074;
    48: op1_10_in17 = reg_0140;
    49: op1_10_in17 = reg_0003;
    50: op1_10_in17 = reg_0535;
    52: op1_10_in17 = reg_0427;
    53: op1_10_in17 = reg_0363;
    54: op1_10_in17 = reg_0796;
    55: op1_10_in17 = reg_0138;
    56: op1_10_in17 = reg_0256;
    57: op1_10_in17 = reg_0371;
    58: op1_10_in17 = imem07_in[83:80];
    59: op1_10_in17 = imem07_in[91:88];
    61: op1_10_in17 = reg_0479;
    62: op1_10_in17 = imem04_in[119:116];
    63: op1_10_in17 = reg_0547;
    64: op1_10_in17 = imem05_in[107:104];
    66: op1_10_in17 = reg_0489;
    67: op1_10_in17 = imem01_in[115:112];
    68: op1_10_in17 = reg_0666;
    69: op1_10_in17 = imem07_in[43:40];
    70: op1_10_in17 = reg_0158;
    71: op1_10_in17 = reg_0262;
    72: op1_10_in17 = imem07_in[47:44];
    73: op1_10_in17 = reg_0624;
    75: op1_10_in17 = imem01_in[127:124];
    76: op1_10_in17 = reg_0586;
    77: op1_10_in17 = reg_0527;
    78: op1_10_in17 = reg_0056;
    79: op1_10_in17 = reg_0657;
    80: op1_10_in17 = reg_0444;
    81: op1_10_in17 = reg_0291;
    82: op1_10_in17 = reg_0809;
    83: op1_10_in17 = reg_0469;
    84: op1_10_in17 = imem06_in[7:4];
    86: op1_10_in17 = reg_0096;
    87: op1_10_in17 = reg_0254;
    88: op1_10_in17 = imem03_in[91:88];
    89: op1_10_in17 = reg_0144;
    90: op1_10_in17 = reg_0788;
    91: op1_10_in17 = reg_0295;
    93: op1_10_in17 = reg_0196;
    94: op1_10_in17 = reg_0237;
    95: op1_10_in17 = reg_0424;
    default: op1_10_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_10_inv17 = 1;
    7: op1_10_inv17 = 1;
    9: op1_10_inv17 = 1;
    11: op1_10_inv17 = 1;
    12: op1_10_inv17 = 1;
    15: op1_10_inv17 = 1;
    19: op1_10_inv17 = 1;
    20: op1_10_inv17 = 1;
    21: op1_10_inv17 = 1;
    23: op1_10_inv17 = 1;
    25: op1_10_inv17 = 1;
    27: op1_10_inv17 = 1;
    28: op1_10_inv17 = 1;
    34: op1_10_inv17 = 1;
    38: op1_10_inv17 = 1;
    39: op1_10_inv17 = 1;
    40: op1_10_inv17 = 1;
    42: op1_10_inv17 = 1;
    44: op1_10_inv17 = 1;
    46: op1_10_inv17 = 1;
    48: op1_10_inv17 = 1;
    49: op1_10_inv17 = 1;
    50: op1_10_inv17 = 1;
    52: op1_10_inv17 = 1;
    53: op1_10_inv17 = 1;
    55: op1_10_inv17 = 1;
    57: op1_10_inv17 = 1;
    58: op1_10_inv17 = 1;
    59: op1_10_inv17 = 1;
    62: op1_10_inv17 = 1;
    65: op1_10_inv17 = 1;
    66: op1_10_inv17 = 1;
    67: op1_10_inv17 = 1;
    68: op1_10_inv17 = 1;
    71: op1_10_inv17 = 1;
    75: op1_10_inv17 = 1;
    76: op1_10_inv17 = 1;
    77: op1_10_inv17 = 1;
    82: op1_10_inv17 = 1;
    87: op1_10_inv17 = 1;
    88: op1_10_inv17 = 1;
    89: op1_10_inv17 = 1;
    91: op1_10_inv17 = 1;
    92: op1_10_inv17 = 1;
    94: op1_10_inv17 = 1;
    default: op1_10_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in18 = reg_0196;
    5: op1_10_in18 = reg_0211;
    23: op1_10_in18 = reg_0211;
    6: op1_10_in18 = reg_0369;
    7: op1_10_in18 = reg_0628;
    8: op1_10_in18 = reg_0517;
    9: op1_10_in18 = reg_0749;
    10: op1_10_in18 = imem03_in[99:96];
    11: op1_10_in18 = reg_0706;
    12: op1_10_in18 = reg_0533;
    13: op1_10_in18 = reg_0129;
    14: op1_10_in18 = reg_0717;
    15: op1_10_in18 = reg_0342;
    16: op1_10_in18 = reg_0069;
    57: op1_10_in18 = reg_0069;
    17: op1_10_in18 = reg_0088;
    78: op1_10_in18 = reg_0088;
    18: op1_10_in18 = reg_0059;
    62: op1_10_in18 = reg_0059;
    19: op1_10_in18 = reg_0334;
    20: op1_10_in18 = reg_0789;
    21: op1_10_in18 = reg_0192;
    22: op1_10_in18 = reg_0778;
    24: op1_10_in18 = reg_0355;
    25: op1_10_in18 = imem07_in[55:52];
    26: op1_10_in18 = reg_0500;
    27: op1_10_in18 = reg_0315;
    28: op1_10_in18 = reg_0123;
    29: op1_10_in18 = reg_0639;
    30: op1_10_in18 = reg_0079;
    31: op1_10_in18 = reg_0726;
    33: op1_10_in18 = reg_0531;
    34: op1_10_in18 = reg_0762;
    73: op1_10_in18 = reg_0762;
    35: op1_10_in18 = reg_0408;
    37: op1_10_in18 = reg_0775;
    38: op1_10_in18 = imem01_in[11:8];
    39: op1_10_in18 = reg_0638;
    40: op1_10_in18 = reg_0092;
    41: op1_10_in18 = imem07_in[15:12];
    42: op1_10_in18 = reg_0161;
    43: op1_10_in18 = imem01_in[67:64];
    44: op1_10_in18 = reg_0493;
    45: op1_10_in18 = imem06_in[43:40];
    46: op1_10_in18 = imem01_in[47:44];
    47: op1_10_in18 = reg_0610;
    48: op1_10_in18 = imem06_in[7:4];
    49: op1_10_in18 = reg_0803;
    50: op1_10_in18 = imem03_in[43:40];
    51: op1_10_in18 = imem01_in[19:16];
    52: op1_10_in18 = reg_0336;
    53: op1_10_in18 = reg_0527;
    54: op1_10_in18 = reg_0484;
    55: op1_10_in18 = reg_0289;
    56: op1_10_in18 = reg_0742;
    58: op1_10_in18 = imem07_in[103:100];
    59: op1_10_in18 = imem07_in[119:116];
    61: op1_10_in18 = imem01_in[3:0];
    63: op1_10_in18 = reg_0432;
    64: op1_10_in18 = imem05_in[111:108];
    65: op1_10_in18 = reg_0346;
    66: op1_10_in18 = reg_0103;
    67: op1_10_in18 = imem01_in[119:116];
    68: op1_10_in18 = reg_0739;
    69: op1_10_in18 = imem07_in[67:64];
    80: op1_10_in18 = imem07_in[67:64];
    71: op1_10_in18 = reg_0542;
    72: op1_10_in18 = imem07_in[79:76];
    75: op1_10_in18 = reg_0772;
    76: op1_10_in18 = reg_0414;
    77: op1_10_in18 = reg_0590;
    79: op1_10_in18 = reg_0818;
    81: op1_10_in18 = reg_0814;
    82: op1_10_in18 = reg_0530;
    83: op1_10_in18 = reg_0474;
    84: op1_10_in18 = imem06_in[23:20];
    86: op1_10_in18 = reg_0097;
    87: op1_10_in18 = reg_0257;
    88: op1_10_in18 = imem03_in[127:124];
    89: op1_10_in18 = reg_0583;
    90: op1_10_in18 = reg_0146;
    91: op1_10_in18 = reg_0636;
    92: op1_10_in18 = reg_0107;
    93: op1_10_in18 = reg_0197;
    94: op1_10_in18 = reg_0235;
    95: op1_10_in18 = reg_0498;
    default: op1_10_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv18 = 1;
    5: op1_10_inv18 = 1;
    6: op1_10_inv18 = 1;
    7: op1_10_inv18 = 1;
    11: op1_10_inv18 = 1;
    15: op1_10_inv18 = 1;
    16: op1_10_inv18 = 1;
    17: op1_10_inv18 = 1;
    18: op1_10_inv18 = 1;
    20: op1_10_inv18 = 1;
    21: op1_10_inv18 = 1;
    22: op1_10_inv18 = 1;
    23: op1_10_inv18 = 1;
    24: op1_10_inv18 = 1;
    27: op1_10_inv18 = 1;
    34: op1_10_inv18 = 1;
    42: op1_10_inv18 = 1;
    43: op1_10_inv18 = 1;
    44: op1_10_inv18 = 1;
    45: op1_10_inv18 = 1;
    49: op1_10_inv18 = 1;
    50: op1_10_inv18 = 1;
    51: op1_10_inv18 = 1;
    54: op1_10_inv18 = 1;
    55: op1_10_inv18 = 1;
    56: op1_10_inv18 = 1;
    57: op1_10_inv18 = 1;
    58: op1_10_inv18 = 1;
    59: op1_10_inv18 = 1;
    61: op1_10_inv18 = 1;
    62: op1_10_inv18 = 1;
    64: op1_10_inv18 = 1;
    66: op1_10_inv18 = 1;
    67: op1_10_inv18 = 1;
    75: op1_10_inv18 = 1;
    76: op1_10_inv18 = 1;
    77: op1_10_inv18 = 1;
    79: op1_10_inv18 = 1;
    81: op1_10_inv18 = 1;
    82: op1_10_inv18 = 1;
    84: op1_10_inv18 = 1;
    86: op1_10_inv18 = 1;
    87: op1_10_inv18 = 1;
    88: op1_10_inv18 = 1;
    89: op1_10_inv18 = 1;
    93: op1_10_inv18 = 1;
    95: op1_10_inv18 = 1;
    default: op1_10_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in19 = reg_0195;
    5: op1_10_in19 = reg_0201;
    6: op1_10_in19 = reg_0322;
    7: op1_10_in19 = reg_0621;
    8: op1_10_in19 = reg_0506;
    9: op1_10_in19 = imem07_in[7:4];
    10: op1_10_in19 = imem03_in[119:116];
    11: op1_10_in19 = reg_0429;
    12: op1_10_in19 = reg_0531;
    13: op1_10_in19 = reg_0131;
    14: op1_10_in19 = reg_0712;
    31: op1_10_in19 = reg_0712;
    15: op1_10_in19 = reg_0086;
    16: op1_10_in19 = reg_0074;
    17: op1_10_in19 = reg_0080;
    18: op1_10_in19 = reg_0058;
    19: op1_10_in19 = reg_0359;
    20: op1_10_in19 = reg_0494;
    21: op1_10_in19 = reg_0197;
    22: op1_10_in19 = reg_0776;
    23: op1_10_in19 = reg_0186;
    24: op1_10_in19 = reg_0092;
    25: op1_10_in19 = imem07_in[63:60];
    26: op1_10_in19 = reg_0556;
    27: op1_10_in19 = reg_0552;
    82: op1_10_in19 = reg_0552;
    28: op1_10_in19 = reg_0105;
    29: op1_10_in19 = reg_0647;
    30: op1_10_in19 = reg_0075;
    33: op1_10_in19 = reg_0098;
    34: op1_10_in19 = reg_0773;
    37: op1_10_in19 = reg_0773;
    35: op1_10_in19 = reg_0377;
    38: op1_10_in19 = imem01_in[35:32];
    39: op1_10_in19 = reg_0644;
    40: op1_10_in19 = reg_0314;
    41: op1_10_in19 = imem07_in[31:28];
    42: op1_10_in19 = reg_0159;
    43: op1_10_in19 = imem01_in[127:124];
    44: op1_10_in19 = reg_0780;
    45: op1_10_in19 = imem06_in[95:92];
    46: op1_10_in19 = imem01_in[83:80];
    47: op1_10_in19 = reg_0585;
    48: op1_10_in19 = imem06_in[23:20];
    49: op1_10_in19 = imem04_in[39:36];
    50: op1_10_in19 = imem03_in[47:44];
    51: op1_10_in19 = imem01_in[87:84];
    52: op1_10_in19 = reg_0341;
    53: op1_10_in19 = reg_0743;
    54: op1_10_in19 = reg_0495;
    55: op1_10_in19 = reg_0625;
    56: op1_10_in19 = reg_0070;
    57: op1_10_in19 = reg_0622;
    58: op1_10_in19 = imem07_in[119:116];
    59: op1_10_in19 = reg_0723;
    61: op1_10_in19 = imem01_in[15:12];
    62: op1_10_in19 = reg_0262;
    63: op1_10_in19 = reg_0305;
    64: op1_10_in19 = reg_0245;
    65: op1_10_in19 = reg_0408;
    66: op1_10_in19 = reg_0229;
    67: op1_10_in19 = imem01_in[123:120];
    68: op1_10_in19 = reg_0657;
    69: op1_10_in19 = reg_0716;
    71: op1_10_in19 = reg_0537;
    72: op1_10_in19 = imem07_in[83:80];
    73: op1_10_in19 = reg_0817;
    75: op1_10_in19 = reg_0102;
    76: op1_10_in19 = reg_0096;
    77: op1_10_in19 = reg_0343;
    78: op1_10_in19 = reg_0055;
    79: op1_10_in19 = reg_0752;
    80: op1_10_in19 = imem07_in[71:68];
    81: op1_10_in19 = reg_0339;
    83: op1_10_in19 = reg_0459;
    84: op1_10_in19 = imem06_in[63:60];
    86: op1_10_in19 = reg_0526;
    87: op1_10_in19 = reg_0761;
    88: op1_10_in19 = reg_0573;
    89: op1_10_in19 = reg_0491;
    90: op1_10_in19 = reg_0550;
    91: op1_10_in19 = reg_0051;
    92: op1_10_in19 = reg_0019;
    94: op1_10_in19 = reg_0019;
    93: op1_10_in19 = reg_0421;
    95: op1_10_in19 = reg_0123;
    default: op1_10_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv19 = 1;
    5: op1_10_inv19 = 1;
    6: op1_10_inv19 = 1;
    7: op1_10_inv19 = 1;
    9: op1_10_inv19 = 1;
    10: op1_10_inv19 = 1;
    13: op1_10_inv19 = 1;
    16: op1_10_inv19 = 1;
    18: op1_10_inv19 = 1;
    19: op1_10_inv19 = 1;
    23: op1_10_inv19 = 1;
    24: op1_10_inv19 = 1;
    28: op1_10_inv19 = 1;
    30: op1_10_inv19 = 1;
    33: op1_10_inv19 = 1;
    34: op1_10_inv19 = 1;
    37: op1_10_inv19 = 1;
    39: op1_10_inv19 = 1;
    43: op1_10_inv19 = 1;
    44: op1_10_inv19 = 1;
    45: op1_10_inv19 = 1;
    48: op1_10_inv19 = 1;
    49: op1_10_inv19 = 1;
    50: op1_10_inv19 = 1;
    51: op1_10_inv19 = 1;
    52: op1_10_inv19 = 1;
    53: op1_10_inv19 = 1;
    55: op1_10_inv19 = 1;
    62: op1_10_inv19 = 1;
    63: op1_10_inv19 = 1;
    67: op1_10_inv19 = 1;
    69: op1_10_inv19 = 1;
    72: op1_10_inv19 = 1;
    73: op1_10_inv19 = 1;
    81: op1_10_inv19 = 1;
    82: op1_10_inv19 = 1;
    89: op1_10_inv19 = 1;
    91: op1_10_inv19 = 1;
    92: op1_10_inv19 = 1;
    93: op1_10_inv19 = 1;
    default: op1_10_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in20 = imem01_in[51:48];
    5: op1_10_in20 = reg_0197;
    6: op1_10_in20 = reg_0374;
    7: op1_10_in20 = reg_0616;
    8: op1_10_in20 = reg_0508;
    9: op1_10_in20 = imem07_in[43:40];
    10: op1_10_in20 = reg_0569;
    11: op1_10_in20 = reg_0419;
    12: op1_10_in20 = reg_0303;
    13: op1_10_in20 = reg_0144;
    14: op1_10_in20 = reg_0708;
    15: op1_10_in20 = reg_0084;
    16: op1_10_in20 = imem05_in[19:16];
    17: op1_10_in20 = reg_0085;
    18: op1_10_in20 = reg_0552;
    19: op1_10_in20 = reg_0330;
    20: op1_10_in20 = reg_0486;
    21: op1_10_in20 = imem01_in[55:52];
    22: op1_10_in20 = reg_0241;
    23: op1_10_in20 = reg_0196;
    24: op1_10_in20 = reg_0540;
    25: op1_10_in20 = reg_0723;
    26: op1_10_in20 = reg_0273;
    27: op1_10_in20 = reg_0087;
    28: op1_10_in20 = reg_0103;
    29: op1_10_in20 = reg_0648;
    30: op1_10_in20 = imem05_in[7:4];
    31: op1_10_in20 = reg_0707;
    33: op1_10_in20 = reg_0498;
    34: op1_10_in20 = reg_0329;
    35: op1_10_in20 = reg_0319;
    37: op1_10_in20 = reg_0270;
    38: op1_10_in20 = reg_0336;
    39: op1_10_in20 = reg_0667;
    65: op1_10_in20 = reg_0667;
    40: op1_10_in20 = reg_0538;
    41: op1_10_in20 = imem07_in[119:116];
    42: op1_10_in20 = reg_0182;
    43: op1_10_in20 = reg_0501;
    44: op1_10_in20 = reg_0794;
    45: op1_10_in20 = imem06_in[103:100];
    46: op1_10_in20 = reg_0496;
    47: op1_10_in20 = reg_0640;
    48: op1_10_in20 = imem06_in[43:40];
    49: op1_10_in20 = imem04_in[55:52];
    50: op1_10_in20 = imem03_in[67:64];
    51: op1_10_in20 = imem01_in[91:88];
    52: op1_10_in20 = reg_0360;
    53: op1_10_in20 = reg_0740;
    54: op1_10_in20 = reg_0790;
    55: op1_10_in20 = reg_0606;
    56: op1_10_in20 = reg_0102;
    57: op1_10_in20 = reg_0311;
    58: op1_10_in20 = reg_0728;
    59: op1_10_in20 = reg_0726;
    69: op1_10_in20 = reg_0726;
    61: op1_10_in20 = imem01_in[35:32];
    62: op1_10_in20 = reg_0316;
    63: op1_10_in20 = reg_0615;
    64: op1_10_in20 = reg_0276;
    66: op1_10_in20 = reg_0249;
    67: op1_10_in20 = reg_0668;
    68: op1_10_in20 = reg_0483;
    71: op1_10_in20 = reg_0510;
    72: op1_10_in20 = imem07_in[87:84];
    80: op1_10_in20 = imem07_in[87:84];
    73: op1_10_in20 = reg_0619;
    75: op1_10_in20 = reg_0131;
    76: op1_10_in20 = reg_0756;
    77: op1_10_in20 = reg_0566;
    78: op1_10_in20 = reg_0558;
    79: op1_10_in20 = imem07_in[35:32];
    81: op1_10_in20 = reg_0773;
    82: op1_10_in20 = reg_0043;
    83: op1_10_in20 = reg_0191;
    84: op1_10_in20 = imem06_in[91:88];
    86: op1_10_in20 = imem03_in[15:12];
    87: op1_10_in20 = reg_0828;
    88: op1_10_in20 = reg_0801;
    89: op1_10_in20 = reg_0407;
    90: op1_10_in20 = reg_0793;
    91: op1_10_in20 = reg_0110;
    92: op1_10_in20 = reg_0188;
    93: op1_10_in20 = imem01_in[27:24];
    94: op1_10_in20 = reg_0645;
    95: op1_10_in20 = reg_0073;
    default: op1_10_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv20 = 1;
    5: op1_10_inv20 = 1;
    13: op1_10_inv20 = 1;
    18: op1_10_inv20 = 1;
    19: op1_10_inv20 = 1;
    22: op1_10_inv20 = 1;
    24: op1_10_inv20 = 1;
    25: op1_10_inv20 = 1;
    26: op1_10_inv20 = 1;
    27: op1_10_inv20 = 1;
    28: op1_10_inv20 = 1;
    29: op1_10_inv20 = 1;
    30: op1_10_inv20 = 1;
    33: op1_10_inv20 = 1;
    34: op1_10_inv20 = 1;
    35: op1_10_inv20 = 1;
    37: op1_10_inv20 = 1;
    38: op1_10_inv20 = 1;
    41: op1_10_inv20 = 1;
    44: op1_10_inv20 = 1;
    45: op1_10_inv20 = 1;
    46: op1_10_inv20 = 1;
    51: op1_10_inv20 = 1;
    52: op1_10_inv20 = 1;
    53: op1_10_inv20 = 1;
    57: op1_10_inv20 = 1;
    62: op1_10_inv20 = 1;
    64: op1_10_inv20 = 1;
    66: op1_10_inv20 = 1;
    67: op1_10_inv20 = 1;
    68: op1_10_inv20 = 1;
    72: op1_10_inv20 = 1;
    73: op1_10_inv20 = 1;
    76: op1_10_inv20 = 1;
    77: op1_10_inv20 = 1;
    78: op1_10_inv20 = 1;
    80: op1_10_inv20 = 1;
    81: op1_10_inv20 = 1;
    82: op1_10_inv20 = 1;
    83: op1_10_inv20 = 1;
    84: op1_10_inv20 = 1;
    86: op1_10_inv20 = 1;
    87: op1_10_inv20 = 1;
    88: op1_10_inv20 = 1;
    89: op1_10_inv20 = 1;
    91: op1_10_inv20 = 1;
    92: op1_10_inv20 = 1;
    94: op1_10_inv20 = 1;
    95: op1_10_inv20 = 1;
    default: op1_10_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in21 = imem01_in[91:88];
    5: op1_10_in21 = imem01_in[75:72];
    21: op1_10_in21 = imem01_in[75:72];
    6: op1_10_in21 = reg_0804;
    7: op1_10_in21 = reg_0626;
    8: op1_10_in21 = reg_0233;
    9: op1_10_in21 = imem07_in[51:48];
    10: op1_10_in21 = reg_0591;
    11: op1_10_in21 = reg_0437;
    12: op1_10_in21 = reg_0281;
    13: op1_10_in21 = imem06_in[19:16];
    14: op1_10_in21 = reg_0715;
    15: op1_10_in21 = reg_0087;
    16: op1_10_in21 = imem05_in[23:20];
    17: op1_10_in21 = reg_0086;
    18: op1_10_in21 = reg_0537;
    19: op1_10_in21 = reg_0346;
    20: op1_10_in21 = reg_0085;
    22: op1_10_in21 = reg_0218;
    23: op1_10_in21 = reg_0192;
    24: op1_10_in21 = imem03_in[27:24];
    25: op1_10_in21 = reg_0703;
    26: op1_10_in21 = reg_0290;
    27: op1_10_in21 = reg_0088;
    28: op1_10_in21 = reg_0111;
    29: op1_10_in21 = reg_0644;
    30: op1_10_in21 = imem05_in[43:40];
    31: op1_10_in21 = reg_0700;
    33: op1_10_in21 = reg_0093;
    34: op1_10_in21 = reg_0371;
    35: op1_10_in21 = reg_0338;
    37: op1_10_in21 = reg_0372;
    38: op1_10_in21 = reg_0520;
    43: op1_10_in21 = reg_0520;
    65: op1_10_in21 = reg_0520;
    39: op1_10_in21 = reg_0341;
    40: op1_10_in21 = imem03_in[3:0];
    41: op1_10_in21 = reg_0723;
    42: op1_10_in21 = reg_0164;
    44: op1_10_in21 = reg_0742;
    45: op1_10_in21 = imem06_in[115:112];
    46: op1_10_in21 = reg_0820;
    47: op1_10_in21 = reg_0255;
    48: op1_10_in21 = imem06_in[83:80];
    49: op1_10_in21 = imem04_in[87:84];
    50: op1_10_in21 = imem03_in[79:76];
    51: op1_10_in21 = reg_0735;
    52: op1_10_in21 = reg_0540;
    53: op1_10_in21 = reg_0063;
    54: op1_10_in21 = reg_0486;
    55: op1_10_in21 = reg_0608;
    56: op1_10_in21 = reg_0148;
    57: op1_10_in21 = reg_0289;
    84: op1_10_in21 = reg_0289;
    58: op1_10_in21 = reg_0702;
    59: op1_10_in21 = reg_0714;
    61: op1_10_in21 = imem01_in[39:36];
    62: op1_10_in21 = reg_0542;
    63: op1_10_in21 = reg_0431;
    64: op1_10_in21 = reg_0128;
    66: op1_10_in21 = reg_0783;
    67: op1_10_in21 = reg_0772;
    68: op1_10_in21 = reg_0753;
    69: op1_10_in21 = reg_0725;
    71: op1_10_in21 = reg_0429;
    72: op1_10_in21 = reg_0716;
    73: op1_10_in21 = reg_0031;
    75: op1_10_in21 = reg_0394;
    76: op1_10_in21 = reg_0526;
    77: op1_10_in21 = reg_0092;
    78: op1_10_in21 = reg_0510;
    79: op1_10_in21 = imem07_in[39:36];
    80: op1_10_in21 = imem07_in[99:96];
    81: op1_10_in21 = reg_0512;
    82: op1_10_in21 = reg_0083;
    83: op1_10_in21 = reg_0187;
    86: op1_10_in21 = imem03_in[55:52];
    87: op1_10_in21 = reg_0734;
    88: op1_10_in21 = reg_0015;
    89: op1_10_in21 = reg_0285;
    90: op1_10_in21 = reg_0090;
    91: op1_10_in21 = reg_0228;
    92: op1_10_in21 = reg_0225;
    93: op1_10_in21 = imem01_in[31:28];
    94: op1_10_in21 = reg_0217;
    95: op1_10_in21 = reg_0125;
    default: op1_10_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv21 = 1;
    6: op1_10_inv21 = 1;
    8: op1_10_inv21 = 1;
    12: op1_10_inv21 = 1;
    13: op1_10_inv21 = 1;
    14: op1_10_inv21 = 1;
    15: op1_10_inv21 = 1;
    17: op1_10_inv21 = 1;
    18: op1_10_inv21 = 1;
    19: op1_10_inv21 = 1;
    20: op1_10_inv21 = 1;
    21: op1_10_inv21 = 1;
    22: op1_10_inv21 = 1;
    26: op1_10_inv21 = 1;
    28: op1_10_inv21 = 1;
    30: op1_10_inv21 = 1;
    31: op1_10_inv21 = 1;
    33: op1_10_inv21 = 1;
    34: op1_10_inv21 = 1;
    38: op1_10_inv21 = 1;
    40: op1_10_inv21 = 1;
    41: op1_10_inv21 = 1;
    43: op1_10_inv21 = 1;
    44: op1_10_inv21 = 1;
    46: op1_10_inv21 = 1;
    48: op1_10_inv21 = 1;
    49: op1_10_inv21 = 1;
    50: op1_10_inv21 = 1;
    55: op1_10_inv21 = 1;
    56: op1_10_inv21 = 1;
    57: op1_10_inv21 = 1;
    58: op1_10_inv21 = 1;
    62: op1_10_inv21 = 1;
    64: op1_10_inv21 = 1;
    66: op1_10_inv21 = 1;
    67: op1_10_inv21 = 1;
    68: op1_10_inv21 = 1;
    69: op1_10_inv21 = 1;
    71: op1_10_inv21 = 1;
    72: op1_10_inv21 = 1;
    78: op1_10_inv21 = 1;
    80: op1_10_inv21 = 1;
    83: op1_10_inv21 = 1;
    87: op1_10_inv21 = 1;
    89: op1_10_inv21 = 1;
    92: op1_10_inv21 = 1;
    95: op1_10_inv21 = 1;
    default: op1_10_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in22 = imem01_in[95:92];
    5: op1_10_in22 = imem01_in[87:84];
    6: op1_10_in22 = reg_0802;
    7: op1_10_in22 = reg_0618;
    8: op1_10_in22 = reg_0242;
    9: op1_10_in22 = imem07_in[75:72];
    10: op1_10_in22 = reg_0584;
    11: op1_10_in22 = reg_0158;
    12: op1_10_in22 = reg_0305;
    13: op1_10_in22 = imem06_in[47:44];
    14: op1_10_in22 = reg_0706;
    15: op1_10_in22 = reg_0094;
    16: op1_10_in22 = imem05_in[59:56];
    17: op1_10_in22 = imem03_in[31:28];
    18: op1_10_in22 = imem04_in[19:16];
    19: op1_10_in22 = reg_0324;
    20: op1_10_in22 = reg_0147;
    21: op1_10_in22 = imem01_in[91:88];
    22: op1_10_in22 = reg_0249;
    23: op1_10_in22 = imem01_in[47:44];
    93: op1_10_in22 = imem01_in[47:44];
    24: op1_10_in22 = imem03_in[43:40];
    25: op1_10_in22 = reg_0712;
    58: op1_10_in22 = reg_0712;
    26: op1_10_in22 = reg_0291;
    57: op1_10_in22 = reg_0291;
    27: op1_10_in22 = reg_0510;
    28: op1_10_in22 = reg_0112;
    29: op1_10_in22 = reg_0354;
    53: op1_10_in22 = reg_0354;
    30: op1_10_in22 = imem05_in[63:60];
    31: op1_10_in22 = reg_0429;
    78: op1_10_in22 = reg_0429;
    33: op1_10_in22 = imem03_in[35:32];
    34: op1_10_in22 = reg_0368;
    35: op1_10_in22 = reg_0368;
    37: op1_10_in22 = reg_0338;
    38: op1_10_in22 = reg_0824;
    39: op1_10_in22 = reg_0355;
    40: op1_10_in22 = imem03_in[23:20];
    76: op1_10_in22 = imem03_in[23:20];
    41: op1_10_in22 = reg_0708;
    42: op1_10_in22 = reg_0170;
    43: op1_10_in22 = reg_0822;
    44: op1_10_in22 = reg_0226;
    45: op1_10_in22 = reg_0247;
    46: op1_10_in22 = reg_0825;
    47: op1_10_in22 = reg_0643;
    48: op1_10_in22 = reg_0416;
    49: op1_10_in22 = imem04_in[95:92];
    50: op1_10_in22 = imem03_in[83:80];
    51: op1_10_in22 = reg_0085;
    52: op1_10_in22 = reg_0757;
    54: op1_10_in22 = reg_0309;
    55: op1_10_in22 = reg_0766;
    56: op1_10_in22 = reg_0151;
    59: op1_10_in22 = reg_0703;
    61: op1_10_in22 = imem01_in[55:52];
    62: op1_10_in22 = reg_0523;
    63: op1_10_in22 = reg_0508;
    71: op1_10_in22 = reg_0508;
    64: op1_10_in22 = reg_0129;
    65: op1_10_in22 = reg_0812;
    66: op1_10_in22 = reg_0790;
    67: op1_10_in22 = reg_0765;
    68: op1_10_in22 = reg_0484;
    69: op1_10_in22 = reg_0702;
    72: op1_10_in22 = reg_0729;
    73: op1_10_in22 = reg_0773;
    75: op1_10_in22 = reg_0759;
    77: op1_10_in22 = reg_0540;
    79: op1_10_in22 = imem07_in[47:44];
    80: op1_10_in22 = imem07_in[107:104];
    81: op1_10_in22 = reg_0573;
    82: op1_10_in22 = reg_0086;
    83: op1_10_in22 = reg_0204;
    84: op1_10_in22 = reg_0624;
    86: op1_10_in22 = imem03_in[67:64];
    87: op1_10_in22 = imem06_in[19:16];
    88: op1_10_in22 = reg_0589;
    89: op1_10_in22 = reg_0149;
    90: op1_10_in22 = reg_0027;
    91: op1_10_in22 = reg_0185;
    92: op1_10_in22 = reg_0497;
    94: op1_10_in22 = reg_0518;
    95: op1_10_in22 = reg_0670;
    default: op1_10_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv22 = 1;
    6: op1_10_inv22 = 1;
    7: op1_10_inv22 = 1;
    9: op1_10_inv22 = 1;
    12: op1_10_inv22 = 1;
    13: op1_10_inv22 = 1;
    15: op1_10_inv22 = 1;
    17: op1_10_inv22 = 1;
    18: op1_10_inv22 = 1;
    19: op1_10_inv22 = 1;
    21: op1_10_inv22 = 1;
    23: op1_10_inv22 = 1;
    24: op1_10_inv22 = 1;
    28: op1_10_inv22 = 1;
    29: op1_10_inv22 = 1;
    30: op1_10_inv22 = 1;
    33: op1_10_inv22 = 1;
    34: op1_10_inv22 = 1;
    37: op1_10_inv22 = 1;
    38: op1_10_inv22 = 1;
    39: op1_10_inv22 = 1;
    41: op1_10_inv22 = 1;
    43: op1_10_inv22 = 1;
    44: op1_10_inv22 = 1;
    45: op1_10_inv22 = 1;
    49: op1_10_inv22 = 1;
    58: op1_10_inv22 = 1;
    59: op1_10_inv22 = 1;
    64: op1_10_inv22 = 1;
    65: op1_10_inv22 = 1;
    67: op1_10_inv22 = 1;
    69: op1_10_inv22 = 1;
    71: op1_10_inv22 = 1;
    72: op1_10_inv22 = 1;
    75: op1_10_inv22 = 1;
    77: op1_10_inv22 = 1;
    78: op1_10_inv22 = 1;
    80: op1_10_inv22 = 1;
    81: op1_10_inv22 = 1;
    82: op1_10_inv22 = 1;
    84: op1_10_inv22 = 1;
    88: op1_10_inv22 = 1;
    89: op1_10_inv22 = 1;
    90: op1_10_inv22 = 1;
    95: op1_10_inv22 = 1;
    default: op1_10_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in23 = imem01_in[111:108];
    5: op1_10_in23 = imem01_in[123:120];
    6: op1_10_in23 = reg_0799;
    7: op1_10_in23 = reg_0402;
    8: op1_10_in23 = reg_0247;
    9: op1_10_in23 = imem07_in[119:116];
    10: op1_10_in23 = reg_0580;
    12: op1_10_in23 = reg_0277;
    13: op1_10_in23 = imem06_in[67:64];
    14: op1_10_in23 = reg_0422;
    15: op1_10_in23 = reg_0079;
    16: op1_10_in23 = imem05_in[107:104];
    17: op1_10_in23 = imem03_in[35:32];
    40: op1_10_in23 = imem03_in[35:32];
    18: op1_10_in23 = imem04_in[87:84];
    19: op1_10_in23 = reg_0365;
    20: op1_10_in23 = reg_0148;
    21: op1_10_in23 = imem01_in[95:92];
    22: op1_10_in23 = reg_0104;
    23: op1_10_in23 = imem01_in[99:96];
    24: op1_10_in23 = imem03_in[75:72];
    25: op1_10_in23 = reg_0729;
    26: op1_10_in23 = reg_0295;
    27: op1_10_in23 = reg_0516;
    28: op1_10_in23 = reg_0114;
    29: op1_10_in23 = reg_0341;
    30: op1_10_in23 = imem05_in[75:72];
    31: op1_10_in23 = reg_0432;
    33: op1_10_in23 = imem03_in[39:36];
    34: op1_10_in23 = reg_0818;
    35: op1_10_in23 = reg_0375;
    37: op1_10_in23 = imem07_in[3:0];
    38: op1_10_in23 = reg_0563;
    39: op1_10_in23 = reg_0347;
    41: op1_10_in23 = reg_0709;
    42: op1_10_in23 = reg_0157;
    43: op1_10_in23 = reg_0337;
    44: op1_10_in23 = reg_0269;
    45: op1_10_in23 = reg_0618;
    46: op1_10_in23 = reg_0760;
    47: op1_10_in23 = imem05_in[59:56];
    48: op1_10_in23 = reg_0609;
    49: op1_10_in23 = imem04_in[119:116];
    50: op1_10_in23 = imem03_in[103:100];
    51: op1_10_in23 = reg_0668;
    52: op1_10_in23 = imem03_in[3:0];
    53: op1_10_in23 = reg_0401;
    54: op1_10_in23 = reg_0226;
    55: op1_10_in23 = reg_0763;
    56: op1_10_in23 = reg_0142;
    57: op1_10_in23 = reg_0577;
    58: op1_10_in23 = reg_0724;
    59: op1_10_in23 = reg_0724;
    61: op1_10_in23 = reg_0761;
    62: op1_10_in23 = reg_0547;
    63: op1_10_in23 = reg_0301;
    64: op1_10_in23 = reg_0130;
    65: op1_10_in23 = reg_0218;
    66: op1_10_in23 = reg_0236;
    67: op1_10_in23 = reg_0778;
    68: op1_10_in23 = reg_0655;
    69: op1_10_in23 = reg_0703;
    71: op1_10_in23 = reg_0679;
    72: op1_10_in23 = reg_0715;
    73: op1_10_in23 = reg_0638;
    75: op1_10_in23 = reg_0388;
    76: op1_10_in23 = imem03_in[31:28];
    77: op1_10_in23 = reg_0756;
    78: op1_10_in23 = reg_0631;
    79: op1_10_in23 = imem07_in[71:68];
    80: op1_10_in23 = imem07_in[115:112];
    81: op1_10_in23 = reg_0039;
    82: op1_10_in23 = reg_0057;
    83: op1_10_in23 = reg_0194;
    84: op1_10_in23 = reg_0762;
    86: op1_10_in23 = imem03_in[99:96];
    87: op1_10_in23 = imem06_in[35:32];
    88: op1_10_in23 = reg_0010;
    89: op1_10_in23 = reg_0827;
    90: op1_10_in23 = reg_0144;
    92: op1_10_in23 = reg_0759;
    93: op1_10_in23 = imem01_in[79:76];
    94: op1_10_in23 = reg_0419;
    95: op1_10_in23 = reg_0675;
    default: op1_10_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv23 = 1;
    5: op1_10_inv23 = 1;
    7: op1_10_inv23 = 1;
    8: op1_10_inv23 = 1;
    12: op1_10_inv23 = 1;
    13: op1_10_inv23 = 1;
    14: op1_10_inv23 = 1;
    18: op1_10_inv23 = 1;
    22: op1_10_inv23 = 1;
    25: op1_10_inv23 = 1;
    26: op1_10_inv23 = 1;
    27: op1_10_inv23 = 1;
    29: op1_10_inv23 = 1;
    30: op1_10_inv23 = 1;
    31: op1_10_inv23 = 1;
    34: op1_10_inv23 = 1;
    40: op1_10_inv23 = 1;
    42: op1_10_inv23 = 1;
    45: op1_10_inv23 = 1;
    46: op1_10_inv23 = 1;
    50: op1_10_inv23 = 1;
    52: op1_10_inv23 = 1;
    53: op1_10_inv23 = 1;
    55: op1_10_inv23 = 1;
    58: op1_10_inv23 = 1;
    59: op1_10_inv23 = 1;
    62: op1_10_inv23 = 1;
    63: op1_10_inv23 = 1;
    66: op1_10_inv23 = 1;
    69: op1_10_inv23 = 1;
    71: op1_10_inv23 = 1;
    72: op1_10_inv23 = 1;
    73: op1_10_inv23 = 1;
    79: op1_10_inv23 = 1;
    82: op1_10_inv23 = 1;
    83: op1_10_inv23 = 1;
    84: op1_10_inv23 = 1;
    86: op1_10_inv23 = 1;
    87: op1_10_inv23 = 1;
    88: op1_10_inv23 = 1;
    89: op1_10_inv23 = 1;
    92: op1_10_inv23 = 1;
    93: op1_10_inv23 = 1;
    94: op1_10_inv23 = 1;
    default: op1_10_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in24 = reg_0503;
    5: op1_10_in24 = imem01_in[127:124];
    6: op1_10_in24 = imem04_in[3:0];
    7: op1_10_in24 = reg_0356;
    8: op1_10_in24 = reg_0236;
    9: op1_10_in24 = reg_0704;
    10: op1_10_in24 = reg_0576;
    12: op1_10_in24 = reg_0276;
    13: op1_10_in24 = reg_0611;
    14: op1_10_in24 = reg_0433;
    15: op1_10_in24 = imem03_in[11:8];
    16: op1_10_in24 = imem05_in[111:108];
    17: op1_10_in24 = imem03_in[83:80];
    18: op1_10_in24 = imem04_in[99:96];
    19: op1_10_in24 = reg_0355;
    68: op1_10_in24 = reg_0355;
    20: op1_10_in24 = reg_0136;
    21: op1_10_in24 = imem01_in[111:108];
    22: op1_10_in24 = reg_0120;
    23: op1_10_in24 = imem01_in[107:104];
    24: op1_10_in24 = imem03_in[99:96];
    25: op1_10_in24 = reg_0713;
    58: op1_10_in24 = reg_0713;
    26: op1_10_in24 = reg_0298;
    27: op1_10_in24 = reg_0556;
    28: op1_10_in24 = reg_0100;
    29: op1_10_in24 = reg_0361;
    30: op1_10_in24 = imem05_in[119:116];
    31: op1_10_in24 = reg_0436;
    33: op1_10_in24 = imem03_in[59:56];
    34: op1_10_in24 = reg_0605;
    35: op1_10_in24 = imem07_in[11:8];
    37: op1_10_in24 = imem07_in[71:68];
    38: op1_10_in24 = reg_0487;
    39: op1_10_in24 = reg_0092;
    40: op1_10_in24 = imem03_in[51:48];
    41: op1_10_in24 = reg_0441;
    43: op1_10_in24 = reg_0519;
    44: op1_10_in24 = reg_0277;
    45: op1_10_in24 = reg_0405;
    46: op1_10_in24 = reg_0241;
    47: op1_10_in24 = imem05_in[63:60];
    48: op1_10_in24 = reg_0293;
    49: op1_10_in24 = reg_0262;
    50: op1_10_in24 = imem03_in[107:104];
    51: op1_10_in24 = reg_0496;
    52: op1_10_in24 = imem03_in[47:44];
    53: op1_10_in24 = reg_0311;
    54: op1_10_in24 = reg_0307;
    55: op1_10_in24 = reg_0776;
    56: op1_10_in24 = reg_0146;
    57: op1_10_in24 = reg_0409;
    59: op1_10_in24 = reg_0708;
    61: op1_10_in24 = reg_0649;
    62: op1_10_in24 = reg_0429;
    63: op1_10_in24 = reg_0640;
    64: op1_10_in24 = reg_0140;
    65: op1_10_in24 = reg_0787;
    66: op1_10_in24 = reg_0142;
    67: op1_10_in24 = reg_0737;
    69: op1_10_in24 = reg_0724;
    71: op1_10_in24 = reg_0062;
    72: op1_10_in24 = reg_0711;
    73: op1_10_in24 = reg_0039;
    75: op1_10_in24 = reg_0225;
    76: op1_10_in24 = imem03_in[55:52];
    77: op1_10_in24 = reg_0531;
    78: op1_10_in24 = reg_0431;
    79: op1_10_in24 = imem07_in[99:96];
    81: op1_10_in24 = reg_0322;
    82: op1_10_in24 = reg_0075;
    83: op1_10_in24 = reg_0196;
    84: op1_10_in24 = reg_0404;
    86: op1_10_in24 = reg_0589;
    87: op1_10_in24 = imem06_in[71:68];
    88: op1_10_in24 = reg_0595;
    89: op1_10_in24 = reg_0152;
    90: op1_10_in24 = reg_0797;
    92: op1_10_in24 = reg_0397;
    93: op1_10_in24 = imem01_in[103:100];
    94: op1_10_in24 = imem01_in[19:16];
    95: op1_10_in24 = reg_0671;
    default: op1_10_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv24 = 1;
    5: op1_10_inv24 = 1;
    6: op1_10_inv24 = 1;
    7: op1_10_inv24 = 1;
    9: op1_10_inv24 = 1;
    10: op1_10_inv24 = 1;
    13: op1_10_inv24 = 1;
    14: op1_10_inv24 = 1;
    15: op1_10_inv24 = 1;
    17: op1_10_inv24 = 1;
    20: op1_10_inv24 = 1;
    21: op1_10_inv24 = 1;
    22: op1_10_inv24 = 1;
    23: op1_10_inv24 = 1;
    26: op1_10_inv24 = 1;
    27: op1_10_inv24 = 1;
    30: op1_10_inv24 = 1;
    31: op1_10_inv24 = 1;
    35: op1_10_inv24 = 1;
    39: op1_10_inv24 = 1;
    41: op1_10_inv24 = 1;
    45: op1_10_inv24 = 1;
    46: op1_10_inv24 = 1;
    49: op1_10_inv24 = 1;
    52: op1_10_inv24 = 1;
    54: op1_10_inv24 = 1;
    55: op1_10_inv24 = 1;
    56: op1_10_inv24 = 1;
    57: op1_10_inv24 = 1;
    59: op1_10_inv24 = 1;
    61: op1_10_inv24 = 1;
    62: op1_10_inv24 = 1;
    64: op1_10_inv24 = 1;
    65: op1_10_inv24 = 1;
    66: op1_10_inv24 = 1;
    67: op1_10_inv24 = 1;
    71: op1_10_inv24 = 1;
    77: op1_10_inv24 = 1;
    79: op1_10_inv24 = 1;
    82: op1_10_inv24 = 1;
    83: op1_10_inv24 = 1;
    84: op1_10_inv24 = 1;
    86: op1_10_inv24 = 1;
    90: op1_10_inv24 = 1;
    93: op1_10_inv24 = 1;
    94: op1_10_inv24 = 1;
    default: op1_10_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in25 = reg_0517;
    5: op1_10_in25 = reg_0520;
    6: op1_10_in25 = imem04_in[71:68];
    7: op1_10_in25 = reg_0407;
    8: op1_10_in25 = reg_0248;
    9: op1_10_in25 = reg_0712;
    10: op1_10_in25 = reg_0394;
    12: op1_10_in25 = reg_0291;
    13: op1_10_in25 = reg_0577;
    14: op1_10_in25 = reg_0423;
    31: op1_10_in25 = reg_0423;
    15: op1_10_in25 = imem03_in[31:28];
    16: op1_10_in25 = reg_0798;
    17: op1_10_in25 = imem03_in[103:100];
    40: op1_10_in25 = imem03_in[103:100];
    18: op1_10_in25 = reg_0257;
    89: op1_10_in25 = reg_0257;
    19: op1_10_in25 = reg_0314;
    20: op1_10_in25 = reg_0152;
    21: op1_10_in25 = imem01_in[127:124];
    22: op1_10_in25 = reg_0126;
    23: op1_10_in25 = imem01_in[123:120];
    24: op1_10_in25 = imem03_in[115:112];
    25: op1_10_in25 = reg_0425;
    26: op1_10_in25 = reg_0253;
    58: op1_10_in25 = reg_0253;
    27: op1_10_in25 = reg_0301;
    28: op1_10_in25 = reg_0106;
    29: op1_10_in25 = reg_0363;
    30: op1_10_in25 = reg_0495;
    33: op1_10_in25 = imem03_in[91:88];
    34: op1_10_in25 = reg_0766;
    35: op1_10_in25 = imem07_in[31:28];
    37: op1_10_in25 = imem07_in[99:96];
    38: op1_10_in25 = reg_0235;
    43: op1_10_in25 = reg_0235;
    39: op1_10_in25 = reg_0769;
    41: op1_10_in25 = reg_0447;
    44: op1_10_in25 = reg_0734;
    45: op1_10_in25 = reg_0775;
    46: op1_10_in25 = reg_0504;
    47: op1_10_in25 = imem05_in[75:72];
    48: op1_10_in25 = reg_0265;
    49: op1_10_in25 = reg_0316;
    50: op1_10_in25 = reg_0601;
    51: op1_10_in25 = reg_0820;
    52: op1_10_in25 = reg_0579;
    53: op1_10_in25 = imem03_in[3:0];
    54: op1_10_in25 = reg_0136;
    55: op1_10_in25 = reg_0404;
    56: op1_10_in25 = reg_0156;
    57: op1_10_in25 = reg_0238;
    59: op1_10_in25 = reg_0718;
    61: op1_10_in25 = reg_0237;
    62: op1_10_in25 = reg_0071;
    63: op1_10_in25 = reg_0776;
    64: op1_10_in25 = reg_0134;
    65: op1_10_in25 = reg_0029;
    66: op1_10_in25 = reg_0146;
    67: op1_10_in25 = reg_0502;
    68: op1_10_in25 = reg_0372;
    69: op1_10_in25 = reg_0708;
    71: op1_10_in25 = reg_0644;
    72: op1_10_in25 = reg_0727;
    73: op1_10_in25 = reg_0025;
    75: op1_10_in25 = reg_0574;
    76: op1_10_in25 = reg_0602;
    77: op1_10_in25 = reg_0498;
    78: op1_10_in25 = reg_0050;
    79: op1_10_in25 = reg_0721;
    81: op1_10_in25 = reg_0777;
    82: op1_10_in25 = reg_0533;
    83: op1_10_in25 = reg_0205;
    84: op1_10_in25 = reg_0618;
    86: op1_10_in25 = reg_0604;
    87: op1_10_in25 = imem06_in[75:72];
    88: op1_10_in25 = reg_0486;
    90: op1_10_in25 = reg_0583;
    92: op1_10_in25 = imem01_in[51:48];
    93: op1_10_in25 = reg_0085;
    94: op1_10_in25 = imem01_in[63:60];
    95: op1_10_in25 = reg_0674;
    default: op1_10_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv25 = 1;
    8: op1_10_inv25 = 1;
    9: op1_10_inv25 = 1;
    10: op1_10_inv25 = 1;
    12: op1_10_inv25 = 1;
    13: op1_10_inv25 = 1;
    14: op1_10_inv25 = 1;
    15: op1_10_inv25 = 1;
    16: op1_10_inv25 = 1;
    17: op1_10_inv25 = 1;
    19: op1_10_inv25 = 1;
    22: op1_10_inv25 = 1;
    23: op1_10_inv25 = 1;
    26: op1_10_inv25 = 1;
    28: op1_10_inv25 = 1;
    30: op1_10_inv25 = 1;
    33: op1_10_inv25 = 1;
    35: op1_10_inv25 = 1;
    37: op1_10_inv25 = 1;
    39: op1_10_inv25 = 1;
    41: op1_10_inv25 = 1;
    44: op1_10_inv25 = 1;
    45: op1_10_inv25 = 1;
    46: op1_10_inv25 = 1;
    54: op1_10_inv25 = 1;
    55: op1_10_inv25 = 1;
    58: op1_10_inv25 = 1;
    61: op1_10_inv25 = 1;
    62: op1_10_inv25 = 1;
    63: op1_10_inv25 = 1;
    65: op1_10_inv25 = 1;
    66: op1_10_inv25 = 1;
    67: op1_10_inv25 = 1;
    69: op1_10_inv25 = 1;
    71: op1_10_inv25 = 1;
    72: op1_10_inv25 = 1;
    76: op1_10_inv25 = 1;
    78: op1_10_inv25 = 1;
    82: op1_10_inv25 = 1;
    83: op1_10_inv25 = 1;
    89: op1_10_inv25 = 1;
    92: op1_10_inv25 = 1;
    93: op1_10_inv25 = 1;
    94: op1_10_inv25 = 1;
    default: op1_10_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in26 = reg_0518;
    5: op1_10_in26 = reg_0521;
    6: op1_10_in26 = imem04_in[75:72];
    7: op1_10_in26 = reg_0405;
    8: op1_10_in26 = reg_0234;
    9: op1_10_in26 = reg_0729;
    10: op1_10_in26 = reg_0360;
    12: op1_10_in26 = reg_0297;
    13: op1_10_in26 = reg_0615;
    14: op1_10_in26 = reg_0439;
    15: op1_10_in26 = imem03_in[43:40];
    16: op1_10_in26 = reg_0781;
    17: op1_10_in26 = reg_0602;
    18: op1_10_in26 = reg_0078;
    19: op1_10_in26 = reg_0092;
    20: op1_10_in26 = imem06_in[79:76];
    21: op1_10_in26 = reg_0497;
    22: op1_10_in26 = imem02_in[27:24];
    23: op1_10_in26 = reg_0512;
    24: op1_10_in26 = reg_0598;
    40: op1_10_in26 = reg_0598;
    25: op1_10_in26 = reg_0441;
    26: op1_10_in26 = reg_0299;
    27: op1_10_in26 = reg_0052;
    28: op1_10_in26 = reg_0101;
    29: op1_10_in26 = reg_0346;
    30: op1_10_in26 = reg_0790;
    31: op1_10_in26 = reg_0448;
    33: op1_10_in26 = imem03_in[107:104];
    34: op1_10_in26 = imem07_in[11:8];
    35: op1_10_in26 = imem07_in[43:40];
    37: op1_10_in26 = imem07_in[111:108];
    38: op1_10_in26 = reg_0240;
    39: op1_10_in26 = reg_0535;
    41: op1_10_in26 = reg_0434;
    43: op1_10_in26 = reg_0574;
    44: op1_10_in26 = reg_0147;
    45: op1_10_in26 = reg_0763;
    46: op1_10_in26 = reg_0116;
    47: op1_10_in26 = imem05_in[95:92];
    48: op1_10_in26 = reg_0025;
    49: op1_10_in26 = reg_0552;
    50: op1_10_in26 = reg_0599;
    76: op1_10_in26 = reg_0599;
    51: op1_10_in26 = reg_0322;
    52: op1_10_in26 = reg_0589;
    53: op1_10_in26 = imem03_in[7:4];
    54: op1_10_in26 = reg_0144;
    55: op1_10_in26 = reg_0038;
    56: op1_10_in26 = reg_0062;
    57: op1_10_in26 = reg_0404;
    58: op1_10_in26 = reg_0266;
    59: op1_10_in26 = reg_0706;
    61: op1_10_in26 = reg_0760;
    62: op1_10_in26 = reg_0629;
    63: op1_10_in26 = imem05_in[7:4];
    64: op1_10_in26 = imem06_in[15:12];
    65: op1_10_in26 = imem07_in[3:0];
    66: op1_10_in26 = reg_0138;
    67: op1_10_in26 = reg_0216;
    68: op1_10_in26 = reg_0356;
    69: op1_10_in26 = reg_0635;
    71: op1_10_in26 = reg_0109;
    72: op1_10_in26 = reg_0067;
    73: op1_10_in26 = reg_0794;
    75: op1_10_in26 = reg_0220;
    77: op1_10_in26 = imem03_in[11:8];
    78: op1_10_in26 = reg_0679;
    79: op1_10_in26 = reg_0163;
    81: op1_10_in26 = reg_0818;
    82: op1_10_in26 = reg_0547;
    83: op1_10_in26 = reg_0197;
    84: op1_10_in26 = reg_0260;
    86: op1_10_in26 = reg_0493;
    87: op1_10_in26 = reg_0289;
    88: op1_10_in26 = reg_0648;
    89: op1_10_in26 = reg_0796;
    90: op1_10_in26 = reg_0252;
    92: op1_10_in26 = imem01_in[95:92];
    94: op1_10_in26 = imem01_in[95:92];
    93: op1_10_in26 = reg_0007;
    95: op1_10_in26 = reg_0121;
    default: op1_10_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_10_inv26 = 1;
    7: op1_10_inv26 = 1;
    8: op1_10_inv26 = 1;
    12: op1_10_inv26 = 1;
    13: op1_10_inv26 = 1;
    15: op1_10_inv26 = 1;
    17: op1_10_inv26 = 1;
    18: op1_10_inv26 = 1;
    21: op1_10_inv26 = 1;
    22: op1_10_inv26 = 1;
    23: op1_10_inv26 = 1;
    24: op1_10_inv26 = 1;
    26: op1_10_inv26 = 1;
    31: op1_10_inv26 = 1;
    33: op1_10_inv26 = 1;
    34: op1_10_inv26 = 1;
    37: op1_10_inv26 = 1;
    39: op1_10_inv26 = 1;
    43: op1_10_inv26 = 1;
    44: op1_10_inv26 = 1;
    45: op1_10_inv26 = 1;
    50: op1_10_inv26 = 1;
    51: op1_10_inv26 = 1;
    52: op1_10_inv26 = 1;
    53: op1_10_inv26 = 1;
    54: op1_10_inv26 = 1;
    56: op1_10_inv26 = 1;
    61: op1_10_inv26 = 1;
    64: op1_10_inv26 = 1;
    65: op1_10_inv26 = 1;
    66: op1_10_inv26 = 1;
    69: op1_10_inv26 = 1;
    71: op1_10_inv26 = 1;
    72: op1_10_inv26 = 1;
    75: op1_10_inv26 = 1;
    76: op1_10_inv26 = 1;
    81: op1_10_inv26 = 1;
    83: op1_10_inv26 = 1;
    87: op1_10_inv26 = 1;
    90: op1_10_inv26 = 1;
    92: op1_10_inv26 = 1;
    93: op1_10_inv26 = 1;
    default: op1_10_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in27 = reg_0506;
    5: op1_10_in27 = reg_0499;
    6: op1_10_in27 = imem04_in[79:76];
    7: op1_10_in27 = reg_0406;
    8: op1_10_in27 = reg_0245;
    9: op1_10_in27 = reg_0709;
    10: op1_10_in27 = reg_0343;
    29: op1_10_in27 = reg_0343;
    12: op1_10_in27 = reg_0298;
    13: op1_10_in27 = reg_0348;
    14: op1_10_in27 = reg_0446;
    15: op1_10_in27 = imem03_in[51:48];
    16: op1_10_in27 = reg_0490;
    17: op1_10_in27 = reg_0572;
    18: op1_10_in27 = reg_0299;
    19: op1_10_in27 = reg_0095;
    20: op1_10_in27 = imem06_in[127:124];
    21: op1_10_in27 = reg_0227;
    22: op1_10_in27 = imem02_in[91:88];
    23: op1_10_in27 = reg_0514;
    24: op1_10_in27 = reg_0571;
    25: op1_10_in27 = reg_0422;
    26: op1_10_in27 = reg_0289;
    27: op1_10_in27 = reg_0274;
    28: op1_10_in27 = reg_0115;
    30: op1_10_in27 = reg_0489;
    31: op1_10_in27 = reg_0431;
    33: op1_10_in27 = reg_0586;
    34: op1_10_in27 = imem07_in[63:60];
    35: op1_10_in27 = imem07_in[59:56];
    37: op1_10_in27 = imem07_in[115:112];
    38: op1_10_in27 = reg_0504;
    39: op1_10_in27 = reg_0094;
    40: op1_10_in27 = reg_0601;
    41: op1_10_in27 = reg_0440;
    43: op1_10_in27 = reg_0603;
    44: op1_10_in27 = reg_0136;
    45: op1_10_in27 = reg_0403;
    46: op1_10_in27 = reg_0104;
    47: op1_10_in27 = reg_0491;
    90: op1_10_in27 = reg_0491;
    48: op1_10_in27 = reg_0369;
    56: op1_10_in27 = reg_0369;
    49: op1_10_in27 = reg_0542;
    50: op1_10_in27 = reg_0579;
    76: op1_10_in27 = reg_0579;
    51: op1_10_in27 = reg_0734;
    52: op1_10_in27 = reg_0384;
    53: op1_10_in27 = imem03_in[23:20];
    54: op1_10_in27 = imem06_in[7:4];
    55: op1_10_in27 = reg_0368;
    57: op1_10_in27 = reg_0339;
    58: op1_10_in27 = reg_0436;
    59: op1_10_in27 = reg_0700;
    61: op1_10_in27 = reg_0232;
    62: op1_10_in27 = reg_0050;
    63: op1_10_in27 = imem05_in[39:36];
    64: op1_10_in27 = imem06_in[47:44];
    65: op1_10_in27 = imem07_in[7:4];
    66: op1_10_in27 = reg_0153;
    67: op1_10_in27 = reg_0290;
    68: op1_10_in27 = reg_0363;
    69: op1_10_in27 = reg_0439;
    71: op1_10_in27 = imem05_in[7:4];
    72: op1_10_in27 = reg_0239;
    73: op1_10_in27 = reg_0651;
    75: op1_10_in27 = reg_0219;
    77: op1_10_in27 = imem03_in[19:16];
    78: op1_10_in27 = reg_0062;
    79: op1_10_in27 = reg_0711;
    81: op1_10_in27 = reg_0787;
    82: op1_10_in27 = imem04_in[3:0];
    83: op1_10_in27 = imem01_in[7:4];
    84: op1_10_in27 = reg_0628;
    86: op1_10_in27 = reg_0318;
    87: op1_10_in27 = reg_0577;
    88: op1_10_in27 = reg_0637;
    89: op1_10_in27 = reg_0137;
    92: op1_10_in27 = imem01_in[107:104];
    93: op1_10_in27 = reg_0425;
    94: op1_10_in27 = reg_0125;
    95: op1_10_in27 = reg_0678;
    default: op1_10_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    14: op1_10_inv27 = 1;
    16: op1_10_inv27 = 1;
    17: op1_10_inv27 = 1;
    19: op1_10_inv27 = 1;
    22: op1_10_inv27 = 1;
    25: op1_10_inv27 = 1;
    28: op1_10_inv27 = 1;
    29: op1_10_inv27 = 1;
    30: op1_10_inv27 = 1;
    33: op1_10_inv27 = 1;
    34: op1_10_inv27 = 1;
    37: op1_10_inv27 = 1;
    38: op1_10_inv27 = 1;
    39: op1_10_inv27 = 1;
    40: op1_10_inv27 = 1;
    43: op1_10_inv27 = 1;
    46: op1_10_inv27 = 1;
    47: op1_10_inv27 = 1;
    48: op1_10_inv27 = 1;
    49: op1_10_inv27 = 1;
    50: op1_10_inv27 = 1;
    53: op1_10_inv27 = 1;
    54: op1_10_inv27 = 1;
    56: op1_10_inv27 = 1;
    57: op1_10_inv27 = 1;
    59: op1_10_inv27 = 1;
    61: op1_10_inv27 = 1;
    65: op1_10_inv27 = 1;
    66: op1_10_inv27 = 1;
    68: op1_10_inv27 = 1;
    72: op1_10_inv27 = 1;
    76: op1_10_inv27 = 1;
    77: op1_10_inv27 = 1;
    78: op1_10_inv27 = 1;
    87: op1_10_inv27 = 1;
    88: op1_10_inv27 = 1;
    89: op1_10_inv27 = 1;
    93: op1_10_inv27 = 1;
    94: op1_10_inv27 = 1;
    default: op1_10_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in28 = reg_0507;
    5: op1_10_in28 = reg_0518;
    6: op1_10_in28 = imem04_in[107:104];
    7: op1_10_in28 = reg_0032;
    8: op1_10_in28 = reg_0238;
    9: op1_10_in28 = reg_0701;
    10: op1_10_in28 = reg_0319;
    12: op1_10_in28 = reg_0288;
    13: op1_10_in28 = reg_0332;
    14: op1_10_in28 = reg_0449;
    15: op1_10_in28 = imem03_in[91:88];
    16: op1_10_in28 = reg_0484;
    17: op1_10_in28 = reg_0592;
    18: op1_10_in28 = reg_0066;
    19: op1_10_in28 = reg_0098;
    20: op1_10_in28 = reg_0610;
    21: op1_10_in28 = reg_0519;
    22: op1_10_in28 = reg_0642;
    23: op1_10_in28 = reg_0227;
    24: op1_10_in28 = reg_0596;
    25: op1_10_in28 = reg_0421;
    61: op1_10_in28 = reg_0421;
    26: op1_10_in28 = reg_0255;
    27: op1_10_in28 = reg_0295;
    28: op1_10_in28 = reg_0121;
    29: op1_10_in28 = reg_0092;
    30: op1_10_in28 = reg_0091;
    78: op1_10_in28 = reg_0091;
    31: op1_10_in28 = reg_0165;
    33: op1_10_in28 = reg_0582;
    34: op1_10_in28 = imem07_in[111:108];
    35: op1_10_in28 = imem07_in[71:68];
    37: op1_10_in28 = reg_0717;
    38: op1_10_in28 = reg_0124;
    43: op1_10_in28 = reg_0124;
    39: op1_10_in28 = imem03_in[3:0];
    40: op1_10_in28 = reg_0750;
    41: op1_10_in28 = reg_0442;
    44: op1_10_in28 = reg_0138;
    45: op1_10_in28 = reg_0819;
    46: op1_10_in28 = reg_0114;
    47: op1_10_in28 = reg_0795;
    48: op1_10_in28 = reg_0370;
    49: op1_10_in28 = reg_0055;
    50: op1_10_in28 = reg_0593;
    51: op1_10_in28 = reg_0306;
    52: op1_10_in28 = reg_0387;
    53: op1_10_in28 = imem03_in[51:48];
    54: op1_10_in28 = imem06_in[19:16];
    55: op1_10_in28 = reg_0037;
    56: op1_10_in28 = reg_0405;
    57: op1_10_in28 = reg_0293;
    58: op1_10_in28 = reg_0447;
    59: op1_10_in28 = reg_0441;
    62: op1_10_in28 = reg_0644;
    63: op1_10_in28 = imem05_in[51:48];
    64: op1_10_in28 = imem06_in[71:68];
    65: op1_10_in28 = imem07_in[23:20];
    66: op1_10_in28 = reg_0141;
    67: op1_10_in28 = reg_0425;
    68: op1_10_in28 = reg_0351;
    69: op1_10_in28 = reg_0446;
    71: op1_10_in28 = imem05_in[11:8];
    72: op1_10_in28 = reg_0174;
    81: op1_10_in28 = reg_0174;
    73: op1_10_in28 = reg_0787;
    75: op1_10_in28 = reg_0105;
    76: op1_10_in28 = reg_0595;
    77: op1_10_in28 = imem03_in[71:68];
    79: op1_10_in28 = reg_0727;
    82: op1_10_in28 = imem04_in[15:12];
    83: op1_10_in28 = imem01_in[11:8];
    84: op1_10_in28 = reg_0242;
    86: op1_10_in28 = reg_0528;
    87: op1_10_in28 = reg_0349;
    88: op1_10_in28 = reg_0396;
    89: op1_10_in28 = imem06_in[39:36];
    90: op1_10_in28 = reg_0531;
    92: op1_10_in28 = imem01_in[119:116];
    93: op1_10_in28 = reg_0755;
    94: op1_10_in28 = reg_0104;
    95: op1_10_in28 = imem02_in[3:0];
    default: op1_10_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_10_inv28 = 1;
    8: op1_10_inv28 = 1;
    12: op1_10_inv28 = 1;
    13: op1_10_inv28 = 1;
    15: op1_10_inv28 = 1;
    17: op1_10_inv28 = 1;
    18: op1_10_inv28 = 1;
    19: op1_10_inv28 = 1;
    24: op1_10_inv28 = 1;
    27: op1_10_inv28 = 1;
    28: op1_10_inv28 = 1;
    31: op1_10_inv28 = 1;
    33: op1_10_inv28 = 1;
    34: op1_10_inv28 = 1;
    40: op1_10_inv28 = 1;
    45: op1_10_inv28 = 1;
    47: op1_10_inv28 = 1;
    48: op1_10_inv28 = 1;
    50: op1_10_inv28 = 1;
    51: op1_10_inv28 = 1;
    52: op1_10_inv28 = 1;
    54: op1_10_inv28 = 1;
    56: op1_10_inv28 = 1;
    57: op1_10_inv28 = 1;
    61: op1_10_inv28 = 1;
    62: op1_10_inv28 = 1;
    66: op1_10_inv28 = 1;
    67: op1_10_inv28 = 1;
    69: op1_10_inv28 = 1;
    77: op1_10_inv28 = 1;
    78: op1_10_inv28 = 1;
    81: op1_10_inv28 = 1;
    82: op1_10_inv28 = 1;
    84: op1_10_inv28 = 1;
    86: op1_10_inv28 = 1;
    94: op1_10_inv28 = 1;
    95: op1_10_inv28 = 1;
    default: op1_10_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in29 = reg_0235;
    5: op1_10_in29 = reg_0515;
    6: op1_10_in29 = reg_0555;
    7: op1_10_in29 = reg_0029;
    8: op1_10_in29 = reg_0119;
    67: op1_10_in29 = reg_0119;
    75: op1_10_in29 = reg_0119;
    9: op1_10_in29 = reg_0706;
    10: op1_10_in29 = reg_0006;
    12: op1_10_in29 = reg_0059;
    13: op1_10_in29 = reg_0344;
    14: op1_10_in29 = reg_0431;
    15: op1_10_in29 = imem03_in[95:92];
    77: op1_10_in29 = imem03_in[95:92];
    16: op1_10_in29 = reg_0794;
    17: op1_10_in29 = reg_0597;
    18: op1_10_in29 = reg_0289;
    19: op1_10_in29 = reg_0094;
    20: op1_10_in29 = reg_0621;
    21: op1_10_in29 = reg_0521;
    22: op1_10_in29 = reg_0650;
    23: op1_10_in29 = reg_0519;
    24: op1_10_in29 = reg_0568;
    25: op1_10_in29 = reg_0449;
    26: op1_10_in29 = reg_0075;
    27: op1_10_in29 = reg_0065;
    28: op1_10_in29 = imem02_in[107:104];
    29: op1_10_in29 = reg_0314;
    30: op1_10_in29 = reg_0742;
    31: op1_10_in29 = reg_0162;
    33: op1_10_in29 = reg_0395;
    34: op1_10_in29 = reg_0721;
    35: op1_10_in29 = imem07_in[87:84];
    37: op1_10_in29 = reg_0725;
    38: op1_10_in29 = reg_0100;
    39: op1_10_in29 = imem03_in[35:32];
    40: op1_10_in29 = reg_0590;
    41: op1_10_in29 = reg_0435;
    43: op1_10_in29 = reg_0104;
    44: op1_10_in29 = reg_0155;
    45: op1_10_in29 = reg_0375;
    56: op1_10_in29 = reg_0375;
    46: op1_10_in29 = imem02_in[7:4];
    95: op1_10_in29 = imem02_in[7:4];
    47: op1_10_in29 = reg_0486;
    48: op1_10_in29 = reg_0762;
    49: op1_10_in29 = reg_0516;
    50: op1_10_in29 = reg_0391;
    51: op1_10_in29 = reg_0511;
    52: op1_10_in29 = reg_0517;
    53: op1_10_in29 = imem03_in[67:64];
    54: op1_10_in29 = imem06_in[35:32];
    55: op1_10_in29 = imem07_in[83:80];
    57: op1_10_in29 = imem06_in[19:16];
    58: op1_10_in29 = reg_0434;
    59: op1_10_in29 = reg_0439;
    61: op1_10_in29 = reg_0306;
    62: op1_10_in29 = imem05_in[15:12];
    63: op1_10_in29 = imem05_in[63:60];
    64: op1_10_in29 = reg_0291;
    65: op1_10_in29 = imem07_in[31:28];
    66: op1_10_in29 = reg_0140;
    68: op1_10_in29 = reg_0323;
    69: op1_10_in29 = reg_0438;
    71: op1_10_in29 = imem05_in[23:20];
    72: op1_10_in29 = reg_0179;
    81: op1_10_in29 = reg_0179;
    73: op1_10_in29 = reg_0367;
    76: op1_10_in29 = reg_0588;
    78: op1_10_in29 = reg_0797;
    79: op1_10_in29 = reg_0253;
    82: op1_10_in29 = imem04_in[23:20];
    83: op1_10_in29 = reg_0224;
    84: op1_10_in29 = reg_0270;
    86: op1_10_in29 = reg_0483;
    87: op1_10_in29 = reg_0817;
    88: op1_10_in29 = reg_0811;
    89: op1_10_in29 = imem06_in[47:44];
    90: op1_10_in29 = reg_0393;
    92: op1_10_in29 = reg_0123;
    93: op1_10_in29 = reg_0673;
    94: op1_10_in29 = reg_0108;
    default: op1_10_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv29 = 1;
    7: op1_10_inv29 = 1;
    8: op1_10_inv29 = 1;
    9: op1_10_inv29 = 1;
    12: op1_10_inv29 = 1;
    13: op1_10_inv29 = 1;
    16: op1_10_inv29 = 1;
    17: op1_10_inv29 = 1;
    20: op1_10_inv29 = 1;
    22: op1_10_inv29 = 1;
    23: op1_10_inv29 = 1;
    25: op1_10_inv29 = 1;
    27: op1_10_inv29 = 1;
    29: op1_10_inv29 = 1;
    33: op1_10_inv29 = 1;
    37: op1_10_inv29 = 1;
    40: op1_10_inv29 = 1;
    44: op1_10_inv29 = 1;
    45: op1_10_inv29 = 1;
    47: op1_10_inv29 = 1;
    49: op1_10_inv29 = 1;
    50: op1_10_inv29 = 1;
    56: op1_10_inv29 = 1;
    57: op1_10_inv29 = 1;
    58: op1_10_inv29 = 1;
    59: op1_10_inv29 = 1;
    62: op1_10_inv29 = 1;
    63: op1_10_inv29 = 1;
    65: op1_10_inv29 = 1;
    71: op1_10_inv29 = 1;
    73: op1_10_inv29 = 1;
    76: op1_10_inv29 = 1;
    78: op1_10_inv29 = 1;
    79: op1_10_inv29 = 1;
    82: op1_10_inv29 = 1;
    83: op1_10_inv29 = 1;
    84: op1_10_inv29 = 1;
    88: op1_10_inv29 = 1;
    89: op1_10_inv29 = 1;
    90: op1_10_inv29 = 1;
    default: op1_10_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_10_in30 = reg_0239;
    5: op1_10_in30 = reg_0233;
    6: op1_10_in30 = reg_0281;
    7: op1_10_in30 = imem07_in[3:0];
    8: op1_10_in30 = reg_0108;
    9: op1_10_in30 = reg_0425;
    10: op1_10_in30 = reg_0003;
    12: op1_10_in30 = reg_0046;
    13: op1_10_in30 = reg_0383;
    14: op1_10_in30 = reg_0180;
    15: op1_10_in30 = imem03_in[115:112];
    16: op1_10_in30 = reg_0498;
    17: op1_10_in30 = reg_0395;
    18: op1_10_in30 = reg_0077;
    19: op1_10_in30 = reg_0093;
    20: op1_10_in30 = reg_0626;
    21: op1_10_in30 = reg_0515;
    22: op1_10_in30 = reg_0666;
    23: op1_10_in30 = reg_0507;
    24: op1_10_in30 = reg_0587;
    25: op1_10_in30 = reg_0444;
    26: op1_10_in30 = reg_0070;
    27: op1_10_in30 = reg_0289;
    28: op1_10_in30 = imem02_in[111:108];
    29: op1_10_in30 = reg_0530;
    30: op1_10_in30 = reg_0527;
    31: op1_10_in30 = imem06_in[71:68];
    33: op1_10_in30 = reg_0517;
    34: op1_10_in30 = reg_0703;
    35: op1_10_in30 = reg_0728;
    37: op1_10_in30 = reg_0709;
    38: op1_10_in30 = reg_0110;
    39: op1_10_in30 = imem03_in[55:52];
    40: op1_10_in30 = reg_0573;
    50: op1_10_in30 = reg_0573;
    41: op1_10_in30 = reg_0175;
    59: op1_10_in30 = reg_0175;
    43: op1_10_in30 = reg_0126;
    44: op1_10_in30 = imem06_in[7:4];
    45: op1_10_in30 = reg_0037;
    46: op1_10_in30 = imem02_in[15:12];
    47: op1_10_in30 = reg_0225;
    48: op1_10_in30 = reg_0621;
    49: op1_10_in30 = reg_0308;
    51: op1_10_in30 = reg_0567;
    52: op1_10_in30 = reg_0006;
    53: op1_10_in30 = imem03_in[87:84];
    54: op1_10_in30 = reg_0291;
    55: op1_10_in30 = reg_0730;
    56: op1_10_in30 = reg_0068;
    57: op1_10_in30 = imem06_in[63:60];
    58: op1_10_in30 = reg_0161;
    61: op1_10_in30 = reg_0502;
    62: op1_10_in30 = imem05_in[35:32];
    63: op1_10_in30 = imem05_in[67:64];
    64: op1_10_in30 = reg_0624;
    65: op1_10_in30 = imem07_in[43:40];
    66: op1_10_in30 = imem06_in[15:12];
    67: op1_10_in30 = reg_0672;
    68: op1_10_in30 = reg_0533;
    69: op1_10_in30 = reg_0172;
    71: op1_10_in30 = imem05_in[31:28];
    72: op1_10_in30 = reg_0162;
    73: op1_10_in30 = imem07_in[51:48];
    75: op1_10_in30 = reg_0120;
    76: op1_10_in30 = reg_0571;
    77: op1_10_in30 = reg_0589;
    78: op1_10_in30 = reg_0048;
    79: op1_10_in30 = reg_0445;
    81: op1_10_in30 = reg_0165;
    82: op1_10_in30 = imem04_in[79:76];
    83: op1_10_in30 = reg_0394;
    84: op1_10_in30 = reg_0218;
    86: op1_10_in30 = reg_0372;
    87: op1_10_in30 = reg_0370;
    88: op1_10_in30 = reg_0013;
    89: op1_10_in30 = imem06_in[91:88];
    90: op1_10_in30 = reg_0152;
    92: op1_10_in30 = reg_0124;
    93: op1_10_in30 = reg_0592;
    94: op1_10_in30 = reg_0675;
    95: op1_10_in30 = imem02_in[79:76];
    default: op1_10_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_10_inv30 = 1;
    7: op1_10_inv30 = 1;
    8: op1_10_inv30 = 1;
    12: op1_10_inv30 = 1;
    14: op1_10_inv30 = 1;
    15: op1_10_inv30 = 1;
    16: op1_10_inv30 = 1;
    17: op1_10_inv30 = 1;
    18: op1_10_inv30 = 1;
    20: op1_10_inv30 = 1;
    21: op1_10_inv30 = 1;
    26: op1_10_inv30 = 1;
    27: op1_10_inv30 = 1;
    30: op1_10_inv30 = 1;
    31: op1_10_inv30 = 1;
    33: op1_10_inv30 = 1;
    34: op1_10_inv30 = 1;
    37: op1_10_inv30 = 1;
    38: op1_10_inv30 = 1;
    40: op1_10_inv30 = 1;
    43: op1_10_inv30 = 1;
    44: op1_10_inv30 = 1;
    45: op1_10_inv30 = 1;
    46: op1_10_inv30 = 1;
    47: op1_10_inv30 = 1;
    53: op1_10_inv30 = 1;
    56: op1_10_inv30 = 1;
    59: op1_10_inv30 = 1;
    61: op1_10_inv30 = 1;
    62: op1_10_inv30 = 1;
    63: op1_10_inv30 = 1;
    66: op1_10_inv30 = 1;
    67: op1_10_inv30 = 1;
    68: op1_10_inv30 = 1;
    72: op1_10_inv30 = 1;
    77: op1_10_inv30 = 1;
    78: op1_10_inv30 = 1;
    81: op1_10_inv30 = 1;
    88: op1_10_inv30 = 1;
    92: op1_10_inv30 = 1;
    94: op1_10_inv30 = 1;
    default: op1_10_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_10_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_10_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in00 = reg_0240;
    5: op1_11_in00 = reg_0236;
    78: op1_11_in00 = reg_0236;
    6: op1_11_in00 = reg_0301;
    7: op1_11_in00 = imem07_in[7:4];
    8: op1_11_in00 = reg_0100;
    9: op1_11_in00 = imem00_in[59:56];
    10: op1_11_in00 = reg_0804;
    11: op1_11_in00 = imem00_in[19:16];
    12: op1_11_in00 = reg_0058;
    13: op1_11_in00 = reg_0367;
    14: op1_11_in00 = imem00_in[15:12];
    15: op1_11_in00 = imem03_in[119:116];
    16: op1_11_in00 = reg_0262;
    17: op1_11_in00 = reg_0384;
    18: op1_11_in00 = reg_0075;
    19: op1_11_in00 = imem03_in[15:12];
    3: op1_11_in00 = imem07_in[55:52];
    20: op1_11_in00 = reg_0632;
    21: op1_11_in00 = reg_0525;
    22: op1_11_in00 = reg_0637;
    23: op1_11_in00 = reg_0505;
    24: op1_11_in00 = reg_0592;
    2: op1_11_in00 = imem07_in[99:96];
    25: op1_11_in00 = imem00_in[3:0];
    26: op1_11_in00 = imem05_in[63:60];
    27: op1_11_in00 = reg_0077;
    28: op1_11_in00 = imem02_in[115:112];
    29: op1_11_in00 = reg_0540;
    30: op1_11_in00 = reg_0226;
    1: op1_11_in00 = imem07_in[31:28];
    31: op1_11_in00 = imem00_in[7:4];
    32: op1_11_in00 = imem00_in[7:4];
    60: op1_11_in00 = imem00_in[7:4];
    85: op1_11_in00 = imem00_in[7:4];
    33: op1_11_in00 = reg_0562;
    34: op1_11_in00 = reg_0432;
    35: op1_11_in00 = reg_0430;
    36: op1_11_in00 = imem00_in[123:120];
    37: op1_11_in00 = reg_0707;
    38: op1_11_in00 = imem02_in[15:12];
    39: op1_11_in00 = imem03_in[59:56];
    40: op1_11_in00 = reg_0383;
    41: op1_11_in00 = reg_0181;
    69: op1_11_in00 = reg_0181;
    42: op1_11_in00 = imem00_in[39:36];
    91: op1_11_in00 = imem00_in[39:36];
    43: op1_11_in00 = imem02_in[7:4];
    44: op1_11_in00 = imem06_in[19:16];
    45: op1_11_in00 = imem07_in[103:100];
    46: op1_11_in00 = imem02_in[55:52];
    47: op1_11_in00 = reg_0741;
    48: op1_11_in00 = reg_0375;
    49: op1_11_in00 = reg_0280;
    50: op1_11_in00 = reg_0561;
    51: op1_11_in00 = reg_0216;
    52: op1_11_in00 = reg_0001;
    53: op1_11_in00 = imem03_in[99:96];
    54: op1_11_in00 = reg_0613;
    55: op1_11_in00 = reg_0703;
    56: op1_11_in00 = imem06_in[55:52];
    57: op1_11_in00 = imem06_in[91:88];
    58: op1_11_in00 = reg_0162;
    59: op1_11_in00 = reg_0180;
    61: op1_11_in00 = reg_0603;
    62: op1_11_in00 = imem05_in[67:64];
    63: op1_11_in00 = imem05_in[71:68];
    64: op1_11_in00 = reg_0762;
    65: op1_11_in00 = imem07_in[51:48];
    66: op1_11_in00 = imem06_in[47:44];
    67: op1_11_in00 = reg_0127;
    68: op1_11_in00 = reg_0096;
    70: op1_11_in00 = imem00_in[51:48];
    71: op1_11_in00 = imem05_in[43:40];
    72: op1_11_in00 = reg_0166;
    73: op1_11_in00 = imem07_in[63:60];
    74: op1_11_in00 = imem00_in[75:72];
    75: op1_11_in00 = imem02_in[31:28];
    76: op1_11_in00 = reg_0321;
    77: op1_11_in00 = reg_0350;
    79: op1_11_in00 = reg_0434;
    80: op1_11_in00 = imem00_in[23:20];
    81: op1_11_in00 = reg_0249;
    82: op1_11_in00 = imem04_in[87:84];
    83: op1_11_in00 = reg_0759;
    84: op1_11_in00 = reg_0484;
    86: op1_11_in00 = reg_0003;
    87: op1_11_in00 = reg_0260;
    88: op1_11_in00 = reg_0007;
    89: op1_11_in00 = reg_0289;
    90: op1_11_in00 = imem06_in[15:12];
    92: op1_11_in00 = reg_0125;
    93: op1_11_in00 = reg_0108;
    94: op1_11_in00 = reg_0674;
    95: op1_11_in00 = imem02_in[87:84];
    default: op1_11_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv00 = 1;
    8: op1_11_inv00 = 1;
    10: op1_11_inv00 = 1;
    11: op1_11_inv00 = 1;
    12: op1_11_inv00 = 1;
    14: op1_11_inv00 = 1;
    19: op1_11_inv00 = 1;
    3: op1_11_inv00 = 1;
    20: op1_11_inv00 = 1;
    23: op1_11_inv00 = 1;
    24: op1_11_inv00 = 1;
    25: op1_11_inv00 = 1;
    1: op1_11_inv00 = 1;
    35: op1_11_inv00 = 1;
    38: op1_11_inv00 = 1;
    39: op1_11_inv00 = 1;
    41: op1_11_inv00 = 1;
    46: op1_11_inv00 = 1;
    47: op1_11_inv00 = 1;
    49: op1_11_inv00 = 1;
    50: op1_11_inv00 = 1;
    51: op1_11_inv00 = 1;
    56: op1_11_inv00 = 1;
    58: op1_11_inv00 = 1;
    59: op1_11_inv00 = 1;
    60: op1_11_inv00 = 1;
    61: op1_11_inv00 = 1;
    63: op1_11_inv00 = 1;
    64: op1_11_inv00 = 1;
    65: op1_11_inv00 = 1;
    66: op1_11_inv00 = 1;
    67: op1_11_inv00 = 1;
    68: op1_11_inv00 = 1;
    71: op1_11_inv00 = 1;
    72: op1_11_inv00 = 1;
    73: op1_11_inv00 = 1;
    74: op1_11_inv00 = 1;
    75: op1_11_inv00 = 1;
    76: op1_11_inv00 = 1;
    77: op1_11_inv00 = 1;
    78: op1_11_inv00 = 1;
    79: op1_11_inv00 = 1;
    80: op1_11_inv00 = 1;
    83: op1_11_inv00 = 1;
    84: op1_11_inv00 = 1;
    87: op1_11_inv00 = 1;
    88: op1_11_inv00 = 1;
    91: op1_11_inv00 = 1;
    93: op1_11_inv00 = 1;
    95: op1_11_inv00 = 1;
    default: op1_11_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in01 = reg_0234;
    5: op1_11_in01 = reg_0245;
    6: op1_11_in01 = reg_0294;
    7: op1_11_in01 = imem07_in[43:40];
    8: op1_11_in01 = reg_0101;
    9: op1_11_in01 = imem00_in[63:60];
    91: op1_11_in01 = imem00_in[63:60];
    10: op1_11_in01 = reg_0806;
    11: op1_11_in01 = imem00_in[27:24];
    60: op1_11_in01 = imem00_in[27:24];
    80: op1_11_in01 = imem00_in[27:24];
    85: op1_11_in01 = imem00_in[27:24];
    12: op1_11_in01 = imem05_in[7:4];
    27: op1_11_in01 = imem05_in[7:4];
    13: op1_11_in01 = reg_0812;
    14: op1_11_in01 = imem00_in[31:28];
    31: op1_11_in01 = imem00_in[31:28];
    15: op1_11_in01 = imem03_in[123:120];
    16: op1_11_in01 = reg_0259;
    17: op1_11_in01 = reg_0317;
    18: op1_11_in01 = imem05_in[55:52];
    71: op1_11_in01 = imem05_in[55:52];
    19: op1_11_in01 = imem03_in[39:36];
    3: op1_11_in01 = reg_0441;
    37: op1_11_in01 = reg_0441;
    20: op1_11_in01 = reg_0601;
    21: op1_11_in01 = reg_0505;
    22: op1_11_in01 = reg_0639;
    23: op1_11_in01 = reg_0506;
    24: op1_11_in01 = reg_0589;
    2: op1_11_in01 = imem07_in[111:108];
    25: op1_11_in01 = imem00_in[15:12];
    26: op1_11_in01 = imem05_in[75:72];
    28: op1_11_in01 = imem02_in[123:120];
    29: op1_11_in01 = reg_0498;
    68: op1_11_in01 = reg_0498;
    30: op1_11_in01 = reg_0307;
    1: op1_11_in01 = imem07_in[35:32];
    32: op1_11_in01 = imem00_in[71:68];
    42: op1_11_in01 = imem00_in[71:68];
    33: op1_11_in01 = reg_0499;
    34: op1_11_in01 = reg_0421;
    35: op1_11_in01 = reg_0433;
    36: op1_11_in01 = reg_0693;
    38: op1_11_in01 = imem02_in[43:40];
    39: op1_11_in01 = imem03_in[83:80];
    40: op1_11_in01 = reg_0385;
    41: op1_11_in01 = reg_0160;
    43: op1_11_in01 = imem02_in[39:36];
    44: op1_11_in01 = imem06_in[39:36];
    45: op1_11_in01 = reg_0716;
    46: op1_11_in01 = imem02_in[59:56];
    47: op1_11_in01 = reg_0276;
    48: op1_11_in01 = reg_0367;
    49: op1_11_in01 = reg_0529;
    50: op1_11_in01 = reg_0373;
    51: op1_11_in01 = reg_0290;
    52: op1_11_in01 = reg_0013;
    53: op1_11_in01 = imem03_in[107:104];
    54: op1_11_in01 = reg_0371;
    55: op1_11_in01 = reg_0707;
    56: op1_11_in01 = imem06_in[83:80];
    57: op1_11_in01 = imem06_in[127:124];
    58: op1_11_in01 = reg_0177;
    59: op1_11_in01 = reg_0169;
    61: op1_11_in01 = reg_0219;
    62: op1_11_in01 = imem05_in[71:68];
    63: op1_11_in01 = imem05_in[103:100];
    64: op1_11_in01 = reg_0298;
    65: op1_11_in01 = imem07_in[71:68];
    73: op1_11_in01 = imem07_in[71:68];
    66: op1_11_in01 = reg_0291;
    67: op1_11_in01 = reg_0676;
    69: op1_11_in01 = reg_0162;
    70: op1_11_in01 = imem00_in[59:56];
    72: op1_11_in01 = reg_0168;
    74: op1_11_in01 = imem00_in[79:76];
    75: op1_11_in01 = imem02_in[35:32];
    76: op1_11_in01 = reg_0572;
    77: op1_11_in01 = reg_0600;
    78: op1_11_in01 = reg_0666;
    79: op1_11_in01 = reg_0437;
    81: op1_11_in01 = reg_0717;
    82: op1_11_in01 = imem04_in[115:112];
    83: op1_11_in01 = reg_0388;
    84: op1_11_in01 = reg_0501;
    86: op1_11_in01 = reg_0803;
    87: op1_11_in01 = reg_0628;
    88: op1_11_in01 = reg_0807;
    89: op1_11_in01 = reg_0346;
    90: op1_11_in01 = imem06_in[19:16];
    92: op1_11_in01 = reg_0660;
    93: op1_11_in01 = imem02_in[3:0];
    94: op1_11_in01 = imem02_in[23:20];
    95: op1_11_in01 = reg_0057;
    default: op1_11_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv01 = 1;
    5: op1_11_inv01 = 1;
    6: op1_11_inv01 = 1;
    7: op1_11_inv01 = 1;
    8: op1_11_inv01 = 1;
    11: op1_11_inv01 = 1;
    13: op1_11_inv01 = 1;
    14: op1_11_inv01 = 1;
    17: op1_11_inv01 = 1;
    18: op1_11_inv01 = 1;
    20: op1_11_inv01 = 1;
    21: op1_11_inv01 = 1;
    23: op1_11_inv01 = 1;
    26: op1_11_inv01 = 1;
    27: op1_11_inv01 = 1;
    29: op1_11_inv01 = 1;
    30: op1_11_inv01 = 1;
    1: op1_11_inv01 = 1;
    31: op1_11_inv01 = 1;
    32: op1_11_inv01 = 1;
    36: op1_11_inv01 = 1;
    37: op1_11_inv01 = 1;
    38: op1_11_inv01 = 1;
    41: op1_11_inv01 = 1;
    44: op1_11_inv01 = 1;
    48: op1_11_inv01 = 1;
    49: op1_11_inv01 = 1;
    55: op1_11_inv01 = 1;
    56: op1_11_inv01 = 1;
    58: op1_11_inv01 = 1;
    59: op1_11_inv01 = 1;
    60: op1_11_inv01 = 1;
    61: op1_11_inv01 = 1;
    63: op1_11_inv01 = 1;
    64: op1_11_inv01 = 1;
    65: op1_11_inv01 = 1;
    66: op1_11_inv01 = 1;
    68: op1_11_inv01 = 1;
    71: op1_11_inv01 = 1;
    73: op1_11_inv01 = 1;
    78: op1_11_inv01 = 1;
    80: op1_11_inv01 = 1;
    82: op1_11_inv01 = 1;
    85: op1_11_inv01 = 1;
    86: op1_11_inv01 = 1;
    89: op1_11_inv01 = 1;
    90: op1_11_inv01 = 1;
    92: op1_11_inv01 = 1;
    93: op1_11_inv01 = 1;
    94: op1_11_inv01 = 1;
    default: op1_11_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in02 = reg_0101;
    5: op1_11_in02 = reg_0221;
    6: op1_11_in02 = reg_0276;
    7: op1_11_in02 = imem07_in[51:48];
    8: op1_11_in02 = reg_0121;
    67: op1_11_in02 = reg_0121;
    9: op1_11_in02 = imem00_in[71:68];
    10: op1_11_in02 = reg_0810;
    88: op1_11_in02 = reg_0810;
    11: op1_11_in02 = imem00_in[67:64];
    25: op1_11_in02 = imem00_in[67:64];
    12: op1_11_in02 = imem05_in[15:12];
    13: op1_11_in02 = reg_0747;
    14: op1_11_in02 = imem00_in[35:32];
    80: op1_11_in02 = imem00_in[35:32];
    15: op1_11_in02 = reg_0579;
    16: op1_11_in02 = reg_0270;
    17: op1_11_in02 = reg_0343;
    18: op1_11_in02 = imem05_in[103:100];
    19: op1_11_in02 = imem03_in[95:92];
    3: op1_11_in02 = reg_0432;
    20: op1_11_in02 = reg_0349;
    66: op1_11_in02 = reg_0349;
    21: op1_11_in02 = reg_0511;
    22: op1_11_in02 = reg_0665;
    23: op1_11_in02 = reg_0216;
    24: op1_11_in02 = reg_0593;
    2: op1_11_in02 = imem07_in[115:112];
    26: op1_11_in02 = imem05_in[99:96];
    27: op1_11_in02 = imem05_in[19:16];
    28: op1_11_in02 = reg_0658;
    29: op1_11_in02 = imem03_in[27:24];
    30: op1_11_in02 = reg_0132;
    1: op1_11_in02 = imem07_in[43:40];
    31: op1_11_in02 = imem00_in[59:56];
    32: op1_11_in02 = imem00_in[75:72];
    33: op1_11_in02 = reg_0570;
    50: op1_11_in02 = reg_0570;
    34: op1_11_in02 = reg_0426;
    35: op1_11_in02 = reg_0440;
    36: op1_11_in02 = reg_0674;
    37: op1_11_in02 = reg_0429;
    38: op1_11_in02 = reg_0645;
    39: op1_11_in02 = imem03_in[103:100];
    40: op1_11_in02 = reg_0562;
    41: op1_11_in02 = reg_0158;
    42: op1_11_in02 = imem00_in[123:120];
    43: op1_11_in02 = imem02_in[51:48];
    44: op1_11_in02 = imem06_in[43:40];
    45: op1_11_in02 = reg_0725;
    46: op1_11_in02 = imem02_in[87:84];
    47: op1_11_in02 = reg_0269;
    48: op1_11_in02 = imem07_in[39:36];
    49: op1_11_in02 = reg_0611;
    51: op1_11_in02 = reg_0119;
    61: op1_11_in02 = reg_0119;
    52: op1_11_in02 = reg_0007;
    86: op1_11_in02 = reg_0007;
    53: op1_11_in02 = reg_0395;
    54: op1_11_in02 = reg_0606;
    55: op1_11_in02 = reg_0084;
    56: op1_11_in02 = imem06_in[123:120];
    57: op1_11_in02 = reg_0028;
    58: op1_11_in02 = reg_0170;
    59: op1_11_in02 = reg_0168;
    60: op1_11_in02 = imem00_in[111:108];
    62: op1_11_in02 = imem05_in[123:120];
    63: op1_11_in02 = reg_0791;
    64: op1_11_in02 = reg_0619;
    65: op1_11_in02 = imem07_in[79:76];
    68: op1_11_in02 = imem03_in[3:0];
    69: op1_11_in02 = reg_0159;
    70: op1_11_in02 = imem00_in[127:124];
    71: op1_11_in02 = imem05_in[71:68];
    72: op1_11_in02 = reg_0173;
    73: op1_11_in02 = imem07_in[103:100];
    74: op1_11_in02 = imem00_in[83:80];
    75: op1_11_in02 = imem02_in[39:36];
    76: op1_11_in02 = reg_0549;
    77: op1_11_in02 = reg_0595;
    78: op1_11_in02 = reg_0489;
    79: op1_11_in02 = reg_0267;
    81: op1_11_in02 = reg_0177;
    82: op1_11_in02 = imem04_in[127:124];
    83: op1_11_in02 = reg_0418;
    84: op1_11_in02 = reg_0787;
    85: op1_11_in02 = imem00_in[31:28];
    87: op1_11_in02 = reg_0630;
    89: op1_11_in02 = reg_0618;
    90: op1_11_in02 = imem06_in[27:24];
    91: op1_11_in02 = imem00_in[79:76];
    92: op1_11_in02 = reg_0601;
    93: op1_11_in02 = imem02_in[11:8];
    94: op1_11_in02 = reg_0264;
    95: op1_11_in02 = reg_0081;
    default: op1_11_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv02 = 1;
    6: op1_11_inv02 = 1;
    8: op1_11_inv02 = 1;
    11: op1_11_inv02 = 1;
    13: op1_11_inv02 = 1;
    15: op1_11_inv02 = 1;
    16: op1_11_inv02 = 1;
    17: op1_11_inv02 = 1;
    18: op1_11_inv02 = 1;
    19: op1_11_inv02 = 1;
    22: op1_11_inv02 = 1;
    24: op1_11_inv02 = 1;
    2: op1_11_inv02 = 1;
    25: op1_11_inv02 = 1;
    27: op1_11_inv02 = 1;
    31: op1_11_inv02 = 1;
    32: op1_11_inv02 = 1;
    33: op1_11_inv02 = 1;
    37: op1_11_inv02 = 1;
    38: op1_11_inv02 = 1;
    42: op1_11_inv02 = 1;
    43: op1_11_inv02 = 1;
    48: op1_11_inv02 = 1;
    54: op1_11_inv02 = 1;
    55: op1_11_inv02 = 1;
    56: op1_11_inv02 = 1;
    57: op1_11_inv02 = 1;
    59: op1_11_inv02 = 1;
    60: op1_11_inv02 = 1;
    61: op1_11_inv02 = 1;
    67: op1_11_inv02 = 1;
    69: op1_11_inv02 = 1;
    71: op1_11_inv02 = 1;
    76: op1_11_inv02 = 1;
    79: op1_11_inv02 = 1;
    80: op1_11_inv02 = 1;
    81: op1_11_inv02 = 1;
    82: op1_11_inv02 = 1;
    84: op1_11_inv02 = 1;
    87: op1_11_inv02 = 1;
    88: op1_11_inv02 = 1;
    91: op1_11_inv02 = 1;
    92: op1_11_inv02 = 1;
    94: op1_11_inv02 = 1;
    95: op1_11_inv02 = 1;
    default: op1_11_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in03 = reg_0659;
    5: op1_11_in03 = reg_0105;
    6: op1_11_in03 = reg_0295;
    7: op1_11_in03 = imem07_in[55:52];
    8: op1_11_in03 = reg_0650;
    9: op1_11_in03 = imem00_in[87:84];
    10: op1_11_in03 = imem04_in[11:8];
    11: op1_11_in03 = imem00_in[75:72];
    12: op1_11_in03 = imem05_in[35:32];
    13: op1_11_in03 = reg_0040;
    14: op1_11_in03 = imem00_in[83:80];
    32: op1_11_in03 = imem00_in[83:80];
    85: op1_11_in03 = imem00_in[83:80];
    15: op1_11_in03 = reg_0580;
    16: op1_11_in03 = reg_0264;
    17: op1_11_in03 = reg_0388;
    18: op1_11_in03 = reg_0792;
    62: op1_11_in03 = reg_0792;
    19: op1_11_in03 = imem03_in[99:96];
    3: op1_11_in03 = reg_0445;
    20: op1_11_in03 = reg_0403;
    21: op1_11_in03 = reg_0217;
    22: op1_11_in03 = reg_0667;
    23: op1_11_in03 = reg_0247;
    24: op1_11_in03 = reg_0576;
    2: op1_11_in03 = imem07_in[127:124];
    25: op1_11_in03 = reg_0694;
    26: op1_11_in03 = reg_0483;
    27: op1_11_in03 = imem05_in[31:28];
    28: op1_11_in03 = reg_0664;
    38: op1_11_in03 = reg_0664;
    29: op1_11_in03 = imem03_in[51:48];
    30: op1_11_in03 = reg_0133;
    1: op1_11_in03 = imem07_in[87:84];
    31: op1_11_in03 = reg_0681;
    42: op1_11_in03 = reg_0681;
    33: op1_11_in03 = reg_0003;
    34: op1_11_in03 = reg_0423;
    35: op1_11_in03 = reg_0444;
    36: op1_11_in03 = reg_0680;
    37: op1_11_in03 = reg_0440;
    39: op1_11_in03 = imem03_in[127:124];
    40: op1_11_in03 = reg_0397;
    43: op1_11_in03 = imem02_in[75:72];
    44: op1_11_in03 = imem06_in[75:72];
    45: op1_11_in03 = reg_0724;
    46: op1_11_in03 = imem02_in[107:104];
    47: op1_11_in03 = reg_0272;
    48: op1_11_in03 = imem07_in[67:64];
    49: op1_11_in03 = reg_0077;
    50: op1_11_in03 = reg_0012;
    51: op1_11_in03 = reg_0120;
    61: op1_11_in03 = reg_0120;
    52: op1_11_in03 = reg_0807;
    53: op1_11_in03 = reg_0384;
    54: op1_11_in03 = reg_0339;
    89: op1_11_in03 = reg_0339;
    55: op1_11_in03 = reg_0268;
    56: op1_11_in03 = reg_0025;
    57: op1_11_in03 = reg_0777;
    58: op1_11_in03 = reg_0157;
    59: op1_11_in03 = reg_0157;
    60: op1_11_in03 = imem00_in[119:116];
    63: op1_11_in03 = reg_0490;
    64: op1_11_in03 = reg_0260;
    65: op1_11_in03 = reg_0728;
    66: op1_11_in03 = reg_0409;
    67: op1_11_in03 = reg_0678;
    92: op1_11_in03 = reg_0678;
    68: op1_11_in03 = imem03_in[11:8];
    69: op1_11_in03 = reg_0169;
    70: op1_11_in03 = reg_0697;
    71: op1_11_in03 = imem05_in[103:100];
    73: op1_11_in03 = reg_0719;
    74: op1_11_in03 = imem00_in[123:120];
    75: op1_11_in03 = imem02_in[55:52];
    76: op1_11_in03 = reg_0637;
    77: op1_11_in03 = reg_0751;
    78: op1_11_in03 = imem05_in[11:8];
    79: op1_11_in03 = reg_0438;
    80: op1_11_in03 = imem00_in[47:44];
    81: op1_11_in03 = reg_0173;
    82: op1_11_in03 = reg_0429;
    83: op1_11_in03 = reg_0502;
    84: op1_11_in03 = imem07_in[7:4];
    86: op1_11_in03 = reg_0801;
    87: op1_11_in03 = reg_0270;
    88: op1_11_in03 = imem04_in[15:12];
    90: op1_11_in03 = imem06_in[35:32];
    91: op1_11_in03 = imem00_in[99:96];
    93: op1_11_in03 = imem02_in[15:12];
    94: op1_11_in03 = reg_0656;
    95: op1_11_in03 = reg_0080;
    default: op1_11_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv03 = 1;
    7: op1_11_inv03 = 1;
    8: op1_11_inv03 = 1;
    9: op1_11_inv03 = 1;
    13: op1_11_inv03 = 1;
    16: op1_11_inv03 = 1;
    18: op1_11_inv03 = 1;
    3: op1_11_inv03 = 1;
    20: op1_11_inv03 = 1;
    24: op1_11_inv03 = 1;
    30: op1_11_inv03 = 1;
    32: op1_11_inv03 = 1;
    34: op1_11_inv03 = 1;
    35: op1_11_inv03 = 1;
    37: op1_11_inv03 = 1;
    39: op1_11_inv03 = 1;
    40: op1_11_inv03 = 1;
    42: op1_11_inv03 = 1;
    43: op1_11_inv03 = 1;
    44: op1_11_inv03 = 1;
    45: op1_11_inv03 = 1;
    47: op1_11_inv03 = 1;
    56: op1_11_inv03 = 1;
    62: op1_11_inv03 = 1;
    68: op1_11_inv03 = 1;
    69: op1_11_inv03 = 1;
    73: op1_11_inv03 = 1;
    74: op1_11_inv03 = 1;
    75: op1_11_inv03 = 1;
    76: op1_11_inv03 = 1;
    77: op1_11_inv03 = 1;
    78: op1_11_inv03 = 1;
    81: op1_11_inv03 = 1;
    82: op1_11_inv03 = 1;
    84: op1_11_inv03 = 1;
    85: op1_11_inv03 = 1;
    86: op1_11_inv03 = 1;
    87: op1_11_inv03 = 1;
    94: op1_11_inv03 = 1;
    95: op1_11_inv03 = 1;
    default: op1_11_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in04 = reg_0334;
    5: op1_11_in04 = reg_0116;
    6: op1_11_in04 = reg_0307;
    7: op1_11_in04 = imem07_in[83:80];
    48: op1_11_in04 = imem07_in[83:80];
    8: op1_11_in04 = reg_0653;
    9: op1_11_in04 = reg_0679;
    10: op1_11_in04 = imem04_in[15:12];
    11: op1_11_in04 = imem00_in[95:92];
    32: op1_11_in04 = imem00_in[95:92];
    12: op1_11_in04 = imem05_in[67:64];
    13: op1_11_in04 = reg_0029;
    14: op1_11_in04 = reg_0682;
    15: op1_11_in04 = reg_0578;
    16: op1_11_in04 = reg_0147;
    17: op1_11_in04 = reg_0362;
    18: op1_11_in04 = reg_0796;
    62: op1_11_in04 = reg_0796;
    19: op1_11_in04 = imem03_in[107:104];
    3: op1_11_in04 = reg_0437;
    34: op1_11_in04 = reg_0437;
    20: op1_11_in04 = reg_0406;
    21: op1_11_in04 = reg_0503;
    22: op1_11_in04 = reg_0325;
    23: op1_11_in04 = reg_0236;
    24: op1_11_in04 = reg_0391;
    2: op1_11_in04 = reg_0159;
    25: op1_11_in04 = reg_0688;
    26: op1_11_in04 = reg_0797;
    27: op1_11_in04 = imem05_in[59:56];
    28: op1_11_in04 = reg_0639;
    29: op1_11_in04 = imem03_in[71:68];
    30: op1_11_in04 = reg_0156;
    31: op1_11_in04 = reg_0676;
    33: op1_11_in04 = reg_0803;
    35: op1_11_in04 = reg_0442;
    36: op1_11_in04 = reg_0699;
    37: op1_11_in04 = reg_0169;
    38: op1_11_in04 = reg_0661;
    39: op1_11_in04 = reg_0583;
    40: op1_11_in04 = reg_0396;
    42: op1_11_in04 = reg_0696;
    43: op1_11_in04 = imem02_in[87:84];
    44: op1_11_in04 = imem06_in[83:80];
    45: op1_11_in04 = reg_0441;
    46: op1_11_in04 = reg_0654;
    47: op1_11_in04 = reg_0149;
    49: op1_11_in04 = reg_0616;
    50: op1_11_in04 = reg_0001;
    51: op1_11_in04 = reg_0121;
    52: op1_11_in04 = reg_0800;
    53: op1_11_in04 = reg_0561;
    54: op1_11_in04 = reg_0622;
    56: op1_11_in04 = reg_0408;
    57: op1_11_in04 = reg_0040;
    58: op1_11_in04 = reg_0158;
    59: op1_11_in04 = reg_0184;
    60: op1_11_in04 = reg_0695;
    74: op1_11_in04 = reg_0695;
    61: op1_11_in04 = reg_0674;
    63: op1_11_in04 = reg_0489;
    64: op1_11_in04 = reg_0242;
    65: op1_11_in04 = reg_0704;
    66: op1_11_in04 = reg_0609;
    67: op1_11_in04 = imem02_in[7:4];
    68: op1_11_in04 = imem03_in[63:60];
    69: op1_11_in04 = reg_0182;
    70: op1_11_in04 = reg_0690;
    71: op1_11_in04 = imem05_in[119:116];
    73: op1_11_in04 = reg_0724;
    75: op1_11_in04 = imem02_in[67:64];
    76: op1_11_in04 = reg_0623;
    77: op1_11_in04 = reg_0564;
    78: op1_11_in04 = imem05_in[51:48];
    79: op1_11_in04 = reg_0183;
    80: op1_11_in04 = imem00_in[51:48];
    81: op1_11_in04 = reg_0171;
    82: op1_11_in04 = reg_0529;
    83: op1_11_in04 = reg_0104;
    84: op1_11_in04 = imem07_in[11:8];
    85: op1_11_in04 = imem00_in[107:104];
    86: op1_11_in04 = reg_0014;
    87: op1_11_in04 = reg_0750;
    88: op1_11_in04 = imem04_in[23:20];
    89: op1_11_in04 = reg_0265;
    90: op1_11_in04 = imem06_in[87:84];
    91: op1_11_in04 = imem00_in[115:112];
    92: op1_11_in04 = imem02_in[11:8];
    93: op1_11_in04 = imem02_in[39:36];
    94: op1_11_in04 = reg_0087;
    95: op1_11_in04 = reg_0392;
    default: op1_11_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv04 = 1;
    5: op1_11_inv04 = 1;
    7: op1_11_inv04 = 1;
    9: op1_11_inv04 = 1;
    11: op1_11_inv04 = 1;
    13: op1_11_inv04 = 1;
    14: op1_11_inv04 = 1;
    15: op1_11_inv04 = 1;
    16: op1_11_inv04 = 1;
    19: op1_11_inv04 = 1;
    20: op1_11_inv04 = 1;
    22: op1_11_inv04 = 1;
    25: op1_11_inv04 = 1;
    30: op1_11_inv04 = 1;
    31: op1_11_inv04 = 1;
    33: op1_11_inv04 = 1;
    34: op1_11_inv04 = 1;
    37: op1_11_inv04 = 1;
    39: op1_11_inv04 = 1;
    40: op1_11_inv04 = 1;
    46: op1_11_inv04 = 1;
    47: op1_11_inv04 = 1;
    48: op1_11_inv04 = 1;
    49: op1_11_inv04 = 1;
    50: op1_11_inv04 = 1;
    52: op1_11_inv04 = 1;
    53: op1_11_inv04 = 1;
    54: op1_11_inv04 = 1;
    56: op1_11_inv04 = 1;
    57: op1_11_inv04 = 1;
    58: op1_11_inv04 = 1;
    60: op1_11_inv04 = 1;
    61: op1_11_inv04 = 1;
    63: op1_11_inv04 = 1;
    65: op1_11_inv04 = 1;
    66: op1_11_inv04 = 1;
    68: op1_11_inv04 = 1;
    77: op1_11_inv04 = 1;
    78: op1_11_inv04 = 1;
    79: op1_11_inv04 = 1;
    81: op1_11_inv04 = 1;
    82: op1_11_inv04 = 1;
    83: op1_11_inv04 = 1;
    84: op1_11_inv04 = 1;
    85: op1_11_inv04 = 1;
    88: op1_11_inv04 = 1;
    90: op1_11_inv04 = 1;
    91: op1_11_inv04 = 1;
    92: op1_11_inv04 = 1;
    default: op1_11_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in05 = reg_0350;
    5: op1_11_in05 = reg_0119;
    6: op1_11_in05 = reg_0054;
    7: op1_11_in05 = imem07_in[119:116];
    8: op1_11_in05 = reg_0656;
    95: op1_11_in05 = reg_0656;
    9: op1_11_in05 = reg_0688;
    10: op1_11_in05 = imem04_in[51:48];
    11: op1_11_in05 = reg_0693;
    12: op1_11_in05 = imem05_in[75:72];
    27: op1_11_in05 = imem05_in[75:72];
    13: op1_11_in05 = imem07_in[11:8];
    14: op1_11_in05 = reg_0681;
    15: op1_11_in05 = reg_0576;
    16: op1_11_in05 = reg_0149;
    17: op1_11_in05 = reg_0385;
    18: op1_11_in05 = reg_0493;
    19: op1_11_in05 = reg_0585;
    3: op1_11_in05 = reg_0420;
    20: op1_11_in05 = reg_0337;
    21: op1_11_in05 = reg_0236;
    22: op1_11_in05 = reg_0345;
    23: op1_11_in05 = reg_0238;
    66: op1_11_in05 = reg_0238;
    24: op1_11_in05 = reg_0360;
    25: op1_11_in05 = reg_0465;
    26: op1_11_in05 = reg_0484;
    28: op1_11_in05 = reg_0651;
    29: op1_11_in05 = imem03_in[87:84];
    30: op1_11_in05 = imem06_in[11:8];
    31: op1_11_in05 = reg_0671;
    32: op1_11_in05 = reg_0697;
    33: op1_11_in05 = reg_0807;
    34: op1_11_in05 = reg_0431;
    35: op1_11_in05 = reg_0160;
    36: op1_11_in05 = reg_0470;
    37: op1_11_in05 = reg_0178;
    38: op1_11_in05 = reg_0358;
    39: op1_11_in05 = reg_0594;
    40: op1_11_in05 = reg_0000;
    42: op1_11_in05 = reg_0676;
    43: op1_11_in05 = imem02_in[111:108];
    44: op1_11_in05 = imem06_in[87:84];
    45: op1_11_in05 = reg_0061;
    46: op1_11_in05 = reg_0657;
    47: op1_11_in05 = reg_0135;
    48: op1_11_in05 = reg_0722;
    49: op1_11_in05 = reg_0292;
    50: op1_11_in05 = reg_0803;
    51: op1_11_in05 = reg_0349;
    52: op1_11_in05 = imem04_in[7:4];
    53: op1_11_in05 = reg_0755;
    54: op1_11_in05 = reg_0405;
    56: op1_11_in05 = reg_0773;
    57: op1_11_in05 = reg_0621;
    60: op1_11_in05 = reg_0683;
    61: op1_11_in05 = imem02_in[23:20];
    62: op1_11_in05 = reg_0797;
    63: op1_11_in05 = reg_0215;
    64: op1_11_in05 = reg_0369;
    65: op1_11_in05 = reg_0720;
    67: op1_11_in05 = imem02_in[15:12];
    68: op1_11_in05 = imem03_in[67:64];
    69: op1_11_in05 = reg_0183;
    70: op1_11_in05 = reg_0699;
    71: op1_11_in05 = imem05_in[127:124];
    73: op1_11_in05 = reg_0636;
    74: op1_11_in05 = reg_0694;
    75: op1_11_in05 = imem02_in[87:84];
    76: op1_11_in05 = reg_0019;
    77: op1_11_in05 = reg_0568;
    78: op1_11_in05 = imem05_in[111:108];
    79: op1_11_in05 = reg_0185;
    80: op1_11_in05 = imem00_in[55:52];
    81: op1_11_in05 = reg_0132;
    82: op1_11_in05 = reg_0508;
    83: op1_11_in05 = reg_0675;
    84: op1_11_in05 = imem07_in[43:40];
    85: op1_11_in05 = imem00_in[111:108];
    86: op1_11_in05 = reg_0802;
    87: op1_11_in05 = reg_0608;
    88: op1_11_in05 = imem04_in[43:40];
    89: op1_11_in05 = reg_0260;
    90: op1_11_in05 = imem06_in[119:116];
    91: op1_11_in05 = reg_0189;
    92: op1_11_in05 = imem02_in[39:36];
    93: op1_11_in05 = imem02_in[43:40];
    94: op1_11_in05 = reg_0705;
    default: op1_11_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_11_inv05 = 1;
    8: op1_11_inv05 = 1;
    9: op1_11_inv05 = 1;
    11: op1_11_inv05 = 1;
    12: op1_11_inv05 = 1;
    13: op1_11_inv05 = 1;
    14: op1_11_inv05 = 1;
    16: op1_11_inv05 = 1;
    17: op1_11_inv05 = 1;
    18: op1_11_inv05 = 1;
    23: op1_11_inv05 = 1;
    24: op1_11_inv05 = 1;
    26: op1_11_inv05 = 1;
    28: op1_11_inv05 = 1;
    33: op1_11_inv05 = 1;
    35: op1_11_inv05 = 1;
    36: op1_11_inv05 = 1;
    37: op1_11_inv05 = 1;
    39: op1_11_inv05 = 1;
    40: op1_11_inv05 = 1;
    44: op1_11_inv05 = 1;
    45: op1_11_inv05 = 1;
    46: op1_11_inv05 = 1;
    47: op1_11_inv05 = 1;
    48: op1_11_inv05 = 1;
    49: op1_11_inv05 = 1;
    50: op1_11_inv05 = 1;
    51: op1_11_inv05 = 1;
    57: op1_11_inv05 = 1;
    61: op1_11_inv05 = 1;
    63: op1_11_inv05 = 1;
    65: op1_11_inv05 = 1;
    66: op1_11_inv05 = 1;
    67: op1_11_inv05 = 1;
    68: op1_11_inv05 = 1;
    70: op1_11_inv05 = 1;
    71: op1_11_inv05 = 1;
    73: op1_11_inv05 = 1;
    75: op1_11_inv05 = 1;
    77: op1_11_inv05 = 1;
    78: op1_11_inv05 = 1;
    79: op1_11_inv05 = 1;
    80: op1_11_inv05 = 1;
    82: op1_11_inv05 = 1;
    83: op1_11_inv05 = 1;
    85: op1_11_inv05 = 1;
    87: op1_11_inv05 = 1;
    89: op1_11_inv05 = 1;
    94: op1_11_inv05 = 1;
    default: op1_11_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in06 = reg_0085;
    5: op1_11_in06 = reg_0106;
    51: op1_11_in06 = reg_0106;
    6: op1_11_in06 = reg_0041;
    7: op1_11_in06 = reg_0719;
    48: op1_11_in06 = reg_0719;
    8: op1_11_in06 = reg_0639;
    46: op1_11_in06 = reg_0639;
    9: op1_11_in06 = reg_0699;
    10: op1_11_in06 = imem04_in[87:84];
    11: op1_11_in06 = reg_0694;
    12: op1_11_in06 = imem05_in[115:112];
    27: op1_11_in06 = imem05_in[115:112];
    13: op1_11_in06 = imem07_in[75:72];
    14: op1_11_in06 = reg_0685;
    15: op1_11_in06 = reg_0388;
    53: op1_11_in06 = reg_0388;
    16: op1_11_in06 = reg_0133;
    17: op1_11_in06 = reg_0396;
    18: op1_11_in06 = reg_0793;
    19: op1_11_in06 = reg_0362;
    3: op1_11_in06 = reg_0179;
    20: op1_11_in06 = reg_0747;
    21: op1_11_in06 = reg_0234;
    22: op1_11_in06 = reg_0339;
    23: op1_11_in06 = reg_0125;
    24: op1_11_in06 = reg_0361;
    25: op1_11_in06 = reg_0476;
    26: op1_11_in06 = reg_0491;
    28: op1_11_in06 = reg_0643;
    29: op1_11_in06 = imem03_in[95:92];
    30: op1_11_in06 = imem06_in[15:12];
    31: op1_11_in06 = reg_0668;
    32: op1_11_in06 = reg_0683;
    33: op1_11_in06 = reg_0801;
    34: op1_11_in06 = reg_0175;
    35: op1_11_in06 = reg_0163;
    36: op1_11_in06 = reg_0471;
    38: op1_11_in06 = reg_0354;
    39: op1_11_in06 = reg_0573;
    40: op1_11_in06 = reg_0013;
    42: op1_11_in06 = reg_0689;
    43: op1_11_in06 = reg_0664;
    44: op1_11_in06 = imem06_in[115:112];
    45: op1_11_in06 = reg_0442;
    47: op1_11_in06 = reg_0139;
    49: op1_11_in06 = reg_0520;
    50: op1_11_in06 = reg_0805;
    52: op1_11_in06 = imem04_in[27:24];
    54: op1_11_in06 = reg_0821;
    56: op1_11_in06 = reg_0777;
    87: op1_11_in06 = reg_0777;
    57: op1_11_in06 = reg_0231;
    60: op1_11_in06 = reg_0696;
    61: op1_11_in06 = imem02_in[55:52];
    62: op1_11_in06 = reg_0490;
    77: op1_11_in06 = reg_0490;
    63: op1_11_in06 = reg_0304;
    64: op1_11_in06 = reg_0775;
    65: op1_11_in06 = reg_0702;
    66: op1_11_in06 = reg_0265;
    67: op1_11_in06 = imem02_in[23:20];
    68: op1_11_in06 = reg_0488;
    69: op1_11_in06 = reg_0173;
    70: op1_11_in06 = reg_0454;
    71: op1_11_in06 = reg_0736;
    73: op1_11_in06 = reg_0434;
    74: op1_11_in06 = reg_0690;
    75: op1_11_in06 = imem02_in[95:92];
    76: op1_11_in06 = reg_0003;
    78: op1_11_in06 = reg_0812;
    80: op1_11_in06 = imem00_in[71:68];
    81: op1_11_in06 = reg_0168;
    82: op1_11_in06 = reg_0614;
    83: op1_11_in06 = reg_0107;
    84: op1_11_in06 = imem07_in[51:48];
    85: op1_11_in06 = reg_0695;
    86: op1_11_in06 = reg_0009;
    88: op1_11_in06 = imem04_in[47:44];
    89: op1_11_in06 = reg_0630;
    90: op1_11_in06 = reg_0346;
    91: op1_11_in06 = reg_0077;
    92: op1_11_in06 = imem02_in[43:40];
    93: op1_11_in06 = imem02_in[51:48];
    94: op1_11_in06 = reg_0256;
    95: op1_11_in06 = reg_0374;
    default: op1_11_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv06 = 1;
    5: op1_11_inv06 = 1;
    7: op1_11_inv06 = 1;
    8: op1_11_inv06 = 1;
    9: op1_11_inv06 = 1;
    11: op1_11_inv06 = 1;
    13: op1_11_inv06 = 1;
    14: op1_11_inv06 = 1;
    15: op1_11_inv06 = 1;
    3: op1_11_inv06 = 1;
    20: op1_11_inv06 = 1;
    21: op1_11_inv06 = 1;
    23: op1_11_inv06 = 1;
    24: op1_11_inv06 = 1;
    25: op1_11_inv06 = 1;
    26: op1_11_inv06 = 1;
    27: op1_11_inv06 = 1;
    31: op1_11_inv06 = 1;
    33: op1_11_inv06 = 1;
    34: op1_11_inv06 = 1;
    35: op1_11_inv06 = 1;
    36: op1_11_inv06 = 1;
    43: op1_11_inv06 = 1;
    48: op1_11_inv06 = 1;
    49: op1_11_inv06 = 1;
    50: op1_11_inv06 = 1;
    51: op1_11_inv06 = 1;
    53: op1_11_inv06 = 1;
    57: op1_11_inv06 = 1;
    61: op1_11_inv06 = 1;
    64: op1_11_inv06 = 1;
    65: op1_11_inv06 = 1;
    71: op1_11_inv06 = 1;
    74: op1_11_inv06 = 1;
    77: op1_11_inv06 = 1;
    80: op1_11_inv06 = 1;
    81: op1_11_inv06 = 1;
    83: op1_11_inv06 = 1;
    85: op1_11_inv06 = 1;
    87: op1_11_inv06 = 1;
    88: op1_11_inv06 = 1;
    89: op1_11_inv06 = 1;
    91: op1_11_inv06 = 1;
    92: op1_11_inv06 = 1;
    93: op1_11_inv06 = 1;
    default: op1_11_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in07 = reg_0052;
    5: op1_11_in07 = reg_0101;
    6: op1_11_in07 = reg_0053;
    7: op1_11_in07 = reg_0713;
    8: op1_11_in07 = reg_0357;
    9: op1_11_in07 = reg_0476;
    10: op1_11_in07 = reg_0535;
    11: op1_11_in07 = reg_0676;
    83: op1_11_in07 = reg_0676;
    12: op1_11_in07 = reg_0483;
    13: op1_11_in07 = imem07_in[103:100];
    14: op1_11_in07 = reg_0689;
    60: op1_11_in07 = reg_0689;
    15: op1_11_in07 = reg_0369;
    66: op1_11_in07 = reg_0369;
    16: op1_11_in07 = reg_0152;
    17: op1_11_in07 = reg_0374;
    24: op1_11_in07 = reg_0374;
    18: op1_11_in07 = reg_0790;
    19: op1_11_in07 = reg_0312;
    20: op1_11_in07 = reg_0816;
    21: op1_11_in07 = reg_0238;
    22: op1_11_in07 = reg_0355;
    23: op1_11_in07 = reg_0104;
    25: op1_11_in07 = reg_0480;
    26: op1_11_in07 = reg_0780;
    27: op1_11_in07 = reg_0791;
    28: op1_11_in07 = reg_0652;
    29: op1_11_in07 = imem03_in[123:120];
    30: op1_11_in07 = imem06_in[51:48];
    31: op1_11_in07 = reg_0687;
    32: op1_11_in07 = reg_0672;
    33: op1_11_in07 = reg_0800;
    34: op1_11_in07 = reg_0162;
    35: op1_11_in07 = reg_0183;
    36: op1_11_in07 = reg_0468;
    38: op1_11_in07 = reg_0356;
    39: op1_11_in07 = reg_0755;
    40: op1_11_in07 = reg_0801;
    42: op1_11_in07 = reg_0684;
    43: op1_11_in07 = reg_0661;
    44: op1_11_in07 = reg_0624;
    45: op1_11_in07 = reg_0174;
    73: op1_11_in07 = reg_0174;
    46: op1_11_in07 = reg_0548;
    47: op1_11_in07 = reg_0140;
    48: op1_11_in07 = reg_0710;
    49: op1_11_in07 = reg_0585;
    50: op1_11_in07 = reg_0806;
    51: op1_11_in07 = reg_0107;
    52: op1_11_in07 = imem04_in[35:32];
    53: op1_11_in07 = reg_0383;
    54: op1_11_in07 = reg_0748;
    56: op1_11_in07 = reg_0620;
    57: op1_11_in07 = imem07_in[7:4];
    61: op1_11_in07 = reg_0650;
    62: op1_11_in07 = reg_0786;
    63: op1_11_in07 = reg_0102;
    64: op1_11_in07 = reg_0821;
    65: op1_11_in07 = reg_0709;
    67: op1_11_in07 = imem02_in[35:32];
    68: op1_11_in07 = reg_0588;
    69: op1_11_in07 = reg_0184;
    70: op1_11_in07 = reg_0452;
    71: op1_11_in07 = reg_0231;
    74: op1_11_in07 = reg_0691;
    75: op1_11_in07 = reg_0642;
    76: op1_11_in07 = reg_0015;
    77: op1_11_in07 = reg_0496;
    78: op1_11_in07 = reg_0147;
    80: op1_11_in07 = reg_0694;
    81: op1_11_in07 = reg_0721;
    82: op1_11_in07 = reg_0779;
    84: op1_11_in07 = imem07_in[59:56];
    85: op1_11_in07 = reg_0693;
    86: op1_11_in07 = imem04_in[83:80];
    87: op1_11_in07 = reg_0664;
    88: op1_11_in07 = imem04_in[51:48];
    89: op1_11_in07 = reg_0613;
    90: op1_11_in07 = reg_0291;
    91: op1_11_in07 = reg_0145;
    92: op1_11_in07 = imem02_in[83:80];
    93: op1_11_in07 = imem02_in[99:96];
    94: op1_11_in07 = reg_0361;
    95: op1_11_in07 = reg_0256;
    default: op1_11_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_11_inv07 = 1;
    8: op1_11_inv07 = 1;
    10: op1_11_inv07 = 1;
    13: op1_11_inv07 = 1;
    16: op1_11_inv07 = 1;
    17: op1_11_inv07 = 1;
    21: op1_11_inv07 = 1;
    24: op1_11_inv07 = 1;
    26: op1_11_inv07 = 1;
    27: op1_11_inv07 = 1;
    28: op1_11_inv07 = 1;
    30: op1_11_inv07 = 1;
    32: op1_11_inv07 = 1;
    35: op1_11_inv07 = 1;
    36: op1_11_inv07 = 1;
    38: op1_11_inv07 = 1;
    39: op1_11_inv07 = 1;
    40: op1_11_inv07 = 1;
    44: op1_11_inv07 = 1;
    45: op1_11_inv07 = 1;
    51: op1_11_inv07 = 1;
    52: op1_11_inv07 = 1;
    53: op1_11_inv07 = 1;
    56: op1_11_inv07 = 1;
    62: op1_11_inv07 = 1;
    64: op1_11_inv07 = 1;
    65: op1_11_inv07 = 1;
    67: op1_11_inv07 = 1;
    68: op1_11_inv07 = 1;
    71: op1_11_inv07 = 1;
    81: op1_11_inv07 = 1;
    82: op1_11_inv07 = 1;
    83: op1_11_inv07 = 1;
    85: op1_11_inv07 = 1;
    87: op1_11_inv07 = 1;
    88: op1_11_inv07 = 1;
    92: op1_11_inv07 = 1;
    93: op1_11_inv07 = 1;
    94: op1_11_inv07 = 1;
    95: op1_11_inv07 = 1;
    default: op1_11_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in08 = reg_0084;
    5: op1_11_in08 = reg_0121;
    6: op1_11_in08 = reg_0048;
    7: op1_11_in08 = reg_0423;
    8: op1_11_in08 = reg_0318;
    9: op1_11_in08 = reg_0473;
    10: op1_11_in08 = reg_0540;
    11: op1_11_in08 = reg_0689;
    12: op1_11_in08 = reg_0781;
    13: op1_11_in08 = reg_0716;
    14: op1_11_in08 = reg_0692;
    31: op1_11_in08 = reg_0692;
    15: op1_11_in08 = reg_0322;
    16: op1_11_in08 = reg_0142;
    17: op1_11_in08 = reg_0807;
    18: op1_11_in08 = reg_0737;
    19: op1_11_in08 = reg_0374;
    20: op1_11_in08 = reg_0750;
    21: op1_11_in08 = reg_0243;
    22: op1_11_in08 = reg_0094;
    23: op1_11_in08 = reg_0114;
    24: op1_11_in08 = reg_0001;
    25: op1_11_in08 = reg_0203;
    26: op1_11_in08 = reg_0495;
    27: op1_11_in08 = reg_0483;
    28: op1_11_in08 = reg_0349;
    29: op1_11_in08 = imem03_in[127:124];
    30: op1_11_in08 = imem06_in[91:88];
    32: op1_11_in08 = reg_0694;
    33: op1_11_in08 = reg_0802;
    34: op1_11_in08 = reg_0160;
    35: op1_11_in08 = reg_0168;
    36: op1_11_in08 = reg_0189;
    38: op1_11_in08 = reg_0346;
    39: op1_11_in08 = reg_0568;
    40: op1_11_in08 = reg_0805;
    42: op1_11_in08 = reg_0690;
    43: op1_11_in08 = reg_0665;
    44: op1_11_in08 = reg_0218;
    45: op1_11_in08 = reg_0180;
    46: op1_11_in08 = reg_0336;
    47: op1_11_in08 = reg_0131;
    48: op1_11_in08 = reg_0712;
    49: op1_11_in08 = reg_0515;
    50: op1_11_in08 = reg_0004;
    51: op1_11_in08 = reg_0348;
    52: op1_11_in08 = imem04_in[55:52];
    53: op1_11_in08 = reg_0397;
    54: op1_11_in08 = reg_0403;
    56: op1_11_in08 = reg_0819;
    57: op1_11_in08 = imem07_in[19:16];
    60: op1_11_in08 = reg_0477;
    61: op1_11_in08 = reg_0584;
    62: op1_11_in08 = reg_0489;
    63: op1_11_in08 = reg_0276;
    64: op1_11_in08 = reg_0583;
    65: op1_11_in08 = reg_0436;
    66: op1_11_in08 = reg_0613;
    67: op1_11_in08 = imem02_in[47:44];
    68: op1_11_in08 = reg_0509;
    70: op1_11_in08 = reg_0478;
    71: op1_11_in08 = reg_0742;
    73: op1_11_in08 = reg_0181;
    74: op1_11_in08 = reg_0688;
    75: op1_11_in08 = reg_0141;
    76: op1_11_in08 = imem04_in[31:28];
    77: op1_11_in08 = reg_0747;
    78: op1_11_in08 = reg_0148;
    80: op1_11_in08 = reg_0758;
    81: op1_11_in08 = reg_0167;
    82: op1_11_in08 = reg_0223;
    83: op1_11_in08 = reg_0126;
    84: op1_11_in08 = imem07_in[71:68];
    85: op1_11_in08 = reg_0492;
    86: op1_11_in08 = reg_0542;
    87: op1_11_in08 = imem07_in[7:4];
    88: op1_11_in08 = imem04_in[59:56];
    89: op1_11_in08 = reg_0654;
    90: op1_11_in08 = reg_0354;
    91: op1_11_in08 = reg_0451;
    92: op1_11_in08 = imem02_in[91:88];
    93: op1_11_in08 = imem02_in[103:100];
    94: op1_11_in08 = reg_0356;
    95: op1_11_in08 = reg_0587;
    default: op1_11_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv08 = 1;
    6: op1_11_inv08 = 1;
    8: op1_11_inv08 = 1;
    10: op1_11_inv08 = 1;
    12: op1_11_inv08 = 1;
    15: op1_11_inv08 = 1;
    16: op1_11_inv08 = 1;
    17: op1_11_inv08 = 1;
    18: op1_11_inv08 = 1;
    19: op1_11_inv08 = 1;
    22: op1_11_inv08 = 1;
    24: op1_11_inv08 = 1;
    25: op1_11_inv08 = 1;
    28: op1_11_inv08 = 1;
    33: op1_11_inv08 = 1;
    34: op1_11_inv08 = 1;
    35: op1_11_inv08 = 1;
    39: op1_11_inv08 = 1;
    42: op1_11_inv08 = 1;
    44: op1_11_inv08 = 1;
    46: op1_11_inv08 = 1;
    48: op1_11_inv08 = 1;
    49: op1_11_inv08 = 1;
    52: op1_11_inv08 = 1;
    53: op1_11_inv08 = 1;
    60: op1_11_inv08 = 1;
    66: op1_11_inv08 = 1;
    67: op1_11_inv08 = 1;
    68: op1_11_inv08 = 1;
    71: op1_11_inv08 = 1;
    73: op1_11_inv08 = 1;
    76: op1_11_inv08 = 1;
    81: op1_11_inv08 = 1;
    84: op1_11_inv08 = 1;
    85: op1_11_inv08 = 1;
    87: op1_11_inv08 = 1;
    88: op1_11_inv08 = 1;
    89: op1_11_inv08 = 1;
    95: op1_11_inv08 = 1;
    default: op1_11_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in09 = reg_0094;
    5: op1_11_in09 = reg_0110;
    6: op1_11_in09 = reg_0074;
    7: op1_11_in09 = reg_0175;
    8: op1_11_in09 = reg_0330;
    9: op1_11_in09 = reg_0467;
    10: op1_11_in09 = reg_0301;
    11: op1_11_in09 = reg_0686;
    12: op1_11_in09 = reg_0488;
    13: op1_11_in09 = reg_0731;
    14: op1_11_in09 = reg_0463;
    31: op1_11_in09 = reg_0463;
    15: op1_11_in09 = reg_0323;
    16: op1_11_in09 = reg_0154;
    17: op1_11_in09 = reg_0804;
    18: op1_11_in09 = reg_0735;
    19: op1_11_in09 = reg_0001;
    20: op1_11_in09 = imem07_in[11:8];
    21: op1_11_in09 = reg_0508;
    22: op1_11_in09 = imem03_in[7:4];
    23: op1_11_in09 = reg_0101;
    24: op1_11_in09 = reg_0801;
    25: op1_11_in09 = reg_0193;
    26: op1_11_in09 = reg_0783;
    27: op1_11_in09 = reg_0788;
    28: op1_11_in09 = reg_0344;
    29: op1_11_in09 = reg_0589;
    30: op1_11_in09 = imem06_in[107:104];
    32: op1_11_in09 = reg_0676;
    33: op1_11_in09 = reg_0016;
    34: op1_11_in09 = reg_0183;
    36: op1_11_in09 = imem01_in[3:0];
    38: op1_11_in09 = reg_0092;
    39: op1_11_in09 = reg_0517;
    40: op1_11_in09 = imem04_in[27:24];
    42: op1_11_in09 = reg_0465;
    43: op1_11_in09 = reg_0667;
    44: op1_11_in09 = reg_0606;
    45: op1_11_in09 = reg_0161;
    73: op1_11_in09 = reg_0161;
    46: op1_11_in09 = reg_0364;
    47: op1_11_in09 = imem06_in[7:4];
    48: op1_11_in09 = reg_0708;
    49: op1_11_in09 = reg_0549;
    50: op1_11_in09 = imem04_in[39:36];
    77: op1_11_in09 = imem04_in[39:36];
    51: op1_11_in09 = reg_0108;
    52: op1_11_in09 = imem04_in[127:124];
    53: op1_11_in09 = reg_0396;
    68: op1_11_in09 = reg_0396;
    54: op1_11_in09 = reg_0404;
    90: op1_11_in09 = reg_0404;
    56: op1_11_in09 = reg_0632;
    57: op1_11_in09 = imem07_in[39:36];
    60: op1_11_in09 = reg_0469;
    61: op1_11_in09 = reg_0639;
    62: op1_11_in09 = reg_0486;
    63: op1_11_in09 = reg_0307;
    64: op1_11_in09 = reg_0515;
    65: op1_11_in09 = reg_0447;
    66: op1_11_in09 = reg_0654;
    67: op1_11_in09 = imem02_in[79:76];
    70: op1_11_in09 = reg_0208;
    71: op1_11_in09 = reg_0227;
    74: op1_11_in09 = reg_0462;
    75: op1_11_in09 = reg_0139;
    76: op1_11_in09 = imem04_in[51:48];
    78: op1_11_in09 = reg_0149;
    80: op1_11_in09 = reg_0680;
    81: op1_11_in09 = reg_0166;
    82: op1_11_in09 = reg_0062;
    83: op1_11_in09 = reg_0678;
    84: op1_11_in09 = imem07_in[91:88];
    85: op1_11_in09 = reg_0658;
    86: op1_11_in09 = reg_0534;
    87: op1_11_in09 = imem07_in[15:12];
    88: op1_11_in09 = imem04_in[63:60];
    89: op1_11_in09 = reg_0242;
    91: op1_11_in09 = reg_0464;
    92: op1_11_in09 = imem02_in[99:96];
    93: op1_11_in09 = imem02_in[115:112];
    94: op1_11_in09 = reg_0360;
    95: op1_11_in09 = reg_0362;
    default: op1_11_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv09 = 1;
    10: op1_11_inv09 = 1;
    11: op1_11_inv09 = 1;
    12: op1_11_inv09 = 1;
    13: op1_11_inv09 = 1;
    14: op1_11_inv09 = 1;
    15: op1_11_inv09 = 1;
    18: op1_11_inv09 = 1;
    19: op1_11_inv09 = 1;
    20: op1_11_inv09 = 1;
    23: op1_11_inv09 = 1;
    27: op1_11_inv09 = 1;
    29: op1_11_inv09 = 1;
    36: op1_11_inv09 = 1;
    38: op1_11_inv09 = 1;
    39: op1_11_inv09 = 1;
    42: op1_11_inv09 = 1;
    43: op1_11_inv09 = 1;
    45: op1_11_inv09 = 1;
    48: op1_11_inv09 = 1;
    51: op1_11_inv09 = 1;
    52: op1_11_inv09 = 1;
    54: op1_11_inv09 = 1;
    56: op1_11_inv09 = 1;
    57: op1_11_inv09 = 1;
    60: op1_11_inv09 = 1;
    62: op1_11_inv09 = 1;
    63: op1_11_inv09 = 1;
    65: op1_11_inv09 = 1;
    66: op1_11_inv09 = 1;
    74: op1_11_inv09 = 1;
    75: op1_11_inv09 = 1;
    76: op1_11_inv09 = 1;
    80: op1_11_inv09 = 1;
    81: op1_11_inv09 = 1;
    83: op1_11_inv09 = 1;
    84: op1_11_inv09 = 1;
    85: op1_11_inv09 = 1;
    86: op1_11_inv09 = 1;
    87: op1_11_inv09 = 1;
    89: op1_11_inv09 = 1;
    92: op1_11_inv09 = 1;
    93: op1_11_inv09 = 1;
    default: op1_11_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in10 = imem03_in[27:24];
    5: op1_11_in10 = imem02_in[39:36];
    6: op1_11_in10 = imem05_in[67:64];
    7: op1_11_in10 = reg_0180;
    8: op1_11_in10 = reg_0314;
    9: op1_11_in10 = reg_0470;
    74: op1_11_in10 = reg_0470;
    10: op1_11_in10 = reg_0300;
    11: op1_11_in10 = reg_0679;
    12: op1_11_in10 = reg_0491;
    27: op1_11_in10 = reg_0491;
    13: op1_11_in10 = reg_0702;
    14: op1_11_in10 = reg_0450;
    15: op1_11_in10 = reg_0002;
    19: op1_11_in10 = reg_0002;
    16: op1_11_in10 = reg_0143;
    17: op1_11_in10 = reg_0800;
    24: op1_11_in10 = reg_0800;
    18: op1_11_in10 = reg_0733;
    20: op1_11_in10 = imem07_in[19:16];
    21: op1_11_in10 = reg_0111;
    22: op1_11_in10 = imem03_in[15:12];
    23: op1_11_in10 = reg_0121;
    25: op1_11_in10 = reg_0201;
    26: op1_11_in10 = reg_0790;
    28: op1_11_in10 = reg_0345;
    29: op1_11_in10 = reg_0600;
    30: op1_11_in10 = reg_0605;
    31: op1_11_in10 = reg_0465;
    32: op1_11_in10 = reg_0670;
    33: op1_11_in10 = imem04_in[59:56];
    34: op1_11_in10 = reg_0177;
    73: op1_11_in10 = reg_0177;
    36: op1_11_in10 = imem01_in[11:8];
    38: op1_11_in10 = reg_0080;
    39: op1_11_in10 = reg_0003;
    40: op1_11_in10 = imem04_in[39:36];
    42: op1_11_in10 = reg_0457;
    43: op1_11_in10 = reg_0663;
    44: op1_11_in10 = reg_0293;
    90: op1_11_in10 = reg_0293;
    45: op1_11_in10 = reg_0167;
    46: op1_11_in10 = reg_0354;
    47: op1_11_in10 = imem06_in[11:8];
    48: op1_11_in10 = reg_0705;
    49: op1_11_in10 = reg_0323;
    50: op1_11_in10 = imem04_in[63:60];
    51: op1_11_in10 = reg_0230;
    52: op1_11_in10 = reg_0560;
    53: op1_11_in10 = reg_0804;
    54: op1_11_in10 = reg_0614;
    56: op1_11_in10 = imem07_in[7:4];
    57: op1_11_in10 = imem07_in[47:44];
    60: op1_11_in10 = reg_0456;
    61: op1_11_in10 = reg_0548;
    62: op1_11_in10 = reg_0066;
    63: op1_11_in10 = reg_0277;
    64: op1_11_in10 = reg_0534;
    65: op1_11_in10 = reg_0084;
    66: op1_11_in10 = reg_0377;
    67: op1_11_in10 = imem02_in[87:84];
    68: op1_11_in10 = reg_0811;
    70: op1_11_in10 = reg_0187;
    71: op1_11_in10 = reg_0499;
    75: op1_11_in10 = reg_0704;
    76: op1_11_in10 = imem04_in[55:52];
    77: op1_11_in10 = imem04_in[43:40];
    78: op1_11_in10 = reg_0785;
    80: op1_11_in10 = reg_0453;
    81: op1_11_in10 = reg_0708;
    82: op1_11_in10 = reg_0585;
    83: op1_11_in10 = reg_0532;
    84: op1_11_in10 = imem07_in[111:108];
    85: op1_11_in10 = reg_0758;
    86: op1_11_in10 = reg_0536;
    87: op1_11_in10 = imem07_in[23:20];
    88: op1_11_in10 = imem04_in[71:68];
    89: op1_11_in10 = reg_0515;
    91: op1_11_in10 = reg_0191;
    92: op1_11_in10 = imem02_in[119:116];
    93: op1_11_in10 = reg_0081;
    94: op1_11_in10 = reg_0353;
    95: op1_11_in10 = reg_0341;
    default: op1_11_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv10 = 1;
    8: op1_11_inv10 = 1;
    13: op1_11_inv10 = 1;
    15: op1_11_inv10 = 1;
    17: op1_11_inv10 = 1;
    18: op1_11_inv10 = 1;
    19: op1_11_inv10 = 1;
    25: op1_11_inv10 = 1;
    27: op1_11_inv10 = 1;
    28: op1_11_inv10 = 1;
    29: op1_11_inv10 = 1;
    32: op1_11_inv10 = 1;
    33: op1_11_inv10 = 1;
    36: op1_11_inv10 = 1;
    39: op1_11_inv10 = 1;
    42: op1_11_inv10 = 1;
    43: op1_11_inv10 = 1;
    44: op1_11_inv10 = 1;
    45: op1_11_inv10 = 1;
    47: op1_11_inv10 = 1;
    49: op1_11_inv10 = 1;
    50: op1_11_inv10 = 1;
    51: op1_11_inv10 = 1;
    56: op1_11_inv10 = 1;
    57: op1_11_inv10 = 1;
    62: op1_11_inv10 = 1;
    63: op1_11_inv10 = 1;
    67: op1_11_inv10 = 1;
    70: op1_11_inv10 = 1;
    71: op1_11_inv10 = 1;
    73: op1_11_inv10 = 1;
    74: op1_11_inv10 = 1;
    82: op1_11_inv10 = 1;
    85: op1_11_inv10 = 1;
    86: op1_11_inv10 = 1;
    87: op1_11_inv10 = 1;
    92: op1_11_inv10 = 1;
    95: op1_11_inv10 = 1;
    default: op1_11_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in11 = imem03_in[47:44];
    5: op1_11_in11 = imem02_in[71:68];
    6: op1_11_in11 = imem05_in[79:76];
    7: op1_11_in11 = reg_0161;
    8: op1_11_in11 = reg_0347;
    9: op1_11_in11 = reg_0479;
    10: op1_11_in11 = reg_0302;
    11: op1_11_in11 = reg_0453;
    12: op1_11_in11 = reg_0793;
    13: op1_11_in11 = reg_0729;
    14: op1_11_in11 = reg_0451;
    15: op1_11_in11 = reg_0015;
    17: op1_11_in11 = reg_0015;
    16: op1_11_in11 = reg_0144;
    18: op1_11_in11 = reg_0272;
    19: op1_11_in11 = reg_0008;
    20: op1_11_in11 = imem07_in[35:32];
    21: op1_11_in11 = reg_0119;
    22: op1_11_in11 = imem03_in[19:16];
    23: op1_11_in11 = reg_0110;
    24: op1_11_in11 = reg_0016;
    25: op1_11_in11 = reg_0190;
    26: op1_11_in11 = reg_0485;
    61: op1_11_in11 = reg_0485;
    75: op1_11_in11 = reg_0485;
    27: op1_11_in11 = reg_0795;
    28: op1_11_in11 = reg_0348;
    29: op1_11_in11 = reg_0597;
    30: op1_11_in11 = reg_0626;
    31: op1_11_in11 = reg_0457;
    32: op1_11_in11 = reg_0687;
    33: op1_11_in11 = imem04_in[79:76];
    36: op1_11_in11 = imem01_in[79:76];
    38: op1_11_in11 = reg_0769;
    39: op1_11_in11 = reg_0801;
    68: op1_11_in11 = reg_0801;
    40: op1_11_in11 = imem04_in[51:48];
    42: op1_11_in11 = reg_0481;
    43: op1_11_in11 = reg_0320;
    44: op1_11_in11 = reg_0612;
    46: op1_11_in11 = reg_0359;
    47: op1_11_in11 = imem06_in[23:20];
    48: op1_11_in11 = reg_0718;
    49: op1_11_in11 = reg_0798;
    50: op1_11_in11 = imem04_in[87:84];
    51: op1_11_in11 = reg_0346;
    52: op1_11_in11 = reg_0552;
    53: op1_11_in11 = reg_0800;
    54: op1_11_in11 = reg_0031;
    56: op1_11_in11 = imem07_in[31:28];
    57: op1_11_in11 = imem07_in[63:60];
    60: op1_11_in11 = reg_0191;
    62: op1_11_in11 = reg_0257;
    63: op1_11_in11 = reg_0145;
    64: op1_11_in11 = reg_0700;
    65: op1_11_in11 = reg_0268;
    66: op1_11_in11 = reg_0405;
    67: op1_11_in11 = imem02_in[91:88];
    70: op1_11_in11 = reg_0203;
    71: op1_11_in11 = reg_0489;
    73: op1_11_in11 = reg_0178;
    74: op1_11_in11 = reg_0468;
    76: op1_11_in11 = reg_0262;
    77: op1_11_in11 = imem04_in[47:44];
    78: op1_11_in11 = reg_0781;
    80: op1_11_in11 = reg_0454;
    81: op1_11_in11 = reg_0713;
    82: op1_11_in11 = reg_0065;
    83: op1_11_in11 = imem02_in[19:16];
    84: op1_11_in11 = reg_0721;
    85: op1_11_in11 = reg_0494;
    86: op1_11_in11 = reg_0516;
    87: op1_11_in11 = imem07_in[27:24];
    88: op1_11_in11 = imem04_in[75:72];
    89: op1_11_in11 = reg_0163;
    90: op1_11_in11 = reg_0039;
    91: op1_11_in11 = reg_0194;
    92: op1_11_in11 = reg_0057;
    93: op1_11_in11 = reg_0264;
    94: op1_11_in11 = reg_0343;
    95: op1_11_in11 = reg_0565;
    default: op1_11_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv11 = 1;
    5: op1_11_inv11 = 1;
    6: op1_11_inv11 = 1;
    7: op1_11_inv11 = 1;
    9: op1_11_inv11 = 1;
    15: op1_11_inv11 = 1;
    17: op1_11_inv11 = 1;
    19: op1_11_inv11 = 1;
    21: op1_11_inv11 = 1;
    23: op1_11_inv11 = 1;
    24: op1_11_inv11 = 1;
    25: op1_11_inv11 = 1;
    27: op1_11_inv11 = 1;
    28: op1_11_inv11 = 1;
    30: op1_11_inv11 = 1;
    33: op1_11_inv11 = 1;
    36: op1_11_inv11 = 1;
    42: op1_11_inv11 = 1;
    44: op1_11_inv11 = 1;
    46: op1_11_inv11 = 1;
    47: op1_11_inv11 = 1;
    48: op1_11_inv11 = 1;
    49: op1_11_inv11 = 1;
    52: op1_11_inv11 = 1;
    62: op1_11_inv11 = 1;
    63: op1_11_inv11 = 1;
    64: op1_11_inv11 = 1;
    65: op1_11_inv11 = 1;
    70: op1_11_inv11 = 1;
    73: op1_11_inv11 = 1;
    75: op1_11_inv11 = 1;
    77: op1_11_inv11 = 1;
    80: op1_11_inv11 = 1;
    81: op1_11_inv11 = 1;
    82: op1_11_inv11 = 1;
    85: op1_11_inv11 = 1;
    87: op1_11_inv11 = 1;
    91: op1_11_inv11 = 1;
    94: op1_11_inv11 = 1;
    default: op1_11_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in12 = imem03_in[111:108];
    5: op1_11_in12 = imem02_in[111:108];
    67: op1_11_in12 = imem02_in[111:108];
    6: op1_11_in12 = imem05_in[87:84];
    7: op1_11_in12 = reg_0167;
    8: op1_11_in12 = reg_0092;
    9: op1_11_in12 = reg_0459;
    10: op1_11_in12 = reg_0293;
    11: op1_11_in12 = reg_0469;
    12: op1_11_in12 = reg_0495;
    13: op1_11_in12 = reg_0707;
    14: op1_11_in12 = reg_0455;
    15: op1_11_in12 = reg_0010;
    16: op1_11_in12 = imem06_in[19:16];
    17: op1_11_in12 = reg_0809;
    24: op1_11_in12 = reg_0809;
    18: op1_11_in12 = reg_0744;
    19: op1_11_in12 = imem04_in[15:12];
    20: op1_11_in12 = imem07_in[51:48];
    21: op1_11_in12 = reg_0102;
    22: op1_11_in12 = imem03_in[71:68];
    23: op1_11_in12 = imem02_in[11:8];
    25: op1_11_in12 = reg_0195;
    26: op1_11_in12 = reg_0225;
    27: op1_11_in12 = reg_0793;
    28: op1_11_in12 = reg_0363;
    29: op1_11_in12 = reg_0590;
    30: op1_11_in12 = reg_0632;
    31: op1_11_in12 = reg_0461;
    32: op1_11_in12 = reg_0463;
    33: op1_11_in12 = imem04_in[115:112];
    36: op1_11_in12 = imem01_in[127:124];
    38: op1_11_in12 = reg_0540;
    39: op1_11_in12 = reg_0004;
    40: op1_11_in12 = imem04_in[79:76];
    42: op1_11_in12 = reg_0201;
    43: op1_11_in12 = reg_0353;
    44: op1_11_in12 = reg_0318;
    46: op1_11_in12 = reg_0348;
    47: op1_11_in12 = imem06_in[55:52];
    48: op1_11_in12 = reg_0701;
    49: op1_11_in12 = reg_0490;
    50: op1_11_in12 = reg_0303;
    51: op1_11_in12 = reg_0548;
    52: op1_11_in12 = reg_0554;
    53: op1_11_in12 = reg_0015;
    54: op1_11_in12 = reg_0037;
    56: op1_11_in12 = imem07_in[67:64];
    57: op1_11_in12 = imem07_in[103:100];
    60: op1_11_in12 = reg_0210;
    61: op1_11_in12 = reg_0358;
    75: op1_11_in12 = reg_0358;
    62: op1_11_in12 = reg_0101;
    63: op1_11_in12 = reg_0136;
    64: op1_11_in12 = reg_0794;
    65: op1_11_in12 = reg_0174;
    66: op1_11_in12 = reg_0775;
    68: op1_11_in12 = reg_0016;
    70: op1_11_in12 = reg_0194;
    71: op1_11_in12 = reg_0326;
    73: op1_11_in12 = reg_0158;
    74: op1_11_in12 = reg_0478;
    76: op1_11_in12 = reg_0544;
    77: op1_11_in12 = reg_0552;
    78: op1_11_in12 = reg_0150;
    80: op1_11_in12 = reg_0450;
    81: op1_11_in12 = reg_0711;
    82: op1_11_in12 = reg_0069;
    83: op1_11_in12 = imem02_in[43:40];
    84: op1_11_in12 = reg_0382;
    85: op1_11_in12 = reg_0699;
    86: op1_11_in12 = reg_0615;
    87: op1_11_in12 = imem07_in[87:84];
    88: op1_11_in12 = imem04_in[87:84];
    89: op1_11_in12 = reg_0700;
    90: op1_11_in12 = reg_0578;
    91: op1_11_in12 = reg_0212;
    92: op1_11_in12 = reg_0541;
    93: op1_11_in12 = reg_0498;
    94: op1_11_in12 = reg_0030;
    95: op1_11_in12 = reg_0361;
    default: op1_11_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv12 = 1;
    7: op1_11_inv12 = 1;
    8: op1_11_inv12 = 1;
    9: op1_11_inv12 = 1;
    10: op1_11_inv12 = 1;
    16: op1_11_inv12 = 1;
    17: op1_11_inv12 = 1;
    24: op1_11_inv12 = 1;
    26: op1_11_inv12 = 1;
    27: op1_11_inv12 = 1;
    28: op1_11_inv12 = 1;
    30: op1_11_inv12 = 1;
    31: op1_11_inv12 = 1;
    38: op1_11_inv12 = 1;
    42: op1_11_inv12 = 1;
    46: op1_11_inv12 = 1;
    47: op1_11_inv12 = 1;
    49: op1_11_inv12 = 1;
    50: op1_11_inv12 = 1;
    51: op1_11_inv12 = 1;
    52: op1_11_inv12 = 1;
    62: op1_11_inv12 = 1;
    63: op1_11_inv12 = 1;
    64: op1_11_inv12 = 1;
    65: op1_11_inv12 = 1;
    66: op1_11_inv12 = 1;
    68: op1_11_inv12 = 1;
    70: op1_11_inv12 = 1;
    73: op1_11_inv12 = 1;
    74: op1_11_inv12 = 1;
    75: op1_11_inv12 = 1;
    76: op1_11_inv12 = 1;
    78: op1_11_inv12 = 1;
    81: op1_11_inv12 = 1;
    82: op1_11_inv12 = 1;
    83: op1_11_inv12 = 1;
    92: op1_11_inv12 = 1;
    94: op1_11_inv12 = 1;
    default: op1_11_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in13 = reg_0586;
    5: op1_11_in13 = reg_0655;
    6: op1_11_in13 = imem05_in[107:104];
    7: op1_11_in13 = reg_0163;
    8: op1_11_in13 = reg_0090;
    9: op1_11_in13 = reg_0210;
    10: op1_11_in13 = reg_0296;
    11: op1_11_in13 = reg_0473;
    12: op1_11_in13 = reg_0787;
    13: op1_11_in13 = reg_0430;
    14: op1_11_in13 = reg_0457;
    15: op1_11_in13 = imem04_in[15:12];
    16: op1_11_in13 = imem06_in[63:60];
    17: op1_11_in13 = reg_0052;
    18: op1_11_in13 = reg_0734;
    19: op1_11_in13 = imem04_in[19:16];
    20: op1_11_in13 = imem07_in[107:104];
    21: op1_11_in13 = reg_0126;
    22: op1_11_in13 = imem03_in[119:116];
    23: op1_11_in13 = imem02_in[27:24];
    24: op1_11_in13 = imem04_in[39:36];
    25: op1_11_in13 = reg_0199;
    26: op1_11_in13 = reg_0735;
    27: op1_11_in13 = reg_0495;
    28: op1_11_in13 = reg_0324;
    29: op1_11_in13 = reg_0573;
    30: op1_11_in13 = reg_0627;
    31: op1_11_in13 = reg_0472;
    32: op1_11_in13 = reg_0477;
    85: op1_11_in13 = reg_0477;
    33: op1_11_in13 = imem04_in[119:116];
    36: op1_11_in13 = reg_0514;
    38: op1_11_in13 = reg_0498;
    39: op1_11_in13 = imem04_in[27:24];
    40: op1_11_in13 = imem04_in[83:80];
    42: op1_11_in13 = imem01_in[83:80];
    43: op1_11_in13 = reg_0342;
    44: op1_11_in13 = reg_0377;
    46: op1_11_in13 = reg_0365;
    47: op1_11_in13 = reg_0289;
    48: op1_11_in13 = reg_0706;
    49: op1_11_in13 = reg_0789;
    50: op1_11_in13 = reg_0631;
    51: op1_11_in13 = imem02_in[7:4];
    52: op1_11_in13 = reg_0523;
    53: op1_11_in13 = reg_0809;
    54: op1_11_in13 = reg_0818;
    56: op1_11_in13 = imem07_in[75:72];
    57: op1_11_in13 = reg_0730;
    60: op1_11_in13 = reg_0187;
    61: op1_11_in13 = reg_0362;
    62: op1_11_in13 = reg_0148;
    63: op1_11_in13 = reg_0133;
    64: op1_11_in13 = reg_0368;
    65: op1_11_in13 = reg_0175;
    66: op1_11_in13 = reg_0620;
    89: op1_11_in13 = reg_0620;
    67: op1_11_in13 = reg_0785;
    68: op1_11_in13 = reg_0810;
    70: op1_11_in13 = reg_0202;
    71: op1_11_in13 = reg_0249;
    74: op1_11_in13 = reg_0200;
    75: op1_11_in13 = reg_0565;
    76: op1_11_in13 = reg_0537;
    77: op1_11_in13 = reg_0087;
    78: op1_11_in13 = reg_0761;
    80: op1_11_in13 = reg_0455;
    81: op1_11_in13 = reg_0724;
    82: op1_11_in13 = reg_0311;
    83: op1_11_in13 = imem02_in[51:48];
    84: op1_11_in13 = reg_0725;
    86: op1_11_in13 = reg_0503;
    87: op1_11_in13 = reg_0728;
    88: op1_11_in13 = imem04_in[95:92];
    90: op1_11_in13 = reg_0408;
    91: op1_11_in13 = reg_0205;
    92: op1_11_in13 = reg_0533;
    93: op1_11_in13 = reg_0587;
    94: op1_11_in13 = reg_0043;
    95: op1_11_in13 = reg_0527;
    default: op1_11_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv13 = 1;
    6: op1_11_inv13 = 1;
    8: op1_11_inv13 = 1;
    9: op1_11_inv13 = 1;
    13: op1_11_inv13 = 1;
    14: op1_11_inv13 = 1;
    17: op1_11_inv13 = 1;
    20: op1_11_inv13 = 1;
    21: op1_11_inv13 = 1;
    22: op1_11_inv13 = 1;
    23: op1_11_inv13 = 1;
    24: op1_11_inv13 = 1;
    26: op1_11_inv13 = 1;
    28: op1_11_inv13 = 1;
    31: op1_11_inv13 = 1;
    33: op1_11_inv13 = 1;
    39: op1_11_inv13 = 1;
    40: op1_11_inv13 = 1;
    42: op1_11_inv13 = 1;
    48: op1_11_inv13 = 1;
    50: op1_11_inv13 = 1;
    51: op1_11_inv13 = 1;
    52: op1_11_inv13 = 1;
    53: op1_11_inv13 = 1;
    56: op1_11_inv13 = 1;
    57: op1_11_inv13 = 1;
    61: op1_11_inv13 = 1;
    67: op1_11_inv13 = 1;
    68: op1_11_inv13 = 1;
    70: op1_11_inv13 = 1;
    76: op1_11_inv13 = 1;
    77: op1_11_inv13 = 1;
    80: op1_11_inv13 = 1;
    81: op1_11_inv13 = 1;
    82: op1_11_inv13 = 1;
    83: op1_11_inv13 = 1;
    84: op1_11_inv13 = 1;
    85: op1_11_inv13 = 1;
    91: op1_11_inv13 = 1;
    92: op1_11_inv13 = 1;
    93: op1_11_inv13 = 1;
    default: op1_11_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in14 = reg_0587;
    5: op1_11_in14 = reg_0654;
    6: op1_11_in14 = imem05_in[111:108];
    8: op1_11_in14 = imem03_in[39:36];
    9: op1_11_in14 = reg_0189;
    10: op1_11_in14 = reg_0278;
    11: op1_11_in14 = reg_0459;
    12: op1_11_in14 = reg_0259;
    82: op1_11_in14 = reg_0259;
    13: op1_11_in14 = reg_0429;
    14: op1_11_in14 = reg_0480;
    32: op1_11_in14 = reg_0480;
    15: op1_11_in14 = imem04_in[23:20];
    68: op1_11_in14 = imem04_in[23:20];
    16: op1_11_in14 = reg_0613;
    17: op1_11_in14 = reg_0043;
    76: op1_11_in14 = reg_0043;
    18: op1_11_in14 = reg_0135;
    19: op1_11_in14 = imem04_in[43:40];
    20: op1_11_in14 = reg_0730;
    21: op1_11_in14 = reg_0110;
    22: op1_11_in14 = reg_0598;
    23: op1_11_in14 = imem02_in[123:120];
    24: op1_11_in14 = imem04_in[83:80];
    25: op1_11_in14 = reg_0197;
    26: op1_11_in14 = reg_0276;
    90: op1_11_in14 = reg_0276;
    27: op1_11_in14 = reg_0782;
    28: op1_11_in14 = reg_0343;
    29: op1_11_in14 = reg_0575;
    30: op1_11_in14 = reg_0369;
    31: op1_11_in14 = reg_0473;
    33: op1_11_in14 = imem04_in[127:124];
    36: op1_11_in14 = reg_0557;
    38: op1_11_in14 = reg_0757;
    39: op1_11_in14 = imem04_in[31:28];
    40: op1_11_in14 = reg_0059;
    42: op1_11_in14 = imem01_in[95:92];
    43: op1_11_in14 = reg_0322;
    46: op1_11_in14 = reg_0322;
    44: op1_11_in14 = reg_0409;
    47: op1_11_in14 = reg_0218;
    66: op1_11_in14 = reg_0218;
    48: op1_11_in14 = reg_0064;
    49: op1_11_in14 = reg_0491;
    50: op1_11_in14 = reg_0529;
    51: op1_11_in14 = imem02_in[11:8];
    52: op1_11_in14 = reg_0551;
    53: op1_11_in14 = imem04_in[3:0];
    54: op1_11_in14 = reg_0632;
    56: op1_11_in14 = imem07_in[83:80];
    57: op1_11_in14 = reg_0721;
    60: op1_11_in14 = reg_0209;
    61: op1_11_in14 = reg_0586;
    62: op1_11_in14 = reg_0151;
    63: op1_11_in14 = reg_0151;
    64: op1_11_in14 = reg_0787;
    65: op1_11_in14 = reg_0159;
    67: op1_11_in14 = reg_0621;
    70: op1_11_in14 = imem01_in[19:16];
    71: op1_11_in14 = reg_0153;
    74: op1_11_in14 = reg_0210;
    75: op1_11_in14 = reg_0594;
    77: op1_11_in14 = reg_0616;
    78: op1_11_in14 = reg_0828;
    80: op1_11_in14 = reg_0475;
    81: op1_11_in14 = reg_0727;
    83: op1_11_in14 = imem02_in[55:52];
    84: op1_11_in14 = reg_0724;
    85: op1_11_in14 = reg_0469;
    86: op1_11_in14 = reg_0610;
    87: op1_11_in14 = reg_0710;
    88: op1_11_in14 = reg_0316;
    89: op1_11_in14 = reg_0351;
    91: op1_11_in14 = reg_0199;
    92: op1_11_in14 = reg_0080;
    93: op1_11_in14 = reg_0320;
    94: op1_11_in14 = reg_0487;
    95: op1_11_in14 = reg_0590;
    default: op1_11_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv14 = 1;
    6: op1_11_inv14 = 1;
    8: op1_11_inv14 = 1;
    9: op1_11_inv14 = 1;
    11: op1_11_inv14 = 1;
    12: op1_11_inv14 = 1;
    13: op1_11_inv14 = 1;
    14: op1_11_inv14 = 1;
    16: op1_11_inv14 = 1;
    17: op1_11_inv14 = 1;
    19: op1_11_inv14 = 1;
    21: op1_11_inv14 = 1;
    23: op1_11_inv14 = 1;
    24: op1_11_inv14 = 1;
    26: op1_11_inv14 = 1;
    30: op1_11_inv14 = 1;
    33: op1_11_inv14 = 1;
    38: op1_11_inv14 = 1;
    40: op1_11_inv14 = 1;
    42: op1_11_inv14 = 1;
    47: op1_11_inv14 = 1;
    50: op1_11_inv14 = 1;
    52: op1_11_inv14 = 1;
    57: op1_11_inv14 = 1;
    60: op1_11_inv14 = 1;
    61: op1_11_inv14 = 1;
    64: op1_11_inv14 = 1;
    67: op1_11_inv14 = 1;
    68: op1_11_inv14 = 1;
    70: op1_11_inv14 = 1;
    76: op1_11_inv14 = 1;
    78: op1_11_inv14 = 1;
    80: op1_11_inv14 = 1;
    81: op1_11_inv14 = 1;
    82: op1_11_inv14 = 1;
    83: op1_11_inv14 = 1;
    87: op1_11_inv14 = 1;
    88: op1_11_inv14 = 1;
    90: op1_11_inv14 = 1;
    91: op1_11_inv14 = 1;
    92: op1_11_inv14 = 1;
    93: op1_11_inv14 = 1;
    default: op1_11_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in15 = reg_0588;
    5: op1_11_in15 = reg_0656;
    6: op1_11_in15 = imem05_in[115:112];
    8: op1_11_in15 = imem03_in[43:40];
    9: op1_11_in15 = reg_0186;
    10: op1_11_in15 = reg_0046;
    11: op1_11_in15 = reg_0452;
    12: op1_11_in15 = reg_0273;
    13: op1_11_in15 = reg_0432;
    14: op1_11_in15 = reg_0473;
    15: op1_11_in15 = imem04_in[27:24];
    16: op1_11_in15 = reg_0617;
    17: op1_11_in15 = reg_0055;
    18: op1_11_in15 = reg_0156;
    19: op1_11_in15 = imem04_in[67:64];
    20: op1_11_in15 = reg_0731;
    21: op1_11_in15 = imem02_in[11:8];
    22: op1_11_in15 = reg_0582;
    23: op1_11_in15 = reg_0650;
    24: op1_11_in15 = imem04_in[91:88];
    25: op1_11_in15 = imem01_in[19:16];
    26: op1_11_in15 = reg_0260;
    27: op1_11_in15 = reg_0783;
    28: op1_11_in15 = reg_0097;
    29: op1_11_in15 = reg_0568;
    30: op1_11_in15 = reg_0408;
    31: op1_11_in15 = reg_0467;
    32: op1_11_in15 = reg_0468;
    33: op1_11_in15 = reg_0542;
    36: op1_11_in15 = reg_0760;
    38: op1_11_in15 = imem03_in[39:36];
    39: op1_11_in15 = imem04_in[51:48];
    40: op1_11_in15 = reg_0056;
    42: op1_11_in15 = imem01_in[111:108];
    43: op1_11_in15 = reg_0343;
    44: op1_11_in15 = reg_0329;
    46: op1_11_in15 = reg_0518;
    47: op1_11_in15 = reg_0020;
    48: op1_11_in15 = reg_0439;
    49: op1_11_in15 = reg_0793;
    50: op1_11_in15 = reg_0430;
    51: op1_11_in15 = imem02_in[15:12];
    52: op1_11_in15 = reg_0556;
    53: op1_11_in15 = imem04_in[7:4];
    54: op1_11_in15 = reg_0623;
    56: op1_11_in15 = reg_0720;
    57: op1_11_in15 = reg_0717;
    60: op1_11_in15 = reg_0194;
    61: op1_11_in15 = reg_0324;
    62: op1_11_in15 = reg_0128;
    63: op1_11_in15 = reg_0142;
    64: op1_11_in15 = reg_0752;
    65: op1_11_in15 = reg_0169;
    66: op1_11_in15 = reg_0794;
    67: op1_11_in15 = reg_0657;
    89: op1_11_in15 = reg_0657;
    68: op1_11_in15 = imem04_in[75:72];
    70: op1_11_in15 = imem01_in[47:44];
    71: op1_11_in15 = reg_0144;
    74: op1_11_in15 = reg_0189;
    75: op1_11_in15 = reg_0342;
    76: op1_11_in15 = reg_0088;
    77: op1_11_in15 = reg_0614;
    86: op1_11_in15 = reg_0614;
    78: op1_11_in15 = imem06_in[7:4];
    80: op1_11_in15 = reg_0462;
    81: op1_11_in15 = reg_0334;
    82: op1_11_in15 = reg_0296;
    83: op1_11_in15 = imem02_in[67:64];
    84: op1_11_in15 = reg_0103;
    85: op1_11_in15 = reg_0476;
    87: op1_11_in15 = reg_0161;
    88: op1_11_in15 = reg_0544;
    90: op1_11_in15 = reg_0748;
    91: op1_11_in15 = reg_0192;
    92: op1_11_in15 = reg_0341;
    93: op1_11_in15 = reg_0361;
    94: op1_11_in15 = reg_0136;
    95: op1_11_in15 = reg_0514;
    default: op1_11_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv15 = 1;
    8: op1_11_inv15 = 1;
    10: op1_11_inv15 = 1;
    11: op1_11_inv15 = 1;
    14: op1_11_inv15 = 1;
    15: op1_11_inv15 = 1;
    16: op1_11_inv15 = 1;
    18: op1_11_inv15 = 1;
    23: op1_11_inv15 = 1;
    24: op1_11_inv15 = 1;
    27: op1_11_inv15 = 1;
    30: op1_11_inv15 = 1;
    32: op1_11_inv15 = 1;
    36: op1_11_inv15 = 1;
    38: op1_11_inv15 = 1;
    43: op1_11_inv15 = 1;
    44: op1_11_inv15 = 1;
    46: op1_11_inv15 = 1;
    47: op1_11_inv15 = 1;
    48: op1_11_inv15 = 1;
    49: op1_11_inv15 = 1;
    50: op1_11_inv15 = 1;
    54: op1_11_inv15 = 1;
    57: op1_11_inv15 = 1;
    61: op1_11_inv15 = 1;
    67: op1_11_inv15 = 1;
    70: op1_11_inv15 = 1;
    74: op1_11_inv15 = 1;
    77: op1_11_inv15 = 1;
    82: op1_11_inv15 = 1;
    84: op1_11_inv15 = 1;
    85: op1_11_inv15 = 1;
    86: op1_11_inv15 = 1;
    88: op1_11_inv15 = 1;
    89: op1_11_inv15 = 1;
    92: op1_11_inv15 = 1;
    93: op1_11_inv15 = 1;
    94: op1_11_inv15 = 1;
    95: op1_11_inv15 = 1;
    default: op1_11_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in16 = reg_0311;
    5: op1_11_in16 = reg_0640;
    6: op1_11_in16 = reg_0792;
    8: op1_11_in16 = imem03_in[83:80];
    9: op1_11_in16 = reg_0739;
    10: op1_11_in16 = reg_0047;
    11: op1_11_in16 = reg_0189;
    12: op1_11_in16 = reg_0527;
    13: op1_11_in16 = reg_0433;
    14: op1_11_in16 = reg_0474;
    15: op1_11_in16 = imem04_in[51:48];
    16: op1_11_in16 = reg_0616;
    17: op1_11_in16 = reg_0553;
    18: op1_11_in16 = reg_0131;
    19: op1_11_in16 = imem04_in[99:96];
    20: op1_11_in16 = reg_0721;
    21: op1_11_in16 = imem02_in[31:28];
    22: op1_11_in16 = reg_0596;
    23: op1_11_in16 = reg_0645;
    24: op1_11_in16 = reg_0545;
    25: op1_11_in16 = imem01_in[47:44];
    26: op1_11_in16 = reg_0732;
    27: op1_11_in16 = reg_0786;
    28: op1_11_in16 = reg_0757;
    29: op1_11_in16 = reg_0569;
    30: op1_11_in16 = reg_0407;
    31: op1_11_in16 = reg_0479;
    32: op1_11_in16 = reg_0458;
    33: op1_11_in16 = reg_0083;
    36: op1_11_in16 = reg_0217;
    38: op1_11_in16 = imem03_in[47:44];
    39: op1_11_in16 = imem04_in[71:68];
    40: op1_11_in16 = reg_0555;
    42: op1_11_in16 = reg_0497;
    43: op1_11_in16 = reg_0096;
    44: op1_11_in16 = reg_0406;
    46: op1_11_in16 = reg_0081;
    47: op1_11_in16 = reg_0339;
    48: op1_11_in16 = reg_0181;
    49: op1_11_in16 = imem05_in[67:64];
    50: op1_11_in16 = reg_0077;
    51: op1_11_in16 = imem02_in[43:40];
    52: op1_11_in16 = reg_0547;
    53: op1_11_in16 = imem04_in[15:12];
    54: op1_11_in16 = imem07_in[7:4];
    56: op1_11_in16 = reg_0700;
    57: op1_11_in16 = reg_0709;
    60: op1_11_in16 = reg_0202;
    61: op1_11_in16 = reg_0097;
    62: op1_11_in16 = reg_0141;
    63: op1_11_in16 = reg_0153;
    64: op1_11_in16 = reg_0495;
    65: op1_11_in16 = reg_0182;
    66: op1_11_in16 = reg_0656;
    67: op1_11_in16 = reg_0639;
    68: op1_11_in16 = imem04_in[87:84];
    70: op1_11_in16 = imem01_in[51:48];
    71: op1_11_in16 = imem06_in[15:12];
    74: op1_11_in16 = reg_0204;
    75: op1_11_in16 = reg_0566;
    76: op1_11_in16 = reg_0055;
    77: op1_11_in16 = reg_0622;
    78: op1_11_in16 = imem06_in[51:48];
    80: op1_11_in16 = reg_0472;
    81: op1_11_in16 = reg_0253;
    82: op1_11_in16 = reg_0776;
    83: op1_11_in16 = imem02_in[87:84];
    84: op1_11_in16 = reg_0447;
    85: op1_11_in16 = reg_0475;
    86: op1_11_in16 = reg_0078;
    87: op1_11_in16 = reg_0789;
    88: op1_11_in16 = reg_0173;
    89: op1_11_in16 = reg_0609;
    90: op1_11_in16 = reg_0169;
    91: op1_11_in16 = imem01_in[59:56];
    92: op1_11_in16 = reg_0359;
    93: op1_11_in16 = reg_0356;
    94: op1_11_in16 = reg_0117;
    95: op1_11_in16 = reg_0092;
    default: op1_11_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv16 = 1;
    6: op1_11_inv16 = 1;
    11: op1_11_inv16 = 1;
    16: op1_11_inv16 = 1;
    17: op1_11_inv16 = 1;
    18: op1_11_inv16 = 1;
    19: op1_11_inv16 = 1;
    23: op1_11_inv16 = 1;
    25: op1_11_inv16 = 1;
    27: op1_11_inv16 = 1;
    30: op1_11_inv16 = 1;
    31: op1_11_inv16 = 1;
    32: op1_11_inv16 = 1;
    44: op1_11_inv16 = 1;
    46: op1_11_inv16 = 1;
    47: op1_11_inv16 = 1;
    48: op1_11_inv16 = 1;
    49: op1_11_inv16 = 1;
    50: op1_11_inv16 = 1;
    51: op1_11_inv16 = 1;
    53: op1_11_inv16 = 1;
    60: op1_11_inv16 = 1;
    62: op1_11_inv16 = 1;
    64: op1_11_inv16 = 1;
    67: op1_11_inv16 = 1;
    68: op1_11_inv16 = 1;
    74: op1_11_inv16 = 1;
    76: op1_11_inv16 = 1;
    77: op1_11_inv16 = 1;
    78: op1_11_inv16 = 1;
    84: op1_11_inv16 = 1;
    85: op1_11_inv16 = 1;
    88: op1_11_inv16 = 1;
    89: op1_11_inv16 = 1;
    91: op1_11_inv16 = 1;
    93: op1_11_inv16 = 1;
    94: op1_11_inv16 = 1;
    default: op1_11_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in17 = reg_0317;
    5: op1_11_in17 = reg_0648;
    6: op1_11_in17 = reg_0796;
    8: op1_11_in17 = reg_0583;
    9: op1_11_in17 = reg_0500;
    10: op1_11_in17 = imem05_in[35:32];
    11: op1_11_in17 = reg_0203;
    12: op1_11_in17 = reg_0526;
    13: op1_11_in17 = reg_0440;
    14: op1_11_in17 = reg_0478;
    15: op1_11_in17 = imem04_in[63:60];
    16: op1_11_in17 = reg_0611;
    17: op1_11_in17 = reg_0542;
    18: op1_11_in17 = reg_0134;
    62: op1_11_in17 = reg_0134;
    19: op1_11_in17 = imem04_in[111:108];
    20: op1_11_in17 = reg_0723;
    21: op1_11_in17 = imem02_in[79:76];
    22: op1_11_in17 = reg_0591;
    23: op1_11_in17 = reg_0666;
    24: op1_11_in17 = reg_0315;
    25: op1_11_in17 = imem01_in[63:60];
    91: op1_11_in17 = imem01_in[63:60];
    26: op1_11_in17 = reg_0734;
    27: op1_11_in17 = reg_0784;
    28: op1_11_in17 = imem03_in[3:0];
    29: op1_11_in17 = reg_0499;
    30: op1_11_in17 = reg_0748;
    31: op1_11_in17 = reg_0452;
    32: op1_11_in17 = reg_0191;
    33: op1_11_in17 = reg_0555;
    36: op1_11_in17 = reg_0503;
    38: op1_11_in17 = imem03_in[67:64];
    39: op1_11_in17 = imem04_in[91:88];
    68: op1_11_in17 = imem04_in[91:88];
    40: op1_11_in17 = reg_0547;
    42: op1_11_in17 = reg_0820;
    43: op1_11_in17 = reg_0540;
    61: op1_11_in17 = reg_0540;
    44: op1_11_in17 = reg_0038;
    46: op1_11_in17 = imem03_in[11:8];
    47: op1_11_in17 = reg_0331;
    48: op1_11_in17 = reg_0179;
    49: op1_11_in17 = imem05_in[87:84];
    50: op1_11_in17 = reg_0071;
    51: op1_11_in17 = reg_0770;
    52: op1_11_in17 = reg_0303;
    53: op1_11_in17 = imem04_in[51:48];
    54: op1_11_in17 = imem07_in[15:12];
    56: op1_11_in17 = reg_0053;
    57: op1_11_in17 = reg_0705;
    60: op1_11_in17 = imem01_in[7:4];
    63: op1_11_in17 = imem06_in[11:8];
    64: op1_11_in17 = imem07_in[51:48];
    65: op1_11_in17 = reg_0170;
    66: op1_11_in17 = reg_0368;
    67: op1_11_in17 = reg_0587;
    70: op1_11_in17 = reg_0336;
    71: op1_11_in17 = imem06_in[59:56];
    78: op1_11_in17 = imem06_in[59:56];
    74: op1_11_in17 = reg_0211;
    75: op1_11_in17 = reg_0514;
    76: op1_11_in17 = reg_0516;
    77: op1_11_in17 = imem05_in[23:20];
    80: op1_11_in17 = reg_0459;
    81: op1_11_in17 = reg_0447;
    82: op1_11_in17 = reg_0644;
    83: op1_11_in17 = imem02_in[103:100];
    84: op1_11_in17 = reg_0448;
    85: op1_11_in17 = reg_0480;
    86: op1_11_in17 = reg_0065;
    87: op1_11_in17 = reg_0158;
    88: op1_11_in17 = reg_0261;
    89: op1_11_in17 = reg_0633;
    90: op1_11_in17 = reg_0650;
    92: op1_11_in17 = reg_0565;
    93: op1_11_in17 = reg_0360;
    94: op1_11_in17 = reg_0255;
    95: op1_11_in17 = reg_0757;
    default: op1_11_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv17 = 1;
    6: op1_11_inv17 = 1;
    8: op1_11_inv17 = 1;
    9: op1_11_inv17 = 1;
    10: op1_11_inv17 = 1;
    12: op1_11_inv17 = 1;
    14: op1_11_inv17 = 1;
    15: op1_11_inv17 = 1;
    16: op1_11_inv17 = 1;
    17: op1_11_inv17 = 1;
    20: op1_11_inv17 = 1;
    21: op1_11_inv17 = 1;
    22: op1_11_inv17 = 1;
    23: op1_11_inv17 = 1;
    24: op1_11_inv17 = 1;
    26: op1_11_inv17 = 1;
    28: op1_11_inv17 = 1;
    33: op1_11_inv17 = 1;
    36: op1_11_inv17 = 1;
    39: op1_11_inv17 = 1;
    43: op1_11_inv17 = 1;
    44: op1_11_inv17 = 1;
    46: op1_11_inv17 = 1;
    49: op1_11_inv17 = 1;
    54: op1_11_inv17 = 1;
    60: op1_11_inv17 = 1;
    61: op1_11_inv17 = 1;
    63: op1_11_inv17 = 1;
    65: op1_11_inv17 = 1;
    66: op1_11_inv17 = 1;
    68: op1_11_inv17 = 1;
    74: op1_11_inv17 = 1;
    75: op1_11_inv17 = 1;
    76: op1_11_inv17 = 1;
    77: op1_11_inv17 = 1;
    80: op1_11_inv17 = 1;
    83: op1_11_inv17 = 1;
    86: op1_11_inv17 = 1;
    87: op1_11_inv17 = 1;
    88: op1_11_inv17 = 1;
    90: op1_11_inv17 = 1;
    91: op1_11_inv17 = 1;
    93: op1_11_inv17 = 1;
    94: op1_11_inv17 = 1;
    default: op1_11_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in18 = reg_0012;
    5: op1_11_in18 = reg_0662;
    6: op1_11_in18 = reg_0797;
    8: op1_11_in18 = reg_0587;
    9: op1_11_in18 = reg_0227;
    10: op1_11_in18 = imem05_in[39:36];
    11: op1_11_in18 = reg_0193;
    12: op1_11_in18 = reg_0733;
    13: op1_11_in18 = reg_0442;
    14: op1_11_in18 = reg_0214;
    15: op1_11_in18 = imem04_in[95:92];
    16: op1_11_in18 = reg_0577;
    17: op1_11_in18 = reg_0540;
    18: op1_11_in18 = imem06_in[7:4];
    19: op1_11_in18 = imem04_in[123:120];
    20: op1_11_in18 = reg_0702;
    21: op1_11_in18 = imem02_in[115:112];
    22: op1_11_in18 = reg_0563;
    23: op1_11_in18 = reg_0654;
    24: op1_11_in18 = reg_0542;
    25: op1_11_in18 = imem01_in[67:64];
    26: op1_11_in18 = reg_0285;
    27: op1_11_in18 = reg_0489;
    28: op1_11_in18 = imem03_in[35:32];
    29: op1_11_in18 = reg_0396;
    30: op1_11_in18 = imem07_in[7:4];
    31: op1_11_in18 = reg_0188;
    32: op1_11_in18 = reg_0188;
    33: op1_11_in18 = reg_0516;
    36: op1_11_in18 = reg_0041;
    38: op1_11_in18 = imem03_in[83:80];
    39: op1_11_in18 = imem04_in[107:104];
    40: op1_11_in18 = reg_0303;
    42: op1_11_in18 = reg_0771;
    43: op1_11_in18 = reg_0526;
    44: op1_11_in18 = reg_0777;
    46: op1_11_in18 = imem03_in[91:88];
    47: op1_11_in18 = reg_0821;
    48: op1_11_in18 = reg_0169;
    49: op1_11_in18 = imem05_in[91:88];
    50: op1_11_in18 = reg_0431;
    51: op1_11_in18 = reg_0082;
    52: op1_11_in18 = reg_0077;
    53: op1_11_in18 = imem04_in[59:56];
    54: op1_11_in18 = imem07_in[47:44];
    56: op1_11_in18 = reg_0635;
    57: op1_11_in18 = reg_0707;
    60: op1_11_in18 = imem01_in[75:72];
    61: op1_11_in18 = reg_0757;
    62: op1_11_in18 = imem06_in[43:40];
    63: op1_11_in18 = imem06_in[35:32];
    64: op1_11_in18 = imem07_in[63:60];
    66: op1_11_in18 = reg_0021;
    67: op1_11_in18 = reg_0358;
    68: op1_11_in18 = reg_0059;
    70: op1_11_in18 = reg_0111;
    71: op1_11_in18 = imem06_in[67:64];
    74: op1_11_in18 = reg_0186;
    75: op1_11_in18 = reg_0080;
    76: op1_11_in18 = reg_0631;
    77: op1_11_in18 = imem05_in[55:52];
    78: op1_11_in18 = imem06_in[87:84];
    80: op1_11_in18 = reg_0478;
    81: op1_11_in18 = imem07_in[19:16];
    82: op1_11_in18 = imem05_in[3:0];
    83: op1_11_in18 = reg_0344;
    84: op1_11_in18 = reg_0142;
    85: op1_11_in18 = reg_0473;
    86: op1_11_in18 = reg_0687;
    87: op1_11_in18 = reg_0334;
    88: op1_11_in18 = reg_0523;
    89: op1_11_in18 = reg_0661;
    90: op1_11_in18 = reg_0224;
    91: op1_11_in18 = imem01_in[91:88];
    92: op1_11_in18 = reg_0356;
    93: op1_11_in18 = reg_0594;
    94: op1_11_in18 = imem03_in[7:4];
    95: op1_11_in18 = imem03_in[47:44];
    default: op1_11_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv18 = 1;
    9: op1_11_inv18 = 1;
    10: op1_11_inv18 = 1;
    12: op1_11_inv18 = 1;
    13: op1_11_inv18 = 1;
    17: op1_11_inv18 = 1;
    20: op1_11_inv18 = 1;
    24: op1_11_inv18 = 1;
    25: op1_11_inv18 = 1;
    27: op1_11_inv18 = 1;
    29: op1_11_inv18 = 1;
    32: op1_11_inv18 = 1;
    33: op1_11_inv18 = 1;
    39: op1_11_inv18 = 1;
    42: op1_11_inv18 = 1;
    46: op1_11_inv18 = 1;
    47: op1_11_inv18 = 1;
    51: op1_11_inv18 = 1;
    52: op1_11_inv18 = 1;
    56: op1_11_inv18 = 1;
    57: op1_11_inv18 = 1;
    60: op1_11_inv18 = 1;
    62: op1_11_inv18 = 1;
    70: op1_11_inv18 = 1;
    71: op1_11_inv18 = 1;
    75: op1_11_inv18 = 1;
    77: op1_11_inv18 = 1;
    80: op1_11_inv18 = 1;
    81: op1_11_inv18 = 1;
    82: op1_11_inv18 = 1;
    84: op1_11_inv18 = 1;
    85: op1_11_inv18 = 1;
    87: op1_11_inv18 = 1;
    88: op1_11_inv18 = 1;
    90: op1_11_inv18 = 1;
    92: op1_11_inv18 = 1;
    default: op1_11_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in19 = reg_0002;
    5: op1_11_in19 = reg_0644;
    6: op1_11_in19 = reg_0783;
    8: op1_11_in19 = reg_0388;
    9: op1_11_in19 = reg_0734;
    10: op1_11_in19 = imem05_in[123:120];
    11: op1_11_in19 = reg_0207;
    12: op1_11_in19 = reg_0152;
    13: op1_11_in19 = reg_0437;
    14: op1_11_in19 = reg_0191;
    15: op1_11_in19 = imem04_in[115:112];
    16: op1_11_in19 = reg_0408;
    17: op1_11_in19 = reg_0558;
    18: op1_11_in19 = imem06_in[47:44];
    19: op1_11_in19 = reg_0553;
    20: op1_11_in19 = reg_0709;
    21: op1_11_in19 = imem02_in[123:120];
    22: op1_11_in19 = reg_0595;
    23: op1_11_in19 = reg_0646;
    24: op1_11_in19 = reg_0043;
    25: op1_11_in19 = reg_0514;
    26: op1_11_in19 = reg_0140;
    27: op1_11_in19 = reg_0309;
    28: op1_11_in19 = imem03_in[63:60];
    29: op1_11_in19 = reg_0013;
    30: op1_11_in19 = imem07_in[43:40];
    31: op1_11_in19 = reg_0211;
    32: op1_11_in19 = imem01_in[23:20];
    33: op1_11_in19 = reg_0273;
    36: op1_11_in19 = reg_0219;
    38: op1_11_in19 = reg_0039;
    39: op1_11_in19 = reg_0059;
    40: op1_11_in19 = reg_0308;
    42: op1_11_in19 = reg_0487;
    43: op1_11_in19 = imem03_in[27:24];
    94: op1_11_in19 = imem03_in[27:24];
    44: op1_11_in19 = reg_0368;
    46: op1_11_in19 = imem03_in[127:124];
    47: op1_11_in19 = reg_0270;
    48: op1_11_in19 = reg_0170;
    49: op1_11_in19 = reg_0150;
    50: op1_11_in19 = reg_0520;
    51: op1_11_in19 = imem03_in[11:8];
    52: op1_11_in19 = reg_0616;
    53: op1_11_in19 = imem04_in[91:88];
    54: op1_11_in19 = imem07_in[83:80];
    56: op1_11_in19 = reg_0440;
    57: op1_11_in19 = reg_0706;
    60: op1_11_in19 = imem01_in[79:76];
    61: op1_11_in19 = imem03_in[59:56];
    62: op1_11_in19 = imem06_in[67:64];
    63: op1_11_in19 = imem06_in[39:36];
    64: op1_11_in19 = imem07_in[67:64];
    66: op1_11_in19 = reg_0029;
    67: op1_11_in19 = reg_0364;
    68: op1_11_in19 = reg_0056;
    70: op1_11_in19 = reg_0394;
    71: op1_11_in19 = imem06_in[71:68];
    74: op1_11_in19 = reg_0196;
    75: op1_11_in19 = reg_0530;
    76: op1_11_in19 = reg_0529;
    77: op1_11_in19 = imem05_in[83:80];
    78: op1_11_in19 = imem06_in[107:104];
    80: op1_11_in19 = reg_0203;
    81: op1_11_in19 = imem07_in[27:24];
    82: op1_11_in19 = imem05_in[59:56];
    83: op1_11_in19 = reg_0587;
    84: op1_11_in19 = reg_0066;
    85: op1_11_in19 = reg_0470;
    86: op1_11_in19 = reg_0622;
    87: op1_11_in19 = reg_0067;
    88: op1_11_in19 = reg_0052;
    89: op1_11_in19 = reg_0224;
    90: op1_11_in19 = imem07_in[19:16];
    91: op1_11_in19 = imem01_in[119:116];
    92: op1_11_in19 = reg_0324;
    93: op1_11_in19 = reg_0414;
    95: op1_11_in19 = imem03_in[75:72];
    default: op1_11_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv19 = 1;
    6: op1_11_inv19 = 1;
    10: op1_11_inv19 = 1;
    11: op1_11_inv19 = 1;
    12: op1_11_inv19 = 1;
    15: op1_11_inv19 = 1;
    16: op1_11_inv19 = 1;
    17: op1_11_inv19 = 1;
    20: op1_11_inv19 = 1;
    22: op1_11_inv19 = 1;
    26: op1_11_inv19 = 1;
    27: op1_11_inv19 = 1;
    33: op1_11_inv19 = 1;
    38: op1_11_inv19 = 1;
    43: op1_11_inv19 = 1;
    44: op1_11_inv19 = 1;
    47: op1_11_inv19 = 1;
    48: op1_11_inv19 = 1;
    49: op1_11_inv19 = 1;
    50: op1_11_inv19 = 1;
    51: op1_11_inv19 = 1;
    52: op1_11_inv19 = 1;
    54: op1_11_inv19 = 1;
    56: op1_11_inv19 = 1;
    57: op1_11_inv19 = 1;
    61: op1_11_inv19 = 1;
    68: op1_11_inv19 = 1;
    70: op1_11_inv19 = 1;
    74: op1_11_inv19 = 1;
    75: op1_11_inv19 = 1;
    76: op1_11_inv19 = 1;
    77: op1_11_inv19 = 1;
    80: op1_11_inv19 = 1;
    81: op1_11_inv19 = 1;
    84: op1_11_inv19 = 1;
    87: op1_11_inv19 = 1;
    88: op1_11_inv19 = 1;
    92: op1_11_inv19 = 1;
    94: op1_11_inv19 = 1;
    95: op1_11_inv19 = 1;
    default: op1_11_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in20 = reg_0013;
    5: op1_11_in20 = reg_0643;
    6: op1_11_in20 = reg_0790;
    8: op1_11_in20 = reg_0327;
    9: op1_11_in20 = reg_0519;
    25: op1_11_in20 = reg_0519;
    10: op1_11_in20 = reg_0798;
    11: op1_11_in20 = reg_0198;
    31: op1_11_in20 = reg_0198;
    12: op1_11_in20 = reg_0142;
    13: op1_11_in20 = reg_0179;
    14: op1_11_in20 = reg_0204;
    15: op1_11_in20 = imem04_in[119:116];
    53: op1_11_in20 = imem04_in[119:116];
    16: op1_11_in20 = reg_0349;
    17: op1_11_in20 = reg_0556;
    68: op1_11_in20 = reg_0556;
    18: op1_11_in20 = imem06_in[63:60];
    19: op1_11_in20 = reg_0546;
    20: op1_11_in20 = reg_0713;
    21: op1_11_in20 = reg_0655;
    22: op1_11_in20 = reg_0384;
    23: op1_11_in20 = reg_0657;
    24: op1_11_in20 = reg_0060;
    26: op1_11_in20 = imem06_in[15:12];
    27: op1_11_in20 = reg_0735;
    28: op1_11_in20 = imem03_in[67:64];
    29: op1_11_in20 = reg_0007;
    30: op1_11_in20 = imem07_in[63:60];
    32: op1_11_in20 = imem01_in[31:28];
    33: op1_11_in20 = reg_0293;
    36: op1_11_in20 = reg_0508;
    38: op1_11_in20 = reg_0751;
    39: op1_11_in20 = reg_0262;
    40: op1_11_in20 = reg_0302;
    42: op1_11_in20 = reg_0760;
    43: op1_11_in20 = imem03_in[71:68];
    44: op1_11_in20 = reg_0367;
    46: op1_11_in20 = reg_0586;
    47: op1_11_in20 = reg_0812;
    48: op1_11_in20 = reg_0158;
    49: op1_11_in20 = reg_0154;
    50: op1_11_in20 = reg_0513;
    51: op1_11_in20 = imem03_in[23:20];
    52: op1_11_in20 = reg_0050;
    54: op1_11_in20 = reg_0719;
    56: op1_11_in20 = reg_0443;
    57: op1_11_in20 = reg_0700;
    60: op1_11_in20 = imem01_in[107:104];
    61: op1_11_in20 = imem03_in[123:120];
    62: op1_11_in20 = imem06_in[123:120];
    63: op1_11_in20 = imem06_in[43:40];
    64: op1_11_in20 = imem07_in[71:68];
    66: op1_11_in20 = imem07_in[23:20];
    67: op1_11_in20 = reg_0345;
    83: op1_11_in20 = reg_0345;
    70: op1_11_in20 = reg_0737;
    71: op1_11_in20 = imem06_in[75:72];
    74: op1_11_in20 = imem01_in[7:4];
    75: op1_11_in20 = reg_0094;
    76: op1_11_in20 = reg_0614;
    77: op1_11_in20 = reg_0145;
    78: op1_11_in20 = imem06_in[111:108];
    80: op1_11_in20 = reg_0212;
    81: op1_11_in20 = imem07_in[79:76];
    82: op1_11_in20 = imem05_in[71:68];
    85: op1_11_in20 = reg_0459;
    86: op1_11_in20 = reg_0311;
    87: op1_11_in20 = reg_0051;
    88: op1_11_in20 = reg_0631;
    89: op1_11_in20 = imem07_in[3:0];
    90: op1_11_in20 = imem07_in[75:72];
    91: op1_11_in20 = reg_0668;
    92: op1_11_in20 = reg_0353;
    93: op1_11_in20 = reg_0514;
    94: op1_11_in20 = imem03_in[63:60];
    95: op1_11_in20 = imem03_in[103:100];
    default: op1_11_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv20 = 1;
    5: op1_11_inv20 = 1;
    8: op1_11_inv20 = 1;
    11: op1_11_inv20 = 1;
    13: op1_11_inv20 = 1;
    14: op1_11_inv20 = 1;
    15: op1_11_inv20 = 1;
    16: op1_11_inv20 = 1;
    17: op1_11_inv20 = 1;
    18: op1_11_inv20 = 1;
    20: op1_11_inv20 = 1;
    21: op1_11_inv20 = 1;
    22: op1_11_inv20 = 1;
    26: op1_11_inv20 = 1;
    27: op1_11_inv20 = 1;
    28: op1_11_inv20 = 1;
    30: op1_11_inv20 = 1;
    31: op1_11_inv20 = 1;
    32: op1_11_inv20 = 1;
    33: op1_11_inv20 = 1;
    36: op1_11_inv20 = 1;
    38: op1_11_inv20 = 1;
    39: op1_11_inv20 = 1;
    43: op1_11_inv20 = 1;
    50: op1_11_inv20 = 1;
    51: op1_11_inv20 = 1;
    52: op1_11_inv20 = 1;
    61: op1_11_inv20 = 1;
    63: op1_11_inv20 = 1;
    66: op1_11_inv20 = 1;
    67: op1_11_inv20 = 1;
    68: op1_11_inv20 = 1;
    76: op1_11_inv20 = 1;
    80: op1_11_inv20 = 1;
    85: op1_11_inv20 = 1;
    86: op1_11_inv20 = 1;
    87: op1_11_inv20 = 1;
    90: op1_11_inv20 = 1;
    91: op1_11_inv20 = 1;
    92: op1_11_inv20 = 1;
    93: op1_11_inv20 = 1;
    default: op1_11_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in21 = reg_0014;
    5: op1_11_in21 = reg_0663;
    6: op1_11_in21 = reg_0250;
    8: op1_11_in21 = reg_0396;
    9: op1_11_in21 = reg_0517;
    10: op1_11_in21 = reg_0492;
    11: op1_11_in21 = reg_0201;
    31: op1_11_in21 = reg_0201;
    12: op1_11_in21 = reg_0146;
    13: op1_11_in21 = reg_0161;
    14: op1_11_in21 = reg_0188;
    15: op1_11_in21 = imem04_in[127:124];
    16: op1_11_in21 = reg_0409;
    17: op1_11_in21 = reg_0308;
    68: op1_11_in21 = reg_0308;
    18: op1_11_in21 = imem06_in[91:88];
    19: op1_11_in21 = reg_0540;
    20: op1_11_in21 = reg_0430;
    21: op1_11_in21 = reg_0654;
    22: op1_11_in21 = reg_0373;
    23: op1_11_in21 = reg_0656;
    24: op1_11_in21 = reg_0516;
    25: op1_11_in21 = reg_0825;
    26: op1_11_in21 = imem06_in[75:72];
    27: op1_11_in21 = reg_0260;
    28: op1_11_in21 = imem03_in[75:72];
    43: op1_11_in21 = imem03_in[75:72];
    29: op1_11_in21 = reg_0008;
    30: op1_11_in21 = imem07_in[107:104];
    32: op1_11_in21 = imem01_in[59:56];
    33: op1_11_in21 = reg_0079;
    36: op1_11_in21 = reg_0105;
    38: op1_11_in21 = reg_0590;
    39: op1_11_in21 = reg_0545;
    40: op1_11_in21 = reg_0050;
    42: op1_11_in21 = reg_0241;
    44: op1_11_in21 = imem07_in[3:0];
    46: op1_11_in21 = reg_0582;
    47: op1_11_in21 = reg_0778;
    49: op1_11_in21 = reg_0143;
    50: op1_11_in21 = reg_0585;
    51: op1_11_in21 = imem03_in[47:44];
    52: op1_11_in21 = reg_0617;
    53: op1_11_in21 = reg_0059;
    54: op1_11_in21 = reg_0714;
    56: op1_11_in21 = reg_0437;
    57: op1_11_in21 = reg_0266;
    60: op1_11_in21 = imem01_in[111:108];
    61: op1_11_in21 = reg_0579;
    62: op1_11_in21 = reg_0291;
    63: op1_11_in21 = imem06_in[71:68];
    64: op1_11_in21 = imem07_in[75:72];
    66: op1_11_in21 = imem07_in[87:84];
    67: op1_11_in21 = reg_0361;
    83: op1_11_in21 = reg_0361;
    70: op1_11_in21 = reg_0507;
    71: op1_11_in21 = imem06_in[79:76];
    74: op1_11_in21 = imem01_in[43:40];
    75: op1_11_in21 = imem03_in[19:16];
    76: op1_11_in21 = reg_0679;
    77: op1_11_in21 = reg_0144;
    78: op1_11_in21 = imem06_in[123:120];
    80: op1_11_in21 = reg_0202;
    81: op1_11_in21 = imem07_in[111:108];
    82: op1_11_in21 = imem05_in[79:76];
    85: op1_11_in21 = reg_0209;
    86: op1_11_in21 = reg_0776;
    87: op1_11_in21 = reg_0439;
    88: op1_11_in21 = reg_0616;
    89: op1_11_in21 = imem07_in[7:4];
    90: op1_11_in21 = imem07_in[103:100];
    91: op1_11_in21 = reg_0520;
    92: op1_11_in21 = reg_0343;
    93: op1_11_in21 = reg_0092;
    94: op1_11_in21 = imem03_in[67:64];
    95: op1_11_in21 = imem03_in[127:124];
    default: op1_11_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv21 = 1;
    13: op1_11_inv21 = 1;
    14: op1_11_inv21 = 1;
    15: op1_11_inv21 = 1;
    17: op1_11_inv21 = 1;
    18: op1_11_inv21 = 1;
    19: op1_11_inv21 = 1;
    20: op1_11_inv21 = 1;
    23: op1_11_inv21 = 1;
    24: op1_11_inv21 = 1;
    26: op1_11_inv21 = 1;
    27: op1_11_inv21 = 1;
    28: op1_11_inv21 = 1;
    32: op1_11_inv21 = 1;
    36: op1_11_inv21 = 1;
    40: op1_11_inv21 = 1;
    42: op1_11_inv21 = 1;
    46: op1_11_inv21 = 1;
    47: op1_11_inv21 = 1;
    51: op1_11_inv21 = 1;
    56: op1_11_inv21 = 1;
    57: op1_11_inv21 = 1;
    60: op1_11_inv21 = 1;
    61: op1_11_inv21 = 1;
    62: op1_11_inv21 = 1;
    64: op1_11_inv21 = 1;
    66: op1_11_inv21 = 1;
    67: op1_11_inv21 = 1;
    68: op1_11_inv21 = 1;
    71: op1_11_inv21 = 1;
    74: op1_11_inv21 = 1;
    77: op1_11_inv21 = 1;
    81: op1_11_inv21 = 1;
    87: op1_11_inv21 = 1;
    88: op1_11_inv21 = 1;
    89: op1_11_inv21 = 1;
    91: op1_11_inv21 = 1;
    92: op1_11_inv21 = 1;
    93: op1_11_inv21 = 1;
    95: op1_11_inv21 = 1;
    default: op1_11_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in22 = reg_0015;
    86: op1_11_in22 = reg_0015;
    5: op1_11_in22 = reg_0359;
    6: op1_11_in22 = reg_0152;
    8: op1_11_in22 = reg_0389;
    9: op1_11_in22 = reg_0515;
    10: op1_11_in22 = reg_0780;
    11: op1_11_in22 = reg_0197;
    80: op1_11_in22 = reg_0197;
    12: op1_11_in22 = reg_0137;
    13: op1_11_in22 = reg_0160;
    14: op1_11_in22 = reg_0212;
    15: op1_11_in22 = reg_0543;
    16: op1_11_in22 = reg_0375;
    17: op1_11_in22 = reg_0301;
    18: op1_11_in22 = imem06_in[99:96];
    19: op1_11_in22 = reg_0558;
    20: op1_11_in22 = reg_0426;
    21: op1_11_in22 = reg_0637;
    22: op1_11_in22 = reg_0396;
    23: op1_11_in22 = reg_0649;
    24: op1_11_in22 = reg_0547;
    25: op1_11_in22 = reg_0759;
    26: op1_11_in22 = imem06_in[107:104];
    27: op1_11_in22 = reg_0269;
    28: op1_11_in22 = imem03_in[99:96];
    43: op1_11_in22 = imem03_in[99:96];
    29: op1_11_in22 = reg_0802;
    30: op1_11_in22 = reg_0721;
    31: op1_11_in22 = reg_0213;
    32: op1_11_in22 = imem01_in[83:80];
    33: op1_11_in22 = reg_0255;
    36: op1_11_in22 = reg_0124;
    38: op1_11_in22 = reg_0007;
    39: op1_11_in22 = reg_0552;
    40: op1_11_in22 = reg_0257;
    42: op1_11_in22 = reg_0418;
    44: op1_11_in22 = imem07_in[103:100];
    46: op1_11_in22 = reg_0599;
    47: op1_11_in22 = imem07_in[47:44];
    49: op1_11_in22 = reg_0153;
    50: op1_11_in22 = reg_0233;
    51: op1_11_in22 = imem03_in[55:52];
    52: op1_11_in22 = reg_0078;
    53: op1_11_in22 = reg_0058;
    54: op1_11_in22 = reg_0729;
    56: op1_11_in22 = reg_0180;
    57: op1_11_in22 = reg_0333;
    60: op1_11_in22 = reg_0820;
    61: op1_11_in22 = reg_0493;
    62: op1_11_in22 = reg_0577;
    63: op1_11_in22 = imem06_in[83:80];
    64: op1_11_in22 = imem07_in[83:80];
    66: op1_11_in22 = imem07_in[111:108];
    67: op1_11_in22 = reg_0356;
    68: op1_11_in22 = reg_0283;
    70: op1_11_in22 = reg_0511;
    71: op1_11_in22 = reg_0348;
    74: op1_11_in22 = reg_0111;
    75: op1_11_in22 = imem03_in[35:32];
    76: op1_11_in22 = reg_0644;
    77: op1_11_in22 = reg_0226;
    78: op1_11_in22 = reg_0624;
    82: op1_11_in22 = imem05_in[95:92];
    83: op1_11_in22 = reg_0324;
    85: op1_11_in22 = reg_0207;
    87: op1_11_in22 = reg_0139;
    88: op1_11_in22 = reg_0292;
    89: op1_11_in22 = imem07_in[23:20];
    90: op1_11_in22 = imem07_in[107:104];
    91: op1_11_in22 = reg_0394;
    92: op1_11_in22 = reg_0514;
    93: op1_11_in22 = reg_0743;
    94: op1_11_in22 = imem03_in[79:76];
    95: op1_11_in22 = reg_0582;
    default: op1_11_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv22 = 1;
    5: op1_11_inv22 = 1;
    9: op1_11_inv22 = 1;
    16: op1_11_inv22 = 1;
    18: op1_11_inv22 = 1;
    19: op1_11_inv22 = 1;
    20: op1_11_inv22 = 1;
    22: op1_11_inv22 = 1;
    23: op1_11_inv22 = 1;
    24: op1_11_inv22 = 1;
    27: op1_11_inv22 = 1;
    28: op1_11_inv22 = 1;
    29: op1_11_inv22 = 1;
    31: op1_11_inv22 = 1;
    32: op1_11_inv22 = 1;
    33: op1_11_inv22 = 1;
    39: op1_11_inv22 = 1;
    40: op1_11_inv22 = 1;
    46: op1_11_inv22 = 1;
    47: op1_11_inv22 = 1;
    49: op1_11_inv22 = 1;
    50: op1_11_inv22 = 1;
    51: op1_11_inv22 = 1;
    52: op1_11_inv22 = 1;
    54: op1_11_inv22 = 1;
    56: op1_11_inv22 = 1;
    60: op1_11_inv22 = 1;
    63: op1_11_inv22 = 1;
    66: op1_11_inv22 = 1;
    68: op1_11_inv22 = 1;
    70: op1_11_inv22 = 1;
    75: op1_11_inv22 = 1;
    77: op1_11_inv22 = 1;
    85: op1_11_inv22 = 1;
    86: op1_11_inv22 = 1;
    89: op1_11_inv22 = 1;
    90: op1_11_inv22 = 1;
    91: op1_11_inv22 = 1;
    92: op1_11_inv22 = 1;
    95: op1_11_inv22 = 1;
    default: op1_11_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in23 = reg_0016;
    5: op1_11_in23 = reg_0083;
    6: op1_11_in23 = reg_0130;
    8: op1_11_in23 = reg_0012;
    9: op1_11_in23 = imem01_in[7:4];
    31: op1_11_in23 = imem01_in[7:4];
    80: op1_11_in23 = imem01_in[7:4];
    10: op1_11_in23 = reg_0495;
    11: op1_11_in23 = imem01_in[27:24];
    12: op1_11_in23 = reg_0134;
    13: op1_11_in23 = reg_0164;
    14: op1_11_in23 = reg_0195;
    15: op1_11_in23 = reg_0529;
    16: op1_11_in23 = reg_0404;
    17: op1_11_in23 = reg_0305;
    18: op1_11_in23 = imem06_in[127:124];
    19: op1_11_in23 = reg_0541;
    20: op1_11_in23 = reg_0423;
    21: op1_11_in23 = reg_0656;
    22: op1_11_in23 = reg_0811;
    23: op1_11_in23 = reg_0641;
    24: op1_11_in23 = reg_0303;
    25: op1_11_in23 = reg_0333;
    26: op1_11_in23 = imem06_in[111:108];
    27: op1_11_in23 = reg_0142;
    28: op1_11_in23 = reg_0602;
    29: op1_11_in23 = reg_0810;
    38: op1_11_in23 = reg_0810;
    30: op1_11_in23 = reg_0718;
    32: op1_11_in23 = reg_0501;
    33: op1_11_in23 = reg_0075;
    77: op1_11_in23 = reg_0075;
    36: op1_11_in23 = reg_0116;
    39: op1_11_in23 = reg_0088;
    40: op1_11_in23 = reg_0068;
    42: op1_11_in23 = reg_0511;
    43: op1_11_in23 = imem03_in[127:124];
    44: op1_11_in23 = imem07_in[111:108];
    46: op1_11_in23 = reg_0579;
    47: op1_11_in23 = imem07_in[51:48];
    49: op1_11_in23 = reg_0140;
    50: op1_11_in23 = reg_0644;
    51: op1_11_in23 = imem03_in[63:60];
    52: op1_11_in23 = reg_0296;
    53: op1_11_in23 = reg_0283;
    54: op1_11_in23 = reg_0713;
    56: op1_11_in23 = reg_0178;
    57: op1_11_in23 = reg_0446;
    60: op1_11_in23 = reg_0765;
    61: op1_11_in23 = reg_0331;
    62: op1_11_in23 = reg_0265;
    63: op1_11_in23 = imem06_in[87:84];
    64: op1_11_in23 = imem07_in[123:120];
    66: op1_11_in23 = reg_0719;
    67: op1_11_in23 = reg_0527;
    68: op1_11_in23 = reg_0076;
    70: op1_11_in23 = reg_0290;
    71: op1_11_in23 = reg_0291;
    74: op1_11_in23 = reg_0102;
    75: op1_11_in23 = imem03_in[59:56];
    76: op1_11_in23 = reg_0416;
    78: op1_11_in23 = reg_0762;
    82: op1_11_in23 = imem05_in[107:104];
    83: op1_11_in23 = reg_0514;
    85: op1_11_in23 = reg_0194;
    86: op1_11_in23 = reg_0486;
    87: op1_11_in23 = reg_0089;
    88: op1_11_in23 = reg_0627;
    89: op1_11_in23 = imem07_in[27:24];
    90: op1_11_in23 = imem07_in[115:112];
    91: op1_11_in23 = reg_0101;
    92: op1_11_in23 = reg_0743;
    93: op1_11_in23 = reg_0136;
    94: op1_11_in23 = imem03_in[95:92];
    95: op1_11_in23 = reg_0383;
    default: op1_11_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv23 = 1;
    5: op1_11_inv23 = 1;
    8: op1_11_inv23 = 1;
    15: op1_11_inv23 = 1;
    16: op1_11_inv23 = 1;
    18: op1_11_inv23 = 1;
    20: op1_11_inv23 = 1;
    21: op1_11_inv23 = 1;
    22: op1_11_inv23 = 1;
    23: op1_11_inv23 = 1;
    24: op1_11_inv23 = 1;
    27: op1_11_inv23 = 1;
    28: op1_11_inv23 = 1;
    30: op1_11_inv23 = 1;
    32: op1_11_inv23 = 1;
    38: op1_11_inv23 = 1;
    39: op1_11_inv23 = 1;
    42: op1_11_inv23 = 1;
    51: op1_11_inv23 = 1;
    52: op1_11_inv23 = 1;
    53: op1_11_inv23 = 1;
    56: op1_11_inv23 = 1;
    60: op1_11_inv23 = 1;
    62: op1_11_inv23 = 1;
    63: op1_11_inv23 = 1;
    64: op1_11_inv23 = 1;
    67: op1_11_inv23 = 1;
    68: op1_11_inv23 = 1;
    70: op1_11_inv23 = 1;
    74: op1_11_inv23 = 1;
    77: op1_11_inv23 = 1;
    80: op1_11_inv23 = 1;
    91: op1_11_inv23 = 1;
    92: op1_11_inv23 = 1;
    95: op1_11_inv23 = 1;
    default: op1_11_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in24 = imem04_in[23:20];
    5: op1_11_in24 = reg_0095;
    92: op1_11_in24 = reg_0095;
    6: op1_11_in24 = imem06_in[27:24];
    8: op1_11_in24 = reg_0803;
    22: op1_11_in24 = reg_0803;
    9: op1_11_in24 = imem01_in[27:24];
    10: op1_11_in24 = reg_0786;
    11: op1_11_in24 = imem01_in[39:36];
    12: op1_11_in24 = imem06_in[3:0];
    14: op1_11_in24 = imem01_in[35:32];
    15: op1_11_in24 = reg_0555;
    16: op1_11_in24 = reg_0406;
    67: op1_11_in24 = reg_0406;
    17: op1_11_in24 = reg_0306;
    18: op1_11_in24 = reg_0624;
    19: op1_11_in24 = reg_0053;
    20: op1_11_in24 = reg_0446;
    21: op1_11_in24 = reg_0636;
    23: op1_11_in24 = reg_0341;
    24: op1_11_in24 = reg_0054;
    42: op1_11_in24 = reg_0054;
    25: op1_11_in24 = reg_0515;
    26: op1_11_in24 = imem06_in[127:124];
    27: op1_11_in24 = reg_0139;
    28: op1_11_in24 = reg_0586;
    29: op1_11_in24 = reg_0009;
    30: op1_11_in24 = reg_0424;
    31: op1_11_in24 = imem01_in[11:8];
    32: op1_11_in24 = reg_0519;
    52: op1_11_in24 = reg_0519;
    33: op1_11_in24 = reg_0256;
    36: op1_11_in24 = reg_0104;
    38: op1_11_in24 = imem04_in[11:8];
    39: op1_11_in24 = reg_0060;
    40: op1_11_in24 = reg_0077;
    43: op1_11_in24 = reg_0259;
    44: op1_11_in24 = reg_0716;
    46: op1_11_in24 = reg_0589;
    47: op1_11_in24 = imem07_in[127:124];
    49: op1_11_in24 = reg_0137;
    50: op1_11_in24 = imem05_in[51:48];
    51: op1_11_in24 = imem03_in[87:84];
    53: op1_11_in24 = reg_0631;
    54: op1_11_in24 = reg_0718;
    57: op1_11_in24 = reg_0175;
    60: op1_11_in24 = reg_0322;
    61: op1_11_in24 = reg_0575;
    62: op1_11_in24 = reg_0260;
    63: op1_11_in24 = imem06_in[99:96];
    64: op1_11_in24 = reg_0719;
    66: op1_11_in24 = reg_0726;
    68: op1_11_in24 = reg_0297;
    70: op1_11_in24 = reg_0248;
    71: op1_11_in24 = reg_0605;
    74: op1_11_in24 = reg_0759;
    75: op1_11_in24 = imem03_in[115:112];
    76: op1_11_in24 = imem05_in[71:68];
    77: op1_11_in24 = reg_0789;
    78: op1_11_in24 = reg_0354;
    80: op1_11_in24 = reg_0111;
    82: op1_11_in24 = imem05_in[119:116];
    83: op1_11_in24 = reg_0743;
    85: op1_11_in24 = reg_0198;
    86: op1_11_in24 = reg_0735;
    87: op1_11_in24 = reg_0181;
    88: op1_11_in24 = reg_0062;
    89: op1_11_in24 = imem07_in[35:32];
    90: op1_11_in24 = reg_0722;
    91: op1_11_in24 = reg_0778;
    93: op1_11_in24 = reg_0703;
    94: op1_11_in24 = imem03_in[119:116];
    95: op1_11_in24 = reg_0801;
    default: op1_11_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv24 = 1;
    8: op1_11_inv24 = 1;
    9: op1_11_inv24 = 1;
    11: op1_11_inv24 = 1;
    14: op1_11_inv24 = 1;
    15: op1_11_inv24 = 1;
    16: op1_11_inv24 = 1;
    17: op1_11_inv24 = 1;
    22: op1_11_inv24 = 1;
    25: op1_11_inv24 = 1;
    27: op1_11_inv24 = 1;
    30: op1_11_inv24 = 1;
    33: op1_11_inv24 = 1;
    36: op1_11_inv24 = 1;
    40: op1_11_inv24 = 1;
    42: op1_11_inv24 = 1;
    43: op1_11_inv24 = 1;
    44: op1_11_inv24 = 1;
    46: op1_11_inv24 = 1;
    49: op1_11_inv24 = 1;
    51: op1_11_inv24 = 1;
    52: op1_11_inv24 = 1;
    53: op1_11_inv24 = 1;
    61: op1_11_inv24 = 1;
    64: op1_11_inv24 = 1;
    68: op1_11_inv24 = 1;
    74: op1_11_inv24 = 1;
    77: op1_11_inv24 = 1;
    80: op1_11_inv24 = 1;
    82: op1_11_inv24 = 1;
    83: op1_11_inv24 = 1;
    85: op1_11_inv24 = 1;
    86: op1_11_inv24 = 1;
    92: op1_11_inv24 = 1;
    94: op1_11_inv24 = 1;
    default: op1_11_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in25 = reg_0543;
    5: op1_11_in25 = reg_0090;
    6: op1_11_in25 = imem06_in[39:36];
    8: op1_11_in25 = reg_0013;
    9: op1_11_in25 = imem01_in[35:32];
    10: op1_11_in25 = reg_0268;
    11: op1_11_in25 = imem01_in[47:44];
    12: op1_11_in25 = imem06_in[43:40];
    14: op1_11_in25 = imem01_in[43:40];
    15: op1_11_in25 = reg_0551;
    16: op1_11_in25 = reg_0367;
    17: op1_11_in25 = reg_0302;
    18: op1_11_in25 = reg_0613;
    19: op1_11_in25 = reg_0305;
    24: op1_11_in25 = reg_0305;
    20: op1_11_in25 = reg_0438;
    21: op1_11_in25 = reg_0352;
    22: op1_11_in25 = reg_0806;
    23: op1_11_in25 = reg_0329;
    25: op1_11_in25 = reg_0232;
    26: op1_11_in25 = reg_0610;
    27: op1_11_in25 = reg_0129;
    28: op1_11_in25 = reg_0579;
    29: op1_11_in25 = reg_0004;
    30: op1_11_in25 = reg_0421;
    31: op1_11_in25 = imem01_in[51:48];
    32: op1_11_in25 = reg_0218;
    33: op1_11_in25 = imem05_in[23:20];
    52: op1_11_in25 = imem05_in[23:20];
    36: op1_11_in25 = reg_0119;
    38: op1_11_in25 = imem04_in[19:16];
    39: op1_11_in25 = reg_0057;
    40: op1_11_in25 = reg_0071;
    42: op1_11_in25 = reg_0219;
    43: op1_11_in25 = reg_0591;
    44: op1_11_in25 = reg_0719;
    46: op1_11_in25 = reg_0600;
    47: op1_11_in25 = reg_0723;
    49: op1_11_in25 = reg_0131;
    50: op1_11_in25 = imem05_in[103:100];
    51: op1_11_in25 = imem03_in[119:116];
    53: op1_11_in25 = reg_0078;
    54: op1_11_in25 = reg_0701;
    57: op1_11_in25 = reg_0161;
    60: op1_11_in25 = reg_0652;
    61: op1_11_in25 = reg_0561;
    62: op1_11_in25 = reg_0405;
    63: op1_11_in25 = imem06_in[127:124];
    64: op1_11_in25 = reg_0730;
    66: op1_11_in25 = reg_0717;
    67: op1_11_in25 = reg_0314;
    68: op1_11_in25 = reg_0050;
    70: op1_11_in25 = reg_0243;
    71: op1_11_in25 = reg_0609;
    74: op1_11_in25 = reg_0737;
    75: op1_11_in25 = imem03_in[123:120];
    94: op1_11_in25 = imem03_in[123:120];
    76: op1_11_in25 = reg_0736;
    77: op1_11_in25 = reg_0491;
    78: op1_11_in25 = reg_0293;
    80: op1_11_in25 = reg_0385;
    82: op1_11_in25 = imem05_in[127:124];
    83: op1_11_in25 = reg_0769;
    85: op1_11_in25 = reg_0196;
    86: op1_11_in25 = reg_0165;
    87: op1_11_in25 = reg_0091;
    88: op1_11_in25 = reg_0598;
    89: op1_11_in25 = imem07_in[43:40];
    90: op1_11_in25 = reg_0716;
    91: op1_11_in25 = reg_0511;
    92: op1_11_in25 = reg_0756;
    93: op1_11_in25 = imem03_in[43:40];
    95: op1_11_in25 = reg_0528;
    default: op1_11_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_11_inv25 = 1;
    8: op1_11_inv25 = 1;
    10: op1_11_inv25 = 1;
    11: op1_11_inv25 = 1;
    15: op1_11_inv25 = 1;
    16: op1_11_inv25 = 1;
    17: op1_11_inv25 = 1;
    19: op1_11_inv25 = 1;
    21: op1_11_inv25 = 1;
    22: op1_11_inv25 = 1;
    23: op1_11_inv25 = 1;
    28: op1_11_inv25 = 1;
    29: op1_11_inv25 = 1;
    30: op1_11_inv25 = 1;
    31: op1_11_inv25 = 1;
    36: op1_11_inv25 = 1;
    38: op1_11_inv25 = 1;
    39: op1_11_inv25 = 1;
    40: op1_11_inv25 = 1;
    50: op1_11_inv25 = 1;
    51: op1_11_inv25 = 1;
    53: op1_11_inv25 = 1;
    57: op1_11_inv25 = 1;
    64: op1_11_inv25 = 1;
    83: op1_11_inv25 = 1;
    86: op1_11_inv25 = 1;
    87: op1_11_inv25 = 1;
    88: op1_11_inv25 = 1;
    90: op1_11_inv25 = 1;
    92: op1_11_inv25 = 1;
    93: op1_11_inv25 = 1;
    default: op1_11_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in26 = reg_0545;
    5: op1_11_in26 = reg_0051;
    6: op1_11_in26 = imem06_in[55:52];
    8: op1_11_in26 = reg_0010;
    9: op1_11_in26 = imem01_in[87:84];
    10: op1_11_in26 = reg_0271;
    11: op1_11_in26 = imem01_in[67:64];
    12: op1_11_in26 = imem06_in[51:48];
    14: op1_11_in26 = imem01_in[51:48];
    15: op1_11_in26 = reg_0559;
    16: op1_11_in26 = reg_0401;
    17: op1_11_in26 = reg_0307;
    18: op1_11_in26 = reg_0633;
    19: op1_11_in26 = reg_0273;
    20: op1_11_in26 = reg_0181;
    21: op1_11_in26 = reg_0358;
    22: op1_11_in26 = imem04_in[11:8];
    23: op1_11_in26 = reg_0339;
    24: op1_11_in26 = reg_0274;
    25: op1_11_in26 = reg_0235;
    74: op1_11_in26 = reg_0235;
    26: op1_11_in26 = reg_0620;
    27: op1_11_in26 = reg_0153;
    28: op1_11_in26 = reg_0583;
    62: op1_11_in26 = reg_0583;
    29: op1_11_in26 = imem04_in[51:48];
    30: op1_11_in26 = reg_0447;
    31: op1_11_in26 = imem01_in[59:56];
    32: op1_11_in26 = reg_0506;
    33: op1_11_in26 = reg_0797;
    36: op1_11_in26 = reg_0114;
    38: op1_11_in26 = imem04_in[47:44];
    39: op1_11_in26 = reg_0516;
    40: op1_11_in26 = reg_0074;
    42: op1_11_in26 = reg_0420;
    43: op1_11_in26 = reg_0578;
    44: op1_11_in26 = reg_0730;
    46: op1_11_in26 = reg_0595;
    47: op1_11_in26 = reg_0702;
    49: op1_11_in26 = reg_0134;
    50: op1_11_in26 = reg_0798;
    51: op1_11_in26 = reg_0601;
    52: op1_11_in26 = imem05_in[55:52];
    53: op1_11_in26 = reg_0501;
    54: op1_11_in26 = reg_0700;
    57: op1_11_in26 = reg_0162;
    60: op1_11_in26 = reg_0737;
    61: op1_11_in26 = reg_0517;
    76: op1_11_in26 = reg_0517;
    63: op1_11_in26 = reg_0289;
    64: op1_11_in26 = reg_0726;
    66: op1_11_in26 = reg_0712;
    67: op1_11_in26 = reg_0096;
    68: op1_11_in26 = reg_0679;
    70: op1_11_in26 = reg_0108;
    71: op1_11_in26 = reg_0238;
    75: op1_11_in26 = reg_0338;
    77: op1_11_in26 = reg_0495;
    78: op1_11_in26 = reg_0377;
    80: op1_11_in26 = reg_0759;
    82: op1_11_in26 = reg_0146;
    83: op1_11_in26 = reg_0756;
    85: op1_11_in26 = reg_0212;
    86: op1_11_in26 = reg_0383;
    88: op1_11_in26 = reg_0069;
    89: op1_11_in26 = imem07_in[83:80];
    90: op1_11_in26 = reg_0721;
    91: op1_11_in26 = reg_0502;
    92: op1_11_in26 = reg_0740;
    93: op1_11_in26 = imem03_in[71:68];
    94: op1_11_in26 = reg_0582;
    95: op1_11_in26 = reg_0507;
    default: op1_11_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv26 = 1;
    8: op1_11_inv26 = 1;
    9: op1_11_inv26 = 1;
    11: op1_11_inv26 = 1;
    12: op1_11_inv26 = 1;
    14: op1_11_inv26 = 1;
    17: op1_11_inv26 = 1;
    19: op1_11_inv26 = 1;
    20: op1_11_inv26 = 1;
    22: op1_11_inv26 = 1;
    23: op1_11_inv26 = 1;
    25: op1_11_inv26 = 1;
    26: op1_11_inv26 = 1;
    27: op1_11_inv26 = 1;
    36: op1_11_inv26 = 1;
    39: op1_11_inv26 = 1;
    40: op1_11_inv26 = 1;
    42: op1_11_inv26 = 1;
    47: op1_11_inv26 = 1;
    52: op1_11_inv26 = 1;
    54: op1_11_inv26 = 1;
    57: op1_11_inv26 = 1;
    60: op1_11_inv26 = 1;
    62: op1_11_inv26 = 1;
    64: op1_11_inv26 = 1;
    66: op1_11_inv26 = 1;
    67: op1_11_inv26 = 1;
    75: op1_11_inv26 = 1;
    77: op1_11_inv26 = 1;
    78: op1_11_inv26 = 1;
    82: op1_11_inv26 = 1;
    85: op1_11_inv26 = 1;
    88: op1_11_inv26 = 1;
    89: op1_11_inv26 = 1;
    90: op1_11_inv26 = 1;
    92: op1_11_inv26 = 1;
    95: op1_11_inv26 = 1;
    default: op1_11_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in27 = reg_0550;
    60: op1_11_in27 = reg_0550;
    5: op1_11_in27 = reg_0055;
    6: op1_11_in27 = imem06_in[71:68];
    8: op1_11_in27 = reg_0004;
    9: op1_11_in27 = imem01_in[119:116];
    10: op1_11_in27 = reg_0260;
    11: op1_11_in27 = reg_0501;
    12: op1_11_in27 = imem06_in[95:92];
    14: op1_11_in27 = imem01_in[71:68];
    15: op1_11_in27 = reg_0308;
    16: op1_11_in27 = reg_0028;
    17: op1_11_in27 = imem04_in[55:52];
    29: op1_11_in27 = imem04_in[55:52];
    18: op1_11_in27 = reg_0608;
    19: op1_11_in27 = reg_0529;
    20: op1_11_in27 = reg_0166;
    21: op1_11_in27 = reg_0354;
    22: op1_11_in27 = imem04_in[19:16];
    23: op1_11_in27 = reg_0346;
    24: op1_11_in27 = reg_0286;
    25: op1_11_in27 = reg_0506;
    26: op1_11_in27 = reg_0402;
    27: op1_11_in27 = reg_0140;
    28: op1_11_in27 = reg_0587;
    30: op1_11_in27 = reg_0419;
    31: op1_11_in27 = imem01_in[127:124];
    32: op1_11_in27 = reg_0239;
    33: op1_11_in27 = reg_0491;
    36: op1_11_in27 = reg_0100;
    38: op1_11_in27 = imem04_in[63:60];
    39: op1_11_in27 = reg_0547;
    40: op1_11_in27 = imem05_in[11:8];
    42: op1_11_in27 = reg_0124;
    43: op1_11_in27 = reg_0581;
    44: op1_11_in27 = reg_0721;
    46: op1_11_in27 = reg_0588;
    47: op1_11_in27 = reg_0724;
    49: op1_11_in27 = reg_0144;
    50: op1_11_in27 = reg_0781;
    51: op1_11_in27 = reg_0592;
    52: op1_11_in27 = imem05_in[67:64];
    53: op1_11_in27 = reg_0598;
    54: op1_11_in27 = reg_0295;
    57: op1_11_in27 = reg_0182;
    61: op1_11_in27 = reg_0385;
    62: op1_11_in27 = reg_0593;
    63: op1_11_in27 = reg_0625;
    64: op1_11_in27 = reg_0717;
    66: op1_11_in27 = reg_0705;
    67: op1_11_in27 = reg_0756;
    68: op1_11_in27 = reg_0223;
    70: op1_11_in27 = reg_0785;
    71: op1_11_in27 = reg_0369;
    74: op1_11_in27 = reg_0241;
    75: op1_11_in27 = reg_0559;
    76: op1_11_in27 = reg_0386;
    77: op1_11_in27 = reg_0285;
    78: op1_11_in27 = reg_0583;
    80: op1_11_in27 = reg_0388;
    82: op1_11_in27 = reg_0795;
    83: op1_11_in27 = reg_0098;
    85: op1_11_in27 = reg_0190;
    86: op1_11_in27 = reg_0389;
    95: op1_11_in27 = reg_0389;
    88: op1_11_in27 = reg_0296;
    89: op1_11_in27 = imem07_in[127:124];
    90: op1_11_in27 = reg_0161;
    91: op1_11_in27 = reg_0504;
    92: op1_11_in27 = imem03_in[7:4];
    93: op1_11_in27 = imem03_in[91:88];
    94: op1_11_in27 = reg_0573;
    default: op1_11_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv27 = 1;
    5: op1_11_inv27 = 1;
    8: op1_11_inv27 = 1;
    9: op1_11_inv27 = 1;
    10: op1_11_inv27 = 1;
    11: op1_11_inv27 = 1;
    12: op1_11_inv27 = 1;
    14: op1_11_inv27 = 1;
    16: op1_11_inv27 = 1;
    17: op1_11_inv27 = 1;
    18: op1_11_inv27 = 1;
    20: op1_11_inv27 = 1;
    23: op1_11_inv27 = 1;
    24: op1_11_inv27 = 1;
    25: op1_11_inv27 = 1;
    26: op1_11_inv27 = 1;
    28: op1_11_inv27 = 1;
    29: op1_11_inv27 = 1;
    30: op1_11_inv27 = 1;
    31: op1_11_inv27 = 1;
    32: op1_11_inv27 = 1;
    39: op1_11_inv27 = 1;
    43: op1_11_inv27 = 1;
    44: op1_11_inv27 = 1;
    46: op1_11_inv27 = 1;
    47: op1_11_inv27 = 1;
    52: op1_11_inv27 = 1;
    54: op1_11_inv27 = 1;
    60: op1_11_inv27 = 1;
    64: op1_11_inv27 = 1;
    66: op1_11_inv27 = 1;
    67: op1_11_inv27 = 1;
    68: op1_11_inv27 = 1;
    70: op1_11_inv27 = 1;
    71: op1_11_inv27 = 1;
    74: op1_11_inv27 = 1;
    75: op1_11_inv27 = 1;
    76: op1_11_inv27 = 1;
    80: op1_11_inv27 = 1;
    82: op1_11_inv27 = 1;
    86: op1_11_inv27 = 1;
    89: op1_11_inv27 = 1;
    92: op1_11_inv27 = 1;
    93: op1_11_inv27 = 1;
    default: op1_11_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in28 = reg_0529;
    5: op1_11_in28 = reg_0738;
    6: op1_11_in28 = imem06_in[75:72];
    8: op1_11_in28 = imem04_in[7:4];
    9: op1_11_in28 = reg_0118;
    10: op1_11_in28 = reg_0265;
    11: op1_11_in28 = reg_0513;
    12: op1_11_in28 = imem06_in[103:100];
    14: op1_11_in28 = imem01_in[91:88];
    15: op1_11_in28 = reg_0283;
    16: op1_11_in28 = reg_0753;
    17: op1_11_in28 = imem04_in[67:64];
    18: op1_11_in28 = reg_0623;
    19: op1_11_in28 = reg_0302;
    21: op1_11_in28 = reg_0359;
    22: op1_11_in28 = imem04_in[27:24];
    23: op1_11_in28 = reg_0336;
    24: op1_11_in28 = reg_0065;
    68: op1_11_in28 = reg_0065;
    25: op1_11_in28 = reg_0240;
    26: op1_11_in28 = reg_0386;
    27: op1_11_in28 = imem06_in[39:36];
    28: op1_11_in28 = reg_0593;
    51: op1_11_in28 = reg_0593;
    78: op1_11_in28 = reg_0593;
    29: op1_11_in28 = imem04_in[79:76];
    30: op1_11_in28 = reg_0420;
    31: op1_11_in28 = reg_0759;
    32: op1_11_in28 = reg_0508;
    33: op1_11_in28 = reg_0787;
    36: op1_11_in28 = reg_0109;
    38: op1_11_in28 = imem04_in[95:92];
    39: op1_11_in28 = reg_0273;
    40: op1_11_in28 = imem05_in[23:20];
    42: op1_11_in28 = reg_0112;
    43: op1_11_in28 = reg_0387;
    44: op1_11_in28 = reg_0723;
    46: op1_11_in28 = reg_0590;
    47: op1_11_in28 = reg_0718;
    66: op1_11_in28 = reg_0718;
    49: op1_11_in28 = imem06_in[15:12];
    50: op1_11_in28 = reg_0490;
    52: op1_11_in28 = imem05_in[95:92];
    53: op1_11_in28 = reg_0075;
    54: op1_11_in28 = reg_0053;
    57: op1_11_in28 = reg_0183;
    60: op1_11_in28 = reg_0241;
    61: op1_11_in28 = reg_0572;
    62: op1_11_in28 = reg_0520;
    63: op1_11_in28 = reg_0298;
    64: op1_11_in28 = reg_0711;
    67: op1_11_in28 = reg_0098;
    70: op1_11_in28 = reg_0584;
    71: op1_11_in28 = reg_0578;
    74: op1_11_in28 = reg_0423;
    75: op1_11_in28 = reg_0319;
    76: op1_11_in28 = reg_0309;
    77: op1_11_in28 = reg_0812;
    80: op1_11_in28 = reg_0421;
    82: op1_11_in28 = reg_0550;
    83: op1_11_in28 = reg_0094;
    85: op1_11_in28 = imem01_in[7:4];
    86: op1_11_in28 = reg_0337;
    88: op1_11_in28 = imem05_in[7:4];
    89: op1_11_in28 = reg_0716;
    90: op1_11_in28 = reg_0441;
    91: op1_11_in28 = reg_0673;
    92: op1_11_in28 = imem03_in[23:20];
    93: op1_11_in28 = imem03_in[123:120];
    94: op1_11_in28 = reg_0015;
    95: op1_11_in28 = reg_0395;
    default: op1_11_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_11_inv28 = 1;
    8: op1_11_inv28 = 1;
    10: op1_11_inv28 = 1;
    11: op1_11_inv28 = 1;
    12: op1_11_inv28 = 1;
    14: op1_11_inv28 = 1;
    15: op1_11_inv28 = 1;
    17: op1_11_inv28 = 1;
    24: op1_11_inv28 = 1;
    25: op1_11_inv28 = 1;
    26: op1_11_inv28 = 1;
    27: op1_11_inv28 = 1;
    29: op1_11_inv28 = 1;
    30: op1_11_inv28 = 1;
    32: op1_11_inv28 = 1;
    38: op1_11_inv28 = 1;
    42: op1_11_inv28 = 1;
    44: op1_11_inv28 = 1;
    46: op1_11_inv28 = 1;
    47: op1_11_inv28 = 1;
    49: op1_11_inv28 = 1;
    50: op1_11_inv28 = 1;
    51: op1_11_inv28 = 1;
    53: op1_11_inv28 = 1;
    54: op1_11_inv28 = 1;
    57: op1_11_inv28 = 1;
    60: op1_11_inv28 = 1;
    62: op1_11_inv28 = 1;
    64: op1_11_inv28 = 1;
    67: op1_11_inv28 = 1;
    68: op1_11_inv28 = 1;
    70: op1_11_inv28 = 1;
    71: op1_11_inv28 = 1;
    76: op1_11_inv28 = 1;
    80: op1_11_inv28 = 1;
    82: op1_11_inv28 = 1;
    83: op1_11_inv28 = 1;
    85: op1_11_inv28 = 1;
    86: op1_11_inv28 = 1;
    88: op1_11_inv28 = 1;
    90: op1_11_inv28 = 1;
    94: op1_11_inv28 = 1;
    default: op1_11_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in29 = reg_0539;
    5: op1_11_in29 = reg_0732;
    6: op1_11_in29 = imem06_in[91:88];
    8: op1_11_in29 = imem04_in[47:44];
    9: op1_11_in29 = reg_0120;
    10: op1_11_in29 = reg_0272;
    11: op1_11_in29 = reg_0521;
    12: op1_11_in29 = reg_0629;
    14: op1_11_in29 = imem01_in[99:96];
    15: op1_11_in29 = reg_0289;
    16: op1_11_in29 = reg_0040;
    17: op1_11_in29 = imem04_in[95:92];
    18: op1_11_in29 = reg_0402;
    19: op1_11_in29 = reg_0293;
    21: op1_11_in29 = reg_0329;
    22: op1_11_in29 = imem04_in[59:56];
    23: op1_11_in29 = reg_0092;
    24: op1_11_in29 = reg_0068;
    25: op1_11_in29 = reg_0216;
    26: op1_11_in29 = reg_0399;
    27: op1_11_in29 = imem06_in[55:52];
    28: op1_11_in29 = reg_0597;
    93: op1_11_in29 = reg_0597;
    29: op1_11_in29 = imem04_in[87:84];
    30: op1_11_in29 = reg_0175;
    31: op1_11_in29 = reg_0515;
    53: op1_11_in29 = reg_0515;
    32: op1_11_in29 = reg_0122;
    33: op1_11_in29 = reg_0486;
    36: op1_11_in29 = imem02_in[11:8];
    38: op1_11_in29 = imem04_in[115:112];
    39: op1_11_in29 = reg_0274;
    40: op1_11_in29 = imem05_in[35:32];
    88: op1_11_in29 = imem05_in[35:32];
    42: op1_11_in29 = reg_0102;
    43: op1_11_in29 = reg_0571;
    44: op1_11_in29 = reg_0714;
    46: op1_11_in29 = reg_0391;
    47: op1_11_in29 = reg_0700;
    49: op1_11_in29 = imem06_in[27:24];
    50: op1_11_in29 = reg_0788;
    51: op1_11_in29 = reg_0595;
    52: op1_11_in29 = imem05_in[115:112];
    54: op1_11_in29 = reg_0051;
    57: op1_11_in29 = reg_0170;
    60: op1_11_in29 = reg_0054;
    80: op1_11_in29 = reg_0054;
    61: op1_11_in29 = reg_0000;
    62: op1_11_in29 = reg_0620;
    63: op1_11_in29 = reg_0038;
    64: op1_11_in29 = reg_0707;
    66: op1_11_in29 = reg_0711;
    67: op1_11_in29 = reg_0498;
    68: op1_11_in29 = reg_0622;
    70: op1_11_in29 = reg_0639;
    71: op1_11_in29 = reg_0630;
    74: op1_11_in29 = reg_0574;
    75: op1_11_in29 = reg_0591;
    76: op1_11_in29 = reg_0812;
    77: op1_11_in29 = reg_0148;
    78: op1_11_in29 = reg_0035;
    82: op1_11_in29 = reg_0113;
    83: op1_11_in29 = reg_0093;
    85: op1_11_in29 = imem01_in[11:8];
    86: op1_11_in29 = reg_0227;
    89: op1_11_in29 = reg_0710;
    90: op1_11_in29 = reg_0266;
    91: op1_11_in29 = reg_0592;
    92: op1_11_in29 = imem03_in[27:24];
    94: op1_11_in29 = reg_0799;
    95: op1_11_in29 = reg_0396;
    default: op1_11_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_11_inv29 = 1;
    10: op1_11_inv29 = 1;
    11: op1_11_inv29 = 1;
    15: op1_11_inv29 = 1;
    16: op1_11_inv29 = 1;
    18: op1_11_inv29 = 1;
    21: op1_11_inv29 = 1;
    23: op1_11_inv29 = 1;
    24: op1_11_inv29 = 1;
    31: op1_11_inv29 = 1;
    32: op1_11_inv29 = 1;
    33: op1_11_inv29 = 1;
    36: op1_11_inv29 = 1;
    40: op1_11_inv29 = 1;
    42: op1_11_inv29 = 1;
    43: op1_11_inv29 = 1;
    44: op1_11_inv29 = 1;
    50: op1_11_inv29 = 1;
    51: op1_11_inv29 = 1;
    52: op1_11_inv29 = 1;
    54: op1_11_inv29 = 1;
    57: op1_11_inv29 = 1;
    60: op1_11_inv29 = 1;
    61: op1_11_inv29 = 1;
    63: op1_11_inv29 = 1;
    64: op1_11_inv29 = 1;
    70: op1_11_inv29 = 1;
    74: op1_11_inv29 = 1;
    76: op1_11_inv29 = 1;
    80: op1_11_inv29 = 1;
    82: op1_11_inv29 = 1;
    83: op1_11_inv29 = 1;
    86: op1_11_inv29 = 1;
    90: op1_11_inv29 = 1;
    92: op1_11_inv29 = 1;
    93: op1_11_inv29 = 1;
    94: op1_11_inv29 = 1;
    95: op1_11_inv29 = 1;
    default: op1_11_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_11_in30 = reg_0548;
    5: op1_11_in30 = reg_0735;
    6: op1_11_in30 = imem06_in[99:96];
    8: op1_11_in30 = imem04_in[63:60];
    9: op1_11_in30 = reg_0121;
    10: op1_11_in30 = reg_0261;
    11: op1_11_in30 = reg_0499;
    12: op1_11_in30 = reg_0607;
    14: op1_11_in30 = imem01_in[119:116];
    15: op1_11_in30 = reg_0285;
    16: op1_11_in30 = reg_0038;
    17: op1_11_in30 = imem05_in[11:8];
    18: op1_11_in30 = reg_0381;
    19: op1_11_in30 = reg_0268;
    21: op1_11_in30 = reg_0342;
    22: op1_11_in30 = imem04_in[67:64];
    23: op1_11_in30 = reg_0314;
    24: op1_11_in30 = reg_0071;
    25: op1_11_in30 = reg_0220;
    26: op1_11_in30 = reg_0404;
    27: op1_11_in30 = reg_0628;
    28: op1_11_in30 = reg_0581;
    29: op1_11_in30 = imem04_in[91:88];
    30: op1_11_in30 = reg_0181;
    31: op1_11_in30 = reg_0232;
    32: op1_11_in30 = reg_0118;
    33: op1_11_in30 = reg_0091;
    36: op1_11_in30 = imem02_in[15:12];
    38: op1_11_in30 = imem04_in[119:116];
    39: op1_11_in30 = reg_0306;
    40: op1_11_in30 = imem05_in[43:40];
    42: op1_11_in30 = reg_0114;
    43: op1_11_in30 = reg_0562;
    44: op1_11_in30 = reg_0703;
    46: op1_11_in30 = reg_0568;
    47: op1_11_in30 = reg_0169;
    49: op1_11_in30 = imem06_in[35:32];
    50: op1_11_in30 = reg_0491;
    51: op1_11_in30 = reg_0588;
    52: op1_11_in30 = reg_0483;
    53: op1_11_in30 = reg_0069;
    54: op1_11_in30 = reg_0635;
    57: op1_11_in30 = reg_0158;
    60: op1_11_in30 = reg_0217;
    74: op1_11_in30 = reg_0217;
    80: op1_11_in30 = reg_0217;
    61: op1_11_in30 = reg_0019;
    62: op1_11_in30 = reg_0218;
    63: op1_11_in30 = reg_0260;
    64: op1_11_in30 = reg_0266;
    66: op1_11_in30 = reg_0706;
    67: op1_11_in30 = reg_0093;
    68: op1_11_in30 = reg_0311;
    70: op1_11_in30 = reg_0647;
    71: op1_11_in30 = reg_0654;
    75: op1_11_in30 = reg_0528;
    76: op1_11_in30 = reg_0742;
    77: op1_11_in30 = reg_0150;
    78: op1_11_in30 = reg_0025;
    82: op1_11_in30 = reg_0231;
    83: op1_11_in30 = imem03_in[11:8];
    85: op1_11_in30 = imem01_in[19:16];
    86: op1_11_in30 = reg_0788;
    88: op1_11_in30 = imem05_in[107:104];
    89: op1_11_in30 = reg_0159;
    90: op1_11_in30 = reg_0436;
    91: op1_11_in30 = reg_0675;
    92: op1_11_in30 = imem03_in[31:28];
    93: op1_11_in30 = reg_0367;
    94: op1_11_in30 = reg_0010;
    95: op1_11_in30 = reg_0557;
    default: op1_11_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_11_inv30 = 1;
    5: op1_11_inv30 = 1;
    6: op1_11_inv30 = 1;
    9: op1_11_inv30 = 1;
    15: op1_11_inv30 = 1;
    17: op1_11_inv30 = 1;
    19: op1_11_inv30 = 1;
    22: op1_11_inv30 = 1;
    23: op1_11_inv30 = 1;
    27: op1_11_inv30 = 1;
    28: op1_11_inv30 = 1;
    31: op1_11_inv30 = 1;
    36: op1_11_inv30 = 1;
    38: op1_11_inv30 = 1;
    39: op1_11_inv30 = 1;
    43: op1_11_inv30 = 1;
    46: op1_11_inv30 = 1;
    47: op1_11_inv30 = 1;
    49: op1_11_inv30 = 1;
    50: op1_11_inv30 = 1;
    52: op1_11_inv30 = 1;
    53: op1_11_inv30 = 1;
    57: op1_11_inv30 = 1;
    60: op1_11_inv30 = 1;
    61: op1_11_inv30 = 1;
    62: op1_11_inv30 = 1;
    64: op1_11_inv30 = 1;
    66: op1_11_inv30 = 1;
    68: op1_11_inv30 = 1;
    71: op1_11_inv30 = 1;
    74: op1_11_inv30 = 1;
    75: op1_11_inv30 = 1;
    76: op1_11_inv30 = 1;
    77: op1_11_inv30 = 1;
    82: op1_11_inv30 = 1;
    88: op1_11_inv30 = 1;
    95: op1_11_inv30 = 1;
    default: op1_11_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_11_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_11_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in00 = reg_0531;
    5: op1_12_in00 = reg_0748;
    6: op1_12_in00 = imem06_in[111:108];
    7: op1_12_in00 = imem00_in[67:64];
    8: op1_12_in00 = imem04_in[71:68];
    9: op1_12_in00 = reg_0110;
    10: op1_12_in00 = reg_0142;
    11: op1_12_in00 = reg_0778;
    12: op1_12_in00 = reg_0613;
    13: op1_12_in00 = imem00_in[7:4];
    20: op1_12_in00 = imem00_in[7:4];
    34: op1_12_in00 = imem00_in[7:4];
    35: op1_12_in00 = imem00_in[7:4];
    56: op1_12_in00 = imem00_in[7:4];
    65: op1_12_in00 = imem00_in[7:4];
    14: op1_12_in00 = reg_0496;
    15: op1_12_in00 = reg_0307;
    16: op1_12_in00 = reg_0749;
    17: op1_12_in00 = imem05_in[67:64];
    18: op1_12_in00 = reg_0371;
    19: op1_12_in00 = reg_0286;
    21: op1_12_in00 = reg_0355;
    22: op1_12_in00 = imem04_in[75:72];
    23: op1_12_in00 = reg_0526;
    24: op1_12_in00 = reg_0063;
    3: op1_12_in00 = imem07_in[19:16];
    25: op1_12_in00 = reg_0245;
    2: op1_12_in00 = imem07_in[11:8];
    26: op1_12_in00 = reg_0035;
    27: op1_12_in00 = reg_0604;
    28: op1_12_in00 = reg_0575;
    29: op1_12_in00 = imem04_in[119:116];
    30: op1_12_in00 = imem00_in[11:8];
    37: op1_12_in00 = imem00_in[11:8];
    73: op1_12_in00 = imem00_in[11:8];
    1: op1_12_in00 = imem07_in[39:36];
    31: op1_12_in00 = reg_0505;
    32: op1_12_in00 = reg_0120;
    33: op1_12_in00 = reg_0304;
    50: op1_12_in00 = reg_0304;
    36: op1_12_in00 = imem02_in[23:20];
    38: op1_12_in00 = reg_0552;
    39: op1_12_in00 = reg_0050;
    40: op1_12_in00 = imem05_in[51:48];
    41: op1_12_in00 = imem00_in[27:24];
    69: op1_12_in00 = imem00_in[27:24];
    42: op1_12_in00 = imem02_in[27:24];
    43: op1_12_in00 = reg_0572;
    44: op1_12_in00 = reg_0729;
    45: op1_12_in00 = imem00_in[31:28];
    46: op1_12_in00 = reg_0385;
    47: op1_12_in00 = reg_0173;
    48: op1_12_in00 = reg_0680;
    49: op1_12_in00 = imem06_in[55:52];
    51: op1_12_in00 = reg_0751;
    52: op1_12_in00 = reg_0797;
    53: op1_12_in00 = reg_0288;
    54: op1_12_in00 = reg_0267;
    55: op1_12_in00 = imem00_in[59:56];
    57: op1_12_in00 = reg_0184;
    58: op1_12_in00 = imem00_in[23:20];
    59: op1_12_in00 = imem00_in[43:40];
    60: op1_12_in00 = reg_0234;
    80: op1_12_in00 = reg_0234;
    61: op1_12_in00 = reg_0807;
    62: op1_12_in00 = reg_0368;
    63: op1_12_in00 = reg_0402;
    64: op1_12_in00 = reg_0333;
    90: op1_12_in00 = reg_0333;
    66: op1_12_in00 = reg_0636;
    67: op1_12_in00 = imem03_in[11:8];
    68: op1_12_in00 = reg_0296;
    70: op1_12_in00 = reg_0426;
    71: op1_12_in00 = reg_0775;
    72: op1_12_in00 = imem00_in[15:12];
    87: op1_12_in00 = imem00_in[15:12];
    74: op1_12_in00 = reg_0216;
    75: op1_12_in00 = reg_0357;
    76: op1_12_in00 = reg_0152;
    77: op1_12_in00 = reg_0137;
    78: op1_12_in00 = reg_0663;
    79: op1_12_in00 = imem00_in[35:32];
    81: op1_12_in00 = imem00_in[3:0];
    82: op1_12_in00 = reg_0090;
    83: op1_12_in00 = imem03_in[59:56];
    84: op1_12_in00 = imem00_in[19:16];
    85: op1_12_in00 = imem01_in[67:64];
    86: op1_12_in00 = reg_0146;
    88: op1_12_in00 = imem05_in[111:108];
    89: op1_12_in00 = reg_0166;
    91: op1_12_in00 = reg_0121;
    92: op1_12_in00 = imem03_in[43:40];
    93: op1_12_in00 = reg_0338;
    94: op1_12_in00 = reg_0595;
    95: op1_12_in00 = reg_0418;
    default: op1_12_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv00 = 1;
    5: op1_12_inv00 = 1;
    6: op1_12_inv00 = 1;
    7: op1_12_inv00 = 1;
    9: op1_12_inv00 = 1;
    10: op1_12_inv00 = 1;
    14: op1_12_inv00 = 1;
    16: op1_12_inv00 = 1;
    19: op1_12_inv00 = 1;
    20: op1_12_inv00 = 1;
    21: op1_12_inv00 = 1;
    22: op1_12_inv00 = 1;
    24: op1_12_inv00 = 1;
    2: op1_12_inv00 = 1;
    27: op1_12_inv00 = 1;
    29: op1_12_inv00 = 1;
    1: op1_12_inv00 = 1;
    33: op1_12_inv00 = 1;
    35: op1_12_inv00 = 1;
    36: op1_12_inv00 = 1;
    37: op1_12_inv00 = 1;
    40: op1_12_inv00 = 1;
    42: op1_12_inv00 = 1;
    43: op1_12_inv00 = 1;
    44: op1_12_inv00 = 1;
    45: op1_12_inv00 = 1;
    46: op1_12_inv00 = 1;
    47: op1_12_inv00 = 1;
    51: op1_12_inv00 = 1;
    52: op1_12_inv00 = 1;
    55: op1_12_inv00 = 1;
    56: op1_12_inv00 = 1;
    58: op1_12_inv00 = 1;
    63: op1_12_inv00 = 1;
    66: op1_12_inv00 = 1;
    69: op1_12_inv00 = 1;
    71: op1_12_inv00 = 1;
    73: op1_12_inv00 = 1;
    74: op1_12_inv00 = 1;
    77: op1_12_inv00 = 1;
    78: op1_12_inv00 = 1;
    79: op1_12_inv00 = 1;
    80: op1_12_inv00 = 1;
    81: op1_12_inv00 = 1;
    82: op1_12_inv00 = 1;
    84: op1_12_inv00 = 1;
    85: op1_12_inv00 = 1;
    89: op1_12_inv00 = 1;
    93: op1_12_inv00 = 1;
    94: op1_12_inv00 = 1;
    default: op1_12_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in01 = reg_0303;
    5: op1_12_in01 = reg_0740;
    6: op1_12_in01 = reg_0631;
    7: op1_12_in01 = reg_0693;
    8: op1_12_in01 = imem04_in[75:72];
    9: op1_12_in01 = imem02_in[7:4];
    10: op1_12_in01 = reg_0131;
    11: op1_12_in01 = reg_0515;
    12: op1_12_in01 = reg_0620;
    27: op1_12_in01 = reg_0620;
    78: op1_12_in01 = reg_0620;
    13: op1_12_in01 = imem00_in[11:8];
    14: op1_12_in01 = reg_0520;
    15: op1_12_in01 = reg_0059;
    29: op1_12_in01 = reg_0059;
    16: op1_12_in01 = imem07_in[7:4];
    17: op1_12_in01 = reg_0792;
    18: op1_12_in01 = reg_0375;
    19: op1_12_in01 = reg_0258;
    20: op1_12_in01 = imem00_in[59:56];
    35: op1_12_in01 = imem00_in[59:56];
    21: op1_12_in01 = reg_0347;
    22: op1_12_in01 = imem04_in[79:76];
    23: op1_12_in01 = imem03_in[3:0];
    24: op1_12_in01 = reg_0069;
    3: op1_12_in01 = imem07_in[47:44];
    25: op1_12_in01 = reg_0238;
    2: op1_12_in01 = imem07_in[23:20];
    26: op1_12_in01 = reg_0816;
    28: op1_12_in01 = reg_0568;
    30: op1_12_in01 = imem00_in[23:20];
    72: op1_12_in01 = imem00_in[23:20];
    1: op1_12_in01 = imem07_in[75:72];
    31: op1_12_in01 = reg_0218;
    32: op1_12_in01 = reg_0102;
    33: op1_12_in01 = reg_0279;
    34: op1_12_in01 = imem00_in[27:24];
    37: op1_12_in01 = imem00_in[27:24];
    36: op1_12_in01 = imem02_in[107:104];
    38: op1_12_in01 = reg_0536;
    39: op1_12_in01 = reg_0257;
    40: op1_12_in01 = imem05_in[59:56];
    41: op1_12_in01 = imem00_in[39:36];
    65: op1_12_in01 = imem00_in[39:36];
    73: op1_12_in01 = imem00_in[39:36];
    84: op1_12_in01 = imem00_in[39:36];
    87: op1_12_in01 = imem00_in[39:36];
    42: op1_12_in01 = imem02_in[39:36];
    43: op1_12_in01 = reg_0396;
    44: op1_12_in01 = reg_0718;
    45: op1_12_in01 = imem00_in[35:32];
    46: op1_12_in01 = reg_0392;
    48: op1_12_in01 = reg_0688;
    49: op1_12_in01 = imem06_in[67:64];
    50: op1_12_in01 = reg_0309;
    51: op1_12_in01 = reg_0749;
    52: op1_12_in01 = reg_0788;
    53: op1_12_in01 = imem05_in[7:4];
    54: op1_12_in01 = reg_0448;
    55: op1_12_in01 = imem00_in[63:60];
    56: op1_12_in01 = imem00_in[55:52];
    58: op1_12_in01 = imem00_in[87:84];
    59: op1_12_in01 = imem00_in[67:64];
    60: op1_12_in01 = reg_0105;
    61: op1_12_in01 = reg_0802;
    62: op1_12_in01 = imem07_in[27:24];
    63: op1_12_in01 = reg_0630;
    64: op1_12_in01 = reg_0434;
    66: op1_12_in01 = reg_0438;
    67: op1_12_in01 = imem03_in[15:12];
    68: op1_12_in01 = imem05_in[19:16];
    69: op1_12_in01 = imem00_in[51:48];
    70: op1_12_in01 = reg_0356;
    71: op1_12_in01 = reg_0748;
    74: op1_12_in01 = reg_0220;
    75: op1_12_in01 = reg_0751;
    76: op1_12_in01 = reg_0825;
    77: op1_12_in01 = imem06_in[51:48];
    79: op1_12_in01 = imem00_in[71:68];
    80: op1_12_in01 = reg_0424;
    81: op1_12_in01 = imem00_in[7:4];
    82: op1_12_in01 = reg_0782;
    83: op1_12_in01 = reg_0582;
    85: op1_12_in01 = imem01_in[87:84];
    86: op1_12_in01 = reg_0113;
    88: op1_12_in01 = imem05_in[127:124];
    89: op1_12_in01 = reg_0295;
    90: op1_12_in01 = reg_0446;
    91: op1_12_in01 = imem02_in[19:16];
    92: op1_12_in01 = imem03_in[59:56];
    93: op1_12_in01 = reg_0559;
    94: op1_12_in01 = reg_0028;
    95: op1_12_in01 = reg_0290;
    default: op1_12_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv01 = 1;
    5: op1_12_inv01 = 1;
    6: op1_12_inv01 = 1;
    7: op1_12_inv01 = 1;
    10: op1_12_inv01 = 1;
    11: op1_12_inv01 = 1;
    13: op1_12_inv01 = 1;
    14: op1_12_inv01 = 1;
    16: op1_12_inv01 = 1;
    17: op1_12_inv01 = 1;
    18: op1_12_inv01 = 1;
    19: op1_12_inv01 = 1;
    22: op1_12_inv01 = 1;
    24: op1_12_inv01 = 1;
    25: op1_12_inv01 = 1;
    2: op1_12_inv01 = 1;
    26: op1_12_inv01 = 1;
    27: op1_12_inv01 = 1;
    29: op1_12_inv01 = 1;
    30: op1_12_inv01 = 1;
    33: op1_12_inv01 = 1;
    38: op1_12_inv01 = 1;
    40: op1_12_inv01 = 1;
    41: op1_12_inv01 = 1;
    46: op1_12_inv01 = 1;
    50: op1_12_inv01 = 1;
    54: op1_12_inv01 = 1;
    55: op1_12_inv01 = 1;
    56: op1_12_inv01 = 1;
    58: op1_12_inv01 = 1;
    63: op1_12_inv01 = 1;
    67: op1_12_inv01 = 1;
    71: op1_12_inv01 = 1;
    73: op1_12_inv01 = 1;
    75: op1_12_inv01 = 1;
    77: op1_12_inv01 = 1;
    78: op1_12_inv01 = 1;
    80: op1_12_inv01 = 1;
    82: op1_12_inv01 = 1;
    83: op1_12_inv01 = 1;
    84: op1_12_inv01 = 1;
    87: op1_12_inv01 = 1;
    89: op1_12_inv01 = 1;
    90: op1_12_inv01 = 1;
    91: op1_12_inv01 = 1;
    94: op1_12_inv01 = 1;
    95: op1_12_inv01 = 1;
    default: op1_12_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in02 = reg_0304;
    5: op1_12_in02 = reg_0733;
    6: op1_12_in02 = reg_0577;
    12: op1_12_in02 = reg_0577;
    7: op1_12_in02 = reg_0676;
    8: op1_12_in02 = imem04_in[91:88];
    9: op1_12_in02 = imem02_in[15:12];
    10: op1_12_in02 = imem06_in[19:16];
    11: op1_12_in02 = reg_0510;
    13: op1_12_in02 = imem00_in[35:32];
    14: op1_12_in02 = reg_0515;
    15: op1_12_in02 = reg_0061;
    39: op1_12_in02 = reg_0061;
    16: op1_12_in02 = imem07_in[47:44];
    17: op1_12_in02 = reg_0796;
    18: op1_12_in02 = reg_0028;
    19: op1_12_in02 = reg_0062;
    20: op1_12_in02 = imem00_in[63:60];
    21: op1_12_in02 = reg_0092;
    22: op1_12_in02 = imem04_in[95:92];
    23: op1_12_in02 = imem03_in[27:24];
    24: op1_12_in02 = imem05_in[39:36];
    3: op1_12_in02 = imem07_in[103:100];
    25: op1_12_in02 = reg_0508;
    2: op1_12_in02 = reg_0175;
    26: op1_12_in02 = reg_0036;
    27: op1_12_in02 = reg_0608;
    28: op1_12_in02 = reg_0388;
    29: op1_12_in02 = reg_0545;
    30: op1_12_in02 = imem00_in[51:48];
    41: op1_12_in02 = imem00_in[51:48];
    87: op1_12_in02 = imem00_in[51:48];
    1: op1_12_in02 = imem07_in[95:92];
    31: op1_12_in02 = reg_0240;
    32: op1_12_in02 = imem02_in[11:8];
    33: op1_12_in02 = reg_0742;
    34: op1_12_in02 = imem00_in[31:28];
    72: op1_12_in02 = imem00_in[31:28];
    35: op1_12_in02 = imem00_in[107:104];
    36: op1_12_in02 = imem02_in[111:108];
    37: op1_12_in02 = imem00_in[43:40];
    38: op1_12_in02 = reg_0523;
    40: op1_12_in02 = imem05_in[83:80];
    42: op1_12_in02 = imem02_in[63:60];
    43: op1_12_in02 = reg_0374;
    44: op1_12_in02 = reg_0707;
    45: op1_12_in02 = imem00_in[59:56];
    46: op1_12_in02 = reg_0562;
    48: op1_12_in02 = reg_0687;
    49: op1_12_in02 = reg_0299;
    50: op1_12_in02 = reg_0732;
    86: op1_12_in02 = reg_0732;
    51: op1_12_in02 = reg_0373;
    52: op1_12_in02 = reg_0492;
    53: op1_12_in02 = imem05_in[11:8];
    54: op1_12_in02 = reg_0435;
    55: op1_12_in02 = imem00_in[95:92];
    56: op1_12_in02 = imem00_in[83:80];
    58: op1_12_in02 = reg_0681;
    59: op1_12_in02 = imem00_in[75:72];
    79: op1_12_in02 = imem00_in[75:72];
    60: op1_12_in02 = reg_0108;
    61: op1_12_in02 = imem04_in[63:60];
    62: op1_12_in02 = imem07_in[35:32];
    63: op1_12_in02 = reg_0580;
    64: op1_12_in02 = reg_0440;
    65: op1_12_in02 = imem00_in[55:52];
    69: op1_12_in02 = imem00_in[55:52];
    66: op1_12_in02 = reg_0161;
    67: op1_12_in02 = imem03_in[35:32];
    68: op1_12_in02 = imem05_in[27:24];
    70: op1_12_in02 = reg_0363;
    71: op1_12_in02 = reg_0035;
    73: op1_12_in02 = imem00_in[87:84];
    74: op1_12_in02 = reg_0425;
    75: op1_12_in02 = reg_0398;
    76: op1_12_in02 = imem06_in[79:76];
    77: op1_12_in02 = imem06_in[119:116];
    78: op1_12_in02 = reg_0657;
    80: op1_12_in02 = reg_0243;
    81: op1_12_in02 = imem00_in[15:12];
    82: op1_12_in02 = reg_0517;
    83: op1_12_in02 = reg_0751;
    84: op1_12_in02 = imem00_in[47:44];
    85: op1_12_in02 = imem01_in[91:88];
    88: op1_12_in02 = reg_0736;
    89: op1_12_in02 = reg_0447;
    90: op1_12_in02 = reg_0084;
    91: op1_12_in02 = imem02_in[99:96];
    92: op1_12_in02 = imem03_in[79:76];
    93: op1_12_in02 = reg_0494;
    94: op1_12_in02 = reg_0564;
    95: op1_12_in02 = reg_0806;
    default: op1_12_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv02 = 1;
    6: op1_12_inv02 = 1;
    8: op1_12_inv02 = 1;
    9: op1_12_inv02 = 1;
    10: op1_12_inv02 = 1;
    11: op1_12_inv02 = 1;
    13: op1_12_inv02 = 1;
    15: op1_12_inv02 = 1;
    18: op1_12_inv02 = 1;
    19: op1_12_inv02 = 1;
    21: op1_12_inv02 = 1;
    25: op1_12_inv02 = 1;
    2: op1_12_inv02 = 1;
    26: op1_12_inv02 = 1;
    27: op1_12_inv02 = 1;
    29: op1_12_inv02 = 1;
    31: op1_12_inv02 = 1;
    33: op1_12_inv02 = 1;
    38: op1_12_inv02 = 1;
    39: op1_12_inv02 = 1;
    40: op1_12_inv02 = 1;
    41: op1_12_inv02 = 1;
    43: op1_12_inv02 = 1;
    44: op1_12_inv02 = 1;
    46: op1_12_inv02 = 1;
    49: op1_12_inv02 = 1;
    50: op1_12_inv02 = 1;
    51: op1_12_inv02 = 1;
    53: op1_12_inv02 = 1;
    54: op1_12_inv02 = 1;
    55: op1_12_inv02 = 1;
    56: op1_12_inv02 = 1;
    58: op1_12_inv02 = 1;
    59: op1_12_inv02 = 1;
    61: op1_12_inv02 = 1;
    62: op1_12_inv02 = 1;
    64: op1_12_inv02 = 1;
    69: op1_12_inv02 = 1;
    73: op1_12_inv02 = 1;
    74: op1_12_inv02 = 1;
    77: op1_12_inv02 = 1;
    79: op1_12_inv02 = 1;
    84: op1_12_inv02 = 1;
    85: op1_12_inv02 = 1;
    87: op1_12_inv02 = 1;
    89: op1_12_inv02 = 1;
    90: op1_12_inv02 = 1;
    default: op1_12_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in03 = reg_0293;
    5: op1_12_in03 = reg_0582;
    6: op1_12_in03 = reg_0379;
    7: op1_12_in03 = reg_0689;
    8: op1_12_in03 = imem04_in[95:92];
    9: op1_12_in03 = imem02_in[31:28];
    10: op1_12_in03 = imem06_in[75:72];
    11: op1_12_in03 = reg_0755;
    12: op1_12_in03 = reg_0332;
    13: op1_12_in03 = imem00_in[51:48];
    14: op1_12_in03 = reg_0232;
    15: op1_12_in03 = reg_0062;
    16: op1_12_in03 = imem07_in[51:48];
    17: op1_12_in03 = reg_0493;
    18: op1_12_in03 = reg_0753;
    19: op1_12_in03 = reg_0067;
    20: op1_12_in03 = imem00_in[71:68];
    37: op1_12_in03 = imem00_in[71:68];
    72: op1_12_in03 = imem00_in[71:68];
    87: op1_12_in03 = imem00_in[71:68];
    21: op1_12_in03 = reg_0541;
    22: op1_12_in03 = imem04_in[127:124];
    23: op1_12_in03 = imem03_in[107:104];
    24: op1_12_in03 = imem05_in[47:44];
    3: op1_12_in03 = imem07_in[127:124];
    25: op1_12_in03 = reg_0105;
    2: op1_12_in03 = reg_0161;
    26: op1_12_in03 = reg_0749;
    27: op1_12_in03 = reg_0622;
    28: op1_12_in03 = reg_0517;
    29: op1_12_in03 = reg_0316;
    30: op1_12_in03 = imem00_in[67:64];
    1: op1_12_in03 = imem07_in[111:108];
    31: op1_12_in03 = reg_0503;
    32: op1_12_in03 = imem02_in[15:12];
    33: op1_12_in03 = reg_0527;
    34: op1_12_in03 = imem00_in[47:44];
    35: op1_12_in03 = reg_0676;
    36: op1_12_in03 = reg_0653;
    38: op1_12_in03 = reg_0556;
    39: op1_12_in03 = imem05_in[55:52];
    40: op1_12_in03 = reg_0488;
    41: op1_12_in03 = imem00_in[55:52];
    84: op1_12_in03 = imem00_in[55:52];
    42: op1_12_in03 = imem02_in[79:76];
    43: op1_12_in03 = reg_0001;
    44: op1_12_in03 = reg_0334;
    45: op1_12_in03 = imem00_in[75:72];
    69: op1_12_in03 = imem00_in[75:72];
    46: op1_12_in03 = reg_0376;
    48: op1_12_in03 = reg_0453;
    49: op1_12_in03 = reg_0624;
    50: op1_12_in03 = reg_0277;
    51: op1_12_in03 = reg_0392;
    52: op1_12_in03 = reg_0795;
    53: op1_12_in03 = imem05_in[23:20];
    54: op1_12_in03 = reg_0181;
    55: op1_12_in03 = reg_0682;
    56: op1_12_in03 = imem00_in[119:116];
    58: op1_12_in03 = reg_0694;
    59: op1_12_in03 = imem00_in[79:76];
    60: op1_12_in03 = reg_0674;
    61: op1_12_in03 = imem04_in[103:100];
    62: op1_12_in03 = imem07_in[59:56];
    63: op1_12_in03 = reg_0764;
    64: op1_12_in03 = reg_0444;
    65: op1_12_in03 = imem00_in[95:92];
    66: op1_12_in03 = reg_0162;
    67: op1_12_in03 = imem03_in[55:52];
    68: op1_12_in03 = imem05_in[91:88];
    70: op1_12_in03 = reg_0590;
    71: op1_12_in03 = reg_0515;
    73: op1_12_in03 = imem00_in[115:112];
    74: op1_12_in03 = reg_0506;
    75: op1_12_in03 = reg_0747;
    76: op1_12_in03 = reg_0299;
    77: op1_12_in03 = reg_0404;
    78: op1_12_in03 = reg_0664;
    79: op1_12_in03 = reg_0696;
    80: op1_12_in03 = reg_0120;
    81: op1_12_in03 = imem00_in[23:20];
    82: op1_12_in03 = reg_0245;
    83: op1_12_in03 = reg_0417;
    85: op1_12_in03 = imem01_in[119:116];
    86: op1_12_in03 = imem05_in[11:8];
    88: op1_12_in03 = reg_0135;
    89: op1_12_in03 = reg_0439;
    90: op1_12_in03 = reg_0267;
    91: op1_12_in03 = imem02_in[119:116];
    92: op1_12_in03 = reg_0597;
    93: op1_12_in03 = reg_0595;
    94: op1_12_in03 = reg_0568;
    95: op1_12_in03 = imem04_in[11:8];
    default: op1_12_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv03 = 1;
    7: op1_12_inv03 = 1;
    8: op1_12_inv03 = 1;
    11: op1_12_inv03 = 1;
    12: op1_12_inv03 = 1;
    14: op1_12_inv03 = 1;
    15: op1_12_inv03 = 1;
    16: op1_12_inv03 = 1;
    17: op1_12_inv03 = 1;
    19: op1_12_inv03 = 1;
    21: op1_12_inv03 = 1;
    23: op1_12_inv03 = 1;
    3: op1_12_inv03 = 1;
    26: op1_12_inv03 = 1;
    27: op1_12_inv03 = 1;
    1: op1_12_inv03 = 1;
    31: op1_12_inv03 = 1;
    34: op1_12_inv03 = 1;
    35: op1_12_inv03 = 1;
    36: op1_12_inv03 = 1;
    41: op1_12_inv03 = 1;
    42: op1_12_inv03 = 1;
    43: op1_12_inv03 = 1;
    46: op1_12_inv03 = 1;
    48: op1_12_inv03 = 1;
    49: op1_12_inv03 = 1;
    59: op1_12_inv03 = 1;
    60: op1_12_inv03 = 1;
    64: op1_12_inv03 = 1;
    65: op1_12_inv03 = 1;
    68: op1_12_inv03 = 1;
    74: op1_12_inv03 = 1;
    75: op1_12_inv03 = 1;
    77: op1_12_inv03 = 1;
    79: op1_12_inv03 = 1;
    82: op1_12_inv03 = 1;
    83: op1_12_inv03 = 1;
    84: op1_12_inv03 = 1;
    87: op1_12_inv03 = 1;
    89: op1_12_inv03 = 1;
    93: op1_12_inv03 = 1;
    94: op1_12_inv03 = 1;
    95: op1_12_inv03 = 1;
    default: op1_12_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in04 = reg_0290;
    5: op1_12_in04 = reg_0579;
    6: op1_12_in04 = reg_0371;
    7: op1_12_in04 = reg_0684;
    8: op1_12_in04 = reg_0530;
    21: op1_12_in04 = reg_0530;
    9: op1_12_in04 = imem02_in[47:44];
    10: op1_12_in04 = reg_0614;
    11: op1_12_in04 = reg_0507;
    93: op1_12_in04 = reg_0507;
    12: op1_12_in04 = reg_0375;
    13: op1_12_in04 = imem00_in[111:108];
    72: op1_12_in04 = imem00_in[111:108];
    14: op1_12_in04 = reg_0216;
    15: op1_12_in04 = reg_0065;
    16: op1_12_in04 = imem07_in[95:92];
    17: op1_12_in04 = reg_0782;
    18: op1_12_in04 = reg_0815;
    19: op1_12_in04 = reg_0289;
    20: op1_12_in04 = imem00_in[83:80];
    22: op1_12_in04 = reg_0059;
    23: op1_12_in04 = imem03_in[119:116];
    24: op1_12_in04 = imem05_in[59:56];
    3: op1_12_in04 = reg_0424;
    25: op1_12_in04 = reg_0116;
    2: op1_12_in04 = reg_0167;
    26: op1_12_in04 = imem07_in[47:44];
    27: op1_12_in04 = reg_0615;
    28: op1_12_in04 = reg_0747;
    29: op1_12_in04 = reg_0544;
    30: op1_12_in04 = imem00_in[75:72];
    87: op1_12_in04 = imem00_in[75:72];
    31: op1_12_in04 = reg_0237;
    32: op1_12_in04 = imem02_in[63:60];
    33: op1_12_in04 = reg_0086;
    34: op1_12_in04 = imem00_in[99:96];
    35: op1_12_in04 = reg_0463;
    36: op1_12_in04 = reg_0639;
    37: op1_12_in04 = imem00_in[79:76];
    38: op1_12_in04 = reg_0303;
    39: op1_12_in04 = imem05_in[123:120];
    40: op1_12_in04 = reg_0789;
    41: op1_12_in04 = imem00_in[107:104];
    42: op1_12_in04 = imem02_in[83:80];
    43: op1_12_in04 = reg_0013;
    44: op1_12_in04 = reg_0441;
    45: op1_12_in04 = imem00_in[91:88];
    46: op1_12_in04 = reg_0393;
    48: op1_12_in04 = reg_0455;
    49: op1_12_in04 = reg_0817;
    50: op1_12_in04 = reg_0149;
    51: op1_12_in04 = reg_0006;
    52: op1_12_in04 = reg_0494;
    53: op1_12_in04 = imem05_in[27:24];
    54: op1_12_in04 = reg_0161;
    55: op1_12_in04 = reg_0685;
    56: op1_12_in04 = imem00_in[123:120];
    58: op1_12_in04 = reg_0680;
    59: op1_12_in04 = imem00_in[87:84];
    60: op1_12_in04 = imem02_in[55:52];
    61: op1_12_in04 = imem04_in[107:104];
    62: op1_12_in04 = imem07_in[107:104];
    63: op1_12_in04 = reg_0028;
    64: op1_12_in04 = reg_0437;
    65: op1_12_in04 = imem00_in[115:112];
    66: op1_12_in04 = reg_0183;
    67: op1_12_in04 = imem03_in[59:56];
    68: op1_12_in04 = imem05_in[107:104];
    69: op1_12_in04 = reg_0695;
    73: op1_12_in04 = reg_0695;
    70: op1_12_in04 = reg_0314;
    71: op1_12_in04 = reg_0573;
    74: op1_12_in04 = reg_0073;
    75: op1_12_in04 = reg_0623;
    76: op1_12_in04 = reg_0577;
    77: op1_12_in04 = reg_0618;
    78: op1_12_in04 = reg_0787;
    79: op1_12_in04 = reg_0612;
    80: op1_12_in04 = reg_0108;
    81: op1_12_in04 = imem00_in[27:24];
    82: op1_12_in04 = reg_0138;
    83: op1_12_in04 = reg_0396;
    84: op1_12_in04 = imem00_in[71:68];
    85: op1_12_in04 = reg_0497;
    86: op1_12_in04 = imem05_in[39:36];
    88: op1_12_in04 = reg_0090;
    89: op1_12_in04 = reg_0442;
    90: op1_12_in04 = reg_0268;
    91: op1_12_in04 = imem02_in[123:120];
    92: op1_12_in04 = reg_0575;
    94: op1_12_in04 = reg_0483;
    95: op1_12_in04 = imem04_in[39:36];
    default: op1_12_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv04 = 1;
    8: op1_12_inv04 = 1;
    10: op1_12_inv04 = 1;
    12: op1_12_inv04 = 1;
    14: op1_12_inv04 = 1;
    15: op1_12_inv04 = 1;
    17: op1_12_inv04 = 1;
    21: op1_12_inv04 = 1;
    22: op1_12_inv04 = 1;
    23: op1_12_inv04 = 1;
    3: op1_12_inv04 = 1;
    2: op1_12_inv04 = 1;
    26: op1_12_inv04 = 1;
    30: op1_12_inv04 = 1;
    38: op1_12_inv04 = 1;
    39: op1_12_inv04 = 1;
    41: op1_12_inv04 = 1;
    43: op1_12_inv04 = 1;
    46: op1_12_inv04 = 1;
    48: op1_12_inv04 = 1;
    49: op1_12_inv04 = 1;
    50: op1_12_inv04 = 1;
    55: op1_12_inv04 = 1;
    58: op1_12_inv04 = 1;
    59: op1_12_inv04 = 1;
    60: op1_12_inv04 = 1;
    61: op1_12_inv04 = 1;
    62: op1_12_inv04 = 1;
    64: op1_12_inv04 = 1;
    68: op1_12_inv04 = 1;
    70: op1_12_inv04 = 1;
    74: op1_12_inv04 = 1;
    76: op1_12_inv04 = 1;
    78: op1_12_inv04 = 1;
    80: op1_12_inv04 = 1;
    81: op1_12_inv04 = 1;
    82: op1_12_inv04 = 1;
    83: op1_12_inv04 = 1;
    84: op1_12_inv04 = 1;
    85: op1_12_inv04 = 1;
    87: op1_12_inv04 = 1;
    88: op1_12_inv04 = 1;
    89: op1_12_inv04 = 1;
    90: op1_12_inv04 = 1;
    91: op1_12_inv04 = 1;
    93: op1_12_inv04 = 1;
    94: op1_12_inv04 = 1;
    default: op1_12_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in05 = reg_0291;
    5: op1_12_in05 = reg_0569;
    6: op1_12_in05 = reg_0375;
    7: op1_12_in05 = reg_0690;
    8: op1_12_in05 = reg_0539;
    9: op1_12_in05 = imem02_in[75:72];
    10: op1_12_in05 = reg_0610;
    11: op1_12_in05 = reg_0241;
    12: op1_12_in05 = reg_0315;
    13: op1_12_in05 = reg_0670;
    14: op1_12_in05 = reg_0236;
    15: op1_12_in05 = reg_0067;
    16: op1_12_in05 = imem07_in[107:104];
    17: op1_12_in05 = reg_0267;
    89: op1_12_in05 = reg_0267;
    18: op1_12_in05 = reg_0748;
    19: op1_12_in05 = reg_0255;
    20: op1_12_in05 = imem00_in[107:104];
    21: op1_12_in05 = reg_0096;
    22: op1_12_in05 = reg_0544;
    23: op1_12_in05 = reg_0582;
    24: op1_12_in05 = imem05_in[119:116];
    3: op1_12_in05 = reg_0430;
    25: op1_12_in05 = reg_0102;
    2: op1_12_in05 = reg_0163;
    26: op1_12_in05 = imem07_in[79:76];
    27: op1_12_in05 = reg_0409;
    28: op1_12_in05 = reg_0386;
    29: op1_12_in05 = reg_0328;
    30: op1_12_in05 = imem00_in[91:88];
    31: op1_12_in05 = reg_0245;
    32: op1_12_in05 = imem02_in[95:92];
    33: op1_12_in05 = reg_0148;
    34: op1_12_in05 = imem00_in[127:124];
    87: op1_12_in05 = imem00_in[127:124];
    35: op1_12_in05 = reg_0455;
    36: op1_12_in05 = reg_0648;
    37: op1_12_in05 = imem00_in[87:84];
    38: op1_12_in05 = reg_0294;
    39: op1_12_in05 = reg_0798;
    40: op1_12_in05 = reg_0785;
    52: op1_12_in05 = reg_0785;
    41: op1_12_in05 = imem00_in[123:120];
    45: op1_12_in05 = imem00_in[123:120];
    42: op1_12_in05 = imem02_in[87:84];
    43: op1_12_in05 = reg_0805;
    44: op1_12_in05 = reg_0061;
    46: op1_12_in05 = reg_0389;
    48: op1_12_in05 = reg_0476;
    49: op1_12_in05 = reg_0020;
    50: op1_12_in05 = reg_0136;
    51: op1_12_in05 = reg_0811;
    83: op1_12_in05 = reg_0811;
    53: op1_12_in05 = imem05_in[87:84];
    54: op1_12_in05 = reg_0159;
    55: op1_12_in05 = reg_0698;
    56: op1_12_in05 = reg_0685;
    58: op1_12_in05 = reg_0454;
    59: op1_12_in05 = imem00_in[111:108];
    60: op1_12_in05 = imem02_in[71:68];
    61: op1_12_in05 = imem04_in[115:112];
    62: op1_12_in05 = reg_0720;
    63: op1_12_in05 = reg_0534;
    64: op1_12_in05 = reg_0448;
    65: op1_12_in05 = imem00_in[119:116];
    66: op1_12_in05 = reg_0168;
    67: op1_12_in05 = imem03_in[63:60];
    68: op1_12_in05 = imem05_in[115:112];
    69: op1_12_in05 = reg_0697;
    70: op1_12_in05 = reg_0770;
    71: op1_12_in05 = reg_0787;
    72: op1_12_in05 = reg_0682;
    73: op1_12_in05 = reg_0612;
    74: op1_12_in05 = reg_0601;
    75: op1_12_in05 = reg_0649;
    76: op1_12_in05 = reg_0762;
    77: op1_12_in05 = reg_0242;
    78: op1_12_in05 = reg_0661;
    79: op1_12_in05 = reg_0658;
    80: op1_12_in05 = reg_0660;
    81: op1_12_in05 = imem00_in[31:28];
    82: op1_12_in05 = reg_0257;
    84: op1_12_in05 = imem00_in[75:72];
    85: op1_12_in05 = reg_0668;
    86: op1_12_in05 = imem05_in[59:56];
    88: op1_12_in05 = reg_0326;
    90: op1_12_in05 = reg_0175;
    91: op1_12_in05 = reg_0642;
    92: op1_12_in05 = reg_0568;
    93: op1_12_in05 = reg_0321;
    94: op1_12_in05 = reg_0490;
    95: op1_12_in05 = imem04_in[43:40];
    default: op1_12_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv05 = 1;
    5: op1_12_inv05 = 1;
    6: op1_12_inv05 = 1;
    7: op1_12_inv05 = 1;
    8: op1_12_inv05 = 1;
    9: op1_12_inv05 = 1;
    10: op1_12_inv05 = 1;
    11: op1_12_inv05 = 1;
    14: op1_12_inv05 = 1;
    15: op1_12_inv05 = 1;
    16: op1_12_inv05 = 1;
    18: op1_12_inv05 = 1;
    19: op1_12_inv05 = 1;
    22: op1_12_inv05 = 1;
    23: op1_12_inv05 = 1;
    27: op1_12_inv05 = 1;
    28: op1_12_inv05 = 1;
    29: op1_12_inv05 = 1;
    30: op1_12_inv05 = 1;
    31: op1_12_inv05 = 1;
    32: op1_12_inv05 = 1;
    33: op1_12_inv05 = 1;
    34: op1_12_inv05 = 1;
    36: op1_12_inv05 = 1;
    37: op1_12_inv05 = 1;
    39: op1_12_inv05 = 1;
    41: op1_12_inv05 = 1;
    43: op1_12_inv05 = 1;
    46: op1_12_inv05 = 1;
    48: op1_12_inv05 = 1;
    49: op1_12_inv05 = 1;
    51: op1_12_inv05 = 1;
    55: op1_12_inv05 = 1;
    56: op1_12_inv05 = 1;
    63: op1_12_inv05 = 1;
    64: op1_12_inv05 = 1;
    66: op1_12_inv05 = 1;
    69: op1_12_inv05 = 1;
    71: op1_12_inv05 = 1;
    73: op1_12_inv05 = 1;
    74: op1_12_inv05 = 1;
    76: op1_12_inv05 = 1;
    78: op1_12_inv05 = 1;
    80: op1_12_inv05 = 1;
    83: op1_12_inv05 = 1;
    84: op1_12_inv05 = 1;
    87: op1_12_inv05 = 1;
    88: op1_12_inv05 = 1;
    89: op1_12_inv05 = 1;
    95: op1_12_inv05 = 1;
    default: op1_12_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in06 = reg_0062;
    5: op1_12_in06 = reg_0592;
    6: op1_12_in06 = reg_0367;
    12: op1_12_in06 = reg_0367;
    7: op1_12_in06 = reg_0671;
    8: op1_12_in06 = reg_0555;
    9: op1_12_in06 = imem02_in[95:92];
    10: op1_12_in06 = reg_0613;
    11: op1_12_in06 = reg_0216;
    13: op1_12_in06 = reg_0690;
    14: op1_12_in06 = reg_0504;
    15: op1_12_in06 = reg_0057;
    16: op1_12_in06 = reg_0728;
    17: op1_12_in06 = reg_0262;
    18: op1_12_in06 = imem07_in[55:52];
    19: op1_12_in06 = reg_0288;
    20: op1_12_in06 = imem00_in[115:112];
    21: op1_12_in06 = reg_0540;
    22: op1_12_in06 = reg_0545;
    61: op1_12_in06 = reg_0545;
    23: op1_12_in06 = reg_0573;
    24: op1_12_in06 = imem05_in[127:124];
    68: op1_12_in06 = imem05_in[127:124];
    3: op1_12_in06 = reg_0447;
    25: op1_12_in06 = reg_0114;
    2: op1_12_in06 = reg_0164;
    26: op1_12_in06 = imem07_in[87:84];
    27: op1_12_in06 = reg_0401;
    28: op1_12_in06 = reg_0006;
    29: op1_12_in06 = reg_0556;
    30: op1_12_in06 = imem00_in[103:100];
    31: op1_12_in06 = reg_0508;
    32: op1_12_in06 = imem02_in[103:100];
    33: op1_12_in06 = reg_0143;
    34: op1_12_in06 = reg_0682;
    59: op1_12_in06 = reg_0682;
    65: op1_12_in06 = reg_0682;
    35: op1_12_in06 = reg_0464;
    36: op1_12_in06 = reg_0636;
    37: op1_12_in06 = imem00_in[95:92];
    38: op1_12_in06 = reg_0274;
    39: op1_12_in06 = reg_0797;
    40: op1_12_in06 = reg_0737;
    41: op1_12_in06 = reg_0683;
    42: op1_12_in06 = imem02_in[119:116];
    43: op1_12_in06 = reg_0009;
    44: op1_12_in06 = reg_0180;
    90: op1_12_in06 = reg_0180;
    45: op1_12_in06 = reg_0697;
    46: op1_12_in06 = reg_0000;
    48: op1_12_in06 = reg_0467;
    49: op1_12_in06 = reg_0286;
    50: op1_12_in06 = reg_0128;
    51: op1_12_in06 = reg_0001;
    52: op1_12_in06 = reg_0304;
    53: op1_12_in06 = imem05_in[91:88];
    54: op1_12_in06 = reg_0182;
    55: op1_12_in06 = reg_0494;
    56: op1_12_in06 = reg_0686;
    58: op1_12_in06 = reg_0480;
    60: op1_12_in06 = imem02_in[79:76];
    62: op1_12_in06 = reg_0721;
    63: op1_12_in06 = reg_0368;
    64: op1_12_in06 = reg_0175;
    67: op1_12_in06 = imem03_in[67:64];
    69: op1_12_in06 = reg_0492;
    70: op1_12_in06 = reg_0082;
    71: op1_12_in06 = reg_0752;
    72: op1_12_in06 = reg_0698;
    73: op1_12_in06 = reg_0684;
    74: op1_12_in06 = reg_0678;
    75: op1_12_in06 = reg_0570;
    76: op1_12_in06 = reg_0815;
    77: op1_12_in06 = reg_0369;
    78: op1_12_in06 = reg_0256;
    79: op1_12_in06 = reg_0255;
    80: op1_12_in06 = reg_0677;
    81: op1_12_in06 = imem00_in[43:40];
    82: op1_12_in06 = reg_0824;
    83: op1_12_in06 = imem04_in[3:0];
    84: op1_12_in06 = imem00_in[87:84];
    85: op1_12_in06 = reg_0772;
    86: op1_12_in06 = imem05_in[67:64];
    87: op1_12_in06 = reg_0612;
    88: op1_12_in06 = reg_0538;
    89: op1_12_in06 = reg_0438;
    91: op1_12_in06 = reg_0392;
    92: op1_12_in06 = reg_0002;
    93: op1_12_in06 = reg_0646;
    94: op1_12_in06 = reg_0562;
    95: op1_12_in06 = imem04_in[59:56];
    default: op1_12_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv06 = 1;
    7: op1_12_inv06 = 1;
    8: op1_12_inv06 = 1;
    9: op1_12_inv06 = 1;
    13: op1_12_inv06 = 1;
    14: op1_12_inv06 = 1;
    16: op1_12_inv06 = 1;
    17: op1_12_inv06 = 1;
    18: op1_12_inv06 = 1;
    19: op1_12_inv06 = 1;
    20: op1_12_inv06 = 1;
    21: op1_12_inv06 = 1;
    22: op1_12_inv06 = 1;
    23: op1_12_inv06 = 1;
    3: op1_12_inv06 = 1;
    2: op1_12_inv06 = 1;
    28: op1_12_inv06 = 1;
    34: op1_12_inv06 = 1;
    35: op1_12_inv06 = 1;
    39: op1_12_inv06 = 1;
    41: op1_12_inv06 = 1;
    43: op1_12_inv06 = 1;
    44: op1_12_inv06 = 1;
    45: op1_12_inv06 = 1;
    46: op1_12_inv06 = 1;
    48: op1_12_inv06 = 1;
    56: op1_12_inv06 = 1;
    59: op1_12_inv06 = 1;
    61: op1_12_inv06 = 1;
    62: op1_12_inv06 = 1;
    67: op1_12_inv06 = 1;
    69: op1_12_inv06 = 1;
    70: op1_12_inv06 = 1;
    72: op1_12_inv06 = 1;
    75: op1_12_inv06 = 1;
    77: op1_12_inv06 = 1;
    80: op1_12_inv06 = 1;
    81: op1_12_inv06 = 1;
    82: op1_12_inv06 = 1;
    83: op1_12_inv06 = 1;
    86: op1_12_inv06 = 1;
    88: op1_12_inv06 = 1;
    92: op1_12_inv06 = 1;
    94: op1_12_inv06 = 1;
    default: op1_12_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in07 = reg_0041;
    5: op1_12_in07 = reg_0584;
    6: op1_12_in07 = imem07_in[3:0];
    7: op1_12_in07 = reg_0678;
    80: op1_12_in07 = reg_0678;
    8: op1_12_in07 = reg_0549;
    9: op1_12_in07 = reg_0656;
    10: op1_12_in07 = reg_0619;
    11: op1_12_in07 = reg_0247;
    12: op1_12_in07 = reg_0368;
    13: op1_12_in07 = reg_0668;
    14: op1_12_in07 = reg_0245;
    15: op1_12_in07 = imem05_in[23:20];
    16: op1_12_in07 = reg_0730;
    17: op1_12_in07 = reg_0259;
    19: op1_12_in07 = reg_0259;
    18: op1_12_in07 = imem07_in[75:72];
    20: op1_12_in07 = reg_0689;
    21: op1_12_in07 = imem03_in[3:0];
    22: op1_12_in07 = reg_0315;
    23: op1_12_in07 = reg_0587;
    24: op1_12_in07 = reg_0488;
    3: op1_12_in07 = reg_0445;
    25: op1_12_in07 = reg_0329;
    2: op1_12_in07 = reg_0185;
    26: op1_12_in07 = imem07_in[119:116];
    27: op1_12_in07 = reg_0813;
    28: op1_12_in07 = reg_0808;
    46: op1_12_in07 = reg_0808;
    29: op1_12_in07 = reg_0293;
    30: op1_12_in07 = imem00_in[119:116];
    37: op1_12_in07 = imem00_in[119:116];
    31: op1_12_in07 = reg_0125;
    32: op1_12_in07 = imem02_in[123:120];
    42: op1_12_in07 = imem02_in[123:120];
    33: op1_12_in07 = reg_0140;
    34: op1_12_in07 = reg_0679;
    45: op1_12_in07 = reg_0679;
    35: op1_12_in07 = reg_0476;
    36: op1_12_in07 = reg_0357;
    38: op1_12_in07 = reg_0257;
    39: op1_12_in07 = reg_0492;
    40: op1_12_in07 = reg_0085;
    41: op1_12_in07 = reg_0696;
    43: op1_12_in07 = reg_0004;
    44: op1_12_in07 = reg_0167;
    48: op1_12_in07 = reg_0459;
    49: op1_12_in07 = reg_0609;
    50: op1_12_in07 = reg_0134;
    51: op1_12_in07 = reg_0805;
    52: op1_12_in07 = reg_0102;
    53: op1_12_in07 = imem05_in[111:108];
    54: op1_12_in07 = reg_0160;
    55: op1_12_in07 = reg_0680;
    56: op1_12_in07 = reg_0255;
    58: op1_12_in07 = reg_0210;
    59: op1_12_in07 = reg_0697;
    60: op1_12_in07 = imem02_in[91:88];
    61: op1_12_in07 = reg_0516;
    62: op1_12_in07 = reg_0703;
    63: op1_12_in07 = imem07_in[15:12];
    64: op1_12_in07 = reg_0161;
    65: op1_12_in07 = reg_0683;
    67: op1_12_in07 = imem03_in[71:68];
    68: op1_12_in07 = reg_0091;
    69: op1_12_in07 = reg_0684;
    70: op1_12_in07 = reg_0539;
    71: op1_12_in07 = imem07_in[67:64];
    72: op1_12_in07 = reg_0686;
    73: op1_12_in07 = reg_0633;
    74: op1_12_in07 = imem02_in[95:92];
    75: op1_12_in07 = reg_0019;
    76: op1_12_in07 = reg_0817;
    77: op1_12_in07 = reg_0377;
    78: op1_12_in07 = reg_0089;
    90: op1_12_in07 = reg_0089;
    79: op1_12_in07 = reg_0467;
    81: op1_12_in07 = imem00_in[47:44];
    82: op1_12_in07 = imem06_in[71:68];
    83: op1_12_in07 = imem04_in[115:112];
    84: op1_12_in07 = imem00_in[99:96];
    85: op1_12_in07 = reg_0741;
    86: op1_12_in07 = imem05_in[99:96];
    87: op1_12_in07 = reg_0698;
    88: op1_12_in07 = reg_0552;
    89: op1_12_in07 = reg_0268;
    91: op1_12_in07 = reg_0086;
    92: op1_12_in07 = reg_0319;
    93: op1_12_in07 = reg_0747;
    94: op1_12_in07 = reg_0637;
    95: op1_12_in07 = imem04_in[71:68];
    default: op1_12_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv07 = 1;
    9: op1_12_inv07 = 1;
    10: op1_12_inv07 = 1;
    12: op1_12_inv07 = 1;
    14: op1_12_inv07 = 1;
    16: op1_12_inv07 = 1;
    18: op1_12_inv07 = 1;
    19: op1_12_inv07 = 1;
    25: op1_12_inv07 = 1;
    2: op1_12_inv07 = 1;
    26: op1_12_inv07 = 1;
    27: op1_12_inv07 = 1;
    28: op1_12_inv07 = 1;
    30: op1_12_inv07 = 1;
    31: op1_12_inv07 = 1;
    32: op1_12_inv07 = 1;
    33: op1_12_inv07 = 1;
    37: op1_12_inv07 = 1;
    40: op1_12_inv07 = 1;
    46: op1_12_inv07 = 1;
    49: op1_12_inv07 = 1;
    51: op1_12_inv07 = 1;
    52: op1_12_inv07 = 1;
    53: op1_12_inv07 = 1;
    54: op1_12_inv07 = 1;
    55: op1_12_inv07 = 1;
    56: op1_12_inv07 = 1;
    64: op1_12_inv07 = 1;
    65: op1_12_inv07 = 1;
    67: op1_12_inv07 = 1;
    68: op1_12_inv07 = 1;
    69: op1_12_inv07 = 1;
    70: op1_12_inv07 = 1;
    72: op1_12_inv07 = 1;
    74: op1_12_inv07 = 1;
    75: op1_12_inv07 = 1;
    77: op1_12_inv07 = 1;
    80: op1_12_inv07 = 1;
    82: op1_12_inv07 = 1;
    83: op1_12_inv07 = 1;
    84: op1_12_inv07 = 1;
    92: op1_12_inv07 = 1;
    93: op1_12_inv07 = 1;
    94: op1_12_inv07 = 1;
    95: op1_12_inv07 = 1;
    default: op1_12_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in08 = imem05_in[3:0];
    5: op1_12_in08 = reg_0593;
    6: op1_12_in08 = imem07_in[27:24];
    7: op1_12_in08 = reg_0476;
    8: op1_12_in08 = reg_0533;
    9: op1_12_in08 = reg_0639;
    10: op1_12_in08 = reg_0608;
    11: op1_12_in08 = reg_0118;
    12: op1_12_in08 = reg_0039;
    13: op1_12_in08 = reg_0675;
    14: op1_12_in08 = reg_0238;
    15: op1_12_in08 = imem05_in[47:44];
    16: op1_12_in08 = reg_0731;
    17: op1_12_in08 = reg_0526;
    18: op1_12_in08 = imem07_in[99:96];
    71: op1_12_in08 = imem07_in[99:96];
    19: op1_12_in08 = reg_0262;
    20: op1_12_in08 = reg_0686;
    21: op1_12_in08 = imem03_in[23:20];
    22: op1_12_in08 = reg_0087;
    23: op1_12_in08 = reg_0360;
    24: op1_12_in08 = reg_0785;
    39: op1_12_in08 = reg_0785;
    3: op1_12_in08 = reg_0443;
    25: op1_12_in08 = reg_0335;
    2: op1_12_in08 = reg_0168;
    26: op1_12_in08 = reg_0710;
    27: op1_12_in08 = reg_0819;
    28: op1_12_in08 = reg_0804;
    29: op1_12_in08 = reg_0295;
    30: op1_12_in08 = reg_0695;
    31: op1_12_in08 = reg_0114;
    32: op1_12_in08 = reg_0645;
    33: op1_12_in08 = imem06_in[15:12];
    34: op1_12_in08 = reg_0674;
    35: op1_12_in08 = reg_0472;
    36: op1_12_in08 = reg_0361;
    37: op1_12_in08 = reg_0685;
    38: op1_12_in08 = reg_0074;
    40: op1_12_in08 = reg_0260;
    41: op1_12_in08 = reg_0698;
    42: op1_12_in08 = reg_0650;
    43: op1_12_in08 = imem04_in[15:12];
    44: op1_12_in08 = reg_0159;
    45: op1_12_in08 = reg_0669;
    46: op1_12_in08 = reg_0810;
    48: op1_12_in08 = reg_0452;
    49: op1_12_in08 = reg_0298;
    76: op1_12_in08 = reg_0298;
    50: op1_12_in08 = reg_0144;
    51: op1_12_in08 = reg_0802;
    52: op1_12_in08 = reg_0276;
    53: op1_12_in08 = reg_0798;
    54: op1_12_in08 = reg_0164;
    55: op1_12_in08 = reg_0688;
    56: op1_12_in08 = reg_0117;
    72: op1_12_in08 = reg_0117;
    58: op1_12_in08 = reg_0193;
    59: op1_12_in08 = reg_0658;
    60: op1_12_in08 = imem02_in[95:92];
    61: op1_12_in08 = reg_0615;
    62: op1_12_in08 = reg_0713;
    63: op1_12_in08 = imem07_in[123:120];
    64: op1_12_in08 = reg_0162;
    65: op1_12_in08 = reg_0492;
    67: op1_12_in08 = imem03_in[111:108];
    68: op1_12_in08 = reg_0792;
    69: op1_12_in08 = reg_0749;
    70: op1_12_in08 = imem03_in[31:28];
    73: op1_12_in08 = reg_0450;
    74: op1_12_in08 = imem02_in[115:112];
    75: op1_12_in08 = reg_0013;
    77: op1_12_in08 = reg_0563;
    78: op1_12_in08 = reg_0165;
    79: op1_12_in08 = reg_0470;
    80: op1_12_in08 = imem02_in[11:8];
    81: op1_12_in08 = imem00_in[51:48];
    82: op1_12_in08 = imem06_in[87:84];
    83: op1_12_in08 = reg_0537;
    84: op1_12_in08 = imem00_in[103:100];
    85: op1_12_in08 = reg_0385;
    86: op1_12_in08 = imem05_in[123:120];
    87: op1_12_in08 = reg_0684;
    88: op1_12_in08 = reg_0309;
    89: op1_12_in08 = reg_0175;
    90: op1_12_in08 = reg_0182;
    91: op1_12_in08 = reg_0656;
    92: op1_12_in08 = reg_0294;
    93: op1_12_in08 = reg_0319;
    94: op1_12_in08 = reg_0649;
    95: op1_12_in08 = imem04_in[79:76];
    default: op1_12_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv08 = 1;
    5: op1_12_inv08 = 1;
    6: op1_12_inv08 = 1;
    7: op1_12_inv08 = 1;
    11: op1_12_inv08 = 1;
    19: op1_12_inv08 = 1;
    21: op1_12_inv08 = 1;
    23: op1_12_inv08 = 1;
    24: op1_12_inv08 = 1;
    25: op1_12_inv08 = 1;
    2: op1_12_inv08 = 1;
    26: op1_12_inv08 = 1;
    31: op1_12_inv08 = 1;
    33: op1_12_inv08 = 1;
    35: op1_12_inv08 = 1;
    36: op1_12_inv08 = 1;
    39: op1_12_inv08 = 1;
    44: op1_12_inv08 = 1;
    45: op1_12_inv08 = 1;
    49: op1_12_inv08 = 1;
    50: op1_12_inv08 = 1;
    51: op1_12_inv08 = 1;
    52: op1_12_inv08 = 1;
    53: op1_12_inv08 = 1;
    54: op1_12_inv08 = 1;
    55: op1_12_inv08 = 1;
    58: op1_12_inv08 = 1;
    59: op1_12_inv08 = 1;
    60: op1_12_inv08 = 1;
    61: op1_12_inv08 = 1;
    62: op1_12_inv08 = 1;
    64: op1_12_inv08 = 1;
    65: op1_12_inv08 = 1;
    68: op1_12_inv08 = 1;
    70: op1_12_inv08 = 1;
    76: op1_12_inv08 = 1;
    78: op1_12_inv08 = 1;
    79: op1_12_inv08 = 1;
    83: op1_12_inv08 = 1;
    86: op1_12_inv08 = 1;
    87: op1_12_inv08 = 1;
    88: op1_12_inv08 = 1;
    89: op1_12_inv08 = 1;
    90: op1_12_inv08 = 1;
    93: op1_12_inv08 = 1;
    94: op1_12_inv08 = 1;
    95: op1_12_inv08 = 1;
    default: op1_12_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in09 = imem05_in[15:12];
    5: op1_12_in09 = reg_0580;
    6: op1_12_in09 = imem07_in[47:44];
    7: op1_12_in09 = reg_0466;
    8: op1_12_in09 = reg_0301;
    9: op1_12_in09 = reg_0651;
    10: op1_12_in09 = reg_0627;
    11: op1_12_in09 = reg_0119;
    12: op1_12_in09 = reg_0035;
    13: op1_12_in09 = reg_0687;
    14: op1_12_in09 = reg_0243;
    15: op1_12_in09 = imem05_in[51:48];
    16: op1_12_in09 = reg_0714;
    17: op1_12_in09 = reg_0734;
    18: op1_12_in09 = imem07_in[103:100];
    19: op1_12_in09 = reg_0264;
    20: op1_12_in09 = reg_0679;
    21: op1_12_in09 = imem03_in[87:84];
    22: op1_12_in09 = reg_0056;
    23: op1_12_in09 = reg_0343;
    24: op1_12_in09 = reg_0495;
    3: op1_12_in09 = reg_0448;
    25: op1_12_in09 = reg_0330;
    2: op1_12_in09 = reg_0171;
    26: op1_12_in09 = reg_0726;
    27: op1_12_in09 = reg_0816;
    28: op1_12_in09 = reg_0009;
    29: op1_12_in09 = reg_0050;
    30: op1_12_in09 = reg_0697;
    31: op1_12_in09 = reg_0109;
    32: op1_12_in09 = reg_0655;
    33: op1_12_in09 = imem06_in[43:40];
    34: op1_12_in09 = reg_0450;
    35: op1_12_in09 = reg_0456;
    36: op1_12_in09 = reg_0351;
    37: op1_12_in09 = reg_0690;
    38: op1_12_in09 = reg_0792;
    39: op1_12_in09 = reg_0794;
    40: op1_12_in09 = reg_0132;
    41: op1_12_in09 = reg_0684;
    42: op1_12_in09 = reg_0654;
    43: op1_12_in09 = imem04_in[35:32];
    44: op1_12_in09 = reg_0157;
    45: op1_12_in09 = reg_0454;
    46: op1_12_in09 = imem04_in[3:0];
    48: op1_12_in09 = reg_0214;
    49: op1_12_in09 = reg_0265;
    50: op1_12_in09 = imem06_in[15:12];
    51: op1_12_in09 = imem04_in[19:16];
    52: op1_12_in09 = reg_0744;
    65: op1_12_in09 = reg_0744;
    53: op1_12_in09 = reg_0491;
    88: op1_12_in09 = reg_0491;
    55: op1_12_in09 = reg_0461;
    56: op1_12_in09 = reg_0680;
    59: op1_12_in09 = reg_0680;
    58: op1_12_in09 = reg_0194;
    60: op1_12_in09 = imem02_in[111:108];
    61: op1_12_in09 = reg_0431;
    62: op1_12_in09 = reg_0267;
    63: op1_12_in09 = imem07_in[127:124];
    64: op1_12_in09 = reg_0167;
    67: op1_12_in09 = imem03_in[127:124];
    68: op1_12_in09 = reg_0256;
    69: op1_12_in09 = reg_0691;
    70: op1_12_in09 = imem03_in[79:76];
    71: op1_12_in09 = imem07_in[123:120];
    72: op1_12_in09 = reg_0407;
    73: op1_12_in09 = reg_0469;
    74: op1_12_in09 = reg_0584;
    75: op1_12_in09 = reg_0807;
    76: op1_12_in09 = reg_0404;
    77: op1_12_in09 = reg_0818;
    78: op1_12_in09 = reg_0717;
    79: op1_12_in09 = reg_0478;
    80: op1_12_in09 = imem02_in[43:40];
    81: op1_12_in09 = imem00_in[63:60];
    82: op1_12_in09 = imem06_in[91:88];
    83: op1_12_in09 = reg_0060;
    84: op1_12_in09 = imem00_in[123:120];
    85: op1_12_in09 = reg_0102;
    86: op1_12_in09 = reg_0149;
    87: op1_12_in09 = reg_0686;
    89: op1_12_in09 = reg_0116;
    90: op1_12_in09 = reg_0228;
    91: op1_12_in09 = reg_0059;
    92: op1_12_in09 = reg_0290;
    93: op1_12_in09 = reg_0244;
    94: op1_12_in09 = reg_0271;
    95: op1_12_in09 = imem04_in[87:84];
    default: op1_12_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv09 = 1;
    11: op1_12_inv09 = 1;
    12: op1_12_inv09 = 1;
    13: op1_12_inv09 = 1;
    14: op1_12_inv09 = 1;
    16: op1_12_inv09 = 1;
    17: op1_12_inv09 = 1;
    18: op1_12_inv09 = 1;
    21: op1_12_inv09 = 1;
    22: op1_12_inv09 = 1;
    23: op1_12_inv09 = 1;
    24: op1_12_inv09 = 1;
    25: op1_12_inv09 = 1;
    2: op1_12_inv09 = 1;
    26: op1_12_inv09 = 1;
    28: op1_12_inv09 = 1;
    29: op1_12_inv09 = 1;
    32: op1_12_inv09 = 1;
    33: op1_12_inv09 = 1;
    36: op1_12_inv09 = 1;
    37: op1_12_inv09 = 1;
    39: op1_12_inv09 = 1;
    43: op1_12_inv09 = 1;
    50: op1_12_inv09 = 1;
    51: op1_12_inv09 = 1;
    53: op1_12_inv09 = 1;
    56: op1_12_inv09 = 1;
    61: op1_12_inv09 = 1;
    62: op1_12_inv09 = 1;
    65: op1_12_inv09 = 1;
    69: op1_12_inv09 = 1;
    70: op1_12_inv09 = 1;
    72: op1_12_inv09 = 1;
    73: op1_12_inv09 = 1;
    74: op1_12_inv09 = 1;
    76: op1_12_inv09 = 1;
    77: op1_12_inv09 = 1;
    78: op1_12_inv09 = 1;
    81: op1_12_inv09 = 1;
    87: op1_12_inv09 = 1;
    88: op1_12_inv09 = 1;
    89: op1_12_inv09 = 1;
    94: op1_12_inv09 = 1;
    default: op1_12_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in10 = imem05_in[55:52];
    5: op1_12_in10 = reg_0578;
    6: op1_12_in10 = imem07_in[63:60];
    7: op1_12_in10 = reg_0471;
    8: op1_12_in10 = reg_0305;
    9: op1_12_in10 = reg_0648;
    10: op1_12_in10 = reg_0601;
    11: op1_12_in10 = reg_0108;
    12: op1_12_in10 = reg_0040;
    13: op1_12_in10 = reg_0460;
    73: op1_12_in10 = reg_0460;
    14: op1_12_in10 = reg_0219;
    15: op1_12_in10 = imem05_in[83:80];
    16: op1_12_in10 = reg_0715;
    17: op1_12_in10 = reg_0132;
    18: op1_12_in10 = imem07_in[111:108];
    19: op1_12_in10 = reg_0488;
    20: op1_12_in10 = reg_0691;
    87: op1_12_in10 = reg_0691;
    21: op1_12_in10 = imem03_in[127:124];
    22: op1_12_in10 = reg_0083;
    23: op1_12_in10 = reg_0808;
    24: op1_12_in10 = reg_0787;
    3: op1_12_in10 = reg_0180;
    25: op1_12_in10 = reg_0655;
    26: op1_12_in10 = reg_0714;
    27: op1_12_in10 = reg_0748;
    28: op1_12_in10 = imem04_in[27:24];
    51: op1_12_in10 = imem04_in[27:24];
    29: op1_12_in10 = reg_0284;
    30: op1_12_in10 = reg_0679;
    31: op1_12_in10 = reg_0117;
    32: op1_12_in10 = reg_0637;
    33: op1_12_in10 = imem06_in[79:76];
    34: op1_12_in10 = reg_0451;
    35: op1_12_in10 = reg_0191;
    36: op1_12_in10 = reg_0343;
    37: op1_12_in10 = reg_0699;
    38: op1_12_in10 = reg_0490;
    39: op1_12_in10 = reg_0783;
    40: op1_12_in10 = reg_0140;
    41: op1_12_in10 = reg_0670;
    42: op1_12_in10 = reg_0660;
    43: op1_12_in10 = imem04_in[67:64];
    45: op1_12_in10 = reg_0466;
    46: op1_12_in10 = imem04_in[15:12];
    48: op1_12_in10 = reg_0187;
    49: op1_12_in10 = reg_0278;
    50: op1_12_in10 = imem06_in[27:24];
    52: op1_12_in10 = reg_0145;
    53: op1_12_in10 = reg_0795;
    55: op1_12_in10 = reg_0477;
    56: op1_12_in10 = reg_0476;
    58: op1_12_in10 = reg_0205;
    59: op1_12_in10 = reg_0465;
    60: op1_12_in10 = imem02_in[115:112];
    61: op1_12_in10 = reg_0610;
    62: op1_12_in10 = reg_0165;
    63: op1_12_in10 = reg_0704;
    64: op1_12_in10 = reg_0168;
    65: op1_12_in10 = reg_0658;
    67: op1_12_in10 = reg_0596;
    68: op1_12_in10 = reg_0226;
    69: op1_12_in10 = reg_0692;
    72: op1_12_in10 = reg_0692;
    70: op1_12_in10 = reg_0589;
    71: op1_12_in10 = reg_0721;
    74: op1_12_in10 = reg_0656;
    75: op1_12_in10 = reg_0800;
    76: op1_12_in10 = reg_0293;
    77: op1_12_in10 = reg_0767;
    78: op1_12_in10 = reg_0100;
    79: op1_12_in10 = reg_0214;
    80: op1_12_in10 = imem02_in[55:52];
    81: op1_12_in10 = imem00_in[67:64];
    82: op1_12_in10 = imem06_in[127:124];
    83: op1_12_in10 = reg_0536;
    84: op1_12_in10 = reg_0689;
    85: op1_12_in10 = reg_0131;
    86: op1_12_in10 = reg_0742;
    88: op1_12_in10 = reg_0229;
    89: op1_12_in10 = reg_0236;
    90: op1_12_in10 = reg_0325;
    91: op1_12_in10 = reg_0594;
    92: op1_12_in10 = reg_0004;
    93: op1_12_in10 = imem04_in[11:8];
    94: op1_12_in10 = reg_0002;
    95: op1_12_in10 = imem04_in[91:88];
    default: op1_12_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv10 = 1;
    5: op1_12_inv10 = 1;
    6: op1_12_inv10 = 1;
    11: op1_12_inv10 = 1;
    12: op1_12_inv10 = 1;
    15: op1_12_inv10 = 1;
    17: op1_12_inv10 = 1;
    18: op1_12_inv10 = 1;
    19: op1_12_inv10 = 1;
    23: op1_12_inv10 = 1;
    24: op1_12_inv10 = 1;
    3: op1_12_inv10 = 1;
    25: op1_12_inv10 = 1;
    26: op1_12_inv10 = 1;
    30: op1_12_inv10 = 1;
    31: op1_12_inv10 = 1;
    32: op1_12_inv10 = 1;
    33: op1_12_inv10 = 1;
    37: op1_12_inv10 = 1;
    40: op1_12_inv10 = 1;
    41: op1_12_inv10 = 1;
    42: op1_12_inv10 = 1;
    45: op1_12_inv10 = 1;
    49: op1_12_inv10 = 1;
    50: op1_12_inv10 = 1;
    51: op1_12_inv10 = 1;
    55: op1_12_inv10 = 1;
    56: op1_12_inv10 = 1;
    61: op1_12_inv10 = 1;
    62: op1_12_inv10 = 1;
    63: op1_12_inv10 = 1;
    65: op1_12_inv10 = 1;
    68: op1_12_inv10 = 1;
    69: op1_12_inv10 = 1;
    72: op1_12_inv10 = 1;
    75: op1_12_inv10 = 1;
    76: op1_12_inv10 = 1;
    77: op1_12_inv10 = 1;
    78: op1_12_inv10 = 1;
    79: op1_12_inv10 = 1;
    82: op1_12_inv10 = 1;
    84: op1_12_inv10 = 1;
    86: op1_12_inv10 = 1;
    87: op1_12_inv10 = 1;
    91: op1_12_inv10 = 1;
    93: op1_12_inv10 = 1;
    94: op1_12_inv10 = 1;
    default: op1_12_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in11 = imem05_in[79:76];
    5: op1_12_in11 = reg_0360;
    6: op1_12_in11 = imem07_in[111:108];
    7: op1_12_in11 = reg_0452;
    8: op1_12_in11 = reg_0282;
    9: op1_12_in11 = reg_0638;
    10: op1_12_in11 = reg_0382;
    11: op1_12_in11 = reg_0102;
    12: op1_12_in11 = reg_0817;
    13: op1_12_in11 = reg_0471;
    14: op1_12_in11 = reg_0103;
    15: op1_12_in11 = imem05_in[95:92];
    16: op1_12_in11 = reg_0442;
    17: op1_12_in11 = reg_0145;
    18: op1_12_in11 = imem07_in[119:116];
    19: op1_12_in11 = reg_0790;
    20: op1_12_in11 = reg_0669;
    21: op1_12_in11 = reg_0598;
    22: op1_12_in11 = reg_0305;
    23: op1_12_in11 = reg_0004;
    24: op1_12_in11 = reg_0279;
    3: op1_12_in11 = reg_0161;
    62: op1_12_in11 = reg_0161;
    25: op1_12_in11 = reg_0656;
    26: op1_12_in11 = reg_0702;
    27: op1_12_in11 = reg_0037;
    28: op1_12_in11 = imem04_in[31:28];
    29: op1_12_in11 = reg_0278;
    30: op1_12_in11 = reg_0476;
    34: op1_12_in11 = reg_0476;
    31: op1_12_in11 = imem02_in[7:4];
    32: op1_12_in11 = reg_0358;
    33: op1_12_in11 = reg_0631;
    35: op1_12_in11 = reg_0189;
    36: op1_12_in11 = reg_0347;
    37: op1_12_in11 = reg_0455;
    59: op1_12_in11 = reg_0455;
    38: op1_12_in11 = reg_0484;
    39: op1_12_in11 = reg_0784;
    40: op1_12_in11 = reg_0137;
    86: op1_12_in11 = reg_0137;
    41: op1_12_in11 = reg_0668;
    42: op1_12_in11 = reg_0657;
    43: op1_12_in11 = imem04_in[75:72];
    45: op1_12_in11 = reg_0470;
    55: op1_12_in11 = reg_0470;
    72: op1_12_in11 = reg_0470;
    46: op1_12_in11 = imem04_in[23:20];
    48: op1_12_in11 = reg_0193;
    49: op1_12_in11 = reg_0317;
    50: op1_12_in11 = imem06_in[31:28];
    51: op1_12_in11 = imem04_in[63:60];
    52: op1_12_in11 = reg_0138;
    53: op1_12_in11 = reg_0493;
    56: op1_12_in11 = reg_0462;
    58: op1_12_in11 = reg_0190;
    60: op1_12_in11 = reg_0651;
    61: op1_12_in11 = reg_0078;
    63: op1_12_in11 = reg_0708;
    65: op1_12_in11 = reg_0688;
    87: op1_12_in11 = reg_0688;
    67: op1_12_in11 = reg_0331;
    68: op1_12_in11 = reg_0793;
    69: op1_12_in11 = reg_0463;
    70: op1_12_in11 = reg_0597;
    71: op1_12_in11 = reg_0714;
    73: op1_12_in11 = reg_0467;
    74: op1_12_in11 = reg_0753;
    75: op1_12_in11 = reg_0008;
    76: op1_12_in11 = reg_0265;
    77: op1_12_in11 = reg_0661;
    78: op1_12_in11 = reg_0729;
    79: op1_12_in11 = reg_0188;
    80: op1_12_in11 = imem02_in[67:64];
    81: op1_12_in11 = imem00_in[71:68];
    82: op1_12_in11 = reg_0625;
    83: op1_12_in11 = reg_0249;
    84: op1_12_in11 = reg_0634;
    85: op1_12_in11 = reg_0388;
    88: op1_12_in11 = reg_0288;
    89: op1_12_in11 = reg_0426;
    90: op1_12_in11 = reg_0178;
    91: op1_12_in11 = reg_0365;
    92: op1_12_in11 = imem04_in[19:16];
    93: op1_12_in11 = imem04_in[43:40];
    94: op1_12_in11 = reg_0418;
    95: op1_12_in11 = imem04_in[107:104];
    default: op1_12_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv11 = 1;
    7: op1_12_inv11 = 1;
    8: op1_12_inv11 = 1;
    9: op1_12_inv11 = 1;
    12: op1_12_inv11 = 1;
    13: op1_12_inv11 = 1;
    21: op1_12_inv11 = 1;
    22: op1_12_inv11 = 1;
    25: op1_12_inv11 = 1;
    26: op1_12_inv11 = 1;
    28: op1_12_inv11 = 1;
    29: op1_12_inv11 = 1;
    31: op1_12_inv11 = 1;
    33: op1_12_inv11 = 1;
    34: op1_12_inv11 = 1;
    35: op1_12_inv11 = 1;
    36: op1_12_inv11 = 1;
    38: op1_12_inv11 = 1;
    42: op1_12_inv11 = 1;
    46: op1_12_inv11 = 1;
    48: op1_12_inv11 = 1;
    51: op1_12_inv11 = 1;
    52: op1_12_inv11 = 1;
    53: op1_12_inv11 = 1;
    56: op1_12_inv11 = 1;
    60: op1_12_inv11 = 1;
    62: op1_12_inv11 = 1;
    65: op1_12_inv11 = 1;
    67: op1_12_inv11 = 1;
    68: op1_12_inv11 = 1;
    69: op1_12_inv11 = 1;
    71: op1_12_inv11 = 1;
    75: op1_12_inv11 = 1;
    78: op1_12_inv11 = 1;
    79: op1_12_inv11 = 1;
    80: op1_12_inv11 = 1;
    81: op1_12_inv11 = 1;
    84: op1_12_inv11 = 1;
    85: op1_12_inv11 = 1;
    86: op1_12_inv11 = 1;
    87: op1_12_inv11 = 1;
    88: op1_12_inv11 = 1;
    91: op1_12_inv11 = 1;
    94: op1_12_inv11 = 1;
    default: op1_12_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in12 = imem05_in[119:116];
    15: op1_12_in12 = imem05_in[119:116];
    5: op1_12_in12 = reg_0370;
    6: op1_12_in12 = reg_0728;
    7: op1_12_in12 = reg_0187;
    72: op1_12_in12 = reg_0187;
    8: op1_12_in12 = reg_0285;
    9: op1_12_in12 = reg_0667;
    10: op1_12_in12 = reg_0403;
    11: op1_12_in12 = reg_0101;
    12: op1_12_in12 = reg_0037;
    13: op1_12_in12 = reg_0468;
    14: op1_12_in12 = reg_0118;
    16: op1_12_in12 = reg_0443;
    17: op1_12_in12 = reg_0142;
    18: op1_12_in12 = imem07_in[127:124];
    19: op1_12_in12 = imem05_in[63:60];
    20: op1_12_in12 = reg_0454;
    84: op1_12_in12 = reg_0454;
    21: op1_12_in12 = reg_0572;
    22: op1_12_in12 = reg_0290;
    23: op1_12_in12 = reg_0548;
    24: op1_12_in12 = reg_0735;
    3: op1_12_in12 = reg_0169;
    25: op1_12_in12 = reg_0639;
    26: op1_12_in12 = reg_0715;
    27: op1_12_in12 = reg_0029;
    28: op1_12_in12 = imem04_in[43:40];
    29: op1_12_in12 = reg_0257;
    30: op1_12_in12 = reg_0466;
    34: op1_12_in12 = reg_0466;
    31: op1_12_in12 = imem02_in[15:12];
    32: op1_12_in12 = reg_0320;
    33: op1_12_in12 = reg_0622;
    35: op1_12_in12 = reg_0204;
    36: op1_12_in12 = reg_0518;
    37: op1_12_in12 = reg_0462;
    38: op1_12_in12 = reg_0789;
    39: op1_12_in12 = reg_0742;
    40: op1_12_in12 = imem06_in[55:52];
    41: op1_12_in12 = reg_0450;
    42: op1_12_in12 = reg_0349;
    43: op1_12_in12 = imem04_in[83:80];
    45: op1_12_in12 = reg_0456;
    46: op1_12_in12 = imem04_in[67:64];
    48: op1_12_in12 = reg_0207;
    49: op1_12_in12 = reg_0405;
    50: op1_12_in12 = imem06_in[35:32];
    86: op1_12_in12 = imem06_in[35:32];
    51: op1_12_in12 = imem04_in[75:72];
    52: op1_12_in12 = reg_0130;
    53: op1_12_in12 = reg_0494;
    55: op1_12_in12 = reg_0459;
    73: op1_12_in12 = reg_0459;
    56: op1_12_in12 = reg_0480;
    58: op1_12_in12 = imem01_in[55:52];
    59: op1_12_in12 = reg_0464;
    60: op1_12_in12 = reg_0647;
    61: op1_12_in12 = reg_0644;
    62: op1_12_in12 = reg_0162;
    63: op1_12_in12 = reg_0439;
    65: op1_12_in12 = reg_0453;
    67: op1_12_in12 = reg_0564;
    68: op1_12_in12 = reg_0499;
    69: op1_12_in12 = reg_0457;
    70: op1_12_in12 = reg_0600;
    71: op1_12_in12 = reg_0729;
    74: op1_12_in12 = reg_0703;
    75: op1_12_in12 = reg_0016;
    76: op1_12_in12 = reg_0628;
    77: op1_12_in12 = reg_0256;
    78: op1_12_in12 = reg_0714;
    79: op1_12_in12 = reg_0201;
    80: op1_12_in12 = imem02_in[103:100];
    81: op1_12_in12 = imem00_in[103:100];
    82: op1_12_in12 = reg_0409;
    83: op1_12_in12 = reg_0308;
    85: op1_12_in12 = reg_0507;
    87: op1_12_in12 = reg_0633;
    88: op1_12_in12 = reg_0824;
    89: op1_12_in12 = reg_0066;
    91: op1_12_in12 = reg_0342;
    92: op1_12_in12 = imem04_in[55:52];
    93: op1_12_in12 = imem04_in[51:48];
    94: op1_12_in12 = reg_0319;
    95: op1_12_in12 = reg_0544;
    default: op1_12_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_12_inv12 = 1;
    10: op1_12_inv12 = 1;
    11: op1_12_inv12 = 1;
    12: op1_12_inv12 = 1;
    15: op1_12_inv12 = 1;
    17: op1_12_inv12 = 1;
    18: op1_12_inv12 = 1;
    20: op1_12_inv12 = 1;
    21: op1_12_inv12 = 1;
    24: op1_12_inv12 = 1;
    25: op1_12_inv12 = 1;
    28: op1_12_inv12 = 1;
    29: op1_12_inv12 = 1;
    30: op1_12_inv12 = 1;
    31: op1_12_inv12 = 1;
    32: op1_12_inv12 = 1;
    33: op1_12_inv12 = 1;
    37: op1_12_inv12 = 1;
    38: op1_12_inv12 = 1;
    40: op1_12_inv12 = 1;
    45: op1_12_inv12 = 1;
    53: op1_12_inv12 = 1;
    56: op1_12_inv12 = 1;
    62: op1_12_inv12 = 1;
    67: op1_12_inv12 = 1;
    68: op1_12_inv12 = 1;
    69: op1_12_inv12 = 1;
    70: op1_12_inv12 = 1;
    72: op1_12_inv12 = 1;
    74: op1_12_inv12 = 1;
    78: op1_12_inv12 = 1;
    79: op1_12_inv12 = 1;
    80: op1_12_inv12 = 1;
    83: op1_12_inv12 = 1;
    84: op1_12_inv12 = 1;
    88: op1_12_inv12 = 1;
    89: op1_12_inv12 = 1;
    91: op1_12_inv12 = 1;
    92: op1_12_inv12 = 1;
    default: op1_12_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in13 = reg_0490;
    5: op1_12_in13 = reg_0312;
    6: op1_12_in13 = reg_0719;
    18: op1_12_in13 = reg_0719;
    7: op1_12_in13 = reg_0203;
    8: op1_12_in13 = reg_0275;
    95: op1_12_in13 = reg_0275;
    9: op1_12_in13 = reg_0352;
    10: op1_12_in13 = reg_0315;
    11: op1_12_in13 = reg_0109;
    12: op1_12_in13 = reg_0750;
    13: op1_12_in13 = reg_0452;
    14: op1_12_in13 = reg_0116;
    15: op1_12_in13 = reg_0781;
    16: op1_12_in13 = reg_0420;
    17: op1_12_in13 = reg_0139;
    19: op1_12_in13 = imem05_in[75:72];
    20: op1_12_in13 = reg_0477;
    41: op1_12_in13 = reg_0477;
    21: op1_12_in13 = reg_0587;
    22: op1_12_in13 = reg_0051;
    23: op1_12_in13 = reg_0259;
    24: op1_12_in13 = reg_0527;
    91: op1_12_in13 = reg_0527;
    3: op1_12_in13 = reg_0177;
    25: op1_12_in13 = reg_0644;
    26: op1_12_in13 = reg_0701;
    27: op1_12_in13 = imem07_in[3:0];
    28: op1_12_in13 = imem04_in[59:56];
    92: op1_12_in13 = imem04_in[59:56];
    29: op1_12_in13 = reg_0062;
    30: op1_12_in13 = reg_0462;
    34: op1_12_in13 = reg_0462;
    31: op1_12_in13 = imem02_in[55:52];
    32: op1_12_in13 = reg_0229;
    33: op1_12_in13 = reg_0405;
    35: op1_12_in13 = reg_0188;
    36: op1_12_in13 = reg_0092;
    37: op1_12_in13 = reg_0471;
    38: op1_12_in13 = reg_0493;
    39: op1_12_in13 = reg_0735;
    40: op1_12_in13 = imem06_in[87:84];
    42: op1_12_in13 = reg_0360;
    43: op1_12_in13 = imem04_in[87:84];
    45: op1_12_in13 = reg_0193;
    46: op1_12_in13 = reg_0544;
    48: op1_12_in13 = reg_0186;
    49: op1_12_in13 = reg_0404;
    50: op1_12_in13 = imem06_in[39:36];
    51: op1_12_in13 = imem04_in[111:108];
    52: op1_12_in13 = reg_0131;
    53: op1_12_in13 = reg_0786;
    55: op1_12_in13 = reg_0208;
    56: op1_12_in13 = reg_0189;
    58: op1_12_in13 = reg_0496;
    59: op1_12_in13 = reg_0466;
    60: op1_12_in13 = reg_0355;
    61: op1_12_in13 = reg_0416;
    62: op1_12_in13 = reg_0169;
    63: op1_12_in13 = reg_0239;
    65: op1_12_in13 = reg_0455;
    67: op1_12_in13 = reg_0385;
    68: op1_12_in13 = reg_0732;
    69: op1_12_in13 = reg_0464;
    70: op1_12_in13 = reg_0595;
    71: op1_12_in13 = reg_0708;
    72: op1_12_in13 = reg_0211;
    73: op1_12_in13 = reg_0200;
    74: op1_12_in13 = reg_0607;
    75: op1_12_in13 = reg_0810;
    76: op1_12_in13 = reg_0242;
    77: op1_12_in13 = imem07_in[23:20];
    78: op1_12_in13 = imem07_in[43:40];
    79: op1_12_in13 = reg_0202;
    80: op1_12_in13 = reg_0142;
    81: op1_12_in13 = imem00_in[107:104];
    82: op1_12_in13 = reg_0354;
    83: op1_12_in13 = reg_0431;
    84: op1_12_in13 = reg_0457;
    85: op1_12_in13 = reg_0760;
    86: op1_12_in13 = imem06_in[71:68];
    87: op1_12_in13 = reg_0465;
    88: op1_12_in13 = reg_0029;
    89: op1_12_in13 = reg_0183;
    93: op1_12_in13 = imem04_in[103:100];
    94: op1_12_in13 = imem04_in[43:40];
    default: op1_12_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv13 = 1;
    6: op1_12_inv13 = 1;
    8: op1_12_inv13 = 1;
    10: op1_12_inv13 = 1;
    12: op1_12_inv13 = 1;
    14: op1_12_inv13 = 1;
    16: op1_12_inv13 = 1;
    17: op1_12_inv13 = 1;
    18: op1_12_inv13 = 1;
    22: op1_12_inv13 = 1;
    23: op1_12_inv13 = 1;
    24: op1_12_inv13 = 1;
    3: op1_12_inv13 = 1;
    25: op1_12_inv13 = 1;
    26: op1_12_inv13 = 1;
    29: op1_12_inv13 = 1;
    30: op1_12_inv13 = 1;
    33: op1_12_inv13 = 1;
    35: op1_12_inv13 = 1;
    39: op1_12_inv13 = 1;
    41: op1_12_inv13 = 1;
    42: op1_12_inv13 = 1;
    43: op1_12_inv13 = 1;
    46: op1_12_inv13 = 1;
    48: op1_12_inv13 = 1;
    50: op1_12_inv13 = 1;
    51: op1_12_inv13 = 1;
    52: op1_12_inv13 = 1;
    53: op1_12_inv13 = 1;
    56: op1_12_inv13 = 1;
    59: op1_12_inv13 = 1;
    67: op1_12_inv13 = 1;
    68: op1_12_inv13 = 1;
    72: op1_12_inv13 = 1;
    74: op1_12_inv13 = 1;
    78: op1_12_inv13 = 1;
    81: op1_12_inv13 = 1;
    82: op1_12_inv13 = 1;
    83: op1_12_inv13 = 1;
    84: op1_12_inv13 = 1;
    85: op1_12_inv13 = 1;
    88: op1_12_inv13 = 1;
    91: op1_12_inv13 = 1;
    93: op1_12_inv13 = 1;
    95: op1_12_inv13 = 1;
    default: op1_12_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in14 = reg_0491;
    5: op1_12_in14 = reg_0393;
    6: op1_12_in14 = reg_0707;
    71: op1_12_in14 = reg_0707;
    7: op1_12_in14 = reg_0190;
    8: op1_12_in14 = reg_0065;
    29: op1_12_in14 = reg_0065;
    9: op1_12_in14 = reg_0364;
    10: op1_12_in14 = reg_0813;
    11: op1_12_in14 = reg_0110;
    12: op1_12_in14 = reg_0752;
    13: op1_12_in14 = reg_0478;
    14: op1_12_in14 = reg_0119;
    15: op1_12_in14 = reg_0488;
    16: op1_12_in14 = reg_0448;
    17: op1_12_in14 = reg_0140;
    18: op1_12_in14 = reg_0717;
    19: op1_12_in14 = imem05_in[87:84];
    20: op1_12_in14 = reg_0469;
    21: op1_12_in14 = reg_0589;
    22: op1_12_in14 = reg_0258;
    23: op1_12_in14 = reg_0520;
    24: op1_12_in14 = reg_0085;
    3: op1_12_in14 = reg_0164;
    25: op1_12_in14 = imem02_in[47:44];
    26: op1_12_in14 = reg_0424;
    27: op1_12_in14 = imem07_in[23:20];
    28: op1_12_in14 = imem04_in[83:80];
    92: op1_12_in14 = imem04_in[83:80];
    30: op1_12_in14 = reg_0467;
    34: op1_12_in14 = reg_0467;
    31: op1_12_in14 = imem02_in[59:56];
    32: op1_12_in14 = reg_0354;
    33: op1_12_in14 = reg_0775;
    35: op1_12_in14 = reg_0201;
    36: op1_12_in14 = reg_0743;
    37: op1_12_in14 = reg_0187;
    56: op1_12_in14 = reg_0187;
    38: op1_12_in14 = reg_0784;
    39: op1_12_in14 = reg_0733;
    40: op1_12_in14 = imem06_in[103:100];
    41: op1_12_in14 = reg_0462;
    42: op1_12_in14 = reg_0346;
    43: op1_12_in14 = imem04_in[95:92];
    45: op1_12_in14 = reg_0207;
    46: op1_12_in14 = reg_0560;
    48: op1_12_in14 = reg_0758;
    49: op1_12_in14 = reg_0614;
    50: op1_12_in14 = imem06_in[67:64];
    51: op1_12_in14 = reg_0315;
    52: op1_12_in14 = imem06_in[3:0];
    53: op1_12_in14 = reg_0226;
    55: op1_12_in14 = reg_0191;
    58: op1_12_in14 = reg_0649;
    59: op1_12_in14 = reg_0473;
    60: op1_12_in14 = reg_0344;
    61: op1_12_in14 = imem05_in[47:44];
    62: op1_12_in14 = reg_0168;
    63: op1_12_in14 = reg_0267;
    65: op1_12_in14 = reg_0464;
    67: op1_12_in14 = reg_0569;
    68: op1_12_in14 = reg_0277;
    69: op1_12_in14 = reg_0477;
    84: op1_12_in14 = reg_0477;
    70: op1_12_in14 = reg_0331;
    72: op1_12_in14 = reg_0194;
    73: op1_12_in14 = reg_0208;
    74: op1_12_in14 = reg_0581;
    75: op1_12_in14 = imem04_in[35:32];
    76: op1_12_in14 = reg_0405;
    77: op1_12_in14 = imem07_in[27:24];
    78: op1_12_in14 = imem07_in[47:44];
    79: op1_12_in14 = reg_0206;
    80: op1_12_in14 = reg_0325;
    81: op1_12_in14 = imem00_in[111:108];
    82: op1_12_in14 = reg_0238;
    83: op1_12_in14 = reg_0679;
    85: op1_12_in14 = reg_0232;
    86: op1_12_in14 = reg_0299;
    87: op1_12_in14 = reg_0455;
    88: op1_12_in14 = reg_0816;
    89: op1_12_in14 = reg_0184;
    91: op1_12_in14 = reg_0095;
    93: op1_12_in14 = reg_0316;
    94: op1_12_in14 = imem04_in[111:108];
    95: op1_12_in14 = reg_0177;
    default: op1_12_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv14 = 1;
    5: op1_12_inv14 = 1;
    6: op1_12_inv14 = 1;
    8: op1_12_inv14 = 1;
    9: op1_12_inv14 = 1;
    10: op1_12_inv14 = 1;
    11: op1_12_inv14 = 1;
    12: op1_12_inv14 = 1;
    13: op1_12_inv14 = 1;
    15: op1_12_inv14 = 1;
    20: op1_12_inv14 = 1;
    23: op1_12_inv14 = 1;
    27: op1_12_inv14 = 1;
    32: op1_12_inv14 = 1;
    33: op1_12_inv14 = 1;
    34: op1_12_inv14 = 1;
    35: op1_12_inv14 = 1;
    39: op1_12_inv14 = 1;
    40: op1_12_inv14 = 1;
    41: op1_12_inv14 = 1;
    42: op1_12_inv14 = 1;
    43: op1_12_inv14 = 1;
    51: op1_12_inv14 = 1;
    53: op1_12_inv14 = 1;
    56: op1_12_inv14 = 1;
    58: op1_12_inv14 = 1;
    59: op1_12_inv14 = 1;
    60: op1_12_inv14 = 1;
    68: op1_12_inv14 = 1;
    69: op1_12_inv14 = 1;
    71: op1_12_inv14 = 1;
    74: op1_12_inv14 = 1;
    76: op1_12_inv14 = 1;
    77: op1_12_inv14 = 1;
    78: op1_12_inv14 = 1;
    81: op1_12_inv14 = 1;
    82: op1_12_inv14 = 1;
    84: op1_12_inv14 = 1;
    86: op1_12_inv14 = 1;
    92: op1_12_inv14 = 1;
    93: op1_12_inv14 = 1;
    default: op1_12_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in15 = reg_0492;
    5: op1_12_in15 = reg_0331;
    6: op1_12_in15 = reg_0430;
    7: op1_12_in15 = reg_0202;
    37: op1_12_in15 = reg_0202;
    8: op1_12_in15 = reg_0064;
    9: op1_12_in15 = reg_0341;
    10: op1_12_in15 = imem07_in[11:8];
    11: op1_12_in15 = imem02_in[19:16];
    12: op1_12_in15 = imem07_in[3:0];
    13: op1_12_in15 = reg_0193;
    14: op1_12_in15 = imem02_in[11:8];
    15: op1_12_in15 = reg_0795;
    16: op1_12_in15 = reg_0165;
    17: op1_12_in15 = imem06_in[15:12];
    18: op1_12_in15 = reg_0709;
    19: op1_12_in15 = imem05_in[107:104];
    61: op1_12_in15 = imem05_in[107:104];
    20: op1_12_in15 = reg_0460;
    21: op1_12_in15 = reg_0584;
    91: op1_12_in15 = reg_0584;
    22: op1_12_in15 = reg_0255;
    23: op1_12_in15 = reg_0559;
    24: op1_12_in15 = reg_0224;
    3: op1_12_in15 = reg_0185;
    25: op1_12_in15 = imem02_in[63:60];
    31: op1_12_in15 = imem02_in[63:60];
    26: op1_12_in15 = reg_0426;
    27: op1_12_in15 = imem07_in[39:36];
    28: op1_12_in15 = reg_0262;
    29: op1_12_in15 = reg_0067;
    30: op1_12_in15 = reg_0191;
    41: op1_12_in15 = reg_0191;
    32: op1_12_in15 = reg_0363;
    33: op1_12_in15 = reg_0773;
    34: op1_12_in15 = reg_0459;
    35: op1_12_in15 = reg_0212;
    36: op1_12_in15 = reg_0095;
    38: op1_12_in15 = reg_0736;
    39: op1_12_in15 = reg_0282;
    40: op1_12_in15 = reg_0624;
    42: op1_12_in15 = reg_0347;
    43: op1_12_in15 = reg_0059;
    45: op1_12_in15 = reg_0199;
    46: op1_12_in15 = reg_0555;
    48: op1_12_in15 = reg_0089;
    49: op1_12_in15 = reg_0812;
    50: op1_12_in15 = imem06_in[107:104];
    51: op1_12_in15 = reg_0560;
    52: op1_12_in15 = imem06_in[43:40];
    53: op1_12_in15 = reg_0258;
    55: op1_12_in15 = reg_0187;
    56: op1_12_in15 = reg_0207;
    58: op1_12_in15 = reg_0418;
    59: op1_12_in15 = reg_0474;
    60: op1_12_in15 = reg_0358;
    62: op1_12_in15 = reg_0171;
    63: op1_12_in15 = reg_0448;
    65: op1_12_in15 = reg_0469;
    84: op1_12_in15 = reg_0469;
    67: op1_12_in15 = reg_0001;
    68: op1_12_in15 = reg_0099;
    69: op1_12_in15 = reg_0473;
    70: op1_12_in15 = reg_0569;
    71: op1_12_in15 = reg_0727;
    72: op1_12_in15 = reg_0205;
    73: op1_12_in15 = imem01_in[35:32];
    74: op1_12_in15 = reg_0360;
    75: op1_12_in15 = imem04_in[87:84];
    76: op1_12_in15 = reg_0270;
    77: op1_12_in15 = imem07_in[31:28];
    78: op1_12_in15 = imem07_in[59:56];
    79: op1_12_in15 = reg_0192;
    80: op1_12_in15 = reg_0141;
    81: op1_12_in15 = reg_0695;
    82: op1_12_in15 = reg_0618;
    83: op1_12_in15 = reg_0223;
    85: op1_12_in15 = reg_0423;
    86: op1_12_in15 = reg_0577;
    87: op1_12_in15 = reg_0477;
    88: op1_12_in15 = reg_0794;
    92: op1_12_in15 = imem04_in[127:124];
    93: op1_12_in15 = reg_0553;
    94: op1_12_in15 = imem04_in[115:112];
    95: op1_12_in15 = reg_0542;
    default: op1_12_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv15 = 1;
    5: op1_12_inv15 = 1;
    7: op1_12_inv15 = 1;
    9: op1_12_inv15 = 1;
    11: op1_12_inv15 = 1;
    12: op1_12_inv15 = 1;
    14: op1_12_inv15 = 1;
    15: op1_12_inv15 = 1;
    16: op1_12_inv15 = 1;
    18: op1_12_inv15 = 1;
    19: op1_12_inv15 = 1;
    20: op1_12_inv15 = 1;
    21: op1_12_inv15 = 1;
    3: op1_12_inv15 = 1;
    26: op1_12_inv15 = 1;
    34: op1_12_inv15 = 1;
    36: op1_12_inv15 = 1;
    38: op1_12_inv15 = 1;
    41: op1_12_inv15 = 1;
    42: op1_12_inv15 = 1;
    45: op1_12_inv15 = 1;
    49: op1_12_inv15 = 1;
    50: op1_12_inv15 = 1;
    53: op1_12_inv15 = 1;
    55: op1_12_inv15 = 1;
    59: op1_12_inv15 = 1;
    62: op1_12_inv15 = 1;
    63: op1_12_inv15 = 1;
    65: op1_12_inv15 = 1;
    67: op1_12_inv15 = 1;
    69: op1_12_inv15 = 1;
    70: op1_12_inv15 = 1;
    73: op1_12_inv15 = 1;
    74: op1_12_inv15 = 1;
    79: op1_12_inv15 = 1;
    81: op1_12_inv15 = 1;
    83: op1_12_inv15 = 1;
    85: op1_12_inv15 = 1;
    86: op1_12_inv15 = 1;
    87: op1_12_inv15 = 1;
    88: op1_12_inv15 = 1;
    94: op1_12_inv15 = 1;
    default: op1_12_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in16 = reg_0493;
    5: op1_12_in16 = imem03_in[3:0];
    6: op1_12_in16 = reg_0442;
    7: op1_12_in16 = imem01_in[3:0];
    8: op1_12_in16 = reg_0050;
    9: op1_12_in16 = reg_0359;
    10: op1_12_in16 = imem07_in[39:36];
    11: op1_12_in16 = imem02_in[51:48];
    12: op1_12_in16 = imem07_in[23:20];
    13: op1_12_in16 = reg_0211;
    14: op1_12_in16 = imem02_in[39:36];
    15: op1_12_in16 = reg_0494;
    16: op1_12_in16 = reg_0166;
    17: op1_12_in16 = imem06_in[35:32];
    18: op1_12_in16 = reg_0713;
    19: op1_12_in16 = imem05_in[123:120];
    20: op1_12_in16 = reg_0479;
    21: op1_12_in16 = reg_0588;
    22: op1_12_in16 = reg_0068;
    23: op1_12_in16 = reg_0311;
    24: op1_12_in16 = reg_0260;
    39: op1_12_in16 = reg_0260;
    3: op1_12_in16 = reg_0168;
    25: op1_12_in16 = imem02_in[71:68];
    26: op1_12_in16 = reg_0446;
    27: op1_12_in16 = imem07_in[47:44];
    28: op1_12_in16 = reg_0545;
    29: op1_12_in16 = imem05_in[3:0];
    30: op1_12_in16 = reg_0188;
    31: op1_12_in16 = imem02_in[83:80];
    32: op1_12_in16 = reg_0530;
    33: op1_12_in16 = reg_0763;
    34: op1_12_in16 = reg_0452;
    35: op1_12_in16 = imem01_in[19:16];
    36: op1_12_in16 = reg_0097;
    37: op1_12_in16 = imem01_in[7:4];
    72: op1_12_in16 = imem01_in[7:4];
    79: op1_12_in16 = imem01_in[7:4];
    38: op1_12_in16 = reg_0271;
    40: op1_12_in16 = reg_0605;
    41: op1_12_in16 = reg_0210;
    42: op1_12_in16 = reg_0096;
    91: op1_12_in16 = reg_0096;
    43: op1_12_in16 = reg_0316;
    45: op1_12_in16 = imem01_in[63:60];
    46: op1_12_in16 = reg_0510;
    48: op1_12_in16 = reg_0246;
    49: op1_12_in16 = reg_0819;
    50: op1_12_in16 = imem06_in[111:108];
    51: op1_12_in16 = reg_0087;
    52: op1_12_in16 = imem06_in[59:56];
    53: op1_12_in16 = reg_0249;
    55: op1_12_in16 = reg_0209;
    56: op1_12_in16 = reg_0199;
    58: op1_12_in16 = reg_0504;
    59: op1_12_in16 = reg_0458;
    60: op1_12_in16 = reg_0362;
    61: op1_12_in16 = reg_0114;
    63: op1_12_in16 = reg_0175;
    65: op1_12_in16 = reg_0476;
    84: op1_12_in16 = reg_0476;
    67: op1_12_in16 = reg_0002;
    68: op1_12_in16 = reg_0309;
    69: op1_12_in16 = reg_0194;
    70: op1_12_in16 = reg_0387;
    71: op1_12_in16 = reg_0334;
    73: op1_12_in16 = imem01_in[51:48];
    74: op1_12_in16 = reg_0594;
    75: op1_12_in16 = imem04_in[91:88];
    76: op1_12_in16 = reg_0583;
    77: op1_12_in16 = imem07_in[71:68];
    78: op1_12_in16 = imem07_in[67:64];
    80: op1_12_in16 = reg_0703;
    81: op1_12_in16 = reg_0693;
    82: op1_12_in16 = reg_0035;
    83: op1_12_in16 = reg_0585;
    85: op1_12_in16 = reg_0567;
    86: op1_12_in16 = reg_0762;
    87: op1_12_in16 = reg_0473;
    88: op1_12_in16 = reg_0319;
    92: op1_12_in16 = reg_0247;
    93: op1_12_in16 = reg_0432;
    94: op1_12_in16 = imem04_in[119:116];
    95: op1_12_in16 = reg_0537;
    default: op1_12_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv16 = 1;
    6: op1_12_inv16 = 1;
    7: op1_12_inv16 = 1;
    8: op1_12_inv16 = 1;
    10: op1_12_inv16 = 1;
    11: op1_12_inv16 = 1;
    13: op1_12_inv16 = 1;
    15: op1_12_inv16 = 1;
    17: op1_12_inv16 = 1;
    18: op1_12_inv16 = 1;
    21: op1_12_inv16 = 1;
    3: op1_12_inv16 = 1;
    25: op1_12_inv16 = 1;
    28: op1_12_inv16 = 1;
    29: op1_12_inv16 = 1;
    30: op1_12_inv16 = 1;
    32: op1_12_inv16 = 1;
    34: op1_12_inv16 = 1;
    35: op1_12_inv16 = 1;
    37: op1_12_inv16 = 1;
    38: op1_12_inv16 = 1;
    39: op1_12_inv16 = 1;
    40: op1_12_inv16 = 1;
    48: op1_12_inv16 = 1;
    49: op1_12_inv16 = 1;
    50: op1_12_inv16 = 1;
    52: op1_12_inv16 = 1;
    53: op1_12_inv16 = 1;
    56: op1_12_inv16 = 1;
    58: op1_12_inv16 = 1;
    59: op1_12_inv16 = 1;
    61: op1_12_inv16 = 1;
    65: op1_12_inv16 = 1;
    68: op1_12_inv16 = 1;
    70: op1_12_inv16 = 1;
    71: op1_12_inv16 = 1;
    72: op1_12_inv16 = 1;
    73: op1_12_inv16 = 1;
    75: op1_12_inv16 = 1;
    76: op1_12_inv16 = 1;
    78: op1_12_inv16 = 1;
    81: op1_12_inv16 = 1;
    82: op1_12_inv16 = 1;
    83: op1_12_inv16 = 1;
    84: op1_12_inv16 = 1;
    86: op1_12_inv16 = 1;
    91: op1_12_inv16 = 1;
    92: op1_12_inv16 = 1;
    default: op1_12_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in17 = reg_0494;
    5: op1_12_in17 = imem03_in[23:20];
    6: op1_12_in17 = reg_0172;
    63: op1_12_in17 = reg_0172;
    7: op1_12_in17 = imem01_in[27:24];
    37: op1_12_in17 = imem01_in[27:24];
    8: op1_12_in17 = imem05_in[47:44];
    9: op1_12_in17 = reg_0330;
    10: op1_12_in17 = imem07_in[55:52];
    11: op1_12_in17 = imem02_in[59:56];
    12: op1_12_in17 = imem07_in[35:32];
    13: op1_12_in17 = reg_0205;
    14: op1_12_in17 = imem02_in[47:44];
    15: op1_12_in17 = reg_0780;
    16: op1_12_in17 = reg_0164;
    17: op1_12_in17 = imem06_in[39:36];
    18: op1_12_in17 = reg_0429;
    19: op1_12_in17 = reg_0143;
    20: op1_12_in17 = reg_0459;
    21: op1_12_in17 = reg_0576;
    22: op1_12_in17 = reg_0075;
    23: op1_12_in17 = imem04_in[11:8];
    24: op1_12_in17 = reg_0272;
    3: op1_12_in17 = reg_0178;
    25: op1_12_in17 = imem02_in[103:100];
    26: op1_12_in17 = reg_0438;
    27: op1_12_in17 = imem07_in[59:56];
    28: op1_12_in17 = reg_0544;
    29: op1_12_in17 = imem05_in[35:32];
    30: op1_12_in17 = reg_0186;
    31: op1_12_in17 = imem02_in[111:108];
    32: op1_12_in17 = reg_0769;
    36: op1_12_in17 = reg_0769;
    33: op1_12_in17 = reg_0406;
    34: op1_12_in17 = reg_0210;
    35: op1_12_in17 = imem01_in[31:28];
    38: op1_12_in17 = reg_0304;
    39: op1_12_in17 = reg_0285;
    40: op1_12_in17 = reg_0020;
    41: op1_12_in17 = imem01_in[35:32];
    42: op1_12_in17 = reg_0535;
    43: op1_12_in17 = reg_0043;
    51: op1_12_in17 = reg_0043;
    45: op1_12_in17 = reg_0758;
    46: op1_12_in17 = reg_0516;
    48: op1_12_in17 = reg_0099;
    49: op1_12_in17 = reg_0238;
    50: op1_12_in17 = reg_0291;
    52: op1_12_in17 = imem06_in[83:80];
    53: op1_12_in17 = reg_0086;
    55: op1_12_in17 = reg_0188;
    56: op1_12_in17 = imem01_in[15:12];
    58: op1_12_in17 = reg_0670;
    59: op1_12_in17 = reg_0214;
    60: op1_12_in17 = reg_0359;
    61: op1_12_in17 = reg_0113;
    65: op1_12_in17 = reg_0470;
    67: op1_12_in17 = reg_0808;
    68: op1_12_in17 = reg_0245;
    69: op1_12_in17 = reg_0202;
    70: op1_12_in17 = reg_0623;
    71: op1_12_in17 = reg_0441;
    72: op1_12_in17 = imem01_in[23:20];
    73: op1_12_in17 = imem01_in[71:68];
    74: op1_12_in17 = reg_0590;
    75: op1_12_in17 = imem04_in[107:104];
    76: op1_12_in17 = reg_0638;
    77: op1_12_in17 = imem07_in[107:104];
    78: op1_12_in17 = imem07_in[71:68];
    79: op1_12_in17 = imem01_in[11:8];
    80: op1_12_in17 = reg_0587;
    81: op1_12_in17 = reg_0681;
    82: op1_12_in17 = reg_0515;
    83: op1_12_in17 = reg_0065;
    84: op1_12_in17 = reg_0466;
    85: op1_12_in17 = reg_0290;
    86: op1_12_in17 = reg_0401;
    87: op1_12_in17 = reg_0200;
    88: op1_12_in17 = reg_0354;
    91: op1_12_in17 = reg_0487;
    92: op1_12_in17 = reg_0262;
    93: op1_12_in17 = reg_0076;
    94: op1_12_in17 = imem04_in[127:124];
    95: op1_12_in17 = reg_0060;
    default: op1_12_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv17 = 1;
    8: op1_12_inv17 = 1;
    10: op1_12_inv17 = 1;
    14: op1_12_inv17 = 1;
    17: op1_12_inv17 = 1;
    19: op1_12_inv17 = 1;
    24: op1_12_inv17 = 1;
    27: op1_12_inv17 = 1;
    28: op1_12_inv17 = 1;
    31: op1_12_inv17 = 1;
    32: op1_12_inv17 = 1;
    33: op1_12_inv17 = 1;
    35: op1_12_inv17 = 1;
    36: op1_12_inv17 = 1;
    39: op1_12_inv17 = 1;
    41: op1_12_inv17 = 1;
    46: op1_12_inv17 = 1;
    48: op1_12_inv17 = 1;
    49: op1_12_inv17 = 1;
    50: op1_12_inv17 = 1;
    52: op1_12_inv17 = 1;
    53: op1_12_inv17 = 1;
    60: op1_12_inv17 = 1;
    63: op1_12_inv17 = 1;
    67: op1_12_inv17 = 1;
    68: op1_12_inv17 = 1;
    69: op1_12_inv17 = 1;
    70: op1_12_inv17 = 1;
    71: op1_12_inv17 = 1;
    72: op1_12_inv17 = 1;
    73: op1_12_inv17 = 1;
    77: op1_12_inv17 = 1;
    78: op1_12_inv17 = 1;
    79: op1_12_inv17 = 1;
    81: op1_12_inv17 = 1;
    82: op1_12_inv17 = 1;
    84: op1_12_inv17 = 1;
    87: op1_12_inv17 = 1;
    91: op1_12_inv17 = 1;
    93: op1_12_inv17 = 1;
    94: op1_12_inv17 = 1;
    95: op1_12_inv17 = 1;
    default: op1_12_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in18 = reg_0495;
    5: op1_12_in18 = imem03_in[35:32];
    6: op1_12_in18 = reg_0161;
    7: op1_12_in18 = imem01_in[39:36];
    35: op1_12_in18 = imem01_in[39:36];
    41: op1_12_in18 = imem01_in[39:36];
    8: op1_12_in18 = imem05_in[75:72];
    9: op1_12_in18 = reg_0092;
    10: op1_12_in18 = imem07_in[63:60];
    11: op1_12_in18 = imem02_in[95:92];
    12: op1_12_in18 = imem07_in[39:36];
    13: op1_12_in18 = reg_0199;
    14: op1_12_in18 = imem02_in[51:48];
    15: op1_12_in18 = reg_0782;
    16: op1_12_in18 = reg_0176;
    17: op1_12_in18 = imem06_in[99:96];
    18: op1_12_in18 = reg_0436;
    19: op1_12_in18 = reg_0153;
    20: op1_12_in18 = reg_0214;
    21: op1_12_in18 = reg_0360;
    22: op1_12_in18 = reg_0072;
    23: op1_12_in18 = imem04_in[47:44];
    24: op1_12_in18 = reg_0086;
    25: op1_12_in18 = reg_0743;
    26: op1_12_in18 = reg_0431;
    27: op1_12_in18 = imem07_in[71:68];
    28: op1_12_in18 = reg_0328;
    29: op1_12_in18 = reg_0791;
    30: op1_12_in18 = reg_0196;
    31: op1_12_in18 = reg_0647;
    32: op1_12_in18 = reg_0539;
    33: op1_12_in18 = reg_0028;
    34: op1_12_in18 = reg_0211;
    36: op1_12_in18 = reg_0540;
    37: op1_12_in18 = imem01_in[119:116];
    38: op1_12_in18 = reg_0309;
    39: op1_12_in18 = reg_0135;
    40: op1_12_in18 = reg_0286;
    42: op1_12_in18 = reg_0531;
    43: op1_12_in18 = reg_0555;
    45: op1_12_in18 = reg_0514;
    74: op1_12_in18 = reg_0514;
    46: op1_12_in18 = reg_0280;
    48: op1_12_in18 = reg_0824;
    49: op1_12_in18 = imem07_in[87:84];
    50: op1_12_in18 = reg_0613;
    51: op1_12_in18 = reg_0088;
    52: op1_12_in18 = reg_0619;
    53: op1_12_in18 = reg_0152;
    55: op1_12_in18 = reg_0203;
    56: op1_12_in18 = imem01_in[35:32];
    58: op1_12_in18 = reg_0675;
    59: op1_12_in18 = reg_0201;
    60: op1_12_in18 = reg_0356;
    61: op1_12_in18 = reg_0278;
    63: op1_12_in18 = reg_0167;
    65: op1_12_in18 = reg_0458;
    67: op1_12_in18 = reg_0015;
    68: op1_12_in18 = reg_0103;
    69: op1_12_in18 = imem01_in[11:8];
    70: op1_12_in18 = reg_0649;
    71: op1_12_in18 = reg_0439;
    72: op1_12_in18 = imem01_in[51:48];
    73: op1_12_in18 = imem01_in[75:72];
    75: op1_12_in18 = imem04_in[127:124];
    76: op1_12_in18 = reg_0576;
    77: op1_12_in18 = reg_0389;
    78: op1_12_in18 = imem07_in[83:80];
    79: op1_12_in18 = imem01_in[47:44];
    80: op1_12_in18 = reg_0345;
    81: op1_12_in18 = reg_0685;
    82: op1_12_in18 = reg_0039;
    83: op1_12_in18 = reg_0780;
    84: op1_12_in18 = reg_0205;
    85: op1_12_in18 = reg_0073;
    86: op1_12_in18 = reg_0032;
    87: op1_12_in18 = reg_0189;
    88: op1_12_in18 = reg_0618;
    91: op1_12_in18 = reg_0117;
    92: op1_12_in18 = reg_0058;
    93: op1_12_in18 = reg_0529;
    94: op1_12_in18 = reg_0275;
    95: op1_12_in18 = reg_0551;
    default: op1_12_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv18 = 1;
    10: op1_12_inv18 = 1;
    11: op1_12_inv18 = 1;
    12: op1_12_inv18 = 1;
    13: op1_12_inv18 = 1;
    16: op1_12_inv18 = 1;
    17: op1_12_inv18 = 1;
    21: op1_12_inv18 = 1;
    22: op1_12_inv18 = 1;
    23: op1_12_inv18 = 1;
    24: op1_12_inv18 = 1;
    28: op1_12_inv18 = 1;
    32: op1_12_inv18 = 1;
    33: op1_12_inv18 = 1;
    34: op1_12_inv18 = 1;
    35: op1_12_inv18 = 1;
    36: op1_12_inv18 = 1;
    37: op1_12_inv18 = 1;
    38: op1_12_inv18 = 1;
    40: op1_12_inv18 = 1;
    42: op1_12_inv18 = 1;
    46: op1_12_inv18 = 1;
    48: op1_12_inv18 = 1;
    49: op1_12_inv18 = 1;
    50: op1_12_inv18 = 1;
    52: op1_12_inv18 = 1;
    53: op1_12_inv18 = 1;
    59: op1_12_inv18 = 1;
    61: op1_12_inv18 = 1;
    63: op1_12_inv18 = 1;
    67: op1_12_inv18 = 1;
    68: op1_12_inv18 = 1;
    69: op1_12_inv18 = 1;
    71: op1_12_inv18 = 1;
    72: op1_12_inv18 = 1;
    73: op1_12_inv18 = 1;
    74: op1_12_inv18 = 1;
    75: op1_12_inv18 = 1;
    76: op1_12_inv18 = 1;
    77: op1_12_inv18 = 1;
    78: op1_12_inv18 = 1;
    79: op1_12_inv18 = 1;
    80: op1_12_inv18 = 1;
    82: op1_12_inv18 = 1;
    87: op1_12_inv18 = 1;
    92: op1_12_inv18 = 1;
    default: op1_12_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in19 = reg_0262;
    5: op1_12_in19 = imem04_in[7:4];
    6: op1_12_in19 = reg_0163;
    7: op1_12_in19 = imem01_in[83:80];
    8: op1_12_in19 = imem05_in[127:124];
    9: op1_12_in19 = reg_0088;
    10: op1_12_in19 = imem07_in[103:100];
    11: op1_12_in19 = imem02_in[123:120];
    12: op1_12_in19 = imem07_in[75:72];
    13: op1_12_in19 = imem01_in[27:24];
    14: op1_12_in19 = reg_0642;
    15: op1_12_in19 = reg_0786;
    17: op1_12_in19 = reg_0611;
    18: op1_12_in19 = reg_0447;
    19: op1_12_in19 = reg_0155;
    20: op1_12_in19 = reg_0210;
    21: op1_12_in19 = reg_0343;
    22: op1_12_in19 = imem05_in[71:68];
    23: op1_12_in19 = imem04_in[55:52];
    24: op1_12_in19 = reg_0147;
    25: op1_12_in19 = reg_0096;
    26: op1_12_in19 = reg_0179;
    27: op1_12_in19 = imem07_in[83:80];
    28: op1_12_in19 = reg_0087;
    29: op1_12_in19 = reg_0792;
    30: op1_12_in19 = reg_0205;
    31: op1_12_in19 = reg_0640;
    32: op1_12_in19 = reg_0526;
    33: op1_12_in19 = reg_0819;
    34: op1_12_in19 = reg_0201;
    35: op1_12_in19 = imem01_in[71:68];
    36: op1_12_in19 = reg_0535;
    92: op1_12_in19 = reg_0535;
    37: op1_12_in19 = reg_0337;
    38: op1_12_in19 = reg_0135;
    39: op1_12_in19 = reg_0133;
    40: op1_12_in19 = reg_0215;
    41: op1_12_in19 = imem01_in[103:100];
    72: op1_12_in19 = imem01_in[103:100];
    42: op1_12_in19 = imem03_in[79:76];
    43: op1_12_in19 = reg_0433;
    45: op1_12_in19 = reg_0515;
    46: op1_12_in19 = reg_0297;
    48: op1_12_in19 = reg_0245;
    49: op1_12_in19 = imem07_in[107:104];
    50: op1_12_in19 = reg_0286;
    51: op1_12_in19 = reg_0536;
    52: op1_12_in19 = reg_0633;
    53: op1_12_in19 = reg_0154;
    55: op1_12_in19 = reg_0196;
    56: op1_12_in19 = imem01_in[55:52];
    58: op1_12_in19 = reg_0676;
    59: op1_12_in19 = reg_0190;
    60: op1_12_in19 = reg_0406;
    61: op1_12_in19 = reg_0277;
    63: op1_12_in19 = reg_0182;
    65: op1_12_in19 = reg_0207;
    67: op1_12_in19 = reg_0806;
    68: op1_12_in19 = reg_0236;
    69: op1_12_in19 = imem01_in[23:20];
    70: op1_12_in19 = reg_0012;
    71: op1_12_in19 = reg_0442;
    73: op1_12_in19 = reg_0497;
    74: op1_12_in19 = reg_0323;
    75: op1_12_in19 = reg_0545;
    76: op1_12_in19 = reg_0512;
    77: op1_12_in19 = reg_0393;
    78: op1_12_in19 = imem07_in[115:112];
    79: op1_12_in19 = reg_0336;
    80: op1_12_in19 = reg_0363;
    81: op1_12_in19 = reg_0492;
    82: op1_12_in19 = reg_0484;
    83: op1_12_in19 = reg_0311;
    84: op1_12_in19 = reg_0195;
    85: op1_12_in19 = reg_0108;
    86: op1_12_in19 = reg_0593;
    87: op1_12_in19 = reg_0187;
    88: op1_12_in19 = reg_0408;
    91: op1_12_in19 = reg_0055;
    93: op1_12_in19 = reg_0431;
    94: op1_12_in19 = reg_0534;
    95: op1_12_in19 = reg_0516;
    default: op1_12_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_12_inv19 = 1;
    10: op1_12_inv19 = 1;
    11: op1_12_inv19 = 1;
    12: op1_12_inv19 = 1;
    13: op1_12_inv19 = 1;
    17: op1_12_inv19 = 1;
    18: op1_12_inv19 = 1;
    19: op1_12_inv19 = 1;
    20: op1_12_inv19 = 1;
    21: op1_12_inv19 = 1;
    23: op1_12_inv19 = 1;
    24: op1_12_inv19 = 1;
    25: op1_12_inv19 = 1;
    28: op1_12_inv19 = 1;
    30: op1_12_inv19 = 1;
    32: op1_12_inv19 = 1;
    33: op1_12_inv19 = 1;
    36: op1_12_inv19 = 1;
    37: op1_12_inv19 = 1;
    39: op1_12_inv19 = 1;
    41: op1_12_inv19 = 1;
    42: op1_12_inv19 = 1;
    46: op1_12_inv19 = 1;
    53: op1_12_inv19 = 1;
    55: op1_12_inv19 = 1;
    59: op1_12_inv19 = 1;
    60: op1_12_inv19 = 1;
    65: op1_12_inv19 = 1;
    68: op1_12_inv19 = 1;
    71: op1_12_inv19 = 1;
    73: op1_12_inv19 = 1;
    75: op1_12_inv19 = 1;
    76: op1_12_inv19 = 1;
    77: op1_12_inv19 = 1;
    80: op1_12_inv19 = 1;
    81: op1_12_inv19 = 1;
    82: op1_12_inv19 = 1;
    83: op1_12_inv19 = 1;
    84: op1_12_inv19 = 1;
    86: op1_12_inv19 = 1;
    87: op1_12_inv19 = 1;
    88: op1_12_inv19 = 1;
    91: op1_12_inv19 = 1;
    94: op1_12_inv19 = 1;
    default: op1_12_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in20 = reg_0250;
    5: op1_12_in20 = imem04_in[11:8];
    6: op1_12_in20 = reg_0164;
    7: op1_12_in20 = imem01_in[91:88];
    8: op1_12_in20 = reg_0482;
    9: op1_12_in20 = reg_0095;
    10: op1_12_in20 = reg_0712;
    11: op1_12_in20 = reg_0666;
    14: op1_12_in20 = reg_0666;
    12: op1_12_in20 = imem07_in[91:88];
    13: op1_12_in20 = imem01_in[31:28];
    15: op1_12_in20 = reg_0486;
    17: op1_12_in20 = reg_0608;
    18: op1_12_in20 = reg_0444;
    19: op1_12_in20 = reg_0134;
    20: op1_12_in20 = reg_0207;
    21: op1_12_in20 = reg_0369;
    22: op1_12_in20 = imem05_in[107:104];
    23: op1_12_in20 = imem04_in[107:104];
    24: op1_12_in20 = reg_0135;
    25: op1_12_in20 = reg_0770;
    36: op1_12_in20 = reg_0770;
    26: op1_12_in20 = reg_0168;
    27: op1_12_in20 = imem07_in[119:116];
    28: op1_12_in20 = reg_0055;
    29: op1_12_in20 = reg_0798;
    30: op1_12_in20 = reg_0190;
    31: op1_12_in20 = reg_0349;
    32: op1_12_in20 = imem03_in[15:12];
    33: op1_12_in20 = reg_0779;
    34: op1_12_in20 = reg_0213;
    35: op1_12_in20 = imem01_in[83:80];
    37: op1_12_in20 = reg_0824;
    38: op1_12_in20 = reg_0133;
    39: op1_12_in20 = reg_0150;
    40: op1_12_in20 = reg_0278;
    52: op1_12_in20 = reg_0278;
    41: op1_12_in20 = imem01_in[107:104];
    42: op1_12_in20 = reg_0583;
    43: op1_12_in20 = reg_0631;
    45: op1_12_in20 = reg_0550;
    46: op1_12_in20 = reg_0508;
    48: op1_12_in20 = reg_0559;
    49: op1_12_in20 = reg_0720;
    50: op1_12_in20 = reg_0618;
    51: op1_12_in20 = reg_0551;
    53: op1_12_in20 = reg_0143;
    55: op1_12_in20 = reg_0205;
    56: op1_12_in20 = imem01_in[79:76];
    58: op1_12_in20 = imem02_in[119:116];
    59: op1_12_in20 = imem01_in[23:20];
    60: op1_12_in20 = reg_0518;
    61: op1_12_in20 = reg_0145;
    68: op1_12_in20 = reg_0145;
    63: op1_12_in20 = reg_0176;
    65: op1_12_in20 = imem01_in[3:0];
    67: op1_12_in20 = reg_0010;
    69: op1_12_in20 = imem01_in[43:40];
    70: op1_12_in20 = reg_0810;
    71: op1_12_in20 = reg_0180;
    72: op1_12_in20 = imem01_in[111:108];
    73: op1_12_in20 = reg_0820;
    74: op1_12_in20 = reg_0092;
    75: op1_12_in20 = reg_0553;
    76: op1_12_in20 = reg_0218;
    77: op1_12_in20 = reg_0253;
    78: op1_12_in20 = reg_0334;
    79: op1_12_in20 = reg_0225;
    80: op1_12_in20 = reg_0342;
    81: op1_12_in20 = reg_0612;
    82: op1_12_in20 = reg_0752;
    83: op1_12_in20 = reg_0776;
    84: op1_12_in20 = reg_0192;
    85: op1_12_in20 = reg_0106;
    86: op1_12_in20 = reg_0651;
    87: op1_12_in20 = reg_0201;
    88: op1_12_in20 = reg_0328;
    91: op1_12_in20 = imem03_in[7:4];
    92: op1_12_in20 = reg_0537;
    93: op1_12_in20 = reg_0301;
    94: op1_12_in20 = reg_0535;
    95: op1_12_in20 = reg_0556;
    default: op1_12_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv20 = 1;
    5: op1_12_inv20 = 1;
    6: op1_12_inv20 = 1;
    7: op1_12_inv20 = 1;
    10: op1_12_inv20 = 1;
    11: op1_12_inv20 = 1;
    17: op1_12_inv20 = 1;
    18: op1_12_inv20 = 1;
    24: op1_12_inv20 = 1;
    25: op1_12_inv20 = 1;
    30: op1_12_inv20 = 1;
    31: op1_12_inv20 = 1;
    32: op1_12_inv20 = 1;
    33: op1_12_inv20 = 1;
    35: op1_12_inv20 = 1;
    36: op1_12_inv20 = 1;
    37: op1_12_inv20 = 1;
    38: op1_12_inv20 = 1;
    41: op1_12_inv20 = 1;
    46: op1_12_inv20 = 1;
    48: op1_12_inv20 = 1;
    50: op1_12_inv20 = 1;
    51: op1_12_inv20 = 1;
    56: op1_12_inv20 = 1;
    58: op1_12_inv20 = 1;
    67: op1_12_inv20 = 1;
    70: op1_12_inv20 = 1;
    72: op1_12_inv20 = 1;
    75: op1_12_inv20 = 1;
    76: op1_12_inv20 = 1;
    77: op1_12_inv20 = 1;
    78: op1_12_inv20 = 1;
    83: op1_12_inv20 = 1;
    88: op1_12_inv20 = 1;
    93: op1_12_inv20 = 1;
    default: op1_12_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in21 = reg_0251;
    5: op1_12_in21 = imem04_in[15:12];
    7: op1_12_in21 = reg_0500;
    8: op1_12_in21 = reg_0488;
    9: op1_12_in21 = reg_0052;
    10: op1_12_in21 = reg_0701;
    11: op1_12_in21 = reg_0637;
    12: op1_12_in21 = imem07_in[111:108];
    13: op1_12_in21 = imem01_in[43:40];
    14: op1_12_in21 = reg_0654;
    15: op1_12_in21 = reg_0262;
    17: op1_12_in21 = reg_0618;
    18: op1_12_in21 = reg_0435;
    19: op1_12_in21 = imem06_in[87:84];
    20: op1_12_in21 = reg_0211;
    21: op1_12_in21 = reg_0385;
    22: op1_12_in21 = imem05_in[111:108];
    23: op1_12_in21 = imem04_in[111:108];
    24: op1_12_in21 = reg_0128;
    25: op1_12_in21 = reg_0098;
    26: op1_12_in21 = reg_0157;
    27: op1_12_in21 = imem07_in[123:120];
    28: op1_12_in21 = reg_0556;
    29: op1_12_in21 = reg_0797;
    30: op1_12_in21 = reg_0197;
    31: op1_12_in21 = reg_0361;
    32: op1_12_in21 = imem03_in[87:84];
    33: op1_12_in21 = reg_0380;
    34: op1_12_in21 = reg_0212;
    35: op1_12_in21 = imem01_in[95:92];
    69: op1_12_in21 = imem01_in[95:92];
    36: op1_12_in21 = imem03_in[23:20];
    37: op1_12_in21 = reg_0759;
    38: op1_12_in21 = reg_0151;
    39: op1_12_in21 = reg_0153;
    53: op1_12_in21 = reg_0153;
    40: op1_12_in21 = reg_0408;
    41: op1_12_in21 = reg_0820;
    42: op1_12_in21 = reg_0565;
    43: op1_12_in21 = reg_0431;
    45: op1_12_in21 = reg_0760;
    46: op1_12_in21 = reg_0257;
    48: op1_12_in21 = imem01_in[47:44];
    49: op1_12_in21 = reg_0729;
    50: op1_12_in21 = reg_0402;
    51: op1_12_in21 = reg_0280;
    52: op1_12_in21 = reg_0612;
    55: op1_12_in21 = reg_0202;
    56: op1_12_in21 = imem01_in[119:116];
    58: op1_12_in21 = reg_0337;
    59: op1_12_in21 = imem01_in[35:32];
    60: op1_12_in21 = reg_0533;
    61: op1_12_in21 = reg_0136;
    63: op1_12_in21 = reg_0184;
    65: op1_12_in21 = imem01_in[23:20];
    67: op1_12_in21 = imem04_in[7:4];
    68: op1_12_in21 = reg_0134;
    70: op1_12_in21 = imem04_in[59:56];
    71: op1_12_in21 = reg_0172;
    72: op1_12_in21 = reg_0376;
    73: op1_12_in21 = reg_0130;
    74: op1_12_in21 = reg_0541;
    75: op1_12_in21 = reg_0537;
    76: op1_12_in21 = reg_0794;
    77: op1_12_in21 = reg_0239;
    78: op1_12_in21 = reg_0635;
    79: op1_12_in21 = reg_0423;
    80: op1_12_in21 = reg_0527;
    81: op1_12_in21 = reg_0698;
    82: op1_12_in21 = imem07_in[3:0];
    83: op1_12_in21 = reg_0416;
    84: op1_12_in21 = imem01_in[19:16];
    85: op1_12_in21 = reg_0669;
    86: op1_12_in21 = reg_0652;
    87: op1_12_in21 = reg_0213;
    88: op1_12_in21 = imem06_in[35:32];
    91: op1_12_in21 = reg_0528;
    92: op1_12_in21 = reg_0555;
    93: op1_12_in21 = reg_0643;
    94: op1_12_in21 = reg_0548;
    95: op1_12_in21 = reg_0308;
    default: op1_12_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv21 = 1;
    5: op1_12_inv21 = 1;
    7: op1_12_inv21 = 1;
    11: op1_12_inv21 = 1;
    13: op1_12_inv21 = 1;
    14: op1_12_inv21 = 1;
    18: op1_12_inv21 = 1;
    20: op1_12_inv21 = 1;
    21: op1_12_inv21 = 1;
    24: op1_12_inv21 = 1;
    25: op1_12_inv21 = 1;
    26: op1_12_inv21 = 1;
    29: op1_12_inv21 = 1;
    33: op1_12_inv21 = 1;
    34: op1_12_inv21 = 1;
    35: op1_12_inv21 = 1;
    37: op1_12_inv21 = 1;
    38: op1_12_inv21 = 1;
    39: op1_12_inv21 = 1;
    41: op1_12_inv21 = 1;
    42: op1_12_inv21 = 1;
    45: op1_12_inv21 = 1;
    46: op1_12_inv21 = 1;
    48: op1_12_inv21 = 1;
    50: op1_12_inv21 = 1;
    53: op1_12_inv21 = 1;
    60: op1_12_inv21 = 1;
    61: op1_12_inv21 = 1;
    63: op1_12_inv21 = 1;
    65: op1_12_inv21 = 1;
    67: op1_12_inv21 = 1;
    68: op1_12_inv21 = 1;
    69: op1_12_inv21 = 1;
    71: op1_12_inv21 = 1;
    73: op1_12_inv21 = 1;
    74: op1_12_inv21 = 1;
    75: op1_12_inv21 = 1;
    76: op1_12_inv21 = 1;
    77: op1_12_inv21 = 1;
    81: op1_12_inv21 = 1;
    83: op1_12_inv21 = 1;
    85: op1_12_inv21 = 1;
    94: op1_12_inv21 = 1;
    default: op1_12_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in22 = reg_0263;
    5: op1_12_in22 = imem04_in[43:40];
    7: op1_12_in22 = reg_0524;
    8: op1_12_in22 = reg_0484;
    9: op1_12_in22 = reg_0098;
    10: op1_12_in22 = reg_0424;
    11: op1_12_in22 = reg_0646;
    12: op1_12_in22 = reg_0722;
    13: op1_12_in22 = imem01_in[51:48];
    14: op1_12_in22 = reg_0358;
    15: op1_12_in22 = reg_0270;
    17: op1_12_in22 = reg_0623;
    18: op1_12_in22 = reg_0180;
    19: op1_12_in22 = reg_0614;
    20: op1_12_in22 = reg_0198;
    21: op1_12_in22 = reg_0398;
    22: op1_12_in22 = reg_0781;
    23: op1_12_in22 = imem04_in[115:112];
    24: op1_12_in22 = reg_0153;
    25: op1_12_in22 = reg_0498;
    26: op1_12_in22 = reg_0173;
    27: op1_12_in22 = reg_0716;
    28: op1_12_in22 = reg_0305;
    29: op1_12_in22 = reg_0488;
    30: op1_12_in22 = imem01_in[99:96];
    31: op1_12_in22 = reg_0365;
    32: op1_12_in22 = imem03_in[123:120];
    33: op1_12_in22 = imem07_in[3:0];
    34: op1_12_in22 = reg_0199;
    35: op1_12_in22 = imem01_in[123:120];
    36: op1_12_in22 = imem03_in[59:56];
    37: op1_12_in22 = reg_0333;
    38: op1_12_in22 = reg_0152;
    39: op1_12_in22 = reg_0137;
    40: op1_12_in22 = reg_0762;
    41: op1_12_in22 = reg_0334;
    42: op1_12_in22 = reg_0039;
    43: op1_12_in22 = reg_0050;
    45: op1_12_in22 = reg_0559;
    46: op1_12_in22 = reg_0066;
    48: op1_12_in22 = imem01_in[63:60];
    84: op1_12_in22 = imem01_in[63:60];
    49: op1_12_in22 = reg_0718;
    50: op1_12_in22 = reg_0318;
    51: op1_12_in22 = reg_0052;
    52: op1_12_in22 = reg_0407;
    53: op1_12_in22 = reg_0140;
    55: op1_12_in22 = reg_0206;
    56: op1_12_in22 = reg_0085;
    58: op1_12_in22 = reg_0417;
    59: op1_12_in22 = imem01_in[39:36];
    60: op1_12_in22 = reg_0082;
    61: op1_12_in22 = reg_0129;
    65: op1_12_in22 = imem01_in[35:32];
    67: op1_12_in22 = imem04_in[23:20];
    68: op1_12_in22 = imem06_in[15:12];
    69: op1_12_in22 = imem01_in[103:100];
    70: op1_12_in22 = imem04_in[95:92];
    71: op1_12_in22 = reg_0165;
    72: op1_12_in22 = reg_0668;
    73: op1_12_in22 = reg_0258;
    74: op1_12_in22 = reg_0314;
    75: op1_12_in22 = reg_0055;
    76: op1_12_in22 = reg_0501;
    77: op1_12_in22 = reg_0448;
    78: op1_12_in22 = reg_0449;
    79: op1_12_in22 = reg_0054;
    80: op1_12_in22 = reg_0539;
    81: op1_12_in22 = reg_0658;
    82: op1_12_in22 = imem07_in[23:20];
    83: op1_12_in22 = reg_0109;
    85: op1_12_in22 = reg_0601;
    86: op1_12_in22 = reg_0818;
    87: op1_12_in22 = reg_0192;
    88: op1_12_in22 = imem06_in[51:48];
    91: op1_12_in22 = reg_0010;
    92: op1_12_in22 = reg_0554;
    94: op1_12_in22 = reg_0554;
    93: op1_12_in22 = reg_0640;
    95: op1_12_in22 = reg_0079;
    default: op1_12_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv22 = 1;
    10: op1_12_inv22 = 1;
    13: op1_12_inv22 = 1;
    14: op1_12_inv22 = 1;
    15: op1_12_inv22 = 1;
    21: op1_12_inv22 = 1;
    23: op1_12_inv22 = 1;
    24: op1_12_inv22 = 1;
    25: op1_12_inv22 = 1;
    26: op1_12_inv22 = 1;
    28: op1_12_inv22 = 1;
    29: op1_12_inv22 = 1;
    30: op1_12_inv22 = 1;
    31: op1_12_inv22 = 1;
    33: op1_12_inv22 = 1;
    36: op1_12_inv22 = 1;
    39: op1_12_inv22 = 1;
    41: op1_12_inv22 = 1;
    42: op1_12_inv22 = 1;
    46: op1_12_inv22 = 1;
    48: op1_12_inv22 = 1;
    51: op1_12_inv22 = 1;
    52: op1_12_inv22 = 1;
    58: op1_12_inv22 = 1;
    59: op1_12_inv22 = 1;
    65: op1_12_inv22 = 1;
    68: op1_12_inv22 = 1;
    72: op1_12_inv22 = 1;
    73: op1_12_inv22 = 1;
    74: op1_12_inv22 = 1;
    77: op1_12_inv22 = 1;
    78: op1_12_inv22 = 1;
    79: op1_12_inv22 = 1;
    80: op1_12_inv22 = 1;
    81: op1_12_inv22 = 1;
    82: op1_12_inv22 = 1;
    86: op1_12_inv22 = 1;
    87: op1_12_inv22 = 1;
    92: op1_12_inv22 = 1;
    93: op1_12_inv22 = 1;
    95: op1_12_inv22 = 1;
    default: op1_12_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in23 = reg_0145;
    5: op1_12_in23 = imem04_in[55:52];
    7: op1_12_in23 = reg_0517;
    8: op1_12_in23 = reg_0793;
    9: op1_12_in23 = imem03_in[3:0];
    10: op1_12_in23 = reg_0432;
    92: op1_12_in23 = reg_0432;
    11: op1_12_in23 = reg_0664;
    12: op1_12_in23 = reg_0728;
    13: op1_12_in23 = imem01_in[63:60];
    14: op1_12_in23 = reg_0359;
    15: op1_12_in23 = reg_0230;
    17: op1_12_in23 = reg_0601;
    18: op1_12_in23 = reg_0172;
    19: op1_12_in23 = reg_0633;
    20: op1_12_in23 = imem01_in[23:20];
    34: op1_12_in23 = imem01_in[23:20];
    21: op1_12_in23 = reg_0396;
    22: op1_12_in23 = reg_0488;
    23: op1_12_in23 = imem04_in[127:124];
    24: op1_12_in23 = reg_0137;
    53: op1_12_in23 = reg_0137;
    25: op1_12_in23 = reg_0757;
    26: op1_12_in23 = reg_0184;
    27: op1_12_in23 = reg_0704;
    28: op1_12_in23 = reg_0534;
    29: op1_12_in23 = reg_0491;
    30: op1_12_in23 = reg_0758;
    31: op1_12_in23 = reg_0355;
    32: op1_12_in23 = imem03_in[127:124];
    33: op1_12_in23 = imem07_in[11:8];
    35: op1_12_in23 = reg_0520;
    72: op1_12_in23 = reg_0520;
    36: op1_12_in23 = imem03_in[87:84];
    37: op1_12_in23 = reg_0103;
    38: op1_12_in23 = reg_0134;
    39: op1_12_in23 = imem06_in[11:8];
    40: op1_12_in23 = reg_0821;
    41: op1_12_in23 = reg_0824;
    42: op1_12_in23 = reg_0584;
    43: op1_12_in23 = reg_0257;
    45: op1_12_in23 = reg_0502;
    46: op1_12_in23 = reg_0258;
    48: op1_12_in23 = imem01_in[71:68];
    49: op1_12_in23 = reg_0334;
    50: op1_12_in23 = reg_0317;
    51: op1_12_in23 = reg_0076;
    52: op1_12_in23 = reg_0763;
    55: op1_12_in23 = imem01_in[83:80];
    56: op1_12_in23 = reg_0496;
    58: op1_12_in23 = reg_0485;
    59: op1_12_in23 = imem01_in[51:48];
    60: op1_12_in23 = imem03_in[31:28];
    61: op1_12_in23 = imem06_in[31:28];
    65: op1_12_in23 = imem01_in[47:44];
    67: op1_12_in23 = imem04_in[59:56];
    68: op1_12_in23 = imem06_in[19:16];
    69: op1_12_in23 = imem01_in[107:104];
    70: op1_12_in23 = imem04_in[99:96];
    71: op1_12_in23 = reg_0169;
    73: op1_12_in23 = reg_0235;
    74: op1_12_in23 = reg_0080;
    75: op1_12_in23 = reg_0058;
    76: op1_12_in23 = reg_0767;
    86: op1_12_in23 = reg_0767;
    77: op1_12_in23 = reg_0175;
    78: op1_12_in23 = reg_0267;
    79: op1_12_in23 = reg_0216;
    80: op1_12_in23 = reg_0756;
    81: op1_12_in23 = reg_0255;
    82: op1_12_in23 = imem07_in[55:52];
    83: op1_12_in23 = imem05_in[31:28];
    84: op1_12_in23 = imem01_in[91:88];
    85: op1_12_in23 = reg_0671;
    87: op1_12_in23 = imem01_in[15:12];
    88: op1_12_in23 = imem06_in[55:52];
    91: op1_12_in23 = reg_0384;
    93: op1_12_in23 = reg_0296;
    94: op1_12_in23 = reg_0516;
    95: op1_12_in23 = reg_0052;
    default: op1_12_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv23 = 1;
    5: op1_12_inv23 = 1;
    8: op1_12_inv23 = 1;
    11: op1_12_inv23 = 1;
    12: op1_12_inv23 = 1;
    14: op1_12_inv23 = 1;
    15: op1_12_inv23 = 1;
    17: op1_12_inv23 = 1;
    19: op1_12_inv23 = 1;
    23: op1_12_inv23 = 1;
    24: op1_12_inv23 = 1;
    26: op1_12_inv23 = 1;
    30: op1_12_inv23 = 1;
    31: op1_12_inv23 = 1;
    32: op1_12_inv23 = 1;
    34: op1_12_inv23 = 1;
    35: op1_12_inv23 = 1;
    36: op1_12_inv23 = 1;
    37: op1_12_inv23 = 1;
    43: op1_12_inv23 = 1;
    46: op1_12_inv23 = 1;
    49: op1_12_inv23 = 1;
    50: op1_12_inv23 = 1;
    53: op1_12_inv23 = 1;
    55: op1_12_inv23 = 1;
    56: op1_12_inv23 = 1;
    59: op1_12_inv23 = 1;
    61: op1_12_inv23 = 1;
    65: op1_12_inv23 = 1;
    67: op1_12_inv23 = 1;
    68: op1_12_inv23 = 1;
    69: op1_12_inv23 = 1;
    73: op1_12_inv23 = 1;
    75: op1_12_inv23 = 1;
    76: op1_12_inv23 = 1;
    79: op1_12_inv23 = 1;
    85: op1_12_inv23 = 1;
    86: op1_12_inv23 = 1;
    87: op1_12_inv23 = 1;
    92: op1_12_inv23 = 1;
    94: op1_12_inv23 = 1;
    95: op1_12_inv23 = 1;
    default: op1_12_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in24 = reg_0133;
    5: op1_12_in24 = imem04_in[75:72];
    7: op1_12_in24 = reg_0508;
    8: op1_12_in24 = reg_0787;
    9: op1_12_in24 = imem03_in[7:4];
    10: op1_12_in24 = reg_0419;
    45: op1_12_in24 = reg_0419;
    11: op1_12_in24 = reg_0656;
    12: op1_12_in24 = reg_0719;
    27: op1_12_in24 = reg_0719;
    13: op1_12_in24 = imem01_in[87:84];
    59: op1_12_in24 = imem01_in[87:84];
    14: op1_12_in24 = reg_0363;
    15: op1_12_in24 = reg_0732;
    17: op1_12_in24 = reg_0381;
    18: op1_12_in24 = reg_0178;
    19: op1_12_in24 = reg_0348;
    20: op1_12_in24 = imem01_in[47:44];
    21: op1_12_in24 = reg_0389;
    22: op1_12_in24 = reg_0780;
    29: op1_12_in24 = reg_0780;
    23: op1_12_in24 = reg_0308;
    24: op1_12_in24 = reg_0144;
    25: op1_12_in24 = reg_0532;
    28: op1_12_in24 = reg_0297;
    30: op1_12_in24 = reg_0520;
    31: op1_12_in24 = reg_0323;
    32: op1_12_in24 = reg_0565;
    33: op1_12_in24 = imem07_in[71:68];
    34: op1_12_in24 = imem01_in[39:36];
    87: op1_12_in24 = imem01_in[39:36];
    35: op1_12_in24 = reg_0337;
    36: op1_12_in24 = imem03_in[119:116];
    37: op1_12_in24 = reg_0102;
    38: op1_12_in24 = reg_0610;
    39: op1_12_in24 = imem06_in[59:56];
    40: op1_12_in24 = reg_0748;
    41: op1_12_in24 = reg_0227;
    42: op1_12_in24 = reg_0755;
    43: op1_12_in24 = reg_0281;
    46: op1_12_in24 = reg_0070;
    48: op1_12_in24 = imem01_in[79:76];
    65: op1_12_in24 = imem01_in[79:76];
    49: op1_12_in24 = reg_0266;
    50: op1_12_in24 = reg_0369;
    51: op1_12_in24 = reg_0302;
    52: op1_12_in24 = reg_0038;
    53: op1_12_in24 = reg_0134;
    55: op1_12_in24 = imem01_in[107:104];
    56: op1_12_in24 = reg_0820;
    72: op1_12_in24 = reg_0820;
    58: op1_12_in24 = reg_0358;
    60: op1_12_in24 = imem03_in[67:64];
    61: op1_12_in24 = imem06_in[63:60];
    67: op1_12_in24 = imem04_in[111:108];
    68: op1_12_in24 = imem06_in[43:40];
    69: op1_12_in24 = imem01_in[127:124];
    70: op1_12_in24 = imem04_in[103:100];
    73: op1_12_in24 = reg_0241;
    74: op1_12_in24 = reg_0540;
    75: op1_12_in24 = reg_0547;
    76: op1_12_in24 = reg_0256;
    77: op1_12_in24 = reg_0166;
    78: op1_12_in24 = reg_0179;
    79: op1_12_in24 = reg_0425;
    80: op1_12_in24 = reg_0531;
    81: op1_12_in24 = reg_0692;
    82: op1_12_in24 = imem07_in[75:72];
    83: op1_12_in24 = imem05_in[55:52];
    84: op1_12_in24 = imem01_in[111:108];
    85: op1_12_in24 = reg_0678;
    86: op1_12_in24 = reg_0011;
    88: op1_12_in24 = imem06_in[87:84];
    91: op1_12_in24 = reg_0564;
    92: op1_12_in24 = reg_0280;
    93: op1_12_in24 = reg_0233;
    94: op1_12_in24 = reg_0249;
    95: op1_12_in24 = reg_0629;
    default: op1_12_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_12_inv24 = 1;
    10: op1_12_inv24 = 1;
    11: op1_12_inv24 = 1;
    12: op1_12_inv24 = 1;
    14: op1_12_inv24 = 1;
    15: op1_12_inv24 = 1;
    17: op1_12_inv24 = 1;
    23: op1_12_inv24 = 1;
    24: op1_12_inv24 = 1;
    28: op1_12_inv24 = 1;
    31: op1_12_inv24 = 1;
    33: op1_12_inv24 = 1;
    35: op1_12_inv24 = 1;
    40: op1_12_inv24 = 1;
    41: op1_12_inv24 = 1;
    42: op1_12_inv24 = 1;
    43: op1_12_inv24 = 1;
    45: op1_12_inv24 = 1;
    48: op1_12_inv24 = 1;
    51: op1_12_inv24 = 1;
    53: op1_12_inv24 = 1;
    59: op1_12_inv24 = 1;
    60: op1_12_inv24 = 1;
    61: op1_12_inv24 = 1;
    65: op1_12_inv24 = 1;
    68: op1_12_inv24 = 1;
    72: op1_12_inv24 = 1;
    76: op1_12_inv24 = 1;
    77: op1_12_inv24 = 1;
    79: op1_12_inv24 = 1;
    80: op1_12_inv24 = 1;
    84: op1_12_inv24 = 1;
    85: op1_12_inv24 = 1;
    87: op1_12_inv24 = 1;
    91: op1_12_inv24 = 1;
    94: op1_12_inv24 = 1;
    default: op1_12_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in25 = reg_0151;
    5: op1_12_in25 = imem04_in[107:104];
    7: op1_12_in25 = reg_0230;
    8: op1_12_in25 = reg_0256;
    9: op1_12_in25 = imem03_in[15:12];
    10: op1_12_in25 = reg_0434;
    11: op1_12_in25 = reg_0640;
    12: op1_12_in25 = reg_0730;
    13: op1_12_in25 = imem01_in[115:112];
    55: op1_12_in25 = imem01_in[115:112];
    14: op1_12_in25 = reg_0338;
    15: op1_12_in25 = reg_0744;
    17: op1_12_in25 = reg_0349;
    19: op1_12_in25 = reg_0379;
    20: op1_12_in25 = imem01_in[67:64];
    34: op1_12_in25 = imem01_in[67:64];
    21: op1_12_in25 = reg_0000;
    22: op1_12_in25 = reg_0794;
    23: op1_12_in25 = reg_0301;
    24: op1_12_in25 = reg_0607;
    25: op1_12_in25 = imem03_in[3:0];
    27: op1_12_in25 = reg_0723;
    28: op1_12_in25 = reg_0286;
    29: op1_12_in25 = reg_0785;
    30: op1_12_in25 = reg_0563;
    31: op1_12_in25 = reg_0518;
    32: op1_12_in25 = reg_0592;
    33: op1_12_in25 = imem07_in[83:80];
    35: op1_12_in25 = reg_0549;
    36: op1_12_in25 = reg_0599;
    37: op1_12_in25 = imem02_in[39:36];
    38: op1_12_in25 = reg_0629;
    39: op1_12_in25 = imem06_in[79:76];
    40: op1_12_in25 = reg_0406;
    41: op1_12_in25 = reg_0825;
    42: op1_12_in25 = reg_0571;
    43: op1_12_in25 = reg_0078;
    45: op1_12_in25 = reg_0420;
    46: op1_12_in25 = reg_0353;
    48: op1_12_in25 = imem01_in[95:92];
    49: op1_12_in25 = reg_0333;
    50: op1_12_in25 = reg_0748;
    51: op1_12_in25 = reg_0071;
    52: op1_12_in25 = reg_0753;
    53: op1_12_in25 = imem06_in[15:12];
    56: op1_12_in25 = reg_0761;
    58: op1_12_in25 = reg_0586;
    59: op1_12_in25 = imem01_in[99:96];
    60: op1_12_in25 = imem03_in[75:72];
    61: op1_12_in25 = imem06_in[99:96];
    65: op1_12_in25 = imem01_in[83:80];
    67: op1_12_in25 = reg_0537;
    68: op1_12_in25 = imem06_in[59:56];
    69: op1_12_in25 = reg_0376;
    70: op1_12_in25 = imem04_in[111:108];
    72: op1_12_in25 = reg_0397;
    73: op1_12_in25 = reg_0418;
    74: op1_12_in25 = reg_0526;
    75: op1_12_in25 = reg_0308;
    76: op1_12_in25 = imem07_in[11:8];
    78: op1_12_in25 = reg_0168;
    79: op1_12_in25 = reg_0505;
    80: op1_12_in25 = reg_0532;
    81: op1_12_in25 = reg_0699;
    82: op1_12_in25 = imem07_in[95:92];
    83: op1_12_in25 = imem05_in[63:60];
    84: op1_12_in25 = reg_0336;
    85: op1_12_in25 = imem02_in[7:4];
    86: op1_12_in25 = imem07_in[39:36];
    87: op1_12_in25 = imem01_in[43:40];
    88: op1_12_in25 = imem06_in[103:100];
    91: op1_12_in25 = reg_0490;
    92: op1_12_in25 = reg_0631;
    93: op1_12_in25 = imem05_in[3:0];
    94: op1_12_in25 = reg_0079;
    95: op1_12_in25 = reg_0617;
    default: op1_12_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv25 = 1;
    7: op1_12_inv25 = 1;
    8: op1_12_inv25 = 1;
    10: op1_12_inv25 = 1;
    11: op1_12_inv25 = 1;
    12: op1_12_inv25 = 1;
    14: op1_12_inv25 = 1;
    17: op1_12_inv25 = 1;
    24: op1_12_inv25 = 1;
    28: op1_12_inv25 = 1;
    30: op1_12_inv25 = 1;
    31: op1_12_inv25 = 1;
    35: op1_12_inv25 = 1;
    37: op1_12_inv25 = 1;
    39: op1_12_inv25 = 1;
    41: op1_12_inv25 = 1;
    45: op1_12_inv25 = 1;
    46: op1_12_inv25 = 1;
    49: op1_12_inv25 = 1;
    50: op1_12_inv25 = 1;
    51: op1_12_inv25 = 1;
    52: op1_12_inv25 = 1;
    53: op1_12_inv25 = 1;
    55: op1_12_inv25 = 1;
    56: op1_12_inv25 = 1;
    58: op1_12_inv25 = 1;
    59: op1_12_inv25 = 1;
    61: op1_12_inv25 = 1;
    70: op1_12_inv25 = 1;
    73: op1_12_inv25 = 1;
    74: op1_12_inv25 = 1;
    76: op1_12_inv25 = 1;
    84: op1_12_inv25 = 1;
    88: op1_12_inv25 = 1;
    91: op1_12_inv25 = 1;
    default: op1_12_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in26 = reg_0138;
    5: op1_12_in26 = reg_0548;
    7: op1_12_in26 = reg_0247;
    8: op1_12_in26 = reg_0241;
    9: op1_12_in26 = imem03_in[39:36];
    10: op1_12_in26 = reg_0446;
    11: op1_12_in26 = reg_0665;
    12: op1_12_in26 = reg_0434;
    13: op1_12_in26 = reg_0523;
    67: op1_12_in26 = reg_0523;
    14: op1_12_in26 = reg_0049;
    15: op1_12_in26 = reg_0132;
    17: op1_12_in26 = reg_0405;
    19: op1_12_in26 = reg_0351;
    20: op1_12_in26 = imem01_in[91:88];
    34: op1_12_in26 = imem01_in[91:88];
    21: op1_12_in26 = reg_0012;
    22: op1_12_in26 = reg_0276;
    23: op1_12_in26 = reg_0306;
    24: op1_12_in26 = reg_0613;
    25: op1_12_in26 = imem03_in[27:24];
    27: op1_12_in26 = reg_0726;
    28: op1_12_in26 = reg_0298;
    29: op1_12_in26 = reg_0794;
    30: op1_12_in26 = reg_0761;
    59: op1_12_in26 = reg_0761;
    31: op1_12_in26 = reg_0541;
    32: op1_12_in26 = reg_0584;
    33: op1_12_in26 = reg_0728;
    35: op1_12_in26 = reg_0333;
    41: op1_12_in26 = reg_0333;
    36: op1_12_in26 = reg_0596;
    37: op1_12_in26 = imem02_in[51:48];
    38: op1_12_in26 = reg_0219;
    39: op1_12_in26 = imem06_in[83:80];
    40: op1_12_in26 = reg_0620;
    42: op1_12_in26 = reg_0385;
    43: op1_12_in26 = imem05_in[3:0];
    46: op1_12_in26 = imem05_in[3:0];
    45: op1_12_in26 = reg_0124;
    48: op1_12_in26 = imem01_in[115:112];
    49: op1_12_in26 = reg_0084;
    50: op1_12_in26 = reg_0401;
    51: op1_12_in26 = reg_0508;
    52: op1_12_in26 = reg_0607;
    53: op1_12_in26 = imem06_in[47:44];
    55: op1_12_in26 = reg_0735;
    56: op1_12_in26 = reg_0737;
    72: op1_12_in26 = reg_0737;
    58: op1_12_in26 = reg_0590;
    60: op1_12_in26 = imem03_in[79:76];
    61: op1_12_in26 = imem06_in[119:116];
    65: op1_12_in26 = imem01_in[95:92];
    68: op1_12_in26 = imem06_in[127:124];
    69: op1_12_in26 = reg_0114;
    70: op1_12_in26 = imem04_in[123:120];
    73: op1_12_in26 = reg_0511;
    74: op1_12_in26 = reg_0093;
    75: op1_12_in26 = reg_0615;
    76: op1_12_in26 = imem07_in[39:36];
    78: op1_12_in26 = reg_0178;
    79: op1_12_in26 = reg_0122;
    80: op1_12_in26 = imem03_in[7:4];
    81: op1_12_in26 = reg_0453;
    82: op1_12_in26 = reg_0710;
    83: op1_12_in26 = imem05_in[75:72];
    84: op1_12_in26 = reg_0423;
    85: op1_12_in26 = imem02_in[23:20];
    86: op1_12_in26 = imem07_in[51:48];
    87: op1_12_in26 = imem01_in[79:76];
    88: op1_12_in26 = imem06_in[107:104];
    91: op1_12_in26 = reg_0387;
    92: op1_12_in26 = reg_0068;
    93: op1_12_in26 = imem05_in[11:8];
    94: op1_12_in26 = reg_0529;
    95: op1_12_in26 = reg_0779;
    default: op1_12_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_12_inv26 = 1;
    9: op1_12_inv26 = 1;
    10: op1_12_inv26 = 1;
    11: op1_12_inv26 = 1;
    15: op1_12_inv26 = 1;
    19: op1_12_inv26 = 1;
    24: op1_12_inv26 = 1;
    25: op1_12_inv26 = 1;
    33: op1_12_inv26 = 1;
    34: op1_12_inv26 = 1;
    35: op1_12_inv26 = 1;
    36: op1_12_inv26 = 1;
    40: op1_12_inv26 = 1;
    42: op1_12_inv26 = 1;
    45: op1_12_inv26 = 1;
    49: op1_12_inv26 = 1;
    50: op1_12_inv26 = 1;
    51: op1_12_inv26 = 1;
    52: op1_12_inv26 = 1;
    55: op1_12_inv26 = 1;
    56: op1_12_inv26 = 1;
    58: op1_12_inv26 = 1;
    61: op1_12_inv26 = 1;
    67: op1_12_inv26 = 1;
    68: op1_12_inv26 = 1;
    73: op1_12_inv26 = 1;
    75: op1_12_inv26 = 1;
    79: op1_12_inv26 = 1;
    83: op1_12_inv26 = 1;
    84: op1_12_inv26 = 1;
    85: op1_12_inv26 = 1;
    86: op1_12_inv26 = 1;
    87: op1_12_inv26 = 1;
    88: op1_12_inv26 = 1;
    91: op1_12_inv26 = 1;
    94: op1_12_inv26 = 1;
    default: op1_12_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in27 = imem06_in[11:8];
    5: op1_12_in27 = reg_0537;
    7: op1_12_in27 = reg_0122;
    8: op1_12_in27 = reg_0257;
    9: op1_12_in27 = imem03_in[79:76];
    10: op1_12_in27 = reg_0440;
    11: op1_12_in27 = reg_0667;
    12: op1_12_in27 = reg_0444;
    13: op1_12_in27 = reg_0820;
    14: op1_12_in27 = reg_0087;
    15: op1_12_in27 = reg_0145;
    17: op1_12_in27 = reg_0313;
    19: op1_12_in27 = reg_0313;
    20: op1_12_in27 = imem01_in[107:104];
    21: op1_12_in27 = reg_0003;
    22: op1_12_in27 = reg_0260;
    23: op1_12_in27 = reg_0265;
    24: op1_12_in27 = reg_0631;
    25: op1_12_in27 = imem03_in[43:40];
    27: op1_12_in27 = reg_0717;
    28: op1_12_in27 = reg_0051;
    29: op1_12_in27 = reg_0787;
    30: op1_12_in27 = reg_0507;
    31: op1_12_in27 = reg_0533;
    32: op1_12_in27 = reg_0751;
    33: op1_12_in27 = reg_0710;
    34: op1_12_in27 = reg_0497;
    55: op1_12_in27 = reg_0497;
    35: op1_12_in27 = reg_0235;
    41: op1_12_in27 = reg_0235;
    36: op1_12_in27 = reg_0585;
    37: op1_12_in27 = imem02_in[67:64];
    38: op1_12_in27 = reg_0626;
    39: op1_12_in27 = imem06_in[103:100];
    40: op1_12_in27 = reg_0815;
    42: op1_12_in27 = reg_0562;
    43: op1_12_in27 = imem05_in[35:32];
    45: op1_12_in27 = reg_0109;
    46: op1_12_in27 = imem05_in[71:68];
    48: op1_12_in27 = reg_0423;
    49: op1_12_in27 = reg_0267;
    50: op1_12_in27 = reg_0028;
    51: op1_12_in27 = reg_0065;
    95: op1_12_in27 = reg_0065;
    52: op1_12_in27 = reg_0620;
    53: op1_12_in27 = imem06_in[59:56];
    56: op1_12_in27 = reg_0418;
    58: op1_12_in27 = reg_0566;
    59: op1_12_in27 = reg_0649;
    60: op1_12_in27 = imem03_in[127:124];
    61: op1_12_in27 = imem06_in[123:120];
    65: op1_12_in27 = reg_0663;
    67: op1_12_in27 = reg_0556;
    68: op1_12_in27 = reg_0115;
    69: op1_12_in27 = reg_0131;
    70: op1_12_in27 = reg_0059;
    72: op1_12_in27 = reg_0422;
    73: op1_12_in27 = reg_0422;
    74: op1_12_in27 = imem03_in[75:72];
    75: op1_12_in27 = reg_0050;
    76: op1_12_in27 = imem07_in[59:56];
    78: op1_12_in27 = reg_0176;
    79: op1_12_in27 = reg_0672;
    80: op1_12_in27 = imem03_in[27:24];
    81: op1_12_in27 = reg_0464;
    82: op1_12_in27 = reg_0167;
    83: op1_12_in27 = imem05_in[91:88];
    84: op1_12_in27 = reg_0421;
    85: op1_12_in27 = imem02_in[27:24];
    86: op1_12_in27 = imem07_in[71:68];
    87: op1_12_in27 = imem01_in[87:84];
    88: op1_12_in27 = imem06_in[111:108];
    91: op1_12_in27 = reg_0001;
    92: op1_12_in27 = reg_0644;
    93: op1_12_in27 = imem05_in[31:28];
    94: op1_12_in27 = reg_0614;
    default: op1_12_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv27 = 1;
    12: op1_12_inv27 = 1;
    13: op1_12_inv27 = 1;
    14: op1_12_inv27 = 1;
    15: op1_12_inv27 = 1;
    17: op1_12_inv27 = 1;
    20: op1_12_inv27 = 1;
    21: op1_12_inv27 = 1;
    25: op1_12_inv27 = 1;
    30: op1_12_inv27 = 1;
    33: op1_12_inv27 = 1;
    34: op1_12_inv27 = 1;
    37: op1_12_inv27 = 1;
    42: op1_12_inv27 = 1;
    45: op1_12_inv27 = 1;
    46: op1_12_inv27 = 1;
    49: op1_12_inv27 = 1;
    51: op1_12_inv27 = 1;
    52: op1_12_inv27 = 1;
    53: op1_12_inv27 = 1;
    58: op1_12_inv27 = 1;
    59: op1_12_inv27 = 1;
    67: op1_12_inv27 = 1;
    68: op1_12_inv27 = 1;
    69: op1_12_inv27 = 1;
    72: op1_12_inv27 = 1;
    74: op1_12_inv27 = 1;
    75: op1_12_inv27 = 1;
    76: op1_12_inv27 = 1;
    79: op1_12_inv27 = 1;
    84: op1_12_inv27 = 1;
    85: op1_12_inv27 = 1;
    93: op1_12_inv27 = 1;
    default: op1_12_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in28 = imem06_in[19:16];
    5: op1_12_in28 = reg_0549;
    7: op1_12_in28 = reg_0103;
    8: op1_12_in28 = reg_0258;
    9: op1_12_in28 = reg_0582;
    10: op1_12_in28 = reg_0159;
    11: op1_12_in28 = reg_0341;
    12: op1_12_in28 = reg_0437;
    13: op1_12_in28 = reg_0825;
    14: op1_12_in28 = imem03_in[47:44];
    15: op1_12_in28 = reg_0152;
    17: op1_12_in28 = reg_0404;
    19: op1_12_in28 = reg_0404;
    20: op1_12_in28 = reg_0512;
    21: op1_12_in28 = reg_0804;
    22: op1_12_in28 = reg_0089;
    23: op1_12_in28 = reg_0253;
    24: op1_12_in28 = reg_0633;
    25: op1_12_in28 = reg_0602;
    27: op1_12_in28 = reg_0714;
    28: op1_12_in28 = reg_0278;
    29: op1_12_in28 = reg_0091;
    30: op1_12_in28 = reg_0505;
    31: op1_12_in28 = reg_0094;
    32: op1_12_in28 = reg_0395;
    33: op1_12_in28 = reg_0709;
    34: op1_12_in28 = reg_0824;
    35: op1_12_in28 = reg_0242;
    36: op1_12_in28 = reg_0600;
    37: op1_12_in28 = imem02_in[99:96];
    38: op1_12_in28 = reg_0615;
    39: op1_12_in28 = imem06_in[115:112];
    53: op1_12_in28 = imem06_in[115:112];
    40: op1_12_in28 = reg_0040;
    41: op1_12_in28 = reg_0306;
    56: op1_12_in28 = reg_0306;
    42: op1_12_in28 = reg_0811;
    43: op1_12_in28 = imem05_in[39:36];
    45: op1_12_in28 = imem02_in[63:60];
    46: op1_12_in28 = imem05_in[103:100];
    48: op1_12_in28 = reg_0421;
    49: op1_12_in28 = reg_0174;
    50: op1_12_in28 = reg_0368;
    51: op1_12_in28 = reg_0507;
    52: op1_12_in28 = reg_0236;
    55: op1_12_in28 = reg_0668;
    58: op1_12_in28 = reg_0518;
    59: op1_12_in28 = reg_0237;
    60: op1_12_in28 = reg_0347;
    61: op1_12_in28 = reg_0577;
    65: op1_12_in28 = reg_0100;
    67: op1_12_in28 = reg_0433;
    68: op1_12_in28 = reg_0291;
    69: op1_12_in28 = reg_0737;
    70: op1_12_in28 = reg_0087;
    72: op1_12_in28 = reg_0217;
    73: op1_12_in28 = reg_0506;
    74: op1_12_in28 = imem03_in[91:88];
    75: op1_12_in28 = reg_0617;
    76: op1_12_in28 = imem07_in[67:64];
    79: op1_12_in28 = reg_0676;
    80: op1_12_in28 = imem03_in[75:72];
    81: op1_12_in28 = reg_0469;
    82: op1_12_in28 = reg_0726;
    83: op1_12_in28 = imem05_in[95:92];
    93: op1_12_in28 = imem05_in[95:92];
    84: op1_12_in28 = reg_0511;
    85: op1_12_in28 = imem02_in[55:52];
    86: op1_12_in28 = imem07_in[87:84];
    87: op1_12_in28 = reg_0497;
    88: op1_12_in28 = imem07_in[27:24];
    91: op1_12_in28 = reg_0418;
    92: op1_12_in28 = imem05_in[63:60];
    94: op1_12_in28 = reg_0371;
    95: op1_12_in28 = reg_0598;
    default: op1_12_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_12_inv28 = 1;
    8: op1_12_inv28 = 1;
    13: op1_12_inv28 = 1;
    14: op1_12_inv28 = 1;
    15: op1_12_inv28 = 1;
    17: op1_12_inv28 = 1;
    19: op1_12_inv28 = 1;
    20: op1_12_inv28 = 1;
    23: op1_12_inv28 = 1;
    24: op1_12_inv28 = 1;
    25: op1_12_inv28 = 1;
    28: op1_12_inv28 = 1;
    31: op1_12_inv28 = 1;
    34: op1_12_inv28 = 1;
    35: op1_12_inv28 = 1;
    38: op1_12_inv28 = 1;
    39: op1_12_inv28 = 1;
    40: op1_12_inv28 = 1;
    41: op1_12_inv28 = 1;
    42: op1_12_inv28 = 1;
    45: op1_12_inv28 = 1;
    46: op1_12_inv28 = 1;
    49: op1_12_inv28 = 1;
    53: op1_12_inv28 = 1;
    55: op1_12_inv28 = 1;
    60: op1_12_inv28 = 1;
    61: op1_12_inv28 = 1;
    65: op1_12_inv28 = 1;
    68: op1_12_inv28 = 1;
    73: op1_12_inv28 = 1;
    74: op1_12_inv28 = 1;
    76: op1_12_inv28 = 1;
    79: op1_12_inv28 = 1;
    83: op1_12_inv28 = 1;
    85: op1_12_inv28 = 1;
    86: op1_12_inv28 = 1;
    87: op1_12_inv28 = 1;
    92: op1_12_inv28 = 1;
    94: op1_12_inv28 = 1;
    default: op1_12_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in29 = imem06_in[27:24];
    5: op1_12_in29 = reg_0554;
    7: op1_12_in29 = reg_0125;
    8: op1_12_in29 = reg_0253;
    9: op1_12_in29 = reg_0571;
    10: op1_12_in29 = reg_0169;
    11: op1_12_in29 = reg_0359;
    12: op1_12_in29 = reg_0420;
    13: op1_12_in29 = reg_0510;
    14: op1_12_in29 = imem03_in[79:76];
    15: op1_12_in29 = imem06_in[39:36];
    17: op1_12_in29 = reg_0406;
    19: op1_12_in29 = reg_0315;
    20: op1_12_in29 = reg_0227;
    21: op1_12_in29 = reg_0008;
    22: op1_12_in29 = reg_0148;
    23: op1_12_in29 = reg_0065;
    24: op1_12_in29 = reg_0632;
    25: op1_12_in29 = reg_0586;
    27: op1_12_in29 = reg_0702;
    28: op1_12_in29 = reg_0071;
    29: op1_12_in29 = reg_0741;
    30: op1_12_in29 = reg_0511;
    31: op1_12_in29 = imem03_in[3:0];
    32: op1_12_in29 = reg_0385;
    33: op1_12_in29 = reg_0711;
    34: op1_12_in29 = reg_0825;
    35: op1_12_in29 = reg_0245;
    36: op1_12_in29 = reg_0597;
    37: op1_12_in29 = imem02_in[103:100];
    38: op1_12_in29 = imem06_in[31:28];
    39: op1_12_in29 = imem06_in[119:116];
    40: op1_12_in29 = reg_0368;
    41: op1_12_in29 = reg_0054;
    42: op1_12_in29 = reg_0803;
    43: op1_12_in29 = imem05_in[123:120];
    45: op1_12_in29 = imem02_in[87:84];
    46: op1_12_in29 = reg_0791;
    48: op1_12_in29 = reg_0422;
    49: op1_12_in29 = reg_0167;
    50: op1_12_in29 = reg_0037;
    51: op1_12_in29 = reg_0068;
    52: op1_12_in29 = imem07_in[27:24];
    53: op1_12_in29 = reg_0299;
    55: op1_12_in29 = reg_0765;
    56: op1_12_in29 = reg_0217;
    69: op1_12_in29 = reg_0217;
    58: op1_12_in29 = reg_0541;
    59: op1_12_in29 = reg_0557;
    60: op1_12_in29 = reg_0559;
    61: op1_12_in29 = reg_0409;
    65: op1_12_in29 = reg_0734;
    67: op1_12_in29 = reg_0069;
    95: op1_12_in29 = reg_0069;
    68: op1_12_in29 = reg_0339;
    70: op1_12_in29 = reg_0523;
    72: op1_12_in29 = reg_0567;
    73: op1_12_in29 = reg_0243;
    74: op1_12_in29 = reg_0599;
    75: op1_12_in29 = reg_0614;
    76: op1_12_in29 = imem07_in[83:80];
    79: op1_12_in29 = imem02_in[47:44];
    80: op1_12_in29 = imem03_in[95:92];
    81: op1_12_in29 = reg_0481;
    82: op1_12_in29 = reg_0784;
    83: op1_12_in29 = reg_0641;
    84: op1_12_in29 = reg_0502;
    85: op1_12_in29 = imem02_in[67:64];
    86: op1_12_in29 = imem07_in[99:96];
    87: op1_12_in29 = reg_0225;
    88: op1_12_in29 = imem07_in[79:76];
    91: op1_12_in29 = reg_0807;
    92: op1_12_in29 = imem05_in[107:104];
    93: op1_12_in29 = imem05_in[119:116];
    94: op1_12_in29 = reg_0774;
    default: op1_12_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_12_inv29 = 1;
    5: op1_12_inv29 = 1;
    8: op1_12_inv29 = 1;
    9: op1_12_inv29 = 1;
    10: op1_12_inv29 = 1;
    13: op1_12_inv29 = 1;
    15: op1_12_inv29 = 1;
    17: op1_12_inv29 = 1;
    20: op1_12_inv29 = 1;
    21: op1_12_inv29 = 1;
    23: op1_12_inv29 = 1;
    24: op1_12_inv29 = 1;
    25: op1_12_inv29 = 1;
    30: op1_12_inv29 = 1;
    31: op1_12_inv29 = 1;
    33: op1_12_inv29 = 1;
    35: op1_12_inv29 = 1;
    36: op1_12_inv29 = 1;
    37: op1_12_inv29 = 1;
    38: op1_12_inv29 = 1;
    39: op1_12_inv29 = 1;
    41: op1_12_inv29 = 1;
    43: op1_12_inv29 = 1;
    46: op1_12_inv29 = 1;
    48: op1_12_inv29 = 1;
    49: op1_12_inv29 = 1;
    52: op1_12_inv29 = 1;
    55: op1_12_inv29 = 1;
    56: op1_12_inv29 = 1;
    60: op1_12_inv29 = 1;
    61: op1_12_inv29 = 1;
    65: op1_12_inv29 = 1;
    69: op1_12_inv29 = 1;
    73: op1_12_inv29 = 1;
    75: op1_12_inv29 = 1;
    76: op1_12_inv29 = 1;
    80: op1_12_inv29 = 1;
    81: op1_12_inv29 = 1;
    83: op1_12_inv29 = 1;
    84: op1_12_inv29 = 1;
    85: op1_12_inv29 = 1;
    86: op1_12_inv29 = 1;
    88: op1_12_inv29 = 1;
    92: op1_12_inv29 = 1;
    94: op1_12_inv29 = 1;
    default: op1_12_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_12_in30 = imem06_in[55:52];
    5: op1_12_in30 = reg_0540;
    7: op1_12_in30 = reg_0101;
    8: op1_12_in30 = reg_0136;
    9: op1_12_in30 = reg_0573;
    10: op1_12_in30 = reg_0185;
    11: op1_12_in30 = reg_0328;
    12: op1_12_in30 = imem07_in[23:20];
    13: op1_12_in30 = reg_0507;
    14: op1_12_in30 = imem03_in[127:124];
    15: op1_12_in30 = imem06_in[95:92];
    17: op1_12_in30 = reg_0028;
    19: op1_12_in30 = imem07_in[55:52];
    20: op1_12_in30 = reg_0499;
    21: op1_12_in30 = reg_0015;
    22: op1_12_in30 = reg_0133;
    23: op1_12_in30 = reg_0071;
    24: op1_12_in30 = reg_0622;
    25: op1_12_in30 = reg_0599;
    27: op1_12_in30 = reg_0729;
    28: op1_12_in30 = reg_0075;
    29: op1_12_in30 = reg_0304;
    30: op1_12_in30 = reg_0240;
    31: op1_12_in30 = imem03_in[23:20];
    32: op1_12_in30 = reg_0572;
    33: op1_12_in30 = reg_0706;
    34: op1_12_in30 = reg_0550;
    35: op1_12_in30 = reg_0238;
    36: op1_12_in30 = reg_0590;
    37: op1_12_in30 = imem02_in[107:104];
    38: op1_12_in30 = imem06_in[47:44];
    39: op1_12_in30 = imem06_in[123:120];
    40: op1_12_in30 = reg_0236;
    41: op1_12_in30 = reg_0216;
    42: op1_12_in30 = reg_0809;
    43: op1_12_in30 = reg_0791;
    45: op1_12_in30 = reg_0642;
    46: op1_12_in30 = reg_0788;
    48: op1_12_in30 = reg_0574;
    87: op1_12_in30 = reg_0574;
    50: op1_12_in30 = reg_0367;
    51: op1_12_in30 = reg_0069;
    52: op1_12_in30 = imem07_in[91:88];
    53: op1_12_in30 = reg_0291;
    55: op1_12_in30 = reg_0100;
    56: op1_12_in30 = reg_0567;
    58: op1_12_in30 = reg_0743;
    59: op1_12_in30 = reg_0321;
    60: op1_12_in30 = reg_0596;
    61: op1_12_in30 = reg_0298;
    65: op1_12_in30 = reg_0737;
    67: op1_12_in30 = reg_0233;
    94: op1_12_in30 = reg_0233;
    68: op1_12_in30 = reg_0630;
    69: op1_12_in30 = reg_0234;
    70: op1_12_in30 = reg_0558;
    72: op1_12_in30 = reg_0124;
    73: op1_12_in30 = reg_0125;
    74: op1_12_in30 = reg_0073;
    75: op1_12_in30 = reg_0585;
    76: op1_12_in30 = reg_0252;
    79: op1_12_in30 = imem02_in[111:108];
    80: op1_12_in30 = imem03_in[119:116];
    81: op1_12_in30 = reg_0474;
    82: op1_12_in30 = reg_0715;
    83: op1_12_in30 = reg_0027;
    84: op1_12_in30 = reg_0244;
    85: op1_12_in30 = imem02_in[91:88];
    86: op1_12_in30 = imem07_in[119:116];
    88: op1_12_in30 = imem07_in[107:104];
    91: op1_12_in30 = reg_0368;
    92: op1_12_in30 = reg_0792;
    93: op1_12_in30 = reg_0227;
    95: op1_12_in30 = reg_0774;
    default: op1_12_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    10: op1_12_inv30 = 1;
    13: op1_12_inv30 = 1;
    15: op1_12_inv30 = 1;
    19: op1_12_inv30 = 1;
    20: op1_12_inv30 = 1;
    24: op1_12_inv30 = 1;
    25: op1_12_inv30 = 1;
    27: op1_12_inv30 = 1;
    29: op1_12_inv30 = 1;
    30: op1_12_inv30 = 1;
    31: op1_12_inv30 = 1;
    32: op1_12_inv30 = 1;
    33: op1_12_inv30 = 1;
    35: op1_12_inv30 = 1;
    36: op1_12_inv30 = 1;
    37: op1_12_inv30 = 1;
    40: op1_12_inv30 = 1;
    43: op1_12_inv30 = 1;
    46: op1_12_inv30 = 1;
    51: op1_12_inv30 = 1;
    52: op1_12_inv30 = 1;
    53: op1_12_inv30 = 1;
    55: op1_12_inv30 = 1;
    56: op1_12_inv30 = 1;
    61: op1_12_inv30 = 1;
    65: op1_12_inv30 = 1;
    67: op1_12_inv30 = 1;
    68: op1_12_inv30 = 1;
    69: op1_12_inv30 = 1;
    72: op1_12_inv30 = 1;
    73: op1_12_inv30 = 1;
    74: op1_12_inv30 = 1;
    75: op1_12_inv30 = 1;
    76: op1_12_inv30 = 1;
    79: op1_12_inv30 = 1;
    82: op1_12_inv30 = 1;
    83: op1_12_inv30 = 1;
    84: op1_12_inv30 = 1;
    85: op1_12_inv30 = 1;
    87: op1_12_inv30 = 1;
    91: op1_12_inv30 = 1;
    default: op1_12_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_12_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_12_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in00 = imem06_in[59:56];
    5: op1_13_in00 = reg_0541;
    6: op1_13_in00 = imem00_in[15:12];
    7: op1_13_in00 = reg_0109;
    54: op1_13_in00 = reg_0109;
    67: op1_13_in00 = reg_0109;
    8: op1_13_in00 = reg_0146;
    92: op1_13_in00 = reg_0146;
    9: op1_13_in00 = reg_0572;
    10: op1_13_in00 = imem00_in[3:0];
    44: op1_13_in00 = imem00_in[3:0];
    11: op1_13_in00 = reg_0045;
    12: op1_13_in00 = imem00_in[47:44];
    27: op1_13_in00 = imem00_in[47:44];
    13: op1_13_in00 = reg_0821;
    14: op1_13_in00 = reg_0598;
    15: op1_13_in00 = imem06_in[103:100];
    16: op1_13_in00 = imem00_in[55:52];
    17: op1_13_in00 = reg_0747;
    18: op1_13_in00 = imem00_in[75:72];
    19: op1_13_in00 = imem07_in[83:80];
    20: op1_13_in00 = reg_0511;
    21: op1_13_in00 = reg_0270;
    22: op1_13_in00 = reg_0150;
    23: op1_13_in00 = imem05_in[39:36];
    24: op1_13_in00 = reg_0348;
    25: op1_13_in00 = reg_0579;
    3: op1_13_in00 = imem07_in[91:88];
    26: op1_13_in00 = imem00_in[23:20];
    49: op1_13_in00 = imem00_in[23:20];
    64: op1_13_in00 = imem00_in[23:20];
    89: op1_13_in00 = imem00_in[23:20];
    2: op1_13_in00 = imem07_in[19:16];
    28: op1_13_in00 = reg_0070;
    29: op1_13_in00 = reg_0309;
    30: op1_13_in00 = reg_0248;
    84: op1_13_in00 = reg_0248;
    31: op1_13_in00 = imem03_in[67:64];
    1: op1_13_in00 = imem07_in[43:40];
    32: op1_13_in00 = reg_0499;
    33: op1_13_in00 = imem00_in[63:60];
    34: op1_13_in00 = reg_0507;
    35: op1_13_in00 = reg_0219;
    36: op1_13_in00 = reg_0387;
    37: op1_13_in00 = reg_0661;
    38: op1_13_in00 = imem06_in[51:48];
    39: op1_13_in00 = reg_0289;
    40: op1_13_in00 = imem07_in[3:0];
    41: op1_13_in00 = reg_0234;
    42: op1_13_in00 = imem04_in[11:8];
    43: op1_13_in00 = reg_0491;
    45: op1_13_in00 = reg_0654;
    68: op1_13_in00 = reg_0654;
    46: op1_13_in00 = reg_0794;
    47: op1_13_in00 = imem00_in[59:56];
    48: op1_13_in00 = reg_0294;
    50: op1_13_in00 = imem07_in[7:4];
    51: op1_13_in00 = imem05_in[3:0];
    52: op1_13_in00 = imem07_in[99:96];
    53: op1_13_in00 = reg_0613;
    55: op1_13_in00 = reg_0825;
    56: op1_13_in00 = reg_0502;
    57: op1_13_in00 = imem00_in[7:4];
    66: op1_13_in00 = imem00_in[7:4];
    78: op1_13_in00 = imem00_in[7:4];
    58: op1_13_in00 = reg_0535;
    59: op1_13_in00 = reg_0423;
    60: op1_13_in00 = reg_0750;
    61: op1_13_in00 = reg_0606;
    62: op1_13_in00 = imem00_in[39:36];
    63: op1_13_in00 = imem00_in[27:24];
    65: op1_13_in00 = reg_0760;
    69: op1_13_in00 = reg_0506;
    70: op1_13_in00 = reg_0500;
    71: op1_13_in00 = imem00_in[19:16];
    72: op1_13_in00 = reg_0119;
    73: op1_13_in00 = reg_0660;
    74: op1_13_in00 = reg_0493;
    75: op1_13_in00 = reg_0065;
    76: op1_13_in00 = reg_0276;
    77: op1_13_in00 = imem00_in[35:32];
    79: op1_13_in00 = imem02_in[123:120];
    80: op1_13_in00 = reg_0329;
    81: op1_13_in00 = reg_0459;
    82: op1_13_in00 = reg_0158;
    83: op1_13_in00 = reg_0246;
    85: op1_13_in00 = imem02_in[107:104];
    86: op1_13_in00 = reg_0708;
    87: op1_13_in00 = reg_0220;
    88: op1_13_in00 = imem07_in[115:112];
    90: op1_13_in00 = reg_0696;
    91: op1_13_in00 = reg_0244;
    93: op1_13_in00 = reg_0128;
    94: op1_13_in00 = imem05_in[23:20];
    95: op1_13_in00 = reg_0640;
    default: op1_13_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv00 = 1;
    7: op1_13_inv00 = 1;
    8: op1_13_inv00 = 1;
    12: op1_13_inv00 = 1;
    13: op1_13_inv00 = 1;
    15: op1_13_inv00 = 1;
    16: op1_13_inv00 = 1;
    17: op1_13_inv00 = 1;
    20: op1_13_inv00 = 1;
    21: op1_13_inv00 = 1;
    24: op1_13_inv00 = 1;
    3: op1_13_inv00 = 1;
    28: op1_13_inv00 = 1;
    30: op1_13_inv00 = 1;
    31: op1_13_inv00 = 1;
    1: op1_13_inv00 = 1;
    32: op1_13_inv00 = 1;
    33: op1_13_inv00 = 1;
    34: op1_13_inv00 = 1;
    36: op1_13_inv00 = 1;
    38: op1_13_inv00 = 1;
    40: op1_13_inv00 = 1;
    42: op1_13_inv00 = 1;
    43: op1_13_inv00 = 1;
    44: op1_13_inv00 = 1;
    46: op1_13_inv00 = 1;
    48: op1_13_inv00 = 1;
    49: op1_13_inv00 = 1;
    50: op1_13_inv00 = 1;
    51: op1_13_inv00 = 1;
    52: op1_13_inv00 = 1;
    53: op1_13_inv00 = 1;
    55: op1_13_inv00 = 1;
    56: op1_13_inv00 = 1;
    60: op1_13_inv00 = 1;
    61: op1_13_inv00 = 1;
    62: op1_13_inv00 = 1;
    63: op1_13_inv00 = 1;
    64: op1_13_inv00 = 1;
    65: op1_13_inv00 = 1;
    66: op1_13_inv00 = 1;
    67: op1_13_inv00 = 1;
    71: op1_13_inv00 = 1;
    72: op1_13_inv00 = 1;
    74: op1_13_inv00 = 1;
    76: op1_13_inv00 = 1;
    77: op1_13_inv00 = 1;
    79: op1_13_inv00 = 1;
    80: op1_13_inv00 = 1;
    81: op1_13_inv00 = 1;
    84: op1_13_inv00 = 1;
    86: op1_13_inv00 = 1;
    88: op1_13_inv00 = 1;
    89: op1_13_inv00 = 1;
    90: op1_13_inv00 = 1;
    93: op1_13_inv00 = 1;
    95: op1_13_inv00 = 1;
    default: op1_13_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in01 = imem06_in[83:80];
    5: op1_13_in01 = reg_0281;
    6: op1_13_in01 = imem00_in[55:52];
    7: op1_13_in01 = reg_0107;
    8: op1_13_in01 = reg_0143;
    9: op1_13_in01 = reg_0395;
    10: op1_13_in01 = imem00_in[23:20];
    11: op1_13_in01 = reg_0089;
    12: op1_13_in01 = imem00_in[79:76];
    13: op1_13_in01 = reg_0511;
    14: op1_13_in01 = reg_0572;
    15: op1_13_in01 = reg_0620;
    16: op1_13_in01 = imem00_in[103:100];
    17: op1_13_in01 = reg_0005;
    18: op1_13_in01 = imem00_in[115:112];
    19: op1_13_in01 = reg_0726;
    20: op1_13_in01 = reg_0218;
    53: op1_13_in01 = reg_0218;
    21: op1_13_in01 = reg_0537;
    22: op1_13_in01 = reg_0152;
    23: op1_13_in01 = imem05_in[59:56];
    24: op1_13_in01 = reg_0372;
    25: op1_13_in01 = reg_0568;
    3: op1_13_in01 = imem07_in[111:108];
    26: op1_13_in01 = imem00_in[63:60];
    62: op1_13_in01 = imem00_in[63:60];
    27: op1_13_in01 = imem00_in[95:92];
    2: op1_13_in01 = imem07_in[23:20];
    28: op1_13_in01 = imem05_in[19:16];
    29: op1_13_in01 = reg_0744;
    30: op1_13_in01 = reg_0122;
    69: op1_13_in01 = reg_0122;
    31: op1_13_in01 = reg_0566;
    32: op1_13_in01 = reg_0807;
    33: op1_13_in01 = imem00_in[107:104];
    34: op1_13_in01 = reg_0232;
    65: op1_13_in01 = reg_0232;
    35: op1_13_in01 = reg_0123;
    36: op1_13_in01 = reg_0373;
    37: op1_13_in01 = reg_0651;
    38: op1_13_in01 = imem06_in[59:56];
    39: op1_13_in01 = reg_0605;
    40: op1_13_in01 = imem07_in[39:36];
    50: op1_13_in01 = imem07_in[39:36];
    41: op1_13_in01 = reg_0424;
    42: op1_13_in01 = imem04_in[39:36];
    91: op1_13_in01 = imem04_in[39:36];
    43: op1_13_in01 = reg_0793;
    44: op1_13_in01 = imem00_in[15:12];
    45: op1_13_in01 = reg_0661;
    46: op1_13_in01 = reg_0485;
    47: op1_13_in01 = reg_0685;
    48: op1_13_in01 = reg_0425;
    87: op1_13_in01 = reg_0425;
    49: op1_13_in01 = imem00_in[47:44];
    64: op1_13_in01 = imem00_in[47:44];
    51: op1_13_in01 = imem05_in[15:12];
    52: op1_13_in01 = imem07_in[127:124];
    88: op1_13_in01 = imem07_in[127:124];
    54: op1_13_in01 = reg_0687;
    55: op1_13_in01 = reg_0759;
    56: op1_13_in01 = reg_0248;
    57: op1_13_in01 = imem00_in[59:56];
    58: op1_13_in01 = reg_0098;
    59: op1_13_in01 = reg_0054;
    60: op1_13_in01 = reg_0329;
    61: op1_13_in01 = reg_0401;
    63: op1_13_in01 = imem00_in[39:36];
    66: op1_13_in01 = imem00_in[27:24];
    67: op1_13_in01 = reg_0070;
    68: op1_13_in01 = reg_0512;
    70: op1_13_in01 = reg_0432;
    71: op1_13_in01 = imem00_in[35:32];
    72: op1_13_in01 = reg_0677;
    73: op1_13_in01 = reg_0677;
    74: op1_13_in01 = reg_0596;
    75: op1_13_in01 = reg_0068;
    76: op1_13_in01 = reg_0279;
    77: op1_13_in01 = imem00_in[75:72];
    78: op1_13_in01 = imem00_in[11:8];
    79: op1_13_in01 = reg_0642;
    80: op1_13_in01 = reg_0399;
    81: op1_13_in01 = reg_0452;
    82: op1_13_in01 = reg_0157;
    83: op1_13_in01 = reg_0486;
    84: op1_13_in01 = reg_0504;
    85: op1_13_in01 = reg_0057;
    86: op1_13_in01 = reg_0103;
    89: op1_13_in01 = imem00_in[51:48];
    90: op1_13_in01 = reg_0684;
    92: op1_13_in01 = reg_0517;
    93: op1_13_in01 = reg_0138;
    94: op1_13_in01 = imem05_in[31:28];
    95: op1_13_in01 = imem05_in[3:0];
    default: op1_13_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv01 = 1;
    8: op1_13_inv01 = 1;
    10: op1_13_inv01 = 1;
    11: op1_13_inv01 = 1;
    15: op1_13_inv01 = 1;
    18: op1_13_inv01 = 1;
    20: op1_13_inv01 = 1;
    22: op1_13_inv01 = 1;
    24: op1_13_inv01 = 1;
    26: op1_13_inv01 = 1;
    27: op1_13_inv01 = 1;
    2: op1_13_inv01 = 1;
    28: op1_13_inv01 = 1;
    29: op1_13_inv01 = 1;
    30: op1_13_inv01 = 1;
    32: op1_13_inv01 = 1;
    33: op1_13_inv01 = 1;
    36: op1_13_inv01 = 1;
    38: op1_13_inv01 = 1;
    40: op1_13_inv01 = 1;
    41: op1_13_inv01 = 1;
    42: op1_13_inv01 = 1;
    46: op1_13_inv01 = 1;
    48: op1_13_inv01 = 1;
    49: op1_13_inv01 = 1;
    52: op1_13_inv01 = 1;
    53: op1_13_inv01 = 1;
    54: op1_13_inv01 = 1;
    58: op1_13_inv01 = 1;
    62: op1_13_inv01 = 1;
    66: op1_13_inv01 = 1;
    70: op1_13_inv01 = 1;
    73: op1_13_inv01 = 1;
    81: op1_13_inv01 = 1;
    82: op1_13_inv01 = 1;
    84: op1_13_inv01 = 1;
    85: op1_13_inv01 = 1;
    86: op1_13_inv01 = 1;
    88: op1_13_inv01 = 1;
    89: op1_13_inv01 = 1;
    90: op1_13_inv01 = 1;
    94: op1_13_inv01 = 1;
    95: op1_13_inv01 = 1;
    default: op1_13_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in02 = imem06_in[95:92];
    5: op1_13_in02 = reg_0294;
    6: op1_13_in02 = imem00_in[79:76];
    7: op1_13_in02 = reg_0126;
    8: op1_13_in02 = reg_0153;
    9: op1_13_in02 = reg_0387;
    60: op1_13_in02 = reg_0387;
    10: op1_13_in02 = imem00_in[35:32];
    11: op1_13_in02 = reg_0073;
    12: op1_13_in02 = imem00_in[83:80];
    77: op1_13_in02 = imem00_in[83:80];
    13: op1_13_in02 = reg_0239;
    14: op1_13_in02 = reg_0597;
    15: op1_13_in02 = reg_0621;
    16: op1_13_in02 = reg_0695;
    17: op1_13_in02 = reg_0751;
    18: op1_13_in02 = reg_0684;
    47: op1_13_in02 = reg_0684;
    19: op1_13_in02 = reg_0717;
    20: op1_13_in02 = reg_0506;
    21: op1_13_in02 = reg_0259;
    31: op1_13_in02 = reg_0259;
    22: op1_13_in02 = reg_0143;
    23: op1_13_in02 = imem05_in[63:60];
    24: op1_13_in02 = reg_0349;
    25: op1_13_in02 = reg_0578;
    3: op1_13_in02 = reg_0425;
    26: op1_13_in02 = imem00_in[71:68];
    49: op1_13_in02 = imem00_in[71:68];
    62: op1_13_in02 = imem00_in[71:68];
    27: op1_13_in02 = imem00_in[127:124];
    2: op1_13_in02 = imem07_in[59:56];
    28: op1_13_in02 = imem05_in[27:24];
    29: op1_13_in02 = reg_0148;
    30: op1_13_in02 = reg_0125;
    32: op1_13_in02 = reg_0800;
    33: op1_13_in02 = reg_0690;
    34: op1_13_in02 = reg_0246;
    35: op1_13_in02 = reg_0105;
    36: op1_13_in02 = reg_0747;
    37: op1_13_in02 = reg_0638;
    38: op1_13_in02 = imem06_in[91:88];
    39: op1_13_in02 = reg_0817;
    40: op1_13_in02 = imem07_in[87:84];
    41: op1_13_in02 = reg_0099;
    42: op1_13_in02 = imem04_in[55:52];
    43: op1_13_in02 = reg_0485;
    44: op1_13_in02 = reg_0672;
    45: op1_13_in02 = reg_0647;
    46: op1_13_in02 = reg_0309;
    48: op1_13_in02 = reg_0111;
    50: op1_13_in02 = imem07_in[67:64];
    51: op1_13_in02 = imem05_in[43:40];
    52: op1_13_in02 = reg_0727;
    53: op1_13_in02 = reg_0020;
    54: op1_13_in02 = imem00_in[15:12];
    78: op1_13_in02 = imem00_in[15:12];
    55: op1_13_in02 = reg_0237;
    56: op1_13_in02 = reg_0419;
    57: op1_13_in02 = imem00_in[67:64];
    71: op1_13_in02 = imem00_in[67:64];
    58: op1_13_in02 = reg_0757;
    59: op1_13_in02 = reg_0567;
    61: op1_13_in02 = reg_0405;
    63: op1_13_in02 = imem00_in[43:40];
    64: op1_13_in02 = reg_0492;
    65: op1_13_in02 = reg_0418;
    66: op1_13_in02 = imem00_in[59:56];
    67: op1_13_in02 = reg_0102;
    68: op1_13_in02 = reg_0534;
    69: op1_13_in02 = reg_0673;
    70: op1_13_in02 = reg_0077;
    72: op1_13_in02 = reg_0674;
    73: op1_13_in02 = reg_0674;
    74: op1_13_in02 = reg_0528;
    75: op1_13_in02 = reg_0513;
    76: op1_13_in02 = reg_0393;
    79: op1_13_in02 = reg_0254;
    80: op1_13_in02 = reg_0648;
    81: op1_13_in02 = reg_0208;
    82: op1_13_in02 = reg_0447;
    83: op1_13_in02 = reg_0278;
    84: op1_13_in02 = reg_0592;
    85: op1_13_in02 = reg_0533;
    86: op1_13_in02 = reg_0061;
    87: op1_13_in02 = reg_0234;
    88: op1_13_in02 = reg_0723;
    89: op1_13_in02 = imem00_in[91:88];
    90: op1_13_in02 = reg_0165;
    91: op1_13_in02 = imem04_in[67:64];
    92: op1_13_in02 = reg_0538;
    93: op1_13_in02 = reg_0285;
    94: op1_13_in02 = imem05_in[67:64];
    95: op1_13_in02 = imem05_in[71:68];
    default: op1_13_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv02 = 1;
    8: op1_13_inv02 = 1;
    10: op1_13_inv02 = 1;
    18: op1_13_inv02 = 1;
    19: op1_13_inv02 = 1;
    21: op1_13_inv02 = 1;
    23: op1_13_inv02 = 1;
    26: op1_13_inv02 = 1;
    27: op1_13_inv02 = 1;
    2: op1_13_inv02 = 1;
    28: op1_13_inv02 = 1;
    29: op1_13_inv02 = 1;
    30: op1_13_inv02 = 1;
    34: op1_13_inv02 = 1;
    35: op1_13_inv02 = 1;
    37: op1_13_inv02 = 1;
    39: op1_13_inv02 = 1;
    41: op1_13_inv02 = 1;
    43: op1_13_inv02 = 1;
    44: op1_13_inv02 = 1;
    45: op1_13_inv02 = 1;
    47: op1_13_inv02 = 1;
    48: op1_13_inv02 = 1;
    53: op1_13_inv02 = 1;
    54: op1_13_inv02 = 1;
    55: op1_13_inv02 = 1;
    58: op1_13_inv02 = 1;
    59: op1_13_inv02 = 1;
    60: op1_13_inv02 = 1;
    61: op1_13_inv02 = 1;
    63: op1_13_inv02 = 1;
    65: op1_13_inv02 = 1;
    66: op1_13_inv02 = 1;
    67: op1_13_inv02 = 1;
    68: op1_13_inv02 = 1;
    72: op1_13_inv02 = 1;
    75: op1_13_inv02 = 1;
    79: op1_13_inv02 = 1;
    82: op1_13_inv02 = 1;
    83: op1_13_inv02 = 1;
    86: op1_13_inv02 = 1;
    88: op1_13_inv02 = 1;
    91: op1_13_inv02 = 1;
    92: op1_13_inv02 = 1;
    94: op1_13_inv02 = 1;
    95: op1_13_inv02 = 1;
    default: op1_13_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in03 = imem06_in[111:108];
    5: op1_13_in03 = reg_0277;
    6: op1_13_in03 = reg_0670;
    7: op1_13_in03 = imem02_in[7:4];
    8: op1_13_in03 = reg_0141;
    9: op1_13_in03 = reg_0312;
    10: op1_13_in03 = imem00_in[47:44];
    11: op1_13_in03 = imem03_in[3:0];
    12: op1_13_in03 = imem00_in[95:92];
    13: op1_13_in03 = reg_0220;
    14: op1_13_in03 = reg_0360;
    15: op1_13_in03 = reg_0619;
    16: op1_13_in03 = reg_0696;
    17: op1_13_in03 = imem07_in[3:0];
    18: op1_13_in03 = reg_0679;
    19: op1_13_in03 = reg_0714;
    20: op1_13_in03 = reg_0234;
    21: op1_13_in03 = reg_0311;
    22: op1_13_in03 = imem06_in[7:4];
    23: op1_13_in03 = imem05_in[87:84];
    24: op1_13_in03 = reg_0383;
    25: op1_13_in03 = reg_0590;
    3: op1_13_in03 = reg_0424;
    26: op1_13_in03 = imem00_in[79:76];
    62: op1_13_in03 = imem00_in[79:76];
    66: op1_13_in03 = imem00_in[79:76];
    27: op1_13_in03 = reg_0693;
    2: op1_13_in03 = imem07_in[83:80];
    28: op1_13_in03 = imem05_in[75:72];
    29: op1_13_in03 = reg_0139;
    30: op1_13_in03 = reg_0112;
    31: op1_13_in03 = reg_0565;
    32: op1_13_in03 = reg_0014;
    33: op1_13_in03 = reg_0451;
    34: op1_13_in03 = reg_0217;
    35: op1_13_in03 = reg_0124;
    36: op1_13_in03 = reg_0012;
    37: op1_13_in03 = reg_0662;
    38: op1_13_in03 = imem06_in[99:96];
    39: op1_13_in03 = reg_0215;
    40: op1_13_in03 = imem07_in[95:92];
    41: op1_13_in03 = reg_0115;
    42: op1_13_in03 = imem04_in[123:120];
    43: op1_13_in03 = reg_0489;
    44: op1_13_in03 = reg_0677;
    45: op1_13_in03 = reg_0346;
    46: op1_13_in03 = reg_0226;
    47: op1_13_in03 = reg_0686;
    48: op1_13_in03 = reg_0104;
    49: op1_13_in03 = reg_0683;
    50: op1_13_in03 = imem07_in[99:96];
    51: op1_13_in03 = imem05_in[47:44];
    52: op1_13_in03 = reg_0441;
    53: op1_13_in03 = reg_0371;
    54: op1_13_in03 = imem00_in[87:84];
    55: op1_13_in03 = reg_0423;
    56: op1_13_in03 = reg_0105;
    87: op1_13_in03 = reg_0105;
    57: op1_13_in03 = imem00_in[71:68];
    71: op1_13_in03 = imem00_in[71:68];
    78: op1_13_in03 = imem00_in[71:68];
    58: op1_13_in03 = reg_0740;
    59: op1_13_in03 = reg_0123;
    60: op1_13_in03 = reg_0564;
    61: op1_13_in03 = reg_0375;
    63: op1_13_in03 = imem00_in[55:52];
    64: op1_13_in03 = reg_0694;
    65: op1_13_in03 = reg_0306;
    67: op1_13_in03 = reg_0225;
    68: op1_13_in03 = reg_0620;
    69: op1_13_in03 = reg_0125;
    70: op1_13_in03 = reg_0071;
    72: op1_13_in03 = reg_0121;
    73: op1_13_in03 = imem02_in[75:72];
    74: op1_13_in03 = reg_0488;
    75: op1_13_in03 = reg_0416;
    76: op1_13_in03 = reg_0334;
    77: op1_13_in03 = imem00_in[115:112];
    79: op1_13_in03 = reg_0392;
    80: op1_13_in03 = reg_0575;
    81: op1_13_in03 = reg_0204;
    82: op1_13_in03 = reg_0061;
    83: op1_13_in03 = reg_0285;
    84: op1_13_in03 = reg_0108;
    85: op1_13_in03 = reg_0080;
    86: op1_13_in03 = reg_0439;
    88: op1_13_in03 = reg_0712;
    89: op1_13_in03 = imem00_in[99:96];
    90: op1_13_in03 = reg_0634;
    91: op1_13_in03 = imem04_in[71:68];
    92: op1_13_in03 = reg_0245;
    93: op1_13_in03 = reg_0812;
    94: op1_13_in03 = reg_0736;
    95: op1_13_in03 = imem05_in[91:88];
    default: op1_13_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv03 = 1;
    8: op1_13_inv03 = 1;
    9: op1_13_inv03 = 1;
    13: op1_13_inv03 = 1;
    16: op1_13_inv03 = 1;
    18: op1_13_inv03 = 1;
    19: op1_13_inv03 = 1;
    20: op1_13_inv03 = 1;
    21: op1_13_inv03 = 1;
    23: op1_13_inv03 = 1;
    3: op1_13_inv03 = 1;
    27: op1_13_inv03 = 1;
    2: op1_13_inv03 = 1;
    28: op1_13_inv03 = 1;
    31: op1_13_inv03 = 1;
    32: op1_13_inv03 = 1;
    33: op1_13_inv03 = 1;
    35: op1_13_inv03 = 1;
    38: op1_13_inv03 = 1;
    39: op1_13_inv03 = 1;
    40: op1_13_inv03 = 1;
    41: op1_13_inv03 = 1;
    43: op1_13_inv03 = 1;
    44: op1_13_inv03 = 1;
    45: op1_13_inv03 = 1;
    52: op1_13_inv03 = 1;
    54: op1_13_inv03 = 1;
    55: op1_13_inv03 = 1;
    56: op1_13_inv03 = 1;
    60: op1_13_inv03 = 1;
    61: op1_13_inv03 = 1;
    62: op1_13_inv03 = 1;
    64: op1_13_inv03 = 1;
    65: op1_13_inv03 = 1;
    70: op1_13_inv03 = 1;
    72: op1_13_inv03 = 1;
    74: op1_13_inv03 = 1;
    76: op1_13_inv03 = 1;
    77: op1_13_inv03 = 1;
    78: op1_13_inv03 = 1;
    80: op1_13_inv03 = 1;
    81: op1_13_inv03 = 1;
    83: op1_13_inv03 = 1;
    86: op1_13_inv03 = 1;
    89: op1_13_inv03 = 1;
    91: op1_13_inv03 = 1;
    92: op1_13_inv03 = 1;
    93: op1_13_inv03 = 1;
    94: op1_13_inv03 = 1;
    default: op1_13_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in04 = reg_0610;
    5: op1_13_in04 = reg_0282;
    6: op1_13_in04 = reg_0677;
    7: op1_13_in04 = imem02_in[15:12];
    8: op1_13_in04 = reg_0217;
    9: op1_13_in04 = reg_0331;
    10: op1_13_in04 = imem00_in[75:72];
    71: op1_13_in04 = imem00_in[75:72];
    11: op1_13_in04 = imem03_in[35:32];
    12: op1_13_in04 = imem00_in[107:104];
    13: op1_13_in04 = reg_0243;
    14: op1_13_in04 = reg_0369;
    15: op1_13_in04 = reg_0618;
    16: op1_13_in04 = reg_0676;
    17: op1_13_in04 = imem07_in[43:40];
    18: op1_13_in04 = reg_0671;
    19: op1_13_in04 = reg_0703;
    20: op1_13_in04 = reg_0122;
    21: op1_13_in04 = imem04_in[3:0];
    22: op1_13_in04 = imem06_in[75:72];
    23: op1_13_in04 = reg_0482;
    24: op1_13_in04 = reg_0028;
    25: op1_13_in04 = reg_0576;
    3: op1_13_in04 = reg_0440;
    86: op1_13_in04 = reg_0440;
    26: op1_13_in04 = imem00_in[83:80];
    27: op1_13_in04 = reg_0685;
    2: op1_13_in04 = imem07_in[91:88];
    28: op1_13_in04 = imem05_in[79:76];
    29: op1_13_in04 = reg_0153;
    30: op1_13_in04 = reg_0121;
    31: op1_13_in04 = reg_0591;
    32: op1_13_in04 = reg_0015;
    33: op1_13_in04 = reg_0455;
    34: op1_13_in04 = reg_0240;
    35: op1_13_in04 = reg_0118;
    36: op1_13_in04 = reg_0013;
    37: op1_13_in04 = reg_0665;
    38: op1_13_in04 = imem06_in[111:108];
    39: op1_13_in04 = reg_0577;
    40: op1_13_in04 = imem07_in[107:104];
    41: op1_13_in04 = imem02_in[55:52];
    42: op1_13_in04 = imem04_in[127:124];
    43: op1_13_in04 = reg_0091;
    44: op1_13_in04 = reg_0691;
    45: op1_13_in04 = reg_0417;
    46: op1_13_in04 = reg_0276;
    47: op1_13_in04 = reg_0690;
    48: op1_13_in04 = reg_0106;
    49: op1_13_in04 = reg_0681;
    50: op1_13_in04 = imem07_in[127:124];
    51: op1_13_in04 = imem05_in[111:108];
    52: op1_13_in04 = reg_0253;
    53: op1_13_in04 = reg_0298;
    54: op1_13_in04 = imem00_in[95:92];
    55: op1_13_in04 = reg_0418;
    56: op1_13_in04 = reg_0125;
    57: op1_13_in04 = reg_0683;
    58: op1_13_in04 = imem03_in[23:20];
    59: op1_13_in04 = reg_0124;
    60: op1_13_in04 = reg_0562;
    61: op1_13_in04 = reg_0608;
    62: op1_13_in04 = reg_0697;
    89: op1_13_in04 = reg_0697;
    63: op1_13_in04 = imem00_in[103:100];
    64: op1_13_in04 = reg_0117;
    65: op1_13_in04 = reg_0054;
    66: op1_13_in04 = reg_0698;
    67: op1_13_in04 = reg_0224;
    68: op1_13_in04 = reg_0656;
    69: op1_13_in04 = reg_0108;
    70: op1_13_in04 = reg_0292;
    72: op1_13_in04 = reg_0126;
    73: op1_13_in04 = imem02_in[87:84];
    74: op1_13_in04 = reg_0399;
    75: op1_13_in04 = imem05_in[3:0];
    76: op1_13_in04 = reg_0266;
    77: op1_13_in04 = reg_0695;
    78: op1_13_in04 = imem00_in[87:84];
    79: op1_13_in04 = reg_0584;
    80: op1_13_in04 = reg_0568;
    81: op1_13_in04 = reg_0188;
    82: op1_13_in04 = reg_0333;
    83: op1_13_in04 = reg_0147;
    84: op1_13_in04 = reg_0660;
    85: op1_13_in04 = reg_0530;
    87: op1_13_in04 = reg_0104;
    88: op1_13_in04 = reg_0164;
    90: op1_13_in04 = imem00_in[35:32];
    91: op1_13_in04 = imem04_in[99:96];
    92: op1_13_in04 = reg_0583;
    93: op1_13_in04 = reg_0149;
    94: op1_13_in04 = reg_0135;
    95: op1_13_in04 = imem05_in[127:124];
    default: op1_13_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv04 = 1;
    8: op1_13_inv04 = 1;
    9: op1_13_inv04 = 1;
    11: op1_13_inv04 = 1;
    13: op1_13_inv04 = 1;
    14: op1_13_inv04 = 1;
    18: op1_13_inv04 = 1;
    19: op1_13_inv04 = 1;
    22: op1_13_inv04 = 1;
    25: op1_13_inv04 = 1;
    26: op1_13_inv04 = 1;
    27: op1_13_inv04 = 1;
    2: op1_13_inv04 = 1;
    30: op1_13_inv04 = 1;
    31: op1_13_inv04 = 1;
    32: op1_13_inv04 = 1;
    33: op1_13_inv04 = 1;
    34: op1_13_inv04 = 1;
    35: op1_13_inv04 = 1;
    36: op1_13_inv04 = 1;
    39: op1_13_inv04 = 1;
    41: op1_13_inv04 = 1;
    42: op1_13_inv04 = 1;
    43: op1_13_inv04 = 1;
    44: op1_13_inv04 = 1;
    45: op1_13_inv04 = 1;
    47: op1_13_inv04 = 1;
    48: op1_13_inv04 = 1;
    49: op1_13_inv04 = 1;
    50: op1_13_inv04 = 1;
    52: op1_13_inv04 = 1;
    53: op1_13_inv04 = 1;
    57: op1_13_inv04 = 1;
    60: op1_13_inv04 = 1;
    61: op1_13_inv04 = 1;
    63: op1_13_inv04 = 1;
    64: op1_13_inv04 = 1;
    65: op1_13_inv04 = 1;
    66: op1_13_inv04 = 1;
    67: op1_13_inv04 = 1;
    69: op1_13_inv04 = 1;
    71: op1_13_inv04 = 1;
    72: op1_13_inv04 = 1;
    73: op1_13_inv04 = 1;
    74: op1_13_inv04 = 1;
    79: op1_13_inv04 = 1;
    80: op1_13_inv04 = 1;
    82: op1_13_inv04 = 1;
    83: op1_13_inv04 = 1;
    84: op1_13_inv04 = 1;
    86: op1_13_inv04 = 1;
    87: op1_13_inv04 = 1;
    88: op1_13_inv04 = 1;
    89: op1_13_inv04 = 1;
    90: op1_13_inv04 = 1;
    93: op1_13_inv04 = 1;
    95: op1_13_inv04 = 1;
    default: op1_13_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in05 = reg_0624;
    5: op1_13_in05 = reg_0306;
    6: op1_13_in05 = reg_0678;
    18: op1_13_in05 = reg_0678;
    7: op1_13_in05 = imem02_in[43:40];
    8: op1_13_in05 = reg_0218;
    9: op1_13_in05 = reg_0001;
    10: op1_13_in05 = imem00_in[115:112];
    11: op1_13_in05 = imem03_in[59:56];
    12: op1_13_in05 = reg_0672;
    13: op1_13_in05 = reg_0125;
    14: op1_13_in05 = reg_0385;
    15: op1_13_in05 = reg_0601;
    16: op1_13_in05 = reg_0689;
    17: op1_13_in05 = imem07_in[107:104];
    19: op1_13_in05 = reg_0724;
    20: op1_13_in05 = reg_0111;
    21: op1_13_in05 = imem04_in[47:44];
    22: op1_13_in05 = imem06_in[79:76];
    23: op1_13_in05 = reg_0483;
    24: op1_13_in05 = reg_0815;
    25: op1_13_in05 = reg_0395;
    3: op1_13_in05 = reg_0444;
    26: op1_13_in05 = imem00_in[87:84];
    27: op1_13_in05 = reg_0690;
    62: op1_13_in05 = reg_0690;
    2: op1_13_in05 = imem07_in[95:92];
    28: op1_13_in05 = imem05_in[87:84];
    29: op1_13_in05 = reg_0140;
    30: op1_13_in05 = imem02_in[7:4];
    31: op1_13_in05 = reg_0600;
    32: op1_13_in05 = imem04_in[23:20];
    33: op1_13_in05 = reg_0469;
    34: op1_13_in05 = reg_0238;
    35: op1_13_in05 = reg_0117;
    36: op1_13_in05 = imem04_in[7:4];
    37: op1_13_in05 = reg_0636;
    76: op1_13_in05 = reg_0636;
    38: op1_13_in05 = reg_0402;
    39: op1_13_in05 = reg_0405;
    40: op1_13_in05 = imem07_in[111:108];
    41: op1_13_in05 = imem02_in[71:68];
    42: op1_13_in05 = reg_0328;
    43: op1_13_in05 = reg_0225;
    44: op1_13_in05 = reg_0688;
    45: op1_13_in05 = reg_0349;
    46: op1_13_in05 = reg_0733;
    47: op1_13_in05 = reg_0668;
    48: op1_13_in05 = reg_0115;
    49: op1_13_in05 = reg_0694;
    57: op1_13_in05 = reg_0694;
    50: op1_13_in05 = reg_0730;
    51: op1_13_in05 = reg_0488;
    52: op1_13_in05 = reg_0295;
    53: op1_13_in05 = reg_0408;
    54: op1_13_in05 = reg_0463;
    55: op1_13_in05 = reg_0217;
    56: op1_13_in05 = reg_0104;
    58: op1_13_in05 = imem03_in[35:32];
    59: op1_13_in05 = reg_0127;
    60: op1_13_in05 = reg_0572;
    61: op1_13_in05 = reg_0638;
    63: op1_13_in05 = imem00_in[123:120];
    64: op1_13_in05 = reg_0692;
    65: op1_13_in05 = reg_0567;
    66: op1_13_in05 = reg_0744;
    67: op1_13_in05 = imem05_in[3:0];
    68: op1_13_in05 = reg_0368;
    69: op1_13_in05 = reg_0660;
    87: op1_13_in05 = reg_0660;
    70: op1_13_in05 = reg_0050;
    71: op1_13_in05 = imem00_in[83:80];
    72: op1_13_in05 = imem02_in[3:0];
    73: op1_13_in05 = imem02_in[99:96];
    74: op1_13_in05 = reg_0595;
    75: op1_13_in05 = imem05_in[19:16];
    77: op1_13_in05 = reg_0682;
    78: op1_13_in05 = imem00_in[95:92];
    79: op1_13_in05 = reg_0141;
    80: op1_13_in05 = reg_0396;
    81: op1_13_in05 = reg_0193;
    82: op1_13_in05 = reg_0449;
    83: op1_13_in05 = imem06_in[47:44];
    84: op1_13_in05 = reg_0669;
    85: op1_13_in05 = reg_0639;
    86: op1_13_in05 = reg_0084;
    88: op1_13_in05 = reg_0709;
    89: op1_13_in05 = reg_0685;
    90: op1_13_in05 = imem00_in[51:48];
    91: op1_13_in05 = reg_0262;
    92: op1_13_in05 = reg_0751;
    93: op1_13_in05 = reg_0825;
    94: op1_13_in05 = reg_0788;
    95: op1_13_in05 = reg_0791;
    default: op1_13_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv05 = 1;
    8: op1_13_inv05 = 1;
    9: op1_13_inv05 = 1;
    11: op1_13_inv05 = 1;
    14: op1_13_inv05 = 1;
    15: op1_13_inv05 = 1;
    16: op1_13_inv05 = 1;
    20: op1_13_inv05 = 1;
    21: op1_13_inv05 = 1;
    3: op1_13_inv05 = 1;
    26: op1_13_inv05 = 1;
    27: op1_13_inv05 = 1;
    2: op1_13_inv05 = 1;
    28: op1_13_inv05 = 1;
    29: op1_13_inv05 = 1;
    31: op1_13_inv05 = 1;
    32: op1_13_inv05 = 1;
    33: op1_13_inv05 = 1;
    34: op1_13_inv05 = 1;
    40: op1_13_inv05 = 1;
    42: op1_13_inv05 = 1;
    44: op1_13_inv05 = 1;
    45: op1_13_inv05 = 1;
    46: op1_13_inv05 = 1;
    48: op1_13_inv05 = 1;
    51: op1_13_inv05 = 1;
    53: op1_13_inv05 = 1;
    54: op1_13_inv05 = 1;
    56: op1_13_inv05 = 1;
    58: op1_13_inv05 = 1;
    59: op1_13_inv05 = 1;
    60: op1_13_inv05 = 1;
    61: op1_13_inv05 = 1;
    63: op1_13_inv05 = 1;
    67: op1_13_inv05 = 1;
    68: op1_13_inv05 = 1;
    69: op1_13_inv05 = 1;
    73: op1_13_inv05 = 1;
    74: op1_13_inv05 = 1;
    77: op1_13_inv05 = 1;
    78: op1_13_inv05 = 1;
    79: op1_13_inv05 = 1;
    84: op1_13_inv05 = 1;
    85: op1_13_inv05 = 1;
    87: op1_13_inv05 = 1;
    89: op1_13_inv05 = 1;
    94: op1_13_inv05 = 1;
    default: op1_13_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in06 = reg_0611;
    5: op1_13_in06 = reg_0275;
    6: op1_13_in06 = reg_0450;
    44: op1_13_in06 = reg_0450;
    89: op1_13_in06 = reg_0450;
    7: op1_13_in06 = imem02_in[47:44];
    8: op1_13_in06 = reg_0215;
    9: op1_13_in06 = imem04_in[11:8];
    10: op1_13_in06 = imem00_in[119:116];
    11: op1_13_in06 = imem03_in[103:100];
    12: op1_13_in06 = reg_0698;
    49: op1_13_in06 = reg_0698;
    13: op1_13_in06 = reg_0112;
    20: op1_13_in06 = reg_0112;
    14: op1_13_in06 = reg_0312;
    15: op1_13_in06 = reg_0402;
    16: op1_13_in06 = reg_0677;
    56: op1_13_in06 = reg_0677;
    17: op1_13_in06 = reg_0704;
    40: op1_13_in06 = reg_0704;
    18: op1_13_in06 = reg_0476;
    19: op1_13_in06 = reg_0432;
    21: op1_13_in06 = imem04_in[59:56];
    22: op1_13_in06 = imem06_in[95:92];
    23: op1_13_in06 = reg_0491;
    51: op1_13_in06 = reg_0491;
    24: op1_13_in06 = reg_0814;
    25: op1_13_in06 = reg_0373;
    3: op1_13_in06 = reg_0443;
    26: op1_13_in06 = imem00_in[95:92];
    71: op1_13_in06 = imem00_in[95:92];
    27: op1_13_in06 = reg_0477;
    2: op1_13_in06 = imem07_in[99:96];
    28: op1_13_in06 = reg_0781;
    29: op1_13_in06 = reg_0155;
    30: op1_13_in06 = imem02_in[39:36];
    72: op1_13_in06 = imem02_in[39:36];
    31: op1_13_in06 = reg_0578;
    32: op1_13_in06 = imem04_in[47:44];
    33: op1_13_in06 = reg_0460;
    34: op1_13_in06 = reg_0105;
    35: op1_13_in06 = imem02_in[7:4];
    69: op1_13_in06 = imem02_in[7:4];
    36: op1_13_in06 = imem04_in[31:28];
    37: op1_13_in06 = reg_0663;
    38: op1_13_in06 = reg_0270;
    39: op1_13_in06 = reg_0775;
    41: op1_13_in06 = imem02_in[91:88];
    42: op1_13_in06 = reg_0536;
    43: op1_13_in06 = reg_0736;
    45: op1_13_in06 = reg_0358;
    46: op1_13_in06 = reg_0277;
    47: op1_13_in06 = reg_0680;
    48: op1_13_in06 = reg_0110;
    50: op1_13_in06 = reg_0729;
    52: op1_13_in06 = reg_0067;
    53: op1_13_in06 = reg_0748;
    54: op1_13_in06 = reg_0451;
    55: op1_13_in06 = reg_0603;
    57: op1_13_in06 = reg_0689;
    58: op1_13_in06 = imem03_in[87:84];
    59: op1_13_in06 = reg_0674;
    60: op1_13_in06 = reg_0019;
    61: op1_13_in06 = reg_0580;
    62: op1_13_in06 = reg_0633;
    63: op1_13_in06 = imem00_in[127:124];
    64: op1_13_in06 = reg_0634;
    65: op1_13_in06 = reg_0248;
    66: op1_13_in06 = reg_0658;
    67: op1_13_in06 = imem05_in[7:4];
    68: op1_13_in06 = reg_0752;
    70: op1_13_in06 = reg_0062;
    73: op1_13_in06 = imem02_in[111:108];
    74: op1_13_in06 = reg_0575;
    75: op1_13_in06 = imem05_in[27:24];
    76: op1_13_in06 = reg_0053;
    77: op1_13_in06 = reg_0693;
    78: op1_13_in06 = reg_0697;
    79: op1_13_in06 = reg_0140;
    80: op1_13_in06 = reg_0570;
    81: op1_13_in06 = reg_0207;
    82: op1_13_in06 = reg_0444;
    83: op1_13_in06 = imem06_in[59:56];
    84: op1_13_in06 = reg_0601;
    85: op1_13_in06 = reg_0753;
    86: op1_13_in06 = reg_0437;
    87: op1_13_in06 = reg_0678;
    88: op1_13_in06 = reg_0713;
    90: op1_13_in06 = imem00_in[63:60];
    91: op1_13_in06 = reg_0544;
    92: op1_13_in06 = reg_0579;
    93: op1_13_in06 = reg_0796;
    94: op1_13_in06 = reg_0793;
    95: op1_13_in06 = reg_0133;
    default: op1_13_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv06 = 1;
    5: op1_13_inv06 = 1;
    7: op1_13_inv06 = 1;
    9: op1_13_inv06 = 1;
    11: op1_13_inv06 = 1;
    15: op1_13_inv06 = 1;
    18: op1_13_inv06 = 1;
    20: op1_13_inv06 = 1;
    22: op1_13_inv06 = 1;
    24: op1_13_inv06 = 1;
    25: op1_13_inv06 = 1;
    3: op1_13_inv06 = 1;
    26: op1_13_inv06 = 1;
    27: op1_13_inv06 = 1;
    2: op1_13_inv06 = 1;
    28: op1_13_inv06 = 1;
    34: op1_13_inv06 = 1;
    35: op1_13_inv06 = 1;
    38: op1_13_inv06 = 1;
    39: op1_13_inv06 = 1;
    40: op1_13_inv06 = 1;
    41: op1_13_inv06 = 1;
    43: op1_13_inv06 = 1;
    50: op1_13_inv06 = 1;
    51: op1_13_inv06 = 1;
    53: op1_13_inv06 = 1;
    54: op1_13_inv06 = 1;
    55: op1_13_inv06 = 1;
    58: op1_13_inv06 = 1;
    59: op1_13_inv06 = 1;
    60: op1_13_inv06 = 1;
    61: op1_13_inv06 = 1;
    62: op1_13_inv06 = 1;
    67: op1_13_inv06 = 1;
    68: op1_13_inv06 = 1;
    69: op1_13_inv06 = 1;
    70: op1_13_inv06 = 1;
    73: op1_13_inv06 = 1;
    78: op1_13_inv06 = 1;
    81: op1_13_inv06 = 1;
    85: op1_13_inv06 = 1;
    87: op1_13_inv06 = 1;
    89: op1_13_inv06 = 1;
    94: op1_13_inv06 = 1;
    default: op1_13_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in07 = reg_0623;
    5: op1_13_in07 = reg_0062;
    6: op1_13_in07 = reg_0473;
    7: op1_13_in07 = imem02_in[71:68];
    8: op1_13_in07 = reg_0628;
    9: op1_13_in07 = imem04_in[55:52];
    10: op1_13_in07 = reg_0695;
    11: op1_13_in07 = reg_0583;
    12: op1_13_in07 = reg_0691;
    13: op1_13_in07 = reg_0106;
    14: op1_13_in07 = reg_0006;
    15: op1_13_in07 = reg_0372;
    16: op1_13_in07 = reg_0671;
    17: op1_13_in07 = reg_0719;
    18: op1_13_in07 = reg_0462;
    19: op1_13_in07 = reg_0183;
    20: op1_13_in07 = reg_0114;
    21: op1_13_in07 = imem04_in[67:64];
    22: op1_13_in07 = reg_0626;
    23: op1_13_in07 = reg_0795;
    24: op1_13_in07 = reg_0750;
    25: op1_13_in07 = reg_0376;
    3: op1_13_in07 = reg_0448;
    26: op1_13_in07 = imem00_in[111:108];
    27: op1_13_in07 = reg_0466;
    2: op1_13_in07 = imem07_in[107:104];
    28: op1_13_in07 = reg_0780;
    29: op1_13_in07 = reg_0137;
    93: op1_13_in07 = reg_0137;
    30: op1_13_in07 = imem02_in[43:40];
    31: op1_13_in07 = reg_0588;
    32: op1_13_in07 = imem04_in[51:48];
    33: op1_13_in07 = reg_0458;
    34: op1_13_in07 = reg_0102;
    35: op1_13_in07 = imem02_in[19:16];
    87: op1_13_in07 = imem02_in[19:16];
    36: op1_13_in07 = imem04_in[63:60];
    37: op1_13_in07 = reg_0530;
    38: op1_13_in07 = reg_0776;
    39: op1_13_in07 = reg_0776;
    40: op1_13_in07 = reg_0726;
    41: op1_13_in07 = imem02_in[127:124];
    42: op1_13_in07 = reg_0556;
    43: op1_13_in07 = reg_0737;
    44: op1_13_in07 = reg_0455;
    45: op1_13_in07 = reg_0356;
    46: op1_13_in07 = reg_0285;
    47: op1_13_in07 = reg_0454;
    48: op1_13_in07 = imem02_in[11:8];
    49: op1_13_in07 = reg_0679;
    50: op1_13_in07 = reg_0715;
    51: op1_13_in07 = reg_0493;
    52: op1_13_in07 = reg_0442;
    53: op1_13_in07 = reg_0319;
    54: op1_13_in07 = reg_0464;
    55: op1_13_in07 = reg_0419;
    56: op1_13_in07 = reg_0669;
    57: op1_13_in07 = reg_0744;
    58: op1_13_in07 = imem03_in[119:116];
    59: op1_13_in07 = imem02_in[47:44];
    60: op1_13_in07 = reg_0012;
    80: op1_13_in07 = reg_0012;
    61: op1_13_in07 = reg_0515;
    62: op1_13_in07 = reg_0692;
    63: op1_13_in07 = reg_0683;
    78: op1_13_in07 = reg_0683;
    64: op1_13_in07 = reg_0451;
    65: op1_13_in07 = reg_0603;
    66: op1_13_in07 = reg_0481;
    67: op1_13_in07 = imem05_in[35:32];
    68: op1_13_in07 = imem07_in[3:0];
    69: op1_13_in07 = imem02_in[51:48];
    70: op1_13_in07 = reg_0687;
    71: op1_13_in07 = imem00_in[99:96];
    72: op1_13_in07 = imem02_in[55:52];
    73: op1_13_in07 = imem02_in[115:112];
    74: op1_13_in07 = reg_0562;
    75: op1_13_in07 = imem05_in[31:28];
    76: op1_13_in07 = reg_0439;
    77: op1_13_in07 = reg_0689;
    79: op1_13_in07 = reg_0304;
    81: op1_13_in07 = imem01_in[19:16];
    82: op1_13_in07 = reg_0267;
    83: op1_13_in07 = imem06_in[87:84];
    84: op1_13_in07 = reg_0126;
    85: op1_13_in07 = reg_0083;
    86: op1_13_in07 = reg_0139;
    88: op1_13_in07 = reg_0158;
    89: op1_13_in07 = reg_0460;
    90: op1_13_in07 = imem00_in[67:64];
    91: op1_13_in07 = reg_0177;
    92: op1_13_in07 = reg_0560;
    94: op1_13_in07 = reg_0113;
    95: op1_13_in07 = reg_0666;
    default: op1_13_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv07 = 1;
    5: op1_13_inv07 = 1;
    8: op1_13_inv07 = 1;
    9: op1_13_inv07 = 1;
    10: op1_13_inv07 = 1;
    11: op1_13_inv07 = 1;
    13: op1_13_inv07 = 1;
    14: op1_13_inv07 = 1;
    15: op1_13_inv07 = 1;
    16: op1_13_inv07 = 1;
    19: op1_13_inv07 = 1;
    21: op1_13_inv07 = 1;
    23: op1_13_inv07 = 1;
    25: op1_13_inv07 = 1;
    3: op1_13_inv07 = 1;
    28: op1_13_inv07 = 1;
    34: op1_13_inv07 = 1;
    38: op1_13_inv07 = 1;
    39: op1_13_inv07 = 1;
    40: op1_13_inv07 = 1;
    41: op1_13_inv07 = 1;
    43: op1_13_inv07 = 1;
    44: op1_13_inv07 = 1;
    46: op1_13_inv07 = 1;
    47: op1_13_inv07 = 1;
    48: op1_13_inv07 = 1;
    52: op1_13_inv07 = 1;
    53: op1_13_inv07 = 1;
    54: op1_13_inv07 = 1;
    55: op1_13_inv07 = 1;
    56: op1_13_inv07 = 1;
    57: op1_13_inv07 = 1;
    59: op1_13_inv07 = 1;
    60: op1_13_inv07 = 1;
    61: op1_13_inv07 = 1;
    62: op1_13_inv07 = 1;
    63: op1_13_inv07 = 1;
    65: op1_13_inv07 = 1;
    66: op1_13_inv07 = 1;
    67: op1_13_inv07 = 1;
    70: op1_13_inv07 = 1;
    72: op1_13_inv07 = 1;
    73: op1_13_inv07 = 1;
    75: op1_13_inv07 = 1;
    76: op1_13_inv07 = 1;
    79: op1_13_inv07 = 1;
    82: op1_13_inv07 = 1;
    83: op1_13_inv07 = 1;
    84: op1_13_inv07 = 1;
    89: op1_13_inv07 = 1;
    91: op1_13_inv07 = 1;
    93: op1_13_inv07 = 1;
    94: op1_13_inv07 = 1;
    95: op1_13_inv07 = 1;
    default: op1_13_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in08 = reg_0612;
    5: op1_13_in08 = reg_0067;
    6: op1_13_in08 = reg_0470;
    7: op1_13_in08 = imem02_in[75:72];
    8: op1_13_in08 = reg_0604;
    9: op1_13_in08 = imem04_in[59:56];
    10: op1_13_in08 = reg_0683;
    11: op1_13_in08 = reg_0592;
    12: op1_13_in08 = reg_0678;
    13: op1_13_in08 = reg_0109;
    14: op1_13_in08 = reg_0003;
    15: op1_13_in08 = reg_0368;
    16: op1_13_in08 = reg_0668;
    17: op1_13_in08 = reg_0717;
    18: op1_13_in08 = reg_0481;
    19: op1_13_in08 = reg_0166;
    20: op1_13_in08 = reg_0101;
    21: op1_13_in08 = imem04_in[71:68];
    22: op1_13_in08 = reg_0619;
    23: op1_13_in08 = reg_0780;
    24: op1_13_in08 = reg_0749;
    77: op1_13_in08 = reg_0749;
    25: op1_13_in08 = reg_0019;
    3: op1_13_in08 = reg_0182;
    26: op1_13_in08 = imem00_in[119:116];
    27: op1_13_in08 = reg_0462;
    54: op1_13_in08 = reg_0462;
    2: op1_13_in08 = imem07_in[115:112];
    28: op1_13_in08 = reg_0786;
    29: op1_13_in08 = imem06_in[35:32];
    30: op1_13_in08 = imem02_in[59:56];
    31: op1_13_in08 = reg_0751;
    32: op1_13_in08 = imem04_in[87:84];
    33: op1_13_in08 = reg_0191;
    34: op1_13_in08 = reg_0126;
    35: op1_13_in08 = imem02_in[115:112];
    36: op1_13_in08 = imem04_in[111:108];
    37: op1_13_in08 = reg_0535;
    38: op1_13_in08 = reg_0372;
    39: op1_13_in08 = reg_0404;
    40: op1_13_in08 = reg_0729;
    41: op1_13_in08 = reg_0645;
    42: op1_13_in08 = reg_0429;
    43: op1_13_in08 = reg_0733;
    44: op1_13_in08 = reg_0464;
    45: op1_13_in08 = reg_0363;
    46: op1_13_in08 = reg_0147;
    47: op1_13_in08 = reg_0450;
    48: op1_13_in08 = imem02_in[19:16];
    49: op1_13_in08 = reg_0691;
    57: op1_13_in08 = reg_0691;
    50: op1_13_in08 = reg_0266;
    51: op1_13_in08 = reg_0793;
    52: op1_13_in08 = reg_0443;
    76: op1_13_in08 = reg_0443;
    53: op1_13_in08 = reg_0038;
    55: op1_13_in08 = reg_0243;
    56: op1_13_in08 = reg_0107;
    58: op1_13_in08 = reg_0596;
    59: op1_13_in08 = imem02_in[79:76];
    60: op1_13_in08 = reg_0013;
    61: op1_13_in08 = reg_0819;
    62: op1_13_in08 = reg_0463;
    63: op1_13_in08 = reg_0658;
    64: op1_13_in08 = reg_0477;
    65: op1_13_in08 = reg_0506;
    66: op1_13_in08 = reg_0480;
    67: op1_13_in08 = imem05_in[63:60];
    68: op1_13_in08 = imem07_in[19:16];
    69: op1_13_in08 = imem02_in[87:84];
    70: op1_13_in08 = reg_0513;
    71: op1_13_in08 = reg_0697;
    72: op1_13_in08 = imem02_in[111:108];
    73: op1_13_in08 = reg_0642;
    74: op1_13_in08 = reg_0496;
    75: op1_13_in08 = imem05_in[47:44];
    78: op1_13_in08 = reg_0685;
    79: op1_13_in08 = reg_0548;
    91: op1_13_in08 = reg_0548;
    80: op1_13_in08 = reg_0803;
    81: op1_13_in08 = imem01_in[35:32];
    82: op1_13_in08 = reg_0175;
    83: op1_13_in08 = reg_0625;
    84: op1_13_in08 = reg_0169;
    85: op1_13_in08 = reg_0485;
    86: op1_13_in08 = reg_0327;
    87: op1_13_in08 = imem02_in[71:68];
    88: op1_13_in08 = reg_0053;
    89: op1_13_in08 = reg_0214;
    90: op1_13_in08 = imem00_in[71:68];
    92: op1_13_in08 = reg_0812;
    93: op1_13_in08 = reg_0734;
    94: op1_13_in08 = reg_0782;
    95: op1_13_in08 = reg_0795;
    default: op1_13_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv08 = 1;
    10: op1_13_inv08 = 1;
    11: op1_13_inv08 = 1;
    18: op1_13_inv08 = 1;
    19: op1_13_inv08 = 1;
    21: op1_13_inv08 = 1;
    23: op1_13_inv08 = 1;
    25: op1_13_inv08 = 1;
    3: op1_13_inv08 = 1;
    2: op1_13_inv08 = 1;
    28: op1_13_inv08 = 1;
    29: op1_13_inv08 = 1;
    30: op1_13_inv08 = 1;
    33: op1_13_inv08 = 1;
    34: op1_13_inv08 = 1;
    37: op1_13_inv08 = 1;
    38: op1_13_inv08 = 1;
    39: op1_13_inv08 = 1;
    43: op1_13_inv08 = 1;
    44: op1_13_inv08 = 1;
    45: op1_13_inv08 = 1;
    46: op1_13_inv08 = 1;
    48: op1_13_inv08 = 1;
    52: op1_13_inv08 = 1;
    53: op1_13_inv08 = 1;
    61: op1_13_inv08 = 1;
    63: op1_13_inv08 = 1;
    64: op1_13_inv08 = 1;
    66: op1_13_inv08 = 1;
    67: op1_13_inv08 = 1;
    76: op1_13_inv08 = 1;
    78: op1_13_inv08 = 1;
    79: op1_13_inv08 = 1;
    80: op1_13_inv08 = 1;
    81: op1_13_inv08 = 1;
    82: op1_13_inv08 = 1;
    84: op1_13_inv08 = 1;
    86: op1_13_inv08 = 1;
    88: op1_13_inv08 = 1;
    89: op1_13_inv08 = 1;
    90: op1_13_inv08 = 1;
    default: op1_13_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in09 = reg_0379;
    5: op1_13_in09 = reg_0056;
    6: op1_13_in09 = reg_0479;
    7: op1_13_in09 = imem02_in[119:116];
    8: op1_13_in09 = reg_0607;
    9: op1_13_in09 = imem04_in[115:112];
    10: op1_13_in09 = reg_0690;
    11: op1_13_in09 = reg_0600;
    12: op1_13_in09 = reg_0457;
    13: op1_13_in09 = imem02_in[3:0];
    14: op1_13_in09 = reg_0803;
    15: op1_13_in09 = reg_0813;
    16: op1_13_in09 = reg_0461;
    17: op1_13_in09 = reg_0703;
    18: op1_13_in09 = reg_0472;
    19: op1_13_in09 = reg_0164;
    20: op1_13_in09 = reg_0107;
    21: op1_13_in09 = imem04_in[79:76];
    22: op1_13_in09 = reg_0632;
    23: op1_13_in09 = reg_0785;
    69: op1_13_in09 = reg_0785;
    24: op1_13_in09 = imem07_in[3:0];
    25: op1_13_in09 = reg_0001;
    26: op1_13_in09 = reg_0697;
    27: op1_13_in09 = reg_0200;
    2: op1_13_in09 = reg_0159;
    28: op1_13_in09 = reg_0486;
    29: op1_13_in09 = imem06_in[71:68];
    30: op1_13_in09 = imem02_in[87:84];
    59: op1_13_in09 = imem02_in[87:84];
    87: op1_13_in09 = imem02_in[87:84];
    31: op1_13_in09 = reg_0385;
    32: op1_13_in09 = imem04_in[99:96];
    33: op1_13_in09 = imem01_in[3:0];
    34: op1_13_in09 = imem02_in[19:16];
    56: op1_13_in09 = imem02_in[19:16];
    35: op1_13_in09 = imem02_in[127:124];
    36: op1_13_in09 = reg_0560;
    37: op1_13_in09 = reg_0539;
    38: op1_13_in09 = reg_0777;
    39: op1_13_in09 = reg_0242;
    40: op1_13_in09 = reg_0705;
    41: op1_13_in09 = reg_0653;
    42: op1_13_in09 = reg_0076;
    43: op1_13_in09 = reg_0734;
    44: op1_13_in09 = reg_0460;
    45: op1_13_in09 = reg_0365;
    46: op1_13_in09 = reg_0146;
    47: op1_13_in09 = reg_0474;
    48: op1_13_in09 = imem02_in[43:40];
    49: op1_13_in09 = reg_0671;
    50: op1_13_in09 = reg_0295;
    51: op1_13_in09 = reg_0794;
    52: op1_13_in09 = reg_0438;
    53: op1_13_in09 = reg_0576;
    54: op1_13_in09 = reg_0480;
    55: op1_13_in09 = reg_0675;
    57: op1_13_in09 = reg_0758;
    77: op1_13_in09 = reg_0758;
    58: op1_13_in09 = reg_0384;
    60: op1_13_in09 = reg_0804;
    61: op1_13_in09 = reg_0642;
    62: op1_13_in09 = reg_0450;
    63: op1_13_in09 = reg_0407;
    64: op1_13_in09 = reg_0475;
    65: op1_13_in09 = reg_0243;
    66: op1_13_in09 = reg_0468;
    67: op1_13_in09 = imem05_in[67:64];
    68: op1_13_in09 = imem07_in[23:20];
    70: op1_13_in09 = reg_0640;
    71: op1_13_in09 = reg_0492;
    72: op1_13_in09 = reg_0325;
    73: op1_13_in09 = reg_0702;
    74: op1_13_in09 = reg_0396;
    75: op1_13_in09 = imem05_in[55:52];
    76: op1_13_in09 = reg_0165;
    84: op1_13_in09 = reg_0165;
    78: op1_13_in09 = reg_0694;
    79: op1_13_in09 = reg_0374;
    80: op1_13_in09 = reg_0805;
    81: op1_13_in09 = imem01_in[43:40];
    82: op1_13_in09 = reg_0236;
    83: op1_13_in09 = reg_0349;
    85: op1_13_in09 = reg_0320;
    86: op1_13_in09 = reg_0183;
    88: op1_13_in09 = reg_0445;
    89: op1_13_in09 = reg_0211;
    90: op1_13_in09 = imem00_in[111:108];
    91: op1_13_in09 = reg_0555;
    92: op1_13_in09 = reg_0149;
    93: op1_13_in09 = imem06_in[15:12];
    94: op1_13_in09 = reg_0134;
    95: op1_13_in09 = reg_0793;
    default: op1_13_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv09 = 1;
    5: op1_13_inv09 = 1;
    6: op1_13_inv09 = 1;
    8: op1_13_inv09 = 1;
    9: op1_13_inv09 = 1;
    11: op1_13_inv09 = 1;
    13: op1_13_inv09 = 1;
    17: op1_13_inv09 = 1;
    18: op1_13_inv09 = 1;
    20: op1_13_inv09 = 1;
    22: op1_13_inv09 = 1;
    23: op1_13_inv09 = 1;
    25: op1_13_inv09 = 1;
    27: op1_13_inv09 = 1;
    2: op1_13_inv09 = 1;
    30: op1_13_inv09 = 1;
    31: op1_13_inv09 = 1;
    33: op1_13_inv09 = 1;
    35: op1_13_inv09 = 1;
    37: op1_13_inv09 = 1;
    38: op1_13_inv09 = 1;
    39: op1_13_inv09 = 1;
    41: op1_13_inv09 = 1;
    42: op1_13_inv09 = 1;
    43: op1_13_inv09 = 1;
    47: op1_13_inv09 = 1;
    50: op1_13_inv09 = 1;
    53: op1_13_inv09 = 1;
    54: op1_13_inv09 = 1;
    57: op1_13_inv09 = 1;
    58: op1_13_inv09 = 1;
    59: op1_13_inv09 = 1;
    60: op1_13_inv09 = 1;
    61: op1_13_inv09 = 1;
    63: op1_13_inv09 = 1;
    66: op1_13_inv09 = 1;
    68: op1_13_inv09 = 1;
    70: op1_13_inv09 = 1;
    73: op1_13_inv09 = 1;
    74: op1_13_inv09 = 1;
    75: op1_13_inv09 = 1;
    76: op1_13_inv09 = 1;
    77: op1_13_inv09 = 1;
    78: op1_13_inv09 = 1;
    79: op1_13_inv09 = 1;
    83: op1_13_inv09 = 1;
    84: op1_13_inv09 = 1;
    86: op1_13_inv09 = 1;
    89: op1_13_inv09 = 1;
    91: op1_13_inv09 = 1;
    default: op1_13_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in10 = reg_0381;
    5: op1_13_in10 = reg_0068;
    6: op1_13_in10 = reg_0211;
    7: op1_13_in10 = reg_0658;
    8: op1_13_in10 = reg_0605;
    9: op1_13_in10 = reg_0540;
    10: op1_13_in10 = reg_0678;
    11: op1_13_in10 = reg_0578;
    12: op1_13_in10 = reg_0466;
    13: op1_13_in10 = imem02_in[43:40];
    14: op1_13_in10 = reg_0807;
    15: op1_13_in10 = reg_0815;
    16: op1_13_in10 = reg_0460;
    17: op1_13_in10 = reg_0724;
    18: op1_13_in10 = reg_0204;
    19: op1_13_in10 = reg_0178;
    20: op1_13_in10 = reg_0056;
    21: op1_13_in10 = imem04_in[87:84];
    22: op1_13_in10 = reg_0332;
    23: op1_13_in10 = reg_0794;
    24: op1_13_in10 = imem07_in[23:20];
    25: op1_13_in10 = reg_0003;
    26: op1_13_in10 = reg_0672;
    27: op1_13_in10 = reg_0188;
    2: op1_13_in10 = reg_0160;
    28: op1_13_in10 = reg_0090;
    29: op1_13_in10 = reg_0610;
    30: op1_13_in10 = imem02_in[91:88];
    31: op1_13_in10 = reg_0397;
    32: op1_13_in10 = imem04_in[111:108];
    33: op1_13_in10 = imem01_in[7:4];
    34: op1_13_in10 = imem02_in[35:32];
    35: op1_13_in10 = reg_0646;
    36: op1_13_in10 = reg_0542;
    37: op1_13_in10 = imem03_in[59:56];
    38: op1_13_in10 = reg_0814;
    39: op1_13_in10 = reg_0620;
    40: op1_13_in10 = reg_0718;
    41: op1_13_in10 = reg_0663;
    42: op1_13_in10 = reg_0077;
    43: op1_13_in10 = reg_0132;
    44: op1_13_in10 = reg_0480;
    45: op1_13_in10 = reg_0321;
    46: op1_13_in10 = reg_0139;
    47: op1_13_in10 = reg_0479;
    48: op1_13_in10 = reg_0666;
    49: op1_13_in10 = reg_0688;
    50: op1_13_in10 = reg_0436;
    51: op1_13_in10 = reg_0790;
    52: op1_13_in10 = reg_0165;
    53: op1_13_in10 = reg_0621;
    54: op1_13_in10 = reg_0473;
    55: op1_13_in10 = reg_0669;
    56: op1_13_in10 = imem02_in[63:60];
    57: op1_13_in10 = reg_0633;
    58: op1_13_in10 = reg_0392;
    59: op1_13_in10 = imem02_in[111:108];
    60: op1_13_in10 = reg_0805;
    61: op1_13_in10 = reg_0021;
    62: op1_13_in10 = reg_0455;
    63: op1_13_in10 = reg_0247;
    64: op1_13_in10 = reg_0472;
    65: op1_13_in10 = reg_0420;
    66: op1_13_in10 = reg_0208;
    67: op1_13_in10 = imem05_in[95:92];
    68: op1_13_in10 = imem07_in[39:36];
    69: op1_13_in10 = reg_0563;
    70: op1_13_in10 = imem05_in[19:16];
    71: op1_13_in10 = reg_0698;
    72: op1_13_in10 = reg_0141;
    73: op1_13_in10 = reg_0705;
    74: op1_13_in10 = reg_0811;
    75: op1_13_in10 = imem05_in[75:72];
    76: op1_13_in10 = reg_0162;
    77: op1_13_in10 = reg_0692;
    78: op1_13_in10 = reg_0612;
    79: op1_13_in10 = reg_0426;
    80: op1_13_in10 = reg_0810;
    81: op1_13_in10 = imem01_in[63:60];
    82: op1_13_in10 = reg_0142;
    83: op1_13_in10 = reg_0402;
    84: op1_13_in10 = reg_0531;
    85: op1_13_in10 = reg_0586;
    86: op1_13_in10 = reg_0170;
    87: op1_13_in10 = imem02_in[115:112];
    88: op1_13_in10 = reg_0434;
    89: op1_13_in10 = reg_0198;
    90: op1_13_in10 = reg_0463;
    91: op1_13_in10 = reg_0060;
    92: op1_13_in10 = reg_0765;
    93: op1_13_in10 = imem06_in[35:32];
    94: op1_13_in10 = reg_0538;
    95: op1_13_in10 = reg_0355;
    default: op1_13_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv10 = 1;
    8: op1_13_inv10 = 1;
    12: op1_13_inv10 = 1;
    13: op1_13_inv10 = 1;
    14: op1_13_inv10 = 1;
    15: op1_13_inv10 = 1;
    16: op1_13_inv10 = 1;
    17: op1_13_inv10 = 1;
    19: op1_13_inv10 = 1;
    20: op1_13_inv10 = 1;
    21: op1_13_inv10 = 1;
    22: op1_13_inv10 = 1;
    24: op1_13_inv10 = 1;
    25: op1_13_inv10 = 1;
    26: op1_13_inv10 = 1;
    27: op1_13_inv10 = 1;
    28: op1_13_inv10 = 1;
    29: op1_13_inv10 = 1;
    30: op1_13_inv10 = 1;
    32: op1_13_inv10 = 1;
    35: op1_13_inv10 = 1;
    36: op1_13_inv10 = 1;
    38: op1_13_inv10 = 1;
    40: op1_13_inv10 = 1;
    42: op1_13_inv10 = 1;
    45: op1_13_inv10 = 1;
    46: op1_13_inv10 = 1;
    50: op1_13_inv10 = 1;
    54: op1_13_inv10 = 1;
    55: op1_13_inv10 = 1;
    56: op1_13_inv10 = 1;
    57: op1_13_inv10 = 1;
    58: op1_13_inv10 = 1;
    59: op1_13_inv10 = 1;
    60: op1_13_inv10 = 1;
    66: op1_13_inv10 = 1;
    67: op1_13_inv10 = 1;
    70: op1_13_inv10 = 1;
    75: op1_13_inv10 = 1;
    76: op1_13_inv10 = 1;
    79: op1_13_inv10 = 1;
    82: op1_13_inv10 = 1;
    84: op1_13_inv10 = 1;
    85: op1_13_inv10 = 1;
    88: op1_13_inv10 = 1;
    90: op1_13_inv10 = 1;
    92: op1_13_inv10 = 1;
    93: op1_13_inv10 = 1;
    94: op1_13_inv10 = 1;
    default: op1_13_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in11 = reg_0351;
    5: op1_13_in11 = reg_0071;
    6: op1_13_in11 = reg_0201;
    7: op1_13_in11 = reg_0666;
    8: op1_13_in11 = reg_0408;
    9: op1_13_in11 = reg_0533;
    10: op1_13_in11 = reg_0680;
    11: op1_13_in11 = reg_0581;
    12: op1_13_in11 = reg_0480;
    13: op1_13_in11 = imem02_in[111:108];
    56: op1_13_in11 = imem02_in[111:108];
    14: op1_13_in11 = reg_0801;
    15: op1_13_in11 = reg_0816;
    16: op1_13_in11 = reg_0210;
    17: op1_13_in11 = reg_0708;
    18: op1_13_in11 = reg_0207;
    19: op1_13_in11 = reg_0176;
    20: op1_13_in11 = reg_0060;
    21: op1_13_in11 = imem04_in[119:116];
    22: op1_13_in11 = reg_0344;
    23: op1_13_in11 = reg_0787;
    61: op1_13_in11 = reg_0787;
    24: op1_13_in11 = imem07_in[31:28];
    25: op1_13_in11 = reg_0803;
    26: op1_13_in11 = reg_0694;
    27: op1_13_in11 = reg_0203;
    2: op1_13_in11 = reg_0185;
    52: op1_13_in11 = reg_0185;
    28: op1_13_in11 = reg_0271;
    29: op1_13_in11 = reg_0608;
    30: op1_13_in11 = imem02_in[95:92];
    31: op1_13_in11 = reg_0012;
    32: op1_13_in11 = reg_0059;
    33: op1_13_in11 = imem01_in[11:8];
    34: op1_13_in11 = imem02_in[39:36];
    35: op1_13_in11 = reg_0660;
    36: op1_13_in11 = reg_0056;
    37: op1_13_in11 = imem03_in[79:76];
    38: op1_13_in11 = reg_0238;
    39: op1_13_in11 = reg_0621;
    40: op1_13_in11 = reg_0711;
    41: op1_13_in11 = reg_0349;
    42: op1_13_in11 = reg_0297;
    43: op1_13_in11 = reg_0128;
    44: op1_13_in11 = reg_0459;
    45: op1_13_in11 = reg_0518;
    46: op1_13_in11 = reg_0129;
    47: op1_13_in11 = reg_0458;
    48: op1_13_in11 = reg_0655;
    49: op1_13_in11 = reg_0465;
    63: op1_13_in11 = reg_0465;
    77: op1_13_in11 = reg_0465;
    90: op1_13_in11 = reg_0465;
    50: op1_13_in11 = reg_0442;
    51: op1_13_in11 = reg_0091;
    86: op1_13_in11 = reg_0091;
    53: op1_13_in11 = reg_0814;
    54: op1_13_in11 = reg_0479;
    55: op1_13_in11 = reg_0671;
    57: op1_13_in11 = reg_0455;
    58: op1_13_in11 = reg_0807;
    59: op1_13_in11 = imem02_in[127:124];
    60: op1_13_in11 = reg_0810;
    62: op1_13_in11 = reg_0469;
    64: op1_13_in11 = reg_0468;
    65: op1_13_in11 = reg_0122;
    66: op1_13_in11 = reg_0204;
    67: op1_13_in11 = reg_0246;
    68: op1_13_in11 = reg_0719;
    69: op1_13_in11 = reg_0352;
    70: op1_13_in11 = imem05_in[55:52];
    71: op1_13_in11 = reg_0684;
    72: op1_13_in11 = reg_0138;
    73: op1_13_in11 = reg_0587;
    74: op1_13_in11 = reg_0001;
    75: op1_13_in11 = imem05_in[83:80];
    76: op1_13_in11 = reg_0169;
    78: op1_13_in11 = reg_0634;
    79: op1_13_in11 = reg_0485;
    80: op1_13_in11 = reg_0809;
    81: op1_13_in11 = imem01_in[71:68];
    82: op1_13_in11 = reg_0228;
    83: op1_13_in11 = reg_0519;
    84: op1_13_in11 = reg_0538;
    85: op1_13_in11 = reg_0360;
    87: op1_13_in11 = reg_0642;
    88: op1_13_in11 = reg_0267;
    89: op1_13_in11 = reg_0206;
    91: op1_13_in11 = reg_0558;
    92: op1_13_in11 = reg_0734;
    93: op1_13_in11 = imem06_in[75:72];
    94: op1_13_in11 = reg_0552;
    95: op1_13_in11 = reg_0144;
    default: op1_13_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv11 = 1;
    8: op1_13_inv11 = 1;
    11: op1_13_inv11 = 1;
    12: op1_13_inv11 = 1;
    14: op1_13_inv11 = 1;
    17: op1_13_inv11 = 1;
    18: op1_13_inv11 = 1;
    21: op1_13_inv11 = 1;
    23: op1_13_inv11 = 1;
    25: op1_13_inv11 = 1;
    26: op1_13_inv11 = 1;
    27: op1_13_inv11 = 1;
    2: op1_13_inv11 = 1;
    28: op1_13_inv11 = 1;
    33: op1_13_inv11 = 1;
    34: op1_13_inv11 = 1;
    36: op1_13_inv11 = 1;
    37: op1_13_inv11 = 1;
    38: op1_13_inv11 = 1;
    40: op1_13_inv11 = 1;
    41: op1_13_inv11 = 1;
    43: op1_13_inv11 = 1;
    44: op1_13_inv11 = 1;
    47: op1_13_inv11 = 1;
    49: op1_13_inv11 = 1;
    51: op1_13_inv11 = 1;
    52: op1_13_inv11 = 1;
    55: op1_13_inv11 = 1;
    58: op1_13_inv11 = 1;
    61: op1_13_inv11 = 1;
    62: op1_13_inv11 = 1;
    65: op1_13_inv11 = 1;
    66: op1_13_inv11 = 1;
    67: op1_13_inv11 = 1;
    73: op1_13_inv11 = 1;
    76: op1_13_inv11 = 1;
    77: op1_13_inv11 = 1;
    78: op1_13_inv11 = 1;
    80: op1_13_inv11 = 1;
    82: op1_13_inv11 = 1;
    83: op1_13_inv11 = 1;
    84: op1_13_inv11 = 1;
    85: op1_13_inv11 = 1;
    87: op1_13_inv11 = 1;
    88: op1_13_inv11 = 1;
    90: op1_13_inv11 = 1;
    93: op1_13_inv11 = 1;
    94: op1_13_inv11 = 1;
    default: op1_13_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in12 = reg_0382;
    5: op1_13_in12 = reg_0057;
    87: op1_13_in12 = reg_0057;
    6: op1_13_in12 = reg_0205;
    7: op1_13_in12 = reg_0641;
    8: op1_13_in12 = reg_0351;
    9: op1_13_in12 = reg_0294;
    10: op1_13_in12 = reg_0669;
    11: op1_13_in12 = reg_0360;
    12: op1_13_in12 = reg_0214;
    13: op1_13_in12 = imem02_in[123:120];
    56: op1_13_in12 = imem02_in[123:120];
    14: op1_13_in12 = reg_0015;
    74: op1_13_in12 = reg_0015;
    15: op1_13_in12 = reg_0037;
    16: op1_13_in12 = reg_0204;
    17: op1_13_in12 = reg_0718;
    18: op1_13_in12 = reg_0213;
    20: op1_13_in12 = reg_0083;
    21: op1_13_in12 = reg_0053;
    22: op1_13_in12 = reg_0381;
    23: op1_13_in12 = reg_0304;
    28: op1_13_in12 = reg_0304;
    51: op1_13_in12 = reg_0304;
    24: op1_13_in12 = imem07_in[59:56];
    25: op1_13_in12 = reg_0013;
    26: op1_13_in12 = reg_0676;
    27: op1_13_in12 = reg_0186;
    29: op1_13_in12 = reg_0618;
    30: op1_13_in12 = imem02_in[103:100];
    31: op1_13_in12 = reg_0807;
    32: op1_13_in12 = reg_0316;
    33: op1_13_in12 = imem01_in[15:12];
    34: op1_13_in12 = imem02_in[43:40];
    35: op1_13_in12 = reg_0657;
    36: op1_13_in12 = reg_0088;
    37: op1_13_in12 = imem03_in[99:96];
    38: op1_13_in12 = imem07_in[35:32];
    39: op1_13_in12 = reg_0368;
    40: op1_13_in12 = reg_0429;
    41: op1_13_in12 = reg_0344;
    42: op1_13_in12 = reg_0066;
    43: op1_13_in12 = reg_0152;
    44: op1_13_in12 = reg_0203;
    45: op1_13_in12 = reg_0531;
    46: op1_13_in12 = reg_0141;
    47: op1_13_in12 = reg_0189;
    48: op1_13_in12 = reg_0654;
    49: op1_13_in12 = reg_0475;
    57: op1_13_in12 = reg_0475;
    50: op1_13_in12 = reg_0084;
    52: op1_13_in12 = reg_0168;
    84: op1_13_in12 = reg_0168;
    53: op1_13_in12 = reg_0818;
    54: op1_13_in12 = reg_0459;
    55: op1_13_in12 = imem02_in[23:20];
    58: op1_13_in12 = reg_0507;
    59: op1_13_in12 = reg_0337;
    60: op1_13_in12 = reg_0010;
    61: op1_13_in12 = reg_0632;
    62: op1_13_in12 = reg_0474;
    63: op1_13_in12 = reg_0455;
    64: op1_13_in12 = reg_0458;
    65: op1_13_in12 = reg_0124;
    66: op1_13_in12 = reg_0194;
    67: op1_13_in12 = reg_0128;
    68: op1_13_in12 = reg_0725;
    69: op1_13_in12 = reg_0586;
    73: op1_13_in12 = reg_0586;
    70: op1_13_in12 = imem05_in[59:56];
    71: op1_13_in12 = reg_0749;
    72: op1_13_in12 = reg_0364;
    75: op1_13_in12 = imem05_in[123:120];
    76: op1_13_in12 = reg_0182;
    77: op1_13_in12 = reg_0454;
    90: op1_13_in12 = reg_0454;
    78: op1_13_in12 = reg_0453;
    79: op1_13_in12 = reg_0345;
    80: op1_13_in12 = imem04_in[11:8];
    81: op1_13_in12 = imem01_in[99:96];
    82: op1_13_in12 = reg_0325;
    83: op1_13_in12 = reg_0369;
    85: op1_13_in12 = reg_0342;
    88: op1_13_in12 = reg_0089;
    89: op1_13_in12 = reg_0199;
    91: op1_13_in12 = reg_0551;
    92: op1_13_in12 = imem06_in[3:0];
    93: op1_13_in12 = imem06_in[83:80];
    94: op1_13_in12 = reg_0500;
    95: op1_13_in12 = reg_0489;
    default: op1_13_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv12 = 1;
    9: op1_13_inv12 = 1;
    10: op1_13_inv12 = 1;
    11: op1_13_inv12 = 1;
    12: op1_13_inv12 = 1;
    14: op1_13_inv12 = 1;
    15: op1_13_inv12 = 1;
    20: op1_13_inv12 = 1;
    21: op1_13_inv12 = 1;
    24: op1_13_inv12 = 1;
    25: op1_13_inv12 = 1;
    27: op1_13_inv12 = 1;
    28: op1_13_inv12 = 1;
    30: op1_13_inv12 = 1;
    34: op1_13_inv12 = 1;
    35: op1_13_inv12 = 1;
    36: op1_13_inv12 = 1;
    37: op1_13_inv12 = 1;
    39: op1_13_inv12 = 1;
    40: op1_13_inv12 = 1;
    47: op1_13_inv12 = 1;
    48: op1_13_inv12 = 1;
    49: op1_13_inv12 = 1;
    50: op1_13_inv12 = 1;
    52: op1_13_inv12 = 1;
    55: op1_13_inv12 = 1;
    57: op1_13_inv12 = 1;
    60: op1_13_inv12 = 1;
    61: op1_13_inv12 = 1;
    62: op1_13_inv12 = 1;
    64: op1_13_inv12 = 1;
    66: op1_13_inv12 = 1;
    67: op1_13_inv12 = 1;
    69: op1_13_inv12 = 1;
    71: op1_13_inv12 = 1;
    72: op1_13_inv12 = 1;
    73: op1_13_inv12 = 1;
    74: op1_13_inv12 = 1;
    81: op1_13_inv12 = 1;
    82: op1_13_inv12 = 1;
    84: op1_13_inv12 = 1;
    85: op1_13_inv12 = 1;
    87: op1_13_inv12 = 1;
    88: op1_13_inv12 = 1;
    89: op1_13_inv12 = 1;
    92: op1_13_inv12 = 1;
    94: op1_13_inv12 = 1;
    default: op1_13_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in13 = reg_0383;
    5: op1_13_in13 = reg_0072;
    6: op1_13_in13 = imem01_in[99:96];
    7: op1_13_in13 = reg_0665;
    8: op1_13_in13 = reg_0409;
    9: op1_13_in13 = reg_0297;
    10: op1_13_in13 = reg_0457;
    11: op1_13_in13 = reg_0317;
    12: op1_13_in13 = reg_0194;
    47: op1_13_in13 = reg_0194;
    13: op1_13_in13 = imem02_in[127:124];
    14: op1_13_in13 = reg_0810;
    15: op1_13_in13 = imem07_in[19:16];
    16: op1_13_in13 = reg_0198;
    17: op1_13_in13 = reg_0727;
    18: op1_13_in13 = reg_0196;
    20: op1_13_in13 = reg_0655;
    21: op1_13_in13 = reg_0283;
    91: op1_13_in13 = reg_0283;
    22: op1_13_in13 = reg_0408;
    23: op1_13_in13 = reg_0309;
    28: op1_13_in13 = reg_0309;
    24: op1_13_in13 = imem07_in[71:68];
    25: op1_13_in13 = reg_0007;
    26: op1_13_in13 = reg_0686;
    27: op1_13_in13 = reg_0195;
    29: op1_13_in13 = reg_0622;
    30: op1_13_in13 = reg_0666;
    31: op1_13_in13 = reg_0802;
    32: op1_13_in13 = reg_0536;
    33: op1_13_in13 = imem01_in[31:28];
    34: op1_13_in13 = imem02_in[123:120];
    35: op1_13_in13 = reg_0661;
    36: op1_13_in13 = reg_0555;
    37: op1_13_in13 = imem03_in[119:116];
    38: op1_13_in13 = imem07_in[103:100];
    39: op1_13_in13 = reg_0231;
    40: op1_13_in13 = reg_0448;
    41: op1_13_in13 = reg_0320;
    42: op1_13_in13 = reg_0254;
    43: op1_13_in13 = reg_0142;
    44: op1_13_in13 = reg_0211;
    45: op1_13_in13 = imem03_in[87:84];
    46: op1_13_in13 = imem06_in[3:0];
    48: op1_13_in13 = reg_0660;
    49: op1_13_in13 = reg_0480;
    50: op1_13_in13 = reg_0267;
    51: op1_13_in13 = reg_0070;
    53: op1_13_in13 = imem07_in[23:20];
    54: op1_13_in13 = reg_0193;
    55: op1_13_in13 = imem02_in[43:40];
    56: op1_13_in13 = reg_0650;
    57: op1_13_in13 = reg_0468;
    58: op1_13_in13 = reg_0403;
    59: op1_13_in13 = reg_0584;
    60: op1_13_in13 = imem04_in[19:16];
    61: op1_13_in13 = imem07_in[39:36];
    62: op1_13_in13 = reg_0214;
    63: op1_13_in13 = reg_0477;
    90: op1_13_in13 = reg_0477;
    64: op1_13_in13 = reg_0204;
    65: op1_13_in13 = reg_0672;
    66: op1_13_in13 = reg_0206;
    67: op1_13_in13 = reg_0789;
    68: op1_13_in13 = reg_0718;
    69: op1_13_in13 = reg_0345;
    70: op1_13_in13 = reg_0391;
    71: op1_13_in13 = reg_0634;
    72: op1_13_in13 = reg_0359;
    73: op1_13_in13 = reg_0361;
    74: op1_13_in13 = reg_0799;
    75: op1_13_in13 = reg_0337;
    76: op1_13_in13 = reg_0164;
    77: op1_13_in13 = reg_0451;
    78: op1_13_in13 = reg_0455;
    79: op1_13_in13 = reg_0565;
    80: op1_13_in13 = imem04_in[51:48];
    81: op1_13_in13 = imem01_in[107:104];
    82: op1_13_in13 = reg_0091;
    83: op1_13_in13 = reg_0816;
    84: op1_13_in13 = reg_0639;
    85: op1_13_in13 = reg_0406;
    87: op1_13_in13 = reg_0656;
    88: op1_13_in13 = reg_0730;
    89: op1_13_in13 = imem01_in[19:16];
    92: op1_13_in13 = reg_0291;
    93: op1_13_in13 = imem06_in[103:100];
    94: op1_13_in13 = reg_0492;
    95: op1_13_in13 = reg_0797;
    default: op1_13_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv13 = 1;
    6: op1_13_inv13 = 1;
    7: op1_13_inv13 = 1;
    11: op1_13_inv13 = 1;
    12: op1_13_inv13 = 1;
    14: op1_13_inv13 = 1;
    15: op1_13_inv13 = 1;
    16: op1_13_inv13 = 1;
    18: op1_13_inv13 = 1;
    20: op1_13_inv13 = 1;
    22: op1_13_inv13 = 1;
    23: op1_13_inv13 = 1;
    25: op1_13_inv13 = 1;
    26: op1_13_inv13 = 1;
    27: op1_13_inv13 = 1;
    30: op1_13_inv13 = 1;
    31: op1_13_inv13 = 1;
    35: op1_13_inv13 = 1;
    37: op1_13_inv13 = 1;
    41: op1_13_inv13 = 1;
    45: op1_13_inv13 = 1;
    47: op1_13_inv13 = 1;
    49: op1_13_inv13 = 1;
    50: op1_13_inv13 = 1;
    53: op1_13_inv13 = 1;
    55: op1_13_inv13 = 1;
    58: op1_13_inv13 = 1;
    59: op1_13_inv13 = 1;
    60: op1_13_inv13 = 1;
    61: op1_13_inv13 = 1;
    64: op1_13_inv13 = 1;
    69: op1_13_inv13 = 1;
    70: op1_13_inv13 = 1;
    72: op1_13_inv13 = 1;
    77: op1_13_inv13 = 1;
    78: op1_13_inv13 = 1;
    83: op1_13_inv13 = 1;
    87: op1_13_inv13 = 1;
    89: op1_13_inv13 = 1;
    91: op1_13_inv13 = 1;
    93: op1_13_inv13 = 1;
    95: op1_13_inv13 = 1;
    default: op1_13_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in14 = reg_0315;
    5: op1_13_in14 = reg_0749;
    6: op1_13_in14 = reg_0523;
    7: op1_13_in14 = reg_0652;
    8: op1_13_in14 = reg_0401;
    9: op1_13_in14 = reg_0047;
    10: op1_13_in14 = reg_0459;
    11: op1_13_in14 = reg_0327;
    12: op1_13_in14 = imem01_in[55:52];
    13: op1_13_in14 = reg_0654;
    14: op1_13_in14 = reg_0809;
    15: op1_13_in14 = imem07_in[43:40];
    16: op1_13_in14 = reg_0212;
    17: op1_13_in14 = reg_0425;
    18: op1_13_in14 = reg_0195;
    20: op1_13_in14 = reg_0651;
    21: op1_13_in14 = reg_0529;
    22: op1_13_in14 = reg_0406;
    23: op1_13_in14 = reg_0735;
    28: op1_13_in14 = reg_0735;
    24: op1_13_in14 = imem07_in[79:76];
    25: op1_13_in14 = reg_0804;
    26: op1_13_in14 = reg_0670;
    27: op1_13_in14 = imem01_in[11:8];
    29: op1_13_in14 = reg_0623;
    30: op1_13_in14 = reg_0660;
    31: op1_13_in14 = reg_0015;
    32: op1_13_in14 = reg_0510;
    33: op1_13_in14 = imem01_in[35:32];
    34: op1_13_in14 = reg_0657;
    35: op1_13_in14 = reg_0662;
    36: op1_13_in14 = reg_0536;
    37: op1_13_in14 = reg_0587;
    38: op1_13_in14 = imem07_in[119:116];
    39: op1_13_in14 = reg_0029;
    40: op1_13_in14 = reg_0169;
    41: op1_13_in14 = reg_0342;
    42: op1_13_in14 = reg_0068;
    43: op1_13_in14 = reg_0134;
    44: op1_13_in14 = reg_0186;
    45: op1_13_in14 = reg_0580;
    94: op1_13_in14 = reg_0580;
    46: op1_13_in14 = imem06_in[27:24];
    47: op1_13_in14 = reg_0192;
    66: op1_13_in14 = reg_0192;
    48: op1_13_in14 = reg_0346;
    49: op1_13_in14 = reg_0473;
    50: op1_13_in14 = reg_0164;
    51: op1_13_in14 = reg_0102;
    53: op1_13_in14 = imem07_in[39:36];
    54: op1_13_in14 = reg_0201;
    55: op1_13_in14 = imem02_in[91:88];
    56: op1_13_in14 = reg_0337;
    57: op1_13_in14 = reg_0452;
    58: op1_13_in14 = reg_0262;
    59: op1_13_in14 = reg_0639;
    60: op1_13_in14 = imem04_in[23:20];
    61: op1_13_in14 = imem07_in[67:64];
    62: op1_13_in14 = reg_0200;
    63: op1_13_in14 = reg_0472;
    64: op1_13_in14 = reg_0188;
    65: op1_13_in14 = reg_0671;
    67: op1_13_in14 = reg_0278;
    68: op1_13_in14 = reg_0067;
    69: op1_13_in14 = reg_0361;
    72: op1_13_in14 = reg_0361;
    79: op1_13_in14 = reg_0361;
    70: op1_13_in14 = reg_0487;
    71: op1_13_in14 = reg_0451;
    73: op1_13_in14 = reg_0351;
    74: op1_13_in14 = imem04_in[15:12];
    75: op1_13_in14 = reg_0667;
    76: op1_13_in14 = reg_0170;
    77: op1_13_in14 = reg_0461;
    78: op1_13_in14 = reg_0477;
    80: op1_13_in14 = imem04_in[71:68];
    81: op1_13_in14 = reg_0085;
    82: op1_13_in14 = reg_0176;
    83: op1_13_in14 = reg_0748;
    84: op1_13_in14 = reg_0322;
    85: op1_13_in14 = reg_0281;
    87: op1_13_in14 = reg_0304;
    88: op1_13_in14 = reg_0110;
    89: op1_13_in14 = imem01_in[75:72];
    90: op1_13_in14 = reg_0476;
    91: op1_13_in14 = reg_0071;
    92: op1_13_in14 = reg_0354;
    93: op1_13_in14 = imem06_in[111:108];
    95: op1_13_in14 = reg_0583;
    default: op1_13_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv14 = 1;
    9: op1_13_inv14 = 1;
    11: op1_13_inv14 = 1;
    12: op1_13_inv14 = 1;
    15: op1_13_inv14 = 1;
    16: op1_13_inv14 = 1;
    17: op1_13_inv14 = 1;
    18: op1_13_inv14 = 1;
    23: op1_13_inv14 = 1;
    24: op1_13_inv14 = 1;
    26: op1_13_inv14 = 1;
    27: op1_13_inv14 = 1;
    36: op1_13_inv14 = 1;
    38: op1_13_inv14 = 1;
    41: op1_13_inv14 = 1;
    42: op1_13_inv14 = 1;
    45: op1_13_inv14 = 1;
    46: op1_13_inv14 = 1;
    47: op1_13_inv14 = 1;
    49: op1_13_inv14 = 1;
    53: op1_13_inv14 = 1;
    56: op1_13_inv14 = 1;
    61: op1_13_inv14 = 1;
    63: op1_13_inv14 = 1;
    66: op1_13_inv14 = 1;
    72: op1_13_inv14 = 1;
    74: op1_13_inv14 = 1;
    79: op1_13_inv14 = 1;
    81: op1_13_inv14 = 1;
    82: op1_13_inv14 = 1;
    85: op1_13_inv14 = 1;
    89: op1_13_inv14 = 1;
    90: op1_13_inv14 = 1;
    91: op1_13_inv14 = 1;
    93: op1_13_inv14 = 1;
    default: op1_13_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in15 = reg_0367;
    39: op1_13_in15 = reg_0367;
    5: op1_13_in15 = reg_0736;
    6: op1_13_in15 = reg_0501;
    7: op1_13_in15 = reg_0320;
    8: op1_13_in15 = imem06_in[7:4];
    9: op1_13_in15 = reg_0066;
    10: op1_13_in15 = reg_0186;
    11: op1_13_in15 = reg_0312;
    12: op1_13_in15 = imem01_in[63:60];
    13: op1_13_in15 = reg_0661;
    14: op1_13_in15 = imem04_in[43:40];
    74: op1_13_in15 = imem04_in[43:40];
    15: op1_13_in15 = imem07_in[47:44];
    16: op1_13_in15 = reg_0190;
    17: op1_13_in15 = reg_0441;
    18: op1_13_in15 = reg_0197;
    20: op1_13_in15 = reg_0640;
    21: op1_13_in15 = reg_0302;
    22: op1_13_in15 = reg_0028;
    23: op1_13_in15 = reg_0272;
    24: op1_13_in15 = imem07_in[107:104];
    25: op1_13_in15 = reg_0806;
    26: op1_13_in15 = reg_0679;
    27: op1_13_in15 = imem01_in[27:24];
    28: op1_13_in15 = reg_0527;
    29: op1_13_in15 = reg_0615;
    30: op1_13_in15 = reg_0656;
    31: op1_13_in15 = reg_0016;
    32: op1_13_in15 = reg_0556;
    33: op1_13_in15 = imem01_in[71:68];
    34: op1_13_in15 = reg_0662;
    35: op1_13_in15 = reg_0667;
    36: op1_13_in15 = reg_0551;
    37: op1_13_in15 = reg_0596;
    38: op1_13_in15 = imem07_in[123:120];
    40: op1_13_in15 = reg_0183;
    41: op1_13_in15 = reg_0350;
    42: op1_13_in15 = reg_0070;
    43: op1_13_in15 = reg_0144;
    44: op1_13_in15 = reg_0198;
    45: op1_13_in15 = reg_0578;
    46: op1_13_in15 = imem06_in[39:36];
    47: op1_13_in15 = reg_0085;
    48: op1_13_in15 = reg_0638;
    49: op1_13_in15 = reg_0470;
    63: op1_13_in15 = reg_0470;
    50: op1_13_in15 = reg_0168;
    51: op1_13_in15 = reg_0285;
    53: op1_13_in15 = imem07_in[51:48];
    54: op1_13_in15 = reg_0205;
    55: op1_13_in15 = imem02_in[119:116];
    56: op1_13_in15 = reg_0666;
    57: op1_13_in15 = reg_0458;
    58: op1_13_in15 = reg_0315;
    59: op1_13_in15 = reg_0427;
    60: op1_13_in15 = imem04_in[55:52];
    61: op1_13_in15 = imem07_in[83:80];
    62: op1_13_in15 = reg_0210;
    64: op1_13_in15 = reg_0207;
    65: op1_13_in15 = reg_0127;
    66: op1_13_in15 = imem01_in[15:12];
    67: op1_13_in15 = reg_0786;
    68: op1_13_in15 = reg_0635;
    69: op1_13_in15 = reg_0342;
    70: op1_13_in15 = reg_0374;
    71: op1_13_in15 = reg_0455;
    72: op1_13_in15 = reg_0363;
    73: op1_13_in15 = reg_0365;
    75: op1_13_in15 = reg_0133;
    77: op1_13_in15 = reg_0466;
    90: op1_13_in15 = reg_0466;
    78: op1_13_in15 = reg_0469;
    79: op1_13_in15 = reg_0360;
    80: op1_13_in15 = imem04_in[75:72];
    81: op1_13_in15 = reg_0497;
    83: op1_13_in15 = reg_0270;
    84: op1_13_in15 = reg_0059;
    85: op1_13_in15 = reg_0132;
    87: op1_13_in15 = reg_0587;
    88: op1_13_in15 = reg_0236;
    89: op1_13_in15 = imem01_in[83:80];
    91: op1_13_in15 = reg_0598;
    92: op1_13_in15 = reg_0038;
    93: op1_13_in15 = reg_0348;
    94: op1_13_in15 = reg_0751;
    95: op1_13_in15 = reg_0288;
    default: op1_13_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv15 = 1;
    6: op1_13_inv15 = 1;
    10: op1_13_inv15 = 1;
    11: op1_13_inv15 = 1;
    12: op1_13_inv15 = 1;
    14: op1_13_inv15 = 1;
    15: op1_13_inv15 = 1;
    17: op1_13_inv15 = 1;
    18: op1_13_inv15 = 1;
    23: op1_13_inv15 = 1;
    25: op1_13_inv15 = 1;
    26: op1_13_inv15 = 1;
    27: op1_13_inv15 = 1;
    28: op1_13_inv15 = 1;
    29: op1_13_inv15 = 1;
    30: op1_13_inv15 = 1;
    34: op1_13_inv15 = 1;
    35: op1_13_inv15 = 1;
    36: op1_13_inv15 = 1;
    37: op1_13_inv15 = 1;
    40: op1_13_inv15 = 1;
    43: op1_13_inv15 = 1;
    44: op1_13_inv15 = 1;
    45: op1_13_inv15 = 1;
    46: op1_13_inv15 = 1;
    48: op1_13_inv15 = 1;
    49: op1_13_inv15 = 1;
    50: op1_13_inv15 = 1;
    53: op1_13_inv15 = 1;
    54: op1_13_inv15 = 1;
    58: op1_13_inv15 = 1;
    60: op1_13_inv15 = 1;
    62: op1_13_inv15 = 1;
    64: op1_13_inv15 = 1;
    65: op1_13_inv15 = 1;
    66: op1_13_inv15 = 1;
    67: op1_13_inv15 = 1;
    70: op1_13_inv15 = 1;
    72: op1_13_inv15 = 1;
    73: op1_13_inv15 = 1;
    74: op1_13_inv15 = 1;
    75: op1_13_inv15 = 1;
    81: op1_13_inv15 = 1;
    84: op1_13_inv15 = 1;
    85: op1_13_inv15 = 1;
    93: op1_13_inv15 = 1;
    default: op1_13_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in16 = reg_0368;
    5: op1_13_in16 = reg_0750;
    6: op1_13_in16 = reg_0502;
    7: op1_13_in16 = reg_0330;
    8: op1_13_in16 = imem06_in[19:16];
    9: op1_13_in16 = reg_0076;
    10: op1_13_in16 = reg_0196;
    11: op1_13_in16 = reg_0397;
    12: op1_13_in16 = imem01_in[119:116];
    13: op1_13_in16 = reg_0665;
    14: op1_13_in16 = imem04_in[47:44];
    15: op1_13_in16 = imem07_in[75:72];
    16: op1_13_in16 = reg_0199;
    17: op1_13_in16 = reg_0428;
    18: op1_13_in16 = imem01_in[3:0];
    20: op1_13_in16 = reg_0334;
    21: op1_13_in16 = reg_0292;
    22: op1_13_in16 = reg_0032;
    23: op1_13_in16 = reg_0734;
    24: op1_13_in16 = imem07_in[119:116];
    25: op1_13_in16 = reg_0810;
    26: op1_13_in16 = reg_0678;
    27: op1_13_in16 = imem01_in[63:60];
    28: op1_13_in16 = reg_0260;
    29: op1_13_in16 = reg_0408;
    30: op1_13_in16 = reg_0638;
    31: op1_13_in16 = reg_0806;
    32: op1_13_in16 = reg_0303;
    33: op1_13_in16 = reg_0336;
    34: op1_13_in16 = reg_0643;
    35: op1_13_in16 = reg_0344;
    36: op1_13_in16 = reg_0308;
    37: op1_13_in16 = reg_0592;
    38: op1_13_in16 = reg_0714;
    39: op1_13_in16 = imem07_in[3:0];
    40: op1_13_in16 = reg_0177;
    41: op1_13_in16 = reg_0518;
    42: op1_13_in16 = imem05_in[3:0];
    43: op1_13_in16 = imem06_in[3:0];
    44: op1_13_in16 = reg_0190;
    45: op1_13_in16 = reg_0590;
    46: op1_13_in16 = imem06_in[43:40];
    47: op1_13_in16 = reg_0233;
    48: op1_13_in16 = reg_0667;
    49: op1_13_in16 = reg_0471;
    50: op1_13_in16 = reg_0178;
    51: op1_13_in16 = reg_0148;
    53: op1_13_in16 = imem07_in[79:76];
    54: op1_13_in16 = imem01_in[35:32];
    55: op1_13_in16 = reg_0637;
    56: op1_13_in16 = reg_0637;
    57: op1_13_in16 = reg_0187;
    62: op1_13_in16 = reg_0187;
    58: op1_13_in16 = reg_0552;
    59: op1_13_in16 = reg_0352;
    60: op1_13_in16 = imem04_in[59:56];
    61: op1_13_in16 = imem07_in[103:100];
    63: op1_13_in16 = reg_0459;
    64: op1_13_in16 = reg_0186;
    65: op1_13_in16 = imem02_in[15:12];
    66: op1_13_in16 = imem01_in[79:76];
    67: op1_13_in16 = reg_0486;
    68: op1_13_in16 = reg_0333;
    69: op1_13_in16 = reg_0414;
    70: op1_13_in16 = reg_0517;
    71: op1_13_in16 = reg_0191;
    72: op1_13_in16 = reg_0353;
    73: op1_13_in16 = reg_0743;
    74: op1_13_in16 = imem04_in[91:88];
    75: op1_13_in16 = reg_0795;
    77: op1_13_in16 = reg_0452;
    78: op1_13_in16 = reg_0480;
    90: op1_13_in16 = reg_0480;
    79: op1_13_in16 = reg_0342;
    80: op1_13_in16 = imem04_in[79:76];
    81: op1_13_in16 = reg_0772;
    83: op1_13_in16 = reg_0764;
    84: op1_13_in16 = reg_0361;
    85: op1_13_in16 = reg_0540;
    87: op1_13_in16 = reg_0345;
    88: op1_13_in16 = reg_0182;
    89: op1_13_in16 = imem01_in[87:84];
    91: op1_13_in16 = reg_0371;
    92: op1_13_in16 = reg_0265;
    93: op1_13_in16 = reg_0578;
    94: op1_13_in16 = reg_0288;
    95: op1_13_in16 = reg_0393;
    default: op1_13_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv16 = 1;
    5: op1_13_inv16 = 1;
    9: op1_13_inv16 = 1;
    13: op1_13_inv16 = 1;
    15: op1_13_inv16 = 1;
    16: op1_13_inv16 = 1;
    17: op1_13_inv16 = 1;
    18: op1_13_inv16 = 1;
    20: op1_13_inv16 = 1;
    23: op1_13_inv16 = 1;
    24: op1_13_inv16 = 1;
    25: op1_13_inv16 = 1;
    26: op1_13_inv16 = 1;
    29: op1_13_inv16 = 1;
    30: op1_13_inv16 = 1;
    32: op1_13_inv16 = 1;
    33: op1_13_inv16 = 1;
    36: op1_13_inv16 = 1;
    40: op1_13_inv16 = 1;
    41: op1_13_inv16 = 1;
    42: op1_13_inv16 = 1;
    43: op1_13_inv16 = 1;
    44: op1_13_inv16 = 1;
    47: op1_13_inv16 = 1;
    51: op1_13_inv16 = 1;
    55: op1_13_inv16 = 1;
    56: op1_13_inv16 = 1;
    58: op1_13_inv16 = 1;
    60: op1_13_inv16 = 1;
    63: op1_13_inv16 = 1;
    66: op1_13_inv16 = 1;
    67: op1_13_inv16 = 1;
    68: op1_13_inv16 = 1;
    70: op1_13_inv16 = 1;
    71: op1_13_inv16 = 1;
    79: op1_13_inv16 = 1;
    84: op1_13_inv16 = 1;
    85: op1_13_inv16 = 1;
    87: op1_13_inv16 = 1;
    92: op1_13_inv16 = 1;
    94: op1_13_inv16 = 1;
    default: op1_13_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in17 = reg_0031;
    5: op1_13_in17 = reg_0751;
    6: op1_13_in17 = reg_0515;
    7: op1_13_in17 = reg_0353;
    8: op1_13_in17 = imem06_in[23:20];
    9: op1_13_in17 = reg_0067;
    10: op1_13_in17 = reg_0197;
    11: op1_13_in17 = reg_0361;
    87: op1_13_in17 = reg_0361;
    12: op1_13_in17 = imem01_in[123:120];
    13: op1_13_in17 = reg_0333;
    14: op1_13_in17 = imem04_in[59:56];
    15: op1_13_in17 = imem07_in[107:104];
    16: op1_13_in17 = imem01_in[71:68];
    17: op1_13_in17 = reg_0175;
    18: op1_13_in17 = imem01_in[11:8];
    64: op1_13_in17 = imem01_in[11:8];
    20: op1_13_in17 = reg_0341;
    21: op1_13_in17 = reg_0061;
    22: op1_13_in17 = reg_0040;
    23: op1_13_in17 = reg_0285;
    24: op1_13_in17 = imem07_in[123:120];
    25: op1_13_in17 = reg_0809;
    26: op1_13_in17 = reg_0687;
    27: op1_13_in17 = imem01_in[83:80];
    28: op1_13_in17 = reg_0272;
    29: op1_13_in17 = reg_0762;
    30: op1_13_in17 = reg_0663;
    31: op1_13_in17 = reg_0004;
    32: op1_13_in17 = reg_0308;
    33: op1_13_in17 = reg_0501;
    34: op1_13_in17 = reg_0363;
    35: op1_13_in17 = reg_0343;
    36: op1_13_in17 = reg_0273;
    37: op1_13_in17 = reg_0591;
    38: op1_13_in17 = reg_0715;
    39: op1_13_in17 = imem07_in[87:84];
    53: op1_13_in17 = imem07_in[87:84];
    40: op1_13_in17 = reg_0185;
    41: op1_13_in17 = reg_0092;
    79: op1_13_in17 = reg_0092;
    42: op1_13_in17 = imem05_in[51:48];
    43: op1_13_in17 = imem06_in[123:120];
    44: op1_13_in17 = reg_0195;
    45: op1_13_in17 = reg_0749;
    46: op1_13_in17 = imem06_in[55:52];
    47: op1_13_in17 = reg_0227;
    48: op1_13_in17 = reg_0336;
    89: op1_13_in17 = reg_0336;
    49: op1_13_in17 = reg_0200;
    63: op1_13_in17 = reg_0200;
    50: op1_13_in17 = reg_0173;
    51: op1_13_in17 = reg_0151;
    54: op1_13_in17 = imem01_in[59:56];
    55: op1_13_in17 = reg_0346;
    56: op1_13_in17 = reg_0584;
    57: op1_13_in17 = reg_0193;
    58: op1_13_in17 = reg_0056;
    59: op1_13_in17 = reg_0344;
    60: op1_13_in17 = imem04_in[63:60];
    61: op1_13_in17 = imem07_in[115:112];
    62: op1_13_in17 = reg_0204;
    71: op1_13_in17 = reg_0204;
    65: op1_13_in17 = imem02_in[91:88];
    66: op1_13_in17 = imem01_in[91:88];
    67: op1_13_in17 = reg_0145;
    68: op1_13_in17 = reg_0442;
    69: op1_13_in17 = reg_0323;
    70: op1_13_in17 = reg_0075;
    72: op1_13_in17 = reg_0342;
    73: op1_13_in17 = reg_0080;
    74: op1_13_in17 = imem04_in[111:108];
    75: op1_13_in17 = reg_0732;
    77: op1_13_in17 = reg_0458;
    78: op1_13_in17 = reg_0468;
    80: op1_13_in17 = reg_0043;
    81: op1_13_in17 = reg_0520;
    83: op1_13_in17 = reg_0700;
    84: op1_13_in17 = reg_0365;
    85: op1_13_in17 = reg_0526;
    88: op1_13_in17 = reg_0100;
    90: op1_13_in17 = reg_0473;
    91: op1_13_in17 = imem05_in[23:20];
    92: op1_13_in17 = reg_0628;
    93: op1_13_in17 = reg_0408;
    94: op1_13_in17 = reg_0393;
    95: op1_13_in17 = reg_0579;
    default: op1_13_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv17 = 1;
    5: op1_13_inv17 = 1;
    6: op1_13_inv17 = 1;
    9: op1_13_inv17 = 1;
    11: op1_13_inv17 = 1;
    12: op1_13_inv17 = 1;
    13: op1_13_inv17 = 1;
    15: op1_13_inv17 = 1;
    17: op1_13_inv17 = 1;
    18: op1_13_inv17 = 1;
    20: op1_13_inv17 = 1;
    21: op1_13_inv17 = 1;
    23: op1_13_inv17 = 1;
    24: op1_13_inv17 = 1;
    25: op1_13_inv17 = 1;
    26: op1_13_inv17 = 1;
    27: op1_13_inv17 = 1;
    29: op1_13_inv17 = 1;
    31: op1_13_inv17 = 1;
    32: op1_13_inv17 = 1;
    33: op1_13_inv17 = 1;
    34: op1_13_inv17 = 1;
    35: op1_13_inv17 = 1;
    37: op1_13_inv17 = 1;
    38: op1_13_inv17 = 1;
    39: op1_13_inv17 = 1;
    40: op1_13_inv17 = 1;
    43: op1_13_inv17 = 1;
    44: op1_13_inv17 = 1;
    45: op1_13_inv17 = 1;
    47: op1_13_inv17 = 1;
    54: op1_13_inv17 = 1;
    55: op1_13_inv17 = 1;
    56: op1_13_inv17 = 1;
    61: op1_13_inv17 = 1;
    62: op1_13_inv17 = 1;
    63: op1_13_inv17 = 1;
    68: op1_13_inv17 = 1;
    70: op1_13_inv17 = 1;
    71: op1_13_inv17 = 1;
    74: op1_13_inv17 = 1;
    78: op1_13_inv17 = 1;
    79: op1_13_inv17 = 1;
    87: op1_13_inv17 = 1;
    90: op1_13_inv17 = 1;
    93: op1_13_inv17 = 1;
    94: op1_13_inv17 = 1;
    default: op1_13_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in18 = reg_0032;
    5: op1_13_in18 = reg_0752;
    6: op1_13_in18 = reg_0505;
    7: op1_13_in18 = reg_0310;
    8: op1_13_in18 = imem06_in[71:68];
    9: op1_13_in18 = imem05_in[51:48];
    10: op1_13_in18 = reg_0739;
    11: op1_13_in18 = reg_0309;
    12: op1_13_in18 = reg_0501;
    13: op1_13_in18 = reg_0364;
    14: op1_13_in18 = imem04_in[71:68];
    15: op1_13_in18 = reg_0731;
    16: op1_13_in18 = imem01_in[75:72];
    17: op1_13_in18 = reg_0161;
    68: op1_13_in18 = reg_0161;
    18: op1_13_in18 = imem01_in[31:28];
    20: op1_13_in18 = reg_0359;
    21: op1_13_in18 = reg_0065;
    22: op1_13_in18 = reg_0814;
    23: op1_13_in18 = reg_0132;
    24: op1_13_in18 = reg_0719;
    25: op1_13_in18 = imem04_in[7:4];
    26: op1_13_in18 = reg_0669;
    27: op1_13_in18 = imem01_in[115:112];
    28: op1_13_in18 = reg_0744;
    29: op1_13_in18 = reg_0403;
    30: op1_13_in18 = reg_0358;
    31: op1_13_in18 = imem04_in[11:8];
    32: op1_13_in18 = reg_0291;
    33: op1_13_in18 = reg_0487;
    34: op1_13_in18 = reg_0360;
    35: op1_13_in18 = reg_0092;
    36: op1_13_in18 = reg_0290;
    37: op1_13_in18 = reg_0600;
    38: op1_13_in18 = reg_0436;
    39: op1_13_in18 = imem07_in[111:108];
    53: op1_13_in18 = imem07_in[111:108];
    40: op1_13_in18 = reg_0157;
    41: op1_13_in18 = reg_0769;
    42: op1_13_in18 = imem05_in[63:60];
    43: op1_13_in18 = reg_0218;
    44: op1_13_in18 = reg_0197;
    45: op1_13_in18 = reg_0394;
    46: op1_13_in18 = imem06_in[75:72];
    47: op1_13_in18 = imem01_in[3:0];
    48: op1_13_in18 = reg_0352;
    49: op1_13_in18 = reg_0193;
    51: op1_13_in18 = reg_0138;
    54: op1_13_in18 = imem01_in[71:68];
    55: op1_13_in18 = reg_0548;
    56: op1_13_in18 = reg_0657;
    57: op1_13_in18 = reg_0205;
    58: op1_13_in18 = reg_0055;
    59: op1_13_in18 = reg_0320;
    60: op1_13_in18 = imem04_in[67:64];
    61: op1_13_in18 = imem07_in[127:124];
    62: op1_13_in18 = reg_0186;
    71: op1_13_in18 = reg_0186;
    63: op1_13_in18 = reg_0208;
    77: op1_13_in18 = reg_0208;
    64: op1_13_in18 = imem01_in[63:60];
    65: op1_13_in18 = imem02_in[127:124];
    66: op1_13_in18 = imem01_in[111:108];
    67: op1_13_in18 = reg_0130;
    69: op1_13_in18 = reg_0743;
    70: op1_13_in18 = reg_0229;
    72: op1_13_in18 = reg_0414;
    73: op1_13_in18 = reg_0757;
    74: op1_13_in18 = reg_0059;
    75: op1_13_in18 = reg_0489;
    78: op1_13_in18 = reg_0191;
    79: op1_13_in18 = reg_0541;
    80: op1_13_in18 = reg_0060;
    81: op1_13_in18 = reg_0385;
    83: op1_13_in18 = reg_0651;
    84: op1_13_in18 = reg_0342;
    85: op1_13_in18 = reg_0093;
    87: op1_13_in18 = reg_0343;
    88: op1_13_in18 = reg_0170;
    89: op1_13_in18 = reg_0741;
    90: op1_13_in18 = reg_0467;
    91: op1_13_in18 = imem05_in[35:32];
    92: op1_13_in18 = reg_0578;
    93: op1_13_in18 = reg_0307;
    94: op1_13_in18 = reg_0277;
    95: op1_13_in18 = reg_0547;
    default: op1_13_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv18 = 1;
    6: op1_13_inv18 = 1;
    7: op1_13_inv18 = 1;
    8: op1_13_inv18 = 1;
    14: op1_13_inv18 = 1;
    16: op1_13_inv18 = 1;
    20: op1_13_inv18 = 1;
    21: op1_13_inv18 = 1;
    23: op1_13_inv18 = 1;
    25: op1_13_inv18 = 1;
    26: op1_13_inv18 = 1;
    27: op1_13_inv18 = 1;
    30: op1_13_inv18 = 1;
    34: op1_13_inv18 = 1;
    36: op1_13_inv18 = 1;
    37: op1_13_inv18 = 1;
    39: op1_13_inv18 = 1;
    40: op1_13_inv18 = 1;
    41: op1_13_inv18 = 1;
    42: op1_13_inv18 = 1;
    45: op1_13_inv18 = 1;
    48: op1_13_inv18 = 1;
    49: op1_13_inv18 = 1;
    51: op1_13_inv18 = 1;
    54: op1_13_inv18 = 1;
    56: op1_13_inv18 = 1;
    57: op1_13_inv18 = 1;
    58: op1_13_inv18 = 1;
    59: op1_13_inv18 = 1;
    66: op1_13_inv18 = 1;
    69: op1_13_inv18 = 1;
    72: op1_13_inv18 = 1;
    74: op1_13_inv18 = 1;
    77: op1_13_inv18 = 1;
    78: op1_13_inv18 = 1;
    79: op1_13_inv18 = 1;
    83: op1_13_inv18 = 1;
    89: op1_13_inv18 = 1;
    90: op1_13_inv18 = 1;
    default: op1_13_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in19 = reg_0017;
    5: op1_13_in19 = imem05_in[3:0];
    6: op1_13_in19 = reg_0232;
    7: op1_13_in19 = reg_0355;
    8: op1_13_in19 = imem07_in[23:20];
    9: op1_13_in19 = imem05_in[75:72];
    10: op1_13_in19 = reg_0734;
    28: op1_13_in19 = reg_0734;
    11: op1_13_in19 = reg_0374;
    12: op1_13_in19 = reg_0499;
    13: op1_13_in19 = reg_0320;
    30: op1_13_in19 = reg_0320;
    14: op1_13_in19 = imem04_in[91:88];
    60: op1_13_in19 = imem04_in[91:88];
    15: op1_13_in19 = reg_0714;
    16: op1_13_in19 = imem01_in[95:92];
    17: op1_13_in19 = reg_0169;
    18: op1_13_in19 = imem01_in[47:44];
    20: op1_13_in19 = reg_0329;
    21: op1_13_in19 = reg_0076;
    22: op1_13_in19 = reg_0748;
    23: op1_13_in19 = reg_0136;
    24: op1_13_in19 = reg_0730;
    25: op1_13_in19 = imem04_in[15:12];
    31: op1_13_in19 = imem04_in[15:12];
    26: op1_13_in19 = reg_0453;
    27: op1_13_in19 = reg_0758;
    29: op1_13_in19 = reg_0038;
    32: op1_13_in19 = reg_0268;
    33: op1_13_in19 = reg_0235;
    34: op1_13_in19 = reg_0342;
    35: op1_13_in19 = reg_0080;
    79: op1_13_in19 = reg_0080;
    36: op1_13_in19 = reg_0266;
    37: op1_13_in19 = reg_0391;
    38: op1_13_in19 = reg_0422;
    39: op1_13_in19 = imem07_in[119:116];
    53: op1_13_in19 = imem07_in[119:116];
    40: op1_13_in19 = reg_0158;
    41: op1_13_in19 = reg_0531;
    42: op1_13_in19 = imem05_in[115:112];
    43: op1_13_in19 = reg_0298;
    44: op1_13_in19 = imem01_in[7:4];
    45: op1_13_in19 = reg_0564;
    46: op1_13_in19 = imem06_in[107:104];
    47: op1_13_in19 = imem01_in[79:76];
    48: op1_13_in19 = reg_0341;
    49: op1_13_in19 = reg_0202;
    51: op1_13_in19 = reg_0141;
    54: op1_13_in19 = reg_0735;
    55: op1_13_in19 = reg_0427;
    56: op1_13_in19 = reg_0638;
    57: op1_13_in19 = imem01_in[11:8];
    58: op1_13_in19 = reg_0083;
    59: op1_13_in19 = reg_0581;
    61: op1_13_in19 = reg_0719;
    62: op1_13_in19 = reg_0194;
    63: op1_13_in19 = reg_0203;
    64: op1_13_in19 = imem01_in[91:88];
    65: op1_13_in19 = reg_0657;
    66: op1_13_in19 = imem01_in[115:112];
    67: op1_13_in19 = reg_0140;
    68: op1_13_in19 = reg_0162;
    69: op1_13_in19 = reg_0533;
    70: op1_13_in19 = reg_0278;
    71: op1_13_in19 = reg_0196;
    72: op1_13_in19 = reg_0590;
    73: op1_13_in19 = imem03_in[15:12];
    74: op1_13_in19 = reg_0262;
    75: op1_13_in19 = reg_0099;
    77: op1_13_in19 = reg_0210;
    78: op1_13_in19 = reg_0210;
    80: op1_13_in19 = reg_0536;
    81: op1_13_in19 = reg_0112;
    83: op1_13_in19 = reg_0819;
    84: op1_13_in19 = reg_0414;
    85: op1_13_in19 = reg_0740;
    87: op1_13_in19 = reg_0514;
    89: op1_13_in19 = reg_0385;
    90: op1_13_in19 = reg_0471;
    91: op1_13_in19 = imem05_in[39:36];
    92: op1_13_in19 = reg_0307;
    93: op1_13_in19 = reg_0515;
    94: op1_13_in19 = reg_0579;
    95: op1_13_in19 = reg_0150;
    default: op1_13_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_13_inv19 = 1;
    11: op1_13_inv19 = 1;
    12: op1_13_inv19 = 1;
    13: op1_13_inv19 = 1;
    15: op1_13_inv19 = 1;
    16: op1_13_inv19 = 1;
    17: op1_13_inv19 = 1;
    18: op1_13_inv19 = 1;
    21: op1_13_inv19 = 1;
    22: op1_13_inv19 = 1;
    30: op1_13_inv19 = 1;
    31: op1_13_inv19 = 1;
    34: op1_13_inv19 = 1;
    36: op1_13_inv19 = 1;
    42: op1_13_inv19 = 1;
    43: op1_13_inv19 = 1;
    44: op1_13_inv19 = 1;
    45: op1_13_inv19 = 1;
    48: op1_13_inv19 = 1;
    53: op1_13_inv19 = 1;
    54: op1_13_inv19 = 1;
    55: op1_13_inv19 = 1;
    56: op1_13_inv19 = 1;
    58: op1_13_inv19 = 1;
    59: op1_13_inv19 = 1;
    60: op1_13_inv19 = 1;
    61: op1_13_inv19 = 1;
    63: op1_13_inv19 = 1;
    64: op1_13_inv19 = 1;
    66: op1_13_inv19 = 1;
    67: op1_13_inv19 = 1;
    69: op1_13_inv19 = 1;
    70: op1_13_inv19 = 1;
    72: op1_13_inv19 = 1;
    75: op1_13_inv19 = 1;
    78: op1_13_inv19 = 1;
    80: op1_13_inv19 = 1;
    83: op1_13_inv19 = 1;
    85: op1_13_inv19 = 1;
    90: op1_13_inv19 = 1;
    92: op1_13_inv19 = 1;
    94: op1_13_inv19 = 1;
    default: op1_13_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in20 = reg_0020;
    5: op1_13_in20 = imem05_in[7:4];
    6: op1_13_in20 = reg_0222;
    7: op1_13_in20 = reg_0095;
    8: op1_13_in20 = imem07_in[71:68];
    9: op1_13_in20 = imem05_in[103:100];
    10: op1_13_in20 = imem01_in[7:4];
    11: op1_13_in20 = reg_0389;
    12: op1_13_in20 = reg_0825;
    95: op1_13_in20 = reg_0825;
    13: op1_13_in20 = reg_0346;
    14: op1_13_in20 = reg_0545;
    74: op1_13_in20 = reg_0545;
    15: op1_13_in20 = reg_0724;
    16: op1_13_in20 = imem01_in[103:100];
    47: op1_13_in20 = imem01_in[103:100];
    17: op1_13_in20 = reg_0182;
    18: op1_13_in20 = imem01_in[67:64];
    20: op1_13_in20 = reg_0318;
    21: op1_13_in20 = reg_0070;
    22: op1_13_in20 = imem07_in[11:8];
    23: op1_13_in20 = reg_0129;
    24: op1_13_in20 = reg_0710;
    25: op1_13_in20 = imem04_in[19:16];
    31: op1_13_in20 = imem04_in[19:16];
    26: op1_13_in20 = reg_0469;
    27: op1_13_in20 = reg_0513;
    28: op1_13_in20 = reg_0089;
    29: op1_13_in20 = reg_0039;
    30: op1_13_in20 = reg_0345;
    32: op1_13_in20 = reg_0050;
    33: op1_13_in20 = reg_0511;
    34: op1_13_in20 = reg_0082;
    35: op1_13_in20 = reg_0082;
    36: op1_13_in20 = reg_0066;
    75: op1_13_in20 = reg_0066;
    37: op1_13_in20 = reg_0573;
    38: op1_13_in20 = reg_0447;
    39: op1_13_in20 = imem07_in[127:124];
    41: op1_13_in20 = reg_0094;
    42: op1_13_in20 = reg_0791;
    43: op1_13_in20 = reg_0633;
    44: op1_13_in20 = imem01_in[11:8];
    45: op1_13_in20 = reg_0517;
    46: op1_13_in20 = reg_0604;
    48: op1_13_in20 = reg_0359;
    49: op1_13_in20 = imem01_in[3:0];
    51: op1_13_in20 = reg_0137;
    53: op1_13_in20 = reg_0716;
    54: op1_13_in20 = reg_0496;
    55: op1_13_in20 = reg_0352;
    56: op1_13_in20 = reg_0485;
    57: op1_13_in20 = reg_0761;
    58: op1_13_in20 = reg_0555;
    59: op1_13_in20 = reg_0324;
    60: op1_13_in20 = imem04_in[99:96];
    61: op1_13_in20 = reg_0730;
    62: op1_13_in20 = reg_0213;
    63: op1_13_in20 = reg_0194;
    64: op1_13_in20 = imem01_in[95:92];
    65: op1_13_in20 = reg_0639;
    66: op1_13_in20 = reg_0735;
    67: op1_13_in20 = imem06_in[11:8];
    68: op1_13_in20 = reg_0167;
    69: op1_13_in20 = reg_0096;
    70: op1_13_in20 = reg_0150;
    71: op1_13_in20 = reg_0192;
    72: op1_13_in20 = reg_0518;
    73: op1_13_in20 = imem03_in[83:80];
    77: op1_13_in20 = reg_0189;
    78: op1_13_in20 = reg_0207;
    79: op1_13_in20 = reg_0756;
    80: op1_13_in20 = reg_0551;
    81: op1_13_in20 = reg_0102;
    83: op1_13_in20 = reg_0661;
    84: op1_13_in20 = reg_0527;
    85: op1_13_in20 = imem03_in[3:0];
    87: op1_13_in20 = reg_0043;
    89: op1_13_in20 = reg_0131;
    90: op1_13_in20 = reg_0456;
    91: op1_13_in20 = imem05_in[43:40];
    92: op1_13_in20 = reg_0037;
    93: op1_13_in20 = reg_0681;
    94: op1_13_in20 = reg_0547;
    default: op1_13_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv20 = 1;
    12: op1_13_inv20 = 1;
    14: op1_13_inv20 = 1;
    17: op1_13_inv20 = 1;
    18: op1_13_inv20 = 1;
    24: op1_13_inv20 = 1;
    25: op1_13_inv20 = 1;
    27: op1_13_inv20 = 1;
    35: op1_13_inv20 = 1;
    36: op1_13_inv20 = 1;
    37: op1_13_inv20 = 1;
    38: op1_13_inv20 = 1;
    41: op1_13_inv20 = 1;
    44: op1_13_inv20 = 1;
    46: op1_13_inv20 = 1;
    48: op1_13_inv20 = 1;
    53: op1_13_inv20 = 1;
    54: op1_13_inv20 = 1;
    55: op1_13_inv20 = 1;
    57: op1_13_inv20 = 1;
    60: op1_13_inv20 = 1;
    62: op1_13_inv20 = 1;
    63: op1_13_inv20 = 1;
    65: op1_13_inv20 = 1;
    66: op1_13_inv20 = 1;
    68: op1_13_inv20 = 1;
    69: op1_13_inv20 = 1;
    70: op1_13_inv20 = 1;
    71: op1_13_inv20 = 1;
    73: op1_13_inv20 = 1;
    74: op1_13_inv20 = 1;
    75: op1_13_inv20 = 1;
    78: op1_13_inv20 = 1;
    83: op1_13_inv20 = 1;
    84: op1_13_inv20 = 1;
    87: op1_13_inv20 = 1;
    92: op1_13_inv20 = 1;
    93: op1_13_inv20 = 1;
    94: op1_13_inv20 = 1;
    default: op1_13_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in21 = reg_0018;
    5: op1_13_in21 = imem05_in[71:68];
    6: op1_13_in21 = reg_0246;
    7: op1_13_in21 = reg_0082;
    69: op1_13_in21 = reg_0082;
    8: op1_13_in21 = imem07_in[75:72];
    9: op1_13_in21 = imem05_in[111:108];
    10: op1_13_in21 = imem01_in[11:8];
    11: op1_13_in21 = reg_0000;
    12: op1_13_in21 = reg_0517;
    13: op1_13_in21 = reg_0092;
    72: op1_13_in21 = reg_0092;
    14: op1_13_in21 = reg_0536;
    15: op1_13_in21 = reg_0708;
    16: op1_13_in21 = imem01_in[127:124];
    17: op1_13_in21 = reg_0160;
    18: op1_13_in21 = imem01_in[91:88];
    20: op1_13_in21 = reg_0342;
    21: op1_13_in21 = reg_0256;
    22: op1_13_in21 = imem07_in[23:20];
    23: op1_13_in21 = imem06_in[19:16];
    24: op1_13_in21 = reg_0731;
    53: op1_13_in21 = reg_0731;
    25: op1_13_in21 = imem04_in[43:40];
    26: op1_13_in21 = reg_0472;
    27: op1_13_in21 = reg_0337;
    28: op1_13_in21 = reg_0132;
    29: op1_13_in21 = reg_0753;
    65: op1_13_in21 = reg_0753;
    30: op1_13_in21 = reg_0540;
    31: op1_13_in21 = imem04_in[39:36];
    32: op1_13_in21 = reg_0278;
    33: op1_13_in21 = reg_0248;
    34: op1_13_in21 = reg_0538;
    35: op1_13_in21 = reg_0756;
    36: op1_13_in21 = reg_0067;
    37: op1_13_in21 = reg_0397;
    38: op1_13_in21 = reg_0428;
    39: op1_13_in21 = reg_0728;
    41: op1_13_in21 = imem03_in[11:8];
    79: op1_13_in21 = imem03_in[11:8];
    85: op1_13_in21 = imem03_in[11:8];
    42: op1_13_in21 = reg_0796;
    43: op1_13_in21 = reg_0618;
    44: op1_13_in21 = imem01_in[35:32];
    49: op1_13_in21 = imem01_in[35:32];
    45: op1_13_in21 = reg_0398;
    46: op1_13_in21 = reg_0247;
    47: op1_13_in21 = reg_0422;
    48: op1_13_in21 = reg_0518;
    51: op1_13_in21 = imem06_in[7:4];
    54: op1_13_in21 = reg_0761;
    55: op1_13_in21 = reg_0359;
    56: op1_13_in21 = reg_0358;
    57: op1_13_in21 = reg_0765;
    58: op1_13_in21 = reg_0510;
    59: op1_13_in21 = reg_0365;
    60: op1_13_in21 = imem04_in[111:108];
    61: op1_13_in21 = reg_0717;
    62: op1_13_in21 = imem01_in[31:28];
    63: op1_13_in21 = reg_0202;
    64: op1_13_in21 = imem01_in[115:112];
    66: op1_13_in21 = reg_0550;
    67: op1_13_in21 = imem06_in[67:64];
    68: op1_13_in21 = reg_0170;
    70: op1_13_in21 = reg_0151;
    71: op1_13_in21 = imem01_in[3:0];
    73: op1_13_in21 = imem03_in[107:104];
    74: op1_13_in21 = reg_0544;
    75: op1_13_in21 = reg_0285;
    77: op1_13_in21 = reg_0193;
    78: op1_13_in21 = reg_0186;
    80: op1_13_in21 = reg_0283;
    81: op1_13_in21 = reg_0114;
    83: op1_13_in21 = imem07_in[79:76];
    84: op1_13_in21 = imem02_in[7:4];
    87: op1_13_in21 = reg_0314;
    89: op1_13_in21 = reg_0394;
    90: op1_13_in21 = reg_0458;
    91: op1_13_in21 = imem05_in[99:96];
    92: op1_13_in21 = reg_0633;
    93: op1_13_in21 = reg_0621;
    94: op1_13_in21 = reg_0812;
    95: op1_13_in21 = reg_0829;
    default: op1_13_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv21 = 1;
    12: op1_13_inv21 = 1;
    13: op1_13_inv21 = 1;
    16: op1_13_inv21 = 1;
    17: op1_13_inv21 = 1;
    18: op1_13_inv21 = 1;
    20: op1_13_inv21 = 1;
    22: op1_13_inv21 = 1;
    23: op1_13_inv21 = 1;
    24: op1_13_inv21 = 1;
    29: op1_13_inv21 = 1;
    30: op1_13_inv21 = 1;
    32: op1_13_inv21 = 1;
    34: op1_13_inv21 = 1;
    35: op1_13_inv21 = 1;
    36: op1_13_inv21 = 1;
    38: op1_13_inv21 = 1;
    41: op1_13_inv21 = 1;
    44: op1_13_inv21 = 1;
    45: op1_13_inv21 = 1;
    47: op1_13_inv21 = 1;
    48: op1_13_inv21 = 1;
    54: op1_13_inv21 = 1;
    57: op1_13_inv21 = 1;
    58: op1_13_inv21 = 1;
    59: op1_13_inv21 = 1;
    63: op1_13_inv21 = 1;
    65: op1_13_inv21 = 1;
    73: op1_13_inv21 = 1;
    78: op1_13_inv21 = 1;
    79: op1_13_inv21 = 1;
    87: op1_13_inv21 = 1;
    90: op1_13_inv21 = 1;
    91: op1_13_inv21 = 1;
    92: op1_13_inv21 = 1;
    93: op1_13_inv21 = 1;
    94: op1_13_inv21 = 1;
    default: op1_13_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in22 = imem07_in[3:0];
    93: op1_13_in22 = imem07_in[3:0];
    5: op1_13_in22 = imem05_in[95:92];
    6: op1_13_in22 = reg_0224;
    92: op1_13_in22 = reg_0224;
    7: op1_13_in22 = reg_0055;
    8: op1_13_in22 = imem07_in[79:76];
    9: op1_13_in22 = imem05_in[123:120];
    10: op1_13_in22 = imem01_in[27:24];
    11: op1_13_in22 = reg_0811;
    12: op1_13_in22 = reg_0515;
    13: op1_13_in22 = reg_0084;
    14: op1_13_in22 = reg_0550;
    15: op1_13_in22 = reg_0707;
    16: op1_13_in22 = reg_0522;
    17: op1_13_in22 = reg_0183;
    18: op1_13_in22 = reg_0225;
    20: op1_13_in22 = reg_0336;
    21: op1_13_in22 = imem05_in[35:32];
    22: op1_13_in22 = imem07_in[123:120];
    23: op1_13_in22 = imem06_in[87:84];
    24: op1_13_in22 = reg_0703;
    25: op1_13_in22 = imem04_in[59:56];
    26: op1_13_in22 = reg_0200;
    27: op1_13_in22 = reg_0227;
    28: op1_13_in22 = reg_0145;
    29: op1_13_in22 = reg_0813;
    30: op1_13_in22 = reg_0535;
    31: op1_13_in22 = imem04_in[63:60];
    32: op1_13_in22 = reg_0257;
    33: op1_13_in22 = reg_0111;
    34: op1_13_in22 = reg_0740;
    35: op1_13_in22 = reg_0098;
    36: op1_13_in22 = reg_0072;
    37: op1_13_in22 = reg_0396;
    38: op1_13_in22 = reg_0443;
    39: op1_13_in22 = reg_0719;
    41: op1_13_in22 = imem03_in[71:68];
    42: op1_13_in22 = reg_0488;
    43: op1_13_in22 = reg_0370;
    44: op1_13_in22 = imem01_in[39:36];
    45: op1_13_in22 = reg_0374;
    46: op1_13_in22 = reg_0286;
    47: op1_13_in22 = reg_0574;
    48: op1_13_in22 = reg_0092;
    49: op1_13_in22 = imem01_in[47:44];
    51: op1_13_in22 = imem06_in[47:44];
    53: op1_13_in22 = reg_0713;
    54: op1_13_in22 = reg_0322;
    55: op1_13_in22 = reg_0353;
    56: op1_13_in22 = reg_0581;
    57: op1_13_in22 = reg_0649;
    58: op1_13_in22 = reg_0500;
    59: op1_13_in22 = reg_0527;
    60: op1_13_in22 = reg_0262;
    61: op1_13_in22 = reg_0064;
    62: op1_13_in22 = imem01_in[35:32];
    63: op1_13_in22 = imem01_in[19:16];
    64: op1_13_in22 = reg_0820;
    65: op1_13_in22 = reg_0342;
    66: op1_13_in22 = reg_0422;
    67: op1_13_in22 = imem06_in[75:72];
    69: op1_13_in22 = reg_0539;
    70: op1_13_in22 = reg_0142;
    71: op1_13_in22 = imem01_in[63:60];
    72: op1_13_in22 = reg_0314;
    73: op1_13_in22 = imem03_in[123:120];
    74: op1_13_in22 = reg_0315;
    75: op1_13_in22 = reg_0151;
    77: op1_13_in22 = reg_0194;
    78: op1_13_in22 = reg_0192;
    79: op1_13_in22 = imem03_in[35:32];
    80: op1_13_in22 = reg_0305;
    81: op1_13_in22 = reg_0397;
    83: op1_13_in22 = reg_0712;
    84: op1_13_in22 = imem02_in[91:88];
    85: op1_13_in22 = imem03_in[15:12];
    87: op1_13_in22 = reg_0487;
    89: op1_13_in22 = reg_0388;
    90: op1_13_in22 = reg_0198;
    91: op1_13_in22 = imem05_in[115:112];
    94: op1_13_in22 = reg_0827;
    95: op1_13_in22 = reg_0153;
    default: op1_13_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv22 = 1;
    5: op1_13_inv22 = 1;
    6: op1_13_inv22 = 1;
    8: op1_13_inv22 = 1;
    9: op1_13_inv22 = 1;
    10: op1_13_inv22 = 1;
    13: op1_13_inv22 = 1;
    14: op1_13_inv22 = 1;
    15: op1_13_inv22 = 1;
    16: op1_13_inv22 = 1;
    20: op1_13_inv22 = 1;
    23: op1_13_inv22 = 1;
    24: op1_13_inv22 = 1;
    25: op1_13_inv22 = 1;
    26: op1_13_inv22 = 1;
    31: op1_13_inv22 = 1;
    33: op1_13_inv22 = 1;
    35: op1_13_inv22 = 1;
    36: op1_13_inv22 = 1;
    37: op1_13_inv22 = 1;
    42: op1_13_inv22 = 1;
    44: op1_13_inv22 = 1;
    45: op1_13_inv22 = 1;
    46: op1_13_inv22 = 1;
    53: op1_13_inv22 = 1;
    54: op1_13_inv22 = 1;
    57: op1_13_inv22 = 1;
    58: op1_13_inv22 = 1;
    61: op1_13_inv22 = 1;
    64: op1_13_inv22 = 1;
    65: op1_13_inv22 = 1;
    66: op1_13_inv22 = 1;
    69: op1_13_inv22 = 1;
    70: op1_13_inv22 = 1;
    71: op1_13_inv22 = 1;
    85: op1_13_inv22 = 1;
    87: op1_13_inv22 = 1;
    92: op1_13_inv22 = 1;
    93: op1_13_inv22 = 1;
    94: op1_13_inv22 = 1;
    default: op1_13_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in23 = imem07_in[27:24];
    5: op1_13_in23 = imem05_in[107:104];
    6: op1_13_in23 = reg_0220;
    7: op1_13_in23 = reg_0077;
    8: op1_13_in23 = reg_0719;
    9: op1_13_in23 = imem05_in[127:124];
    91: op1_13_in23 = imem05_in[127:124];
    10: op1_13_in23 = imem01_in[115:112];
    11: op1_13_in23 = reg_0004;
    12: op1_13_in23 = reg_0516;
    13: op1_13_in23 = reg_0098;
    69: op1_13_in23 = reg_0098;
    14: op1_13_in23 = reg_0548;
    15: op1_13_in23 = reg_0700;
    16: op1_13_in23 = reg_0225;
    17: op1_13_in23 = reg_0170;
    18: op1_13_in23 = reg_0241;
    20: op1_13_in23 = imem02_in[27:24];
    21: op1_13_in23 = imem05_in[39:36];
    22: op1_13_in23 = reg_0723;
    23: op1_13_in23 = reg_0625;
    24: op1_13_in23 = reg_0712;
    25: op1_13_in23 = imem04_in[71:68];
    26: op1_13_in23 = reg_0197;
    27: op1_13_in23 = reg_0825;
    28: op1_13_in23 = reg_0135;
    29: op1_13_in23 = reg_0815;
    30: op1_13_in23 = reg_0756;
    31: op1_13_in23 = imem04_in[75:72];
    32: op1_13_in23 = reg_0281;
    33: op1_13_in23 = reg_0118;
    34: op1_13_in23 = imem03_in[3:0];
    35: op1_13_in23 = reg_0757;
    36: op1_13_in23 = imem05_in[7:4];
    37: op1_13_in23 = reg_0003;
    38: op1_13_in23 = reg_0448;
    39: op1_13_in23 = reg_0725;
    41: op1_13_in23 = imem03_in[115:112];
    42: op1_13_in23 = reg_0789;
    43: op1_13_in23 = reg_0409;
    44: op1_13_in23 = imem01_in[47:44];
    45: op1_13_in23 = reg_0006;
    46: op1_13_in23 = reg_0633;
    47: op1_13_in23 = reg_0054;
    48: op1_13_in23 = reg_0081;
    49: op1_13_in23 = reg_0735;
    51: op1_13_in23 = imem06_in[51:48];
    53: op1_13_in23 = reg_0061;
    54: op1_13_in23 = reg_0487;
    55: op1_13_in23 = reg_0414;
    56: op1_13_in23 = reg_0514;
    57: op1_13_in23 = reg_0737;
    58: op1_13_in23 = reg_0547;
    59: op1_13_in23 = reg_0590;
    60: op1_13_in23 = reg_0560;
    61: op1_13_in23 = reg_0253;
    62: op1_13_in23 = imem01_in[39:36];
    63: op1_13_in23 = imem01_in[35:32];
    64: op1_13_in23 = reg_0322;
    65: op1_13_in23 = reg_0092;
    66: op1_13_in23 = reg_0248;
    67: op1_13_in23 = imem06_in[95:92];
    70: op1_13_in23 = reg_0156;
    71: op1_13_in23 = reg_0497;
    72: op1_13_in23 = imem03_in[11:8];
    73: op1_13_in23 = reg_0559;
    74: op1_13_in23 = reg_0552;
    75: op1_13_in23 = reg_0828;
    95: op1_13_in23 = reg_0828;
    77: op1_13_in23 = imem01_in[19:16];
    78: op1_13_in23 = imem01_in[3:0];
    79: op1_13_in23 = imem03_in[39:36];
    80: op1_13_in23 = reg_0631;
    81: op1_13_in23 = reg_0507;
    83: op1_13_in23 = reg_0157;
    84: op1_13_in23 = imem02_in[95:92];
    85: op1_13_in23 = imem03_in[35:32];
    87: op1_13_in23 = reg_0136;
    89: op1_13_in23 = reg_0232;
    90: op1_13_in23 = reg_0190;
    92: op1_13_in23 = reg_0764;
    93: op1_13_in23 = imem07_in[11:8];
    94: op1_13_in23 = reg_0822;
    default: op1_13_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv23 = 1;
    10: op1_13_inv23 = 1;
    12: op1_13_inv23 = 1;
    13: op1_13_inv23 = 1;
    16: op1_13_inv23 = 1;
    20: op1_13_inv23 = 1;
    22: op1_13_inv23 = 1;
    24: op1_13_inv23 = 1;
    27: op1_13_inv23 = 1;
    29: op1_13_inv23 = 1;
    30: op1_13_inv23 = 1;
    31: op1_13_inv23 = 1;
    33: op1_13_inv23 = 1;
    34: op1_13_inv23 = 1;
    35: op1_13_inv23 = 1;
    36: op1_13_inv23 = 1;
    38: op1_13_inv23 = 1;
    39: op1_13_inv23 = 1;
    41: op1_13_inv23 = 1;
    44: op1_13_inv23 = 1;
    45: op1_13_inv23 = 1;
    46: op1_13_inv23 = 1;
    48: op1_13_inv23 = 1;
    58: op1_13_inv23 = 1;
    61: op1_13_inv23 = 1;
    63: op1_13_inv23 = 1;
    65: op1_13_inv23 = 1;
    67: op1_13_inv23 = 1;
    69: op1_13_inv23 = 1;
    70: op1_13_inv23 = 1;
    71: op1_13_inv23 = 1;
    74: op1_13_inv23 = 1;
    77: op1_13_inv23 = 1;
    78: op1_13_inv23 = 1;
    79: op1_13_inv23 = 1;
    80: op1_13_inv23 = 1;
    87: op1_13_inv23 = 1;
    89: op1_13_inv23 = 1;
    90: op1_13_inv23 = 1;
    91: op1_13_inv23 = 1;
    95: op1_13_inv23 = 1;
    default: op1_13_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in24 = reg_0722;
    5: op1_13_in24 = imem05_in[119:116];
    6: op1_13_in24 = reg_0247;
    7: op1_13_in24 = reg_0093;
    8: op1_13_in24 = reg_0726;
    9: op1_13_in24 = reg_0788;
    10: op1_13_in24 = imem01_in[119:116];
    11: op1_13_in24 = imem04_in[55:52];
    12: op1_13_in24 = reg_0505;
    18: op1_13_in24 = reg_0505;
    13: op1_13_in24 = reg_0055;
    14: op1_13_in24 = reg_0558;
    15: op1_13_in24 = reg_0423;
    16: op1_13_in24 = reg_0215;
    17: op1_13_in24 = reg_0176;
    20: op1_13_in24 = imem02_in[47:44];
    21: op1_13_in24 = imem05_in[55:52];
    22: op1_13_in24 = reg_0711;
    23: op1_13_in24 = reg_0604;
    24: op1_13_in24 = reg_0707;
    25: op1_13_in24 = imem04_in[87:84];
    26: op1_13_in24 = imem01_in[7:4];
    27: op1_13_in24 = reg_0333;
    28: op1_13_in24 = reg_0151;
    94: op1_13_in24 = reg_0151;
    29: op1_13_in24 = reg_0814;
    30: op1_13_in24 = reg_0380;
    31: op1_13_in24 = imem04_in[115:112];
    32: op1_13_in24 = reg_0299;
    33: op1_13_in24 = imem02_in[35:32];
    34: op1_13_in24 = imem03_in[15:12];
    35: op1_13_in24 = imem03_in[7:4];
    36: op1_13_in24 = imem05_in[31:28];
    37: op1_13_in24 = reg_0807;
    38: op1_13_in24 = reg_0431;
    39: op1_13_in24 = reg_0706;
    41: op1_13_in24 = imem03_in[127:124];
    42: op1_13_in24 = reg_0492;
    43: op1_13_in24 = reg_0748;
    44: op1_13_in24 = imem01_in[55:52];
    45: op1_13_in24 = reg_0009;
    46: op1_13_in24 = reg_0766;
    47: op1_13_in24 = reg_0502;
    48: op1_13_in24 = reg_0540;
    49: op1_13_in24 = reg_0497;
    51: op1_13_in24 = imem06_in[87:84];
    53: op1_13_in24 = reg_0239;
    54: op1_13_in24 = reg_0217;
    55: op1_13_in24 = reg_0406;
    56: op1_13_in24 = reg_0530;
    57: op1_13_in24 = reg_0422;
    58: op1_13_in24 = reg_0429;
    59: op1_13_in24 = reg_0541;
    60: op1_13_in24 = reg_0552;
    61: op1_13_in24 = reg_0445;
    62: op1_13_in24 = imem01_in[107:104];
    63: op1_13_in24 = imem01_in[59:56];
    64: op1_13_in24 = reg_0550;
    65: op1_13_in24 = reg_0095;
    66: op1_13_in24 = reg_0419;
    67: op1_13_in24 = imem06_in[119:116];
    69: op1_13_in24 = reg_0094;
    70: op1_13_in24 = reg_0154;
    71: op1_13_in24 = reg_0112;
    72: op1_13_in24 = imem03_in[47:44];
    73: op1_13_in24 = reg_0493;
    74: op1_13_in24 = reg_0056;
    75: op1_13_in24 = imem06_in[3:0];
    77: op1_13_in24 = imem01_in[27:24];
    78: op1_13_in24 = imem01_in[23:20];
    79: op1_13_in24 = imem03_in[59:56];
    80: op1_13_in24 = reg_0077;
    81: op1_13_in24 = reg_0232;
    83: op1_13_in24 = reg_0334;
    84: op1_13_in24 = imem02_in[115:112];
    85: op1_13_in24 = imem03_in[39:36];
    87: op1_13_in24 = reg_0757;
    89: op1_13_in24 = reg_0511;
    90: op1_13_in24 = imem01_in[35:32];
    91: op1_13_in24 = reg_0337;
    92: op1_13_in24 = imem07_in[31:28];
    93: op1_13_in24 = imem07_in[71:68];
    95: op1_13_in24 = reg_0824;
    default: op1_13_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_13_inv24 = 1;
    9: op1_13_inv24 = 1;
    14: op1_13_inv24 = 1;
    15: op1_13_inv24 = 1;
    16: op1_13_inv24 = 1;
    22: op1_13_inv24 = 1;
    23: op1_13_inv24 = 1;
    24: op1_13_inv24 = 1;
    25: op1_13_inv24 = 1;
    26: op1_13_inv24 = 1;
    27: op1_13_inv24 = 1;
    28: op1_13_inv24 = 1;
    31: op1_13_inv24 = 1;
    32: op1_13_inv24 = 1;
    33: op1_13_inv24 = 1;
    35: op1_13_inv24 = 1;
    36: op1_13_inv24 = 1;
    37: op1_13_inv24 = 1;
    38: op1_13_inv24 = 1;
    41: op1_13_inv24 = 1;
    45: op1_13_inv24 = 1;
    51: op1_13_inv24 = 1;
    54: op1_13_inv24 = 1;
    56: op1_13_inv24 = 1;
    59: op1_13_inv24 = 1;
    62: op1_13_inv24 = 1;
    64: op1_13_inv24 = 1;
    71: op1_13_inv24 = 1;
    73: op1_13_inv24 = 1;
    77: op1_13_inv24 = 1;
    78: op1_13_inv24 = 1;
    80: op1_13_inv24 = 1;
    85: op1_13_inv24 = 1;
    87: op1_13_inv24 = 1;
    91: op1_13_inv24 = 1;
    92: op1_13_inv24 = 1;
    93: op1_13_inv24 = 1;
    94: op1_13_inv24 = 1;
    default: op1_13_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in25 = reg_0710;
    5: op1_13_in25 = reg_0215;
    6: op1_13_in25 = reg_0236;
    7: op1_13_in25 = imem03_in[15:12];
    8: op1_13_in25 = reg_0725;
    9: op1_13_in25 = reg_0783;
    10: op1_13_in25 = reg_0232;
    11: op1_13_in25 = imem04_in[59:56];
    12: op1_13_in25 = reg_0233;
    13: op1_13_in25 = imem03_in[19:16];
    84: op1_13_in25 = imem03_in[19:16];
    14: op1_13_in25 = reg_0531;
    15: op1_13_in25 = reg_0439;
    16: op1_13_in25 = reg_0246;
    18: op1_13_in25 = reg_0511;
    20: op1_13_in25 = imem02_in[55:52];
    21: op1_13_in25 = imem05_in[79:76];
    22: op1_13_in25 = reg_0425;
    23: op1_13_in25 = reg_0607;
    24: op1_13_in25 = reg_0701;
    25: op1_13_in25 = imem04_in[95:92];
    26: op1_13_in25 = imem01_in[39:36];
    27: op1_13_in25 = reg_0557;
    28: op1_13_in25 = reg_0146;
    29: op1_13_in25 = reg_0036;
    30: op1_13_in25 = reg_0040;
    31: op1_13_in25 = imem04_in[119:116];
    32: op1_13_in25 = reg_0077;
    33: op1_13_in25 = imem02_in[51:48];
    34: op1_13_in25 = imem03_in[35:32];
    35: op1_13_in25 = imem03_in[11:8];
    59: op1_13_in25 = imem03_in[11:8];
    36: op1_13_in25 = imem05_in[67:64];
    37: op1_13_in25 = reg_0809;
    38: op1_13_in25 = reg_0180;
    39: op1_13_in25 = reg_0436;
    41: op1_13_in25 = reg_0395;
    42: op1_13_in25 = reg_0780;
    43: op1_13_in25 = reg_0818;
    44: op1_13_in25 = imem01_in[115:112];
    62: op1_13_in25 = imem01_in[115:112];
    45: op1_13_in25 = reg_0069;
    46: op1_13_in25 = reg_0612;
    47: op1_13_in25 = reg_0244;
    48: op1_13_in25 = reg_0082;
    65: op1_13_in25 = reg_0082;
    49: op1_13_in25 = reg_0496;
    51: op1_13_in25 = imem06_in[103:100];
    53: op1_13_in25 = reg_0167;
    54: op1_13_in25 = reg_0419;
    55: op1_13_in25 = reg_0343;
    56: op1_13_in25 = reg_0498;
    57: op1_13_in25 = reg_0574;
    89: op1_13_in25 = reg_0574;
    58: op1_13_in25 = reg_0631;
    60: op1_13_in25 = reg_0500;
    61: op1_13_in25 = reg_0442;
    63: op1_13_in25 = imem01_in[67:64];
    64: op1_13_in25 = reg_0421;
    66: op1_13_in25 = reg_0424;
    67: op1_13_in25 = imem06_in[123:120];
    69: op1_13_in25 = reg_0039;
    70: op1_13_in25 = reg_0144;
    71: op1_13_in25 = reg_0397;
    72: op1_13_in25 = imem03_in[79:76];
    73: op1_13_in25 = reg_0357;
    74: op1_13_in25 = reg_0516;
    75: op1_13_in25 = imem06_in[23:20];
    77: op1_13_in25 = imem01_in[35:32];
    78: op1_13_in25 = imem01_in[27:24];
    79: op1_13_in25 = imem03_in[123:120];
    80: op1_13_in25 = reg_0071;
    81: op1_13_in25 = reg_0240;
    83: op1_13_in25 = reg_0053;
    85: op1_13_in25 = imem03_in[67:64];
    87: op1_13_in25 = reg_0315;
    90: op1_13_in25 = imem01_in[103:100];
    91: op1_13_in25 = reg_0641;
    92: op1_13_in25 = imem07_in[87:84];
    93: op1_13_in25 = imem07_in[99:96];
    94: op1_13_in25 = reg_0257;
    95: op1_13_in25 = imem06_in[3:0];
    default: op1_13_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv25 = 1;
    5: op1_13_inv25 = 1;
    7: op1_13_inv25 = 1;
    10: op1_13_inv25 = 1;
    11: op1_13_inv25 = 1;
    13: op1_13_inv25 = 1;
    18: op1_13_inv25 = 1;
    23: op1_13_inv25 = 1;
    24: op1_13_inv25 = 1;
    25: op1_13_inv25 = 1;
    26: op1_13_inv25 = 1;
    27: op1_13_inv25 = 1;
    33: op1_13_inv25 = 1;
    34: op1_13_inv25 = 1;
    35: op1_13_inv25 = 1;
    36: op1_13_inv25 = 1;
    37: op1_13_inv25 = 1;
    39: op1_13_inv25 = 1;
    41: op1_13_inv25 = 1;
    44: op1_13_inv25 = 1;
    46: op1_13_inv25 = 1;
    48: op1_13_inv25 = 1;
    49: op1_13_inv25 = 1;
    51: op1_13_inv25 = 1;
    53: op1_13_inv25 = 1;
    59: op1_13_inv25 = 1;
    60: op1_13_inv25 = 1;
    63: op1_13_inv25 = 1;
    64: op1_13_inv25 = 1;
    65: op1_13_inv25 = 1;
    71: op1_13_inv25 = 1;
    81: op1_13_inv25 = 1;
    84: op1_13_inv25 = 1;
    85: op1_13_inv25 = 1;
    89: op1_13_inv25 = 1;
    91: op1_13_inv25 = 1;
    default: op1_13_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in26 = reg_0723;
    5: op1_13_in26 = reg_0259;
    6: op1_13_in26 = reg_0248;
    57: op1_13_in26 = reg_0248;
    7: op1_13_in26 = imem03_in[23:20];
    13: op1_13_in26 = imem03_in[23:20];
    8: op1_13_in26 = reg_0714;
    9: op1_13_in26 = reg_0268;
    10: op1_13_in26 = reg_0217;
    11: op1_13_in26 = imem04_in[63:60];
    12: op1_13_in26 = reg_0246;
    14: op1_13_in26 = reg_0547;
    15: op1_13_in26 = reg_0427;
    16: op1_13_in26 = reg_0506;
    47: op1_13_in26 = reg_0506;
    18: op1_13_in26 = reg_0218;
    20: op1_13_in26 = imem02_in[59:56];
    21: op1_13_in26 = imem05_in[83:80];
    36: op1_13_in26 = imem05_in[83:80];
    22: op1_13_in26 = reg_0424;
    54: op1_13_in26 = reg_0424;
    23: op1_13_in26 = reg_0631;
    24: op1_13_in26 = reg_0706;
    25: op1_13_in26 = imem04_in[119:116];
    26: op1_13_in26 = imem01_in[67:64];
    27: op1_13_in26 = reg_0550;
    28: op1_13_in26 = reg_0154;
    29: op1_13_in26 = reg_0029;
    30: op1_13_in26 = reg_0338;
    31: op1_13_in26 = reg_0544;
    32: op1_13_in26 = reg_0069;
    33: op1_13_in26 = imem02_in[67:64];
    34: op1_13_in26 = imem03_in[39:36];
    35: op1_13_in26 = imem03_in[39:36];
    37: op1_13_in26 = imem04_in[83:80];
    38: op1_13_in26 = reg_0165;
    39: op1_13_in26 = reg_0434;
    41: op1_13_in26 = reg_0387;
    42: op1_13_in26 = reg_0783;
    43: op1_13_in26 = reg_0238;
    44: op1_13_in26 = reg_0497;
    45: op1_13_in26 = reg_0296;
    46: op1_13_in26 = reg_0821;
    48: op1_13_in26 = reg_0526;
    49: op1_13_in26 = reg_0761;
    51: op1_13_in26 = imem06_in[119:116];
    53: op1_13_in26 = reg_0160;
    55: op1_13_in26 = reg_0518;
    56: op1_13_in26 = imem03_in[11:8];
    58: op1_13_in26 = reg_0074;
    59: op1_13_in26 = imem03_in[31:28];
    60: op1_13_in26 = reg_0079;
    61: op1_13_in26 = reg_0267;
    62: op1_13_in26 = imem01_in[119:116];
    63: op1_13_in26 = imem01_in[91:88];
    64: op1_13_in26 = reg_0306;
    65: op1_13_in26 = reg_0098;
    66: op1_13_in26 = reg_0105;
    67: op1_13_in26 = reg_0577;
    69: op1_13_in26 = reg_0090;
    70: op1_13_in26 = reg_0812;
    71: op1_13_in26 = reg_0760;
    72: op1_13_in26 = reg_0602;
    73: op1_13_in26 = reg_0588;
    74: op1_13_in26 = reg_0052;
    75: op1_13_in26 = imem06_in[27:24];
    77: op1_13_in26 = imem01_in[75:72];
    78: op1_13_in26 = imem01_in[39:36];
    79: op1_13_in26 = reg_0347;
    80: op1_13_in26 = reg_0508;
    81: op1_13_in26 = reg_0290;
    83: op1_13_in26 = reg_0061;
    84: op1_13_in26 = imem03_in[99:96];
    85: op1_13_in26 = imem03_in[87:84];
    87: op1_13_in26 = reg_0063;
    89: op1_13_in26 = reg_0567;
    90: op1_13_in26 = imem01_in[111:108];
    91: op1_13_in26 = reg_0231;
    92: op1_13_in26 = imem07_in[99:96];
    93: op1_13_in26 = reg_0726;
    94: op1_13_in26 = reg_0828;
    95: op1_13_in26 = imem06_in[47:44];
    default: op1_13_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv26 = 1;
    12: op1_13_inv26 = 1;
    15: op1_13_inv26 = 1;
    16: op1_13_inv26 = 1;
    18: op1_13_inv26 = 1;
    26: op1_13_inv26 = 1;
    28: op1_13_inv26 = 1;
    29: op1_13_inv26 = 1;
    30: op1_13_inv26 = 1;
    31: op1_13_inv26 = 1;
    32: op1_13_inv26 = 1;
    33: op1_13_inv26 = 1;
    37: op1_13_inv26 = 1;
    42: op1_13_inv26 = 1;
    43: op1_13_inv26 = 1;
    44: op1_13_inv26 = 1;
    47: op1_13_inv26 = 1;
    48: op1_13_inv26 = 1;
    53: op1_13_inv26 = 1;
    54: op1_13_inv26 = 1;
    57: op1_13_inv26 = 1;
    58: op1_13_inv26 = 1;
    60: op1_13_inv26 = 1;
    61: op1_13_inv26 = 1;
    63: op1_13_inv26 = 1;
    64: op1_13_inv26 = 1;
    67: op1_13_inv26 = 1;
    69: op1_13_inv26 = 1;
    72: op1_13_inv26 = 1;
    74: op1_13_inv26 = 1;
    75: op1_13_inv26 = 1;
    77: op1_13_inv26 = 1;
    79: op1_13_inv26 = 1;
    80: op1_13_inv26 = 1;
    83: op1_13_inv26 = 1;
    89: op1_13_inv26 = 1;
    90: op1_13_inv26 = 1;
    91: op1_13_inv26 = 1;
    92: op1_13_inv26 = 1;
    default: op1_13_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in27 = reg_0724;
    5: op1_13_in27 = reg_0270;
    6: op1_13_in27 = reg_0245;
    7: op1_13_in27 = imem03_in[27:24];
    8: op1_13_in27 = reg_0701;
    9: op1_13_in27 = reg_0250;
    10: op1_13_in27 = reg_0504;
    11: op1_13_in27 = imem04_in[83:80];
    12: op1_13_in27 = reg_0218;
    13: op1_13_in27 = imem03_in[111:108];
    14: op1_13_in27 = reg_0281;
    15: op1_13_in27 = reg_0420;
    16: op1_13_in27 = reg_0242;
    18: op1_13_in27 = reg_0506;
    20: op1_13_in27 = imem02_in[67:64];
    21: op1_13_in27 = imem05_in[103:100];
    36: op1_13_in27 = imem05_in[103:100];
    22: op1_13_in27 = reg_0429;
    23: op1_13_in27 = reg_0626;
    24: op1_13_in27 = reg_0424;
    25: op1_13_in27 = imem04_in[127:124];
    26: op1_13_in27 = imem01_in[71:68];
    27: op1_13_in27 = reg_0240;
    71: op1_13_in27 = reg_0240;
    28: op1_13_in27 = reg_0139;
    29: op1_13_in27 = reg_0751;
    30: op1_13_in27 = reg_0368;
    31: op1_13_in27 = reg_0315;
    32: op1_13_in27 = reg_0256;
    33: op1_13_in27 = imem02_in[83:80];
    34: op1_13_in27 = imem03_in[43:40];
    35: op1_13_in27 = imem03_in[67:64];
    37: op1_13_in27 = imem04_in[123:120];
    38: op1_13_in27 = reg_0179;
    39: op1_13_in27 = reg_0438;
    41: op1_13_in27 = reg_0388;
    42: op1_13_in27 = reg_0304;
    43: op1_13_in27 = reg_0367;
    44: op1_13_in27 = reg_0513;
    45: op1_13_in27 = reg_0249;
    46: op1_13_in27 = reg_0776;
    47: op1_13_in27 = reg_0219;
    48: op1_13_in27 = imem03_in[3:0];
    49: op1_13_in27 = reg_0100;
    51: op1_13_in27 = reg_0624;
    53: op1_13_in27 = reg_0163;
    54: op1_13_in27 = reg_0123;
    81: op1_13_in27 = reg_0123;
    55: op1_13_in27 = reg_0092;
    56: op1_13_in27 = imem03_in[15:12];
    57: op1_13_in27 = reg_0505;
    58: op1_13_in27 = imem04_in[11:8];
    59: op1_13_in27 = imem03_in[39:36];
    60: op1_13_in27 = reg_0631;
    61: op1_13_in27 = reg_0161;
    62: op1_13_in27 = reg_0761;
    63: op1_13_in27 = imem01_in[107:104];
    64: op1_13_in27 = reg_0220;
    65: op1_13_in27 = reg_0498;
    66: op1_13_in27 = reg_0675;
    67: op1_13_in27 = reg_0298;
    69: op1_13_in27 = reg_0599;
    70: op1_13_in27 = reg_0032;
    72: op1_13_in27 = reg_0347;
    73: op1_13_in27 = reg_0564;
    74: op1_13_in27 = reg_0529;
    75: op1_13_in27 = imem06_in[63:60];
    77: op1_13_in27 = imem01_in[95:92];
    78: op1_13_in27 = reg_0085;
    79: op1_13_in27 = reg_0317;
    80: op1_13_in27 = reg_0050;
    83: op1_13_in27 = reg_0445;
    84: op1_13_in27 = reg_0582;
    85: op1_13_in27 = imem03_in[103:100];
    87: op1_13_in27 = reg_0329;
    89: op1_13_in27 = reg_0502;
    90: op1_13_in27 = imem01_in[115:112];
    91: op1_13_in27 = reg_0499;
    92: op1_13_in27 = reg_0726;
    93: op1_13_in27 = reg_0164;
    94: op1_13_in27 = imem06_in[75:72];
    95: op1_13_in27 = imem06_in[75:72];
    default: op1_13_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_13_inv27 = 1;
    7: op1_13_inv27 = 1;
    8: op1_13_inv27 = 1;
    10: op1_13_inv27 = 1;
    13: op1_13_inv27 = 1;
    14: op1_13_inv27 = 1;
    16: op1_13_inv27 = 1;
    18: op1_13_inv27 = 1;
    20: op1_13_inv27 = 1;
    21: op1_13_inv27 = 1;
    23: op1_13_inv27 = 1;
    24: op1_13_inv27 = 1;
    29: op1_13_inv27 = 1;
    30: op1_13_inv27 = 1;
    32: op1_13_inv27 = 1;
    33: op1_13_inv27 = 1;
    35: op1_13_inv27 = 1;
    36: op1_13_inv27 = 1;
    37: op1_13_inv27 = 1;
    41: op1_13_inv27 = 1;
    42: op1_13_inv27 = 1;
    43: op1_13_inv27 = 1;
    44: op1_13_inv27 = 1;
    46: op1_13_inv27 = 1;
    47: op1_13_inv27 = 1;
    48: op1_13_inv27 = 1;
    53: op1_13_inv27 = 1;
    55: op1_13_inv27 = 1;
    56: op1_13_inv27 = 1;
    58: op1_13_inv27 = 1;
    59: op1_13_inv27 = 1;
    62: op1_13_inv27 = 1;
    64: op1_13_inv27 = 1;
    65: op1_13_inv27 = 1;
    67: op1_13_inv27 = 1;
    71: op1_13_inv27 = 1;
    72: op1_13_inv27 = 1;
    77: op1_13_inv27 = 1;
    81: op1_13_inv27 = 1;
    83: op1_13_inv27 = 1;
    84: op1_13_inv27 = 1;
    85: op1_13_inv27 = 1;
    87: op1_13_inv27 = 1;
    89: op1_13_inv27 = 1;
    92: op1_13_inv27 = 1;
    93: op1_13_inv27 = 1;
    94: op1_13_inv27 = 1;
    95: op1_13_inv27 = 1;
    default: op1_13_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in28 = reg_0707;
    5: op1_13_in28 = reg_0253;
    9: op1_13_in28 = reg_0253;
    6: op1_13_in28 = reg_0238;
    7: op1_13_in28 = imem03_in[51:48];
    8: op1_13_in28 = reg_0422;
    10: op1_13_in28 = reg_0243;
    11: op1_13_in28 = imem04_in[87:84];
    12: op1_13_in28 = reg_0242;
    13: op1_13_in28 = imem03_in[123:120];
    14: op1_13_in28 = reg_0295;
    15: op1_13_in28 = reg_0169;
    61: op1_13_in28 = reg_0169;
    16: op1_13_in28 = reg_0502;
    18: op1_13_in28 = reg_0239;
    20: op1_13_in28 = imem02_in[83:80];
    21: op1_13_in28 = imem05_in[111:108];
    22: op1_13_in28 = reg_0434;
    23: op1_13_in28 = reg_0615;
    24: op1_13_in28 = reg_0436;
    25: op1_13_in28 = reg_0545;
    45: op1_13_in28 = reg_0545;
    26: op1_13_in28 = imem01_in[111:108];
    27: op1_13_in28 = reg_0118;
    28: op1_13_in28 = reg_0153;
    29: op1_13_in28 = imem07_in[23:20];
    30: op1_13_in28 = reg_0381;
    31: op1_13_in28 = reg_0057;
    32: op1_13_in28 = imem05_in[31:28];
    33: op1_13_in28 = imem02_in[107:104];
    34: op1_13_in28 = imem03_in[47:44];
    59: op1_13_in28 = imem03_in[47:44];
    35: op1_13_in28 = imem03_in[79:76];
    36: op1_13_in28 = reg_0791;
    37: op1_13_in28 = imem04_in[127:124];
    38: op1_13_in28 = reg_0166;
    39: op1_13_in28 = reg_0448;
    41: op1_13_in28 = reg_0373;
    42: op1_13_in28 = reg_0733;
    43: op1_13_in28 = imem07_in[35:32];
    44: op1_13_in28 = reg_0520;
    46: op1_13_in28 = reg_0319;
    79: op1_13_in28 = reg_0319;
    47: op1_13_in28 = reg_0505;
    48: op1_13_in28 = imem03_in[39:36];
    49: op1_13_in28 = reg_0216;
    71: op1_13_in28 = reg_0216;
    51: op1_13_in28 = reg_0613;
    53: op1_13_in28 = reg_0178;
    54: op1_13_in28 = reg_0125;
    55: op1_13_in28 = reg_0080;
    56: op1_13_in28 = imem03_in[31:28];
    57: op1_13_in28 = reg_0124;
    58: op1_13_in28 = imem04_in[67:64];
    60: op1_13_in28 = reg_0627;
    62: op1_13_in28 = reg_0825;
    63: op1_13_in28 = imem01_in[127:124];
    64: op1_13_in28 = reg_0504;
    65: op1_13_in28 = reg_0093;
    66: op1_13_in28 = reg_0121;
    67: op1_13_in28 = reg_0401;
    69: op1_13_in28 = reg_0750;
    70: op1_13_in28 = reg_0275;
    72: op1_13_in28 = reg_0589;
    73: op1_13_in28 = reg_0496;
    74: op1_13_in28 = reg_0508;
    75: op1_13_in28 = imem06_in[95:92];
    77: op1_13_in28 = imem01_in[107:104];
    78: op1_13_in28 = reg_0497;
    80: op1_13_in28 = reg_0610;
    81: op1_13_in28 = reg_0673;
    83: op1_13_in28 = reg_0444;
    84: op1_13_in28 = reg_0350;
    85: op1_13_in28 = imem03_in[107:104];
    87: op1_13_in28 = reg_0163;
    89: op1_13_in28 = reg_0105;
    90: op1_13_in28 = reg_0759;
    91: op1_13_in28 = reg_0488;
    92: op1_13_in28 = reg_0382;
    93: op1_13_in28 = reg_0713;
    94: op1_13_in28 = imem06_in[123:120];
    95: op1_13_in28 = imem06_in[127:124];
    default: op1_13_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv28 = 1;
    7: op1_13_inv28 = 1;
    8: op1_13_inv28 = 1;
    9: op1_13_inv28 = 1;
    11: op1_13_inv28 = 1;
    12: op1_13_inv28 = 1;
    13: op1_13_inv28 = 1;
    16: op1_13_inv28 = 1;
    21: op1_13_inv28 = 1;
    24: op1_13_inv28 = 1;
    27: op1_13_inv28 = 1;
    30: op1_13_inv28 = 1;
    31: op1_13_inv28 = 1;
    32: op1_13_inv28 = 1;
    34: op1_13_inv28 = 1;
    39: op1_13_inv28 = 1;
    41: op1_13_inv28 = 1;
    46: op1_13_inv28 = 1;
    49: op1_13_inv28 = 1;
    51: op1_13_inv28 = 1;
    53: op1_13_inv28 = 1;
    59: op1_13_inv28 = 1;
    65: op1_13_inv28 = 1;
    66: op1_13_inv28 = 1;
    69: op1_13_inv28 = 1;
    70: op1_13_inv28 = 1;
    72: op1_13_inv28 = 1;
    73: op1_13_inv28 = 1;
    74: op1_13_inv28 = 1;
    75: op1_13_inv28 = 1;
    78: op1_13_inv28 = 1;
    79: op1_13_inv28 = 1;
    80: op1_13_inv28 = 1;
    81: op1_13_inv28 = 1;
    83: op1_13_inv28 = 1;
    85: op1_13_inv28 = 1;
    87: op1_13_inv28 = 1;
    89: op1_13_inv28 = 1;
    90: op1_13_inv28 = 1;
    91: op1_13_inv28 = 1;
    92: op1_13_inv28 = 1;
    93: op1_13_inv28 = 1;
    default: op1_13_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in29 = reg_0700;
    5: op1_13_in29 = reg_0263;
    6: op1_13_in29 = reg_0219;
    7: op1_13_in29 = imem03_in[75:72];
    8: op1_13_in29 = reg_0447;
    9: op1_13_in29 = reg_0147;
    10: op1_13_in29 = reg_0112;
    11: op1_13_in29 = imem04_in[99:96];
    12: op1_13_in29 = reg_0502;
    13: op1_13_in29 = reg_0586;
    14: op1_13_in29 = reg_0286;
    15: op1_13_in29 = reg_0163;
    16: op1_13_in29 = reg_0247;
    18: op1_13_in29 = reg_0217;
    20: op1_13_in29 = imem02_in[95:92];
    21: op1_13_in29 = imem05_in[115:112];
    22: op1_13_in29 = reg_0449;
    23: op1_13_in29 = reg_0406;
    24: op1_13_in29 = reg_0421;
    25: op1_13_in29 = reg_0087;
    26: op1_13_in29 = imem01_in[123:120];
    27: op1_13_in29 = reg_0119;
    28: op1_13_in29 = reg_0130;
    29: op1_13_in29 = imem07_in[47:44];
    43: op1_13_in29 = imem07_in[47:44];
    30: op1_13_in29 = imem03_in[19:16];
    31: op1_13_in29 = reg_0500;
    32: op1_13_in29 = imem05_in[75:72];
    33: op1_13_in29 = reg_0650;
    34: op1_13_in29 = imem03_in[67:64];
    35: op1_13_in29 = imem03_in[95:92];
    36: op1_13_in29 = reg_0798;
    37: op1_13_in29 = reg_0542;
    38: op1_13_in29 = reg_0164;
    39: op1_13_in29 = reg_0431;
    41: op1_13_in29 = reg_0385;
    42: op1_13_in29 = reg_0149;
    44: op1_13_in29 = reg_0514;
    45: op1_13_in29 = reg_0055;
    46: op1_13_in29 = reg_0607;
    47: op1_13_in29 = reg_0105;
    48: op1_13_in29 = imem03_in[43:40];
    49: op1_13_in29 = reg_0425;
    51: op1_13_in29 = reg_0606;
    53: op1_13_in29 = reg_0158;
    54: op1_13_in29 = reg_0104;
    55: op1_13_in29 = reg_0531;
    56: op1_13_in29 = imem03_in[39:36];
    57: op1_13_in29 = reg_0125;
    81: op1_13_in29 = reg_0125;
    58: op1_13_in29 = imem04_in[95:92];
    59: op1_13_in29 = imem03_in[51:48];
    60: op1_13_in29 = reg_0626;
    61: op1_13_in29 = reg_0166;
    62: op1_13_in29 = reg_0760;
    63: op1_13_in29 = reg_0733;
    64: op1_13_in29 = reg_0424;
    65: op1_13_in29 = imem03_in[27:24];
    66: op1_13_in29 = imem02_in[7:4];
    67: op1_13_in29 = reg_0260;
    69: op1_13_in29 = reg_0318;
    70: op1_13_in29 = reg_0656;
    71: op1_13_in29 = reg_0123;
    72: op1_13_in29 = reg_0597;
    73: op1_13_in29 = reg_0811;
    74: op1_13_in29 = reg_0779;
    75: op1_13_in29 = reg_0348;
    77: op1_13_in29 = imem01_in[111:108];
    78: op1_13_in29 = reg_0653;
    79: op1_13_in29 = reg_0399;
    80: op1_13_in29 = reg_0585;
    83: op1_13_in29 = reg_0089;
    84: op1_13_in29 = reg_0600;
    85: op1_13_in29 = reg_0063;
    87: op1_13_in29 = reg_0347;
    89: op1_13_in29 = reg_0592;
    90: op1_13_in29 = reg_0235;
    91: op1_13_in29 = reg_0751;
    92: op1_13_in29 = reg_0334;
    93: op1_13_in29 = reg_0711;
    94: op1_13_in29 = reg_0762;
    95: op1_13_in29 = reg_0289;
    default: op1_13_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_13_inv29 = 1;
    7: op1_13_inv29 = 1;
    8: op1_13_inv29 = 1;
    9: op1_13_inv29 = 1;
    10: op1_13_inv29 = 1;
    11: op1_13_inv29 = 1;
    12: op1_13_inv29 = 1;
    18: op1_13_inv29 = 1;
    20: op1_13_inv29 = 1;
    23: op1_13_inv29 = 1;
    24: op1_13_inv29 = 1;
    27: op1_13_inv29 = 1;
    29: op1_13_inv29 = 1;
    30: op1_13_inv29 = 1;
    31: op1_13_inv29 = 1;
    32: op1_13_inv29 = 1;
    33: op1_13_inv29 = 1;
    36: op1_13_inv29 = 1;
    37: op1_13_inv29 = 1;
    38: op1_13_inv29 = 1;
    45: op1_13_inv29 = 1;
    46: op1_13_inv29 = 1;
    47: op1_13_inv29 = 1;
    49: op1_13_inv29 = 1;
    54: op1_13_inv29 = 1;
    55: op1_13_inv29 = 1;
    57: op1_13_inv29 = 1;
    61: op1_13_inv29 = 1;
    63: op1_13_inv29 = 1;
    66: op1_13_inv29 = 1;
    67: op1_13_inv29 = 1;
    69: op1_13_inv29 = 1;
    70: op1_13_inv29 = 1;
    71: op1_13_inv29 = 1;
    72: op1_13_inv29 = 1;
    73: op1_13_inv29 = 1;
    77: op1_13_inv29 = 1;
    78: op1_13_inv29 = 1;
    79: op1_13_inv29 = 1;
    83: op1_13_inv29 = 1;
    85: op1_13_inv29 = 1;
    87: op1_13_inv29 = 1;
    89: op1_13_inv29 = 1;
    90: op1_13_inv29 = 1;
    93: op1_13_inv29 = 1;
    95: op1_13_inv29 = 1;
    default: op1_13_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_13_in30 = reg_0434;
    5: op1_13_in30 = reg_0151;
    6: op1_13_in30 = reg_0225;
    7: op1_13_in30 = imem03_in[87:84];
    8: op1_13_in30 = reg_0419;
    9: op1_13_in30 = reg_0143;
    10: op1_13_in30 = reg_0115;
    11: op1_13_in30 = imem04_in[111:108];
    12: op1_13_in30 = reg_0216;
    13: op1_13_in30 = reg_0587;
    14: op1_13_in30 = reg_0298;
    15: op1_13_in30 = reg_0183;
    16: op1_13_in30 = reg_0237;
    18: op1_13_in30 = reg_0248;
    20: op1_13_in30 = imem03_in[63:60];
    48: op1_13_in30 = imem03_in[63:60];
    21: op1_13_in30 = imem05_in[119:116];
    22: op1_13_in30 = reg_0448;
    23: op1_13_in30 = reg_0367;
    24: op1_13_in30 = reg_0418;
    25: op1_13_in30 = reg_0088;
    26: op1_13_in30 = reg_0501;
    27: op1_13_in30 = reg_0108;
    28: op1_13_in30 = reg_0140;
    29: op1_13_in30 = imem07_in[55:52];
    30: op1_13_in30 = imem03_in[23:20];
    31: op1_13_in30 = reg_0534;
    32: op1_13_in30 = imem05_in[83:80];
    33: op1_13_in30 = reg_0645;
    78: op1_13_in30 = reg_0645;
    34: op1_13_in30 = imem03_in[75:72];
    35: op1_13_in30 = imem03_in[127:124];
    36: op1_13_in30 = reg_0486;
    37: op1_13_in30 = reg_0043;
    38: op1_13_in30 = reg_0185;
    39: op1_13_in30 = reg_0174;
    41: op1_13_in30 = reg_0397;
    42: op1_13_in30 = reg_0145;
    43: op1_13_in30 = imem07_in[71:68];
    44: op1_13_in30 = reg_0519;
    45: op1_13_in30 = reg_0556;
    46: op1_13_in30 = reg_0778;
    47: op1_13_in30 = reg_0122;
    49: op1_13_in30 = reg_0603;
    51: op1_13_in30 = reg_0612;
    54: op1_13_in30 = reg_0669;
    55: op1_13_in30 = reg_0498;
    56: op1_13_in30 = imem03_in[47:44];
    57: op1_13_in30 = reg_0592;
    58: op1_13_in30 = imem04_in[103:100];
    59: op1_13_in30 = imem03_in[67:64];
    60: op1_13_in30 = reg_0062;
    61: op1_13_in30 = reg_0173;
    62: op1_13_in30 = reg_0054;
    63: op1_13_in30 = reg_0772;
    64: op1_13_in30 = reg_0243;
    65: op1_13_in30 = imem03_in[51:48];
    66: op1_13_in30 = imem02_in[11:8];
    67: op1_13_in30 = reg_0369;
    69: op1_13_in30 = reg_0509;
    70: op1_13_in30 = reg_0021;
    71: op1_13_in30 = reg_0118;
    72: op1_13_in30 = reg_0338;
    73: op1_13_in30 = reg_0808;
    74: op1_13_in30 = reg_0078;
    75: op1_13_in30 = reg_0625;
    77: op1_13_in30 = reg_0130;
    79: op1_13_in30 = reg_0595;
    84: op1_13_in30 = reg_0595;
    80: op1_13_in30 = reg_0065;
    81: op1_13_in30 = reg_0120;
    83: op1_13_in30 = reg_0116;
    85: op1_13_in30 = reg_0582;
    87: op1_13_in30 = imem03_in[31:28];
    89: op1_13_in30 = reg_0121;
    90: op1_13_in30 = reg_0506;
    91: op1_13_in30 = reg_0399;
    92: op1_13_in30 = reg_0266;
    93: op1_13_in30 = reg_0724;
    94: op1_13_in30 = reg_0409;
    95: op1_13_in30 = reg_0299;
    default: op1_13_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_13_inv30 = 1;
    7: op1_13_inv30 = 1;
    8: op1_13_inv30 = 1;
    9: op1_13_inv30 = 1;
    11: op1_13_inv30 = 1;
    12: op1_13_inv30 = 1;
    13: op1_13_inv30 = 1;
    16: op1_13_inv30 = 1;
    18: op1_13_inv30 = 1;
    20: op1_13_inv30 = 1;
    21: op1_13_inv30 = 1;
    23: op1_13_inv30 = 1;
    24: op1_13_inv30 = 1;
    25: op1_13_inv30 = 1;
    26: op1_13_inv30 = 1;
    28: op1_13_inv30 = 1;
    29: op1_13_inv30 = 1;
    31: op1_13_inv30 = 1;
    33: op1_13_inv30 = 1;
    34: op1_13_inv30 = 1;
    37: op1_13_inv30 = 1;
    38: op1_13_inv30 = 1;
    39: op1_13_inv30 = 1;
    42: op1_13_inv30 = 1;
    43: op1_13_inv30 = 1;
    44: op1_13_inv30 = 1;
    46: op1_13_inv30 = 1;
    47: op1_13_inv30 = 1;
    58: op1_13_inv30 = 1;
    59: op1_13_inv30 = 1;
    62: op1_13_inv30 = 1;
    64: op1_13_inv30 = 1;
    65: op1_13_inv30 = 1;
    67: op1_13_inv30 = 1;
    72: op1_13_inv30 = 1;
    74: op1_13_inv30 = 1;
    75: op1_13_inv30 = 1;
    77: op1_13_inv30 = 1;
    79: op1_13_inv30 = 1;
    80: op1_13_inv30 = 1;
    81: op1_13_inv30 = 1;
    83: op1_13_inv30 = 1;
    84: op1_13_inv30 = 1;
    85: op1_13_inv30 = 1;
    87: op1_13_inv30 = 1;
    89: op1_13_inv30 = 1;
    91: op1_13_inv30 = 1;
    92: op1_13_inv30 = 1;
    default: op1_13_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_13_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_13_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in00 = imem00_in[3:0];
    19: op1_14_in00 = imem00_in[3:0];
    22: op1_14_in00 = imem00_in[3:0];
    76: op1_14_in00 = imem00_in[3:0];
    5: op1_14_in00 = reg_0142;
    6: op1_14_in00 = reg_0112;
    7: op1_14_in00 = imem03_in[103:100];
    8: op1_14_in00 = imem00_in[7:4];
    82: op1_14_in00 = imem00_in[7:4];
    9: op1_14_in00 = reg_0130;
    10: op1_14_in00 = reg_0117;
    11: op1_14_in00 = imem04_in[119:116];
    12: op1_14_in00 = reg_0243;
    13: op1_14_in00 = reg_0591;
    72: op1_14_in00 = reg_0591;
    14: op1_14_in00 = reg_0061;
    15: op1_14_in00 = imem00_in[27:24];
    16: op1_14_in00 = reg_0504;
    17: op1_14_in00 = imem00_in[23:20];
    18: op1_14_in00 = reg_0237;
    20: op1_14_in00 = imem03_in[99:96];
    21: op1_14_in00 = reg_0488;
    23: op1_14_in00 = reg_0033;
    24: op1_14_in00 = imem00_in[39:36];
    86: op1_14_in00 = imem00_in[39:36];
    25: op1_14_in00 = reg_0555;
    26: op1_14_in00 = reg_0824;
    3: op1_14_in00 = imem07_in[95:92];
    1: op1_14_in00 = imem07_in[95:92];
    27: op1_14_in00 = reg_0114;
    28: op1_14_in00 = reg_0131;
    29: op1_14_in00 = imem00_in[79:76];
    30: op1_14_in00 = imem03_in[67:64];
    65: op1_14_in00 = imem03_in[67:64];
    31: op1_14_in00 = reg_0293;
    32: op1_14_in00 = imem05_in[119:116];
    2: op1_14_in00 = imem07_in[15:12];
    33: op1_14_in00 = reg_0662;
    34: op1_14_in00 = imem03_in[111:108];
    35: op1_14_in00 = reg_0592;
    36: op1_14_in00 = reg_0736;
    37: op1_14_in00 = reg_0054;
    38: op1_14_in00 = reg_0157;
    39: op1_14_in00 = reg_0175;
    40: op1_14_in00 = imem00_in[11:8];
    52: op1_14_in00 = imem00_in[11:8];
    53: op1_14_in00 = imem00_in[11:8];
    41: op1_14_in00 = reg_0000;
    42: op1_14_in00 = reg_0139;
    43: op1_14_in00 = imem07_in[79:76];
    44: op1_14_in00 = reg_0563;
    45: op1_14_in00 = reg_0631;
    46: op1_14_in00 = reg_0621;
    47: op1_14_in00 = reg_0111;
    48: op1_14_in00 = imem03_in[95:92];
    49: op1_14_in00 = reg_0506;
    50: op1_14_in00 = imem00_in[35:32];
    51: op1_14_in00 = reg_0331;
    54: op1_14_in00 = reg_0671;
    55: op1_14_in00 = imem03_in[11:8];
    56: op1_14_in00 = imem03_in[59:56];
    57: op1_14_in00 = reg_0672;
    81: op1_14_in00 = reg_0672;
    58: op1_14_in00 = imem05_in[11:8];
    59: op1_14_in00 = imem03_in[83:80];
    60: op1_14_in00 = reg_0687;
    61: op1_14_in00 = reg_0171;
    62: op1_14_in00 = reg_0567;
    63: op1_14_in00 = reg_0663;
    64: op1_14_in00 = reg_0105;
    66: op1_14_in00 = imem02_in[15:12];
    67: op1_14_in00 = reg_0630;
    68: op1_14_in00 = imem00_in[19:16];
    69: op1_14_in00 = imem03_in[3:0];
    70: op1_14_in00 = reg_0304;
    71: op1_14_in00 = reg_0670;
    73: op1_14_in00 = reg_0805;
    74: op1_14_in00 = reg_0069;
    75: op1_14_in00 = reg_0115;
    77: op1_14_in00 = reg_0760;
    78: op1_14_in00 = reg_0294;
    79: op1_14_in00 = reg_0751;
    80: op1_14_in00 = reg_0622;
    83: op1_14_in00 = reg_0141;
    84: op1_14_in00 = reg_0509;
    85: op1_14_in00 = reg_0317;
    87: op1_14_in00 = imem03_in[39:36];
    88: op1_14_in00 = imem00_in[55:52];
    89: op1_14_in00 = imem02_in[35:32];
    90: op1_14_in00 = reg_0119;
    91: op1_14_in00 = reg_0495;
    92: op1_14_in00 = reg_0053;
    93: op1_14_in00 = reg_0067;
    94: op1_14_in00 = reg_0619;
    95: op1_14_in00 = reg_0625;
    default: op1_14_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv00 = 1;
    9: op1_14_inv00 = 1;
    10: op1_14_inv00 = 1;
    12: op1_14_inv00 = 1;
    15: op1_14_inv00 = 1;
    16: op1_14_inv00 = 1;
    18: op1_14_inv00 = 1;
    20: op1_14_inv00 = 1;
    22: op1_14_inv00 = 1;
    23: op1_14_inv00 = 1;
    3: op1_14_inv00 = 1;
    27: op1_14_inv00 = 1;
    28: op1_14_inv00 = 1;
    31: op1_14_inv00 = 1;
    32: op1_14_inv00 = 1;
    33: op1_14_inv00 = 1;
    36: op1_14_inv00 = 1;
    37: op1_14_inv00 = 1;
    39: op1_14_inv00 = 1;
    43: op1_14_inv00 = 1;
    45: op1_14_inv00 = 1;
    47: op1_14_inv00 = 1;
    49: op1_14_inv00 = 1;
    52: op1_14_inv00 = 1;
    54: op1_14_inv00 = 1;
    57: op1_14_inv00 = 1;
    62: op1_14_inv00 = 1;
    64: op1_14_inv00 = 1;
    67: op1_14_inv00 = 1;
    69: op1_14_inv00 = 1;
    70: op1_14_inv00 = 1;
    73: op1_14_inv00 = 1;
    74: op1_14_inv00 = 1;
    75: op1_14_inv00 = 1;
    77: op1_14_inv00 = 1;
    82: op1_14_inv00 = 1;
    83: op1_14_inv00 = 1;
    84: op1_14_inv00 = 1;
    87: op1_14_inv00 = 1;
    88: op1_14_inv00 = 1;
    89: op1_14_inv00 = 1;
    91: op1_14_inv00 = 1;
    92: op1_14_inv00 = 1;
    93: op1_14_inv00 = 1;
    94: op1_14_inv00 = 1;
    95: op1_14_inv00 = 1;
    default: op1_14_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in01 = imem00_in[55:52];
    5: op1_14_in01 = reg_0141;
    6: op1_14_in01 = reg_0109;
    7: op1_14_in01 = imem03_in[119:116];
    8: op1_14_in01 = imem00_in[47:44];
    22: op1_14_in01 = imem00_in[47:44];
    9: op1_14_in01 = imem06_in[3:0];
    42: op1_14_in01 = imem06_in[3:0];
    10: op1_14_in01 = reg_0113;
    11: op1_14_in01 = reg_0545;
    12: op1_14_in01 = reg_0105;
    13: op1_14_in01 = reg_0563;
    14: op1_14_in01 = reg_0075;
    15: op1_14_in01 = imem00_in[31:28];
    16: op1_14_in01 = reg_0219;
    17: op1_14_in01 = imem00_in[51:48];
    50: op1_14_in01 = imem00_in[51:48];
    18: op1_14_in01 = reg_0245;
    19: op1_14_in01 = imem00_in[99:96];
    20: op1_14_in01 = reg_0573;
    21: op1_14_in01 = reg_0789;
    23: op1_14_in01 = reg_0753;
    24: op1_14_in01 = imem00_in[59:56];
    25: op1_14_in01 = reg_0057;
    26: op1_14_in01 = reg_0559;
    3: op1_14_in01 = reg_0441;
    27: op1_14_in01 = imem02_in[35:32];
    28: op1_14_in01 = reg_0144;
    29: op1_14_in01 = reg_0698;
    30: op1_14_in01 = imem03_in[87:84];
    56: op1_14_in01 = imem03_in[87:84];
    31: op1_14_in01 = reg_0290;
    32: op1_14_in01 = reg_0797;
    2: op1_14_in01 = imem07_in[71:68];
    33: op1_14_in01 = reg_0352;
    34: op1_14_in01 = imem03_in[123:120];
    48: op1_14_in01 = imem03_in[123:120];
    35: op1_14_in01 = reg_0750;
    72: op1_14_in01 = reg_0750;
    36: op1_14_in01 = reg_0737;
    37: op1_14_in01 = reg_0305;
    39: op1_14_in01 = reg_0179;
    40: op1_14_in01 = imem00_in[19:16];
    41: op1_14_in01 = reg_0012;
    43: op1_14_in01 = imem07_in[95:92];
    44: op1_14_in01 = reg_0487;
    45: op1_14_in01 = reg_0503;
    46: op1_14_in01 = imem07_in[63:60];
    47: op1_14_in01 = reg_0100;
    49: op1_14_in01 = reg_0424;
    51: op1_14_in01 = reg_0405;
    52: op1_14_in01 = imem00_in[23:20];
    82: op1_14_in01 = imem00_in[23:20];
    53: op1_14_in01 = imem00_in[27:24];
    54: op1_14_in01 = reg_0676;
    90: op1_14_in01 = reg_0676;
    55: op1_14_in01 = imem03_in[27:24];
    57: op1_14_in01 = reg_0675;
    58: op1_14_in01 = imem05_in[31:28];
    59: op1_14_in01 = imem03_in[91:88];
    60: op1_14_in01 = reg_0640;
    62: op1_14_in01 = reg_0425;
    63: op1_14_in01 = reg_0820;
    64: op1_14_in01 = reg_0592;
    65: op1_14_in01 = reg_0063;
    66: op1_14_in01 = imem02_in[63:60];
    67: op1_14_in01 = reg_0613;
    68: op1_14_in01 = imem00_in[39:36];
    69: op1_14_in01 = imem03_in[15:12];
    70: op1_14_in01 = reg_0605;
    71: op1_14_in01 = reg_0108;
    73: op1_14_in01 = reg_0802;
    74: op1_14_in01 = reg_0774;
    75: op1_14_in01 = reg_0624;
    76: op1_14_in01 = imem00_in[7:4];
    77: op1_14_in01 = reg_0073;
    78: op1_14_in01 = reg_0506;
    79: op1_14_in01 = reg_0331;
    80: op1_14_in01 = reg_0069;
    81: op1_14_in01 = reg_0107;
    83: op1_14_in01 = reg_0185;
    84: op1_14_in01 = reg_0321;
    85: op1_14_in01 = reg_0604;
    86: op1_14_in01 = imem00_in[87:84];
    87: op1_14_in01 = imem03_in[43:40];
    88: op1_14_in01 = imem00_in[83:80];
    89: op1_14_in01 = reg_0541;
    91: op1_14_in01 = reg_0254;
    92: op1_14_in01 = reg_0434;
    93: op1_14_in01 = reg_0333;
    94: op1_14_in01 = reg_0238;
    95: op1_14_in01 = reg_0291;
    default: op1_14_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv01 = 1;
    6: op1_14_inv01 = 1;
    7: op1_14_inv01 = 1;
    9: op1_14_inv01 = 1;
    12: op1_14_inv01 = 1;
    13: op1_14_inv01 = 1;
    15: op1_14_inv01 = 1;
    16: op1_14_inv01 = 1;
    18: op1_14_inv01 = 1;
    25: op1_14_inv01 = 1;
    26: op1_14_inv01 = 1;
    27: op1_14_inv01 = 1;
    28: op1_14_inv01 = 1;
    31: op1_14_inv01 = 1;
    33: op1_14_inv01 = 1;
    34: op1_14_inv01 = 1;
    35: op1_14_inv01 = 1;
    36: op1_14_inv01 = 1;
    37: op1_14_inv01 = 1;
    39: op1_14_inv01 = 1;
    43: op1_14_inv01 = 1;
    44: op1_14_inv01 = 1;
    46: op1_14_inv01 = 1;
    47: op1_14_inv01 = 1;
    50: op1_14_inv01 = 1;
    51: op1_14_inv01 = 1;
    52: op1_14_inv01 = 1;
    53: op1_14_inv01 = 1;
    55: op1_14_inv01 = 1;
    56: op1_14_inv01 = 1;
    58: op1_14_inv01 = 1;
    59: op1_14_inv01 = 1;
    60: op1_14_inv01 = 1;
    65: op1_14_inv01 = 1;
    66: op1_14_inv01 = 1;
    69: op1_14_inv01 = 1;
    70: op1_14_inv01 = 1;
    71: op1_14_inv01 = 1;
    72: op1_14_inv01 = 1;
    73: op1_14_inv01 = 1;
    77: op1_14_inv01 = 1;
    80: op1_14_inv01 = 1;
    82: op1_14_inv01 = 1;
    85: op1_14_inv01 = 1;
    89: op1_14_inv01 = 1;
    93: op1_14_inv01 = 1;
    94: op1_14_inv01 = 1;
    default: op1_14_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in02 = imem00_in[91:88];
    50: op1_14_in02 = imem00_in[91:88];
    86: op1_14_in02 = imem00_in[91:88];
    88: op1_14_in02 = imem00_in[91:88];
    5: op1_14_in02 = reg_0137;
    6: op1_14_in02 = imem02_in[7:4];
    7: op1_14_in02 = reg_0586;
    8: op1_14_in02 = imem00_in[51:48];
    9: op1_14_in02 = imem06_in[7:4];
    10: op1_14_in02 = imem02_in[19:16];
    54: op1_14_in02 = imem02_in[19:16];
    11: op1_14_in02 = reg_0557;
    12: op1_14_in02 = reg_0124;
    13: op1_14_in02 = reg_0373;
    14: op1_14_in02 = imem05_in[43:40];
    15: op1_14_in02 = imem00_in[43:40];
    16: op1_14_in02 = reg_0102;
    17: op1_14_in02 = imem00_in[95:92];
    18: op1_14_in02 = reg_0105;
    19: op1_14_in02 = imem00_in[103:100];
    20: op1_14_in02 = reg_0583;
    34: op1_14_in02 = reg_0583;
    21: op1_14_in02 = reg_0491;
    22: op1_14_in02 = imem00_in[87:84];
    23: op1_14_in02 = reg_0040;
    24: op1_14_in02 = imem00_in[83:80];
    25: op1_14_in02 = reg_0536;
    26: op1_14_in02 = reg_0233;
    3: op1_14_in02 = reg_0419;
    27: op1_14_in02 = imem02_in[47:44];
    28: op1_14_in02 = reg_0381;
    29: op1_14_in02 = reg_0690;
    30: op1_14_in02 = imem03_in[103:100];
    31: op1_14_in02 = reg_0291;
    32: op1_14_in02 = reg_0489;
    2: op1_14_in02 = imem07_in[87:84];
    33: op1_14_in02 = reg_0349;
    95: op1_14_in02 = reg_0349;
    35: op1_14_in02 = reg_0589;
    36: op1_14_in02 = reg_0084;
    37: op1_14_in02 = reg_0294;
    39: op1_14_in02 = reg_0162;
    40: op1_14_in02 = imem00_in[67:64];
    41: op1_14_in02 = reg_0806;
    42: op1_14_in02 = imem06_in[59:56];
    43: op1_14_in02 = imem07_in[107:104];
    46: op1_14_in02 = imem07_in[107:104];
    44: op1_14_in02 = reg_0418;
    45: op1_14_in02 = reg_0050;
    47: op1_14_in02 = reg_0115;
    48: op1_14_in02 = imem03_in[127:124];
    49: op1_14_in02 = reg_0219;
    62: op1_14_in02 = reg_0219;
    51: op1_14_in02 = reg_0821;
    52: op1_14_in02 = imem00_in[35:32];
    53: op1_14_in02 = imem00_in[39:36];
    55: op1_14_in02 = imem03_in[55:52];
    56: op1_14_in02 = imem03_in[91:88];
    57: op1_14_in02 = imem02_in[15:12];
    58: op1_14_in02 = imem05_in[55:52];
    59: op1_14_in02 = imem03_in[107:104];
    60: op1_14_in02 = reg_0109;
    63: op1_14_in02 = reg_0649;
    64: op1_14_in02 = reg_0660;
    65: op1_14_in02 = reg_0604;
    66: op1_14_in02 = imem02_in[103:100];
    67: op1_14_in02 = reg_0816;
    68: op1_14_in02 = imem00_in[55:52];
    69: op1_14_in02 = imem03_in[39:36];
    70: op1_14_in02 = reg_0409;
    71: op1_14_in02 = reg_0671;
    72: op1_14_in02 = reg_0318;
    73: op1_14_in02 = reg_0016;
    74: op1_14_in02 = reg_0416;
    75: op1_14_in02 = reg_0817;
    76: op1_14_in02 = imem00_in[27:24];
    77: op1_14_in02 = reg_0106;
    78: op1_14_in02 = reg_0073;
    79: op1_14_in02 = reg_0395;
    80: op1_14_in02 = reg_0513;
    81: op1_14_in02 = reg_0678;
    82: op1_14_in02 = imem00_in[31:28];
    84: op1_14_in02 = reg_0417;
    85: op1_14_in02 = reg_0338;
    87: op1_14_in02 = imem03_in[79:76];
    89: op1_14_in02 = reg_0530;
    90: op1_14_in02 = imem02_in[23:20];
    91: op1_14_in02 = reg_0547;
    92: op1_14_in02 = reg_0267;
    93: op1_14_in02 = reg_0116;
    94: op1_14_in02 = reg_0618;
    default: op1_14_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv02 = 1;
    8: op1_14_inv02 = 1;
    10: op1_14_inv02 = 1;
    11: op1_14_inv02 = 1;
    12: op1_14_inv02 = 1;
    13: op1_14_inv02 = 1;
    15: op1_14_inv02 = 1;
    16: op1_14_inv02 = 1;
    17: op1_14_inv02 = 1;
    18: op1_14_inv02 = 1;
    19: op1_14_inv02 = 1;
    21: op1_14_inv02 = 1;
    22: op1_14_inv02 = 1;
    25: op1_14_inv02 = 1;
    26: op1_14_inv02 = 1;
    3: op1_14_inv02 = 1;
    27: op1_14_inv02 = 1;
    29: op1_14_inv02 = 1;
    30: op1_14_inv02 = 1;
    31: op1_14_inv02 = 1;
    2: op1_14_inv02 = 1;
    35: op1_14_inv02 = 1;
    37: op1_14_inv02 = 1;
    40: op1_14_inv02 = 1;
    41: op1_14_inv02 = 1;
    42: op1_14_inv02 = 1;
    44: op1_14_inv02 = 1;
    45: op1_14_inv02 = 1;
    46: op1_14_inv02 = 1;
    49: op1_14_inv02 = 1;
    51: op1_14_inv02 = 1;
    53: op1_14_inv02 = 1;
    54: op1_14_inv02 = 1;
    56: op1_14_inv02 = 1;
    58: op1_14_inv02 = 1;
    59: op1_14_inv02 = 1;
    60: op1_14_inv02 = 1;
    62: op1_14_inv02 = 1;
    64: op1_14_inv02 = 1;
    65: op1_14_inv02 = 1;
    66: op1_14_inv02 = 1;
    67: op1_14_inv02 = 1;
    71: op1_14_inv02 = 1;
    72: op1_14_inv02 = 1;
    73: op1_14_inv02 = 1;
    76: op1_14_inv02 = 1;
    77: op1_14_inv02 = 1;
    79: op1_14_inv02 = 1;
    81: op1_14_inv02 = 1;
    82: op1_14_inv02 = 1;
    84: op1_14_inv02 = 1;
    85: op1_14_inv02 = 1;
    89: op1_14_inv02 = 1;
    90: op1_14_inv02 = 1;
    91: op1_14_inv02 = 1;
    93: op1_14_inv02 = 1;
    default: op1_14_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in03 = reg_0670;
    5: op1_14_in03 = imem06_in[35:32];
    6: op1_14_in03 = imem02_in[11:8];
    7: op1_14_in03 = reg_0573;
    8: op1_14_in03 = imem00_in[55:52];
    15: op1_14_in03 = imem00_in[55:52];
    9: op1_14_in03 = imem06_in[11:8];
    10: op1_14_in03 = reg_0655;
    11: op1_14_in03 = reg_0552;
    12: op1_14_in03 = reg_0111;
    13: op1_14_in03 = reg_0322;
    14: op1_14_in03 = imem05_in[51:48];
    16: op1_14_in03 = imem02_in[39:36];
    57: op1_14_in03 = imem02_in[39:36];
    17: op1_14_in03 = reg_0684;
    18: op1_14_in03 = reg_0107;
    19: op1_14_in03 = imem00_in[127:124];
    20: op1_14_in03 = reg_0568;
    84: op1_14_in03 = reg_0568;
    21: op1_14_in03 = reg_0795;
    22: op1_14_in03 = reg_0695;
    86: op1_14_in03 = reg_0695;
    23: op1_14_in03 = reg_0037;
    24: op1_14_in03 = imem00_in[99:96];
    50: op1_14_in03 = imem00_in[99:96];
    25: op1_14_in03 = reg_0500;
    26: op1_14_in03 = reg_0511;
    3: op1_14_in03 = reg_0434;
    27: op1_14_in03 = imem02_in[99:96];
    28: op1_14_in03 = reg_0371;
    29: op1_14_in03 = reg_0668;
    30: op1_14_in03 = imem03_in[127:124];
    87: op1_14_in03 = imem03_in[127:124];
    31: op1_14_in03 = reg_0292;
    32: op1_14_in03 = reg_0741;
    2: op1_14_in03 = imem07_in[107:104];
    33: op1_14_in03 = reg_0359;
    34: op1_14_in03 = reg_0039;
    35: op1_14_in03 = reg_0585;
    36: op1_14_in03 = reg_0086;
    37: op1_14_in03 = reg_0297;
    39: op1_14_in03 = reg_0183;
    40: op1_14_in03 = imem00_in[75:72];
    41: op1_14_in03 = reg_0810;
    42: op1_14_in03 = imem06_in[83:80];
    43: op1_14_in03 = imem07_in[111:108];
    44: op1_14_in03 = reg_0306;
    45: op1_14_in03 = imem04_in[3:0];
    46: op1_14_in03 = imem07_in[123:120];
    47: op1_14_in03 = reg_0109;
    48: op1_14_in03 = reg_0566;
    49: op1_14_in03 = reg_0123;
    51: op1_14_in03 = reg_0270;
    52: op1_14_in03 = imem00_in[47:44];
    53: op1_14_in03 = imem00_in[47:44];
    54: op1_14_in03 = imem02_in[27:24];
    55: op1_14_in03 = imem03_in[99:96];
    56: op1_14_in03 = reg_0317;
    58: op1_14_in03 = reg_0112;
    59: op1_14_in03 = reg_0589;
    60: op1_14_in03 = reg_0484;
    62: op1_14_in03 = reg_0505;
    63: op1_14_in03 = reg_0100;
    64: op1_14_in03 = reg_0106;
    65: op1_14_in03 = reg_0493;
    66: op1_14_in03 = imem02_in[111:108];
    67: op1_14_in03 = reg_0583;
    68: op1_14_in03 = imem00_in[71:68];
    69: op1_14_in03 = imem03_in[47:44];
    70: op1_14_in03 = reg_0578;
    71: op1_14_in03 = reg_0127;
    72: op1_14_in03 = reg_0395;
    73: op1_14_in03 = imem04_in[15:12];
    74: op1_14_in03 = imem05_in[35:32];
    75: op1_14_in03 = reg_0618;
    76: op1_14_in03 = imem00_in[35:32];
    77: op1_14_in03 = reg_0601;
    78: op1_14_in03 = reg_0126;
    79: op1_14_in03 = reg_0384;
    80: op1_14_in03 = reg_0233;
    81: op1_14_in03 = imem02_in[7:4];
    82: op1_14_in03 = imem00_in[43:40];
    85: op1_14_in03 = reg_0591;
    88: op1_14_in03 = imem00_in[115:112];
    89: op1_14_in03 = reg_0656;
    90: op1_14_in03 = imem02_in[35:32];
    91: op1_14_in03 = reg_0149;
    92: op1_14_in03 = reg_0066;
    93: op1_14_in03 = reg_0730;
    94: op1_14_in03 = reg_0293;
    95: op1_14_in03 = reg_0370;
    default: op1_14_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv03 = 1;
    7: op1_14_inv03 = 1;
    9: op1_14_inv03 = 1;
    12: op1_14_inv03 = 1;
    13: op1_14_inv03 = 1;
    14: op1_14_inv03 = 1;
    20: op1_14_inv03 = 1;
    21: op1_14_inv03 = 1;
    24: op1_14_inv03 = 1;
    25: op1_14_inv03 = 1;
    3: op1_14_inv03 = 1;
    27: op1_14_inv03 = 1;
    28: op1_14_inv03 = 1;
    29: op1_14_inv03 = 1;
    2: op1_14_inv03 = 1;
    33: op1_14_inv03 = 1;
    35: op1_14_inv03 = 1;
    36: op1_14_inv03 = 1;
    42: op1_14_inv03 = 1;
    43: op1_14_inv03 = 1;
    45: op1_14_inv03 = 1;
    50: op1_14_inv03 = 1;
    52: op1_14_inv03 = 1;
    55: op1_14_inv03 = 1;
    56: op1_14_inv03 = 1;
    60: op1_14_inv03 = 1;
    66: op1_14_inv03 = 1;
    67: op1_14_inv03 = 1;
    71: op1_14_inv03 = 1;
    73: op1_14_inv03 = 1;
    74: op1_14_inv03 = 1;
    75: op1_14_inv03 = 1;
    76: op1_14_inv03 = 1;
    77: op1_14_inv03 = 1;
    78: op1_14_inv03 = 1;
    85: op1_14_inv03 = 1;
    87: op1_14_inv03 = 1;
    88: op1_14_inv03 = 1;
    90: op1_14_inv03 = 1;
    91: op1_14_inv03 = 1;
    93: op1_14_inv03 = 1;
    default: op1_14_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in04 = reg_0679;
    5: op1_14_in04 = imem06_in[63:60];
    9: op1_14_in04 = imem06_in[63:60];
    6: op1_14_in04 = imem02_in[51:48];
    7: op1_14_in04 = reg_0569;
    8: op1_14_in04 = imem00_in[59:56];
    15: op1_14_in04 = imem00_in[59:56];
    10: op1_14_in04 = reg_0653;
    11: op1_14_in04 = reg_0542;
    12: op1_14_in04 = reg_0125;
    13: op1_14_in04 = reg_0376;
    14: op1_14_in04 = imem05_in[75:72];
    16: op1_14_in04 = imem02_in[43:40];
    17: op1_14_in04 = reg_0691;
    18: op1_14_in04 = imem02_in[23:20];
    19: op1_14_in04 = reg_0683;
    20: op1_14_in04 = reg_0370;
    21: op1_14_in04 = reg_0780;
    22: op1_14_in04 = reg_0690;
    23: op1_14_in04 = reg_0750;
    65: op1_14_in04 = reg_0750;
    24: op1_14_in04 = imem00_in[123:120];
    25: op1_14_in04 = reg_0305;
    26: op1_14_in04 = reg_0242;
    3: op1_14_in04 = reg_0444;
    27: op1_14_in04 = imem02_in[103:100];
    28: op1_14_in04 = reg_0375;
    29: op1_14_in04 = reg_0675;
    30: op1_14_in04 = reg_0398;
    31: op1_14_in04 = reg_0266;
    32: op1_14_in04 = reg_0085;
    2: op1_14_in04 = imem07_in[115:112];
    33: op1_14_in04 = reg_0342;
    34: op1_14_in04 = reg_0591;
    35: op1_14_in04 = reg_0593;
    36: op1_14_in04 = reg_0156;
    37: op1_14_in04 = reg_0298;
    39: op1_14_in04 = reg_0166;
    40: op1_14_in04 = imem00_in[87:84];
    53: op1_14_in04 = imem00_in[87:84];
    41: op1_14_in04 = reg_0268;
    42: op1_14_in04 = imem06_in[95:92];
    43: op1_14_in04 = reg_0720;
    44: op1_14_in04 = reg_0217;
    45: op1_14_in04 = imem04_in[43:40];
    46: op1_14_in04 = reg_0704;
    47: op1_14_in04 = imem02_in[7:4];
    48: op1_14_in04 = reg_0583;
    49: op1_14_in04 = reg_0111;
    50: op1_14_in04 = reg_0693;
    51: op1_14_in04 = reg_0319;
    52: op1_14_in04 = imem00_in[99:96];
    54: op1_14_in04 = imem02_in[47:44];
    55: op1_14_in04 = imem03_in[111:108];
    56: op1_14_in04 = reg_0599;
    57: op1_14_in04 = imem02_in[63:60];
    58: op1_14_in04 = reg_0278;
    59: op1_14_in04 = reg_0338;
    60: op1_14_in04 = reg_0040;
    62: op1_14_in04 = reg_0123;
    63: op1_14_in04 = reg_0778;
    64: op1_14_in04 = reg_0107;
    66: op1_14_in04 = reg_0501;
    67: op1_14_in04 = reg_0035;
    68: op1_14_in04 = imem00_in[119:116];
    88: op1_14_in04 = imem00_in[119:116];
    69: op1_14_in04 = imem03_in[51:48];
    70: op1_14_in04 = reg_0408;
    71: op1_14_in04 = reg_0674;
    72: op1_14_in04 = reg_0755;
    79: op1_14_in04 = reg_0755;
    73: op1_14_in04 = imem04_in[19:16];
    74: op1_14_in04 = imem05_in[55:52];
    75: op1_14_in04 = reg_0628;
    76: op1_14_in04 = imem00_in[47:44];
    77: op1_14_in04 = imem02_in[31:28];
    78: op1_14_in04 = imem02_in[27:24];
    80: op1_14_in04 = reg_0644;
    81: op1_14_in04 = imem02_in[39:36];
    82: op1_14_in04 = imem00_in[63:60];
    84: op1_14_in04 = reg_0368;
    85: op1_14_in04 = reg_0329;
    86: op1_14_in04 = reg_0682;
    87: op1_14_in04 = reg_0028;
    89: op1_14_in04 = reg_0639;
    90: op1_14_in04 = imem02_in[99:96];
    91: op1_14_in04 = reg_0783;
    92: op1_14_in04 = reg_0228;
    93: op1_14_in04 = reg_0426;
    94: op1_14_in04 = reg_0401;
    95: op1_14_in04 = reg_0618;
    default: op1_14_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv04 = 1;
    5: op1_14_inv04 = 1;
    6: op1_14_inv04 = 1;
    9: op1_14_inv04 = 1;
    11: op1_14_inv04 = 1;
    12: op1_14_inv04 = 1;
    14: op1_14_inv04 = 1;
    16: op1_14_inv04 = 1;
    17: op1_14_inv04 = 1;
    18: op1_14_inv04 = 1;
    19: op1_14_inv04 = 1;
    20: op1_14_inv04 = 1;
    21: op1_14_inv04 = 1;
    24: op1_14_inv04 = 1;
    29: op1_14_inv04 = 1;
    36: op1_14_inv04 = 1;
    37: op1_14_inv04 = 1;
    39: op1_14_inv04 = 1;
    40: op1_14_inv04 = 1;
    41: op1_14_inv04 = 1;
    43: op1_14_inv04 = 1;
    45: op1_14_inv04 = 1;
    47: op1_14_inv04 = 1;
    49: op1_14_inv04 = 1;
    51: op1_14_inv04 = 1;
    54: op1_14_inv04 = 1;
    58: op1_14_inv04 = 1;
    59: op1_14_inv04 = 1;
    60: op1_14_inv04 = 1;
    62: op1_14_inv04 = 1;
    63: op1_14_inv04 = 1;
    64: op1_14_inv04 = 1;
    65: op1_14_inv04 = 1;
    68: op1_14_inv04 = 1;
    70: op1_14_inv04 = 1;
    71: op1_14_inv04 = 1;
    75: op1_14_inv04 = 1;
    76: op1_14_inv04 = 1;
    77: op1_14_inv04 = 1;
    78: op1_14_inv04 = 1;
    79: op1_14_inv04 = 1;
    81: op1_14_inv04 = 1;
    84: op1_14_inv04 = 1;
    85: op1_14_inv04 = 1;
    86: op1_14_inv04 = 1;
    87: op1_14_inv04 = 1;
    90: op1_14_inv04 = 1;
    92: op1_14_inv04 = 1;
    93: op1_14_inv04 = 1;
    94: op1_14_inv04 = 1;
    95: op1_14_inv04 = 1;
    default: op1_14_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in05 = reg_0465;
    5: op1_14_in05 = imem06_in[67:64];
    6: op1_14_in05 = imem02_in[79:76];
    7: op1_14_in05 = reg_0591;
    8: op1_14_in05 = imem00_in[115:112];
    40: op1_14_in05 = imem00_in[115:112];
    9: op1_14_in05 = imem06_in[87:84];
    10: op1_14_in05 = reg_0661;
    11: op1_14_in05 = reg_0548;
    12: op1_14_in05 = reg_0116;
    49: op1_14_in05 = reg_0116;
    13: op1_14_in05 = reg_0374;
    14: op1_14_in05 = imem05_in[103:100];
    15: op1_14_in05 = imem00_in[91:88];
    16: op1_14_in05 = imem02_in[75:72];
    17: op1_14_in05 = reg_0674;
    18: op1_14_in05 = imem02_in[47:44];
    77: op1_14_in05 = imem02_in[47:44];
    19: op1_14_in05 = reg_0694;
    20: op1_14_in05 = reg_0362;
    21: op1_14_in05 = reg_0485;
    22: op1_14_in05 = reg_0481;
    23: op1_14_in05 = reg_0029;
    24: op1_14_in05 = reg_0693;
    25: op1_14_in05 = reg_0273;
    26: op1_14_in05 = reg_0245;
    3: op1_14_in05 = reg_0181;
    2: op1_14_in05 = reg_0181;
    27: op1_14_in05 = reg_0647;
    28: op1_14_in05 = reg_0339;
    29: op1_14_in05 = reg_0450;
    30: op1_14_in05 = reg_0747;
    31: op1_14_in05 = reg_0070;
    32: op1_14_in05 = reg_0733;
    33: op1_14_in05 = reg_0322;
    34: op1_14_in05 = reg_0584;
    35: op1_14_in05 = reg_0580;
    36: op1_14_in05 = reg_0130;
    37: op1_14_in05 = reg_0299;
    39: op1_14_in05 = reg_0185;
    41: op1_14_in05 = reg_0553;
    42: op1_14_in05 = reg_0613;
    43: op1_14_in05 = reg_0725;
    44: op1_14_in05 = reg_0220;
    45: op1_14_in05 = imem04_in[59:56];
    46: op1_14_in05 = reg_0730;
    47: op1_14_in05 = imem02_in[19:16];
    48: op1_14_in05 = reg_0565;
    50: op1_14_in05 = reg_0684;
    51: op1_14_in05 = reg_0764;
    52: op1_14_in05 = imem00_in[111:108];
    53: op1_14_in05 = imem00_in[107:104];
    54: op1_14_in05 = imem02_in[55:52];
    55: op1_14_in05 = reg_0559;
    56: op1_14_in05 = reg_0338;
    57: op1_14_in05 = imem02_in[115:112];
    58: op1_14_in05 = reg_0782;
    59: op1_14_in05 = reg_0319;
    60: op1_14_in05 = reg_0785;
    62: op1_14_in05 = reg_0660;
    63: op1_14_in05 = reg_0737;
    64: op1_14_in05 = imem02_in[23:20];
    65: op1_14_in05 = reg_0350;
    66: op1_14_in05 = reg_0045;
    67: op1_14_in05 = reg_0794;
    68: op1_14_in05 = imem00_in[123:120];
    69: op1_14_in05 = imem03_in[99:96];
    70: op1_14_in05 = reg_0270;
    71: op1_14_in05 = reg_0133;
    72: op1_14_in05 = reg_0572;
    73: op1_14_in05 = imem04_in[31:28];
    74: op1_14_in05 = imem05_in[59:56];
    75: op1_14_in05 = reg_0242;
    76: op1_14_in05 = imem00_in[75:72];
    78: op1_14_in05 = imem02_in[35:32];
    79: op1_14_in05 = reg_0403;
    80: op1_14_in05 = imem05_in[19:16];
    81: op1_14_in05 = imem02_in[51:48];
    82: op1_14_in05 = imem00_in[71:68];
    84: op1_14_in05 = reg_0569;
    85: op1_14_in05 = reg_0399;
    86: op1_14_in05 = reg_0685;
    87: op1_14_in05 = reg_0417;
    88: op1_14_in05 = reg_0634;
    89: op1_14_in05 = reg_0087;
    90: op1_14_in05 = reg_0081;
    91: op1_14_in05 = reg_0828;
    92: op1_14_in05 = reg_0100;
    93: op1_14_in05 = reg_0099;
    94: op1_14_in05 = reg_0276;
    95: op1_14_in05 = reg_0766;
    default: op1_14_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv05 = 1;
    5: op1_14_inv05 = 1;
    6: op1_14_inv05 = 1;
    10: op1_14_inv05 = 1;
    11: op1_14_inv05 = 1;
    12: op1_14_inv05 = 1;
    16: op1_14_inv05 = 1;
    18: op1_14_inv05 = 1;
    20: op1_14_inv05 = 1;
    21: op1_14_inv05 = 1;
    29: op1_14_inv05 = 1;
    30: op1_14_inv05 = 1;
    31: op1_14_inv05 = 1;
    34: op1_14_inv05 = 1;
    35: op1_14_inv05 = 1;
    37: op1_14_inv05 = 1;
    39: op1_14_inv05 = 1;
    41: op1_14_inv05 = 1;
    45: op1_14_inv05 = 1;
    47: op1_14_inv05 = 1;
    48: op1_14_inv05 = 1;
    49: op1_14_inv05 = 1;
    50: op1_14_inv05 = 1;
    52: op1_14_inv05 = 1;
    53: op1_14_inv05 = 1;
    54: op1_14_inv05 = 1;
    55: op1_14_inv05 = 1;
    57: op1_14_inv05 = 1;
    58: op1_14_inv05 = 1;
    60: op1_14_inv05 = 1;
    64: op1_14_inv05 = 1;
    66: op1_14_inv05 = 1;
    69: op1_14_inv05 = 1;
    70: op1_14_inv05 = 1;
    71: op1_14_inv05 = 1;
    74: op1_14_inv05 = 1;
    78: op1_14_inv05 = 1;
    80: op1_14_inv05 = 1;
    84: op1_14_inv05 = 1;
    88: op1_14_inv05 = 1;
    90: op1_14_inv05 = 1;
    default: op1_14_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in06 = reg_0455;
    5: op1_14_in06 = imem06_in[83:80];
    6: op1_14_in06 = imem02_in[99:96];
    18: op1_14_in06 = imem02_in[99:96];
    7: op1_14_in06 = reg_0593;
    8: op1_14_in06 = imem00_in[119:116];
    9: op1_14_in06 = reg_0625;
    10: op1_14_in06 = reg_0640;
    27: op1_14_in06 = reg_0640;
    11: op1_14_in06 = reg_0549;
    12: op1_14_in06 = reg_0119;
    13: op1_14_in06 = reg_0389;
    30: op1_14_in06 = reg_0389;
    14: op1_14_in06 = reg_0781;
    15: op1_14_in06 = imem00_in[103:100];
    16: op1_14_in06 = imem02_in[87:84];
    47: op1_14_in06 = imem02_in[87:84];
    17: op1_14_in06 = reg_0699;
    19: op1_14_in06 = reg_0676;
    20: op1_14_in06 = reg_0398;
    21: op1_14_in06 = reg_0787;
    22: op1_14_in06 = reg_0471;
    23: op1_14_in06 = reg_0749;
    35: op1_14_in06 = reg_0749;
    24: op1_14_in06 = reg_0690;
    25: op1_14_in06 = reg_0294;
    26: op1_14_in06 = reg_0238;
    3: op1_14_in06 = reg_0182;
    28: op1_14_in06 = reg_0607;
    29: op1_14_in06 = reg_0464;
    31: op1_14_in06 = reg_0064;
    32: op1_14_in06 = reg_0282;
    2: op1_14_in06 = reg_0162;
    33: op1_14_in06 = reg_0518;
    34: op1_14_in06 = reg_0600;
    36: op1_14_in06 = reg_0813;
    37: op1_14_in06 = reg_0069;
    40: op1_14_in06 = imem00_in[123:120];
    41: op1_14_in06 = reg_0056;
    42: op1_14_in06 = reg_0608;
    43: op1_14_in06 = reg_0703;
    44: op1_14_in06 = reg_0505;
    45: op1_14_in06 = imem04_in[87:84];
    46: op1_14_in06 = reg_0731;
    48: op1_14_in06 = reg_0587;
    49: op1_14_in06 = reg_0104;
    50: op1_14_in06 = reg_0679;
    51: op1_14_in06 = reg_0576;
    52: op1_14_in06 = reg_0693;
    53: op1_14_in06 = reg_0695;
    54: op1_14_in06 = imem02_in[63:60];
    55: op1_14_in06 = reg_0750;
    56: op1_14_in06 = reg_0595;
    57: op1_14_in06 = reg_0337;
    58: op1_14_in06 = reg_0486;
    59: op1_14_in06 = reg_0318;
    60: op1_14_in06 = imem05_in[3:0];
    62: op1_14_in06 = reg_0040;
    63: op1_14_in06 = reg_0240;
    64: op1_14_in06 = imem02_in[35:32];
    65: op1_14_in06 = reg_0329;
    66: op1_14_in06 = reg_0275;
    67: op1_14_in06 = imem07_in[11:8];
    68: op1_14_in06 = reg_0682;
    69: op1_14_in06 = imem03_in[107:104];
    70: op1_14_in06 = reg_0375;
    71: op1_14_in06 = reg_0090;
    72: op1_14_in06 = reg_0372;
    87: op1_14_in06 = reg_0372;
    73: op1_14_in06 = imem04_in[39:36];
    74: op1_14_in06 = imem05_in[71:68];
    75: op1_14_in06 = reg_0031;
    76: op1_14_in06 = imem00_in[79:76];
    77: op1_14_in06 = imem02_in[119:116];
    78: op1_14_in06 = imem02_in[43:40];
    79: op1_14_in06 = reg_0562;
    80: op1_14_in06 = imem05_in[27:24];
    81: op1_14_in06 = imem02_in[67:64];
    82: op1_14_in06 = imem00_in[127:124];
    84: op1_14_in06 = reg_0807;
    85: op1_14_in06 = reg_0751;
    86: op1_14_in06 = reg_0684;
    88: op1_14_in06 = reg_0469;
    89: op1_14_in06 = reg_0251;
    90: op1_14_in06 = reg_0530;
    91: op1_14_in06 = imem06_in[3:0];
    92: op1_14_in06 = reg_0185;
    93: op1_14_in06 = reg_0141;
    94: op1_14_in06 = reg_0748;
    95: op1_14_in06 = reg_0038;
    default: op1_14_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv06 = 1;
    5: op1_14_inv06 = 1;
    6: op1_14_inv06 = 1;
    7: op1_14_inv06 = 1;
    14: op1_14_inv06 = 1;
    16: op1_14_inv06 = 1;
    17: op1_14_inv06 = 1;
    18: op1_14_inv06 = 1;
    19: op1_14_inv06 = 1;
    20: op1_14_inv06 = 1;
    21: op1_14_inv06 = 1;
    22: op1_14_inv06 = 1;
    25: op1_14_inv06 = 1;
    26: op1_14_inv06 = 1;
    27: op1_14_inv06 = 1;
    29: op1_14_inv06 = 1;
    30: op1_14_inv06 = 1;
    32: op1_14_inv06 = 1;
    33: op1_14_inv06 = 1;
    36: op1_14_inv06 = 1;
    37: op1_14_inv06 = 1;
    41: op1_14_inv06 = 1;
    42: op1_14_inv06 = 1;
    44: op1_14_inv06 = 1;
    45: op1_14_inv06 = 1;
    47: op1_14_inv06 = 1;
    48: op1_14_inv06 = 1;
    49: op1_14_inv06 = 1;
    51: op1_14_inv06 = 1;
    53: op1_14_inv06 = 1;
    55: op1_14_inv06 = 1;
    56: op1_14_inv06 = 1;
    60: op1_14_inv06 = 1;
    63: op1_14_inv06 = 1;
    64: op1_14_inv06 = 1;
    65: op1_14_inv06 = 1;
    66: op1_14_inv06 = 1;
    67: op1_14_inv06 = 1;
    68: op1_14_inv06 = 1;
    71: op1_14_inv06 = 1;
    73: op1_14_inv06 = 1;
    74: op1_14_inv06 = 1;
    76: op1_14_inv06 = 1;
    77: op1_14_inv06 = 1;
    78: op1_14_inv06 = 1;
    81: op1_14_inv06 = 1;
    85: op1_14_inv06 = 1;
    86: op1_14_inv06 = 1;
    88: op1_14_inv06 = 1;
    89: op1_14_inv06 = 1;
    92: op1_14_inv06 = 1;
    93: op1_14_inv06 = 1;
    default: op1_14_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in07 = reg_0475;
    5: op1_14_in07 = imem06_in[119:116];
    6: op1_14_in07 = imem02_in[115:112];
    18: op1_14_in07 = imem02_in[115:112];
    7: op1_14_in07 = reg_0384;
    8: op1_14_in07 = reg_0683;
    9: op1_14_in07 = reg_0604;
    10: op1_14_in07 = reg_0352;
    89: op1_14_in07 = reg_0352;
    11: op1_14_in07 = reg_0546;
    12: op1_14_in07 = reg_0102;
    13: op1_14_in07 = reg_0006;
    14: op1_14_in07 = reg_0484;
    15: op1_14_in07 = imem00_in[115:112];
    16: op1_14_in07 = reg_0650;
    17: op1_14_in07 = reg_0454;
    19: op1_14_in07 = reg_0689;
    40: op1_14_in07 = reg_0689;
    52: op1_14_in07 = reg_0689;
    20: op1_14_in07 = reg_0397;
    21: op1_14_in07 = reg_0486;
    22: op1_14_in07 = reg_0479;
    23: op1_14_in07 = imem07_in[39:36];
    24: op1_14_in07 = reg_0674;
    25: op1_14_in07 = reg_0529;
    26: op1_14_in07 = reg_0219;
    3: op1_14_in07 = reg_0160;
    27: op1_14_in07 = reg_0644;
    28: op1_14_in07 = reg_0608;
    29: op1_14_in07 = reg_0477;
    30: op1_14_in07 = reg_0803;
    31: op1_14_in07 = imem05_in[3:0];
    32: op1_14_in07 = reg_0285;
    2: op1_14_in07 = reg_0159;
    33: op1_14_in07 = reg_0530;
    34: op1_14_in07 = reg_0751;
    35: op1_14_in07 = reg_0575;
    36: op1_14_in07 = reg_0416;
    37: op1_14_in07 = imem05_in[7:4];
    41: op1_14_in07 = reg_0551;
    42: op1_14_in07 = reg_0766;
    43: op1_14_in07 = reg_0705;
    44: op1_14_in07 = reg_0105;
    45: op1_14_in07 = imem05_in[47:44];
    80: op1_14_in07 = imem05_in[47:44];
    46: op1_14_in07 = reg_0725;
    47: op1_14_in07 = imem02_in[95:92];
    81: op1_14_in07 = imem02_in[95:92];
    48: op1_14_in07 = reg_0589;
    49: op1_14_in07 = reg_0119;
    50: op1_14_in07 = reg_0690;
    51: op1_14_in07 = reg_0311;
    53: op1_14_in07 = reg_0697;
    54: op1_14_in07 = imem02_in[79:76];
    55: op1_14_in07 = reg_0318;
    56: op1_14_in07 = reg_0588;
    57: op1_14_in07 = reg_0666;
    58: op1_14_in07 = reg_0215;
    59: op1_14_in07 = reg_0116;
    60: op1_14_in07 = imem05_in[75:72];
    62: op1_14_in07 = reg_0091;
    63: op1_14_in07 = reg_0504;
    64: op1_14_in07 = imem02_in[43:40];
    65: op1_14_in07 = reg_0488;
    66: op1_14_in07 = reg_0485;
    67: op1_14_in07 = imem07_in[15:12];
    68: op1_14_in07 = reg_0492;
    69: op1_14_in07 = imem03_in[127:124];
    70: op1_14_in07 = reg_0035;
    71: op1_14_in07 = reg_0134;
    72: op1_14_in07 = reg_0403;
    73: op1_14_in07 = imem04_in[67:64];
    74: op1_14_in07 = imem05_in[79:76];
    75: op1_14_in07 = reg_0578;
    76: op1_14_in07 = imem00_in[91:88];
    77: op1_14_in07 = imem02_in[127:124];
    78: op1_14_in07 = imem02_in[67:64];
    79: op1_14_in07 = reg_0733;
    82: op1_14_in07 = reg_0696;
    84: op1_14_in07 = imem04_in[51:48];
    85: op1_14_in07 = reg_0648;
    86: op1_14_in07 = reg_0692;
    87: op1_14_in07 = reg_0549;
    88: op1_14_in07 = reg_0462;
    90: op1_14_in07 = reg_0656;
    91: op1_14_in07 = imem06_in[59:56];
    92: op1_14_in07 = reg_0427;
    93: op1_14_in07 = reg_0176;
    94: op1_14_in07 = reg_0638;
    95: op1_14_in07 = reg_0265;
    default: op1_14_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv07 = 1;
    5: op1_14_inv07 = 1;
    8: op1_14_inv07 = 1;
    9: op1_14_inv07 = 1;
    11: op1_14_inv07 = 1;
    14: op1_14_inv07 = 1;
    24: op1_14_inv07 = 1;
    26: op1_14_inv07 = 1;
    3: op1_14_inv07 = 1;
    29: op1_14_inv07 = 1;
    30: op1_14_inv07 = 1;
    31: op1_14_inv07 = 1;
    32: op1_14_inv07 = 1;
    2: op1_14_inv07 = 1;
    34: op1_14_inv07 = 1;
    36: op1_14_inv07 = 1;
    43: op1_14_inv07 = 1;
    45: op1_14_inv07 = 1;
    46: op1_14_inv07 = 1;
    48: op1_14_inv07 = 1;
    50: op1_14_inv07 = 1;
    54: op1_14_inv07 = 1;
    55: op1_14_inv07 = 1;
    56: op1_14_inv07 = 1;
    59: op1_14_inv07 = 1;
    71: op1_14_inv07 = 1;
    72: op1_14_inv07 = 1;
    73: op1_14_inv07 = 1;
    74: op1_14_inv07 = 1;
    76: op1_14_inv07 = 1;
    81: op1_14_inv07 = 1;
    82: op1_14_inv07 = 1;
    85: op1_14_inv07 = 1;
    86: op1_14_inv07 = 1;
    89: op1_14_inv07 = 1;
    90: op1_14_inv07 = 1;
    92: op1_14_inv07 = 1;
    93: op1_14_inv07 = 1;
    94: op1_14_inv07 = 1;
    95: op1_14_inv07 = 1;
    default: op1_14_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in08 = reg_0460;
    5: op1_14_in08 = imem06_in[123:120];
    6: op1_14_in08 = imem02_in[127:124];
    7: op1_14_in08 = reg_0362;
    8: op1_14_in08 = reg_0696;
    9: op1_14_in08 = reg_0616;
    10: op1_14_in08 = reg_0357;
    59: op1_14_in08 = reg_0357;
    11: op1_14_in08 = reg_0540;
    12: op1_14_in08 = imem02_in[7:4];
    13: op1_14_in08 = reg_0803;
    14: op1_14_in08 = reg_0493;
    15: op1_14_in08 = reg_0682;
    16: op1_14_in08 = reg_0645;
    17: op1_14_in08 = reg_0455;
    18: op1_14_in08 = reg_0642;
    19: op1_14_in08 = reg_0686;
    20: op1_14_in08 = reg_0393;
    21: op1_14_in08 = reg_0735;
    22: op1_14_in08 = reg_0210;
    23: op1_14_in08 = imem07_in[87:84];
    24: op1_14_in08 = reg_0678;
    25: op1_14_in08 = reg_0293;
    26: op1_14_in08 = reg_0111;
    3: op1_14_in08 = reg_0163;
    2: op1_14_in08 = reg_0163;
    27: op1_14_in08 = reg_0659;
    28: op1_14_in08 = reg_0615;
    29: op1_14_in08 = reg_0480;
    30: op1_14_in08 = reg_0804;
    31: op1_14_in08 = imem05_in[19:16];
    32: op1_14_in08 = reg_0086;
    33: op1_14_in08 = reg_0093;
    34: op1_14_in08 = reg_0384;
    85: op1_14_in08 = reg_0384;
    35: op1_14_in08 = reg_0517;
    36: op1_14_in08 = reg_0619;
    37: op1_14_in08 = imem05_in[87:84];
    40: op1_14_in08 = reg_0668;
    41: op1_14_in08 = reg_0510;
    42: op1_14_in08 = reg_0622;
    43: op1_14_in08 = reg_0053;
    44: op1_14_in08 = reg_0116;
    45: op1_14_in08 = imem05_in[63:60];
    46: op1_14_in08 = reg_0705;
    47: op1_14_in08 = reg_0647;
    48: op1_14_in08 = reg_0578;
    49: op1_14_in08 = reg_0117;
    50: op1_14_in08 = reg_0677;
    51: op1_14_in08 = reg_0614;
    52: op1_14_in08 = reg_0463;
    53: op1_14_in08 = reg_0694;
    54: op1_14_in08 = imem02_in[107:104];
    55: op1_14_in08 = reg_0329;
    56: op1_14_in08 = reg_0751;
    57: op1_14_in08 = reg_0651;
    58: op1_14_in08 = reg_0226;
    60: op1_14_in08 = imem05_in[99:96];
    62: op1_14_in08 = reg_0110;
    63: op1_14_in08 = reg_0506;
    64: op1_14_in08 = reg_0650;
    77: op1_14_in08 = reg_0650;
    65: op1_14_in08 = reg_0399;
    66: op1_14_in08 = reg_0586;
    67: op1_14_in08 = imem07_in[47:44];
    68: op1_14_in08 = reg_0689;
    69: op1_14_in08 = reg_0019;
    70: op1_14_in08 = imem06_in[43:40];
    71: op1_14_in08 = reg_0641;
    72: op1_14_in08 = reg_0549;
    73: op1_14_in08 = imem04_in[103:100];
    74: op1_14_in08 = imem05_in[95:92];
    75: op1_14_in08 = reg_0405;
    76: op1_14_in08 = imem00_in[99:96];
    78: op1_14_in08 = imem02_in[103:100];
    79: op1_14_in08 = reg_0747;
    80: op1_14_in08 = imem05_in[55:52];
    81: op1_14_in08 = imem02_in[115:112];
    82: op1_14_in08 = reg_0658;
    84: op1_14_in08 = imem04_in[79:76];
    86: op1_14_in08 = reg_0451;
    87: op1_14_in08 = reg_0496;
    88: op1_14_in08 = reg_0481;
    89: op1_14_in08 = reg_0358;
    90: op1_14_in08 = reg_0704;
    91: op1_14_in08 = imem06_in[83:80];
    93: op1_14_in08 = reg_0184;
    94: op1_14_in08 = reg_0655;
    95: op1_14_in08 = reg_0039;
    default: op1_14_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv08 = 1;
    5: op1_14_inv08 = 1;
    9: op1_14_inv08 = 1;
    11: op1_14_inv08 = 1;
    12: op1_14_inv08 = 1;
    13: op1_14_inv08 = 1;
    16: op1_14_inv08 = 1;
    18: op1_14_inv08 = 1;
    19: op1_14_inv08 = 1;
    21: op1_14_inv08 = 1;
    22: op1_14_inv08 = 1;
    23: op1_14_inv08 = 1;
    25: op1_14_inv08 = 1;
    27: op1_14_inv08 = 1;
    31: op1_14_inv08 = 1;
    32: op1_14_inv08 = 1;
    33: op1_14_inv08 = 1;
    35: op1_14_inv08 = 1;
    36: op1_14_inv08 = 1;
    40: op1_14_inv08 = 1;
    43: op1_14_inv08 = 1;
    45: op1_14_inv08 = 1;
    48: op1_14_inv08 = 1;
    49: op1_14_inv08 = 1;
    51: op1_14_inv08 = 1;
    53: op1_14_inv08 = 1;
    55: op1_14_inv08 = 1;
    60: op1_14_inv08 = 1;
    62: op1_14_inv08 = 1;
    64: op1_14_inv08 = 1;
    66: op1_14_inv08 = 1;
    71: op1_14_inv08 = 1;
    73: op1_14_inv08 = 1;
    75: op1_14_inv08 = 1;
    76: op1_14_inv08 = 1;
    79: op1_14_inv08 = 1;
    80: op1_14_inv08 = 1;
    81: op1_14_inv08 = 1;
    84: op1_14_inv08 = 1;
    88: op1_14_inv08 = 1;
    93: op1_14_inv08 = 1;
    94: op1_14_inv08 = 1;
    default: op1_14_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in09 = reg_0468;
    52: op1_14_in09 = reg_0468;
    5: op1_14_in09 = reg_0614;
    6: op1_14_in09 = reg_0658;
    7: op1_14_in09 = reg_0373;
    8: op1_14_in09 = reg_0685;
    9: op1_14_in09 = reg_0609;
    10: op1_14_in09 = reg_0338;
    11: op1_14_in09 = reg_0532;
    12: op1_14_in09 = imem02_in[31:28];
    13: op1_14_in09 = reg_0007;
    69: op1_14_in09 = reg_0007;
    14: op1_14_in09 = reg_0793;
    15: op1_14_in09 = reg_0690;
    16: op1_14_in09 = reg_0655;
    17: op1_14_in09 = reg_0469;
    18: op1_14_in09 = reg_0661;
    19: op1_14_in09 = reg_0677;
    20: op1_14_in09 = reg_0019;
    21: op1_14_in09 = reg_0260;
    22: op1_14_in09 = reg_0202;
    23: op1_14_in09 = imem07_in[119:116];
    24: op1_14_in09 = reg_0692;
    25: op1_14_in09 = reg_0290;
    26: op1_14_in09 = reg_0119;
    44: op1_14_in09 = reg_0119;
    3: op1_14_in09 = reg_0183;
    27: op1_14_in09 = reg_0360;
    28: op1_14_in09 = imem06_in[7:4];
    29: op1_14_in09 = reg_0471;
    30: op1_14_in09 = reg_0004;
    31: op1_14_in09 = imem05_in[39:36];
    32: op1_14_in09 = reg_0145;
    33: op1_14_in09 = imem03_in[7:4];
    34: op1_14_in09 = reg_0391;
    65: op1_14_in09 = reg_0391;
    35: op1_14_in09 = reg_0374;
    36: op1_14_in09 = reg_0625;
    37: op1_14_in09 = imem05_in[115:112];
    40: op1_14_in09 = reg_0680;
    41: op1_14_in09 = imem04_in[19:16];
    42: op1_14_in09 = reg_0774;
    43: op1_14_in09 = reg_0635;
    45: op1_14_in09 = imem05_in[71:68];
    46: op1_14_in09 = reg_0706;
    47: op1_14_in09 = reg_0346;
    48: op1_14_in09 = reg_0581;
    49: op1_14_in09 = reg_0126;
    50: op1_14_in09 = reg_0673;
    51: op1_14_in09 = reg_0607;
    53: op1_14_in09 = reg_0698;
    54: op1_14_in09 = reg_0642;
    55: op1_14_in09 = reg_0588;
    59: op1_14_in09 = reg_0588;
    56: op1_14_in09 = reg_0568;
    57: op1_14_in09 = reg_0647;
    58: op1_14_in09 = reg_0279;
    60: op1_14_in09 = reg_0091;
    62: op1_14_in09 = reg_0075;
    63: op1_14_in09 = reg_0104;
    64: op1_14_in09 = reg_0584;
    66: op1_14_in09 = reg_0565;
    67: op1_14_in09 = imem07_in[67:64];
    68: op1_14_in09 = reg_0744;
    70: op1_14_in09 = imem06_in[87:84];
    71: op1_14_in09 = reg_0355;
    72: op1_14_in09 = reg_0747;
    73: op1_14_in09 = reg_0315;
    74: op1_14_in09 = imem05_in[103:100];
    75: op1_14_in09 = reg_0816;
    76: op1_14_in09 = imem00_in[119:116];
    77: op1_14_in09 = reg_0254;
    78: op1_14_in09 = reg_0639;
    79: op1_14_in09 = reg_0000;
    80: op1_14_in09 = imem05_in[59:56];
    81: op1_14_in09 = imem02_in[127:124];
    82: op1_14_in09 = reg_0758;
    84: op1_14_in09 = imem04_in[91:88];
    85: op1_14_in09 = reg_0575;
    86: op1_14_in09 = reg_0477;
    87: op1_14_in09 = reg_0396;
    88: op1_14_in09 = reg_0472;
    89: op1_14_in09 = reg_0363;
    90: op1_14_in09 = reg_0324;
    91: op1_14_in09 = reg_0624;
    94: op1_14_in09 = reg_0335;
    95: op1_14_in09 = reg_0630;
    default: op1_14_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv09 = 1;
    5: op1_14_inv09 = 1;
    6: op1_14_inv09 = 1;
    7: op1_14_inv09 = 1;
    9: op1_14_inv09 = 1;
    10: op1_14_inv09 = 1;
    16: op1_14_inv09 = 1;
    18: op1_14_inv09 = 1;
    19: op1_14_inv09 = 1;
    21: op1_14_inv09 = 1;
    22: op1_14_inv09 = 1;
    23: op1_14_inv09 = 1;
    24: op1_14_inv09 = 1;
    26: op1_14_inv09 = 1;
    27: op1_14_inv09 = 1;
    29: op1_14_inv09 = 1;
    30: op1_14_inv09 = 1;
    32: op1_14_inv09 = 1;
    34: op1_14_inv09 = 1;
    36: op1_14_inv09 = 1;
    40: op1_14_inv09 = 1;
    41: op1_14_inv09 = 1;
    42: op1_14_inv09 = 1;
    44: op1_14_inv09 = 1;
    47: op1_14_inv09 = 1;
    50: op1_14_inv09 = 1;
    52: op1_14_inv09 = 1;
    63: op1_14_inv09 = 1;
    64: op1_14_inv09 = 1;
    65: op1_14_inv09 = 1;
    66: op1_14_inv09 = 1;
    67: op1_14_inv09 = 1;
    68: op1_14_inv09 = 1;
    70: op1_14_inv09 = 1;
    75: op1_14_inv09 = 1;
    76: op1_14_inv09 = 1;
    78: op1_14_inv09 = 1;
    79: op1_14_inv09 = 1;
    82: op1_14_inv09 = 1;
    84: op1_14_inv09 = 1;
    85: op1_14_inv09 = 1;
    89: op1_14_inv09 = 1;
    90: op1_14_inv09 = 1;
    91: op1_14_inv09 = 1;
    94: op1_14_inv09 = 1;
    default: op1_14_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in10 = reg_0192;
    5: op1_14_in10 = reg_0625;
    6: op1_14_in10 = reg_0664;
    7: op1_14_in10 = reg_0322;
    8: op1_14_in10 = reg_0672;
    9: op1_14_in10 = reg_0611;
    10: op1_14_in10 = reg_0350;
    11: op1_14_in10 = reg_0558;
    12: op1_14_in10 = imem02_in[51:48];
    13: op1_14_in10 = reg_0800;
    14: op1_14_in10 = reg_0783;
    15: op1_14_in10 = reg_0671;
    16: op1_14_in10 = reg_0661;
    17: op1_14_in10 = reg_0472;
    18: op1_14_in10 = reg_0647;
    19: op1_14_in10 = reg_0678;
    20: op1_14_in10 = reg_0012;
    21: op1_14_in10 = reg_0269;
    22: op1_14_in10 = reg_0197;
    23: op1_14_in10 = imem07_in[127:124];
    24: op1_14_in10 = reg_0465;
    25: op1_14_in10 = reg_0268;
    26: op1_14_in10 = reg_0115;
    3: op1_14_in10 = reg_0185;
    27: op1_14_in10 = reg_0081;
    28: op1_14_in10 = imem06_in[19:16];
    29: op1_14_in10 = reg_0479;
    30: op1_14_in10 = imem04_in[11:8];
    31: op1_14_in10 = imem05_in[63:60];
    32: op1_14_in10 = imem06_in[11:8];
    33: op1_14_in10 = imem03_in[59:56];
    34: op1_14_in10 = reg_0575;
    35: op1_14_in10 = reg_0389;
    36: op1_14_in10 = reg_0605;
    37: op1_14_in10 = reg_0490;
    40: op1_14_in10 = reg_0455;
    41: op1_14_in10 = imem04_in[43:40];
    42: op1_14_in10 = reg_0318;
    43: op1_14_in10 = reg_0061;
    44: op1_14_in10 = reg_0100;
    45: op1_14_in10 = imem05_in[79:76];
    80: op1_14_in10 = imem05_in[79:76];
    46: op1_14_in10 = reg_0295;
    47: op1_14_in10 = reg_0638;
    48: op1_14_in10 = reg_0595;
    49: op1_14_in10 = reg_0110;
    50: op1_14_in10 = reg_0699;
    53: op1_14_in10 = reg_0699;
    51: op1_14_in10 = reg_0372;
    52: op1_14_in10 = reg_0209;
    54: op1_14_in10 = reg_0657;
    75: op1_14_in10 = reg_0657;
    55: op1_14_in10 = reg_0395;
    56: op1_14_in10 = reg_0386;
    57: op1_14_in10 = reg_0301;
    58: op1_14_in10 = reg_0224;
    59: op1_14_in10 = reg_0509;
    60: op1_14_in10 = reg_0103;
    62: op1_14_in10 = reg_0112;
    63: op1_14_in10 = reg_0677;
    64: op1_14_in10 = reg_0483;
    65: op1_14_in10 = reg_0747;
    66: op1_14_in10 = reg_0414;
    67: op1_14_in10 = imem07_in[71:68];
    68: op1_14_in10 = reg_0470;
    69: op1_14_in10 = reg_0799;
    70: op1_14_in10 = imem06_in[111:108];
    71: op1_14_in10 = reg_0135;
    72: op1_14_in10 = reg_0557;
    73: op1_14_in10 = reg_0060;
    74: op1_14_in10 = imem05_in[107:104];
    76: op1_14_in10 = imem00_in[127:124];
    77: op1_14_in10 = reg_0621;
    78: op1_14_in10 = reg_0753;
    79: op1_14_in10 = reg_0002;
    81: op1_14_in10 = reg_0534;
    82: op1_14_in10 = reg_0463;
    84: op1_14_in10 = imem04_in[103:100];
    85: op1_14_in10 = reg_0568;
    86: op1_14_in10 = reg_0469;
    87: op1_14_in10 = reg_0570;
    88: op1_14_in10 = reg_0474;
    89: op1_14_in10 = reg_0132;
    90: op1_14_in10 = reg_0527;
    91: op1_14_in10 = reg_0405;
    94: op1_14_in10 = reg_0620;
    95: op1_14_in10 = reg_0659;
    default: op1_14_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv10 = 1;
    5: op1_14_inv10 = 1;
    6: op1_14_inv10 = 1;
    8: op1_14_inv10 = 1;
    11: op1_14_inv10 = 1;
    13: op1_14_inv10 = 1;
    14: op1_14_inv10 = 1;
    18: op1_14_inv10 = 1;
    19: op1_14_inv10 = 1;
    20: op1_14_inv10 = 1;
    23: op1_14_inv10 = 1;
    24: op1_14_inv10 = 1;
    25: op1_14_inv10 = 1;
    3: op1_14_inv10 = 1;
    27: op1_14_inv10 = 1;
    30: op1_14_inv10 = 1;
    32: op1_14_inv10 = 1;
    33: op1_14_inv10 = 1;
    34: op1_14_inv10 = 1;
    40: op1_14_inv10 = 1;
    41: op1_14_inv10 = 1;
    42: op1_14_inv10 = 1;
    43: op1_14_inv10 = 1;
    44: op1_14_inv10 = 1;
    46: op1_14_inv10 = 1;
    47: op1_14_inv10 = 1;
    48: op1_14_inv10 = 1;
    50: op1_14_inv10 = 1;
    52: op1_14_inv10 = 1;
    54: op1_14_inv10 = 1;
    56: op1_14_inv10 = 1;
    58: op1_14_inv10 = 1;
    59: op1_14_inv10 = 1;
    60: op1_14_inv10 = 1;
    62: op1_14_inv10 = 1;
    65: op1_14_inv10 = 1;
    68: op1_14_inv10 = 1;
    71: op1_14_inv10 = 1;
    72: op1_14_inv10 = 1;
    75: op1_14_inv10 = 1;
    76: op1_14_inv10 = 1;
    77: op1_14_inv10 = 1;
    78: op1_14_inv10 = 1;
    79: op1_14_inv10 = 1;
    81: op1_14_inv10 = 1;
    85: op1_14_inv10 = 1;
    86: op1_14_inv10 = 1;
    87: op1_14_inv10 = 1;
    90: op1_14_inv10 = 1;
    default: op1_14_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in11 = imem01_in[43:40];
    5: op1_14_in11 = reg_0605;
    6: op1_14_in11 = reg_0661;
    7: op1_14_in11 = reg_0361;
    8: op1_14_in11 = reg_0676;
    9: op1_14_in11 = reg_0618;
    10: op1_14_in11 = reg_0042;
    11: op1_14_in11 = reg_0533;
    12: op1_14_in11 = imem02_in[79:76];
    13: op1_14_in11 = reg_0805;
    14: op1_14_in11 = reg_0786;
    15: op1_14_in11 = reg_0680;
    16: op1_14_in11 = reg_0639;
    77: op1_14_in11 = reg_0639;
    17: op1_14_in11 = reg_0471;
    18: op1_14_in11 = reg_0649;
    72: op1_14_in11 = reg_0649;
    19: op1_14_in11 = reg_0688;
    20: op1_14_in11 = reg_0803;
    21: op1_14_in11 = reg_0277;
    22: op1_14_in11 = imem01_in[63:60];
    23: op1_14_in11 = reg_0716;
    24: op1_14_in11 = reg_0454;
    25: op1_14_in11 = reg_0292;
    26: op1_14_in11 = reg_0121;
    3: op1_14_in11 = reg_0157;
    27: op1_14_in11 = reg_0080;
    28: op1_14_in11 = imem06_in[43:40];
    29: op1_14_in11 = reg_0459;
    30: op1_14_in11 = imem04_in[19:16];
    31: op1_14_in11 = imem05_in[75:72];
    32: op1_14_in11 = imem06_in[47:44];
    33: op1_14_in11 = imem03_in[83:80];
    34: op1_14_in11 = reg_0561;
    35: op1_14_in11 = reg_0001;
    87: op1_14_in11 = reg_0001;
    36: op1_14_in11 = reg_0633;
    37: op1_14_in11 = reg_0495;
    40: op1_14_in11 = reg_0461;
    41: op1_14_in11 = imem04_in[55:52];
    42: op1_14_in11 = reg_0407;
    43: op1_14_in11 = reg_0440;
    44: op1_14_in11 = reg_0101;
    45: op1_14_in11 = imem05_in[95:92];
    46: op1_14_in11 = reg_0636;
    47: op1_14_in11 = reg_0662;
    48: op1_14_in11 = reg_0751;
    49: op1_14_in11 = imem02_in[7:4];
    50: op1_14_in11 = reg_0464;
    51: op1_14_in11 = reg_0819;
    52: op1_14_in11 = reg_0204;
    53: op1_14_in11 = reg_0451;
    54: op1_14_in11 = reg_0647;
    55: op1_14_in11 = reg_0564;
    56: op1_14_in11 = reg_0570;
    57: op1_14_in11 = reg_0485;
    58: op1_14_in11 = reg_0066;
    59: op1_14_in11 = reg_0383;
    60: op1_14_in11 = reg_0070;
    62: op1_14_in11 = reg_0231;
    63: op1_14_in11 = reg_0669;
    64: op1_14_in11 = reg_0417;
    65: op1_14_in11 = reg_0006;
    66: op1_14_in11 = reg_0527;
    67: op1_14_in11 = imem07_in[87:84];
    68: op1_14_in11 = reg_0474;
    69: op1_14_in11 = reg_0004;
    70: op1_14_in11 = imem07_in[39:36];
    71: op1_14_in11 = imem02_in[27:24];
    73: op1_14_in11 = reg_0558;
    74: op1_14_in11 = imem05_in[115:112];
    75: op1_14_in11 = reg_0767;
    76: op1_14_in11 = reg_0744;
    78: op1_14_in11 = reg_0655;
    79: op1_14_in11 = reg_0802;
    80: op1_14_in11 = imem05_in[91:88];
    81: op1_14_in11 = reg_0392;
    82: op1_14_in11 = reg_0450;
    84: op1_14_in11 = imem04_in[107:104];
    85: op1_14_in11 = reg_0398;
    86: op1_14_in11 = reg_0473;
    88: op1_14_in11 = reg_0479;
    89: op1_14_in11 = reg_0756;
    90: op1_14_in11 = reg_0590;
    91: op1_14_in11 = reg_0246;
    94: op1_14_in11 = reg_0351;
    95: op1_14_in11 = reg_0276;
    default: op1_14_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv11 = 1;
    7: op1_14_inv11 = 1;
    10: op1_14_inv11 = 1;
    11: op1_14_inv11 = 1;
    12: op1_14_inv11 = 1;
    13: op1_14_inv11 = 1;
    16: op1_14_inv11 = 1;
    17: op1_14_inv11 = 1;
    18: op1_14_inv11 = 1;
    24: op1_14_inv11 = 1;
    25: op1_14_inv11 = 1;
    26: op1_14_inv11 = 1;
    29: op1_14_inv11 = 1;
    30: op1_14_inv11 = 1;
    31: op1_14_inv11 = 1;
    34: op1_14_inv11 = 1;
    36: op1_14_inv11 = 1;
    40: op1_14_inv11 = 1;
    41: op1_14_inv11 = 1;
    42: op1_14_inv11 = 1;
    43: op1_14_inv11 = 1;
    44: op1_14_inv11 = 1;
    45: op1_14_inv11 = 1;
    47: op1_14_inv11 = 1;
    49: op1_14_inv11 = 1;
    50: op1_14_inv11 = 1;
    51: op1_14_inv11 = 1;
    54: op1_14_inv11 = 1;
    56: op1_14_inv11 = 1;
    59: op1_14_inv11 = 1;
    60: op1_14_inv11 = 1;
    63: op1_14_inv11 = 1;
    65: op1_14_inv11 = 1;
    66: op1_14_inv11 = 1;
    70: op1_14_inv11 = 1;
    71: op1_14_inv11 = 1;
    72: op1_14_inv11 = 1;
    76: op1_14_inv11 = 1;
    78: op1_14_inv11 = 1;
    79: op1_14_inv11 = 1;
    80: op1_14_inv11 = 1;
    81: op1_14_inv11 = 1;
    84: op1_14_inv11 = 1;
    85: op1_14_inv11 = 1;
    86: op1_14_inv11 = 1;
    87: op1_14_inv11 = 1;
    89: op1_14_inv11 = 1;
    90: op1_14_inv11 = 1;
    default: op1_14_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in12 = imem01_in[59:56];
    5: op1_14_in12 = reg_0626;
    6: op1_14_in12 = reg_0656;
    7: op1_14_in12 = reg_0002;
    8: op1_14_in12 = reg_0698;
    9: op1_14_in12 = reg_0356;
    10: op1_14_in12 = reg_0055;
    11: op1_14_in12 = reg_0556;
    12: op1_14_in12 = reg_0646;
    13: op1_14_in12 = reg_0802;
    14: op1_14_in12 = reg_0489;
    15: op1_14_in12 = reg_0699;
    16: op1_14_in12 = reg_0651;
    95: op1_14_in12 = reg_0651;
    17: op1_14_in12 = reg_0452;
    18: op1_14_in12 = reg_0352;
    19: op1_14_in12 = reg_0669;
    20: op1_14_in12 = reg_0014;
    21: op1_14_in12 = reg_0086;
    22: op1_14_in12 = imem01_in[71:68];
    23: op1_14_in12 = reg_0719;
    24: op1_14_in12 = reg_0451;
    25: op1_14_in12 = reg_0257;
    26: op1_14_in12 = reg_0126;
    3: op1_14_in12 = reg_0173;
    27: op1_14_in12 = reg_0530;
    28: op1_14_in12 = imem06_in[47:44];
    29: op1_14_in12 = reg_0191;
    30: op1_14_in12 = imem04_in[23:20];
    31: op1_14_in12 = imem05_in[103:100];
    32: op1_14_in12 = imem06_in[55:52];
    33: op1_14_in12 = imem03_in[87:84];
    34: op1_14_in12 = reg_0572;
    35: op1_14_in12 = reg_0801;
    36: op1_14_in12 = reg_0380;
    37: op1_14_in12 = reg_0091;
    40: op1_14_in12 = reg_0476;
    53: op1_14_in12 = reg_0476;
    41: op1_14_in12 = imem04_in[59:56];
    79: op1_14_in12 = imem04_in[59:56];
    42: op1_14_in12 = reg_0821;
    43: op1_14_in12 = reg_0442;
    44: op1_14_in12 = reg_0109;
    45: op1_14_in12 = imem05_in[127:124];
    46: op1_14_in12 = reg_0447;
    47: op1_14_in12 = reg_0355;
    48: op1_14_in12 = reg_0590;
    49: op1_14_in12 = imem02_in[27:24];
    50: op1_14_in12 = reg_0466;
    51: op1_14_in12 = reg_0375;
    52: op1_14_in12 = reg_0188;
    54: op1_14_in12 = reg_0427;
    78: op1_14_in12 = reg_0427;
    55: op1_14_in12 = reg_0569;
    56: op1_14_in12 = reg_0006;
    72: op1_14_in12 = reg_0006;
    57: op1_14_in12 = reg_0587;
    58: op1_14_in12 = reg_0135;
    59: op1_14_in12 = reg_0393;
    60: op1_14_in12 = reg_0226;
    62: op1_14_in12 = reg_0224;
    63: op1_14_in12 = imem02_in[23:20];
    64: op1_14_in12 = reg_0344;
    65: op1_14_in12 = reg_0007;
    66: op1_14_in12 = reg_0566;
    67: op1_14_in12 = imem07_in[107:104];
    68: op1_14_in12 = reg_0456;
    69: op1_14_in12 = imem04_in[7:4];
    70: op1_14_in12 = imem07_in[55:52];
    71: op1_14_in12 = imem02_in[47:44];
    73: op1_14_in12 = reg_0308;
    74: op1_14_in12 = reg_0667;
    75: op1_14_in12 = reg_0752;
    76: op1_14_in12 = reg_0247;
    77: op1_14_in12 = reg_0304;
    80: op1_14_in12 = imem05_in[99:96];
    81: op1_14_in12 = reg_0487;
    82: op1_14_in12 = reg_0481;
    84: op1_14_in12 = imem04_in[115:112];
    85: op1_14_in12 = reg_0637;
    86: op1_14_in12 = reg_0459;
    88: op1_14_in12 = reg_0459;
    87: op1_14_in12 = reg_0808;
    89: op1_14_in12 = reg_0098;
    90: op1_14_in12 = reg_0043;
    91: op1_14_in12 = reg_0169;
    94: op1_14_in12 = reg_0664;
    default: op1_14_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv12 = 1;
    6: op1_14_inv12 = 1;
    8: op1_14_inv12 = 1;
    9: op1_14_inv12 = 1;
    10: op1_14_inv12 = 1;
    11: op1_14_inv12 = 1;
    12: op1_14_inv12 = 1;
    15: op1_14_inv12 = 1;
    16: op1_14_inv12 = 1;
    17: op1_14_inv12 = 1;
    19: op1_14_inv12 = 1;
    21: op1_14_inv12 = 1;
    26: op1_14_inv12 = 1;
    3: op1_14_inv12 = 1;
    27: op1_14_inv12 = 1;
    28: op1_14_inv12 = 1;
    32: op1_14_inv12 = 1;
    33: op1_14_inv12 = 1;
    35: op1_14_inv12 = 1;
    37: op1_14_inv12 = 1;
    40: op1_14_inv12 = 1;
    43: op1_14_inv12 = 1;
    44: op1_14_inv12 = 1;
    46: op1_14_inv12 = 1;
    47: op1_14_inv12 = 1;
    51: op1_14_inv12 = 1;
    54: op1_14_inv12 = 1;
    55: op1_14_inv12 = 1;
    57: op1_14_inv12 = 1;
    58: op1_14_inv12 = 1;
    64: op1_14_inv12 = 1;
    65: op1_14_inv12 = 1;
    66: op1_14_inv12 = 1;
    67: op1_14_inv12 = 1;
    69: op1_14_inv12 = 1;
    78: op1_14_inv12 = 1;
    85: op1_14_inv12 = 1;
    87: op1_14_inv12 = 1;
    90: op1_14_inv12 = 1;
    94: op1_14_inv12 = 1;
    default: op1_14_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in13 = imem01_in[67:64];
    5: op1_14_in13 = reg_0618;
    6: op1_14_in13 = reg_0651;
    7: op1_14_in13 = reg_0808;
    8: op1_14_in13 = reg_0679;
    9: op1_14_in13 = reg_0381;
    10: op1_14_in13 = imem03_in[23:20];
    11: op1_14_in13 = reg_0299;
    12: op1_14_in13 = reg_0363;
    13: op1_14_in13 = reg_0799;
    14: op1_14_in13 = reg_0273;
    15: op1_14_in13 = reg_0451;
    16: op1_14_in13 = reg_0640;
    17: op1_14_in13 = reg_0196;
    18: op1_14_in13 = reg_0357;
    19: op1_14_in13 = reg_0464;
    20: op1_14_in13 = reg_0016;
    21: op1_14_in13 = reg_0132;
    22: op1_14_in13 = reg_0822;
    23: op1_14_in13 = reg_0721;
    24: op1_14_in13 = reg_0475;
    25: op1_14_in13 = reg_0065;
    26: op1_14_in13 = reg_0110;
    27: op1_14_in13 = reg_0757;
    28: op1_14_in13 = imem06_in[55:52];
    29: op1_14_in13 = reg_0211;
    30: op1_14_in13 = imem04_in[103:100];
    31: op1_14_in13 = imem05_in[119:116];
    32: op1_14_in13 = imem06_in[95:92];
    33: op1_14_in13 = imem03_in[91:88];
    34: op1_14_in13 = reg_0747;
    59: op1_14_in13 = reg_0747;
    35: op1_14_in13 = imem04_in[3:0];
    36: op1_14_in13 = reg_0612;
    37: op1_14_in13 = reg_0275;
    40: op1_14_in13 = reg_0479;
    41: op1_14_in13 = imem04_in[63:60];
    42: op1_14_in13 = reg_0607;
    43: op1_14_in13 = reg_0267;
    44: op1_14_in13 = reg_0653;
    45: op1_14_in13 = reg_0796;
    46: op1_14_in13 = reg_0635;
    47: op1_14_in13 = reg_0665;
    48: op1_14_in13 = reg_0384;
    49: op1_14_in13 = imem02_in[51:48];
    50: op1_14_in13 = reg_0470;
    51: op1_14_in13 = imem07_in[55:52];
    52: op1_14_in13 = reg_0255;
    53: op1_14_in13 = reg_0466;
    54: op1_14_in13 = reg_0359;
    55: op1_14_in13 = reg_0376;
    56: op1_14_in13 = reg_0013;
    57: op1_14_in13 = reg_0358;
    58: op1_14_in13 = reg_0154;
    60: op1_14_in13 = reg_0258;
    62: op1_14_in13 = reg_0236;
    63: op1_14_in13 = imem02_in[111:108];
    64: op1_14_in13 = reg_0343;
    65: op1_14_in13 = reg_0804;
    66: op1_14_in13 = reg_0081;
    67: op1_14_in13 = reg_0719;
    68: op1_14_in13 = reg_0189;
    69: op1_14_in13 = imem04_in[11:8];
    70: op1_14_in13 = imem07_in[79:76];
    71: op1_14_in13 = imem02_in[63:60];
    72: op1_14_in13 = reg_0002;
    73: op1_14_in13 = reg_0280;
    74: op1_14_in13 = reg_0070;
    75: op1_14_in13 = imem07_in[3:0];
    76: op1_14_in13 = reg_0465;
    77: op1_14_in13 = reg_0702;
    78: op1_14_in13 = reg_0360;
    79: op1_14_in13 = reg_0059;
    80: op1_14_in13 = imem05_in[127:124];
    81: op1_14_in13 = reg_0656;
    82: op1_14_in13 = reg_0456;
    84: op1_14_in13 = imem04_in[119:116];
    85: op1_14_in13 = reg_0019;
    86: op1_14_in13 = reg_0204;
    87: op1_14_in13 = reg_0807;
    88: op1_14_in13 = reg_0188;
    89: op1_14_in13 = reg_0317;
    90: op1_14_in13 = reg_0314;
    91: op1_14_in13 = reg_0663;
    94: op1_14_in13 = reg_0633;
    95: op1_14_in13 = reg_0351;
    default: op1_14_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv13 = 1;
    5: op1_14_inv13 = 1;
    6: op1_14_inv13 = 1;
    7: op1_14_inv13 = 1;
    8: op1_14_inv13 = 1;
    10: op1_14_inv13 = 1;
    13: op1_14_inv13 = 1;
    16: op1_14_inv13 = 1;
    25: op1_14_inv13 = 1;
    26: op1_14_inv13 = 1;
    28: op1_14_inv13 = 1;
    29: op1_14_inv13 = 1;
    30: op1_14_inv13 = 1;
    32: op1_14_inv13 = 1;
    33: op1_14_inv13 = 1;
    36: op1_14_inv13 = 1;
    41: op1_14_inv13 = 1;
    42: op1_14_inv13 = 1;
    43: op1_14_inv13 = 1;
    44: op1_14_inv13 = 1;
    47: op1_14_inv13 = 1;
    48: op1_14_inv13 = 1;
    50: op1_14_inv13 = 1;
    58: op1_14_inv13 = 1;
    59: op1_14_inv13 = 1;
    62: op1_14_inv13 = 1;
    63: op1_14_inv13 = 1;
    66: op1_14_inv13 = 1;
    68: op1_14_inv13 = 1;
    71: op1_14_inv13 = 1;
    72: op1_14_inv13 = 1;
    78: op1_14_inv13 = 1;
    79: op1_14_inv13 = 1;
    81: op1_14_inv13 = 1;
    88: op1_14_inv13 = 1;
    95: op1_14_inv13 = 1;
    default: op1_14_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in14 = imem01_in[75:72];
    5: op1_14_in14 = reg_0356;
    6: op1_14_in14 = reg_0636;
    7: op1_14_in14 = reg_0804;
    8: op1_14_in14 = reg_0677;
    9: op1_14_in14 = reg_0408;
    10: op1_14_in14 = imem03_in[59:56];
    11: op1_14_in14 = reg_0282;
    37: op1_14_in14 = reg_0282;
    12: op1_14_in14 = reg_0328;
    13: op1_14_in14 = reg_0810;
    20: op1_14_in14 = reg_0810;
    14: op1_14_in14 = reg_0226;
    15: op1_14_in14 = reg_0464;
    76: op1_14_in14 = reg_0464;
    16: op1_14_in14 = reg_0663;
    17: op1_14_in14 = reg_0202;
    18: op1_14_in14 = reg_0320;
    19: op1_14_in14 = reg_0461;
    21: op1_14_in14 = reg_0148;
    22: op1_14_in14 = reg_0517;
    23: op1_14_in14 = reg_0717;
    24: op1_14_in14 = reg_0472;
    25: op1_14_in14 = reg_0070;
    26: op1_14_in14 = imem02_in[27:24];
    27: op1_14_in14 = reg_0538;
    28: op1_14_in14 = imem06_in[75:72];
    29: op1_14_in14 = reg_0201;
    30: op1_14_in14 = reg_0262;
    84: op1_14_in14 = reg_0262;
    31: op1_14_in14 = reg_0792;
    32: op1_14_in14 = imem06_in[123:120];
    33: op1_14_in14 = imem03_in[95:92];
    34: op1_14_in14 = reg_0374;
    77: op1_14_in14 = reg_0374;
    35: op1_14_in14 = imem04_in[95:92];
    36: op1_14_in14 = reg_0402;
    40: op1_14_in14 = reg_0452;
    50: op1_14_in14 = reg_0452;
    41: op1_14_in14 = imem04_in[71:68];
    42: op1_14_in14 = reg_0778;
    43: op1_14_in14 = reg_0159;
    44: op1_14_in14 = reg_0646;
    45: op1_14_in14 = reg_0491;
    46: op1_14_in14 = reg_0440;
    47: op1_14_in14 = reg_0427;
    48: op1_14_in14 = reg_0376;
    49: op1_14_in14 = imem02_in[63:60];
    51: op1_14_in14 = imem07_in[67:64];
    52: op1_14_in14 = reg_0260;
    53: op1_14_in14 = reg_0481;
    54: op1_14_in14 = reg_0565;
    55: op1_14_in14 = reg_0499;
    56: op1_14_in14 = reg_0806;
    57: op1_14_in14 = reg_0581;
    58: op1_14_in14 = reg_0141;
    59: op1_14_in14 = reg_0013;
    60: op1_14_in14 = reg_0066;
    62: op1_14_in14 = imem02_in[3:0];
    63: op1_14_in14 = reg_0403;
    64: op1_14_in14 = reg_0323;
    78: op1_14_in14 = reg_0323;
    65: op1_14_in14 = reg_0010;
    66: op1_14_in14 = reg_0080;
    67: op1_14_in14 = reg_0710;
    68: op1_14_in14 = reg_0207;
    69: op1_14_in14 = imem04_in[35:32];
    70: op1_14_in14 = imem07_in[103:100];
    71: op1_14_in14 = imem02_in[75:72];
    72: op1_14_in14 = reg_0803;
    73: op1_14_in14 = reg_0626;
    74: op1_14_in14 = reg_0355;
    75: op1_14_in14 = imem07_in[11:8];
    79: op1_14_in14 = reg_0560;
    80: op1_14_in14 = reg_0337;
    81: op1_14_in14 = reg_0639;
    82: op1_14_in14 = reg_0200;
    85: op1_14_in14 = reg_0001;
    86: op1_14_in14 = reg_0194;
    87: op1_14_in14 = reg_0805;
    88: op1_14_in14 = reg_0211;
    89: op1_14_in14 = reg_0187;
    90: op1_14_in14 = reg_0132;
    91: op1_14_in14 = reg_0609;
    94: op1_14_in14 = reg_0680;
    95: op1_14_in14 = reg_0819;
    default: op1_14_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv14 = 1;
    5: op1_14_inv14 = 1;
    6: op1_14_inv14 = 1;
    8: op1_14_inv14 = 1;
    10: op1_14_inv14 = 1;
    12: op1_14_inv14 = 1;
    13: op1_14_inv14 = 1;
    14: op1_14_inv14 = 1;
    15: op1_14_inv14 = 1;
    16: op1_14_inv14 = 1;
    17: op1_14_inv14 = 1;
    22: op1_14_inv14 = 1;
    24: op1_14_inv14 = 1;
    25: op1_14_inv14 = 1;
    26: op1_14_inv14 = 1;
    30: op1_14_inv14 = 1;
    31: op1_14_inv14 = 1;
    32: op1_14_inv14 = 1;
    33: op1_14_inv14 = 1;
    35: op1_14_inv14 = 1;
    37: op1_14_inv14 = 1;
    40: op1_14_inv14 = 1;
    42: op1_14_inv14 = 1;
    44: op1_14_inv14 = 1;
    45: op1_14_inv14 = 1;
    48: op1_14_inv14 = 1;
    52: op1_14_inv14 = 1;
    53: op1_14_inv14 = 1;
    54: op1_14_inv14 = 1;
    55: op1_14_inv14 = 1;
    57: op1_14_inv14 = 1;
    63: op1_14_inv14 = 1;
    64: op1_14_inv14 = 1;
    65: op1_14_inv14 = 1;
    68: op1_14_inv14 = 1;
    69: op1_14_inv14 = 1;
    70: op1_14_inv14 = 1;
    73: op1_14_inv14 = 1;
    74: op1_14_inv14 = 1;
    77: op1_14_inv14 = 1;
    79: op1_14_inv14 = 1;
    80: op1_14_inv14 = 1;
    81: op1_14_inv14 = 1;
    85: op1_14_inv14 = 1;
    87: op1_14_inv14 = 1;
    89: op1_14_inv14 = 1;
    91: op1_14_inv14 = 1;
    94: op1_14_inv14 = 1;
    95: op1_14_inv14 = 1;
    default: op1_14_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in15 = imem01_in[83:80];
    5: op1_14_in15 = reg_0372;
    6: op1_14_in15 = reg_0333;
    7: op1_14_in15 = reg_0800;
    8: op1_14_in15 = reg_0691;
    9: op1_14_in15 = reg_0392;
    10: op1_14_in15 = imem03_in[87:84];
    11: op1_14_in15 = reg_0296;
    12: op1_14_in15 = reg_0086;
    13: op1_14_in15 = imem04_in[47:44];
    14: op1_14_in15 = reg_0734;
    15: op1_14_in15 = reg_0474;
    16: op1_14_in15 = reg_0334;
    17: op1_14_in15 = reg_0197;
    18: op1_14_in15 = reg_0318;
    19: op1_14_in15 = reg_0472;
    20: op1_14_in15 = imem04_in[27:24];
    56: op1_14_in15 = imem04_in[27:24];
    21: op1_14_in15 = reg_0142;
    22: op1_14_in15 = reg_0510;
    23: op1_14_in15 = reg_0715;
    24: op1_14_in15 = reg_0471;
    25: op1_14_in15 = reg_0288;
    26: op1_14_in15 = imem02_in[47:44];
    27: op1_14_in15 = reg_0038;
    28: op1_14_in15 = imem06_in[79:76];
    29: op1_14_in15 = reg_0196;
    30: op1_14_in15 = reg_0328;
    31: op1_14_in15 = reg_0798;
    32: op1_14_in15 = reg_0610;
    33: op1_14_in15 = imem03_in[103:100];
    34: op1_14_in15 = reg_0389;
    35: op1_14_in15 = imem04_in[111:108];
    36: op1_14_in15 = reg_0774;
    37: op1_14_in15 = reg_0130;
    40: op1_14_in15 = reg_0458;
    41: op1_14_in15 = imem04_in[99:96];
    42: op1_14_in15 = reg_0231;
    43: op1_14_in15 = reg_0160;
    44: op1_14_in15 = reg_0648;
    45: op1_14_in15 = reg_0271;
    46: op1_14_in15 = reg_0437;
    47: op1_14_in15 = reg_0357;
    48: op1_14_in15 = reg_0000;
    49: op1_14_in15 = imem02_in[67:64];
    50: op1_14_in15 = reg_0214;
    51: op1_14_in15 = imem07_in[87:84];
    52: op1_14_in15 = reg_0109;
    53: op1_14_in15 = reg_0459;
    54: op1_14_in15 = reg_0361;
    55: op1_14_in15 = reg_0570;
    57: op1_14_in15 = reg_0363;
    58: op1_14_in15 = reg_0140;
    59: op1_14_in15 = reg_0007;
    60: op1_14_in15 = reg_0732;
    62: op1_14_in15 = imem02_in[19:16];
    63: op1_14_in15 = reg_0666;
    64: op1_14_in15 = reg_0081;
    65: op1_14_in15 = imem04_in[3:0];
    66: op1_14_in15 = reg_0540;
    67: op1_14_in15 = reg_0731;
    68: op1_14_in15 = reg_0028;
    69: op1_14_in15 = imem04_in[115:112];
    70: op1_14_in15 = imem07_in[127:124];
    71: op1_14_in15 = reg_0485;
    72: op1_14_in15 = reg_0805;
    73: op1_14_in15 = reg_0679;
    74: op1_14_in15 = reg_0797;
    75: op1_14_in15 = imem07_in[51:48];
    76: op1_14_in15 = reg_0481;
    77: op1_14_in15 = reg_0594;
    78: op1_14_in15 = reg_0080;
    79: op1_14_in15 = reg_0779;
    80: op1_14_in15 = reg_0146;
    81: op1_14_in15 = reg_0753;
    82: op1_14_in15 = reg_0208;
    84: op1_14_in15 = reg_0545;
    85: op1_14_in15 = reg_0003;
    86: op1_14_in15 = reg_0195;
    87: op1_14_in15 = reg_0016;
    88: op1_14_in15 = reg_0199;
    89: op1_14_in15 = reg_0803;
    90: op1_14_in15 = reg_0584;
    91: op1_14_in15 = imem07_in[7:4];
    94: op1_14_in15 = reg_0650;
    95: op1_14_in15 = reg_0609;
    default: op1_14_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv15 = 1;
    7: op1_14_inv15 = 1;
    8: op1_14_inv15 = 1;
    9: op1_14_inv15 = 1;
    11: op1_14_inv15 = 1;
    13: op1_14_inv15 = 1;
    15: op1_14_inv15 = 1;
    17: op1_14_inv15 = 1;
    18: op1_14_inv15 = 1;
    19: op1_14_inv15 = 1;
    20: op1_14_inv15 = 1;
    21: op1_14_inv15 = 1;
    22: op1_14_inv15 = 1;
    23: op1_14_inv15 = 1;
    29: op1_14_inv15 = 1;
    31: op1_14_inv15 = 1;
    33: op1_14_inv15 = 1;
    34: op1_14_inv15 = 1;
    41: op1_14_inv15 = 1;
    43: op1_14_inv15 = 1;
    44: op1_14_inv15 = 1;
    47: op1_14_inv15 = 1;
    48: op1_14_inv15 = 1;
    52: op1_14_inv15 = 1;
    53: op1_14_inv15 = 1;
    60: op1_14_inv15 = 1;
    65: op1_14_inv15 = 1;
    66: op1_14_inv15 = 1;
    67: op1_14_inv15 = 1;
    68: op1_14_inv15 = 1;
    71: op1_14_inv15 = 1;
    72: op1_14_inv15 = 1;
    74: op1_14_inv15 = 1;
    77: op1_14_inv15 = 1;
    78: op1_14_inv15 = 1;
    81: op1_14_inv15 = 1;
    85: op1_14_inv15 = 1;
    86: op1_14_inv15 = 1;
    87: op1_14_inv15 = 1;
    88: op1_14_inv15 = 1;
    91: op1_14_inv15 = 1;
    94: op1_14_inv15 = 1;
    default: op1_14_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in16 = imem01_in[95:92];
    5: op1_14_in16 = reg_0313;
    6: op1_14_in16 = reg_0326;
    7: op1_14_in16 = reg_0809;
    8: op1_14_in16 = reg_0673;
    9: op1_14_in16 = reg_0409;
    10: op1_14_in16 = imem03_in[99:96];
    11: op1_14_in16 = reg_0286;
    12: op1_14_in16 = reg_0090;
    13: op1_14_in16 = imem04_in[63:60];
    14: op1_14_in16 = reg_0148;
    60: op1_14_in16 = reg_0148;
    15: op1_14_in16 = reg_0189;
    16: op1_14_in16 = reg_0320;
    71: op1_14_in16 = reg_0320;
    17: op1_14_in16 = imem01_in[27:24];
    18: op1_14_in16 = reg_0310;
    19: op1_14_in16 = reg_0467;
    76: op1_14_in16 = reg_0467;
    20: op1_14_in16 = imem04_in[35:32];
    21: op1_14_in16 = reg_0139;
    22: op1_14_in16 = reg_0755;
    23: op1_14_in16 = reg_0701;
    24: op1_14_in16 = reg_0468;
    25: op1_14_in16 = imem05_in[83:80];
    26: op1_14_in16 = imem02_in[51:48];
    27: op1_14_in16 = reg_0264;
    28: op1_14_in16 = imem06_in[87:84];
    29: op1_14_in16 = reg_0212;
    30: op1_14_in16 = reg_0088;
    31: op1_14_in16 = reg_0781;
    32: op1_14_in16 = reg_0613;
    33: op1_14_in16 = imem03_in[115:112];
    34: op1_14_in16 = reg_0012;
    35: op1_14_in16 = reg_0262;
    36: op1_14_in16 = reg_0317;
    37: op1_14_in16 = imem06_in[3:0];
    40: op1_14_in16 = reg_0200;
    41: op1_14_in16 = imem04_in[103:100];
    42: op1_14_in16 = reg_0238;
    43: op1_14_in16 = reg_0183;
    44: op1_14_in16 = reg_0649;
    45: op1_14_in16 = reg_0527;
    46: op1_14_in16 = reg_0448;
    47: op1_14_in16 = reg_0364;
    48: op1_14_in16 = reg_0811;
    49: op1_14_in16 = imem02_in[99:96];
    50: op1_14_in16 = reg_0191;
    51: op1_14_in16 = reg_0720;
    52: op1_14_in16 = reg_0112;
    53: op1_14_in16 = reg_0478;
    54: op1_14_in16 = reg_0323;
    55: op1_14_in16 = reg_0001;
    56: op1_14_in16 = imem04_in[39:36];
    57: op1_14_in16 = reg_0590;
    58: op1_14_in16 = reg_0131;
    59: op1_14_in16 = imem04_in[7:4];
    62: op1_14_in16 = imem02_in[31:28];
    63: op1_14_in16 = reg_0655;
    64: op1_14_in16 = reg_0080;
    65: op1_14_in16 = imem04_in[11:8];
    66: op1_14_in16 = reg_0539;
    67: op1_14_in16 = reg_0708;
    70: op1_14_in16 = reg_0708;
    68: op1_14_in16 = reg_0496;
    69: op1_14_in16 = imem04_in[119:116];
    72: op1_14_in16 = reg_0008;
    73: op1_14_in16 = reg_0687;
    74: op1_14_in16 = reg_0309;
    75: op1_14_in16 = imem07_in[59:56];
    77: op1_14_in16 = reg_0351;
    78: op1_14_in16 = reg_0530;
    79: op1_14_in16 = reg_0774;
    80: op1_14_in16 = reg_0550;
    81: op1_14_in16 = reg_0607;
    82: op1_14_in16 = reg_0186;
    84: op1_14_in16 = reg_0261;
    85: op1_14_in16 = reg_0803;
    86: op1_14_in16 = imem01_in[19:16];
    87: op1_14_in16 = imem04_in[23:20];
    88: op1_14_in16 = imem01_in[7:4];
    89: op1_14_in16 = reg_0347;
    90: op1_14_in16 = reg_0136;
    91: op1_14_in16 = imem07_in[19:16];
    94: op1_14_in16 = reg_0764;
    95: op1_14_in16 = reg_0633;
    default: op1_14_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv16 = 1;
    7: op1_14_inv16 = 1;
    8: op1_14_inv16 = 1;
    12: op1_14_inv16 = 1;
    13: op1_14_inv16 = 1;
    14: op1_14_inv16 = 1;
    15: op1_14_inv16 = 1;
    17: op1_14_inv16 = 1;
    21: op1_14_inv16 = 1;
    23: op1_14_inv16 = 1;
    26: op1_14_inv16 = 1;
    27: op1_14_inv16 = 1;
    28: op1_14_inv16 = 1;
    29: op1_14_inv16 = 1;
    31: op1_14_inv16 = 1;
    32: op1_14_inv16 = 1;
    34: op1_14_inv16 = 1;
    35: op1_14_inv16 = 1;
    36: op1_14_inv16 = 1;
    40: op1_14_inv16 = 1;
    42: op1_14_inv16 = 1;
    45: op1_14_inv16 = 1;
    46: op1_14_inv16 = 1;
    47: op1_14_inv16 = 1;
    50: op1_14_inv16 = 1;
    52: op1_14_inv16 = 1;
    55: op1_14_inv16 = 1;
    59: op1_14_inv16 = 1;
    60: op1_14_inv16 = 1;
    67: op1_14_inv16 = 1;
    68: op1_14_inv16 = 1;
    69: op1_14_inv16 = 1;
    71: op1_14_inv16 = 1;
    73: op1_14_inv16 = 1;
    76: op1_14_inv16 = 1;
    77: op1_14_inv16 = 1;
    78: op1_14_inv16 = 1;
    79: op1_14_inv16 = 1;
    80: op1_14_inv16 = 1;
    84: op1_14_inv16 = 1;
    85: op1_14_inv16 = 1;
    87: op1_14_inv16 = 1;
    88: op1_14_inv16 = 1;
    90: op1_14_inv16 = 1;
    91: op1_14_inv16 = 1;
    94: op1_14_inv16 = 1;
    95: op1_14_inv16 = 1;
    default: op1_14_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in17 = imem01_in[123:120];
    5: op1_14_in17 = reg_0404;
    6: op1_14_in17 = reg_0354;
    7: op1_14_in17 = imem04_in[119:116];
    8: op1_14_in17 = reg_0463;
    9: op1_14_in17 = reg_0315;
    69: op1_14_in17 = reg_0315;
    10: op1_14_in17 = reg_0573;
    11: op1_14_in17 = reg_0250;
    12: op1_14_in17 = reg_0087;
    13: op1_14_in17 = imem04_in[111:108];
    41: op1_14_in17 = imem04_in[111:108];
    14: op1_14_in17 = reg_0149;
    15: op1_14_in17 = reg_0204;
    16: op1_14_in17 = reg_0330;
    17: op1_14_in17 = imem01_in[43:40];
    18: op1_14_in17 = reg_0328;
    35: op1_14_in17 = reg_0328;
    19: op1_14_in17 = reg_0471;
    76: op1_14_in17 = reg_0471;
    20: op1_14_in17 = imem04_in[43:40];
    21: op1_14_in17 = reg_0129;
    22: op1_14_in17 = reg_0821;
    23: op1_14_in17 = reg_0700;
    24: op1_14_in17 = reg_0208;
    25: op1_14_in17 = imem05_in[91:88];
    26: op1_14_in17 = imem02_in[55:52];
    27: op1_14_in17 = reg_0329;
    28: op1_14_in17 = imem06_in[99:96];
    29: op1_14_in17 = imem01_in[3:0];
    30: op1_14_in17 = reg_0523;
    31: op1_14_in17 = reg_0789;
    32: op1_14_in17 = reg_0620;
    33: op1_14_in17 = imem03_in[127:124];
    34: op1_14_in17 = reg_0804;
    85: op1_14_in17 = reg_0804;
    36: op1_14_in17 = reg_0775;
    37: op1_14_in17 = imem06_in[11:8];
    40: op1_14_in17 = reg_0188;
    42: op1_14_in17 = reg_0623;
    43: op1_14_in17 = reg_0166;
    44: op1_14_in17 = reg_0644;
    45: op1_14_in17 = reg_0275;
    46: op1_14_in17 = reg_0175;
    47: op1_14_in17 = reg_0320;
    48: op1_14_in17 = reg_0001;
    49: op1_14_in17 = reg_0254;
    50: op1_14_in17 = reg_0189;
    51: op1_14_in17 = reg_0710;
    52: op1_14_in17 = reg_0668;
    53: op1_14_in17 = reg_0458;
    54: op1_14_in17 = reg_0097;
    55: op1_14_in17 = imem04_in[51:48];
    56: op1_14_in17 = imem04_in[79:76];
    57: op1_14_in17 = reg_0323;
    58: op1_14_in17 = reg_0134;
    59: op1_14_in17 = imem04_in[19:16];
    65: op1_14_in17 = imem04_in[19:16];
    60: op1_14_in17 = reg_0135;
    62: op1_14_in17 = reg_0485;
    63: op1_14_in17 = reg_0114;
    64: op1_14_in17 = reg_0540;
    78: op1_14_in17 = reg_0540;
    66: op1_14_in17 = reg_0094;
    67: op1_14_in17 = reg_0715;
    68: op1_14_in17 = imem01_in[15:12];
    70: op1_14_in17 = reg_0711;
    71: op1_14_in17 = reg_0345;
    81: op1_14_in17 = reg_0345;
    72: op1_14_in17 = reg_0015;
    73: op1_14_in17 = reg_0622;
    74: op1_14_in17 = reg_0786;
    75: op1_14_in17 = imem07_in[67:64];
    77: op1_14_in17 = reg_0533;
    79: op1_14_in17 = reg_0776;
    80: op1_14_in17 = reg_0793;
    82: op1_14_in17 = reg_0198;
    84: op1_14_in17 = reg_0331;
    86: op1_14_in17 = imem01_in[27:24];
    87: op1_14_in17 = imem04_in[59:56];
    88: op1_14_in17 = imem01_in[35:32];
    89: op1_14_in17 = reg_0350;
    90: op1_14_in17 = reg_0756;
    91: op1_14_in17 = imem07_in[35:32];
    94: op1_14_in17 = imem07_in[31:28];
    95: op1_14_in17 = reg_0661;
    default: op1_14_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv17 = 1;
    9: op1_14_inv17 = 1;
    11: op1_14_inv17 = 1;
    12: op1_14_inv17 = 1;
    14: op1_14_inv17 = 1;
    15: op1_14_inv17 = 1;
    16: op1_14_inv17 = 1;
    18: op1_14_inv17 = 1;
    20: op1_14_inv17 = 1;
    22: op1_14_inv17 = 1;
    23: op1_14_inv17 = 1;
    24: op1_14_inv17 = 1;
    25: op1_14_inv17 = 1;
    27: op1_14_inv17 = 1;
    29: op1_14_inv17 = 1;
    31: op1_14_inv17 = 1;
    32: op1_14_inv17 = 1;
    35: op1_14_inv17 = 1;
    36: op1_14_inv17 = 1;
    37: op1_14_inv17 = 1;
    40: op1_14_inv17 = 1;
    41: op1_14_inv17 = 1;
    43: op1_14_inv17 = 1;
    45: op1_14_inv17 = 1;
    47: op1_14_inv17 = 1;
    49: op1_14_inv17 = 1;
    52: op1_14_inv17 = 1;
    55: op1_14_inv17 = 1;
    57: op1_14_inv17 = 1;
    58: op1_14_inv17 = 1;
    59: op1_14_inv17 = 1;
    60: op1_14_inv17 = 1;
    62: op1_14_inv17 = 1;
    65: op1_14_inv17 = 1;
    67: op1_14_inv17 = 1;
    68: op1_14_inv17 = 1;
    69: op1_14_inv17 = 1;
    70: op1_14_inv17 = 1;
    73: op1_14_inv17 = 1;
    77: op1_14_inv17 = 1;
    78: op1_14_inv17 = 1;
    80: op1_14_inv17 = 1;
    81: op1_14_inv17 = 1;
    86: op1_14_inv17 = 1;
    87: op1_14_inv17 = 1;
    89: op1_14_inv17 = 1;
    90: op1_14_inv17 = 1;
    91: op1_14_inv17 = 1;
    94: op1_14_inv17 = 1;
    95: op1_14_inv17 = 1;
    default: op1_14_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in18 = reg_0517;
    5: op1_14_in18 = reg_0315;
    6: op1_14_in18 = reg_0359;
    7: op1_14_in18 = reg_0530;
    8: op1_14_in18 = reg_0465;
    9: op1_14_in18 = reg_0034;
    10: op1_14_in18 = reg_0395;
    11: op1_14_in18 = reg_0256;
    12: op1_14_in18 = reg_0073;
    13: op1_14_in18 = reg_0528;
    14: op1_14_in18 = reg_0145;
    15: op1_14_in18 = reg_0205;
    16: op1_14_in18 = reg_0089;
    17: op1_14_in18 = reg_0229;
    18: op1_14_in18 = reg_0083;
    19: op1_14_in18 = reg_0478;
    20: op1_14_in18 = imem04_in[47:44];
    21: op1_14_in18 = reg_0134;
    22: op1_14_in18 = reg_0511;
    23: op1_14_in18 = reg_0441;
    24: op1_14_in18 = reg_0191;
    25: op1_14_in18 = reg_0781;
    26: op1_14_in18 = imem02_in[91:88];
    27: op1_14_in18 = reg_0311;
    28: op1_14_in18 = imem06_in[103:100];
    29: op1_14_in18 = imem01_in[63:60];
    30: op1_14_in18 = reg_0551;
    31: op1_14_in18 = reg_0494;
    32: op1_14_in18 = reg_0616;
    33: op1_14_in18 = reg_0598;
    34: op1_14_in18 = reg_0810;
    35: op1_14_in18 = reg_0542;
    36: op1_14_in18 = reg_0329;
    37: op1_14_in18 = imem06_in[31:28];
    40: op1_14_in18 = reg_0196;
    76: op1_14_in18 = reg_0196;
    82: op1_14_in18 = reg_0196;
    41: op1_14_in18 = reg_0066;
    42: op1_14_in18 = reg_0233;
    43: op1_14_in18 = reg_0185;
    44: op1_14_in18 = imem02_in[59:56];
    45: op1_14_in18 = reg_0224;
    46: op1_14_in18 = reg_0180;
    47: op1_14_in18 = reg_0343;
    48: op1_14_in18 = reg_0801;
    49: op1_14_in18 = reg_0654;
    50: op1_14_in18 = reg_0211;
    51: op1_14_in18 = reg_0717;
    52: op1_14_in18 = reg_0649;
    53: op1_14_in18 = reg_0210;
    54: op1_14_in18 = reg_0402;
    55: op1_14_in18 = imem04_in[71:68];
    56: op1_14_in18 = reg_0043;
    57: op1_14_in18 = reg_0518;
    71: op1_14_in18 = reg_0518;
    58: op1_14_in18 = imem06_in[7:4];
    59: op1_14_in18 = imem04_in[31:28];
    60: op1_14_in18 = reg_0146;
    62: op1_14_in18 = reg_0358;
    63: op1_14_in18 = reg_0352;
    64: op1_14_in18 = reg_0098;
    90: op1_14_in18 = reg_0098;
    65: op1_14_in18 = imem04_in[39:36];
    66: op1_14_in18 = imem03_in[123:120];
    67: op1_14_in18 = reg_0711;
    68: op1_14_in18 = imem01_in[43:40];
    69: op1_14_in18 = reg_0560;
    70: op1_14_in18 = reg_0067;
    72: op1_14_in18 = reg_0009;
    73: op1_14_in18 = reg_0774;
    74: op1_14_in18 = reg_0236;
    75: op1_14_in18 = imem07_in[87:84];
    77: op1_14_in18 = reg_0081;
    78: op1_14_in18 = reg_0770;
    79: op1_14_in18 = imem05_in[3:0];
    80: op1_14_in18 = reg_0782;
    81: op1_14_in18 = reg_0406;
    84: op1_14_in18 = reg_0303;
    85: op1_14_in18 = reg_0800;
    86: op1_14_in18 = imem01_in[95:92];
    87: op1_14_in18 = imem04_in[67:64];
    88: op1_14_in18 = imem01_in[103:100];
    89: op1_14_in18 = reg_0223;
    91: op1_14_in18 = reg_0391;
    94: op1_14_in18 = imem07_in[95:92];
    95: op1_14_in18 = imem07_in[23:20];
    default: op1_14_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_14_inv18 = 1;
    8: op1_14_inv18 = 1;
    14: op1_14_inv18 = 1;
    15: op1_14_inv18 = 1;
    16: op1_14_inv18 = 1;
    20: op1_14_inv18 = 1;
    21: op1_14_inv18 = 1;
    25: op1_14_inv18 = 1;
    27: op1_14_inv18 = 1;
    28: op1_14_inv18 = 1;
    30: op1_14_inv18 = 1;
    31: op1_14_inv18 = 1;
    33: op1_14_inv18 = 1;
    37: op1_14_inv18 = 1;
    41: op1_14_inv18 = 1;
    44: op1_14_inv18 = 1;
    46: op1_14_inv18 = 1;
    48: op1_14_inv18 = 1;
    49: op1_14_inv18 = 1;
    50: op1_14_inv18 = 1;
    51: op1_14_inv18 = 1;
    52: op1_14_inv18 = 1;
    55: op1_14_inv18 = 1;
    57: op1_14_inv18 = 1;
    58: op1_14_inv18 = 1;
    62: op1_14_inv18 = 1;
    65: op1_14_inv18 = 1;
    71: op1_14_inv18 = 1;
    72: op1_14_inv18 = 1;
    77: op1_14_inv18 = 1;
    78: op1_14_inv18 = 1;
    79: op1_14_inv18 = 1;
    82: op1_14_inv18 = 1;
    85: op1_14_inv18 = 1;
    86: op1_14_inv18 = 1;
    87: op1_14_inv18 = 1;
    89: op1_14_inv18 = 1;
    default: op1_14_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in19 = reg_0518;
    5: op1_14_in19 = reg_0337;
    6: op1_14_in19 = reg_0318;
    7: op1_14_in19 = reg_0528;
    8: op1_14_in19 = reg_0464;
    9: op1_14_in19 = reg_0752;
    10: op1_14_in19 = reg_0360;
    11: op1_14_in19 = reg_0258;
    12: op1_14_in19 = reg_0079;
    13: op1_14_in19 = reg_0555;
    14: op1_14_in19 = reg_0140;
    15: op1_14_in19 = reg_0202;
    16: op1_14_in19 = reg_0085;
    17: op1_14_in19 = reg_0227;
    18: op1_14_in19 = reg_0088;
    56: op1_14_in19 = reg_0088;
    19: op1_14_in19 = reg_0214;
    20: op1_14_in19 = imem04_in[55:52];
    21: op1_14_in19 = imem06_in[39:36];
    22: op1_14_in19 = reg_0237;
    23: op1_14_in19 = reg_0430;
    24: op1_14_in19 = reg_0209;
    25: op1_14_in19 = reg_0309;
    26: op1_14_in19 = imem02_in[107:104];
    27: op1_14_in19 = reg_0586;
    28: op1_14_in19 = imem06_in[127:124];
    29: op1_14_in19 = imem01_in[67:64];
    30: op1_14_in19 = reg_0556;
    31: op1_14_in19 = reg_0780;
    32: op1_14_in19 = reg_0611;
    33: op1_14_in19 = reg_0749;
    34: op1_14_in19 = reg_0004;
    35: op1_14_in19 = reg_0055;
    36: op1_14_in19 = reg_0311;
    37: op1_14_in19 = imem06_in[47:44];
    40: op1_14_in19 = reg_0195;
    82: op1_14_in19 = reg_0195;
    41: op1_14_in19 = reg_0067;
    42: op1_14_in19 = reg_0426;
    44: op1_14_in19 = reg_0362;
    45: op1_14_in19 = reg_0086;
    74: op1_14_in19 = reg_0086;
    46: op1_14_in19 = reg_0177;
    47: op1_14_in19 = reg_0347;
    48: op1_14_in19 = reg_0008;
    49: op1_14_in19 = reg_0660;
    50: op1_14_in19 = reg_0201;
    51: op1_14_in19 = reg_0718;
    52: op1_14_in19 = reg_0322;
    53: op1_14_in19 = reg_0204;
    54: op1_14_in19 = reg_0578;
    55: op1_14_in19 = imem04_in[83:80];
    57: op1_14_in19 = reg_0541;
    58: op1_14_in19 = imem06_in[55:52];
    59: op1_14_in19 = imem04_in[39:36];
    60: op1_14_in19 = reg_0154;
    62: op1_14_in19 = reg_0359;
    63: op1_14_in19 = reg_0345;
    64: op1_14_in19 = reg_0740;
    90: op1_14_in19 = reg_0740;
    65: op1_14_in19 = imem04_in[47:44];
    66: op1_14_in19 = imem03_in[127:124];
    67: op1_14_in19 = reg_0701;
    68: op1_14_in19 = imem01_in[71:68];
    69: op1_14_in19 = reg_0083;
    70: op1_14_in19 = reg_0333;
    71: op1_14_in19 = reg_0082;
    72: op1_14_in19 = reg_0809;
    73: op1_14_in19 = reg_0259;
    75: op1_14_in19 = imem07_in[91:88];
    76: op1_14_in19 = imem01_in[19:16];
    77: op1_14_in19 = reg_0770;
    78: op1_14_in19 = imem03_in[19:16];
    79: op1_14_in19 = imem05_in[23:20];
    80: op1_14_in19 = reg_0326;
    81: op1_14_in19 = reg_0081;
    84: op1_14_in19 = reg_0308;
    85: op1_14_in19 = reg_0810;
    86: op1_14_in19 = reg_0520;
    87: op1_14_in19 = imem04_in[91:88];
    88: op1_14_in19 = imem01_in[127:124];
    89: op1_14_in19 = reg_0338;
    91: op1_14_in19 = reg_0726;
    94: op1_14_in19 = imem07_in[119:116];
    95: op1_14_in19 = imem07_in[79:76];
    default: op1_14_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv19 = 1;
    6: op1_14_inv19 = 1;
    7: op1_14_inv19 = 1;
    9: op1_14_inv19 = 1;
    10: op1_14_inv19 = 1;
    11: op1_14_inv19 = 1;
    14: op1_14_inv19 = 1;
    15: op1_14_inv19 = 1;
    16: op1_14_inv19 = 1;
    20: op1_14_inv19 = 1;
    21: op1_14_inv19 = 1;
    22: op1_14_inv19 = 1;
    24: op1_14_inv19 = 1;
    25: op1_14_inv19 = 1;
    28: op1_14_inv19 = 1;
    29: op1_14_inv19 = 1;
    30: op1_14_inv19 = 1;
    33: op1_14_inv19 = 1;
    36: op1_14_inv19 = 1;
    37: op1_14_inv19 = 1;
    40: op1_14_inv19 = 1;
    41: op1_14_inv19 = 1;
    44: op1_14_inv19 = 1;
    46: op1_14_inv19 = 1;
    47: op1_14_inv19 = 1;
    48: op1_14_inv19 = 1;
    49: op1_14_inv19 = 1;
    50: op1_14_inv19 = 1;
    52: op1_14_inv19 = 1;
    53: op1_14_inv19 = 1;
    56: op1_14_inv19 = 1;
    57: op1_14_inv19 = 1;
    64: op1_14_inv19 = 1;
    65: op1_14_inv19 = 1;
    69: op1_14_inv19 = 1;
    70: op1_14_inv19 = 1;
    71: op1_14_inv19 = 1;
    78: op1_14_inv19 = 1;
    79: op1_14_inv19 = 1;
    82: op1_14_inv19 = 1;
    87: op1_14_inv19 = 1;
    88: op1_14_inv19 = 1;
    89: op1_14_inv19 = 1;
    90: op1_14_inv19 = 1;
    91: op1_14_inv19 = 1;
    default: op1_14_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in20 = reg_0498;
    5: op1_14_in20 = reg_0027;
    6: op1_14_in20 = reg_0330;
    7: op1_14_in20 = reg_0546;
    8: op1_14_in20 = reg_0469;
    9: op1_14_in20 = reg_0038;
    10: op1_14_in20 = reg_0319;
    11: op1_14_in20 = reg_0798;
    12: op1_14_in20 = imem03_in[19:16];
    13: op1_14_in20 = reg_0304;
    14: op1_14_in20 = reg_0134;
    15: op1_14_in20 = reg_0199;
    16: op1_14_in20 = reg_0077;
    17: op1_14_in20 = reg_0516;
    18: op1_14_in20 = reg_0089;
    19: op1_14_in20 = reg_0191;
    20: op1_14_in20 = imem04_in[59:56];
    21: op1_14_in20 = imem06_in[59:56];
    22: op1_14_in20 = reg_0041;
    23: op1_14_in20 = reg_0436;
    24: op1_14_in20 = reg_0207;
    25: op1_14_in20 = reg_0279;
    26: op1_14_in20 = reg_0642;
    27: op1_14_in20 = reg_0592;
    28: op1_14_in20 = reg_0753;
    29: op1_14_in20 = imem01_in[87:84];
    30: op1_14_in20 = reg_0308;
    31: op1_14_in20 = reg_0786;
    32: op1_14_in20 = reg_0627;
    33: op1_14_in20 = reg_0392;
    34: op1_14_in20 = imem04_in[11:8];
    35: op1_14_in20 = reg_0555;
    55: op1_14_in20 = reg_0555;
    56: op1_14_in20 = reg_0555;
    36: op1_14_in20 = imem06_in[3:0];
    37: op1_14_in20 = imem06_in[115:112];
    40: op1_14_in20 = reg_0508;
    41: op1_14_in20 = reg_0070;
    42: op1_14_in20 = reg_0704;
    44: op1_14_in20 = reg_0229;
    45: op1_14_in20 = reg_0132;
    46: op1_14_in20 = reg_0185;
    47: op1_14_in20 = reg_0533;
    48: op1_14_in20 = reg_0257;
    49: op1_14_in20 = reg_0656;
    50: op1_14_in20 = reg_0213;
    53: op1_14_in20 = reg_0213;
    51: op1_14_in20 = reg_0701;
    52: op1_14_in20 = reg_0778;
    86: op1_14_in20 = reg_0778;
    54: op1_14_in20 = reg_0311;
    57: op1_14_in20 = reg_0096;
    81: op1_14_in20 = reg_0096;
    58: op1_14_in20 = imem06_in[79:76];
    59: op1_14_in20 = imem04_in[43:40];
    60: op1_14_in20 = reg_0039;
    62: op1_14_in20 = reg_0342;
    63: op1_14_in20 = reg_0565;
    64: op1_14_in20 = imem03_in[35:32];
    65: op1_14_in20 = imem04_in[79:76];
    66: op1_14_in20 = reg_0599;
    67: op1_14_in20 = reg_0064;
    68: op1_14_in20 = imem01_in[79:76];
    69: op1_14_in20 = reg_0523;
    70: op1_14_in20 = reg_0435;
    71: op1_14_in20 = reg_0740;
    72: op1_14_in20 = imem04_in[15:12];
    73: op1_14_in20 = reg_0640;
    74: op1_14_in20 = reg_0148;
    75: op1_14_in20 = imem07_in[103:100];
    76: op1_14_in20 = imem01_in[39:36];
    77: op1_14_in20 = reg_0757;
    78: op1_14_in20 = imem03_in[43:40];
    79: op1_14_in20 = imem05_in[35:32];
    80: op1_14_in20 = reg_0309;
    82: op1_14_in20 = imem01_in[7:4];
    84: op1_14_in20 = reg_0280;
    85: op1_14_in20 = imem04_in[27:24];
    87: op1_14_in20 = imem04_in[127:124];
    88: op1_14_in20 = reg_0506;
    89: op1_14_in20 = reg_0318;
    90: op1_14_in20 = imem03_in[15:12];
    91: op1_14_in20 = reg_0166;
    94: op1_14_in20 = reg_0167;
    95: op1_14_in20 = imem07_in[111:108];
    default: op1_14_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv20 = 1;
    7: op1_14_inv20 = 1;
    10: op1_14_inv20 = 1;
    11: op1_14_inv20 = 1;
    17: op1_14_inv20 = 1;
    18: op1_14_inv20 = 1;
    19: op1_14_inv20 = 1;
    21: op1_14_inv20 = 1;
    25: op1_14_inv20 = 1;
    26: op1_14_inv20 = 1;
    28: op1_14_inv20 = 1;
    30: op1_14_inv20 = 1;
    33: op1_14_inv20 = 1;
    34: op1_14_inv20 = 1;
    35: op1_14_inv20 = 1;
    37: op1_14_inv20 = 1;
    40: op1_14_inv20 = 1;
    41: op1_14_inv20 = 1;
    44: op1_14_inv20 = 1;
    46: op1_14_inv20 = 1;
    50: op1_14_inv20 = 1;
    52: op1_14_inv20 = 1;
    53: op1_14_inv20 = 1;
    57: op1_14_inv20 = 1;
    58: op1_14_inv20 = 1;
    59: op1_14_inv20 = 1;
    60: op1_14_inv20 = 1;
    62: op1_14_inv20 = 1;
    65: op1_14_inv20 = 1;
    66: op1_14_inv20 = 1;
    67: op1_14_inv20 = 1;
    68: op1_14_inv20 = 1;
    69: op1_14_inv20 = 1;
    70: op1_14_inv20 = 1;
    73: op1_14_inv20 = 1;
    74: op1_14_inv20 = 1;
    78: op1_14_inv20 = 1;
    79: op1_14_inv20 = 1;
    80: op1_14_inv20 = 1;
    81: op1_14_inv20 = 1;
    84: op1_14_inv20 = 1;
    85: op1_14_inv20 = 1;
    86: op1_14_inv20 = 1;
    88: op1_14_inv20 = 1;
    89: op1_14_inv20 = 1;
    90: op1_14_inv20 = 1;
    91: op1_14_inv20 = 1;
    94: op1_14_inv20 = 1;
    default: op1_14_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in21 = reg_0233;
    5: op1_14_in21 = reg_0020;
    6: op1_14_in21 = reg_0363;
    7: op1_14_in21 = reg_0559;
    8: op1_14_in21 = reg_0476;
    9: op1_14_in21 = imem07_in[11:8];
    10: op1_14_in21 = reg_0312;
    11: op1_14_in21 = reg_0488;
    12: op1_14_in21 = imem03_in[31:28];
    16: op1_14_in21 = imem03_in[31:28];
    13: op1_14_in21 = reg_0061;
    14: op1_14_in21 = imem06_in[39:36];
    15: op1_14_in21 = imem01_in[15:12];
    17: op1_14_in21 = reg_0235;
    18: op1_14_in21 = reg_0090;
    19: op1_14_in21 = reg_0189;
    20: op1_14_in21 = imem04_in[87:84];
    65: op1_14_in21 = imem04_in[87:84];
    21: op1_14_in21 = imem06_in[103:100];
    22: op1_14_in21 = reg_0243;
    23: op1_14_in21 = reg_0423;
    24: op1_14_in21 = reg_0197;
    25: op1_14_in21 = reg_0276;
    26: op1_14_in21 = reg_0654;
    27: op1_14_in21 = reg_0591;
    28: op1_14_in21 = reg_0040;
    29: op1_14_in21 = reg_0501;
    30: op1_14_in21 = reg_0054;
    31: op1_14_in21 = reg_0225;
    32: op1_14_in21 = reg_0615;
    33: op1_14_in21 = reg_0376;
    34: op1_14_in21 = imem04_in[19:16];
    35: op1_14_in21 = reg_0308;
    36: op1_14_in21 = imem06_in[51:48];
    37: op1_14_in21 = reg_0604;
    40: op1_14_in21 = reg_0336;
    41: op1_14_in21 = reg_0064;
    42: op1_14_in21 = reg_0726;
    44: op1_14_in21 = reg_0341;
    45: op1_14_in21 = reg_0147;
    46: op1_14_in21 = reg_0176;
    47: op1_14_in21 = reg_0095;
    48: op1_14_in21 = reg_0066;
    49: op1_14_in21 = reg_0346;
    50: op1_14_in21 = reg_0196;
    51: op1_14_in21 = reg_0334;
    52: op1_14_in21 = reg_0550;
    53: op1_14_in21 = reg_0205;
    54: op1_14_in21 = imem03_in[3:0];
    71: op1_14_in21 = imem03_in[3:0];
    55: op1_14_in21 = reg_0500;
    56: op1_14_in21 = reg_0523;
    57: op1_14_in21 = reg_0531;
    58: op1_14_in21 = imem06_in[111:108];
    59: op1_14_in21 = imem04_in[67:64];
    60: op1_14_in21 = reg_0818;
    62: op1_14_in21 = reg_0343;
    63: op1_14_in21 = reg_0514;
    64: op1_14_in21 = imem03_in[39:36];
    66: op1_14_in21 = reg_0338;
    67: op1_14_in21 = reg_0295;
    68: op1_14_in21 = imem01_in[95:92];
    69: op1_14_in21 = reg_0058;
    70: op1_14_in21 = reg_0185;
    72: op1_14_in21 = imem04_in[27:24];
    73: op1_14_in21 = reg_0091;
    74: op1_14_in21 = reg_0785;
    75: op1_14_in21 = imem07_in[107:104];
    76: op1_14_in21 = imem01_in[83:80];
    77: op1_14_in21 = reg_0094;
    78: op1_14_in21 = imem03_in[71:68];
    79: op1_14_in21 = imem05_in[115:112];
    80: op1_14_in21 = reg_0491;
    81: op1_14_in21 = reg_0540;
    82: op1_14_in21 = imem01_in[19:16];
    84: op1_14_in21 = reg_0616;
    85: op1_14_in21 = imem04_in[35:32];
    86: op1_14_in21 = reg_0388;
    87: op1_14_in21 = reg_0060;
    88: op1_14_in21 = reg_0424;
    89: op1_14_in21 = reg_0799;
    90: op1_14_in21 = imem03_in[27:24];
    91: op1_14_in21 = reg_0164;
    94: op1_14_in21 = reg_0382;
    95: op1_14_in21 = imem07_in[115:112];
    default: op1_14_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv21 = 1;
    6: op1_14_inv21 = 1;
    8: op1_14_inv21 = 1;
    10: op1_14_inv21 = 1;
    12: op1_14_inv21 = 1;
    14: op1_14_inv21 = 1;
    15: op1_14_inv21 = 1;
    17: op1_14_inv21 = 1;
    18: op1_14_inv21 = 1;
    19: op1_14_inv21 = 1;
    20: op1_14_inv21 = 1;
    22: op1_14_inv21 = 1;
    23: op1_14_inv21 = 1;
    24: op1_14_inv21 = 1;
    28: op1_14_inv21 = 1;
    29: op1_14_inv21 = 1;
    31: op1_14_inv21 = 1;
    33: op1_14_inv21 = 1;
    34: op1_14_inv21 = 1;
    36: op1_14_inv21 = 1;
    42: op1_14_inv21 = 1;
    47: op1_14_inv21 = 1;
    53: op1_14_inv21 = 1;
    54: op1_14_inv21 = 1;
    55: op1_14_inv21 = 1;
    56: op1_14_inv21 = 1;
    59: op1_14_inv21 = 1;
    60: op1_14_inv21 = 1;
    62: op1_14_inv21 = 1;
    63: op1_14_inv21 = 1;
    64: op1_14_inv21 = 1;
    65: op1_14_inv21 = 1;
    67: op1_14_inv21 = 1;
    68: op1_14_inv21 = 1;
    73: op1_14_inv21 = 1;
    74: op1_14_inv21 = 1;
    75: op1_14_inv21 = 1;
    76: op1_14_inv21 = 1;
    77: op1_14_inv21 = 1;
    78: op1_14_inv21 = 1;
    80: op1_14_inv21 = 1;
    81: op1_14_inv21 = 1;
    82: op1_14_inv21 = 1;
    85: op1_14_inv21 = 1;
    88: op1_14_inv21 = 1;
    90: op1_14_inv21 = 1;
    default: op1_14_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in22 = reg_0228;
    5: op1_14_in22 = reg_0024;
    6: op1_14_in22 = reg_0086;
    7: op1_14_in22 = reg_0531;
    8: op1_14_in22 = reg_0466;
    9: op1_14_in22 = imem07_in[43:40];
    10: op1_14_in22 = reg_0000;
    11: op1_14_in22 = reg_0491;
    12: op1_14_in22 = imem03_in[35:32];
    13: op1_14_in22 = reg_0047;
    14: op1_14_in22 = imem06_in[87:84];
    15: op1_14_in22 = imem01_in[59:56];
    16: op1_14_in22 = imem03_in[87:84];
    17: op1_14_in22 = reg_0505;
    18: op1_14_in22 = reg_0091;
    19: op1_14_in22 = reg_0211;
    20: op1_14_in22 = imem04_in[91:88];
    21: op1_14_in22 = imem06_in[123:120];
    22: op1_14_in22 = reg_0122;
    23: op1_14_in22 = reg_0440;
    24: op1_14_in22 = reg_0499;
    33: op1_14_in22 = reg_0499;
    25: op1_14_in22 = reg_0224;
    48: op1_14_in22 = reg_0224;
    26: op1_14_in22 = reg_0656;
    27: op1_14_in22 = reg_0585;
    28: op1_14_in22 = reg_0036;
    29: op1_14_in22 = reg_0512;
    30: op1_14_in22 = reg_0283;
    31: op1_14_in22 = reg_0309;
    32: op1_14_in22 = reg_0612;
    34: op1_14_in22 = imem04_in[99:96];
    35: op1_14_in22 = reg_0280;
    36: op1_14_in22 = imem07_in[31:28];
    37: op1_14_in22 = reg_0624;
    40: op1_14_in22 = reg_0515;
    41: op1_14_in22 = imem05_in[15:12];
    42: op1_14_in22 = reg_0714;
    44: op1_14_in22 = reg_0359;
    45: op1_14_in22 = reg_0150;
    46: op1_14_in22 = reg_0184;
    47: op1_14_in22 = reg_0769;
    49: op1_14_in22 = reg_0344;
    50: op1_14_in22 = imem01_in[39:36];
    51: op1_14_in22 = reg_0441;
    52: op1_14_in22 = reg_0321;
    53: op1_14_in22 = reg_0192;
    54: op1_14_in22 = imem03_in[7:4];
    55: op1_14_in22 = reg_0303;
    56: op1_14_in22 = reg_0429;
    57: op1_14_in22 = imem03_in[11:8];
    58: op1_14_in22 = reg_0289;
    59: op1_14_in22 = imem04_in[95:92];
    60: op1_14_in22 = reg_0111;
    62: op1_14_in22 = reg_0092;
    63: op1_14_in22 = reg_0314;
    64: op1_14_in22 = imem03_in[43:40];
    65: op1_14_in22 = imem04_in[107:104];
    66: op1_14_in22 = reg_0493;
    67: op1_14_in22 = reg_0446;
    68: op1_14_in22 = reg_0418;
    69: op1_14_in22 = reg_0500;
    70: op1_14_in22 = reg_0171;
    71: op1_14_in22 = imem03_in[83:80];
    78: op1_14_in22 = imem03_in[83:80];
    72: op1_14_in22 = imem04_in[59:56];
    73: op1_14_in22 = reg_0136;
    74: op1_14_in22 = reg_0765;
    75: op1_14_in22 = imem07_in[119:116];
    95: op1_14_in22 = imem07_in[119:116];
    76: op1_14_in22 = imem01_in[115:112];
    77: op1_14_in22 = imem03_in[3:0];
    79: op1_14_in22 = reg_0227;
    80: op1_14_in22 = reg_0276;
    81: op1_14_in22 = reg_0535;
    82: op1_14_in22 = imem01_in[23:20];
    84: op1_14_in22 = reg_0503;
    85: op1_14_in22 = imem04_in[43:40];
    86: op1_14_in22 = reg_0225;
    87: op1_14_in22 = reg_0079;
    88: op1_14_in22 = reg_0243;
    89: op1_14_in22 = reg_0572;
    90: op1_14_in22 = imem03_in[47:44];
    91: op1_14_in22 = reg_0103;
    94: op1_14_in22 = reg_0708;
    default: op1_14_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv22 = 1;
    5: op1_14_inv22 = 1;
    6: op1_14_inv22 = 1;
    9: op1_14_inv22 = 1;
    12: op1_14_inv22 = 1;
    14: op1_14_inv22 = 1;
    16: op1_14_inv22 = 1;
    24: op1_14_inv22 = 1;
    26: op1_14_inv22 = 1;
    29: op1_14_inv22 = 1;
    30: op1_14_inv22 = 1;
    31: op1_14_inv22 = 1;
    34: op1_14_inv22 = 1;
    35: op1_14_inv22 = 1;
    36: op1_14_inv22 = 1;
    45: op1_14_inv22 = 1;
    46: op1_14_inv22 = 1;
    51: op1_14_inv22 = 1;
    52: op1_14_inv22 = 1;
    54: op1_14_inv22 = 1;
    57: op1_14_inv22 = 1;
    60: op1_14_inv22 = 1;
    62: op1_14_inv22 = 1;
    63: op1_14_inv22 = 1;
    64: op1_14_inv22 = 1;
    65: op1_14_inv22 = 1;
    67: op1_14_inv22 = 1;
    69: op1_14_inv22 = 1;
    74: op1_14_inv22 = 1;
    81: op1_14_inv22 = 1;
    87: op1_14_inv22 = 1;
    88: op1_14_inv22 = 1;
    89: op1_14_inv22 = 1;
    90: op1_14_inv22 = 1;
    94: op1_14_inv22 = 1;
    95: op1_14_inv22 = 1;
    default: op1_14_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in23 = reg_0221;
    5: op1_14_in23 = reg_0023;
    6: op1_14_in23 = reg_0090;
    7: op1_14_in23 = reg_0556;
    69: op1_14_in23 = reg_0556;
    8: op1_14_in23 = reg_0472;
    9: op1_14_in23 = imem07_in[55:52];
    10: op1_14_in23 = reg_0800;
    11: op1_14_in23 = reg_0793;
    12: op1_14_in23 = imem03_in[83:80];
    13: op1_14_in23 = reg_0078;
    14: op1_14_in23 = imem06_in[123:120];
    15: op1_14_in23 = imem01_in[63:60];
    16: op1_14_in23 = imem03_in[99:96];
    17: op1_14_in23 = reg_0234;
    18: op1_14_in23 = reg_0084;
    19: op1_14_in23 = reg_0196;
    20: op1_14_in23 = reg_0543;
    21: op1_14_in23 = reg_0614;
    22: op1_14_in23 = reg_0125;
    23: op1_14_in23 = reg_0444;
    67: op1_14_in23 = reg_0444;
    24: op1_14_in23 = reg_0322;
    25: op1_14_in23 = reg_0272;
    26: op1_14_in23 = reg_0640;
    27: op1_14_in23 = reg_0576;
    28: op1_14_in23 = reg_0037;
    29: op1_14_in23 = reg_0557;
    30: op1_14_in23 = reg_0280;
    55: op1_14_in23 = reg_0280;
    31: op1_14_in23 = reg_0226;
    32: op1_14_in23 = reg_0408;
    33: op1_14_in23 = reg_0386;
    34: op1_14_in23 = reg_0316;
    35: op1_14_in23 = reg_0302;
    36: op1_14_in23 = imem07_in[51:48];
    37: op1_14_in23 = reg_0631;
    40: op1_14_in23 = imem01_in[95:92];
    41: op1_14_in23 = imem05_in[35:32];
    42: op1_14_in23 = reg_0707;
    44: op1_14_in23 = reg_0073;
    45: op1_14_in23 = reg_0128;
    46: op1_14_in23 = reg_0437;
    47: op1_14_in23 = reg_0770;
    48: op1_14_in23 = reg_0353;
    49: op1_14_in23 = reg_0358;
    50: op1_14_in23 = imem01_in[43:40];
    51: op1_14_in23 = reg_0443;
    52: op1_14_in23 = reg_0232;
    53: op1_14_in23 = imem01_in[3:0];
    54: op1_14_in23 = imem03_in[15:12];
    56: op1_14_in23 = reg_0432;
    57: op1_14_in23 = imem03_in[23:20];
    58: op1_14_in23 = reg_0401;
    59: op1_14_in23 = imem04_in[119:116];
    60: op1_14_in23 = reg_0005;
    62: op1_14_in23 = reg_0314;
    63: op1_14_in23 = reg_0096;
    64: op1_14_in23 = imem03_in[51:48];
    65: op1_14_in23 = imem04_in[127:124];
    66: op1_14_in23 = reg_0575;
    68: op1_14_in23 = reg_0511;
    71: op1_14_in23 = imem03_in[87:84];
    72: op1_14_in23 = imem04_in[67:64];
    73: op1_14_in23 = reg_0277;
    74: op1_14_in23 = imem06_in[63:60];
    75: op1_14_in23 = imem07_in[123:120];
    95: op1_14_in23 = imem07_in[123:120];
    76: op1_14_in23 = reg_0376;
    77: op1_14_in23 = imem03_in[63:60];
    78: op1_14_in23 = reg_0582;
    79: op1_14_in23 = reg_0641;
    80: op1_14_in23 = reg_0288;
    81: op1_14_in23 = reg_0539;
    82: op1_14_in23 = imem01_in[27:24];
    84: op1_14_in23 = reg_0431;
    85: op1_14_in23 = imem04_in[63:60];
    86: op1_14_in23 = reg_0306;
    87: op1_14_in23 = reg_0297;
    88: op1_14_in23 = reg_0420;
    89: op1_14_in23 = reg_0321;
    90: op1_14_in23 = reg_0573;
    91: op1_14_in23 = reg_0061;
    94: op1_14_in23 = reg_0158;
    default: op1_14_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv23 = 1;
    7: op1_14_inv23 = 1;
    8: op1_14_inv23 = 1;
    10: op1_14_inv23 = 1;
    11: op1_14_inv23 = 1;
    12: op1_14_inv23 = 1;
    13: op1_14_inv23 = 1;
    14: op1_14_inv23 = 1;
    15: op1_14_inv23 = 1;
    16: op1_14_inv23 = 1;
    18: op1_14_inv23 = 1;
    20: op1_14_inv23 = 1;
    26: op1_14_inv23 = 1;
    28: op1_14_inv23 = 1;
    29: op1_14_inv23 = 1;
    32: op1_14_inv23 = 1;
    35: op1_14_inv23 = 1;
    36: op1_14_inv23 = 1;
    40: op1_14_inv23 = 1;
    41: op1_14_inv23 = 1;
    44: op1_14_inv23 = 1;
    50: op1_14_inv23 = 1;
    51: op1_14_inv23 = 1;
    52: op1_14_inv23 = 1;
    54: op1_14_inv23 = 1;
    55: op1_14_inv23 = 1;
    56: op1_14_inv23 = 1;
    57: op1_14_inv23 = 1;
    59: op1_14_inv23 = 1;
    62: op1_14_inv23 = 1;
    63: op1_14_inv23 = 1;
    64: op1_14_inv23 = 1;
    68: op1_14_inv23 = 1;
    69: op1_14_inv23 = 1;
    71: op1_14_inv23 = 1;
    76: op1_14_inv23 = 1;
    78: op1_14_inv23 = 1;
    79: op1_14_inv23 = 1;
    80: op1_14_inv23 = 1;
    82: op1_14_inv23 = 1;
    84: op1_14_inv23 = 1;
    85: op1_14_inv23 = 1;
    87: op1_14_inv23 = 1;
    88: op1_14_inv23 = 1;
    89: op1_14_inv23 = 1;
    90: op1_14_inv23 = 1;
    default: op1_14_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in24 = reg_0219;
    5: op1_14_in24 = imem07_in[3:0];
    6: op1_14_in24 = reg_0051;
    7: op1_14_in24 = reg_0282;
    8: op1_14_in24 = reg_0467;
    9: op1_14_in24 = imem07_in[71:68];
    36: op1_14_in24 = imem07_in[71:68];
    10: op1_14_in24 = reg_0009;
    11: op1_14_in24 = reg_0787;
    12: op1_14_in24 = imem03_in[115:112];
    13: op1_14_in24 = reg_0058;
    14: op1_14_in24 = reg_0617;
    15: op1_14_in24 = imem01_in[91:88];
    16: op1_14_in24 = reg_0579;
    17: op1_14_in24 = reg_0102;
    18: op1_14_in24 = reg_0087;
    19: op1_14_in24 = reg_0199;
    20: op1_14_in24 = reg_0557;
    21: op1_14_in24 = reg_0604;
    90: op1_14_in24 = reg_0604;
    22: op1_14_in24 = reg_0120;
    23: op1_14_in24 = reg_0443;
    24: op1_14_in24 = reg_0517;
    25: op1_14_in24 = reg_0277;
    26: op1_14_in24 = reg_0636;
    27: op1_14_in24 = imem03_in[75:72];
    28: op1_14_in24 = reg_0752;
    29: op1_14_in24 = reg_0507;
    30: op1_14_in24 = reg_0265;
    31: op1_14_in24 = reg_0276;
    32: op1_14_in24 = reg_0405;
    33: op1_14_in24 = reg_0374;
    34: op1_14_in24 = reg_0542;
    35: op1_14_in24 = reg_0267;
    37: op1_14_in24 = reg_0371;
    40: op1_14_in24 = imem01_in[115:112];
    41: op1_14_in24 = imem05_in[47:44];
    42: op1_14_in24 = reg_0701;
    44: op1_14_in24 = reg_0539;
    45: op1_14_in24 = reg_0138;
    47: op1_14_in24 = reg_0756;
    81: op1_14_in24 = reg_0756;
    48: op1_14_in24 = reg_0091;
    49: op1_14_in24 = reg_0354;
    50: op1_14_in24 = imem01_in[95:92];
    51: op1_14_in24 = reg_0448;
    52: op1_14_in24 = reg_0423;
    53: op1_14_in24 = imem01_in[19:16];
    54: op1_14_in24 = imem03_in[35:32];
    55: op1_14_in24 = reg_0052;
    56: op1_14_in24 = reg_0529;
    57: op1_14_in24 = imem03_in[31:28];
    58: op1_14_in24 = reg_0613;
    59: op1_14_in24 = reg_0560;
    60: op1_14_in24 = reg_0289;
    62: op1_14_in24 = reg_0533;
    63: op1_14_in24 = reg_0535;
    64: op1_14_in24 = imem03_in[67:64];
    77: op1_14_in24 = imem03_in[67:64];
    65: op1_14_in24 = reg_0315;
    66: op1_14_in24 = reg_0755;
    89: op1_14_in24 = reg_0755;
    67: op1_14_in24 = reg_0172;
    68: op1_14_in24 = reg_0422;
    86: op1_14_in24 = reg_0422;
    69: op1_14_in24 = reg_0303;
    71: op1_14_in24 = reg_0602;
    72: op1_14_in24 = imem04_in[83:80];
    73: op1_14_in24 = reg_0133;
    74: op1_14_in24 = imem06_in[83:80];
    75: op1_14_in24 = reg_0721;
    76: op1_14_in24 = reg_0111;
    78: op1_14_in24 = reg_0597;
    79: op1_14_in24 = reg_0793;
    80: op1_14_in24 = reg_0719;
    82: op1_14_in24 = imem01_in[51:48];
    84: op1_14_in24 = reg_0622;
    85: op1_14_in24 = imem04_in[75:72];
    87: op1_14_in24 = reg_0585;
    88: op1_14_in24 = reg_0660;
    91: op1_14_in24 = reg_0437;
    94: op1_14_in24 = reg_0724;
    95: op1_14_in24 = reg_0710;
    default: op1_14_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_14_inv24 = 1;
    6: op1_14_inv24 = 1;
    9: op1_14_inv24 = 1;
    11: op1_14_inv24 = 1;
    12: op1_14_inv24 = 1;
    15: op1_14_inv24 = 1;
    17: op1_14_inv24 = 1;
    18: op1_14_inv24 = 1;
    21: op1_14_inv24 = 1;
    23: op1_14_inv24 = 1;
    24: op1_14_inv24 = 1;
    28: op1_14_inv24 = 1;
    29: op1_14_inv24 = 1;
    30: op1_14_inv24 = 1;
    32: op1_14_inv24 = 1;
    33: op1_14_inv24 = 1;
    34: op1_14_inv24 = 1;
    35: op1_14_inv24 = 1;
    37: op1_14_inv24 = 1;
    40: op1_14_inv24 = 1;
    42: op1_14_inv24 = 1;
    45: op1_14_inv24 = 1;
    48: op1_14_inv24 = 1;
    49: op1_14_inv24 = 1;
    50: op1_14_inv24 = 1;
    57: op1_14_inv24 = 1;
    58: op1_14_inv24 = 1;
    59: op1_14_inv24 = 1;
    63: op1_14_inv24 = 1;
    65: op1_14_inv24 = 1;
    72: op1_14_inv24 = 1;
    73: op1_14_inv24 = 1;
    74: op1_14_inv24 = 1;
    75: op1_14_inv24 = 1;
    77: op1_14_inv24 = 1;
    78: op1_14_inv24 = 1;
    80: op1_14_inv24 = 1;
    82: op1_14_inv24 = 1;
    85: op1_14_inv24 = 1;
    86: op1_14_inv24 = 1;
    88: op1_14_inv24 = 1;
    90: op1_14_inv24 = 1;
    91: op1_14_inv24 = 1;
    94: op1_14_inv24 = 1;
    95: op1_14_inv24 = 1;
    default: op1_14_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in25 = reg_0122;
    5: op1_14_in25 = imem07_in[23:20];
    6: op1_14_in25 = reg_0060;
    7: op1_14_in25 = reg_0306;
    8: op1_14_in25 = reg_0471;
    9: op1_14_in25 = imem07_in[95:92];
    10: op1_14_in25 = reg_0010;
    11: op1_14_in25 = imem05_in[15:12];
    12: op1_14_in25 = reg_0583;
    16: op1_14_in25 = reg_0583;
    13: op1_14_in25 = reg_0057;
    14: op1_14_in25 = reg_0612;
    15: op1_14_in25 = imem01_in[103:100];
    17: op1_14_in25 = reg_0101;
    18: op1_14_in25 = reg_0093;
    19: op1_14_in25 = imem01_in[3:0];
    20: op1_14_in25 = reg_0553;
    65: op1_14_in25 = reg_0553;
    21: op1_14_in25 = reg_0630;
    22: op1_14_in25 = reg_0113;
    23: op1_14_in25 = reg_0448;
    24: op1_14_in25 = reg_0778;
    25: op1_14_in25 = reg_0143;
    26: op1_14_in25 = reg_0663;
    27: op1_14_in25 = imem03_in[79:76];
    54: op1_14_in25 = imem03_in[79:76];
    28: op1_14_in25 = imem07_in[7:4];
    29: op1_14_in25 = reg_0760;
    30: op1_14_in25 = reg_0278;
    31: op1_14_in25 = reg_0086;
    32: op1_14_in25 = reg_0773;
    33: op1_14_in25 = reg_0013;
    34: op1_14_in25 = reg_0055;
    35: op1_14_in25 = reg_0050;
    36: op1_14_in25 = imem07_in[79:76];
    37: op1_14_in25 = reg_0606;
    40: op1_14_in25 = reg_0112;
    41: op1_14_in25 = imem05_in[67:64];
    42: op1_14_in25 = reg_0727;
    44: op1_14_in25 = reg_0526;
    45: op1_14_in25 = imem06_in[7:4];
    47: op1_14_in25 = imem03_in[35:32];
    48: op1_14_in25 = reg_0545;
    49: op1_14_in25 = reg_0341;
    50: op1_14_in25 = imem01_in[127:124];
    51: op1_14_in25 = reg_0435;
    52: op1_14_in25 = reg_0511;
    53: op1_14_in25 = imem01_in[55:52];
    55: op1_14_in25 = reg_0302;
    56: op1_14_in25 = reg_0292;
    57: op1_14_in25 = imem03_in[43:40];
    58: op1_14_in25 = reg_0377;
    59: op1_14_in25 = reg_0087;
    60: op1_14_in25 = reg_0260;
    62: op1_14_in25 = reg_0540;
    63: op1_14_in25 = imem03_in[3:0];
    64: op1_14_in25 = imem03_in[75:72];
    66: op1_14_in25 = reg_0568;
    67: op1_14_in25 = reg_0179;
    68: op1_14_in25 = reg_0217;
    69: op1_14_in25 = reg_0283;
    71: op1_14_in25 = reg_0597;
    72: op1_14_in25 = imem04_in[91:88];
    73: op1_14_in25 = reg_0641;
    74: op1_14_in25 = imem06_in[99:96];
    75: op1_14_in25 = reg_0725;
    76: op1_14_in25 = reg_0520;
    77: op1_14_in25 = reg_0579;
    78: op1_14_in25 = reg_0319;
    79: op1_14_in25 = reg_0276;
    80: op1_14_in25 = reg_0285;
    81: op1_14_in25 = imem03_in[7:4];
    82: op1_14_in25 = imem01_in[87:84];
    84: op1_14_in25 = reg_0416;
    85: op1_14_in25 = reg_0247;
    86: op1_14_in25 = reg_0244;
    87: op1_14_in25 = reg_0513;
    88: op1_14_in25 = reg_0669;
    89: op1_14_in25 = reg_0637;
    90: op1_14_in25 = reg_0591;
    91: op1_14_in25 = reg_0116;
    94: op1_14_in25 = reg_0334;
    95: op1_14_in25 = reg_0715;
    default: op1_14_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv25 = 1;
    8: op1_14_inv25 = 1;
    10: op1_14_inv25 = 1;
    11: op1_14_inv25 = 1;
    18: op1_14_inv25 = 1;
    21: op1_14_inv25 = 1;
    22: op1_14_inv25 = 1;
    23: op1_14_inv25 = 1;
    24: op1_14_inv25 = 1;
    25: op1_14_inv25 = 1;
    26: op1_14_inv25 = 1;
    27: op1_14_inv25 = 1;
    29: op1_14_inv25 = 1;
    35: op1_14_inv25 = 1;
    36: op1_14_inv25 = 1;
    40: op1_14_inv25 = 1;
    41: op1_14_inv25 = 1;
    45: op1_14_inv25 = 1;
    47: op1_14_inv25 = 1;
    48: op1_14_inv25 = 1;
    49: op1_14_inv25 = 1;
    50: op1_14_inv25 = 1;
    52: op1_14_inv25 = 1;
    60: op1_14_inv25 = 1;
    64: op1_14_inv25 = 1;
    65: op1_14_inv25 = 1;
    66: op1_14_inv25 = 1;
    68: op1_14_inv25 = 1;
    73: op1_14_inv25 = 1;
    78: op1_14_inv25 = 1;
    79: op1_14_inv25 = 1;
    80: op1_14_inv25 = 1;
    84: op1_14_inv25 = 1;
    89: op1_14_inv25 = 1;
    90: op1_14_inv25 = 1;
    94: op1_14_inv25 = 1;
    default: op1_14_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in26 = reg_0111;
    5: op1_14_in26 = imem07_in[39:36];
    6: op1_14_in26 = reg_0087;
    7: op1_14_in26 = reg_0293;
    8: op1_14_in26 = reg_0478;
    9: op1_14_in26 = reg_0721;
    10: op1_14_in26 = imem04_in[7:4];
    11: op1_14_in26 = imem05_in[31:28];
    84: op1_14_in26 = imem05_in[31:28];
    12: op1_14_in26 = reg_0587;
    13: op1_14_in26 = imem05_in[3:0];
    14: op1_14_in26 = reg_0348;
    15: op1_14_in26 = imem01_in[111:108];
    16: op1_14_in26 = reg_0563;
    17: op1_14_in26 = imem02_in[23:20];
    18: op1_14_in26 = imem03_in[11:8];
    19: op1_14_in26 = imem01_in[19:16];
    20: op1_14_in26 = reg_0550;
    73: op1_14_in26 = reg_0550;
    21: op1_14_in26 = reg_0611;
    22: op1_14_in26 = imem02_in[11:8];
    23: op1_14_in26 = reg_0175;
    24: op1_14_in26 = reg_0324;
    25: op1_14_in26 = reg_0138;
    26: op1_14_in26 = reg_0344;
    27: op1_14_in26 = imem03_in[119:116];
    28: op1_14_in26 = imem07_in[11:8];
    29: op1_14_in26 = reg_0232;
    37: op1_14_in26 = reg_0232;
    30: op1_14_in26 = reg_0281;
    31: op1_14_in26 = reg_0148;
    32: op1_14_in26 = reg_0329;
    33: op1_14_in26 = reg_0802;
    34: op1_14_in26 = reg_0555;
    35: op1_14_in26 = reg_0284;
    36: op1_14_in26 = imem07_in[83:80];
    40: op1_14_in26 = reg_0115;
    41: op1_14_in26 = reg_0492;
    42: op1_14_in26 = imem07_in[15:12];
    44: op1_14_in26 = imem03_in[67:64];
    45: op1_14_in26 = imem06_in[19:16];
    47: op1_14_in26 = imem03_in[71:68];
    48: op1_14_in26 = reg_0328;
    65: op1_14_in26 = reg_0328;
    49: op1_14_in26 = reg_0356;
    50: op1_14_in26 = reg_0735;
    52: op1_14_in26 = reg_0574;
    53: op1_14_in26 = imem01_in[67:64];
    54: op1_14_in26 = imem03_in[103:100];
    55: op1_14_in26 = reg_0071;
    56: op1_14_in26 = reg_0431;
    57: op1_14_in26 = imem03_in[59:56];
    58: op1_14_in26 = reg_0763;
    59: op1_14_in26 = reg_0083;
    60: op1_14_in26 = reg_0242;
    62: op1_14_in26 = reg_0531;
    63: op1_14_in26 = imem03_in[99:96];
    64: op1_14_in26 = imem03_in[115:112];
    66: op1_14_in26 = reg_0562;
    67: op1_14_in26 = reg_0183;
    68: op1_14_in26 = reg_0424;
    69: op1_14_in26 = reg_0076;
    71: op1_14_in26 = reg_0604;
    72: op1_14_in26 = imem04_in[95:92];
    74: op1_14_in26 = imem06_in[103:100];
    75: op1_14_in26 = reg_0132;
    76: op1_14_in26 = reg_0741;
    77: op1_14_in26 = reg_0750;
    78: op1_14_in26 = reg_0591;
    79: op1_14_in26 = reg_0781;
    80: op1_14_in26 = reg_0058;
    81: op1_14_in26 = imem03_in[51:48];
    82: op1_14_in26 = imem01_in[91:88];
    85: op1_14_in26 = reg_0275;
    86: op1_14_in26 = reg_0220;
    87: op1_14_in26 = reg_0640;
    88: op1_14_in26 = reg_0674;
    89: op1_14_in26 = reg_0557;
    90: op1_14_in26 = reg_0318;
    91: op1_14_in26 = reg_0181;
    94: op1_14_in26 = reg_0434;
    95: op1_14_in26 = reg_0441;
    default: op1_14_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv26 = 1;
    5: op1_14_inv26 = 1;
    7: op1_14_inv26 = 1;
    9: op1_14_inv26 = 1;
    10: op1_14_inv26 = 1;
    11: op1_14_inv26 = 1;
    12: op1_14_inv26 = 1;
    16: op1_14_inv26 = 1;
    17: op1_14_inv26 = 1;
    18: op1_14_inv26 = 1;
    19: op1_14_inv26 = 1;
    20: op1_14_inv26 = 1;
    22: op1_14_inv26 = 1;
    23: op1_14_inv26 = 1;
    24: op1_14_inv26 = 1;
    25: op1_14_inv26 = 1;
    26: op1_14_inv26 = 1;
    28: op1_14_inv26 = 1;
    29: op1_14_inv26 = 1;
    30: op1_14_inv26 = 1;
    31: op1_14_inv26 = 1;
    32: op1_14_inv26 = 1;
    36: op1_14_inv26 = 1;
    40: op1_14_inv26 = 1;
    45: op1_14_inv26 = 1;
    48: op1_14_inv26 = 1;
    49: op1_14_inv26 = 1;
    53: op1_14_inv26 = 1;
    55: op1_14_inv26 = 1;
    57: op1_14_inv26 = 1;
    59: op1_14_inv26 = 1;
    64: op1_14_inv26 = 1;
    67: op1_14_inv26 = 1;
    68: op1_14_inv26 = 1;
    69: op1_14_inv26 = 1;
    72: op1_14_inv26 = 1;
    73: op1_14_inv26 = 1;
    74: op1_14_inv26 = 1;
    76: op1_14_inv26 = 1;
    77: op1_14_inv26 = 1;
    80: op1_14_inv26 = 1;
    81: op1_14_inv26 = 1;
    84: op1_14_inv26 = 1;
    87: op1_14_inv26 = 1;
    88: op1_14_inv26 = 1;
    89: op1_14_inv26 = 1;
    91: op1_14_inv26 = 1;
    95: op1_14_inv26 = 1;
    default: op1_14_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in27 = reg_0112;
    5: op1_14_in27 = imem07_in[63:60];
    6: op1_14_in27 = imem03_in[23:20];
    7: op1_14_in27 = reg_0296;
    56: op1_14_in27 = reg_0296;
    8: op1_14_in27 = reg_0200;
    9: op1_14_in27 = reg_0715;
    10: op1_14_in27 = imem04_in[99:96];
    72: op1_14_in27 = imem04_in[99:96];
    11: op1_14_in27 = imem05_in[47:44];
    12: op1_14_in27 = reg_0360;
    13: op1_14_in27 = imem05_in[43:40];
    84: op1_14_in27 = imem05_in[43:40];
    14: op1_14_in27 = reg_0332;
    15: op1_14_in27 = imem01_in[119:116];
    16: op1_14_in27 = reg_0585;
    17: op1_14_in27 = imem02_in[67:64];
    18: op1_14_in27 = imem03_in[27:24];
    19: op1_14_in27 = imem01_in[27:24];
    20: op1_14_in27 = reg_0549;
    21: op1_14_in27 = reg_0622;
    22: op1_14_in27 = imem02_in[19:16];
    88: op1_14_in27 = imem02_in[19:16];
    23: op1_14_in27 = reg_0180;
    24: op1_14_in27 = reg_0755;
    25: op1_14_in27 = reg_0129;
    26: op1_14_in27 = reg_0357;
    27: op1_14_in27 = imem03_in[123:120];
    47: op1_14_in27 = imem03_in[123:120];
    28: op1_14_in27 = imem07_in[19:16];
    42: op1_14_in27 = imem07_in[19:16];
    29: op1_14_in27 = reg_0511;
    30: op1_14_in27 = reg_0076;
    31: op1_14_in27 = reg_0145;
    32: op1_14_in27 = reg_0038;
    33: op1_14_in27 = reg_0016;
    34: op1_14_in27 = reg_0060;
    35: op1_14_in27 = reg_0281;
    36: op1_14_in27 = imem07_in[103:100];
    37: op1_14_in27 = reg_0774;
    40: op1_14_in27 = imem02_in[71:68];
    41: op1_14_in27 = reg_0493;
    44: op1_14_in27 = imem03_in[103:100];
    45: op1_14_in27 = imem06_in[47:44];
    48: op1_14_in27 = reg_0087;
    49: op1_14_in27 = reg_0518;
    50: op1_14_in27 = reg_0733;
    52: op1_14_in27 = reg_0294;
    53: op1_14_in27 = imem01_in[127:124];
    54: op1_14_in27 = imem03_in[115:112];
    55: op1_14_in27 = reg_0503;
    57: op1_14_in27 = imem03_in[71:68];
    58: op1_14_in27 = reg_0270;
    59: op1_14_in27 = reg_0556;
    60: op1_14_in27 = reg_0031;
    62: op1_14_in27 = reg_0098;
    63: op1_14_in27 = imem03_in[127:124];
    64: op1_14_in27 = reg_0602;
    65: op1_14_in27 = reg_0542;
    66: op1_14_in27 = reg_0396;
    67: op1_14_in27 = reg_0176;
    68: op1_14_in27 = reg_0243;
    69: op1_14_in27 = reg_0629;
    71: op1_14_in27 = reg_0596;
    73: op1_14_in27 = reg_0231;
    74: op1_14_in27 = imem06_in[115:112];
    75: op1_14_in27 = reg_0295;
    76: op1_14_in27 = reg_0645;
    77: op1_14_in27 = reg_0318;
    78: op1_14_in27 = reg_0318;
    79: op1_14_in27 = reg_0151;
    80: op1_14_in27 = reg_0148;
    81: op1_14_in27 = imem03_in[55:52];
    82: op1_14_in27 = imem01_in[95:92];
    85: op1_14_in27 = reg_0548;
    86: op1_14_in27 = reg_0425;
    87: op1_14_in27 = reg_0233;
    89: op1_14_in27 = reg_0649;
    90: op1_14_in27 = reg_0572;
    91: op1_14_in27 = reg_0730;
    94: op1_14_in27 = reg_0268;
    95: op1_14_in27 = reg_0266;
    default: op1_14_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv27 = 1;
    5: op1_14_inv27 = 1;
    6: op1_14_inv27 = 1;
    8: op1_14_inv27 = 1;
    10: op1_14_inv27 = 1;
    11: op1_14_inv27 = 1;
    13: op1_14_inv27 = 1;
    15: op1_14_inv27 = 1;
    16: op1_14_inv27 = 1;
    18: op1_14_inv27 = 1;
    20: op1_14_inv27 = 1;
    21: op1_14_inv27 = 1;
    22: op1_14_inv27 = 1;
    23: op1_14_inv27 = 1;
    27: op1_14_inv27 = 1;
    28: op1_14_inv27 = 1;
    30: op1_14_inv27 = 1;
    31: op1_14_inv27 = 1;
    32: op1_14_inv27 = 1;
    33: op1_14_inv27 = 1;
    36: op1_14_inv27 = 1;
    42: op1_14_inv27 = 1;
    44: op1_14_inv27 = 1;
    49: op1_14_inv27 = 1;
    52: op1_14_inv27 = 1;
    54: op1_14_inv27 = 1;
    56: op1_14_inv27 = 1;
    58: op1_14_inv27 = 1;
    59: op1_14_inv27 = 1;
    60: op1_14_inv27 = 1;
    63: op1_14_inv27 = 1;
    64: op1_14_inv27 = 1;
    66: op1_14_inv27 = 1;
    67: op1_14_inv27 = 1;
    68: op1_14_inv27 = 1;
    69: op1_14_inv27 = 1;
    71: op1_14_inv27 = 1;
    72: op1_14_inv27 = 1;
    76: op1_14_inv27 = 1;
    77: op1_14_inv27 = 1;
    81: op1_14_inv27 = 1;
    82: op1_14_inv27 = 1;
    84: op1_14_inv27 = 1;
    85: op1_14_inv27 = 1;
    89: op1_14_inv27 = 1;
    90: op1_14_inv27 = 1;
    91: op1_14_inv27 = 1;
    95: op1_14_inv27 = 1;
    default: op1_14_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in28 = reg_0113;
    5: op1_14_in28 = imem07_in[79:76];
    6: op1_14_in28 = imem03_in[35:32];
    7: op1_14_in28 = reg_0297;
    69: op1_14_in28 = reg_0297;
    8: op1_14_in28 = reg_0208;
    9: op1_14_in28 = reg_0701;
    10: op1_14_in28 = reg_0543;
    11: op1_14_in28 = imem05_in[59:56];
    12: op1_14_in28 = reg_0319;
    13: op1_14_in28 = imem05_in[119:116];
    14: op1_14_in28 = reg_0344;
    15: op1_14_in28 = reg_0821;
    24: op1_14_in28 = reg_0821;
    16: op1_14_in28 = reg_0578;
    17: op1_14_in28 = imem02_in[91:88];
    18: op1_14_in28 = imem03_in[63:60];
    19: op1_14_in28 = imem01_in[55:52];
    20: op1_14_in28 = reg_0554;
    21: op1_14_in28 = reg_0407;
    22: op1_14_in28 = imem02_in[23:20];
    23: op1_14_in28 = reg_0165;
    25: op1_14_in28 = imem06_in[15:12];
    26: op1_14_in28 = reg_0341;
    27: op1_14_in28 = reg_0006;
    28: op1_14_in28 = imem07_in[27:24];
    29: op1_14_in28 = reg_0506;
    30: op1_14_in28 = reg_0255;
    31: op1_14_in28 = reg_0135;
    32: op1_14_in28 = reg_0764;
    33: op1_14_in28 = reg_0009;
    34: op1_14_in28 = reg_0551;
    35: op1_14_in28 = reg_0065;
    36: op1_14_in28 = imem07_in[107:104];
    37: op1_14_in28 = reg_0317;
    40: op1_14_in28 = imem02_in[95:92];
    41: op1_14_in28 = reg_0489;
    42: op1_14_in28 = imem07_in[35:32];
    44: op1_14_in28 = reg_0582;
    45: op1_14_in28 = imem06_in[79:76];
    47: op1_14_in28 = reg_0259;
    48: op1_14_in28 = reg_0542;
    49: op1_14_in28 = reg_0092;
    50: op1_14_in28 = reg_0765;
    52: op1_14_in28 = reg_0248;
    53: op1_14_in28 = reg_0646;
    54: op1_14_in28 = reg_0573;
    55: op1_14_in28 = reg_0431;
    56: op1_14_in28 = reg_0640;
    57: op1_14_in28 = reg_0602;
    58: op1_14_in28 = reg_0753;
    59: op1_14_in28 = reg_0283;
    60: op1_14_in28 = reg_0583;
    62: op1_14_in28 = reg_0526;
    63: op1_14_in28 = reg_0347;
    64: op1_14_in28 = reg_0347;
    65: op1_14_in28 = reg_0537;
    66: op1_14_in28 = reg_0374;
    68: op1_14_in28 = reg_0505;
    71: op1_14_in28 = reg_0528;
    72: op1_14_in28 = imem04_in[119:116];
    73: op1_14_in28 = reg_0090;
    74: op1_14_in28 = reg_0354;
    75: op1_14_in28 = reg_0436;
    76: op1_14_in28 = reg_0112;
    77: op1_14_in28 = reg_0350;
    78: op1_14_in28 = reg_0600;
    79: op1_14_in28 = reg_0742;
    80: op1_14_in28 = reg_0149;
    81: op1_14_in28 = imem03_in[59:56];
    82: op1_14_in28 = imem01_in[99:96];
    84: op1_14_in28 = imem05_in[67:64];
    85: op1_14_in28 = reg_0516;
    86: op1_14_in28 = reg_0234;
    87: op1_14_in28 = imem05_in[7:4];
    88: op1_14_in28 = imem02_in[31:28];
    89: op1_14_in28 = imem03_in[23:20];
    90: op1_14_in28 = reg_0387;
    91: op1_14_in28 = reg_0184;
    94: op1_14_in28 = reg_0182;
    95: op1_14_in28 = reg_0333;
    default: op1_14_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv28 = 1;
    6: op1_14_inv28 = 1;
    7: op1_14_inv28 = 1;
    12: op1_14_inv28 = 1;
    13: op1_14_inv28 = 1;
    16: op1_14_inv28 = 1;
    19: op1_14_inv28 = 1;
    20: op1_14_inv28 = 1;
    21: op1_14_inv28 = 1;
    22: op1_14_inv28 = 1;
    23: op1_14_inv28 = 1;
    25: op1_14_inv28 = 1;
    28: op1_14_inv28 = 1;
    29: op1_14_inv28 = 1;
    32: op1_14_inv28 = 1;
    34: op1_14_inv28 = 1;
    40: op1_14_inv28 = 1;
    44: op1_14_inv28 = 1;
    50: op1_14_inv28 = 1;
    52: op1_14_inv28 = 1;
    53: op1_14_inv28 = 1;
    54: op1_14_inv28 = 1;
    55: op1_14_inv28 = 1;
    58: op1_14_inv28 = 1;
    59: op1_14_inv28 = 1;
    60: op1_14_inv28 = 1;
    63: op1_14_inv28 = 1;
    64: op1_14_inv28 = 1;
    65: op1_14_inv28 = 1;
    66: op1_14_inv28 = 1;
    69: op1_14_inv28 = 1;
    71: op1_14_inv28 = 1;
    73: op1_14_inv28 = 1;
    74: op1_14_inv28 = 1;
    75: op1_14_inv28 = 1;
    77: op1_14_inv28 = 1;
    80: op1_14_inv28 = 1;
    81: op1_14_inv28 = 1;
    85: op1_14_inv28 = 1;
    86: op1_14_inv28 = 1;
    87: op1_14_inv28 = 1;
    88: op1_14_inv28 = 1;
    91: op1_14_inv28 = 1;
    94: op1_14_inv28 = 1;
    default: op1_14_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in29 = reg_0121;
    5: op1_14_in29 = imem07_in[91:88];
    6: op1_14_in29 = imem03_in[47:44];
    7: op1_14_in29 = reg_0275;
    8: op1_14_in29 = reg_0191;
    9: op1_14_in29 = reg_0430;
    10: op1_14_in29 = reg_0552;
    11: op1_14_in29 = imem05_in[107:104];
    12: op1_14_in29 = reg_0385;
    13: op1_14_in29 = reg_0490;
    14: op1_14_in29 = reg_0372;
    15: op1_14_in29 = reg_0216;
    29: op1_14_in29 = reg_0216;
    16: op1_14_in29 = reg_0576;
    17: op1_14_in29 = imem02_in[99:96];
    18: op1_14_in29 = imem03_in[79:76];
    19: op1_14_in29 = imem01_in[59:56];
    20: op1_14_in29 = reg_0556;
    21: op1_14_in29 = reg_0409;
    22: op1_14_in29 = reg_0653;
    23: op1_14_in29 = reg_0162;
    24: op1_14_in29 = imem01_in[15:12];
    25: op1_14_in29 = imem06_in[83:80];
    26: op1_14_in29 = reg_0324;
    27: op1_14_in29 = reg_0811;
    28: op1_14_in29 = imem07_in[31:28];
    30: op1_14_in29 = reg_0068;
    31: op1_14_in29 = reg_0143;
    32: op1_14_in29 = reg_0814;
    33: op1_14_in29 = imem04_in[15:12];
    34: op1_14_in29 = reg_0547;
    35: op1_14_in29 = reg_0288;
    36: op1_14_in29 = imem07_in[115:112];
    37: op1_14_in29 = reg_0242;
    40: op1_14_in29 = reg_0640;
    41: op1_14_in29 = reg_0226;
    42: op1_14_in29 = imem07_in[47:44];
    44: op1_14_in29 = reg_0591;
    45: op1_14_in29 = imem06_in[115:112];
    47: op1_14_in29 = reg_0599;
    48: op1_14_in29 = reg_0055;
    49: op1_14_in29 = reg_0080;
    50: op1_14_in29 = reg_0649;
    52: op1_14_in29 = reg_0243;
    53: op1_14_in29 = reg_0733;
    54: op1_14_in29 = reg_0561;
    55: op1_14_in29 = reg_0508;
    56: op1_14_in29 = imem05_in[35:32];
    57: op1_14_in29 = reg_0347;
    58: op1_14_in29 = reg_0620;
    59: op1_14_in29 = reg_0503;
    60: op1_14_in29 = reg_0593;
    62: op1_14_in29 = reg_0538;
    63: op1_14_in29 = reg_0582;
    64: op1_14_in29 = reg_0604;
    65: op1_14_in29 = reg_0056;
    66: op1_14_in29 = reg_0570;
    68: op1_14_in29 = reg_0677;
    69: op1_14_in29 = reg_0292;
    71: op1_14_in29 = reg_0395;
    72: op1_14_in29 = reg_0059;
    73: op1_14_in29 = reg_0517;
    74: op1_14_in29 = reg_0408;
    75: op1_14_in29 = reg_0635;
    76: op1_14_in29 = reg_0778;
    77: op1_14_in29 = reg_0399;
    78: op1_14_in29 = reg_0488;
    79: op1_14_in29 = reg_0153;
    80: op1_14_in29 = reg_0742;
    81: op1_14_in29 = imem03_in[75:72];
    82: op1_14_in29 = reg_0497;
    84: op1_14_in29 = imem05_in[79:76];
    85: op1_14_in29 = reg_0174;
    86: op1_14_in29 = reg_0506;
    87: op1_14_in29 = imem05_in[55:52];
    88: op1_14_in29 = imem02_in[43:40];
    89: op1_14_in29 = imem03_in[31:28];
    90: op1_14_in29 = reg_0623;
    94: op1_14_in29 = reg_0325;
    95: op1_14_in29 = reg_0239;
    default: op1_14_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_14_inv29 = 1;
    7: op1_14_inv29 = 1;
    8: op1_14_inv29 = 1;
    13: op1_14_inv29 = 1;
    16: op1_14_inv29 = 1;
    17: op1_14_inv29 = 1;
    18: op1_14_inv29 = 1;
    22: op1_14_inv29 = 1;
    26: op1_14_inv29 = 1;
    28: op1_14_inv29 = 1;
    30: op1_14_inv29 = 1;
    32: op1_14_inv29 = 1;
    41: op1_14_inv29 = 1;
    45: op1_14_inv29 = 1;
    49: op1_14_inv29 = 1;
    50: op1_14_inv29 = 1;
    52: op1_14_inv29 = 1;
    53: op1_14_inv29 = 1;
    55: op1_14_inv29 = 1;
    57: op1_14_inv29 = 1;
    59: op1_14_inv29 = 1;
    60: op1_14_inv29 = 1;
    65: op1_14_inv29 = 1;
    68: op1_14_inv29 = 1;
    71: op1_14_inv29 = 1;
    72: op1_14_inv29 = 1;
    73: op1_14_inv29 = 1;
    74: op1_14_inv29 = 1;
    75: op1_14_inv29 = 1;
    76: op1_14_inv29 = 1;
    77: op1_14_inv29 = 1;
    78: op1_14_inv29 = 1;
    79: op1_14_inv29 = 1;
    80: op1_14_inv29 = 1;
    84: op1_14_inv29 = 1;
    85: op1_14_inv29 = 1;
    86: op1_14_inv29 = 1;
    88: op1_14_inv29 = 1;
    89: op1_14_inv29 = 1;
    default: op1_14_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_14_in30 = imem02_in[23:20];
    5: op1_14_in30 = imem07_in[107:104];
    6: op1_14_in30 = imem03_in[51:48];
    7: op1_14_in30 = reg_0278;
    8: op1_14_in30 = reg_0187;
    9: op1_14_in30 = reg_0432;
    10: op1_14_in30 = reg_0548;
    11: op1_14_in30 = reg_0132;
    12: op1_14_in30 = reg_0398;
    13: op1_14_in30 = reg_0488;
    14: op1_14_in30 = reg_0408;
    15: op1_14_in30 = reg_0220;
    16: op1_14_in30 = reg_0319;
    17: op1_14_in30 = imem02_in[127:124];
    18: op1_14_in30 = imem03_in[99:96];
    19: op1_14_in30 = imem01_in[83:80];
    20: op1_14_in30 = reg_0547;
    21: op1_14_in30 = reg_0399;
    22: op1_14_in30 = reg_0661;
    23: op1_14_in30 = reg_0159;
    24: op1_14_in30 = imem01_in[19:16];
    25: op1_14_in30 = imem06_in[115:112];
    26: op1_14_in30 = reg_0322;
    27: op1_14_in30 = reg_0808;
    28: op1_14_in30 = imem07_in[47:44];
    29: op1_14_in30 = reg_0245;
    30: op1_14_in30 = imem05_in[11:8];
    35: op1_14_in30 = imem05_in[11:8];
    31: op1_14_in30 = reg_0153;
    32: op1_14_in30 = reg_0028;
    33: op1_14_in30 = imem04_in[27:24];
    34: op1_14_in30 = reg_0280;
    85: op1_14_in30 = reg_0280;
    36: op1_14_in30 = reg_0722;
    37: op1_14_in30 = reg_0375;
    40: op1_14_in30 = reg_0641;
    41: op1_14_in30 = reg_0282;
    42: op1_14_in30 = reg_0162;
    44: op1_14_in30 = reg_0593;
    45: op1_14_in30 = reg_0625;
    47: op1_14_in30 = reg_0583;
    48: op1_14_in30 = reg_0555;
    49: op1_14_in30 = reg_0097;
    50: op1_14_in30 = reg_0100;
    52: op1_14_in30 = imem01_in[15:12];
    53: op1_14_in30 = reg_0761;
    54: op1_14_in30 = reg_0811;
    55: op1_14_in30 = reg_0626;
    56: op1_14_in30 = imem05_in[39:36];
    57: op1_14_in30 = reg_0589;
    58: op1_14_in30 = reg_0040;
    59: op1_14_in30 = reg_0679;
    60: op1_14_in30 = reg_0576;
    62: op1_14_in30 = reg_0532;
    63: op1_14_in30 = reg_0493;
    64: op1_14_in30 = reg_0493;
    65: op1_14_in30 = reg_0060;
    66: op1_14_in30 = reg_0000;
    68: op1_14_in30 = reg_0674;
    69: op1_14_in30 = reg_0050;
    71: op1_14_in30 = reg_0496;
    72: op1_14_in30 = reg_0537;
    73: op1_14_in30 = reg_0075;
    74: op1_14_in30 = reg_0377;
    75: op1_14_in30 = reg_0239;
    76: op1_14_in30 = reg_0507;
    77: op1_14_in30 = reg_0357;
    78: op1_14_in30 = reg_0648;
    79: op1_14_in30 = reg_0137;
    80: op1_14_in30 = imem06_in[27:24];
    81: op1_14_in30 = imem03_in[79:76];
    82: op1_14_in30 = reg_0520;
    84: op1_14_in30 = imem05_in[83:80];
    86: op1_14_in30 = reg_0419;
    87: op1_14_in30 = imem05_in[99:96];
    88: op1_14_in30 = imem02_in[47:44];
    89: op1_14_in30 = imem03_in[87:84];
    90: op1_14_in30 = reg_0800;
    94: op1_14_in30 = reg_0176;
    95: op1_14_in30 = reg_0444;
    default: op1_14_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_14_inv30 = 1;
    6: op1_14_inv30 = 1;
    7: op1_14_inv30 = 1;
    8: op1_14_inv30 = 1;
    9: op1_14_inv30 = 1;
    10: op1_14_inv30 = 1;
    11: op1_14_inv30 = 1;
    15: op1_14_inv30 = 1;
    18: op1_14_inv30 = 1;
    19: op1_14_inv30 = 1;
    21: op1_14_inv30 = 1;
    23: op1_14_inv30 = 1;
    27: op1_14_inv30 = 1;
    28: op1_14_inv30 = 1;
    36: op1_14_inv30 = 1;
    37: op1_14_inv30 = 1;
    41: op1_14_inv30 = 1;
    44: op1_14_inv30 = 1;
    48: op1_14_inv30 = 1;
    52: op1_14_inv30 = 1;
    54: op1_14_inv30 = 1;
    56: op1_14_inv30 = 1;
    58: op1_14_inv30 = 1;
    62: op1_14_inv30 = 1;
    64: op1_14_inv30 = 1;
    66: op1_14_inv30 = 1;
    69: op1_14_inv30 = 1;
    71: op1_14_inv30 = 1;
    74: op1_14_inv30 = 1;
    76: op1_14_inv30 = 1;
    77: op1_14_inv30 = 1;
    78: op1_14_inv30 = 1;
    81: op1_14_inv30 = 1;
    82: op1_14_inv30 = 1;
    84: op1_14_inv30 = 1;
    85: op1_14_inv30 = 1;
    88: op1_14_inv30 = 1;
    89: op1_14_inv30 = 1;
    90: op1_14_inv30 = 1;
    94: op1_14_inv30 = 1;
    95: op1_14_inv30 = 1;
    default: op1_14_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_14_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_14_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の0番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in00 = imem02_in[31:28];
    5: op1_15_in00 = imem07_in[123:120];
    6: op1_15_in00 = imem03_in[75:72];
    7: op1_15_in00 = reg_0046;
    8: op1_15_in00 = reg_0188;
    90: op1_15_in00 = reg_0188;
    9: op1_15_in00 = imem00_in[35:32];
    51: op1_15_in00 = imem00_in[35:32];
    10: op1_15_in00 = reg_0541;
    11: op1_15_in00 = reg_0148;
    12: op1_15_in00 = reg_0389;
    13: op1_15_in00 = reg_0736;
    87: op1_15_in00 = reg_0736;
    14: op1_15_in00 = reg_0403;
    15: op1_15_in00 = reg_0503;
    16: op1_15_in00 = reg_0327;
    17: op1_15_in00 = reg_0666;
    18: op1_15_in00 = reg_0578;
    19: op1_15_in00 = imem01_in[99:96];
    20: op1_15_in00 = reg_0052;
    21: op1_15_in00 = reg_0367;
    22: op1_15_in00 = reg_0640;
    23: op1_15_in00 = imem00_in[51:48];
    24: op1_15_in00 = imem01_in[39:36];
    25: op1_15_in00 = reg_0610;
    26: op1_15_in00 = reg_0321;
    27: op1_15_in00 = reg_0807;
    28: op1_15_in00 = imem07_in[119:116];
    3: op1_15_in00 = imem07_in[47:44];
    29: op1_15_in00 = reg_0123;
    30: op1_15_in00 = imem05_in[27:24];
    31: op1_15_in00 = reg_0130;
    32: op1_15_in00 = reg_0812;
    1: op1_15_in00 = imem07_in[99:96];
    33: op1_15_in00 = imem04_in[35:32];
    2: op1_15_in00 = reg_0170;
    34: op1_15_in00 = reg_0273;
    35: op1_15_in00 = imem05_in[23:20];
    36: op1_15_in00 = reg_0723;
    37: op1_15_in00 = reg_0037;
    38: op1_15_in00 = imem00_in[67:64];
    39: op1_15_in00 = imem00_in[23:20];
    91: op1_15_in00 = imem00_in[23:20];
    40: op1_15_in00 = reg_0665;
    41: op1_15_in00 = reg_0155;
    42: op1_15_in00 = reg_0169;
    43: op1_15_in00 = imem00_in[3:0];
    67: op1_15_in00 = imem00_in[3:0];
    92: op1_15_in00 = imem00_in[3:0];
    44: op1_15_in00 = reg_0597;
    45: op1_15_in00 = reg_0630;
    46: op1_15_in00 = imem00_in[7:4];
    61: op1_15_in00 = imem00_in[7:4];
    47: op1_15_in00 = reg_0565;
    48: op1_15_in00 = reg_0060;
    49: op1_15_in00 = reg_0540;
    50: op1_15_in00 = reg_0563;
    52: op1_15_in00 = imem01_in[55:52];
    53: op1_15_in00 = reg_0825;
    54: op1_15_in00 = reg_0003;
    55: op1_15_in00 = reg_0227;
    56: op1_15_in00 = imem05_in[71:68];
    57: op1_15_in00 = reg_0599;
    58: op1_15_in00 = reg_0621;
    59: op1_15_in00 = imem05_in[11:8];
    60: op1_15_in00 = imem06_in[27:24];
    62: op1_15_in00 = imem03_in[3:0];
    63: op1_15_in00 = reg_0750;
    64: op1_15_in00 = reg_0357;
    65: op1_15_in00 = reg_0516;
    66: op1_15_in00 = reg_0013;
    68: op1_15_in00 = reg_0121;
    69: op1_15_in00 = reg_0617;
    70: op1_15_in00 = imem00_in[43:40];
    71: op1_15_in00 = reg_0396;
    72: op1_15_in00 = reg_0523;
    73: op1_15_in00 = reg_0245;
    74: op1_15_in00 = reg_0405;
    75: op1_15_in00 = reg_0446;
    76: op1_15_in00 = reg_0232;
    77: op1_15_in00 = reg_0588;
    78: op1_15_in00 = reg_0384;
    79: op1_15_in00 = imem06_in[11:8];
    80: op1_15_in00 = imem06_in[47:44];
    81: op1_15_in00 = imem03_in[83:80];
    82: op1_15_in00 = reg_0224;
    83: op1_15_in00 = imem00_in[31:28];
    84: op1_15_in00 = imem05_in[127:124];
    85: op1_15_in00 = reg_0631;
    86: op1_15_in00 = reg_0420;
    88: op1_15_in00 = reg_0088;
    89: op1_15_in00 = imem03_in[111:108];
    93: op1_15_in00 = imem00_in[15:12];
    94: op1_15_in00 = reg_0140;
    95: op1_15_in00 = reg_0267;
    default: op1_15_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv00 = 1;
    7: op1_15_inv00 = 1;
    10: op1_15_inv00 = 1;
    16: op1_15_inv00 = 1;
    18: op1_15_inv00 = 1;
    20: op1_15_inv00 = 1;
    21: op1_15_inv00 = 1;
    23: op1_15_inv00 = 1;
    24: op1_15_inv00 = 1;
    25: op1_15_inv00 = 1;
    28: op1_15_inv00 = 1;
    3: op1_15_inv00 = 1;
    31: op1_15_inv00 = 1;
    1: op1_15_inv00 = 1;
    33: op1_15_inv00 = 1;
    35: op1_15_inv00 = 1;
    38: op1_15_inv00 = 1;
    40: op1_15_inv00 = 1;
    43: op1_15_inv00 = 1;
    44: op1_15_inv00 = 1;
    45: op1_15_inv00 = 1;
    46: op1_15_inv00 = 1;
    47: op1_15_inv00 = 1;
    48: op1_15_inv00 = 1;
    50: op1_15_inv00 = 1;
    52: op1_15_inv00 = 1;
    53: op1_15_inv00 = 1;
    54: op1_15_inv00 = 1;
    56: op1_15_inv00 = 1;
    57: op1_15_inv00 = 1;
    58: op1_15_inv00 = 1;
    60: op1_15_inv00 = 1;
    62: op1_15_inv00 = 1;
    65: op1_15_inv00 = 1;
    67: op1_15_inv00 = 1;
    69: op1_15_inv00 = 1;
    70: op1_15_inv00 = 1;
    72: op1_15_inv00 = 1;
    74: op1_15_inv00 = 1;
    77: op1_15_inv00 = 1;
    78: op1_15_inv00 = 1;
    79: op1_15_inv00 = 1;
    80: op1_15_inv00 = 1;
    82: op1_15_inv00 = 1;
    83: op1_15_inv00 = 1;
    84: op1_15_inv00 = 1;
    85: op1_15_inv00 = 1;
    86: op1_15_inv00 = 1;
    87: op1_15_inv00 = 1;
    90: op1_15_inv00 = 1;
    91: op1_15_inv00 = 1;
    93: op1_15_inv00 = 1;
    94: op1_15_inv00 = 1;
    default: op1_15_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の1番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in01 = imem02_in[43:40];
    5: op1_15_in01 = reg_0704;
    6: op1_15_in01 = imem03_in[87:84];
    7: op1_15_in01 = imem05_in[3:0];
    8: op1_15_in01 = reg_0203;
    9: op1_15_in01 = imem00_in[47:44];
    51: op1_15_in01 = imem00_in[47:44];
    10: op1_15_in01 = reg_0547;
    11: op1_15_in01 = reg_0136;
    12: op1_15_in01 = reg_0019;
    13: op1_15_in01 = reg_0737;
    14: op1_15_in01 = reg_0390;
    15: op1_15_in01 = reg_0243;
    16: op1_15_in01 = reg_0377;
    17: op1_15_in01 = reg_0664;
    18: op1_15_in01 = reg_0581;
    19: op1_15_in01 = imem01_in[127:124];
    20: op1_15_in01 = reg_0534;
    21: op1_15_in01 = reg_0401;
    22: op1_15_in01 = reg_0667;
    23: op1_15_in01 = imem00_in[83:80];
    24: op1_15_in01 = imem01_in[59:56];
    25: op1_15_in01 = reg_0625;
    26: op1_15_in01 = reg_0323;
    27: op1_15_in01 = imem04_in[31:28];
    28: op1_15_in01 = reg_0720;
    3: op1_15_in01 = imem07_in[51:48];
    29: op1_15_in01 = reg_0105;
    30: op1_15_in01 = imem05_in[67:64];
    31: op1_15_in01 = reg_0131;
    32: op1_15_in01 = reg_0338;
    33: op1_15_in01 = imem04_in[39:36];
    34: op1_15_in01 = reg_0267;
    35: op1_15_in01 = imem05_in[43:40];
    36: op1_15_in01 = reg_0703;
    37: op1_15_in01 = reg_0238;
    38: op1_15_in01 = imem00_in[71:68];
    39: op1_15_in01 = imem00_in[67:64];
    40: op1_15_in01 = reg_0352;
    41: op1_15_in01 = imem06_in[15:12];
    42: op1_15_in01 = reg_0163;
    43: op1_15_in01 = imem00_in[15:12];
    44: op1_15_in01 = reg_0384;
    45: op1_15_in01 = reg_0624;
    46: op1_15_in01 = imem00_in[23:20];
    47: op1_15_in01 = reg_0039;
    48: op1_15_in01 = reg_0516;
    49: op1_15_in01 = reg_0535;
    50: op1_15_in01 = reg_0825;
    52: op1_15_in01 = imem01_in[75:72];
    53: op1_15_in01 = reg_0232;
    54: op1_15_in01 = reg_0807;
    55: op1_15_in01 = reg_0519;
    56: op1_15_in01 = imem05_in[127:124];
    57: op1_15_in01 = reg_0319;
    58: op1_15_in01 = reg_0231;
    59: op1_15_in01 = imem05_in[31:28];
    60: op1_15_in01 = imem06_in[115:112];
    61: op1_15_in01 = imem00_in[51:48];
    70: op1_15_in01 = imem00_in[51:48];
    83: op1_15_in01 = imem00_in[51:48];
    91: op1_15_in01 = imem00_in[51:48];
    62: op1_15_in01 = imem03_in[11:8];
    63: op1_15_in01 = reg_0329;
    64: op1_15_in01 = reg_0331;
    65: op1_15_in01 = reg_0556;
    66: op1_15_in01 = reg_0007;
    67: op1_15_in01 = imem00_in[7:4];
    68: op1_15_in01 = imem02_in[35:32];
    69: op1_15_in01 = reg_0626;
    71: op1_15_in01 = reg_0811;
    72: op1_15_in01 = reg_0551;
    73: op1_15_in01 = reg_0276;
    74: op1_15_in01 = reg_0583;
    75: op1_15_in01 = reg_0442;
    76: op1_15_in01 = reg_0511;
    77: op1_15_in01 = reg_0751;
    78: op1_15_in01 = reg_0417;
    79: op1_15_in01 = imem06_in[35:32];
    80: op1_15_in01 = imem06_in[103:100];
    81: op1_15_in01 = imem03_in[107:104];
    82: op1_15_in01 = reg_0388;
    84: op1_15_in01 = reg_0791;
    85: op1_15_in01 = reg_0074;
    86: op1_15_in01 = reg_0124;
    87: op1_15_in01 = reg_0227;
    88: op1_15_in01 = reg_0530;
    89: op1_15_in01 = imem03_in[115:112];
    90: op1_15_in01 = imem04_in[47:44];
    92: op1_15_in01 = imem00_in[11:8];
    93: op1_15_in01 = imem00_in[63:60];
    95: op1_15_in01 = reg_0438;
    default: op1_15_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv01 = 1;
    8: op1_15_inv01 = 1;
    9: op1_15_inv01 = 1;
    10: op1_15_inv01 = 1;
    11: op1_15_inv01 = 1;
    12: op1_15_inv01 = 1;
    18: op1_15_inv01 = 1;
    19: op1_15_inv01 = 1;
    21: op1_15_inv01 = 1;
    22: op1_15_inv01 = 1;
    24: op1_15_inv01 = 1;
    27: op1_15_inv01 = 1;
    28: op1_15_inv01 = 1;
    3: op1_15_inv01 = 1;
    31: op1_15_inv01 = 1;
    32: op1_15_inv01 = 1;
    33: op1_15_inv01 = 1;
    34: op1_15_inv01 = 1;
    37: op1_15_inv01 = 1;
    39: op1_15_inv01 = 1;
    41: op1_15_inv01 = 1;
    42: op1_15_inv01 = 1;
    46: op1_15_inv01 = 1;
    47: op1_15_inv01 = 1;
    50: op1_15_inv01 = 1;
    52: op1_15_inv01 = 1;
    55: op1_15_inv01 = 1;
    57: op1_15_inv01 = 1;
    58: op1_15_inv01 = 1;
    60: op1_15_inv01 = 1;
    61: op1_15_inv01 = 1;
    62: op1_15_inv01 = 1;
    63: op1_15_inv01 = 1;
    64: op1_15_inv01 = 1;
    65: op1_15_inv01 = 1;
    67: op1_15_inv01 = 1;
    68: op1_15_inv01 = 1;
    72: op1_15_inv01 = 1;
    76: op1_15_inv01 = 1;
    77: op1_15_inv01 = 1;
    79: op1_15_inv01 = 1;
    80: op1_15_inv01 = 1;
    81: op1_15_inv01 = 1;
    84: op1_15_inv01 = 1;
    85: op1_15_inv01 = 1;
    86: op1_15_inv01 = 1;
    88: op1_15_inv01 = 1;
    91: op1_15_inv01 = 1;
    92: op1_15_inv01 = 1;
    93: op1_15_inv01 = 1;
    95: op1_15_inv01 = 1;
    default: op1_15_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の2番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in02 = imem02_in[51:48];
    5: op1_15_in02 = reg_0721;
    6: op1_15_in02 = imem03_in[95:92];
    7: op1_15_in02 = imem05_in[47:44];
    8: op1_15_in02 = reg_0196;
    9: op1_15_in02 = imem00_in[51:48];
    10: op1_15_in02 = reg_0282;
    11: op1_15_in02 = reg_0151;
    12: op1_15_in02 = reg_0811;
    13: op1_15_in02 = reg_0264;
    14: op1_15_in02 = reg_0367;
    15: op1_15_in02 = reg_0508;
    16: op1_15_in02 = reg_0393;
    17: op1_15_in02 = reg_0656;
    18: op1_15_in02 = reg_0588;
    19: op1_15_in02 = reg_0497;
    20: op1_15_in02 = reg_0298;
    80: op1_15_in02 = reg_0298;
    21: op1_15_in02 = reg_0753;
    22: op1_15_in02 = reg_0663;
    23: op1_15_in02 = imem00_in[99:96];
    24: op1_15_in02 = imem01_in[87:84];
    25: op1_15_in02 = reg_0604;
    26: op1_15_in02 = reg_0518;
    27: op1_15_in02 = imem04_in[35:32];
    28: op1_15_in02 = reg_0730;
    3: op1_15_in02 = imem07_in[91:88];
    29: op1_15_in02 = reg_0124;
    30: op1_15_in02 = imem05_in[87:84];
    31: op1_15_in02 = reg_0144;
    32: op1_15_in02 = reg_0030;
    33: op1_15_in02 = imem04_in[127:124];
    34: op1_15_in02 = reg_0299;
    35: op1_15_in02 = imem05_in[71:68];
    36: op1_15_in02 = reg_0440;
    37: op1_15_in02 = imem07_in[27:24];
    38: op1_15_in02 = imem00_in[107:104];
    51: op1_15_in02 = imem00_in[107:104];
    39: op1_15_in02 = imem00_in[71:68];
    40: op1_15_in02 = reg_0365;
    41: op1_15_in02 = imem06_in[23:20];
    42: op1_15_in02 = reg_0183;
    43: op1_15_in02 = imem00_in[91:88];
    44: op1_15_in02 = reg_0575;
    45: op1_15_in02 = reg_0215;
    46: op1_15_in02 = imem00_in[75:72];
    47: op1_15_in02 = reg_0591;
    48: op1_15_in02 = reg_0432;
    49: op1_15_in02 = reg_0770;
    50: op1_15_in02 = reg_0225;
    82: op1_15_in02 = reg_0225;
    52: op1_15_in02 = imem01_in[83:80];
    53: op1_15_in02 = reg_0306;
    54: op1_15_in02 = reg_0810;
    55: op1_15_in02 = imem05_in[3:0];
    56: op1_15_in02 = reg_0792;
    57: op1_15_in02 = reg_0488;
    58: op1_15_in02 = reg_0029;
    59: op1_15_in02 = imem05_in[55:52];
    60: op1_15_in02 = imem07_in[79:76];
    61: op1_15_in02 = imem00_in[67:64];
    62: op1_15_in02 = imem03_in[15:12];
    63: op1_15_in02 = reg_0281;
    64: op1_15_in02 = reg_0385;
    65: op1_15_in02 = reg_0303;
    66: op1_15_in02 = reg_0009;
    67: op1_15_in02 = imem00_in[35:32];
    68: op1_15_in02 = imem02_in[59:56];
    69: op1_15_in02 = reg_0774;
    70: op1_15_in02 = imem00_in[103:100];
    71: op1_15_in02 = reg_0002;
    72: op1_15_in02 = reg_0500;
    73: op1_15_in02 = reg_0307;
    74: op1_15_in02 = reg_0515;
    75: op1_15_in02 = reg_0448;
    76: op1_15_in02 = reg_0574;
    77: op1_15_in02 = reg_0395;
    78: op1_15_in02 = reg_0568;
    79: op1_15_in02 = imem06_in[43:40];
    81: op1_15_in02 = reg_0589;
    83: op1_15_in02 = reg_0684;
    84: op1_15_in02 = reg_0337;
    85: op1_15_in02 = reg_0050;
    86: op1_15_in02 = reg_0120;
    87: op1_15_in02 = reg_0666;
    88: op1_15_in02 = reg_0031;
    89: op1_15_in02 = imem04_in[3:0];
    90: op1_15_in02 = imem04_in[55:52];
    91: op1_15_in02 = imem00_in[115:112];
    92: op1_15_in02 = imem00_in[27:24];
    93: op1_15_in02 = reg_0006;
    95: op1_15_in02 = reg_0268;
    default: op1_15_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv02 = 1;
    5: op1_15_inv02 = 1;
    7: op1_15_inv02 = 1;
    9: op1_15_inv02 = 1;
    10: op1_15_inv02 = 1;
    13: op1_15_inv02 = 1;
    18: op1_15_inv02 = 1;
    19: op1_15_inv02 = 1;
    20: op1_15_inv02 = 1;
    22: op1_15_inv02 = 1;
    23: op1_15_inv02 = 1;
    25: op1_15_inv02 = 1;
    27: op1_15_inv02 = 1;
    3: op1_15_inv02 = 1;
    29: op1_15_inv02 = 1;
    35: op1_15_inv02 = 1;
    37: op1_15_inv02 = 1;
    38: op1_15_inv02 = 1;
    39: op1_15_inv02 = 1;
    42: op1_15_inv02 = 1;
    44: op1_15_inv02 = 1;
    45: op1_15_inv02 = 1;
    47: op1_15_inv02 = 1;
    48: op1_15_inv02 = 1;
    50: op1_15_inv02 = 1;
    52: op1_15_inv02 = 1;
    53: op1_15_inv02 = 1;
    55: op1_15_inv02 = 1;
    56: op1_15_inv02 = 1;
    60: op1_15_inv02 = 1;
    63: op1_15_inv02 = 1;
    64: op1_15_inv02 = 1;
    66: op1_15_inv02 = 1;
    68: op1_15_inv02 = 1;
    71: op1_15_inv02 = 1;
    72: op1_15_inv02 = 1;
    73: op1_15_inv02 = 1;
    74: op1_15_inv02 = 1;
    75: op1_15_inv02 = 1;
    78: op1_15_inv02 = 1;
    79: op1_15_inv02 = 1;
    83: op1_15_inv02 = 1;
    86: op1_15_inv02 = 1;
    89: op1_15_inv02 = 1;
    93: op1_15_inv02 = 1;
    95: op1_15_inv02 = 1;
    default: op1_15_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の3番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in03 = imem02_in[71:68];
    5: op1_15_in03 = reg_0724;
    6: op1_15_in03 = imem03_in[107:104];
    7: op1_15_in03 = imem05_in[51:48];
    8: op1_15_in03 = reg_0205;
    9: op1_15_in03 = imem00_in[83:80];
    39: op1_15_in03 = imem00_in[83:80];
    10: op1_15_in03 = reg_0306;
    11: op1_15_in03 = reg_0152;
    12: op1_15_in03 = reg_0001;
    13: op1_15_in03 = reg_0260;
    14: op1_15_in03 = reg_0039;
    74: op1_15_in03 = reg_0039;
    15: op1_15_in03 = reg_0105;
    16: op1_15_in03 = reg_0361;
    17: op1_15_in03 = reg_0652;
    18: op1_15_in03 = reg_0387;
    19: op1_15_in03 = reg_0229;
    20: op1_15_in03 = reg_0050;
    21: op1_15_in03 = reg_0812;
    22: op1_15_in03 = reg_0320;
    23: op1_15_in03 = reg_0695;
    24: op1_15_in03 = imem01_in[103:100];
    25: op1_15_in03 = reg_0629;
    26: op1_15_in03 = reg_0097;
    27: op1_15_in03 = imem04_in[99:96];
    90: op1_15_in03 = imem04_in[99:96];
    28: op1_15_in03 = reg_0721;
    3: op1_15_in03 = imem07_in[99:96];
    29: op1_15_in03 = reg_0100;
    30: op1_15_in03 = imem05_in[99:96];
    31: op1_15_in03 = reg_0815;
    32: op1_15_in03 = imem07_in[43:40];
    33: op1_15_in03 = reg_0087;
    34: op1_15_in03 = reg_0066;
    73: op1_15_in03 = reg_0066;
    35: op1_15_in03 = reg_0798;
    36: op1_15_in03 = reg_0442;
    37: op1_15_in03 = imem07_in[35:32];
    38: op1_15_in03 = reg_0696;
    40: op1_15_in03 = reg_0342;
    41: op1_15_in03 = imem06_in[31:28];
    42: op1_15_in03 = reg_0166;
    43: op1_15_in03 = reg_0686;
    44: op1_15_in03 = reg_0564;
    45: op1_15_in03 = reg_0265;
    46: op1_15_in03 = imem00_in[79:76];
    61: op1_15_in03 = imem00_in[79:76];
    47: op1_15_in03 = reg_0750;
    48: op1_15_in03 = reg_0305;
    49: op1_15_in03 = reg_0093;
    50: op1_15_in03 = reg_0423;
    82: op1_15_in03 = reg_0423;
    51: op1_15_in03 = reg_0694;
    52: op1_15_in03 = imem02_in[11:8];
    53: op1_15_in03 = reg_0567;
    54: op1_15_in03 = imem04_in[63:60];
    55: op1_15_in03 = imem05_in[87:84];
    56: op1_15_in03 = reg_0781;
    57: op1_15_in03 = reg_0281;
    58: op1_15_in03 = imem07_in[7:4];
    59: op1_15_in03 = imem05_in[103:100];
    60: op1_15_in03 = imem07_in[87:84];
    62: op1_15_in03 = imem03_in[27:24];
    63: op1_15_in03 = reg_0357;
    64: op1_15_in03 = reg_0747;
    65: op1_15_in03 = reg_0280;
    66: op1_15_in03 = imem04_in[11:8];
    67: op1_15_in03 = imem00_in[43:40];
    68: op1_15_in03 = imem02_in[63:60];
    69: op1_15_in03 = reg_0416;
    70: op1_15_in03 = reg_0749;
    91: op1_15_in03 = reg_0749;
    71: op1_15_in03 = reg_0003;
    72: op1_15_in03 = reg_0308;
    75: op1_15_in03 = reg_0167;
    76: op1_15_in03 = reg_0054;
    77: op1_15_in03 = reg_0569;
    78: op1_15_in03 = reg_0572;
    79: op1_15_in03 = imem06_in[63:60];
    80: op1_15_in03 = reg_0354;
    81: op1_15_in03 = reg_0599;
    83: op1_15_in03 = reg_0690;
    84: op1_15_in03 = reg_0736;
    85: op1_15_in03 = reg_0626;
    86: op1_15_in03 = reg_0107;
    87: op1_15_in03 = reg_0128;
    88: op1_15_in03 = reg_0704;
    89: op1_15_in03 = imem04_in[51:48];
    92: op1_15_in03 = imem00_in[47:44];
    93: op1_15_in03 = reg_0693;
    95: op1_15_in03 = reg_0139;
    default: op1_15_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv03 = 1;
    7: op1_15_inv03 = 1;
    8: op1_15_inv03 = 1;
    10: op1_15_inv03 = 1;
    16: op1_15_inv03 = 1;
    18: op1_15_inv03 = 1;
    19: op1_15_inv03 = 1;
    20: op1_15_inv03 = 1;
    24: op1_15_inv03 = 1;
    26: op1_15_inv03 = 1;
    30: op1_15_inv03 = 1;
    32: op1_15_inv03 = 1;
    33: op1_15_inv03 = 1;
    34: op1_15_inv03 = 1;
    35: op1_15_inv03 = 1;
    37: op1_15_inv03 = 1;
    38: op1_15_inv03 = 1;
    39: op1_15_inv03 = 1;
    43: op1_15_inv03 = 1;
    44: op1_15_inv03 = 1;
    45: op1_15_inv03 = 1;
    48: op1_15_inv03 = 1;
    51: op1_15_inv03 = 1;
    52: op1_15_inv03 = 1;
    56: op1_15_inv03 = 1;
    61: op1_15_inv03 = 1;
    63: op1_15_inv03 = 1;
    64: op1_15_inv03 = 1;
    65: op1_15_inv03 = 1;
    72: op1_15_inv03 = 1;
    73: op1_15_inv03 = 1;
    76: op1_15_inv03 = 1;
    77: op1_15_inv03 = 1;
    80: op1_15_inv03 = 1;
    81: op1_15_inv03 = 1;
    82: op1_15_inv03 = 1;
    83: op1_15_inv03 = 1;
    85: op1_15_inv03 = 1;
    87: op1_15_inv03 = 1;
    88: op1_15_inv03 = 1;
    89: op1_15_inv03 = 1;
    91: op1_15_inv03 = 1;
    92: op1_15_inv03 = 1;
    95: op1_15_inv03 = 1;
    default: op1_15_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の4番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in04 = imem02_in[87:84];
    5: op1_15_in04 = reg_0706;
    6: op1_15_in04 = reg_0582;
    7: op1_15_in04 = imem05_in[67:64];
    8: op1_15_in04 = imem01_in[11:8];
    9: op1_15_in04 = imem00_in[107:104];
    61: op1_15_in04 = imem00_in[107:104];
    10: op1_15_in04 = reg_0276;
    11: op1_15_in04 = reg_0144;
    12: op1_15_in04 = reg_0013;
    13: op1_15_in04 = reg_0732;
    14: op1_15_in04 = reg_0753;
    15: op1_15_in04 = reg_0107;
    16: op1_15_in04 = reg_0396;
    17: op1_15_in04 = reg_0325;
    18: op1_15_in04 = reg_0362;
    19: op1_15_in04 = reg_0514;
    20: op1_15_in04 = reg_0065;
    21: op1_15_in04 = reg_0036;
    22: op1_15_in04 = reg_0354;
    23: op1_15_in04 = reg_0682;
    24: op1_15_in04 = imem01_in[123:120];
    25: op1_15_in04 = reg_0607;
    26: op1_15_in04 = reg_0540;
    27: op1_15_in04 = reg_0291;
    28: op1_15_in04 = reg_0714;
    3: op1_15_in04 = imem07_in[107:104];
    29: op1_15_in04 = reg_0101;
    30: op1_15_in04 = reg_0781;
    31: op1_15_in04 = reg_0033;
    32: op1_15_in04 = imem07_in[51:48];
    33: op1_15_in04 = reg_0523;
    34: op1_15_in04 = reg_0289;
    35: op1_15_in04 = reg_0796;
    36: op1_15_in04 = reg_0438;
    37: op1_15_in04 = imem07_in[39:36];
    38: op1_15_in04 = reg_0694;
    39: op1_15_in04 = imem00_in[119:116];
    40: op1_15_in04 = reg_0322;
    41: op1_15_in04 = imem06_in[71:68];
    42: op1_15_in04 = reg_0170;
    43: op1_15_in04 = reg_0691;
    44: op1_15_in04 = reg_0568;
    45: op1_15_in04 = reg_0774;
    46: op1_15_in04 = imem00_in[83:80];
    47: op1_15_in04 = reg_0749;
    48: op1_15_in04 = reg_0616;
    49: op1_15_in04 = reg_0740;
    50: op1_15_in04 = reg_0422;
    51: op1_15_in04 = reg_0689;
    52: op1_15_in04 = imem02_in[31:28];
    53: op1_15_in04 = reg_0123;
    54: op1_15_in04 = imem04_in[75:72];
    55: op1_15_in04 = imem05_in[119:116];
    56: op1_15_in04 = reg_0270;
    57: op1_15_in04 = reg_0588;
    58: op1_15_in04 = imem07_in[15:12];
    59: op1_15_in04 = reg_0113;
    60: op1_15_in04 = imem07_in[127:124];
    62: op1_15_in04 = imem03_in[47:44];
    63: op1_15_in04 = reg_0331;
    64: op1_15_in04 = reg_0570;
    65: op1_15_in04 = reg_0071;
    66: op1_15_in04 = imem04_in[19:16];
    67: op1_15_in04 = imem00_in[75:72];
    68: op1_15_in04 = imem02_in[71:68];
    69: op1_15_in04 = imem05_in[59:56];
    70: op1_15_in04 = reg_0692;
    71: op1_15_in04 = reg_0007;
    72: op1_15_in04 = reg_0280;
    73: op1_15_in04 = imem05_in[55:52];
    74: op1_15_in04 = reg_0700;
    75: op1_15_in04 = reg_0176;
    76: op1_15_in04 = reg_0217;
    77: op1_15_in04 = reg_0387;
    78: op1_15_in04 = reg_0569;
    79: op1_15_in04 = imem06_in[87:84];
    80: op1_15_in04 = reg_0402;
    81: op1_15_in04 = reg_0604;
    82: op1_15_in04 = reg_0306;
    83: op1_15_in04 = reg_0758;
    84: op1_15_in04 = reg_0788;
    85: op1_15_in04 = reg_0614;
    86: op1_15_in04 = reg_0676;
    87: op1_15_in04 = reg_0070;
    88: op1_15_in04 = reg_0075;
    89: op1_15_in04 = imem04_in[59:56];
    90: op1_15_in04 = imem04_in[115:112];
    91: op1_15_in04 = reg_0453;
    92: op1_15_in04 = imem00_in[51:48];
    93: op1_15_in04 = reg_0077;
    95: op1_15_in04 = reg_0175;
    default: op1_15_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv04 = 1;
    6: op1_15_inv04 = 1;
    7: op1_15_inv04 = 1;
    11: op1_15_inv04 = 1;
    13: op1_15_inv04 = 1;
    14: op1_15_inv04 = 1;
    15: op1_15_inv04 = 1;
    19: op1_15_inv04 = 1;
    21: op1_15_inv04 = 1;
    25: op1_15_inv04 = 1;
    26: op1_15_inv04 = 1;
    30: op1_15_inv04 = 1;
    31: op1_15_inv04 = 1;
    33: op1_15_inv04 = 1;
    34: op1_15_inv04 = 1;
    35: op1_15_inv04 = 1;
    37: op1_15_inv04 = 1;
    41: op1_15_inv04 = 1;
    42: op1_15_inv04 = 1;
    44: op1_15_inv04 = 1;
    45: op1_15_inv04 = 1;
    48: op1_15_inv04 = 1;
    51: op1_15_inv04 = 1;
    53: op1_15_inv04 = 1;
    55: op1_15_inv04 = 1;
    56: op1_15_inv04 = 1;
    58: op1_15_inv04 = 1;
    59: op1_15_inv04 = 1;
    61: op1_15_inv04 = 1;
    64: op1_15_inv04 = 1;
    66: op1_15_inv04 = 1;
    70: op1_15_inv04 = 1;
    71: op1_15_inv04 = 1;
    73: op1_15_inv04 = 1;
    74: op1_15_inv04 = 1;
    75: op1_15_inv04 = 1;
    79: op1_15_inv04 = 1;
    80: op1_15_inv04 = 1;
    81: op1_15_inv04 = 1;
    82: op1_15_inv04 = 1;
    84: op1_15_inv04 = 1;
    87: op1_15_inv04 = 1;
    93: op1_15_inv04 = 1;
    default: op1_15_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の5番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in05 = reg_0651;
    5: op1_15_in05 = reg_0436;
    6: op1_15_in05 = reg_0596;
    7: op1_15_in05 = imem05_in[75:72];
    8: op1_15_in05 = imem01_in[23:20];
    9: op1_15_in05 = reg_0672;
    10: op1_15_in05 = reg_0295;
    11: op1_15_in05 = imem06_in[7:4];
    12: op1_15_in05 = reg_0801;
    78: op1_15_in05 = reg_0801;
    13: op1_15_in05 = reg_0132;
    14: op1_15_in05 = reg_0035;
    31: op1_15_in05 = reg_0035;
    15: op1_15_in05 = reg_0126;
    16: op1_15_in05 = reg_0331;
    17: op1_15_in05 = reg_0347;
    18: op1_15_in05 = reg_0369;
    19: op1_15_in05 = reg_0500;
    33: op1_15_in05 = reg_0500;
    20: op1_15_in05 = reg_0076;
    21: op1_15_in05 = imem07_in[15:12];
    22: op1_15_in05 = reg_0324;
    23: op1_15_in05 = reg_0693;
    24: op1_15_in05 = reg_0235;
    25: op1_15_in05 = reg_0620;
    26: op1_15_in05 = reg_0535;
    27: op1_15_in05 = reg_0292;
    28: op1_15_in05 = reg_0703;
    3: op1_15_in05 = reg_0441;
    29: op1_15_in05 = reg_0109;
    30: op1_15_in05 = reg_0490;
    32: op1_15_in05 = imem07_in[95:92];
    34: op1_15_in05 = reg_0254;
    35: op1_15_in05 = reg_0795;
    36: op1_15_in05 = reg_0179;
    37: op1_15_in05 = imem07_in[47:44];
    38: op1_15_in05 = reg_0679;
    51: op1_15_in05 = reg_0679;
    39: op1_15_in05 = imem00_in[127:124];
    40: op1_15_in05 = reg_0355;
    41: op1_15_in05 = imem06_in[87:84];
    43: op1_15_in05 = reg_0668;
    44: op1_15_in05 = reg_0571;
    45: op1_15_in05 = reg_0577;
    46: op1_15_in05 = imem00_in[107:104];
    47: op1_15_in05 = reg_0384;
    63: op1_15_in05 = reg_0384;
    48: op1_15_in05 = reg_0503;
    49: op1_15_in05 = imem03_in[39:36];
    50: op1_15_in05 = reg_0054;
    52: op1_15_in05 = imem02_in[67:64];
    53: op1_15_in05 = reg_0104;
    54: op1_15_in05 = reg_0545;
    55: op1_15_in05 = reg_0215;
    56: op1_15_in05 = reg_0111;
    57: op1_15_in05 = reg_0751;
    58: op1_15_in05 = imem07_in[31:28];
    59: op1_15_in05 = reg_0790;
    60: op1_15_in05 = reg_0718;
    61: op1_15_in05 = reg_0658;
    62: op1_15_in05 = imem03_in[51:48];
    64: op1_15_in05 = reg_0013;
    65: op1_15_in05 = reg_0629;
    66: op1_15_in05 = imem04_in[47:44];
    67: op1_15_in05 = imem00_in[79:76];
    68: op1_15_in05 = imem02_in[91:88];
    69: op1_15_in05 = imem05_in[79:76];
    70: op1_15_in05 = reg_0463;
    71: op1_15_in05 = reg_0804;
    72: op1_15_in05 = reg_0052;
    73: op1_15_in05 = imem05_in[83:80];
    74: op1_15_in05 = reg_0661;
    76: op1_15_in05 = reg_0240;
    77: op1_15_in05 = reg_0396;
    79: op1_15_in05 = imem06_in[99:96];
    80: op1_15_in05 = reg_0519;
    81: op1_15_in05 = reg_0493;
    82: op1_15_in05 = reg_0511;
    83: op1_15_in05 = reg_0457;
    84: op1_15_in05 = reg_0550;
    85: op1_15_in05 = reg_0223;
    86: op1_15_in05 = imem02_in[15:12];
    87: op1_15_in05 = reg_0732;
    88: op1_15_in05 = reg_0374;
    89: op1_15_in05 = reg_0316;
    90: op1_15_in05 = reg_0247;
    91: op1_15_in05 = reg_0451;
    92: op1_15_in05 = imem00_in[75:72];
    93: op1_15_in05 = reg_0000;
    95: op1_15_in05 = reg_0089;
    default: op1_15_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv05 = 1;
    6: op1_15_inv05 = 1;
    8: op1_15_inv05 = 1;
    10: op1_15_inv05 = 1;
    11: op1_15_inv05 = 1;
    12: op1_15_inv05 = 1;
    14: op1_15_inv05 = 1;
    15: op1_15_inv05 = 1;
    17: op1_15_inv05 = 1;
    19: op1_15_inv05 = 1;
    20: op1_15_inv05 = 1;
    21: op1_15_inv05 = 1;
    22: op1_15_inv05 = 1;
    24: op1_15_inv05 = 1;
    25: op1_15_inv05 = 1;
    26: op1_15_inv05 = 1;
    3: op1_15_inv05 = 1;
    29: op1_15_inv05 = 1;
    30: op1_15_inv05 = 1;
    32: op1_15_inv05 = 1;
    34: op1_15_inv05 = 1;
    37: op1_15_inv05 = 1;
    40: op1_15_inv05 = 1;
    41: op1_15_inv05 = 1;
    43: op1_15_inv05 = 1;
    45: op1_15_inv05 = 1;
    47: op1_15_inv05 = 1;
    49: op1_15_inv05 = 1;
    50: op1_15_inv05 = 1;
    51: op1_15_inv05 = 1;
    53: op1_15_inv05 = 1;
    59: op1_15_inv05 = 1;
    61: op1_15_inv05 = 1;
    62: op1_15_inv05 = 1;
    65: op1_15_inv05 = 1;
    66: op1_15_inv05 = 1;
    68: op1_15_inv05 = 1;
    69: op1_15_inv05 = 1;
    73: op1_15_inv05 = 1;
    74: op1_15_inv05 = 1;
    77: op1_15_inv05 = 1;
    79: op1_15_inv05 = 1;
    80: op1_15_inv05 = 1;
    82: op1_15_inv05 = 1;
    83: op1_15_inv05 = 1;
    85: op1_15_inv05 = 1;
    86: op1_15_inv05 = 1;
    87: op1_15_inv05 = 1;
    95: op1_15_inv05 = 1;
    default: op1_15_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の6番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in06 = reg_0636;
    5: op1_15_in06 = reg_0422;
    3: op1_15_in06 = reg_0422;
    6: op1_15_in06 = reg_0583;
    7: op1_15_in06 = imem05_in[99:96];
    8: op1_15_in06 = imem01_in[35:32];
    9: op1_15_in06 = reg_0686;
    93: op1_15_in06 = reg_0686;
    10: op1_15_in06 = reg_0298;
    11: op1_15_in06 = imem06_in[43:40];
    12: op1_15_in06 = reg_0016;
    13: op1_15_in06 = reg_0147;
    14: op1_15_in06 = reg_0816;
    15: op1_15_in06 = imem02_in[11:8];
    16: op1_15_in06 = reg_0803;
    17: op1_15_in06 = reg_0336;
    18: op1_15_in06 = reg_0322;
    19: op1_15_in06 = reg_0824;
    20: op1_15_in06 = reg_0255;
    21: op1_15_in06 = imem07_in[39:36];
    22: op1_15_in06 = reg_0342;
    23: op1_15_in06 = reg_0672;
    24: op1_15_in06 = reg_0216;
    25: op1_15_in06 = reg_0615;
    26: op1_15_in06 = reg_0098;
    27: op1_15_in06 = imem05_in[19:16];
    28: op1_15_in06 = reg_0705;
    29: op1_15_in06 = reg_0127;
    30: op1_15_in06 = reg_0488;
    31: op1_15_in06 = reg_0621;
    32: op1_15_in06 = reg_0702;
    33: op1_15_in06 = reg_0295;
    34: op1_15_in06 = imem05_in[3:0];
    35: op1_15_in06 = reg_0277;
    36: op1_15_in06 = reg_0169;
    37: op1_15_in06 = imem07_in[51:48];
    38: op1_15_in06 = reg_0675;
    39: op1_15_in06 = reg_0695;
    40: op1_15_in06 = imem03_in[35:32];
    41: op1_15_in06 = imem06_in[119:116];
    43: op1_15_in06 = reg_0669;
    44: op1_15_in06 = reg_0385;
    45: op1_15_in06 = reg_0370;
    46: op1_15_in06 = imem00_in[115:112];
    47: op1_15_in06 = reg_0387;
    48: op1_15_in06 = imem04_in[35:32];
    49: op1_15_in06 = imem03_in[63:60];
    50: op1_15_in06 = reg_0217;
    82: op1_15_in06 = reg_0217;
    51: op1_15_in06 = reg_0477;
    52: op1_15_in06 = imem02_in[71:68];
    53: op1_15_in06 = reg_0660;
    54: op1_15_in06 = reg_0043;
    55: op1_15_in06 = reg_0309;
    56: op1_15_in06 = reg_0790;
    57: op1_15_in06 = reg_0331;
    58: op1_15_in06 = imem07_in[67:64];
    59: op1_15_in06 = reg_0218;
    60: op1_15_in06 = reg_0253;
    61: op1_15_in06 = reg_0688;
    62: op1_15_in06 = imem03_in[83:80];
    63: op1_15_in06 = reg_0517;
    84: op1_15_in06 = reg_0517;
    64: op1_15_in06 = reg_0804;
    65: op1_15_in06 = reg_0297;
    72: op1_15_in06 = reg_0297;
    66: op1_15_in06 = imem04_in[63:60];
    67: op1_15_in06 = imem00_in[95:92];
    68: op1_15_in06 = imem02_in[107:104];
    69: op1_15_in06 = reg_0736;
    70: op1_15_in06 = reg_0457;
    71: op1_15_in06 = reg_0802;
    73: op1_15_in06 = imem05_in[87:84];
    74: op1_15_in06 = reg_0367;
    76: op1_15_in06 = reg_0502;
    77: op1_15_in06 = reg_0006;
    78: op1_15_in06 = imem04_in[3:0];
    79: op1_15_in06 = imem06_in[111:108];
    80: op1_15_in06 = reg_0630;
    81: op1_15_in06 = reg_0319;
    83: op1_15_in06 = reg_0475;
    85: op1_15_in06 = reg_0062;
    86: op1_15_in06 = imem02_in[27:24];
    87: op1_15_in06 = reg_0552;
    88: op1_15_in06 = reg_0345;
    89: op1_15_in06 = reg_0544;
    90: op1_15_in06 = reg_0262;
    91: op1_15_in06 = reg_0461;
    92: op1_15_in06 = imem00_in[83:80];
    95: op1_15_in06 = reg_0236;
    default: op1_15_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv06 = 1;
    8: op1_15_inv06 = 1;
    10: op1_15_inv06 = 1;
    11: op1_15_inv06 = 1;
    19: op1_15_inv06 = 1;
    20: op1_15_inv06 = 1;
    22: op1_15_inv06 = 1;
    23: op1_15_inv06 = 1;
    24: op1_15_inv06 = 1;
    26: op1_15_inv06 = 1;
    27: op1_15_inv06 = 1;
    31: op1_15_inv06 = 1;
    32: op1_15_inv06 = 1;
    33: op1_15_inv06 = 1;
    34: op1_15_inv06 = 1;
    35: op1_15_inv06 = 1;
    36: op1_15_inv06 = 1;
    38: op1_15_inv06 = 1;
    39: op1_15_inv06 = 1;
    43: op1_15_inv06 = 1;
    44: op1_15_inv06 = 1;
    45: op1_15_inv06 = 1;
    49: op1_15_inv06 = 1;
    50: op1_15_inv06 = 1;
    51: op1_15_inv06 = 1;
    52: op1_15_inv06 = 1;
    56: op1_15_inv06 = 1;
    58: op1_15_inv06 = 1;
    59: op1_15_inv06 = 1;
    61: op1_15_inv06 = 1;
    62: op1_15_inv06 = 1;
    63: op1_15_inv06 = 1;
    64: op1_15_inv06 = 1;
    66: op1_15_inv06 = 1;
    67: op1_15_inv06 = 1;
    68: op1_15_inv06 = 1;
    70: op1_15_inv06 = 1;
    71: op1_15_inv06 = 1;
    74: op1_15_inv06 = 1;
    76: op1_15_inv06 = 1;
    78: op1_15_inv06 = 1;
    79: op1_15_inv06 = 1;
    80: op1_15_inv06 = 1;
    81: op1_15_inv06 = 1;
    88: op1_15_inv06 = 1;
    95: op1_15_inv06 = 1;
    default: op1_15_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の7番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in07 = reg_0652;
    5: op1_15_in07 = reg_0440;
    6: op1_15_in07 = reg_0568;
    7: op1_15_in07 = reg_0791;
    8: op1_15_in07 = imem01_in[43:40];
    9: op1_15_in07 = reg_0691;
    10: op1_15_in07 = reg_0061;
    11: op1_15_in07 = imem06_in[67:64];
    12: op1_15_in07 = reg_0809;
    13: op1_15_in07 = reg_0149;
    14: op1_15_in07 = reg_0814;
    15: op1_15_in07 = imem02_in[31:28];
    16: op1_15_in07 = reg_0807;
    77: op1_15_in07 = reg_0807;
    17: op1_15_in07 = reg_0097;
    18: op1_15_in07 = reg_0312;
    19: op1_15_in07 = reg_0778;
    20: op1_15_in07 = imem05_in[75:72];
    21: op1_15_in07 = imem07_in[111:108];
    22: op1_15_in07 = reg_0328;
    23: op1_15_in07 = reg_0676;
    24: op1_15_in07 = reg_0247;
    25: op1_15_in07 = reg_0379;
    26: op1_15_in07 = reg_0757;
    27: op1_15_in07 = imem05_in[95:92];
    28: op1_15_in07 = reg_0424;
    3: op1_15_in07 = reg_0433;
    29: op1_15_in07 = imem02_in[35:32];
    86: op1_15_in07 = imem02_in[35:32];
    30: op1_15_in07 = reg_0788;
    31: op1_15_in07 = reg_0616;
    32: op1_15_in07 = reg_0703;
    33: op1_15_in07 = reg_0050;
    72: op1_15_in07 = reg_0050;
    34: op1_15_in07 = imem05_in[15:12];
    35: op1_15_in07 = reg_0132;
    37: op1_15_in07 = imem07_in[79:76];
    38: op1_15_in07 = reg_0688;
    39: op1_15_in07 = reg_0697;
    40: op1_15_in07 = imem03_in[71:68];
    41: op1_15_in07 = reg_0628;
    43: op1_15_in07 = reg_0478;
    44: op1_15_in07 = reg_0376;
    45: op1_15_in07 = reg_0329;
    46: op1_15_in07 = reg_0693;
    47: op1_15_in07 = reg_0396;
    48: op1_15_in07 = imem04_in[43:40];
    49: op1_15_in07 = imem03_in[67:64];
    50: op1_15_in07 = reg_0567;
    82: op1_15_in07 = reg_0567;
    51: op1_15_in07 = reg_0479;
    52: op1_15_in07 = imem02_in[91:88];
    53: op1_15_in07 = reg_0669;
    54: op1_15_in07 = reg_0088;
    55: op1_15_in07 = reg_0226;
    56: op1_15_in07 = reg_0279;
    57: op1_15_in07 = reg_0561;
    58: op1_15_in07 = imem07_in[123:120];
    59: op1_15_in07 = reg_0099;
    60: op1_15_in07 = reg_0266;
    61: op1_15_in07 = reg_0465;
    62: op1_15_in07 = reg_0317;
    63: op1_15_in07 = reg_0398;
    64: op1_15_in07 = reg_0801;
    65: op1_15_in07 = reg_0074;
    66: op1_15_in07 = imem04_in[79:76];
    67: op1_15_in07 = imem00_in[119:116];
    68: op1_15_in07 = imem02_in[119:116];
    69: op1_15_in07 = reg_0782;
    70: op1_15_in07 = reg_0466;
    71: op1_15_in07 = reg_0016;
    73: op1_15_in07 = imem05_in[103:100];
    74: op1_15_in07 = reg_0391;
    76: op1_15_in07 = reg_0248;
    78: op1_15_in07 = imem04_in[11:8];
    79: op1_15_in07 = reg_0265;
    80: op1_15_in07 = reg_0608;
    81: op1_15_in07 = reg_0591;
    83: op1_15_in07 = reg_0458;
    84: op1_15_in07 = reg_0215;
    85: op1_15_in07 = reg_0585;
    87: op1_15_in07 = reg_0245;
    88: op1_15_in07 = reg_0361;
    89: op1_15_in07 = reg_0058;
    90: op1_15_in07 = reg_0535;
    91: op1_15_in07 = reg_0477;
    92: op1_15_in07 = imem00_in[107:104];
    93: op1_15_in07 = reg_0749;
    95: op1_15_in07 = reg_0142;
    default: op1_15_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv07 = 1;
    7: op1_15_inv07 = 1;
    10: op1_15_inv07 = 1;
    17: op1_15_inv07 = 1;
    19: op1_15_inv07 = 1;
    20: op1_15_inv07 = 1;
    21: op1_15_inv07 = 1;
    23: op1_15_inv07 = 1;
    24: op1_15_inv07 = 1;
    27: op1_15_inv07 = 1;
    28: op1_15_inv07 = 1;
    3: op1_15_inv07 = 1;
    30: op1_15_inv07 = 1;
    38: op1_15_inv07 = 1;
    41: op1_15_inv07 = 1;
    43: op1_15_inv07 = 1;
    44: op1_15_inv07 = 1;
    45: op1_15_inv07 = 1;
    47: op1_15_inv07 = 1;
    48: op1_15_inv07 = 1;
    49: op1_15_inv07 = 1;
    50: op1_15_inv07 = 1;
    52: op1_15_inv07 = 1;
    53: op1_15_inv07 = 1;
    55: op1_15_inv07 = 1;
    57: op1_15_inv07 = 1;
    58: op1_15_inv07 = 1;
    59: op1_15_inv07 = 1;
    65: op1_15_inv07 = 1;
    66: op1_15_inv07 = 1;
    68: op1_15_inv07 = 1;
    70: op1_15_inv07 = 1;
    72: op1_15_inv07 = 1;
    78: op1_15_inv07 = 1;
    79: op1_15_inv07 = 1;
    80: op1_15_inv07 = 1;
    82: op1_15_inv07 = 1;
    83: op1_15_inv07 = 1;
    84: op1_15_inv07 = 1;
    86: op1_15_inv07 = 1;
    87: op1_15_inv07 = 1;
    89: op1_15_inv07 = 1;
    93: op1_15_inv07 = 1;
    default: op1_15_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の8番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in08 = reg_0352;
    5: op1_15_in08 = reg_0444;
    6: op1_15_in08 = reg_0587;
    7: op1_15_in08 = reg_0482;
    8: op1_15_in08 = imem01_in[47:44];
    9: op1_15_in08 = reg_0688;
    10: op1_15_in08 = reg_0046;
    11: op1_15_in08 = imem06_in[111:108];
    12: op1_15_in08 = imem04_in[3:0];
    13: op1_15_in08 = reg_0145;
    14: op1_15_in08 = reg_0750;
    15: op1_15_in08 = imem02_in[39:36];
    16: op1_15_in08 = reg_0799;
    17: op1_15_in08 = reg_0087;
    18: op1_15_in08 = reg_0019;
    19: op1_15_in08 = reg_0507;
    20: op1_15_in08 = imem05_in[91:88];
    21: op1_15_in08 = reg_0716;
    22: op1_15_in08 = reg_0336;
    23: op1_15_in08 = reg_0670;
    24: op1_15_in08 = reg_0238;
    25: op1_15_in08 = reg_0405;
    26: op1_15_in08 = reg_0538;
    27: op1_15_in08 = reg_0793;
    28: op1_15_in08 = reg_0432;
    3: op1_15_in08 = reg_0448;
    29: op1_15_in08 = imem02_in[59:56];
    30: op1_15_in08 = reg_0785;
    31: op1_15_in08 = reg_0633;
    32: op1_15_in08 = reg_0709;
    33: op1_15_in08 = reg_0278;
    34: op1_15_in08 = imem05_in[67:64];
    35: op1_15_in08 = reg_0133;
    37: op1_15_in08 = imem07_in[107:104];
    38: op1_15_in08 = reg_0673;
    39: op1_15_in08 = reg_0681;
    46: op1_15_in08 = reg_0681;
    40: op1_15_in08 = imem03_in[95:92];
    41: op1_15_in08 = reg_0613;
    43: op1_15_in08 = reg_0196;
    44: op1_15_in08 = reg_0397;
    45: op1_15_in08 = reg_0753;
    47: op1_15_in08 = reg_0570;
    48: op1_15_in08 = imem04_in[47:44];
    49: op1_15_in08 = imem03_in[83:80];
    50: op1_15_in08 = reg_0244;
    51: op1_15_in08 = reg_0459;
    52: op1_15_in08 = imem02_in[95:92];
    53: op1_15_in08 = reg_0676;
    54: op1_15_in08 = reg_0555;
    55: op1_15_in08 = reg_0224;
    56: op1_15_in08 = reg_0249;
    57: op1_15_in08 = reg_0392;
    58: op1_15_in08 = reg_0720;
    59: op1_15_in08 = reg_0103;
    60: op1_15_in08 = reg_0436;
    61: op1_15_in08 = reg_0451;
    62: op1_15_in08 = reg_0599;
    63: op1_15_in08 = reg_0393;
    64: op1_15_in08 = reg_0004;
    77: op1_15_in08 = reg_0004;
    65: op1_15_in08 = reg_0050;
    66: op1_15_in08 = imem04_in[115:112];
    67: op1_15_in08 = reg_0697;
    68: op1_15_in08 = reg_0650;
    69: op1_15_in08 = reg_0489;
    70: op1_15_in08 = reg_0473;
    71: op1_15_in08 = reg_0010;
    72: op1_15_in08 = reg_0622;
    73: op1_15_in08 = imem06_in[87:84];
    74: op1_15_in08 = reg_0328;
    76: op1_15_in08 = reg_0424;
    78: op1_15_in08 = imem04_in[79:76];
    79: op1_15_in08 = reg_0659;
    80: op1_15_in08 = reg_0583;
    87: op1_15_in08 = reg_0583;
    81: op1_15_in08 = reg_0528;
    82: op1_15_in08 = reg_0502;
    83: op1_15_in08 = reg_0187;
    84: op1_15_in08 = reg_0252;
    85: op1_15_in08 = reg_0065;
    86: op1_15_in08 = imem02_in[43:40];
    88: op1_15_in08 = reg_0356;
    89: op1_15_in08 = reg_0542;
    90: op1_15_in08 = reg_0558;
    91: op1_15_in08 = reg_0469;
    92: op1_15_in08 = imem00_in[115:112];
    93: op1_15_in08 = reg_0658;
    95: op1_15_in08 = reg_0327;
    default: op1_15_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv08 = 1;
    7: op1_15_inv08 = 1;
    12: op1_15_inv08 = 1;
    14: op1_15_inv08 = 1;
    15: op1_15_inv08 = 1;
    16: op1_15_inv08 = 1;
    19: op1_15_inv08 = 1;
    27: op1_15_inv08 = 1;
    30: op1_15_inv08 = 1;
    31: op1_15_inv08 = 1;
    33: op1_15_inv08 = 1;
    34: op1_15_inv08 = 1;
    43: op1_15_inv08 = 1;
    46: op1_15_inv08 = 1;
    47: op1_15_inv08 = 1;
    49: op1_15_inv08 = 1;
    50: op1_15_inv08 = 1;
    51: op1_15_inv08 = 1;
    52: op1_15_inv08 = 1;
    53: op1_15_inv08 = 1;
    55: op1_15_inv08 = 1;
    58: op1_15_inv08 = 1;
    64: op1_15_inv08 = 1;
    67: op1_15_inv08 = 1;
    68: op1_15_inv08 = 1;
    69: op1_15_inv08 = 1;
    70: op1_15_inv08 = 1;
    73: op1_15_inv08 = 1;
    76: op1_15_inv08 = 1;
    79: op1_15_inv08 = 1;
    80: op1_15_inv08 = 1;
    81: op1_15_inv08 = 1;
    82: op1_15_inv08 = 1;
    84: op1_15_inv08 = 1;
    85: op1_15_inv08 = 1;
    86: op1_15_inv08 = 1;
    88: op1_15_inv08 = 1;
    90: op1_15_inv08 = 1;
    91: op1_15_inv08 = 1;
    92: op1_15_inv08 = 1;
    default: op1_15_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の9番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in09 = reg_0324;
    5: op1_15_in09 = reg_0427;
    6: op1_15_in09 = reg_0592;
    7: op1_15_in09 = reg_0797;
    69: op1_15_in09 = reg_0797;
    8: op1_15_in09 = imem01_in[87:84];
    9: op1_15_in09 = reg_0453;
    10: op1_15_in09 = reg_0065;
    11: op1_15_in09 = reg_0630;
    12: op1_15_in09 = imem04_in[7:4];
    13: op1_15_in09 = reg_0136;
    14: op1_15_in09 = imem07_in[23:20];
    15: op1_15_in09 = imem02_in[59:56];
    16: op1_15_in09 = reg_0010;
    17: op1_15_in09 = imem03_in[11:8];
    18: op1_15_in09 = reg_0001;
    19: op1_15_in09 = reg_0215;
    20: op1_15_in09 = reg_0798;
    21: op1_15_in09 = reg_0719;
    22: op1_15_in09 = reg_0081;
    23: op1_15_in09 = reg_0691;
    93: op1_15_in09 = reg_0691;
    24: op1_15_in09 = reg_0219;
    25: op1_15_in09 = reg_0375;
    26: op1_15_in09 = reg_0532;
    27: op1_15_in09 = reg_0782;
    28: op1_15_in09 = reg_0426;
    3: op1_15_in09 = reg_0167;
    29: op1_15_in09 = imem02_in[83:80];
    30: op1_15_in09 = reg_0736;
    31: op1_15_in09 = reg_0632;
    32: op1_15_in09 = reg_0711;
    33: op1_15_in09 = reg_0079;
    34: op1_15_in09 = reg_0483;
    35: op1_15_in09 = reg_0139;
    37: op1_15_in09 = imem07_in[123:120];
    38: op1_15_in09 = reg_0450;
    39: op1_15_in09 = reg_0679;
    40: op1_15_in09 = reg_0039;
    41: op1_15_in09 = reg_0608;
    43: op1_15_in09 = reg_0212;
    44: op1_15_in09 = reg_0386;
    45: op1_15_in09 = reg_0621;
    46: op1_15_in09 = reg_0672;
    47: op1_15_in09 = reg_0016;
    48: op1_15_in09 = imem04_in[55:52];
    49: op1_15_in09 = imem03_in[95:92];
    50: op1_15_in09 = reg_0248;
    51: op1_15_in09 = reg_0200;
    52: op1_15_in09 = imem02_in[99:96];
    53: op1_15_in09 = reg_0121;
    54: op1_15_in09 = reg_0554;
    55: op1_15_in09 = reg_0258;
    56: op1_15_in09 = reg_0086;
    57: op1_15_in09 = reg_0376;
    58: op1_15_in09 = reg_0731;
    59: op1_15_in09 = reg_0279;
    60: op1_15_in09 = reg_0444;
    61: op1_15_in09 = reg_0455;
    62: op1_15_in09 = reg_0319;
    63: op1_15_in09 = reg_0570;
    64: op1_15_in09 = imem04_in[11:8];
    65: op1_15_in09 = reg_0614;
    66: op1_15_in09 = imem04_in[123:120];
    67: op1_15_in09 = reg_0686;
    68: op1_15_in09 = reg_0753;
    70: op1_15_in09 = reg_0474;
    71: op1_15_in09 = imem04_in[35:32];
    72: op1_15_in09 = reg_0259;
    73: op1_15_in09 = imem06_in[115:112];
    74: op1_15_in09 = imem07_in[31:28];
    76: op1_15_in09 = reg_0243;
    77: op1_15_in09 = imem04_in[3:0];
    78: op1_15_in09 = imem04_in[91:88];
    79: op1_15_in09 = reg_0748;
    80: op1_15_in09 = reg_0573;
    81: op1_15_in09 = reg_0350;
    82: op1_15_in09 = reg_0216;
    83: op1_15_in09 = imem01_in[43:40];
    84: op1_15_in09 = reg_0491;
    85: op1_15_in09 = reg_0622;
    86: op1_15_in09 = imem02_in[91:88];
    87: op1_15_in09 = reg_0229;
    88: op1_15_in09 = reg_0594;
    89: op1_15_in09 = reg_0523;
    90: op1_15_in09 = reg_0429;
    91: op1_15_in09 = reg_0466;
    92: op1_15_in09 = reg_0695;
    95: op1_15_in09 = reg_0182;
    default: op1_15_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv09 = 1;
    5: op1_15_inv09 = 1;
    6: op1_15_inv09 = 1;
    7: op1_15_inv09 = 1;
    9: op1_15_inv09 = 1;
    11: op1_15_inv09 = 1;
    13: op1_15_inv09 = 1;
    15: op1_15_inv09 = 1;
    16: op1_15_inv09 = 1;
    19: op1_15_inv09 = 1;
    22: op1_15_inv09 = 1;
    25: op1_15_inv09 = 1;
    27: op1_15_inv09 = 1;
    28: op1_15_inv09 = 1;
    29: op1_15_inv09 = 1;
    31: op1_15_inv09 = 1;
    37: op1_15_inv09 = 1;
    40: op1_15_inv09 = 1;
    43: op1_15_inv09 = 1;
    45: op1_15_inv09 = 1;
    46: op1_15_inv09 = 1;
    50: op1_15_inv09 = 1;
    54: op1_15_inv09 = 1;
    56: op1_15_inv09 = 1;
    57: op1_15_inv09 = 1;
    58: op1_15_inv09 = 1;
    60: op1_15_inv09 = 1;
    64: op1_15_inv09 = 1;
    67: op1_15_inv09 = 1;
    72: op1_15_inv09 = 1;
    77: op1_15_inv09 = 1;
    82: op1_15_inv09 = 1;
    83: op1_15_inv09 = 1;
    84: op1_15_inv09 = 1;
    87: op1_15_inv09 = 1;
    88: op1_15_inv09 = 1;
    89: op1_15_inv09 = 1;
    91: op1_15_inv09 = 1;
    default: op1_15_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の10番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in10 = reg_0353;
    5: op1_15_in10 = reg_0420;
    6: op1_15_in10 = reg_0591;
    7: op1_15_in10 = reg_0789;
    34: op1_15_in10 = reg_0789;
    8: op1_15_in10 = imem01_in[95:92];
    9: op1_15_in10 = reg_0466;
    10: op1_15_in10 = reg_0058;
    11: op1_15_in10 = reg_0624;
    12: op1_15_in10 = imem04_in[55:52];
    71: op1_15_in10 = imem04_in[55:52];
    13: op1_15_in10 = reg_0150;
    14: op1_15_in10 = imem07_in[95:92];
    15: op1_15_in10 = imem02_in[91:88];
    16: op1_15_in10 = reg_0004;
    17: op1_15_in10 = imem03_in[35:32];
    18: op1_15_in10 = reg_0003;
    19: op1_15_in10 = reg_0220;
    82: op1_15_in10 = reg_0220;
    20: op1_15_in10 = reg_0482;
    21: op1_15_in10 = reg_0731;
    22: op1_15_in10 = reg_0532;
    23: op1_15_in10 = reg_0465;
    24: op1_15_in10 = reg_0123;
    25: op1_15_in10 = reg_0399;
    81: op1_15_in10 = reg_0399;
    26: op1_15_in10 = imem03_in[3:0];
    27: op1_15_in10 = reg_0783;
    28: op1_15_in10 = reg_0418;
    3: op1_15_in10 = reg_0183;
    29: op1_15_in10 = imem02_in[87:84];
    30: op1_15_in10 = reg_0285;
    31: op1_15_in10 = reg_0627;
    32: op1_15_in10 = reg_0432;
    90: op1_15_in10 = reg_0432;
    33: op1_15_in10 = reg_0077;
    35: op1_15_in10 = reg_0140;
    37: op1_15_in10 = reg_0730;
    38: op1_15_in10 = reg_0471;
    39: op1_15_in10 = reg_0677;
    40: op1_15_in10 = reg_0755;
    41: op1_15_in10 = reg_0402;
    43: op1_15_in10 = imem01_in[59:56];
    44: op1_15_in10 = reg_0389;
    45: op1_15_in10 = reg_0037;
    46: op1_15_in10 = reg_0680;
    47: op1_15_in10 = reg_0010;
    48: op1_15_in10 = imem04_in[95:92];
    49: op1_15_in10 = imem03_in[99:96];
    50: op1_15_in10 = reg_0234;
    51: op1_15_in10 = reg_0203;
    52: op1_15_in10 = imem02_in[107:104];
    53: op1_15_in10 = imem02_in[47:44];
    54: op1_15_in10 = reg_0057;
    55: op1_15_in10 = reg_0257;
    56: op1_15_in10 = reg_0151;
    57: op1_15_in10 = reg_0803;
    58: op1_15_in10 = reg_0721;
    59: op1_15_in10 = reg_0089;
    60: op1_15_in10 = reg_0267;
    61: op1_15_in10 = reg_0200;
    62: op1_15_in10 = reg_0329;
    63: op1_15_in10 = reg_0801;
    64: op1_15_in10 = imem04_in[79:76];
    65: op1_15_in10 = reg_0301;
    66: op1_15_in10 = reg_0328;
    67: op1_15_in10 = reg_0633;
    68: op1_15_in10 = reg_0352;
    69: op1_15_in10 = reg_0276;
    84: op1_15_in10 = reg_0276;
    70: op1_15_in10 = reg_0478;
    72: op1_15_in10 = reg_0640;
    73: op1_15_in10 = imem06_in[123:120];
    74: op1_15_in10 = imem07_in[83:80];
    76: op1_15_in10 = reg_0122;
    77: op1_15_in10 = imem04_in[7:4];
    78: op1_15_in10 = imem04_in[103:100];
    79: op1_15_in10 = reg_0375;
    80: op1_15_in10 = reg_0029;
    83: op1_15_in10 = imem01_in[63:60];
    85: op1_15_in10 = reg_0774;
    86: op1_15_in10 = imem02_in[95:92];
    87: op1_15_in10 = reg_0393;
    88: op1_15_in10 = reg_0043;
    89: op1_15_in10 = reg_0551;
    91: op1_15_in10 = reg_0475;
    92: op1_15_in10 = reg_0697;
    93: op1_15_in10 = reg_0016;
    95: op1_15_in10 = reg_0066;
    default: op1_15_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv10 = 1;
    7: op1_15_inv10 = 1;
    10: op1_15_inv10 = 1;
    11: op1_15_inv10 = 1;
    12: op1_15_inv10 = 1;
    13: op1_15_inv10 = 1;
    14: op1_15_inv10 = 1;
    15: op1_15_inv10 = 1;
    16: op1_15_inv10 = 1;
    17: op1_15_inv10 = 1;
    19: op1_15_inv10 = 1;
    20: op1_15_inv10 = 1;
    21: op1_15_inv10 = 1;
    25: op1_15_inv10 = 1;
    3: op1_15_inv10 = 1;
    32: op1_15_inv10 = 1;
    33: op1_15_inv10 = 1;
    35: op1_15_inv10 = 1;
    37: op1_15_inv10 = 1;
    38: op1_15_inv10 = 1;
    41: op1_15_inv10 = 1;
    44: op1_15_inv10 = 1;
    45: op1_15_inv10 = 1;
    46: op1_15_inv10 = 1;
    48: op1_15_inv10 = 1;
    49: op1_15_inv10 = 1;
    54: op1_15_inv10 = 1;
    55: op1_15_inv10 = 1;
    56: op1_15_inv10 = 1;
    59: op1_15_inv10 = 1;
    62: op1_15_inv10 = 1;
    64: op1_15_inv10 = 1;
    69: op1_15_inv10 = 1;
    76: op1_15_inv10 = 1;
    78: op1_15_inv10 = 1;
    79: op1_15_inv10 = 1;
    82: op1_15_inv10 = 1;
    83: op1_15_inv10 = 1;
    87: op1_15_inv10 = 1;
    88: op1_15_inv10 = 1;
    89: op1_15_inv10 = 1;
    93: op1_15_inv10 = 1;
    default: op1_15_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の11番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in11 = reg_0342;
    5: op1_15_in11 = reg_0174;
    6: op1_15_in11 = reg_0597;
    7: op1_15_in11 = reg_0492;
    8: op1_15_in11 = imem01_in[111:108];
    9: op1_15_in11 = reg_0480;
    10: op1_15_in11 = reg_0076;
    11: op1_15_in11 = reg_0621;
    12: op1_15_in11 = imem04_in[59:56];
    71: op1_15_in11 = imem04_in[59:56];
    13: op1_15_in11 = reg_0143;
    14: op1_15_in11 = imem07_in[127:124];
    15: op1_15_in11 = imem02_in[111:108];
    16: op1_15_in11 = imem04_in[39:36];
    17: op1_15_in11 = imem03_in[43:40];
    18: op1_15_in11 = reg_0801;
    57: op1_15_in11 = reg_0801;
    19: op1_15_in11 = reg_0236;
    20: op1_15_in11 = reg_0795;
    21: op1_15_in11 = reg_0721;
    22: op1_15_in11 = imem03_in[67:64];
    23: op1_15_in11 = reg_0453;
    24: op1_15_in11 = reg_0105;
    25: op1_15_in11 = reg_0406;
    26: op1_15_in11 = imem03_in[11:8];
    27: op1_15_in11 = reg_0790;
    28: op1_15_in11 = reg_0437;
    3: op1_15_in11 = reg_0166;
    29: op1_15_in11 = imem02_in[95:92];
    30: op1_15_in11 = reg_0136;
    31: op1_15_in11 = reg_0402;
    32: op1_15_in11 = reg_0427;
    33: op1_15_in11 = reg_0288;
    34: op1_15_in11 = reg_0783;
    35: op1_15_in11 = reg_0155;
    37: op1_15_in11 = reg_0710;
    38: op1_15_in11 = reg_0200;
    39: op1_15_in11 = reg_0678;
    40: op1_15_in11 = reg_0373;
    41: op1_15_in11 = reg_0377;
    43: op1_15_in11 = imem01_in[103:100];
    44: op1_15_in11 = reg_0015;
    45: op1_15_in11 = reg_0231;
    46: op1_15_in11 = reg_0673;
    76: op1_15_in11 = reg_0673;
    47: op1_15_in11 = imem04_in[7:4];
    48: op1_15_in11 = imem05_in[27:24];
    49: op1_15_in11 = imem03_in[103:100];
    50: op1_15_in11 = reg_0506;
    51: op1_15_in11 = reg_0201;
    52: op1_15_in11 = imem02_in[119:116];
    53: op1_15_in11 = imem02_in[87:84];
    54: op1_15_in11 = reg_0523;
    55: op1_15_in11 = reg_0148;
    56: op1_15_in11 = reg_0156;
    58: op1_15_in11 = reg_0705;
    59: op1_15_in11 = reg_0133;
    60: op1_15_in11 = reg_0172;
    61: op1_15_in11 = reg_0187;
    62: op1_15_in11 = reg_0281;
    63: op1_15_in11 = reg_0810;
    64: op1_15_in11 = imem04_in[91:88];
    65: op1_15_in11 = reg_0585;
    66: op1_15_in11 = reg_0542;
    67: op1_15_in11 = reg_0247;
    68: op1_15_in11 = reg_0345;
    69: op1_15_in11 = reg_0249;
    70: op1_15_in11 = reg_0211;
    72: op1_15_in11 = reg_0109;
    88: op1_15_in11 = reg_0109;
    73: op1_15_in11 = reg_0346;
    74: op1_15_in11 = reg_0441;
    77: op1_15_in11 = imem04_in[11:8];
    78: op1_15_in11 = imem04_in[107:104];
    79: op1_15_in11 = reg_0035;
    80: op1_15_in11 = reg_0484;
    81: op1_15_in11 = reg_0595;
    82: op1_15_in11 = reg_0504;
    83: op1_15_in11 = imem01_in[119:116];
    84: op1_15_in11 = reg_0781;
    85: op1_15_in11 = reg_0259;
    86: op1_15_in11 = imem02_in[103:100];
    87: op1_15_in11 = reg_0369;
    89: op1_15_in11 = reg_0510;
    90: op1_15_in11 = reg_0079;
    91: op1_15_in11 = reg_0203;
    92: op1_15_in11 = reg_0698;
    93: op1_15_in11 = reg_0171;
    95: op1_15_in11 = reg_0183;
    default: op1_15_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv11 = 1;
    5: op1_15_inv11 = 1;
    6: op1_15_inv11 = 1;
    7: op1_15_inv11 = 1;
    8: op1_15_inv11 = 1;
    9: op1_15_inv11 = 1;
    10: op1_15_inv11 = 1;
    11: op1_15_inv11 = 1;
    13: op1_15_inv11 = 1;
    15: op1_15_inv11 = 1;
    17: op1_15_inv11 = 1;
    21: op1_15_inv11 = 1;
    22: op1_15_inv11 = 1;
    23: op1_15_inv11 = 1;
    25: op1_15_inv11 = 1;
    29: op1_15_inv11 = 1;
    31: op1_15_inv11 = 1;
    32: op1_15_inv11 = 1;
    33: op1_15_inv11 = 1;
    34: op1_15_inv11 = 1;
    37: op1_15_inv11 = 1;
    39: op1_15_inv11 = 1;
    48: op1_15_inv11 = 1;
    50: op1_15_inv11 = 1;
    52: op1_15_inv11 = 1;
    53: op1_15_inv11 = 1;
    54: op1_15_inv11 = 1;
    56: op1_15_inv11 = 1;
    57: op1_15_inv11 = 1;
    60: op1_15_inv11 = 1;
    63: op1_15_inv11 = 1;
    65: op1_15_inv11 = 1;
    66: op1_15_inv11 = 1;
    67: op1_15_inv11 = 1;
    70: op1_15_inv11 = 1;
    73: op1_15_inv11 = 1;
    74: op1_15_inv11 = 1;
    77: op1_15_inv11 = 1;
    78: op1_15_inv11 = 1;
    79: op1_15_inv11 = 1;
    80: op1_15_inv11 = 1;
    81: op1_15_inv11 = 1;
    83: op1_15_inv11 = 1;
    84: op1_15_inv11 = 1;
    85: op1_15_inv11 = 1;
    87: op1_15_inv11 = 1;
    88: op1_15_inv11 = 1;
    90: op1_15_inv11 = 1;
    91: op1_15_inv11 = 1;
    95: op1_15_inv11 = 1;
    default: op1_15_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の12番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in12 = reg_0083;
    5: op1_15_in12 = reg_0181;
    6: op1_15_in12 = reg_0588;
    7: op1_15_in12 = reg_0267;
    8: op1_15_in12 = imem01_in[127:124];
    9: op1_15_in12 = reg_0473;
    10: op1_15_in12 = reg_0043;
    66: op1_15_in12 = reg_0043;
    11: op1_15_in12 = reg_0619;
    12: op1_15_in12 = imem04_in[67:64];
    13: op1_15_in12 = reg_0155;
    14: op1_15_in12 = reg_0719;
    15: op1_15_in12 = reg_0642;
    16: op1_15_in12 = imem04_in[99:96];
    17: op1_15_in12 = imem03_in[91:88];
    18: op1_15_in12 = reg_0279;
    19: op1_15_in12 = reg_0243;
    20: op1_15_in12 = reg_0495;
    21: op1_15_in12 = reg_0729;
    22: op1_15_in12 = imem03_in[119:116];
    23: op1_15_in12 = reg_0469;
    24: op1_15_in12 = reg_0108;
    25: op1_15_in12 = reg_0380;
    26: op1_15_in12 = imem03_in[15:12];
    27: op1_15_in12 = reg_0486;
    28: op1_15_in12 = reg_0420;
    3: op1_15_in12 = reg_0178;
    29: op1_15_in12 = reg_0653;
    30: op1_15_in12 = reg_0133;
    31: op1_15_in12 = reg_0318;
    32: op1_15_in12 = reg_0431;
    33: op1_15_in12 = imem05_in[7:4];
    34: op1_15_in12 = reg_0786;
    35: op1_15_in12 = reg_0137;
    56: op1_15_in12 = reg_0137;
    37: op1_15_in12 = reg_0724;
    38: op1_15_in12 = reg_0210;
    39: op1_15_in12 = reg_0468;
    40: op1_15_in12 = reg_0562;
    41: op1_15_in12 = reg_0329;
    43: op1_15_in12 = imem01_in[111:108];
    44: op1_15_in12 = reg_0799;
    45: op1_15_in12 = reg_0632;
    46: op1_15_in12 = reg_0669;
    47: op1_15_in12 = imem04_in[15:12];
    48: op1_15_in12 = imem05_in[39:36];
    49: op1_15_in12 = reg_0586;
    50: op1_15_in12 = reg_0424;
    82: op1_15_in12 = reg_0424;
    51: op1_15_in12 = reg_0192;
    52: op1_15_in12 = reg_0658;
    92: op1_15_in12 = reg_0658;
    53: op1_15_in12 = imem02_in[91:88];
    54: op1_15_in12 = reg_0058;
    55: op1_15_in12 = reg_0135;
    57: op1_15_in12 = reg_0008;
    58: op1_15_in12 = reg_0436;
    59: op1_15_in12 = reg_0139;
    60: op1_15_in12 = reg_0170;
    61: op1_15_in12 = reg_0194;
    91: op1_15_in12 = reg_0194;
    62: op1_15_in12 = reg_0395;
    63: op1_15_in12 = reg_0009;
    64: op1_15_in12 = imem04_in[111:108];
    65: op1_15_in12 = reg_0065;
    67: op1_15_in12 = reg_0692;
    68: op1_15_in12 = reg_0565;
    69: op1_15_in12 = reg_0307;
    70: op1_15_in12 = reg_0206;
    71: op1_15_in12 = imem04_in[87:84];
    72: op1_15_in12 = reg_0091;
    73: op1_15_in12 = reg_0577;
    74: op1_15_in12 = reg_0064;
    76: op1_15_in12 = reg_0073;
    77: op1_15_in12 = imem04_in[27:24];
    78: op1_15_in12 = reg_0554;
    79: op1_15_in12 = reg_0573;
    80: op1_15_in12 = reg_0787;
    81: op1_15_in12 = reg_0648;
    83: op1_15_in12 = reg_0102;
    84: op1_15_in12 = reg_0830;
    85: op1_15_in12 = imem05_in[11:8];
    86: op1_15_in12 = imem02_in[119:116];
    87: op1_15_in12 = reg_0285;
    88: op1_15_in12 = reg_0136;
    89: op1_15_in12 = reg_0516;
    90: op1_15_in12 = reg_0305;
    93: op1_15_in12 = reg_0455;
    95: op1_15_in12 = reg_0141;
    default: op1_15_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv12 = 1;
    6: op1_15_inv12 = 1;
    9: op1_15_inv12 = 1;
    12: op1_15_inv12 = 1;
    13: op1_15_inv12 = 1;
    14: op1_15_inv12 = 1;
    16: op1_15_inv12 = 1;
    18: op1_15_inv12 = 1;
    19: op1_15_inv12 = 1;
    21: op1_15_inv12 = 1;
    22: op1_15_inv12 = 1;
    23: op1_15_inv12 = 1;
    25: op1_15_inv12 = 1;
    26: op1_15_inv12 = 1;
    3: op1_15_inv12 = 1;
    33: op1_15_inv12 = 1;
    34: op1_15_inv12 = 1;
    35: op1_15_inv12 = 1;
    37: op1_15_inv12 = 1;
    40: op1_15_inv12 = 1;
    47: op1_15_inv12 = 1;
    48: op1_15_inv12 = 1;
    49: op1_15_inv12 = 1;
    53: op1_15_inv12 = 1;
    54: op1_15_inv12 = 1;
    59: op1_15_inv12 = 1;
    61: op1_15_inv12 = 1;
    62: op1_15_inv12 = 1;
    65: op1_15_inv12 = 1;
    67: op1_15_inv12 = 1;
    69: op1_15_inv12 = 1;
    71: op1_15_inv12 = 1;
    72: op1_15_inv12 = 1;
    73: op1_15_inv12 = 1;
    74: op1_15_inv12 = 1;
    76: op1_15_inv12 = 1;
    81: op1_15_inv12 = 1;
    83: op1_15_inv12 = 1;
    84: op1_15_inv12 = 1;
    85: op1_15_inv12 = 1;
    86: op1_15_inv12 = 1;
    87: op1_15_inv12 = 1;
    default: op1_15_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の13番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in13 = reg_0081;
    5: op1_15_in13 = reg_0160;
    6: op1_15_in13 = reg_0384;
    7: op1_15_in13 = reg_0241;
    8: op1_15_in13 = reg_0504;
    9: op1_15_in13 = reg_0470;
    10: op1_15_in13 = reg_0072;
    11: op1_15_in13 = reg_0612;
    12: op1_15_in13 = imem04_in[71:68];
    13: op1_15_in13 = imem06_in[31:28];
    14: op1_15_in13 = reg_0705;
    37: op1_15_in13 = reg_0705;
    15: op1_15_in13 = reg_0658;
    16: op1_15_in13 = imem04_in[119:116];
    77: op1_15_in13 = imem04_in[119:116];
    17: op1_15_in13 = imem03_in[115:112];
    18: op1_15_in13 = reg_0282;
    19: op1_15_in13 = reg_0123;
    20: op1_15_in13 = reg_0787;
    21: op1_15_in13 = reg_0713;
    22: op1_15_in13 = reg_0571;
    23: op1_15_in13 = reg_0473;
    24: op1_15_in13 = reg_0100;
    25: op1_15_in13 = reg_0031;
    26: op1_15_in13 = imem03_in[31:28];
    27: op1_15_in13 = reg_0742;
    28: op1_15_in13 = reg_0172;
    29: op1_15_in13 = reg_0637;
    30: op1_15_in13 = reg_0150;
    31: op1_15_in13 = reg_0370;
    32: op1_15_in13 = reg_0179;
    33: op1_15_in13 = imem05_in[15:12];
    34: op1_15_in13 = reg_0489;
    35: op1_15_in13 = reg_0029;
    38: op1_15_in13 = reg_0187;
    39: op1_15_in13 = reg_0452;
    40: op1_15_in13 = reg_0389;
    41: op1_15_in13 = reg_0401;
    43: op1_15_in13 = reg_0501;
    44: op1_15_in13 = reg_0016;
    45: op1_15_in13 = imem07_in[11:8];
    46: op1_15_in13 = reg_0465;
    47: op1_15_in13 = imem04_in[19:16];
    48: op1_15_in13 = imem05_in[47:44];
    49: op1_15_in13 = reg_0599;
    50: op1_15_in13 = reg_0243;
    51: op1_15_in13 = imem01_in[3:0];
    52: op1_15_in13 = reg_0584;
    53: op1_15_in13 = imem02_in[127:124];
    54: op1_15_in13 = reg_0429;
    55: op1_15_in13 = reg_0128;
    56: op1_15_in13 = reg_0402;
    57: op1_15_in13 = reg_0015;
    58: op1_15_in13 = reg_0051;
    59: op1_15_in13 = reg_0129;
    61: op1_15_in13 = reg_0201;
    62: op1_15_in13 = reg_0575;
    63: op1_15_in13 = reg_0010;
    64: op1_15_in13 = reg_0537;
    65: op1_15_in13 = reg_0069;
    66: op1_15_in13 = reg_0554;
    67: op1_15_in13 = reg_0463;
    68: op1_15_in13 = reg_0356;
    69: op1_15_in13 = reg_0383;
    70: op1_15_in13 = imem01_in[59:56];
    71: op1_15_in13 = imem04_in[111:108];
    72: op1_15_in13 = reg_0735;
    73: op1_15_in13 = reg_0817;
    74: op1_15_in13 = reg_0333;
    76: op1_15_in13 = reg_0675;
    78: op1_15_in13 = reg_0057;
    79: op1_15_in13 = reg_0039;
    80: op1_15_in13 = reg_0661;
    81: op1_15_in13 = reg_0028;
    82: op1_15_in13 = reg_0505;
    83: op1_15_in13 = reg_0101;
    84: op1_15_in13 = reg_0154;
    85: op1_15_in13 = imem05_in[27:24];
    86: op1_15_in13 = reg_0656;
    87: op1_15_in13 = reg_0781;
    88: op1_15_in13 = reg_0757;
    89: op1_15_in13 = reg_0283;
    90: op1_15_in13 = reg_0280;
    91: op1_15_in13 = reg_0213;
    92: op1_15_in13 = reg_0063;
    93: op1_15_in13 = reg_0474;
    95: op1_15_in13 = reg_0178;
    default: op1_15_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv13 = 1;
    9: op1_15_inv13 = 1;
    10: op1_15_inv13 = 1;
    11: op1_15_inv13 = 1;
    12: op1_15_inv13 = 1;
    13: op1_15_inv13 = 1;
    14: op1_15_inv13 = 1;
    15: op1_15_inv13 = 1;
    17: op1_15_inv13 = 1;
    19: op1_15_inv13 = 1;
    20: op1_15_inv13 = 1;
    23: op1_15_inv13 = 1;
    29: op1_15_inv13 = 1;
    31: op1_15_inv13 = 1;
    32: op1_15_inv13 = 1;
    35: op1_15_inv13 = 1;
    37: op1_15_inv13 = 1;
    38: op1_15_inv13 = 1;
    39: op1_15_inv13 = 1;
    43: op1_15_inv13 = 1;
    44: op1_15_inv13 = 1;
    45: op1_15_inv13 = 1;
    46: op1_15_inv13 = 1;
    51: op1_15_inv13 = 1;
    52: op1_15_inv13 = 1;
    54: op1_15_inv13 = 1;
    55: op1_15_inv13 = 1;
    56: op1_15_inv13 = 1;
    57: op1_15_inv13 = 1;
    58: op1_15_inv13 = 1;
    59: op1_15_inv13 = 1;
    61: op1_15_inv13 = 1;
    62: op1_15_inv13 = 1;
    63: op1_15_inv13 = 1;
    64: op1_15_inv13 = 1;
    65: op1_15_inv13 = 1;
    66: op1_15_inv13 = 1;
    67: op1_15_inv13 = 1;
    69: op1_15_inv13 = 1;
    70: op1_15_inv13 = 1;
    71: op1_15_inv13 = 1;
    72: op1_15_inv13 = 1;
    73: op1_15_inv13 = 1;
    76: op1_15_inv13 = 1;
    83: op1_15_inv13 = 1;
    90: op1_15_inv13 = 1;
    91: op1_15_inv13 = 1;
    93: op1_15_inv13 = 1;
    default: op1_15_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の14番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in14 = reg_0086;
    5: op1_15_in14 = reg_0183;
    6: op1_15_in14 = reg_0362;
    7: op1_15_in14 = reg_0148;
    8: op1_15_in14 = reg_0512;
    9: op1_15_in14 = reg_0452;
    10: op1_15_in14 = imem05_in[43:40];
    11: op1_15_in14 = reg_0408;
    12: op1_15_in14 = imem04_in[75:72];
    13: op1_15_in14 = imem06_in[51:48];
    14: op1_15_in14 = reg_0713;
    37: op1_15_in14 = reg_0713;
    15: op1_15_in14 = reg_0653;
    16: op1_15_in14 = reg_0552;
    17: op1_15_in14 = reg_0586;
    18: op1_15_in14 = reg_0285;
    69: op1_15_in14 = reg_0285;
    19: op1_15_in14 = reg_0127;
    20: op1_15_in14 = reg_0736;
    21: op1_15_in14 = reg_0430;
    22: op1_15_in14 = reg_0580;
    23: op1_15_in14 = reg_0456;
    24: op1_15_in14 = reg_0101;
    25: op1_15_in14 = reg_0747;
    26: op1_15_in14 = imem03_in[51:48];
    27: op1_15_in14 = reg_0732;
    28: op1_15_in14 = reg_0160;
    29: op1_15_in14 = reg_0649;
    30: op1_15_in14 = reg_0151;
    87: op1_15_in14 = reg_0151;
    31: op1_15_in14 = reg_0762;
    32: op1_15_in14 = reg_0167;
    33: op1_15_in14 = imem05_in[39:36];
    34: op1_15_in14 = reg_0486;
    35: op1_15_in14 = reg_0031;
    41: op1_15_in14 = reg_0031;
    38: op1_15_in14 = reg_0193;
    39: op1_15_in14 = reg_0200;
    40: op1_15_in14 = reg_0007;
    43: op1_15_in14 = reg_0487;
    44: op1_15_in14 = reg_0810;
    45: op1_15_in14 = imem07_in[23:20];
    46: op1_15_in14 = reg_0461;
    47: op1_15_in14 = imem04_in[23:20];
    48: op1_15_in14 = imem05_in[67:64];
    49: op1_15_in14 = reg_0583;
    50: op1_15_in14 = reg_0111;
    51: op1_15_in14 = imem01_in[55:52];
    52: op1_15_in14 = reg_0346;
    53: op1_15_in14 = reg_0642;
    54: op1_15_in14 = reg_0076;
    55: op1_15_in14 = reg_0140;
    95: op1_15_in14 = reg_0140;
    56: op1_15_in14 = reg_0369;
    57: op1_15_in14 = reg_0016;
    58: op1_15_in14 = reg_0440;
    59: op1_15_in14 = reg_0144;
    61: op1_15_in14 = reg_0213;
    62: op1_15_in14 = reg_0568;
    63: op1_15_in14 = imem04_in[7:4];
    64: op1_15_in14 = reg_0043;
    65: op1_15_in14 = reg_0110;
    66: op1_15_in14 = reg_0551;
    67: op1_15_in14 = reg_0465;
    68: op1_15_in14 = reg_0363;
    70: op1_15_in14 = imem01_in[63:60];
    71: op1_15_in14 = reg_0058;
    72: op1_15_in14 = reg_0143;
    84: op1_15_in14 = reg_0143;
    73: op1_15_in14 = reg_0609;
    74: op1_15_in14 = reg_0267;
    76: op1_15_in14 = reg_0671;
    77: op1_15_in14 = reg_0087;
    78: op1_15_in14 = reg_0516;
    79: op1_15_in14 = reg_0663;
    80: op1_15_in14 = reg_0174;
    81: op1_15_in14 = reg_0575;
    82: op1_15_in14 = reg_0124;
    83: op1_15_in14 = reg_0397;
    85: op1_15_in14 = imem05_in[79:76];
    86: op1_15_in14 = reg_0753;
    88: op1_15_in14 = reg_0740;
    89: op1_15_in14 = reg_0611;
    90: op1_15_in14 = reg_0052;
    91: op1_15_in14 = reg_0190;
    92: op1_15_in14 = reg_0453;
    93: op1_15_in14 = reg_0468;
    default: op1_15_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    5: op1_15_inv14 = 1;
    13: op1_15_inv14 = 1;
    14: op1_15_inv14 = 1;
    16: op1_15_inv14 = 1;
    21: op1_15_inv14 = 1;
    22: op1_15_inv14 = 1;
    26: op1_15_inv14 = 1;
    27: op1_15_inv14 = 1;
    29: op1_15_inv14 = 1;
    30: op1_15_inv14 = 1;
    31: op1_15_inv14 = 1;
    32: op1_15_inv14 = 1;
    33: op1_15_inv14 = 1;
    37: op1_15_inv14 = 1;
    38: op1_15_inv14 = 1;
    39: op1_15_inv14 = 1;
    40: op1_15_inv14 = 1;
    41: op1_15_inv14 = 1;
    44: op1_15_inv14 = 1;
    49: op1_15_inv14 = 1;
    50: op1_15_inv14 = 1;
    54: op1_15_inv14 = 1;
    56: op1_15_inv14 = 1;
    61: op1_15_inv14 = 1;
    62: op1_15_inv14 = 1;
    63: op1_15_inv14 = 1;
    65: op1_15_inv14 = 1;
    66: op1_15_inv14 = 1;
    67: op1_15_inv14 = 1;
    71: op1_15_inv14 = 1;
    72: op1_15_inv14 = 1;
    77: op1_15_inv14 = 1;
    78: op1_15_inv14 = 1;
    79: op1_15_inv14 = 1;
    81: op1_15_inv14 = 1;
    82: op1_15_inv14 = 1;
    84: op1_15_inv14 = 1;
    86: op1_15_inv14 = 1;
    87: op1_15_inv14 = 1;
    88: op1_15_inv14 = 1;
    90: op1_15_inv14 = 1;
    91: op1_15_inv14 = 1;
    92: op1_15_inv14 = 1;
    95: op1_15_inv14 = 1;
    default: op1_15_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の15番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in15 = reg_0087;
    6: op1_15_in15 = reg_0322;
    7: op1_15_in15 = reg_0154;
    8: op1_15_in15 = reg_0511;
    83: op1_15_in15 = reg_0511;
    9: op1_15_in15 = reg_0200;
    10: op1_15_in15 = imem05_in[59:56];
    11: op1_15_in15 = reg_0386;
    12: op1_15_in15 = imem04_in[127:124];
    13: op1_15_in15 = reg_0613;
    14: op1_15_in15 = reg_0707;
    15: op1_15_in15 = reg_0664;
    16: op1_15_in15 = reg_0529;
    17: op1_15_in15 = reg_0585;
    18: op1_15_in15 = reg_0559;
    19: op1_15_in15 = reg_0126;
    20: op1_15_in15 = reg_0304;
    21: op1_15_in15 = reg_0419;
    22: op1_15_in15 = reg_0387;
    23: op1_15_in15 = reg_0214;
    24: op1_15_in15 = reg_0115;
    25: op1_15_in15 = reg_0816;
    26: op1_15_in15 = imem03_in[67:64];
    27: op1_15_in15 = reg_0132;
    28: op1_15_in15 = reg_0163;
    29: op1_15_in15 = reg_0652;
    30: op1_15_in15 = reg_0144;
    31: op1_15_in15 = reg_0377;
    56: op1_15_in15 = reg_0377;
    32: op1_15_in15 = reg_0177;
    33: op1_15_in15 = imem05_in[43:40];
    34: op1_15_in15 = reg_0741;
    35: op1_15_in15 = reg_0812;
    37: op1_15_in15 = reg_0718;
    38: op1_15_in15 = reg_0207;
    39: op1_15_in15 = reg_0210;
    40: op1_15_in15 = reg_0010;
    41: op1_15_in15 = reg_0621;
    43: op1_15_in15 = reg_0548;
    44: op1_15_in15 = imem04_in[35:32];
    45: op1_15_in15 = imem07_in[39:36];
    46: op1_15_in15 = reg_0481;
    47: op1_15_in15 = imem04_in[39:36];
    48: op1_15_in15 = imem05_in[95:92];
    49: op1_15_in15 = reg_0592;
    50: op1_15_in15 = reg_0116;
    51: op1_15_in15 = imem01_in[67:64];
    52: op1_15_in15 = reg_0638;
    53: op1_15_in15 = reg_0666;
    54: op1_15_in15 = reg_0611;
    55: op1_15_in15 = reg_0155;
    57: op1_15_in15 = reg_0004;
    58: op1_15_in15 = reg_0435;
    74: op1_15_in15 = reg_0435;
    59: op1_15_in15 = imem06_in[63:60];
    61: op1_15_in15 = imem01_in[43:40];
    62: op1_15_in15 = reg_0517;
    63: op1_15_in15 = imem04_in[11:8];
    64: op1_15_in15 = reg_0083;
    65: op1_15_in15 = reg_0336;
    66: op1_15_in15 = reg_0516;
    67: op1_15_in15 = reg_0475;
    68: op1_15_in15 = reg_0095;
    69: op1_15_in15 = reg_0151;
    70: op1_15_in15 = imem01_in[111:108];
    71: op1_15_in15 = reg_0556;
    72: op1_15_in15 = reg_0393;
    73: op1_15_in15 = reg_0401;
    76: op1_15_in15 = imem02_in[123:120];
    77: op1_15_in15 = reg_0554;
    78: op1_15_in15 = reg_0547;
    79: op1_15_in15 = reg_0620;
    80: op1_15_in15 = reg_0175;
    81: op1_15_in15 = reg_0417;
    82: op1_15_in15 = reg_0104;
    84: op1_15_in15 = reg_0761;
    85: op1_15_in15 = imem05_in[99:96];
    86: op1_15_in15 = reg_0075;
    87: op1_15_in15 = reg_0152;
    88: op1_15_in15 = imem03_in[43:40];
    89: op1_15_in15 = reg_0503;
    90: op1_15_in15 = reg_0076;
    91: op1_15_in15 = imem01_in[15:12];
    92: op1_15_in15 = reg_0451;
    93: op1_15_in15 = reg_0456;
    default: op1_15_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv15 = 1;
    11: op1_15_inv15 = 1;
    12: op1_15_inv15 = 1;
    14: op1_15_inv15 = 1;
    15: op1_15_inv15 = 1;
    17: op1_15_inv15 = 1;
    18: op1_15_inv15 = 1;
    20: op1_15_inv15 = 1;
    22: op1_15_inv15 = 1;
    24: op1_15_inv15 = 1;
    25: op1_15_inv15 = 1;
    28: op1_15_inv15 = 1;
    30: op1_15_inv15 = 1;
    32: op1_15_inv15 = 1;
    33: op1_15_inv15 = 1;
    35: op1_15_inv15 = 1;
    37: op1_15_inv15 = 1;
    39: op1_15_inv15 = 1;
    44: op1_15_inv15 = 1;
    50: op1_15_inv15 = 1;
    51: op1_15_inv15 = 1;
    52: op1_15_inv15 = 1;
    53: op1_15_inv15 = 1;
    54: op1_15_inv15 = 1;
    55: op1_15_inv15 = 1;
    56: op1_15_inv15 = 1;
    57: op1_15_inv15 = 1;
    58: op1_15_inv15 = 1;
    62: op1_15_inv15 = 1;
    63: op1_15_inv15 = 1;
    66: op1_15_inv15 = 1;
    67: op1_15_inv15 = 1;
    69: op1_15_inv15 = 1;
    70: op1_15_inv15 = 1;
    72: op1_15_inv15 = 1;
    73: op1_15_inv15 = 1;
    76: op1_15_inv15 = 1;
    77: op1_15_inv15 = 1;
    78: op1_15_inv15 = 1;
    80: op1_15_inv15 = 1;
    82: op1_15_inv15 = 1;
    87: op1_15_inv15 = 1;
    90: op1_15_inv15 = 1;
    default: op1_15_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の16番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in16 = imem03_in[3:0];
    6: op1_15_in16 = reg_0396;
    7: op1_15_in16 = reg_0138;
    8: op1_15_in16 = reg_0520;
    9: op1_15_in16 = reg_0208;
    10: op1_15_in16 = imem05_in[63:60];
    11: op1_15_in16 = reg_0406;
    12: op1_15_in16 = reg_0534;
    13: op1_15_in16 = reg_0609;
    14: op1_15_in16 = reg_0706;
    15: op1_15_in16 = reg_0652;
    16: op1_15_in16 = reg_0535;
    17: op1_15_in16 = reg_0595;
    18: op1_15_in16 = imem04_in[7:4];
    19: op1_15_in16 = imem02_in[55:52];
    20: op1_15_in16 = reg_0742;
    21: op1_15_in16 = reg_0446;
    22: op1_15_in16 = reg_0327;
    23: op1_15_in16 = reg_0191;
    24: op1_15_in16 = reg_0117;
    25: op1_15_in16 = reg_0036;
    26: op1_15_in16 = imem03_in[95:92];
    27: op1_15_in16 = reg_0145;
    28: op1_15_in16 = reg_0166;
    29: op1_15_in16 = reg_0357;
    30: op1_15_in16 = imem06_in[15:12];
    31: op1_15_in16 = imem06_in[35:32];
    33: op1_15_in16 = imem05_in[87:84];
    34: op1_15_in16 = reg_0527;
    35: op1_15_in16 = reg_0231;
    37: op1_15_in16 = reg_0711;
    38: op1_15_in16 = reg_0201;
    39: op1_15_in16 = reg_0187;
    40: op1_15_in16 = reg_0809;
    41: op1_15_in16 = imem07_in[27:24];
    43: op1_15_in16 = reg_0235;
    44: op1_15_in16 = imem04_in[51:48];
    45: op1_15_in16 = imem07_in[115:112];
    46: op1_15_in16 = reg_0456;
    47: op1_15_in16 = imem04_in[71:68];
    48: op1_15_in16 = imem05_in[115:112];
    49: op1_15_in16 = reg_0749;
    50: op1_15_in16 = reg_0119;
    51: op1_15_in16 = imem01_in[71:68];
    52: op1_15_in16 = reg_0417;
    53: op1_15_in16 = reg_0637;
    54: op1_15_in16 = reg_0302;
    55: op1_15_in16 = imem06_in[51:48];
    56: op1_15_in16 = reg_0371;
    57: op1_15_in16 = imem04_in[31:28];
    58: op1_15_in16 = reg_0164;
    59: op1_15_in16 = imem06_in[79:76];
    61: op1_15_in16 = imem01_in[47:44];
    62: op1_15_in16 = reg_0571;
    63: op1_15_in16 = imem04_in[35:32];
    64: op1_15_in16 = reg_0305;
    65: op1_15_in16 = reg_0111;
    66: op1_15_in16 = reg_0500;
    67: op1_15_in16 = reg_0462;
    68: op1_15_in16 = reg_0770;
    69: op1_15_in16 = reg_0139;
    70: op1_15_in16 = imem01_in[115:112];
    71: op1_15_in16 = reg_0308;
    72: op1_15_in16 = reg_0137;
    84: op1_15_in16 = reg_0137;
    73: op1_15_in16 = reg_0369;
    74: op1_15_in16 = reg_0175;
    76: op1_15_in16 = reg_0045;
    77: op1_15_in16 = reg_0077;
    78: op1_15_in16 = reg_0303;
    79: op1_15_in16 = reg_0752;
    80: op1_15_in16 = reg_0089;
    81: op1_15_in16 = reg_0572;
    82: op1_15_in16 = reg_0660;
    83: op1_15_in16 = reg_0220;
    85: op1_15_in16 = imem05_in[111:108];
    86: op1_15_in16 = reg_0087;
    87: op1_15_in16 = reg_0257;
    88: op1_15_in16 = imem03_in[115:112];
    89: op1_15_in16 = reg_0431;
    90: op1_15_in16 = reg_0616;
    91: op1_15_in16 = imem01_in[51:48];
    92: op1_15_in16 = reg_0476;
    93: op1_15_in16 = reg_0200;
    default: op1_15_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv16 = 1;
    11: op1_15_inv16 = 1;
    14: op1_15_inv16 = 1;
    15: op1_15_inv16 = 1;
    20: op1_15_inv16 = 1;
    21: op1_15_inv16 = 1;
    22: op1_15_inv16 = 1;
    23: op1_15_inv16 = 1;
    24: op1_15_inv16 = 1;
    25: op1_15_inv16 = 1;
    26: op1_15_inv16 = 1;
    28: op1_15_inv16 = 1;
    30: op1_15_inv16 = 1;
    33: op1_15_inv16 = 1;
    37: op1_15_inv16 = 1;
    39: op1_15_inv16 = 1;
    44: op1_15_inv16 = 1;
    45: op1_15_inv16 = 1;
    47: op1_15_inv16 = 1;
    48: op1_15_inv16 = 1;
    55: op1_15_inv16 = 1;
    56: op1_15_inv16 = 1;
    59: op1_15_inv16 = 1;
    63: op1_15_inv16 = 1;
    64: op1_15_inv16 = 1;
    66: op1_15_inv16 = 1;
    70: op1_15_inv16 = 1;
    71: op1_15_inv16 = 1;
    77: op1_15_inv16 = 1;
    81: op1_15_inv16 = 1;
    84: op1_15_inv16 = 1;
    85: op1_15_inv16 = 1;
    87: op1_15_inv16 = 1;
    90: op1_15_inv16 = 1;
    default: op1_15_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の17番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in17 = imem03_in[87:84];
    6: op1_15_in17 = reg_0374;
    7: op1_15_in17 = reg_0130;
    8: op1_15_in17 = reg_0509;
    9: op1_15_in17 = reg_0204;
    10: op1_15_in17 = imem05_in[75:72];
    11: op1_15_in17 = reg_0028;
    12: op1_15_in17 = reg_0535;
    13: op1_15_in17 = reg_0619;
    14: op1_15_in17 = reg_0423;
    15: op1_15_in17 = reg_0333;
    16: op1_15_in17 = reg_0532;
    17: op1_15_in17 = reg_0394;
    18: op1_15_in17 = imem04_in[15:12];
    19: op1_15_in17 = imem02_in[75:72];
    20: op1_15_in17 = reg_0735;
    21: op1_15_in17 = reg_0443;
    22: op1_15_in17 = reg_0322;
    23: op1_15_in17 = reg_0210;
    24: op1_15_in17 = reg_0121;
    25: op1_15_in17 = reg_0037;
    26: op1_15_in17 = imem03_in[111:108];
    27: op1_15_in17 = reg_0135;
    28: op1_15_in17 = reg_0164;
    29: op1_15_in17 = reg_0364;
    30: op1_15_in17 = imem06_in[23:20];
    31: op1_15_in17 = imem07_in[27:24];
    33: op1_15_in17 = imem05_in[103:100];
    34: op1_15_in17 = reg_0085;
    61: op1_15_in17 = reg_0085;
    35: op1_15_in17 = reg_0293;
    37: op1_15_in17 = reg_0422;
    38: op1_15_in17 = reg_0212;
    39: op1_15_in17 = reg_0198;
    40: op1_15_in17 = imem04_in[47:44];
    41: op1_15_in17 = imem07_in[35:32];
    43: op1_15_in17 = reg_0421;
    44: op1_15_in17 = imem04_in[59:56];
    45: op1_15_in17 = reg_0728;
    46: op1_15_in17 = reg_0458;
    47: op1_15_in17 = imem04_in[83:80];
    48: op1_15_in17 = imem05_in[123:120];
    49: op1_15_in17 = reg_0384;
    50: op1_15_in17 = reg_0112;
    65: op1_15_in17 = reg_0112;
    51: op1_15_in17 = imem01_in[111:108];
    52: op1_15_in17 = reg_0641;
    53: op1_15_in17 = reg_0656;
    54: op1_15_in17 = reg_0297;
    90: op1_15_in17 = reg_0297;
    55: op1_15_in17 = imem06_in[83:80];
    56: op1_15_in17 = reg_0069;
    57: op1_15_in17 = imem04_in[39:36];
    58: op1_15_in17 = reg_0173;
    59: op1_15_in17 = imem06_in[87:84];
    62: op1_15_in17 = reg_0562;
    63: op1_15_in17 = imem04_in[43:40];
    64: op1_15_in17 = reg_0076;
    66: op1_15_in17 = reg_0431;
    67: op1_15_in17 = reg_0472;
    68: op1_15_in17 = reg_0093;
    69: op1_15_in17 = reg_0138;
    70: op1_15_in17 = reg_0759;
    71: op1_15_in17 = reg_0280;
    72: op1_15_in17 = reg_0389;
    73: op1_15_in17 = reg_0578;
    74: op1_15_in17 = reg_0167;
    76: op1_15_in17 = reg_0534;
    77: op1_15_in17 = reg_0050;
    89: op1_15_in17 = reg_0050;
    78: op1_15_in17 = reg_0308;
    79: op1_15_in17 = imem07_in[3:0];
    80: op1_15_in17 = reg_0057;
    81: op1_15_in17 = reg_0403;
    82: op1_15_in17 = reg_0675;
    83: op1_15_in17 = reg_0670;
    84: op1_15_in17 = reg_0734;
    85: op1_15_in17 = reg_0736;
    86: op1_15_in17 = reg_0705;
    87: op1_15_in17 = imem06_in[7:4];
    88: op1_15_in17 = imem03_in[123:120];
    91: op1_15_in17 = imem01_in[55:52];
    92: op1_15_in17 = reg_0460;
    93: op1_15_in17 = reg_0205;
    default: op1_15_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv17 = 1;
    7: op1_15_inv17 = 1;
    8: op1_15_inv17 = 1;
    9: op1_15_inv17 = 1;
    10: op1_15_inv17 = 1;
    15: op1_15_inv17 = 1;
    16: op1_15_inv17 = 1;
    18: op1_15_inv17 = 1;
    21: op1_15_inv17 = 1;
    22: op1_15_inv17 = 1;
    24: op1_15_inv17 = 1;
    26: op1_15_inv17 = 1;
    30: op1_15_inv17 = 1;
    33: op1_15_inv17 = 1;
    38: op1_15_inv17 = 1;
    39: op1_15_inv17 = 1;
    41: op1_15_inv17 = 1;
    44: op1_15_inv17 = 1;
    47: op1_15_inv17 = 1;
    50: op1_15_inv17 = 1;
    51: op1_15_inv17 = 1;
    53: op1_15_inv17 = 1;
    54: op1_15_inv17 = 1;
    55: op1_15_inv17 = 1;
    58: op1_15_inv17 = 1;
    59: op1_15_inv17 = 1;
    62: op1_15_inv17 = 1;
    65: op1_15_inv17 = 1;
    66: op1_15_inv17 = 1;
    69: op1_15_inv17 = 1;
    72: op1_15_inv17 = 1;
    76: op1_15_inv17 = 1;
    77: op1_15_inv17 = 1;
    78: op1_15_inv17 = 1;
    79: op1_15_inv17 = 1;
    80: op1_15_inv17 = 1;
    81: op1_15_inv17 = 1;
    83: op1_15_inv17 = 1;
    84: op1_15_inv17 = 1;
    86: op1_15_inv17 = 1;
    87: op1_15_inv17 = 1;
    88: op1_15_inv17 = 1;
    89: op1_15_inv17 = 1;
    90: op1_15_inv17 = 1;
    91: op1_15_inv17 = 1;
    93: op1_15_inv17 = 1;
    default: op1_15_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の18番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in18 = imem03_in[119:116];
    6: op1_15_in18 = reg_0006;
    7: op1_15_in18 = reg_0155;
    8: op1_15_in18 = reg_0502;
    9: op1_15_in18 = reg_0193;
    10: op1_15_in18 = imem05_in[111:108];
    11: op1_15_in18 = reg_0747;
    12: op1_15_in18 = reg_0549;
    13: op1_15_in18 = reg_0633;
    14: op1_15_in18 = reg_0162;
    15: op1_15_in18 = reg_0088;
    16: op1_15_in18 = reg_0551;
    17: op1_15_in18 = reg_0395;
    18: op1_15_in18 = imem04_in[31:28];
    19: op1_15_in18 = imem02_in[115:112];
    20: op1_15_in18 = reg_0527;
    21: op1_15_in18 = reg_0420;
    22: op1_15_in18 = reg_0389;
    23: op1_15_in18 = reg_0187;
    24: op1_15_in18 = imem02_in[15:12];
    25: op1_15_in18 = reg_0029;
    26: op1_15_in18 = reg_0599;
    27: op1_15_in18 = reg_0136;
    29: op1_15_in18 = reg_0348;
    30: op1_15_in18 = imem06_in[63:60];
    31: op1_15_in18 = imem07_in[95:92];
    33: op1_15_in18 = imem05_in[123:120];
    34: op1_15_in18 = reg_0282;
    35: op1_15_in18 = reg_0615;
    71: op1_15_in18 = reg_0615;
    37: op1_15_in18 = reg_0447;
    38: op1_15_in18 = reg_0205;
    39: op1_15_in18 = reg_0190;
    40: op1_15_in18 = imem04_in[79:76];
    41: op1_15_in18 = imem07_in[43:40];
    43: op1_15_in18 = reg_0574;
    44: op1_15_in18 = imem04_in[63:60];
    45: op1_15_in18 = reg_0635;
    46: op1_15_in18 = reg_0188;
    47: op1_15_in18 = imem04_in[91:88];
    48: op1_15_in18 = reg_0488;
    49: op1_15_in18 = reg_0392;
    50: op1_15_in18 = reg_0114;
    51: op1_15_in18 = imem01_in[123:120];
    52: op1_15_in18 = reg_0362;
    53: op1_15_in18 = reg_0662;
    54: op1_15_in18 = reg_0074;
    55: op1_15_in18 = imem06_in[111:108];
    56: op1_15_in18 = reg_0779;
    57: op1_15_in18 = imem04_in[59:56];
    58: op1_15_in18 = reg_0184;
    59: op1_15_in18 = imem06_in[115:112];
    61: op1_15_in18 = reg_0653;
    62: op1_15_in18 = reg_0397;
    63: op1_15_in18 = imem04_in[55:52];
    64: op1_15_in18 = reg_0611;
    65: op1_15_in18 = reg_0226;
    66: op1_15_in18 = reg_0508;
    67: op1_15_in18 = reg_0474;
    68: op1_15_in18 = imem03_in[7:4];
    69: op1_15_in18 = imem06_in[39:36];
    87: op1_15_in18 = imem06_in[39:36];
    70: op1_15_in18 = reg_0388;
    72: op1_15_in18 = reg_0100;
    73: op1_15_in18 = reg_0748;
    74: op1_15_in18 = reg_0183;
    76: op1_15_in18 = reg_0325;
    77: op1_15_in18 = reg_0078;
    78: op1_15_in18 = reg_0430;
    79: op1_15_in18 = imem07_in[19:16];
    80: op1_15_in18 = reg_0249;
    81: op1_15_in18 = reg_0490;
    82: op1_15_in18 = reg_0106;
    83: op1_15_in18 = reg_0132;
    84: op1_15_in18 = imem06_in[23:20];
    85: op1_15_in18 = reg_0070;
    86: op1_15_in18 = reg_0358;
    88: op1_15_in18 = imem03_in[127:124];
    89: op1_15_in18 = reg_0626;
    90: op1_15_in18 = reg_0679;
    91: op1_15_in18 = imem01_in[71:68];
    92: op1_15_in18 = reg_0481;
    93: op1_15_in18 = reg_0232;
    default: op1_15_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    7: op1_15_inv18 = 1;
    9: op1_15_inv18 = 1;
    11: op1_15_inv18 = 1;
    12: op1_15_inv18 = 1;
    14: op1_15_inv18 = 1;
    15: op1_15_inv18 = 1;
    19: op1_15_inv18 = 1;
    21: op1_15_inv18 = 1;
    22: op1_15_inv18 = 1;
    26: op1_15_inv18 = 1;
    27: op1_15_inv18 = 1;
    29: op1_15_inv18 = 1;
    33: op1_15_inv18 = 1;
    37: op1_15_inv18 = 1;
    40: op1_15_inv18 = 1;
    41: op1_15_inv18 = 1;
    43: op1_15_inv18 = 1;
    44: op1_15_inv18 = 1;
    45: op1_15_inv18 = 1;
    46: op1_15_inv18 = 1;
    48: op1_15_inv18 = 1;
    50: op1_15_inv18 = 1;
    51: op1_15_inv18 = 1;
    52: op1_15_inv18 = 1;
    54: op1_15_inv18 = 1;
    61: op1_15_inv18 = 1;
    62: op1_15_inv18 = 1;
    64: op1_15_inv18 = 1;
    65: op1_15_inv18 = 1;
    66: op1_15_inv18 = 1;
    68: op1_15_inv18 = 1;
    70: op1_15_inv18 = 1;
    71: op1_15_inv18 = 1;
    72: op1_15_inv18 = 1;
    74: op1_15_inv18 = 1;
    79: op1_15_inv18 = 1;
    82: op1_15_inv18 = 1;
    83: op1_15_inv18 = 1;
    90: op1_15_inv18 = 1;
    91: op1_15_inv18 = 1;
    93: op1_15_inv18 = 1;
    default: op1_15_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の19番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in19 = reg_0579;
    6: op1_15_in19 = reg_0012;
    7: op1_15_in19 = imem06_in[23:20];
    8: op1_15_in19 = reg_0524;
    9: op1_15_in19 = reg_0213;
    10: op1_15_in19 = imem05_in[115:112];
    11: op1_15_in19 = reg_0813;
    12: op1_15_in19 = reg_0532;
    13: op1_15_in19 = reg_0349;
    15: op1_15_in19 = reg_0089;
    72: op1_15_in19 = reg_0089;
    16: op1_15_in19 = reg_0531;
    17: op1_15_in19 = reg_0387;
    18: op1_15_in19 = imem04_in[59:56];
    19: op1_15_in19 = reg_0645;
    51: op1_15_in19 = reg_0645;
    20: op1_15_in19 = reg_0085;
    21: op1_15_in19 = reg_0175;
    22: op1_15_in19 = reg_0019;
    49: op1_15_in19 = reg_0019;
    23: op1_15_in19 = reg_0193;
    24: op1_15_in19 = imem02_in[31:28];
    25: op1_15_in19 = reg_0038;
    26: op1_15_in19 = reg_0583;
    27: op1_15_in19 = reg_0138;
    29: op1_15_in19 = reg_0346;
    30: op1_15_in19 = reg_0610;
    54: op1_15_in19 = reg_0610;
    31: op1_15_in19 = reg_0720;
    33: op1_15_in19 = reg_0781;
    34: op1_15_in19 = reg_0269;
    35: op1_15_in19 = imem06_in[7:4];
    37: op1_15_in19 = reg_0439;
    38: op1_15_in19 = reg_0190;
    39: op1_15_in19 = reg_0232;
    40: op1_15_in19 = imem04_in[87:84];
    41: op1_15_in19 = imem07_in[47:44];
    43: op1_15_in19 = reg_0054;
    44: op1_15_in19 = imem04_in[107:104];
    45: op1_15_in19 = reg_0061;
    46: op1_15_in19 = reg_0207;
    47: op1_15_in19 = reg_0315;
    57: op1_15_in19 = reg_0315;
    48: op1_15_in19 = reg_0788;
    50: op1_15_in19 = reg_0109;
    52: op1_15_in19 = reg_0586;
    53: op1_15_in19 = reg_0427;
    55: op1_15_in19 = reg_0630;
    56: op1_15_in19 = reg_0031;
    59: op1_15_in19 = reg_0348;
    61: op1_15_in19 = reg_0778;
    62: op1_15_in19 = reg_0393;
    63: op1_15_in19 = imem04_in[83:80];
    64: op1_15_in19 = reg_0297;
    65: op1_15_in19 = reg_0231;
    66: op1_15_in19 = reg_0301;
    67: op1_15_in19 = reg_0479;
    68: op1_15_in19 = imem03_in[19:16];
    69: op1_15_in19 = imem06_in[115:112];
    70: op1_15_in19 = reg_0397;
    71: op1_15_in19 = reg_0302;
    73: op1_15_in19 = reg_0763;
    76: op1_15_in19 = reg_0656;
    77: op1_15_in19 = reg_0065;
    78: op1_15_in19 = reg_0616;
    79: op1_15_in19 = imem07_in[91:88];
    80: op1_15_in19 = reg_0714;
    81: op1_15_in19 = reg_0396;
    82: op1_15_in19 = reg_0669;
    83: op1_15_in19 = reg_0487;
    84: op1_15_in19 = imem06_in[39:36];
    85: op1_15_in19 = reg_0795;
    86: op1_15_in19 = reg_0345;
    87: op1_15_in19 = imem06_in[71:68];
    88: op1_15_in19 = reg_0591;
    89: op1_15_in19 = reg_0614;
    90: op1_15_in19 = reg_0062;
    91: op1_15_in19 = imem01_in[103:100];
    92: op1_15_in19 = reg_0467;
    93: op1_15_in19 = reg_0421;
    default: op1_15_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv19 = 1;
    7: op1_15_inv19 = 1;
    9: op1_15_inv19 = 1;
    10: op1_15_inv19 = 1;
    11: op1_15_inv19 = 1;
    12: op1_15_inv19 = 1;
    15: op1_15_inv19 = 1;
    17: op1_15_inv19 = 1;
    20: op1_15_inv19 = 1;
    21: op1_15_inv19 = 1;
    23: op1_15_inv19 = 1;
    26: op1_15_inv19 = 1;
    27: op1_15_inv19 = 1;
    29: op1_15_inv19 = 1;
    33: op1_15_inv19 = 1;
    34: op1_15_inv19 = 1;
    35: op1_15_inv19 = 1;
    37: op1_15_inv19 = 1;
    38: op1_15_inv19 = 1;
    39: op1_15_inv19 = 1;
    41: op1_15_inv19 = 1;
    44: op1_15_inv19 = 1;
    45: op1_15_inv19 = 1;
    49: op1_15_inv19 = 1;
    52: op1_15_inv19 = 1;
    53: op1_15_inv19 = 1;
    55: op1_15_inv19 = 1;
    56: op1_15_inv19 = 1;
    57: op1_15_inv19 = 1;
    59: op1_15_inv19 = 1;
    61: op1_15_inv19 = 1;
    62: op1_15_inv19 = 1;
    63: op1_15_inv19 = 1;
    64: op1_15_inv19 = 1;
    66: op1_15_inv19 = 1;
    69: op1_15_inv19 = 1;
    71: op1_15_inv19 = 1;
    73: op1_15_inv19 = 1;
    76: op1_15_inv19 = 1;
    79: op1_15_inv19 = 1;
    80: op1_15_inv19 = 1;
    85: op1_15_inv19 = 1;
    86: op1_15_inv19 = 1;
    90: op1_15_inv19 = 1;
    91: op1_15_inv19 = 1;
    92: op1_15_inv19 = 1;
    default: op1_15_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の20番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in20 = reg_0589;
    6: op1_15_in20 = reg_0013;
    7: op1_15_in20 = imem06_in[43:40];
    84: op1_15_in20 = imem06_in[43:40];
    8: op1_15_in20 = reg_0503;
    71: op1_15_in20 = reg_0503;
    9: op1_15_in20 = reg_0190;
    10: op1_15_in20 = reg_0796;
    11: op1_15_in20 = reg_0035;
    12: op1_15_in20 = reg_0531;
    13: op1_15_in20 = reg_0033;
    15: op1_15_in20 = reg_0095;
    16: op1_15_in20 = reg_0541;
    17: op1_15_in20 = reg_0385;
    18: op1_15_in20 = imem04_in[67:64];
    19: op1_15_in20 = reg_0658;
    20: op1_15_in20 = reg_0224;
    21: op1_15_in20 = reg_0162;
    22: op1_15_in20 = reg_0007;
    23: op1_15_in20 = reg_0198;
    46: op1_15_in20 = reg_0198;
    24: op1_15_in20 = imem02_in[83:80];
    25: op1_15_in20 = imem07_in[3:0];
    26: op1_15_in20 = reg_0572;
    27: op1_15_in20 = reg_0141;
    29: op1_15_in20 = reg_0342;
    86: op1_15_in20 = reg_0342;
    30: op1_15_in20 = reg_0620;
    31: op1_15_in20 = reg_0721;
    33: op1_15_in20 = reg_0490;
    34: op1_15_in20 = reg_0084;
    35: op1_15_in20 = imem06_in[35:32];
    37: op1_15_in20 = reg_0179;
    38: op1_15_in20 = imem01_in[51:48];
    39: op1_15_in20 = reg_0241;
    40: op1_15_in20 = reg_0553;
    41: op1_15_in20 = imem07_in[71:68];
    43: op1_15_in20 = reg_0248;
    44: op1_15_in20 = imem04_in[123:120];
    45: op1_15_in20 = reg_0239;
    47: op1_15_in20 = reg_0537;
    48: op1_15_in20 = reg_0795;
    49: op1_15_in20 = reg_0811;
    50: op1_15_in20 = reg_0117;
    83: op1_15_in20 = reg_0117;
    51: op1_15_in20 = reg_0820;
    52: op1_15_in20 = reg_0356;
    53: op1_15_in20 = reg_0362;
    54: op1_15_in20 = reg_0585;
    55: op1_15_in20 = reg_0624;
    56: op1_15_in20 = imem06_in[31:28];
    57: op1_15_in20 = reg_0087;
    59: op1_15_in20 = reg_0814;
    61: op1_15_in20 = reg_0423;
    62: op1_15_in20 = reg_0006;
    63: op1_15_in20 = imem04_in[115:112];
    64: op1_15_in20 = reg_0292;
    65: op1_15_in20 = reg_0039;
    66: op1_15_in20 = reg_0062;
    67: op1_15_in20 = reg_0214;
    68: op1_15_in20 = imem03_in[23:20];
    69: op1_15_in20 = reg_0817;
    70: op1_15_in20 = reg_0225;
    72: op1_15_in20 = imem05_in[39:36];
    73: op1_15_in20 = reg_0608;
    76: op1_15_in20 = reg_0753;
    77: op1_15_in20 = imem05_in[23:20];
    78: op1_15_in20 = reg_0050;
    79: op1_15_in20 = imem07_in[107:104];
    80: op1_15_in20 = reg_0729;
    81: op1_15_in20 = reg_0557;
    82: op1_15_in20 = reg_0601;
    85: op1_15_in20 = reg_0550;
    87: op1_15_in20 = imem06_in[103:100];
    88: op1_15_in20 = reg_0493;
    89: op1_15_in20 = reg_0679;
    90: op1_15_in20 = imem05_in[47:44];
    91: op1_15_in20 = imem01_in[119:116];
    92: op1_15_in20 = reg_0470;
    93: op1_15_in20 = reg_0098;
    default: op1_15_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv20 = 1;
    10: op1_15_inv20 = 1;
    16: op1_15_inv20 = 1;
    17: op1_15_inv20 = 1;
    19: op1_15_inv20 = 1;
    20: op1_15_inv20 = 1;
    24: op1_15_inv20 = 1;
    25: op1_15_inv20 = 1;
    26: op1_15_inv20 = 1;
    27: op1_15_inv20 = 1;
    30: op1_15_inv20 = 1;
    31: op1_15_inv20 = 1;
    33: op1_15_inv20 = 1;
    34: op1_15_inv20 = 1;
    37: op1_15_inv20 = 1;
    39: op1_15_inv20 = 1;
    40: op1_15_inv20 = 1;
    41: op1_15_inv20 = 1;
    43: op1_15_inv20 = 1;
    45: op1_15_inv20 = 1;
    47: op1_15_inv20 = 1;
    49: op1_15_inv20 = 1;
    50: op1_15_inv20 = 1;
    52: op1_15_inv20 = 1;
    54: op1_15_inv20 = 1;
    55: op1_15_inv20 = 1;
    56: op1_15_inv20 = 1;
    57: op1_15_inv20 = 1;
    61: op1_15_inv20 = 1;
    62: op1_15_inv20 = 1;
    63: op1_15_inv20 = 1;
    64: op1_15_inv20 = 1;
    66: op1_15_inv20 = 1;
    67: op1_15_inv20 = 1;
    68: op1_15_inv20 = 1;
    71: op1_15_inv20 = 1;
    73: op1_15_inv20 = 1;
    77: op1_15_inv20 = 1;
    79: op1_15_inv20 = 1;
    80: op1_15_inv20 = 1;
    82: op1_15_inv20 = 1;
    83: op1_15_inv20 = 1;
    85: op1_15_inv20 = 1;
    88: op1_15_inv20 = 1;
    89: op1_15_inv20 = 1;
    92: op1_15_inv20 = 1;
    default: op1_15_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の21番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in21 = reg_0576;
    6: op1_15_in21 = reg_0801;
    7: op1_15_in21 = imem06_in[91:88];
    8: op1_15_in21 = reg_0515;
    54: op1_15_in21 = reg_0515;
    9: op1_15_in21 = reg_0195;
    10: op1_15_in21 = reg_0797;
    11: op1_15_in21 = reg_0037;
    12: op1_15_in21 = reg_0547;
    13: op1_15_in21 = reg_0813;
    15: op1_15_in21 = reg_0085;
    16: op1_15_in21 = reg_0305;
    17: op1_15_in21 = reg_0396;
    18: op1_15_in21 = reg_0068;
    19: op1_15_in21 = reg_0637;
    20: op1_15_in21 = reg_0277;
    21: op1_15_in21 = reg_0170;
    80: op1_15_in21 = reg_0170;
    22: op1_15_in21 = reg_0004;
    23: op1_15_in21 = reg_0190;
    24: op1_15_in21 = imem02_in[87:84];
    25: op1_15_in21 = imem07_in[39:36];
    26: op1_15_in21 = reg_0592;
    27: op1_15_in21 = reg_0155;
    29: op1_15_in21 = reg_0355;
    30: op1_15_in21 = reg_0626;
    78: op1_15_in21 = reg_0626;
    31: op1_15_in21 = reg_0726;
    33: op1_15_in21 = reg_0785;
    34: op1_15_in21 = reg_0272;
    35: op1_15_in21 = imem06_in[47:44];
    84: op1_15_in21 = imem06_in[47:44];
    37: op1_15_in21 = reg_0161;
    38: op1_15_in21 = imem01_in[115:112];
    39: op1_15_in21 = reg_0248;
    40: op1_15_in21 = reg_0537;
    41: op1_15_in21 = imem07_in[119:116];
    43: op1_15_in21 = reg_0122;
    44: op1_15_in21 = reg_0328;
    45: op1_15_in21 = reg_0444;
    46: op1_15_in21 = reg_0205;
    47: op1_15_in21 = reg_0088;
    48: op1_15_in21 = reg_0793;
    49: op1_15_in21 = reg_0002;
    50: op1_15_in21 = reg_0110;
    51: op1_15_in21 = reg_0563;
    52: op1_15_in21 = reg_0363;
    53: op1_15_in21 = reg_0565;
    55: op1_15_in21 = reg_0298;
    56: op1_15_in21 = imem06_in[39:36];
    57: op1_15_in21 = reg_0056;
    59: op1_15_in21 = reg_0628;
    61: op1_15_in21 = reg_0574;
    62: op1_15_in21 = reg_0013;
    63: op1_15_in21 = reg_0316;
    64: op1_15_in21 = reg_0508;
    65: op1_15_in21 = imem05_in[11:8];
    66: op1_15_in21 = reg_0065;
    67: op1_15_in21 = reg_0200;
    68: op1_15_in21 = imem03_in[35:32];
    69: op1_15_in21 = reg_0814;
    70: op1_15_in21 = reg_0232;
    71: op1_15_in21 = reg_0629;
    72: op1_15_in21 = imem05_in[51:48];
    73: op1_15_in21 = reg_0663;
    76: op1_15_in21 = reg_0655;
    77: op1_15_in21 = imem05_in[99:96];
    79: op1_15_in21 = imem07_in[111:108];
    81: op1_15_in21 = reg_0001;
    82: op1_15_in21 = reg_0678;
    83: op1_15_in21 = imem02_in[7:4];
    85: op1_15_in21 = reg_0113;
    86: op1_15_in21 = reg_0406;
    87: op1_15_in21 = imem06_in[123:120];
    88: op1_15_in21 = reg_0009;
    89: op1_15_in21 = reg_0622;
    90: op1_15_in21 = imem05_in[111:108];
    91: op1_15_in21 = reg_0497;
    92: op1_15_in21 = reg_0479;
    93: op1_15_in21 = reg_0741;
    default: op1_15_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    8: op1_15_inv21 = 1;
    9: op1_15_inv21 = 1;
    13: op1_15_inv21 = 1;
    17: op1_15_inv21 = 1;
    18: op1_15_inv21 = 1;
    20: op1_15_inv21 = 1;
    22: op1_15_inv21 = 1;
    23: op1_15_inv21 = 1;
    24: op1_15_inv21 = 1;
    26: op1_15_inv21 = 1;
    27: op1_15_inv21 = 1;
    29: op1_15_inv21 = 1;
    31: op1_15_inv21 = 1;
    35: op1_15_inv21 = 1;
    38: op1_15_inv21 = 1;
    40: op1_15_inv21 = 1;
    41: op1_15_inv21 = 1;
    43: op1_15_inv21 = 1;
    45: op1_15_inv21 = 1;
    46: op1_15_inv21 = 1;
    47: op1_15_inv21 = 1;
    49: op1_15_inv21 = 1;
    54: op1_15_inv21 = 1;
    55: op1_15_inv21 = 1;
    57: op1_15_inv21 = 1;
    59: op1_15_inv21 = 1;
    65: op1_15_inv21 = 1;
    66: op1_15_inv21 = 1;
    67: op1_15_inv21 = 1;
    72: op1_15_inv21 = 1;
    76: op1_15_inv21 = 1;
    78: op1_15_inv21 = 1;
    81: op1_15_inv21 = 1;
    83: op1_15_inv21 = 1;
    86: op1_15_inv21 = 1;
    89: op1_15_inv21 = 1;
    91: op1_15_inv21 = 1;
    default: op1_15_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の22番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in22 = reg_0384;
    6: op1_15_in22 = reg_0016;
    7: op1_15_in22 = imem06_in[95:92];
    8: op1_15_in22 = reg_0232;
    9: op1_15_in22 = reg_0229;
    10: op1_15_in22 = reg_0491;
    11: op1_15_in22 = reg_0029;
    12: op1_15_in22 = reg_0292;
    13: op1_15_in22 = reg_0034;
    15: op1_15_in22 = reg_0052;
    16: op1_15_in22 = reg_0300;
    17: op1_15_in22 = reg_0309;
    18: op1_15_in22 = reg_0077;
    19: op1_15_in22 = reg_0646;
    20: op1_15_in22 = reg_0145;
    22: op1_15_in22 = imem04_in[59:56];
    23: op1_15_in22 = reg_0206;
    24: op1_15_in22 = imem02_in[115:112];
    25: op1_15_in22 = reg_0730;
    26: op1_15_in22 = reg_0591;
    27: op1_15_in22 = imem06_in[27:24];
    29: op1_15_in22 = reg_0350;
    30: op1_15_in22 = reg_0633;
    31: op1_15_in22 = reg_0715;
    33: op1_15_in22 = reg_0736;
    34: op1_15_in22 = reg_0285;
    35: op1_15_in22 = imem06_in[111:108];
    37: op1_15_in22 = reg_0168;
    38: op1_15_in22 = reg_0758;
    39: op1_15_in22 = reg_0508;
    40: op1_15_in22 = reg_0055;
    57: op1_15_in22 = reg_0055;
    41: op1_15_in22 = imem07_in[127:124];
    79: op1_15_in22 = imem07_in[127:124];
    43: op1_15_in22 = reg_0099;
    44: op1_15_in22 = reg_0542;
    45: op1_15_in22 = reg_0268;
    46: op1_15_in22 = reg_0192;
    47: op1_15_in22 = reg_0058;
    48: op1_15_in22 = reg_0782;
    49: op1_15_in22 = reg_0808;
    50: op1_15_in22 = imem02_in[51:48];
    51: op1_15_in22 = reg_0225;
    52: op1_15_in22 = reg_0096;
    53: op1_15_in22 = reg_0360;
    54: op1_15_in22 = reg_0643;
    55: op1_15_in22 = reg_0619;
    56: op1_15_in22 = imem06_in[47:44];
    59: op1_15_in22 = reg_0369;
    61: op1_15_in22 = reg_0240;
    62: op1_15_in22 = reg_0807;
    63: op1_15_in22 = reg_0553;
    64: op1_15_in22 = reg_0062;
    65: op1_15_in22 = imem05_in[55:52];
    66: op1_15_in22 = reg_0598;
    67: op1_15_in22 = reg_0193;
    68: op1_15_in22 = imem03_in[47:44];
    69: op1_15_in22 = reg_0606;
    70: op1_15_in22 = reg_0054;
    71: op1_15_in22 = reg_0627;
    72: op1_15_in22 = imem05_in[67:64];
    73: op1_15_in22 = reg_0813;
    76: op1_15_in22 = reg_0344;
    77: op1_15_in22 = imem05_in[115:112];
    78: op1_15_in22 = reg_0065;
    80: op1_15_in22 = reg_0091;
    81: op1_15_in22 = reg_0803;
    82: op1_15_in22 = imem02_in[43:40];
    83: op1_15_in22 = imem02_in[59:56];
    84: op1_15_in22 = imem06_in[115:112];
    85: op1_15_in22 = reg_0027;
    86: op1_15_in22 = reg_0514;
    87: op1_15_in22 = reg_0348;
    88: op1_15_in22 = reg_0507;
    89: op1_15_in22 = reg_0780;
    90: op1_15_in22 = reg_0326;
    91: op1_15_in22 = reg_0668;
    92: op1_15_in22 = reg_0459;
    93: op1_15_in22 = reg_0761;
    default: op1_15_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv22 = 1;
    9: op1_15_inv22 = 1;
    10: op1_15_inv22 = 1;
    13: op1_15_inv22 = 1;
    15: op1_15_inv22 = 1;
    18: op1_15_inv22 = 1;
    19: op1_15_inv22 = 1;
    22: op1_15_inv22 = 1;
    23: op1_15_inv22 = 1;
    24: op1_15_inv22 = 1;
    29: op1_15_inv22 = 1;
    33: op1_15_inv22 = 1;
    41: op1_15_inv22 = 1;
    44: op1_15_inv22 = 1;
    45: op1_15_inv22 = 1;
    47: op1_15_inv22 = 1;
    49: op1_15_inv22 = 1;
    54: op1_15_inv22 = 1;
    55: op1_15_inv22 = 1;
    57: op1_15_inv22 = 1;
    61: op1_15_inv22 = 1;
    62: op1_15_inv22 = 1;
    63: op1_15_inv22 = 1;
    64: op1_15_inv22 = 1;
    67: op1_15_inv22 = 1;
    68: op1_15_inv22 = 1;
    69: op1_15_inv22 = 1;
    72: op1_15_inv22 = 1;
    76: op1_15_inv22 = 1;
    77: op1_15_inv22 = 1;
    78: op1_15_inv22 = 1;
    81: op1_15_inv22 = 1;
    84: op1_15_inv22 = 1;
    86: op1_15_inv22 = 1;
    87: op1_15_inv22 = 1;
    88: op1_15_inv22 = 1;
    93: op1_15_inv22 = 1;
    default: op1_15_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の23番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in23 = reg_0343;
    6: op1_15_in23 = reg_0010;
    7: op1_15_in23 = reg_0628;
    8: op1_15_in23 = reg_0235;
    9: op1_15_in23 = reg_0496;
    10: op1_15_in23 = reg_0794;
    11: op1_15_in23 = reg_0752;
    12: op1_15_in23 = reg_0047;
    13: op1_15_in23 = reg_0750;
    15: op1_15_in23 = reg_0086;
    16: op1_15_in23 = reg_0289;
    17: op1_15_in23 = reg_0389;
    18: op1_15_in23 = imem05_in[79:76];
    19: op1_15_in23 = reg_0657;
    20: op1_15_in23 = reg_0152;
    22: op1_15_in23 = imem04_in[63:60];
    23: op1_15_in23 = reg_0199;
    24: op1_15_in23 = reg_0650;
    25: op1_15_in23 = reg_0721;
    26: op1_15_in23 = reg_0581;
    27: op1_15_in23 = imem06_in[103:100];
    29: op1_15_in23 = reg_0540;
    30: op1_15_in23 = reg_0618;
    31: op1_15_in23 = reg_0707;
    33: op1_15_in23 = reg_0279;
    34: op1_15_in23 = reg_0129;
    35: op1_15_in23 = imem06_in[123:120];
    37: op1_15_in23 = reg_0184;
    38: op1_15_in23 = reg_0337;
    39: op1_15_in23 = reg_0758;
    40: op1_15_in23 = reg_0555;
    57: op1_15_in23 = reg_0555;
    41: op1_15_in23 = reg_0702;
    43: op1_15_in23 = reg_0106;
    44: op1_15_in23 = reg_0537;
    45: op1_15_in23 = reg_0167;
    46: op1_15_in23 = imem01_in[19:16];
    47: op1_15_in23 = reg_0280;
    48: op1_15_in23 = reg_0786;
    49: op1_15_in23 = reg_0003;
    50: op1_15_in23 = imem02_in[75:72];
    51: op1_15_in23 = reg_0241;
    52: op1_15_in23 = reg_0094;
    53: op1_15_in23 = reg_0353;
    54: op1_15_in23 = reg_0069;
    55: op1_15_in23 = reg_0408;
    56: op1_15_in23 = imem06_in[59:56];
    59: op1_15_in23 = reg_0659;
    61: op1_15_in23 = reg_0419;
    62: op1_15_in23 = reg_0004;
    63: op1_15_in23 = reg_0071;
    64: op1_15_in23 = reg_0259;
    66: op1_15_in23 = reg_0259;
    65: op1_15_in23 = imem05_in[59:56];
    67: op1_15_in23 = reg_0190;
    68: op1_15_in23 = imem03_in[111:108];
    69: op1_15_in23 = reg_0619;
    70: op1_15_in23 = reg_0217;
    71: op1_15_in23 = reg_0610;
    72: op1_15_in23 = reg_0288;
    73: op1_15_in23 = reg_0501;
    76: op1_15_in23 = reg_0358;
    77: op1_15_in23 = reg_0736;
    78: op1_15_in23 = reg_0068;
    79: op1_15_in23 = reg_0722;
    80: op1_15_in23 = reg_0132;
    81: op1_15_in23 = reg_0804;
    82: op1_15_in23 = imem02_in[67:64];
    83: op1_15_in23 = imem02_in[95:92];
    84: op1_15_in23 = reg_0346;
    85: op1_15_in23 = reg_0134;
    86: op1_15_in23 = reg_0092;
    87: op1_15_in23 = reg_0817;
    88: op1_15_in23 = reg_0571;
    89: op1_15_in23 = reg_0771;
    90: op1_15_in23 = reg_0500;
    91: op1_15_in23 = reg_0385;
    92: op1_15_in23 = reg_0207;
    93: op1_15_in23 = reg_0114;
    default: op1_15_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv23 = 1;
    6: op1_15_inv23 = 1;
    10: op1_15_inv23 = 1;
    12: op1_15_inv23 = 1;
    13: op1_15_inv23 = 1;
    15: op1_15_inv23 = 1;
    20: op1_15_inv23 = 1;
    22: op1_15_inv23 = 1;
    23: op1_15_inv23 = 1;
    25: op1_15_inv23 = 1;
    29: op1_15_inv23 = 1;
    30: op1_15_inv23 = 1;
    31: op1_15_inv23 = 1;
    33: op1_15_inv23 = 1;
    35: op1_15_inv23 = 1;
    39: op1_15_inv23 = 1;
    40: op1_15_inv23 = 1;
    43: op1_15_inv23 = 1;
    44: op1_15_inv23 = 1;
    51: op1_15_inv23 = 1;
    53: op1_15_inv23 = 1;
    54: op1_15_inv23 = 1;
    55: op1_15_inv23 = 1;
    57: op1_15_inv23 = 1;
    59: op1_15_inv23 = 1;
    61: op1_15_inv23 = 1;
    62: op1_15_inv23 = 1;
    63: op1_15_inv23 = 1;
    66: op1_15_inv23 = 1;
    67: op1_15_inv23 = 1;
    69: op1_15_inv23 = 1;
    71: op1_15_inv23 = 1;
    72: op1_15_inv23 = 1;
    73: op1_15_inv23 = 1;
    76: op1_15_inv23 = 1;
    77: op1_15_inv23 = 1;
    82: op1_15_inv23 = 1;
    83: op1_15_inv23 = 1;
    86: op1_15_inv23 = 1;
    91: op1_15_inv23 = 1;
    default: op1_15_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の24番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in24 = reg_0369;
    6: op1_15_in24 = imem04_in[35:32];
    7: op1_15_in24 = reg_0577;
    8: op1_15_in24 = reg_0246;
    9: op1_15_in24 = reg_0500;
    10: op1_15_in24 = reg_0790;
    11: op1_15_in24 = imem07_in[23:20];
    12: op1_15_in24 = reg_0058;
    13: op1_15_in24 = imem07_in[31:28];
    15: op1_15_in24 = reg_0051;
    16: op1_15_in24 = reg_0297;
    47: op1_15_in24 = reg_0297;
    17: op1_15_in24 = reg_0000;
    18: op1_15_in24 = imem05_in[83:80];
    19: op1_15_in24 = reg_0661;
    20: op1_15_in24 = reg_0142;
    22: op1_15_in24 = imem04_in[71:68];
    23: op1_15_in24 = reg_0197;
    24: op1_15_in24 = reg_0666;
    25: op1_15_in24 = reg_0717;
    26: op1_15_in24 = reg_0595;
    27: op1_15_in24 = imem06_in[107:104];
    29: op1_15_in24 = reg_0094;
    30: op1_15_in24 = reg_0370;
    87: op1_15_in24 = reg_0370;
    31: op1_15_in24 = reg_0706;
    33: op1_15_in24 = reg_0089;
    34: op1_15_in24 = reg_0141;
    35: op1_15_in24 = reg_0408;
    38: op1_15_in24 = reg_0519;
    39: op1_15_in24 = reg_0497;
    40: op1_15_in24 = reg_0060;
    57: op1_15_in24 = reg_0060;
    41: op1_15_in24 = reg_0729;
    43: op1_15_in24 = reg_0127;
    44: op1_15_in24 = reg_0088;
    45: op1_15_in24 = reg_0182;
    46: op1_15_in24 = imem01_in[31:28];
    48: op1_15_in24 = reg_0784;
    49: op1_15_in24 = reg_0007;
    50: op1_15_in24 = imem02_in[83:80];
    51: op1_15_in24 = reg_0422;
    52: op1_15_in24 = imem03_in[3:0];
    53: op1_15_in24 = reg_0743;
    86: op1_15_in24 = reg_0743;
    54: op1_15_in24 = reg_0275;
    55: op1_15_in24 = reg_0775;
    59: op1_15_in24 = reg_0775;
    56: op1_15_in24 = imem06_in[71:68];
    61: op1_15_in24 = reg_0104;
    62: op1_15_in24 = imem04_in[3:0];
    63: op1_15_in24 = reg_0292;
    64: op1_15_in24 = reg_0075;
    65: op1_15_in24 = imem05_in[79:76];
    66: op1_15_in24 = reg_0776;
    67: op1_15_in24 = reg_0195;
    68: op1_15_in24 = reg_0604;
    69: op1_15_in24 = reg_0354;
    70: op1_15_in24 = reg_0105;
    71: op1_15_in24 = reg_0223;
    72: op1_15_in24 = reg_0257;
    73: op1_15_in24 = imem07_in[11:8];
    76: op1_15_in24 = reg_0353;
    77: op1_15_in24 = reg_0227;
    78: op1_15_in24 = reg_0513;
    79: op1_15_in24 = reg_0726;
    80: op1_15_in24 = reg_0099;
    81: op1_15_in24 = reg_0809;
    82: op1_15_in24 = imem02_in[71:68];
    83: op1_15_in24 = reg_0356;
    84: op1_15_in24 = reg_0762;
    85: op1_15_in24 = reg_0517;
    88: op1_15_in24 = reg_0564;
    89: op1_15_in24 = reg_0233;
    90: op1_15_in24 = reg_0583;
    91: op1_15_in24 = reg_0102;
    92: op1_15_in24 = reg_0194;
    93: op1_15_in24 = reg_0234;
    default: op1_15_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv24 = 1;
    6: op1_15_inv24 = 1;
    7: op1_15_inv24 = 1;
    8: op1_15_inv24 = 1;
    9: op1_15_inv24 = 1;
    11: op1_15_inv24 = 1;
    12: op1_15_inv24 = 1;
    13: op1_15_inv24 = 1;
    17: op1_15_inv24 = 1;
    19: op1_15_inv24 = 1;
    23: op1_15_inv24 = 1;
    26: op1_15_inv24 = 1;
    27: op1_15_inv24 = 1;
    29: op1_15_inv24 = 1;
    30: op1_15_inv24 = 1;
    38: op1_15_inv24 = 1;
    40: op1_15_inv24 = 1;
    44: op1_15_inv24 = 1;
    48: op1_15_inv24 = 1;
    51: op1_15_inv24 = 1;
    52: op1_15_inv24 = 1;
    53: op1_15_inv24 = 1;
    59: op1_15_inv24 = 1;
    62: op1_15_inv24 = 1;
    65: op1_15_inv24 = 1;
    66: op1_15_inv24 = 1;
    67: op1_15_inv24 = 1;
    68: op1_15_inv24 = 1;
    70: op1_15_inv24 = 1;
    76: op1_15_inv24 = 1;
    79: op1_15_inv24 = 1;
    81: op1_15_inv24 = 1;
    82: op1_15_inv24 = 1;
    83: op1_15_inv24 = 1;
    84: op1_15_inv24 = 1;
    87: op1_15_inv24 = 1;
    88: op1_15_inv24 = 1;
    89: op1_15_inv24 = 1;
    90: op1_15_inv24 = 1;
    92: op1_15_inv24 = 1;
    93: op1_15_inv24 = 1;
    default: op1_15_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の25番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in25 = reg_0385;
    6: op1_15_in25 = imem04_in[43:40];
    7: op1_15_in25 = reg_0622;
    8: op1_15_in25 = reg_0239;
    9: op1_15_in25 = reg_0740;
    10: op1_15_in25 = reg_0267;
    11: op1_15_in25 = imem07_in[55:52];
    12: op1_15_in25 = reg_0066;
    13: op1_15_in25 = imem07_in[71:68];
    15: op1_15_in25 = reg_0084;
    16: op1_15_in25 = reg_0076;
    17: op1_15_in25 = reg_0053;
    18: op1_15_in25 = imem05_in[123:120];
    19: op1_15_in25 = reg_0649;
    20: op1_15_in25 = reg_0138;
    22: op1_15_in25 = imem04_in[115:112];
    23: op1_15_in25 = imem01_in[15:12];
    24: op1_15_in25 = reg_0654;
    25: op1_15_in25 = reg_0703;
    26: op1_15_in25 = reg_0590;
    76: op1_15_in25 = reg_0590;
    27: op1_15_in25 = imem06_in[111:108];
    29: op1_15_in25 = imem03_in[31:28];
    30: op1_15_in25 = reg_0407;
    31: op1_15_in25 = reg_0433;
    33: op1_15_in25 = reg_0128;
    34: op1_15_in25 = reg_0140;
    35: op1_15_in25 = reg_0370;
    38: op1_15_in25 = reg_0333;
    39: op1_15_in25 = reg_0563;
    40: op1_15_in25 = reg_0558;
    41: op1_15_in25 = reg_0708;
    43: op1_15_in25 = reg_0117;
    44: op1_15_in25 = reg_0055;
    45: op1_15_in25 = reg_0166;
    46: op1_15_in25 = imem01_in[67:64];
    47: op1_15_in25 = reg_0617;
    48: op1_15_in25 = reg_0787;
    49: op1_15_in25 = reg_0801;
    50: op1_15_in25 = reg_0337;
    51: op1_15_in25 = reg_0574;
    52: op1_15_in25 = imem03_in[51:48];
    53: op1_15_in25 = reg_0081;
    54: op1_15_in25 = imem05_in[7:4];
    55: op1_15_in25 = reg_0231;
    56: op1_15_in25 = imem06_in[87:84];
    57: op1_15_in25 = reg_0554;
    59: op1_15_in25 = reg_0821;
    61: op1_15_in25 = imem02_in[39:36];
    62: op1_15_in25 = imem04_in[11:8];
    63: op1_15_in25 = reg_0679;
    64: op1_15_in25 = reg_0099;
    65: op1_15_in25 = imem05_in[107:104];
    66: op1_15_in25 = imem05_in[83:80];
    67: op1_15_in25 = imem01_in[7:4];
    68: op1_15_in25 = reg_0319;
    69: op1_15_in25 = reg_0404;
    70: op1_15_in25 = reg_0592;
    71: op1_15_in25 = reg_0069;
    72: op1_15_in25 = reg_0236;
    73: op1_15_in25 = imem07_in[31:28];
    77: op1_15_in25 = reg_0666;
    78: op1_15_in25 = reg_0136;
    79: op1_15_in25 = reg_0158;
    80: op1_15_in25 = reg_0710;
    81: op1_15_in25 = imem04_in[3:0];
    82: op1_15_in25 = imem02_in[103:100];
    83: op1_15_in25 = reg_0363;
    84: op1_15_in25 = reg_0817;
    85: op1_15_in25 = reg_0309;
    86: op1_15_in25 = reg_0526;
    87: op1_15_in25 = reg_0618;
    88: op1_15_in25 = reg_0368;
    89: op1_15_in25 = reg_0416;
    90: op1_15_in25 = reg_0149;
    91: op1_15_in25 = reg_0388;
    92: op1_15_in25 = reg_0201;
    93: op1_15_in25 = imem01_in[11:8];
    default: op1_15_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv25 = 1;
    8: op1_15_inv25 = 1;
    10: op1_15_inv25 = 1;
    12: op1_15_inv25 = 1;
    18: op1_15_inv25 = 1;
    20: op1_15_inv25 = 1;
    24: op1_15_inv25 = 1;
    25: op1_15_inv25 = 1;
    26: op1_15_inv25 = 1;
    31: op1_15_inv25 = 1;
    33: op1_15_inv25 = 1;
    35: op1_15_inv25 = 1;
    38: op1_15_inv25 = 1;
    41: op1_15_inv25 = 1;
    43: op1_15_inv25 = 1;
    44: op1_15_inv25 = 1;
    45: op1_15_inv25 = 1;
    47: op1_15_inv25 = 1;
    49: op1_15_inv25 = 1;
    50: op1_15_inv25 = 1;
    51: op1_15_inv25 = 1;
    54: op1_15_inv25 = 1;
    55: op1_15_inv25 = 1;
    57: op1_15_inv25 = 1;
    59: op1_15_inv25 = 1;
    62: op1_15_inv25 = 1;
    69: op1_15_inv25 = 1;
    70: op1_15_inv25 = 1;
    72: op1_15_inv25 = 1;
    77: op1_15_inv25 = 1;
    81: op1_15_inv25 = 1;
    82: op1_15_inv25 = 1;
    83: op1_15_inv25 = 1;
    84: op1_15_inv25 = 1;
    85: op1_15_inv25 = 1;
    86: op1_15_inv25 = 1;
    88: op1_15_inv25 = 1;
    91: op1_15_inv25 = 1;
    92: op1_15_inv25 = 1;
    default: op1_15_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の26番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in26 = reg_0006;
    6: op1_15_in26 = imem04_in[51:48];
    7: op1_15_in26 = reg_0372;
    88: op1_15_in26 = reg_0372;
    8: op1_15_in26 = reg_0242;
    9: op1_15_in26 = reg_0523;
    10: op1_15_in26 = reg_0262;
    11: op1_15_in26 = imem07_in[59:56];
    12: op1_15_in26 = imem05_in[7:4];
    89: op1_15_in26 = imem05_in[7:4];
    13: op1_15_in26 = imem07_in[111:108];
    15: op1_15_in26 = reg_0094;
    16: op1_15_in26 = reg_0068;
    17: op1_15_in26 = reg_0059;
    18: op1_15_in26 = reg_0488;
    19: op1_15_in26 = reg_0663;
    20: op1_15_in26 = reg_0153;
    22: op1_15_in26 = reg_0316;
    23: op1_15_in26 = reg_0513;
    24: op1_15_in26 = reg_0639;
    50: op1_15_in26 = reg_0639;
    25: op1_15_in26 = reg_0712;
    26: op1_15_in26 = reg_0387;
    27: op1_15_in26 = imem06_in[127:124];
    29: op1_15_in26 = imem03_in[55:52];
    30: op1_15_in26 = reg_0405;
    31: op1_15_in26 = reg_0420;
    33: op1_15_in26 = reg_0139;
    34: op1_15_in26 = imem06_in[15:12];
    35: op1_15_in26 = reg_0821;
    38: op1_15_in26 = reg_0487;
    39: op1_15_in26 = reg_0825;
    40: op1_15_in26 = reg_0058;
    41: op1_15_in26 = reg_0709;
    43: op1_15_in26 = imem02_in[7:4];
    44: op1_15_in26 = reg_0556;
    45: op1_15_in26 = reg_0157;
    46: op1_15_in26 = imem01_in[75:72];
    47: op1_15_in26 = reg_0512;
    48: op1_15_in26 = reg_0304;
    49: op1_15_in26 = imem04_in[19:16];
    62: op1_15_in26 = imem04_in[19:16];
    51: op1_15_in26 = reg_0054;
    52: op1_15_in26 = imem03_in[83:80];
    53: op1_15_in26 = reg_0757;
    54: op1_15_in26 = imem05_in[11:8];
    55: op1_15_in26 = reg_0238;
    56: op1_15_in26 = imem06_in[107:104];
    57: op1_15_in26 = reg_0283;
    59: op1_15_in26 = reg_0375;
    61: op1_15_in26 = imem02_in[43:40];
    63: op1_15_in26 = reg_0223;
    64: op1_15_in26 = reg_0040;
    65: op1_15_in26 = reg_0132;
    66: op1_15_in26 = imem05_in[95:92];
    67: op1_15_in26 = imem01_in[39:36];
    68: op1_15_in26 = reg_0329;
    69: op1_15_in26 = reg_0031;
    70: op1_15_in26 = imem02_in[19:16];
    71: op1_15_in26 = reg_0259;
    72: op1_15_in26 = reg_0148;
    73: op1_15_in26 = imem07_in[55:52];
    76: op1_15_in26 = reg_0080;
    77: op1_15_in26 = reg_0128;
    78: op1_15_in26 = reg_0797;
    79: op1_15_in26 = reg_0711;
    80: op1_15_in26 = reg_0162;
    81: op1_15_in26 = imem04_in[7:4];
    82: op1_15_in26 = imem02_in[119:116];
    83: op1_15_in26 = reg_0594;
    84: op1_15_in26 = reg_0619;
    85: op1_15_in26 = reg_0720;
    86: op1_15_in26 = imem03_in[23:20];
    87: op1_15_in26 = reg_0032;
    90: op1_15_in26 = reg_0827;
    91: op1_15_in26 = reg_0235;
    92: op1_15_in26 = reg_0421;
    93: op1_15_in26 = imem01_in[71:68];
    default: op1_15_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv26 = 1;
    7: op1_15_inv26 = 1;
    9: op1_15_inv26 = 1;
    11: op1_15_inv26 = 1;
    13: op1_15_inv26 = 1;
    15: op1_15_inv26 = 1;
    16: op1_15_inv26 = 1;
    17: op1_15_inv26 = 1;
    19: op1_15_inv26 = 1;
    22: op1_15_inv26 = 1;
    26: op1_15_inv26 = 1;
    27: op1_15_inv26 = 1;
    29: op1_15_inv26 = 1;
    30: op1_15_inv26 = 1;
    31: op1_15_inv26 = 1;
    33: op1_15_inv26 = 1;
    34: op1_15_inv26 = 1;
    39: op1_15_inv26 = 1;
    40: op1_15_inv26 = 1;
    44: op1_15_inv26 = 1;
    48: op1_15_inv26 = 1;
    51: op1_15_inv26 = 1;
    52: op1_15_inv26 = 1;
    53: op1_15_inv26 = 1;
    56: op1_15_inv26 = 1;
    57: op1_15_inv26 = 1;
    63: op1_15_inv26 = 1;
    65: op1_15_inv26 = 1;
    66: op1_15_inv26 = 1;
    67: op1_15_inv26 = 1;
    69: op1_15_inv26 = 1;
    70: op1_15_inv26 = 1;
    76: op1_15_inv26 = 1;
    77: op1_15_inv26 = 1;
    79: op1_15_inv26 = 1;
    80: op1_15_inv26 = 1;
    81: op1_15_inv26 = 1;
    82: op1_15_inv26 = 1;
    84: op1_15_inv26 = 1;
    90: op1_15_inv26 = 1;
    92: op1_15_inv26 = 1;
    default: op1_15_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の27番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in27 = reg_0019;
    6: op1_15_in27 = imem04_in[55:52];
    7: op1_15_in27 = reg_0407;
    8: op1_15_in27 = reg_0240;
    9: op1_15_in27 = reg_0522;
    10: op1_15_in27 = reg_0270;
    11: op1_15_in27 = imem07_in[91:88];
    12: op1_15_in27 = imem05_in[43:40];
    13: op1_15_in27 = imem07_in[115:112];
    15: op1_15_in27 = imem03_in[7:4];
    16: op1_15_in27 = reg_0063;
    17: op1_15_in27 = reg_0051;
    18: op1_15_in27 = reg_0789;
    19: op1_15_in27 = reg_0364;
    20: op1_15_in27 = reg_0131;
    22: op1_15_in27 = reg_0315;
    23: op1_15_in27 = reg_0512;
    24: op1_15_in27 = reg_0641;
    25: op1_15_in27 = reg_0708;
    26: op1_15_in27 = reg_0385;
    27: op1_15_in27 = reg_0628;
    29: op1_15_in27 = imem03_in[99:96];
    30: op1_15_in27 = reg_0409;
    31: op1_15_in27 = reg_0172;
    33: op1_15_in27 = reg_0140;
    34: op1_15_in27 = imem06_in[47:44];
    35: op1_15_in27 = reg_0776;
    38: op1_15_in27 = reg_0506;
    39: op1_15_in27 = reg_0515;
    40: op1_15_in27 = reg_0301;
    41: op1_15_in27 = reg_0718;
    43: op1_15_in27 = imem02_in[27:24];
    44: op1_15_in27 = reg_0071;
    45: op1_15_in27 = reg_0158;
    46: op1_15_in27 = imem01_in[87:84];
    47: op1_15_in27 = reg_0513;
    48: op1_15_in27 = reg_0309;
    49: op1_15_in27 = imem04_in[27:24];
    62: op1_15_in27 = imem04_in[27:24];
    50: op1_15_in27 = reg_0651;
    51: op1_15_in27 = reg_0419;
    52: op1_15_in27 = imem03_in[91:88];
    53: op1_15_in27 = reg_0596;
    54: op1_15_in27 = imem05_in[67:64];
    55: op1_15_in27 = reg_0623;
    56: op1_15_in27 = imem06_in[119:116];
    57: op1_15_in27 = reg_0052;
    59: op1_15_in27 = reg_0764;
    61: op1_15_in27 = imem02_in[51:48];
    63: op1_15_in27 = reg_0069;
    64: op1_15_in27 = reg_0112;
    65: op1_15_in27 = reg_0143;
    66: op1_15_in27 = imem05_in[127:124];
    67: op1_15_in27 = imem01_in[51:48];
    68: op1_15_in27 = reg_0395;
    69: op1_15_in27 = reg_0408;
    70: op1_15_in27 = imem02_in[23:20];
    71: op1_15_in27 = imem05_in[19:16];
    72: op1_15_in27 = reg_0151;
    73: op1_15_in27 = reg_0722;
    76: op1_15_in27 = reg_0530;
    77: op1_15_in27 = reg_0146;
    78: op1_15_in27 = reg_0279;
    79: op1_15_in27 = reg_0447;
    80: op1_15_in27 = reg_0726;
    81: op1_15_in27 = imem04_in[43:40];
    82: op1_15_in27 = imem02_in[127:124];
    83: op1_15_in27 = reg_0343;
    84: op1_15_in27 = reg_0354;
    85: op1_15_in27 = reg_0138;
    86: op1_15_in27 = imem03_in[55:52];
    87: op1_15_in27 = reg_0613;
    88: op1_15_in27 = reg_0646;
    89: op1_15_in27 = imem05_in[95:92];
    90: op1_15_in27 = reg_0781;
    91: op1_15_in27 = reg_0423;
    92: op1_15_in27 = reg_0258;
    93: op1_15_in27 = imem01_in[95:92];
    default: op1_15_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    4: op1_15_inv27 = 1;
    7: op1_15_inv27 = 1;
    8: op1_15_inv27 = 1;
    10: op1_15_inv27 = 1;
    11: op1_15_inv27 = 1;
    13: op1_15_inv27 = 1;
    17: op1_15_inv27 = 1;
    18: op1_15_inv27 = 1;
    19: op1_15_inv27 = 1;
    20: op1_15_inv27 = 1;
    23: op1_15_inv27 = 1;
    24: op1_15_inv27 = 1;
    26: op1_15_inv27 = 1;
    27: op1_15_inv27 = 1;
    29: op1_15_inv27 = 1;
    31: op1_15_inv27 = 1;
    34: op1_15_inv27 = 1;
    38: op1_15_inv27 = 1;
    39: op1_15_inv27 = 1;
    40: op1_15_inv27 = 1;
    41: op1_15_inv27 = 1;
    43: op1_15_inv27 = 1;
    45: op1_15_inv27 = 1;
    46: op1_15_inv27 = 1;
    47: op1_15_inv27 = 1;
    49: op1_15_inv27 = 1;
    50: op1_15_inv27 = 1;
    54: op1_15_inv27 = 1;
    56: op1_15_inv27 = 1;
    57: op1_15_inv27 = 1;
    61: op1_15_inv27 = 1;
    62: op1_15_inv27 = 1;
    63: op1_15_inv27 = 1;
    64: op1_15_inv27 = 1;
    67: op1_15_inv27 = 1;
    68: op1_15_inv27 = 1;
    69: op1_15_inv27 = 1;
    70: op1_15_inv27 = 1;
    71: op1_15_inv27 = 1;
    72: op1_15_inv27 = 1;
    82: op1_15_inv27 = 1;
    83: op1_15_inv27 = 1;
    84: op1_15_inv27 = 1;
    86: op1_15_inv27 = 1;
    88: op1_15_inv27 = 1;
    89: op1_15_inv27 = 1;
    90: op1_15_inv27 = 1;
    default: op1_15_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の28番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in28 = reg_0014;
    6: op1_15_in28 = imem04_in[59:56];
    7: op1_15_in28 = reg_0404;
    35: op1_15_in28 = reg_0404;
    8: op1_15_in28 = reg_0237;
    9: op1_15_in28 = reg_0513;
    10: op1_15_in28 = reg_0274;
    11: op1_15_in28 = imem07_in[107:104];
    12: op1_15_in28 = imem05_in[47:44];
    13: op1_15_in28 = reg_0723;
    15: op1_15_in28 = imem03_in[23:20];
    16: op1_15_in28 = reg_0075;
    17: op1_15_in28 = reg_0284;
    18: op1_15_in28 = reg_0492;
    19: op1_15_in28 = reg_0320;
    20: op1_15_in28 = imem06_in[3:0];
    22: op1_15_in28 = reg_0555;
    23: op1_15_in28 = reg_0824;
    24: op1_15_in28 = reg_0662;
    25: op1_15_in28 = reg_0709;
    26: op1_15_in28 = reg_0398;
    27: op1_15_in28 = reg_0626;
    29: op1_15_in28 = reg_0583;
    30: op1_15_in28 = reg_0776;
    31: op1_15_in28 = reg_0181;
    33: op1_15_in28 = reg_0134;
    34: op1_15_in28 = imem06_in[79:76];
    38: op1_15_in28 = reg_0239;
    39: op1_15_in28 = imem01_in[11:8];
    40: op1_15_in28 = reg_0305;
    41: op1_15_in28 = reg_0706;
    43: op1_15_in28 = imem02_in[51:48];
    44: op1_15_in28 = reg_0292;
    57: op1_15_in28 = reg_0292;
    46: op1_15_in28 = imem01_in[123:120];
    47: op1_15_in28 = reg_0078;
    48: op1_15_in28 = reg_0226;
    49: op1_15_in28 = imem04_in[67:64];
    50: op1_15_in28 = reg_0665;
    51: op1_15_in28 = reg_0243;
    52: op1_15_in28 = imem03_in[103:100];
    53: op1_15_in28 = reg_0281;
    54: op1_15_in28 = imem05_in[107:104];
    55: op1_15_in28 = imem07_in[3:0];
    56: op1_15_in28 = reg_0774;
    59: op1_15_in28 = reg_0515;
    61: op1_15_in28 = imem02_in[59:56];
    62: op1_15_in28 = imem04_in[39:36];
    63: op1_15_in28 = reg_0780;
    64: op1_15_in28 = imem05_in[51:48];
    65: op1_15_in28 = reg_0141;
    66: op1_15_in28 = reg_0791;
    67: op1_15_in28 = imem01_in[55:52];
    68: op1_15_in28 = reg_0575;
    69: op1_15_in28 = reg_0763;
    70: op1_15_in28 = imem02_in[31:28];
    71: op1_15_in28 = imem05_in[119:116];
    72: op1_15_in28 = reg_0152;
    73: op1_15_in28 = reg_0720;
    76: op1_15_in28 = reg_0756;
    77: op1_15_in28 = reg_0641;
    78: op1_15_in28 = reg_0086;
    79: op1_15_in28 = reg_0445;
    80: op1_15_in28 = reg_0784;
    81: op1_15_in28 = imem04_in[55:52];
    82: op1_15_in28 = reg_0650;
    83: op1_15_in28 = reg_0095;
    84: op1_15_in28 = reg_0238;
    85: op1_15_in28 = reg_0288;
    86: op1_15_in28 = imem03_in[59:56];
    87: op1_15_in28 = reg_0307;
    88: op1_15_in28 = reg_0387;
    89: op1_15_in28 = imem05_in[103:100];
    90: op1_15_in28 = reg_0150;
    91: op1_15_in28 = reg_0574;
    92: op1_15_in28 = reg_0741;
    93: op1_15_in28 = imem01_in[111:108];
    default: op1_15_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    6: op1_15_inv28 = 1;
    7: op1_15_inv28 = 1;
    15: op1_15_inv28 = 1;
    16: op1_15_inv28 = 1;
    19: op1_15_inv28 = 1;
    22: op1_15_inv28 = 1;
    23: op1_15_inv28 = 1;
    24: op1_15_inv28 = 1;
    26: op1_15_inv28 = 1;
    27: op1_15_inv28 = 1;
    29: op1_15_inv28 = 1;
    40: op1_15_inv28 = 1;
    41: op1_15_inv28 = 1;
    43: op1_15_inv28 = 1;
    44: op1_15_inv28 = 1;
    46: op1_15_inv28 = 1;
    47: op1_15_inv28 = 1;
    49: op1_15_inv28 = 1;
    53: op1_15_inv28 = 1;
    54: op1_15_inv28 = 1;
    57: op1_15_inv28 = 1;
    61: op1_15_inv28 = 1;
    62: op1_15_inv28 = 1;
    64: op1_15_inv28 = 1;
    68: op1_15_inv28 = 1;
    70: op1_15_inv28 = 1;
    76: op1_15_inv28 = 1;
    79: op1_15_inv28 = 1;
    83: op1_15_inv28 = 1;
    84: op1_15_inv28 = 1;
    85: op1_15_inv28 = 1;
    89: op1_15_inv28 = 1;
    90: op1_15_inv28 = 1;
    93: op1_15_inv28 = 1;
    default: op1_15_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の29番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in29 = reg_0008;
    6: op1_15_in29 = imem04_in[71:68];
    7: op1_15_in29 = reg_0039;
    8: op1_15_in29 = reg_0234;
    9: op1_15_in29 = reg_0514;
    10: op1_15_in29 = reg_0264;
    11: op1_15_in29 = reg_0719;
    12: op1_15_in29 = imem05_in[71:68];
    13: op1_15_in29 = reg_0703;
    15: op1_15_in29 = imem03_in[27:24];
    16: op1_15_in29 = reg_0064;
    17: op1_15_in29 = reg_0535;
    18: op1_15_in29 = reg_0780;
    19: op1_15_in29 = reg_0341;
    20: op1_15_in29 = imem06_in[39:36];
    22: op1_15_in29 = reg_0060;
    23: op1_15_in29 = reg_0519;
    24: op1_15_in29 = reg_0665;
    25: op1_15_in29 = reg_0718;
    26: op1_15_in29 = reg_0396;
    88: op1_15_in29 = reg_0396;
    27: op1_15_in29 = reg_0622;
    29: op1_15_in29 = reg_0584;
    82: op1_15_in29 = reg_0584;
    30: op1_15_in29 = reg_0319;
    31: op1_15_in29 = reg_0162;
    33: op1_15_in29 = imem06_in[7:4];
    34: op1_15_in29 = imem06_in[95:92];
    35: op1_15_in29 = reg_0028;
    38: op1_15_in29 = reg_0240;
    39: op1_15_in29 = imem01_in[43:40];
    40: op1_15_in29 = reg_0280;
    41: op1_15_in29 = reg_0434;
    43: op1_15_in29 = reg_0658;
    44: op1_15_in29 = reg_0508;
    46: op1_15_in29 = reg_0772;
    47: op1_15_in29 = reg_0585;
    48: op1_15_in29 = reg_0276;
    49: op1_15_in29 = imem04_in[87:84];
    62: op1_15_in29 = imem04_in[87:84];
    50: op1_15_in29 = reg_0667;
    51: op1_15_in29 = reg_0123;
    52: op1_15_in29 = reg_0602;
    53: op1_15_in29 = reg_0588;
    54: op1_15_in29 = imem05_in[111:108];
    55: op1_15_in29 = imem07_in[15:12];
    56: op1_15_in29 = reg_0773;
    57: op1_15_in29 = reg_0431;
    59: op1_15_in29 = reg_0812;
    61: op1_15_in29 = imem02_in[75:72];
    63: op1_15_in29 = imem05_in[11:8];
    64: op1_15_in29 = imem05_in[99:96];
    65: op1_15_in29 = reg_0130;
    66: op1_15_in29 = reg_0256;
    67: op1_15_in29 = imem01_in[87:84];
    68: op1_15_in29 = reg_0373;
    69: op1_15_in29 = reg_0515;
    70: op1_15_in29 = reg_0650;
    71: op1_15_in29 = reg_0337;
    72: op1_15_in29 = reg_0154;
    73: op1_15_in29 = reg_0731;
    76: op1_15_in29 = reg_0538;
    77: op1_15_in29 = reg_0144;
    78: op1_15_in29 = reg_0132;
    79: op1_15_in29 = reg_0444;
    80: op1_15_in29 = reg_0789;
    81: op1_15_in29 = imem04_in[107:104];
    83: op1_15_in29 = reg_0096;
    84: op1_15_in29 = reg_0404;
    85: op1_15_in29 = reg_0495;
    86: op1_15_in29 = reg_0597;
    87: op1_15_in29 = reg_0608;
    89: op1_15_in29 = imem05_in[115:112];
    90: op1_15_in29 = reg_0152;
    91: op1_15_in29 = reg_0054;
    92: op1_15_in29 = reg_0820;
    93: op1_15_in29 = reg_0520;
    default: op1_15_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_15_inv29 = 1;
    12: op1_15_inv29 = 1;
    13: op1_15_inv29 = 1;
    16: op1_15_inv29 = 1;
    17: op1_15_inv29 = 1;
    18: op1_15_inv29 = 1;
    20: op1_15_inv29 = 1;
    22: op1_15_inv29 = 1;
    23: op1_15_inv29 = 1;
    29: op1_15_inv29 = 1;
    30: op1_15_inv29 = 1;
    34: op1_15_inv29 = 1;
    35: op1_15_inv29 = 1;
    38: op1_15_inv29 = 1;
    40: op1_15_inv29 = 1;
    46: op1_15_inv29 = 1;
    48: op1_15_inv29 = 1;
    50: op1_15_inv29 = 1;
    53: op1_15_inv29 = 1;
    54: op1_15_inv29 = 1;
    55: op1_15_inv29 = 1;
    61: op1_15_inv29 = 1;
    63: op1_15_inv29 = 1;
    66: op1_15_inv29 = 1;
    71: op1_15_inv29 = 1;
    77: op1_15_inv29 = 1;
    78: op1_15_inv29 = 1;
    80: op1_15_inv29 = 1;
    81: op1_15_inv29 = 1;
    82: op1_15_inv29 = 1;
    84: op1_15_inv29 = 1;
    86: op1_15_inv29 = 1;
    87: op1_15_inv29 = 1;
    88: op1_15_inv29 = 1;
    89: op1_15_inv29 = 1;
    91: op1_15_inv29 = 1;
    92: op1_15_inv29 = 1;
    default: op1_15_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の30番目の入力
  always @ ( * ) begin
    case ( state )
    4: op1_15_in30 = reg_0015;
    6: op1_15_in30 = imem04_in[83:80];
    7: op1_15_in30 = reg_0036;
    8: op1_15_in30 = reg_0245;
    9: op1_15_in30 = reg_0524;
    10: op1_15_in30 = reg_0269;
    11: op1_15_in30 = reg_0710;
    12: op1_15_in30 = imem05_in[87:84];
    13: op1_15_in30 = reg_0708;
    15: op1_15_in30 = imem03_in[39:36];
    16: op1_15_in30 = reg_0072;
    17: op1_15_in30 = reg_0541;
    18: op1_15_in30 = reg_0784;
    19: op1_15_in30 = reg_0329;
    20: op1_15_in30 = imem06_in[71:68];
    22: op1_15_in30 = reg_0058;
    23: op1_15_in30 = reg_0825;
    24: op1_15_in30 = reg_0341;
    25: op1_15_in30 = reg_0711;
    26: op1_15_in30 = reg_0389;
    27: op1_15_in30 = reg_0601;
    29: op1_15_in30 = reg_0585;
    30: op1_15_in30 = reg_0311;
    31: op1_15_in30 = reg_0167;
    33: op1_15_in30 = imem06_in[15:12];
    34: op1_15_in30 = imem06_in[103:100];
    35: op1_15_in30 = reg_0816;
    38: op1_15_in30 = reg_0243;
    39: op1_15_in30 = imem01_in[67:64];
    40: op1_15_in30 = reg_0529;
    41: op1_15_in30 = reg_0440;
    43: op1_15_in30 = reg_0666;
    44: op1_15_in30 = reg_0257;
    90: op1_15_in30 = reg_0257;
    46: op1_15_in30 = reg_0822;
    47: op1_15_in30 = reg_0643;
    48: op1_15_in30 = reg_0307;
    49: op1_15_in30 = imem04_in[91:88];
    50: op1_15_in30 = reg_0320;
    51: op1_15_in30 = reg_0118;
    52: op1_15_in30 = reg_0582;
    53: op1_15_in30 = imem03_in[23:20];
    54: op1_15_in30 = reg_0796;
    55: op1_15_in30 = imem07_in[83:80];
    56: op1_15_in30 = reg_0821;
    57: op1_15_in30 = reg_0598;
    59: op1_15_in30 = reg_0607;
    61: op1_15_in30 = imem02_in[91:88];
    62: op1_15_in30 = imem04_in[95:92];
    63: op1_15_in30 = imem05_in[23:20];
    64: op1_15_in30 = reg_0215;
    65: op1_15_in30 = reg_0131;
    66: op1_15_in30 = reg_0742;
    71: op1_15_in30 = reg_0742;
    67: op1_15_in30 = imem01_in[91:88];
    68: op1_15_in30 = reg_0572;
    69: op1_15_in30 = reg_0819;
    70: op1_15_in30 = reg_0045;
    72: op1_15_in30 = reg_0153;
    73: op1_15_in30 = reg_0721;
    76: op1_15_in30 = reg_0093;
    77: op1_15_in30 = reg_0789;
    78: op1_15_in30 = reg_0786;
    79: op1_15_in30 = reg_0180;
    80: op1_15_in30 = reg_0434;
    81: op1_15_in30 = imem04_in[127:124];
    82: op1_15_in30 = reg_0639;
    83: op1_15_in30 = reg_0097;
    84: op1_15_in30 = reg_0260;
    85: op1_15_in30 = reg_0393;
    86: op1_15_in30 = reg_0338;
    87: op1_15_in30 = reg_0515;
    88: op1_15_in30 = reg_0623;
    89: op1_15_in30 = imem05_in[119:116];
    91: op1_15_in30 = reg_0567;
    93: op1_15_in30 = reg_0567;
    92: op1_15_in30 = reg_0653;
    default: op1_15_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    9: op1_15_inv30 = 1;
    10: op1_15_inv30 = 1;
    11: op1_15_inv30 = 1;
    12: op1_15_inv30 = 1;
    13: op1_15_inv30 = 1;
    15: op1_15_inv30 = 1;
    17: op1_15_inv30 = 1;
    18: op1_15_inv30 = 1;
    20: op1_15_inv30 = 1;
    23: op1_15_inv30 = 1;
    24: op1_15_inv30 = 1;
    26: op1_15_inv30 = 1;
    29: op1_15_inv30 = 1;
    30: op1_15_inv30 = 1;
    31: op1_15_inv30 = 1;
    34: op1_15_inv30 = 1;
    35: op1_15_inv30 = 1;
    41: op1_15_inv30 = 1;
    43: op1_15_inv30 = 1;
    46: op1_15_inv30 = 1;
    47: op1_15_inv30 = 1;
    48: op1_15_inv30 = 1;
    50: op1_15_inv30 = 1;
    51: op1_15_inv30 = 1;
    53: op1_15_inv30 = 1;
    54: op1_15_inv30 = 1;
    55: op1_15_inv30 = 1;
    61: op1_15_inv30 = 1;
    62: op1_15_inv30 = 1;
    70: op1_15_inv30 = 1;
    72: op1_15_inv30 = 1;
    73: op1_15_inv30 = 1;
    76: op1_15_inv30 = 1;
    77: op1_15_inv30 = 1;
    78: op1_15_inv30 = 1;
    84: op1_15_inv30 = 1;
    85: op1_15_inv30 = 1;
    86: op1_15_inv30 = 1;
    90: op1_15_inv30 = 1;
    93: op1_15_inv30 = 1;
    default: op1_15_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_15_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_15_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_00_in00 = reg_0005;
    7: op2_00_in00 = reg_0005;
    33: op2_00_in00 = reg_0005;
    34: op2_00_in00 = reg_0005;
    38: op2_00_in00 = reg_0005;
    39: op2_00_in00 = reg_0005;
    44: op2_00_in00 = reg_0005;
    47: op2_00_in00 = reg_0005;
    62: op2_00_in00 = reg_0005;
    76: op2_00_in00 = reg_0005;
    77: op2_00_in00 = reg_0005;
    96: op2_00_in00 = reg_0005;
    97: op2_00_in00 = reg_0005;
    6: op2_00_in00 = reg_0778;
    8: op2_00_in00 = reg_0777;
    12: op2_00_in00 = reg_0777;
    18: op2_00_in00 = reg_0777;
    28: op2_00_in00 = reg_0777;
    9: op2_00_in00 = reg_0776;
    10: op2_00_in00 = reg_0020;
    17: op2_00_in00 = reg_0020;
    19: op2_00_in00 = reg_0020;
    21: op2_00_in00 = reg_0020;
    24: op2_00_in00 = reg_0020;
    26: op2_00_in00 = reg_0020;
    31: op2_00_in00 = reg_0020;
    70: op2_00_in00 = reg_0020;
    78: op2_00_in00 = reg_0020;
    84: op2_00_in00 = reg_0020;
    88: op2_00_in00 = reg_0020;
    90: op2_00_in00 = reg_0020;
    11: op2_00_in00 = reg_0779;
    25: op2_00_in00 = reg_0779;
    13: op2_00_in00 = reg_0231;
    15: op2_00_in00 = reg_0231;
    16: op2_00_in00 = reg_0231;
    23: op2_00_in00 = reg_0231;
    27: op2_00_in00 = reg_0231;
    30: op2_00_in00 = reg_0231;
    60: op2_00_in00 = reg_0231;
    14: op2_00_in00 = reg_0043;
    20: op2_00_in00 = reg_0043;
    22: op2_00_in00 = reg_0025;
    58: op2_00_in00 = reg_0025;
    61: op2_00_in00 = reg_0025;
    67: op2_00_in00 = reg_0025;
    89: op2_00_in00 = reg_0025;
    29: op2_00_in00 = reg_0766;
    32: op2_00_in00 = reg_0765;
    37: op2_00_in00 = reg_0765;
    71: op2_00_in00 = reg_0765;
    35: op2_00_in00 = reg_0415;
    36: op2_00_in00 = reg_0414;
    43: op2_00_in00 = reg_0414;
    50: op2_00_in00 = reg_0414;
    40: op2_00_in00 = reg_0021;
    45: op2_00_in00 = reg_0021;
    48: op2_00_in00 = reg_0021;
    72: op2_00_in00 = reg_0021;
    94: op2_00_in00 = reg_0021;
    41: op2_00_in00 = reg_0417;
    42: op2_00_in00 = reg_0634;
    46: op2_00_in00 = reg_0032;
    49: op2_00_in00 = reg_0032;
    51: op2_00_in00 = reg_0032;
    56: op2_00_in00 = reg_0032;
    68: op2_00_in00 = reg_0032;
    73: op2_00_in00 = reg_0032;
    79: op2_00_in00 = reg_0032;
    52: op2_00_in00 = reg_0259;
    54: op2_00_in00 = reg_0259;
    53: op2_00_in00 = reg_0768;
    63: op2_00_in00 = reg_0768;
    69: op2_00_in00 = reg_0768;
    85: op2_00_in00 = reg_0768;
    93: op2_00_in00 = reg_0768;
    95: op2_00_in00 = reg_0768;
    55: op2_00_in00 = reg_0416;
    57: op2_00_in00 = reg_0039;
    59: op2_00_in00 = reg_0501;
    64: op2_00_in00 = reg_0037;
    66: op2_00_in00 = reg_0037;
    74: op2_00_in00 = reg_0037;
    80: op2_00_in00 = reg_0037;
    86: op2_00_in00 = reg_0037;
    65: op2_00_in00 = reg_0113;
    75: op2_00_in00 = reg_0136;
    81: op2_00_in00 = reg_0136;
    83: op2_00_in00 = reg_0136;
    82: op2_00_in00 = reg_0413;
    87: op2_00_in00 = reg_0413;
    91: op2_00_in00 = reg_0014;
    92: op2_00_in00 = reg_0046;
    default: op2_00_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_00_in01 = reg_0011;
    7: op2_00_in01 = reg_0011;
    13: op2_00_in01 = reg_0011;
    15: op2_00_in01 = reg_0011;
    16: op2_00_in01 = reg_0011;
    23: op2_00_in01 = reg_0011;
    27: op2_00_in01 = reg_0011;
    30: op2_00_in01 = reg_0011;
    33: op2_00_in01 = reg_0011;
    34: op2_00_in01 = reg_0011;
    38: op2_00_in01 = reg_0011;
    39: op2_00_in01 = reg_0011;
    44: op2_00_in01 = reg_0011;
    47: op2_00_in01 = reg_0011;
    60: op2_00_in01 = reg_0011;
    62: op2_00_in01 = reg_0011;
    96: op2_00_in01 = reg_0011;
    97: op2_00_in01 = reg_0011;
    6: op2_00_in01 = reg_0779;
    8: op2_00_in01 = reg_0778;
    28: op2_00_in01 = reg_0778;
    9: op2_00_in01 = reg_0501;
    57: op2_00_in01 = reg_0501;
    61: op2_00_in01 = reg_0501;
    86: op2_00_in01 = reg_0501;
    10: op2_00_in01 = reg_0021;
    17: op2_00_in01 = reg_0021;
    19: op2_00_in01 = reg_0021;
    21: op2_00_in01 = reg_0021;
    24: op2_00_in01 = reg_0021;
    26: op2_00_in01 = reg_0021;
    31: op2_00_in01 = reg_0021;
    42: op2_00_in01 = reg_0021;
    52: op2_00_in01 = reg_0021;
    54: op2_00_in01 = reg_0021;
    78: op2_00_in01 = reg_0021;
    84: op2_00_in01 = reg_0021;
    88: op2_00_in01 = reg_0021;
    90: op2_00_in01 = reg_0021;
    11: op2_00_in01 = reg_0231;
    25: op2_00_in01 = reg_0231;
    12: op2_00_in01 = reg_0020;
    14: op2_00_in01 = reg_0020;
    35: op2_00_in01 = reg_0020;
    59: op2_00_in01 = reg_0020;
    64: op2_00_in01 = reg_0020;
    66: op2_00_in01 = reg_0020;
    68: op2_00_in01 = reg_0020;
    73: op2_00_in01 = reg_0020;
    80: op2_00_in01 = reg_0020;
    92: op2_00_in01 = reg_0020;
    18: op2_00_in01 = reg_0073;
    20: op2_00_in01 = reg_0073;
    51: op2_00_in01 = reg_0073;
    22: op2_00_in01 = reg_0043;
    29: op2_00_in01 = reg_0259;
    32: op2_00_in01 = reg_0603;
    36: op2_00_in01 = reg_0603;
    37: op2_00_in01 = reg_0415;
    74: op2_00_in01 = reg_0415;
    40: op2_00_in01 = reg_0005;
    41: op2_00_in01 = reg_0005;
    45: op2_00_in01 = reg_0005;
    48: op2_00_in01 = reg_0005;
    53: op2_00_in01 = reg_0005;
    63: op2_00_in01 = reg_0005;
    69: op2_00_in01 = reg_0005;
    72: op2_00_in01 = reg_0005;
    85: op2_00_in01 = reg_0005;
    93: op2_00_in01 = reg_0005;
    94: op2_00_in01 = reg_0005;
    95: op2_00_in01 = reg_0005;
    43: op2_00_in01 = reg_0032;
    58: op2_00_in01 = reg_0032;
    75: op2_00_in01 = reg_0032;
    81: op2_00_in01 = reg_0032;
    83: op2_00_in01 = reg_0032;
    46: op2_00_in01 = reg_0634;
    49: op2_00_in01 = reg_0634;
    50: op2_00_in01 = reg_0063;
    89: op2_00_in01 = reg_0063;
    55: op2_00_in01 = reg_0768;
    56: op2_00_in01 = reg_0767;
    65: op2_00_in01 = reg_0732;
    67: op2_00_in01 = reg_0113;
    71: op2_00_in01 = reg_0113;
    70: op2_00_in01 = reg_0091;
    76: op2_00_in01 = reg_0754;
    77: op2_00_in01 = reg_0754;
    79: op2_00_in01 = reg_0044;
    82: op2_00_in01 = reg_0037;
    87: op2_00_in01 = reg_0350;
    91: op2_00_in01 = reg_0357;
    default: op2_00_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_00_in02 = reg_0017;
    7: op2_00_in02 = reg_0017;
    13: op2_00_in02 = reg_0017;
    15: op2_00_in02 = reg_0017;
    16: op2_00_in02 = reg_0017;
    23: op2_00_in02 = reg_0017;
    27: op2_00_in02 = reg_0017;
    30: op2_00_in02 = reg_0017;
    33: op2_00_in02 = reg_0017;
    34: op2_00_in02 = reg_0017;
    38: op2_00_in02 = reg_0017;
    39: op2_00_in02 = reg_0017;
    44: op2_00_in02 = reg_0017;
    47: op2_00_in02 = reg_0017;
    60: op2_00_in02 = reg_0017;
    62: op2_00_in02 = reg_0017;
    76: op2_00_in02 = reg_0017;
    77: op2_00_in02 = reg_0017;
    96: op2_00_in02 = reg_0017;
    97: op2_00_in02 = reg_0017;
    6: op2_00_in02 = reg_0005;
    42: op2_00_in02 = reg_0005;
    52: op2_00_in02 = reg_0005;
    54: op2_00_in02 = reg_0005;
    55: op2_00_in02 = reg_0005;
    70: op2_00_in02 = reg_0005;
    78: op2_00_in02 = reg_0005;
    84: op2_00_in02 = reg_0005;
    88: op2_00_in02 = reg_0005;
    90: op2_00_in02 = reg_0005;
    8: op2_00_in02 = reg_0021;
    12: op2_00_in02 = reg_0021;
    14: op2_00_in02 = reg_0021;
    28: op2_00_in02 = reg_0021;
    35: op2_00_in02 = reg_0021;
    56: op2_00_in02 = reg_0021;
    68: op2_00_in02 = reg_0021;
    80: op2_00_in02 = reg_0021;
    92: op2_00_in02 = reg_0021;
    9: op2_00_in02 = reg_0732;
    71: op2_00_in02 = reg_0732;
    10: op2_00_in02 = reg_0231;
    17: op2_00_in02 = reg_0231;
    19: op2_00_in02 = reg_0231;
    21: op2_00_in02 = reg_0231;
    24: op2_00_in02 = reg_0231;
    26: op2_00_in02 = reg_0231;
    31: op2_00_in02 = reg_0231;
    11: op2_00_in02 = reg_0011;
    25: op2_00_in02 = reg_0011;
    40: op2_00_in02 = reg_0011;
    41: op2_00_in02 = reg_0011;
    45: op2_00_in02 = reg_0011;
    48: op2_00_in02 = reg_0011;
    53: op2_00_in02 = reg_0011;
    63: op2_00_in02 = reg_0011;
    69: op2_00_in02 = reg_0011;
    93: op2_00_in02 = reg_0011;
    94: op2_00_in02 = reg_0011;
    95: op2_00_in02 = reg_0011;
    18: op2_00_in02 = reg_0779;
    20: op2_00_in02 = reg_0779;
    29: op2_00_in02 = reg_0779;
    22: op2_00_in02 = reg_0073;
    32: op2_00_in02 = reg_0767;
    43: op2_00_in02 = reg_0767;
    50: op2_00_in02 = reg_0767;
    58: op2_00_in02 = reg_0767;
    89: op2_00_in02 = reg_0767;
    36: op2_00_in02 = reg_0634;
    37: op2_00_in02 = reg_0020;
    61: op2_00_in02 = reg_0020;
    75: op2_00_in02 = reg_0020;
    86: op2_00_in02 = reg_0020;
    46: op2_00_in02 = reg_0768;
    49: op2_00_in02 = reg_0768;
    51: op2_00_in02 = reg_0768;
    59: op2_00_in02 = reg_0768;
    65: op2_00_in02 = reg_0768;
    73: op2_00_in02 = reg_0768;
    79: op2_00_in02 = reg_0768;
    91: op2_00_in02 = reg_0768;
    57: op2_00_in02 = reg_0416;
    64: op2_00_in02 = reg_0091;
    66: op2_00_in02 = reg_0091;
    67: op2_00_in02 = reg_0034;
    72: op2_00_in02 = reg_0754;
    74: op2_00_in02 = reg_0715;
    81: op2_00_in02 = reg_0044;
    83: op2_00_in02 = reg_0044;
    82: op2_00_in02 = reg_0088;
    85: op2_00_in02 = reg_0525;
    87: op2_00_in02 = reg_0351;
    default: op2_00_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_00_in03 = reg_0018;
    7: op2_00_in03 = reg_0018;
    13: op2_00_in03 = reg_0018;
    15: op2_00_in03 = reg_0018;
    16: op2_00_in03 = reg_0018;
    23: op2_00_in03 = reg_0018;
    27: op2_00_in03 = reg_0018;
    30: op2_00_in03 = reg_0018;
    33: op2_00_in03 = reg_0018;
    34: op2_00_in03 = reg_0018;
    38: op2_00_in03 = reg_0018;
    39: op2_00_in03 = reg_0018;
    44: op2_00_in03 = reg_0018;
    47: op2_00_in03 = reg_0018;
    60: op2_00_in03 = reg_0018;
    62: op2_00_in03 = reg_0018;
    76: op2_00_in03 = reg_0018;
    77: op2_00_in03 = reg_0018;
    96: op2_00_in03 = reg_0018;
    97: op2_00_in03 = reg_0018;
    6: op2_00_in03 = reg_0011;
    10: op2_00_in03 = reg_0011;
    17: op2_00_in03 = reg_0011;
    19: op2_00_in03 = reg_0011;
    21: op2_00_in03 = reg_0011;
    24: op2_00_in03 = reg_0011;
    26: op2_00_in03 = reg_0011;
    31: op2_00_in03 = reg_0011;
    42: op2_00_in03 = reg_0011;
    52: op2_00_in03 = reg_0011;
    54: op2_00_in03 = reg_0011;
    55: op2_00_in03 = reg_0011;
    90: op2_00_in03 = reg_0011;
    8: op2_00_in03 = reg_0231;
    12: op2_00_in03 = reg_0231;
    14: op2_00_in03 = reg_0231;
    18: op2_00_in03 = reg_0231;
    20: op2_00_in03 = reg_0231;
    28: op2_00_in03 = reg_0231;
    29: op2_00_in03 = reg_0231;
    59: op2_00_in03 = reg_0231;
    9: op2_00_in03 = reg_0779;
    22: op2_00_in03 = reg_0779;
    11: op2_00_in03 = reg_0017;
    25: op2_00_in03 = reg_0017;
    40: op2_00_in03 = reg_0017;
    41: op2_00_in03 = reg_0017;
    45: op2_00_in03 = reg_0017;
    48: op2_00_in03 = reg_0017;
    53: op2_00_in03 = reg_0017;
    63: op2_00_in03 = reg_0017;
    69: op2_00_in03 = reg_0017;
    72: op2_00_in03 = reg_0017;
    93: op2_00_in03 = reg_0017;
    94: op2_00_in03 = reg_0017;
    95: op2_00_in03 = reg_0017;
    32: op2_00_in03 = reg_0768;
    57: op2_00_in03 = reg_0768;
    61: op2_00_in03 = reg_0768;
    67: op2_00_in03 = reg_0768;
    71: op2_00_in03 = reg_0768;
    81: op2_00_in03 = reg_0768;
    83: op2_00_in03 = reg_0768;
    89: op2_00_in03 = reg_0768;
    35: op2_00_in03 = reg_0005;
    46: op2_00_in03 = reg_0005;
    49: op2_00_in03 = reg_0005;
    51: op2_00_in03 = reg_0005;
    56: op2_00_in03 = reg_0005;
    64: op2_00_in03 = reg_0005;
    65: op2_00_in03 = reg_0005;
    66: op2_00_in03 = reg_0005;
    68: op2_00_in03 = reg_0005;
    73: op2_00_in03 = reg_0005;
    79: op2_00_in03 = reg_0005;
    80: op2_00_in03 = reg_0005;
    91: op2_00_in03 = reg_0005;
    92: op2_00_in03 = reg_0005;
    36: op2_00_in03 = reg_0417;
    43: op2_00_in03 = reg_0417;
    37: op2_00_in03 = reg_0021;
    50: op2_00_in03 = reg_0021;
    58: op2_00_in03 = reg_0021;
    74: op2_00_in03 = reg_0021;
    86: op2_00_in03 = reg_0021;
    70: op2_00_in03 = reg_0754;
    78: op2_00_in03 = reg_0754;
    84: op2_00_in03 = reg_0754;
    88: op2_00_in03 = reg_0754;
    75: op2_00_in03 = reg_0091;
    82: op2_00_in03 = reg_0020;
    87: op2_00_in03 = reg_0357;
    default: op2_00_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_00_in04 = reg_0487;
    15: op2_00_in04 = reg_0487;
    23: op2_00_in04 = reg_0487;
    7: op2_00_in04 = reg_0231;
    9: op2_00_in04 = reg_0231;
    22: op2_00_in04 = reg_0231;
    8: op2_00_in04 = reg_0011;
    14: op2_00_in04 = reg_0011;
    28: op2_00_in04 = reg_0011;
    46: op2_00_in04 = reg_0011;
    49: op2_00_in04 = reg_0011;
    51: op2_00_in04 = reg_0011;
    56: op2_00_in04 = reg_0011;
    59: op2_00_in04 = reg_0011;
    64: op2_00_in04 = reg_0011;
    65: op2_00_in04 = reg_0011;
    66: op2_00_in04 = reg_0011;
    68: op2_00_in04 = reg_0011;
    91: op2_00_in04 = reg_0011;
    92: op2_00_in04 = reg_0011;
    10: op2_00_in04 = reg_0017;
    17: op2_00_in04 = reg_0017;
    21: op2_00_in04 = reg_0017;
    26: op2_00_in04 = reg_0017;
    31: op2_00_in04 = reg_0017;
    52: op2_00_in04 = reg_0017;
    54: op2_00_in04 = reg_0017;
    55: op2_00_in04 = reg_0017;
    70: op2_00_in04 = reg_0017;
    78: op2_00_in04 = reg_0017;
    84: op2_00_in04 = reg_0017;
    88: op2_00_in04 = reg_0017;
    11: op2_00_in04 = reg_0018;
    25: op2_00_in04 = reg_0018;
    40: op2_00_in04 = reg_0018;
    41: op2_00_in04 = reg_0018;
    48: op2_00_in04 = reg_0018;
    53: op2_00_in04 = reg_0018;
    69: op2_00_in04 = reg_0018;
    93: op2_00_in04 = reg_0018;
    94: op2_00_in04 = reg_0018;
    95: op2_00_in04 = reg_0018;
    13: op2_00_in04 = reg_0759;
    16: op2_00_in04 = reg_0761;
    18: op2_00_in04 = reg_0538;
    20: op2_00_in04 = reg_0561;
    27: op2_00_in04 = reg_0766;
    30: op2_00_in04 = reg_0340;
    33: op2_00_in04 = reg_0340;
    38: op2_00_in04 = reg_0340;
    39: op2_00_in04 = reg_0340;
    44: op2_00_in04 = reg_0340;
    47: op2_00_in04 = reg_0340;
    60: op2_00_in04 = reg_0340;
    62: op2_00_in04 = reg_0340;
    76: op2_00_in04 = reg_0340;
    77: op2_00_in04 = reg_0340;
    96: op2_00_in04 = reg_0340;
    97: op2_00_in04 = reg_0340;
    32: op2_00_in04 = reg_0005;
    36: op2_00_in04 = reg_0005;
    37: op2_00_in04 = reg_0005;
    43: op2_00_in04 = reg_0005;
    50: op2_00_in04 = reg_0005;
    57: op2_00_in04 = reg_0005;
    58: op2_00_in04 = reg_0005;
    61: op2_00_in04 = reg_0005;
    67: op2_00_in04 = reg_0005;
    71: op2_00_in04 = reg_0005;
    74: op2_00_in04 = reg_0005;
    75: op2_00_in04 = reg_0005;
    81: op2_00_in04 = reg_0005;
    83: op2_00_in04 = reg_0005;
    86: op2_00_in04 = reg_0005;
    89: op2_00_in04 = reg_0005;
    34: op2_00_in04 = reg_0417;
    35: op2_00_in04 = reg_0635;
    73: op2_00_in04 = reg_0754;
    79: op2_00_in04 = reg_0754;
    80: op2_00_in04 = reg_0754;
    82: op2_00_in04 = reg_0021;
    87: op2_00_in04 = reg_0768;
    default: op2_00_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の5番目の入力
  always @ ( * ) begin
    case ( state )
    8: op2_00_in05 = reg_0754;
    74: op2_00_in05 = reg_0754;
    83: op2_00_in05 = reg_0754;
    10: op2_00_in05 = reg_0018;
    52: op2_00_in05 = reg_0018;
    78: op2_00_in05 = reg_0018;
    84: op2_00_in05 = reg_0018;
    11: op2_00_in05 = reg_0487;
    15: op2_00_in05 = reg_0758;
    21: op2_00_in05 = reg_0764;
    22: op2_00_in05 = reg_0564;
    25: op2_00_in05 = reg_0566;
    26: op2_00_in05 = reg_0400;
    28: op2_00_in05 = reg_0017;
    51: op2_00_in05 = reg_0017;
    64: op2_00_in05 = reg_0017;
    33: op2_00_in05 = reg_0416;
    36: op2_00_in05 = reg_0011;
    50: op2_00_in05 = reg_0011;
    67: op2_00_in05 = reg_0011;
    38: op2_00_in05 = reg_0366;
    97: op2_00_in05 = reg_0366;
    41: op2_00_in05 = reg_0340;
    93: op2_00_in05 = reg_0340;
    94: op2_00_in05 = reg_0340;
    95: op2_00_in05 = reg_0340;
    82: op2_00_in05 = reg_0005;
    87: op2_00_in05 = reg_0005;
    default: op2_00_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の6番目の入力
  always @ ( * ) begin
    case ( state )
    10: op2_00_in06 = reg_0487;
    52: op2_00_in06 = reg_0340;
    84: op2_00_in06 = reg_0340;
    83: op2_00_in06 = reg_0017;
    87: op2_00_in06 = reg_0754;
    default: op2_00_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の7番目の入力
  always @ ( * ) begin
    case ( state )
    10: op2_00_in07 = reg_0769;
    83: op2_00_in07 = reg_0018;
    87: op2_00_in07 = reg_0017;
    default: op2_00_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の8番目の入力
  always @ ( * ) begin
    case ( state )
    10: op2_00_in08 = reg_0756;
    default: op2_00_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#0のバイアス入力
  always @ ( * ) begin
    case ( state )
    5: op2_00_bias = 80;
    6: op2_00_bias = 57;
    7: op2_00_bias = 62;
    8: op2_00_bias = 81;
    9: op2_00_bias = 72;
    10: op2_00_bias = 131;
    11: op2_00_bias = 87;
    12: op2_00_bias = 59;
    13: op2_00_bias = 70;
    14: op2_00_bias = 70;
    15: op2_00_bias = 93;
    16: op2_00_bias = 62;
    17: op2_00_bias = 75;
    18: op2_00_bias = 77;
    19: op2_00_bias = 51;
    20: op2_00_bias = 75;
    21: op2_00_bias = 82;
    22: op2_00_bias = 78;
    23: op2_00_bias = 77;
    24: op2_00_bias = 68;
    25: op2_00_bias = 79;
    26: op2_00_bias = 72;
    27: op2_00_bias = 65;
    28: op2_00_bias = 101;
    29: op2_00_bias = 67;
    30: op2_00_bias = 65;
    31: op2_00_bias = 71;
    32: op2_00_bias = 76;
    33: op2_00_bias = 72;
    34: op2_00_bias = 61;
    35: op2_00_bias = 68;
    36: op2_00_bias = 73;
    37: op2_00_bias = 75;
    38: op2_00_bias = 85;
    39: op2_00_bias = 68;
    40: op2_00_bias = 69;
    41: op2_00_bias = 92;
    42: op2_00_bias = 53;
    43: op2_00_bias = 75;
    44: op2_00_bias = 66;
    45: op2_00_bias = 60;
    46: op2_00_bias = 84;
    47: op2_00_bias = 69;
    48: op2_00_bias = 64;
    49: op2_00_bias = 75;
    50: op2_00_bias = 83;
    51: op2_00_bias = 78;
    52: op2_00_bias = 83;
    53: op2_00_bias = 65;
    54: op2_00_bias = 78;
    55: op2_00_bias = 79;
    56: op2_00_bias = 81;
    57: op2_00_bias = 72;
    58: op2_00_bias = 75;
    59: op2_00_bias = 68;
    60: op2_00_bias = 84;
    61: op2_00_bias = 72;
    62: op2_00_bias = 64;
    63: op2_00_bias = 55;
    64: op2_00_bias = 74;
    65: op2_00_bias = 74;
    66: op2_00_bias = 71;
    67: op2_00_bias = 98;
    68: op2_00_bias = 79;
    69: op2_00_bias = 78;
    70: op2_00_bias = 66;
    71: op2_00_bias = 70;
    72: op2_00_bias = 63;
    73: op2_00_bias = 63;
    74: op2_00_bias = 84;
    75: op2_00_bias = 71;
    76: op2_00_bias = 69;
    77: op2_00_bias = 63;
    78: op2_00_bias = 73;
    79: op2_00_bias = 71;
    80: op2_00_bias = 75;
    81: op2_00_bias = 69;
    82: op2_00_bias = 73;
    83: op2_00_bias = 107;
    84: op2_00_bias = 102;
    85: op2_00_bias = 57;
    86: op2_00_bias = 84;
    87: op2_00_bias = 119;
    88: op2_00_bias = 74;
    89: op2_00_bias = 78;
    90: op2_00_bias = 72;
    91: op2_00_bias = 78;
    92: op2_00_bias = 65;
    93: op2_00_bias = 88;
    94: op2_00_bias = 72;
    95: op2_00_bias = 78;
    96: op2_00_bias = 67;
    97: op2_00_bias = 89;
    default: op2_00_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#1の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_01_in00 = reg_0769;
    11: op2_01_in00 = reg_0769;
    6: op2_01_in00 = reg_0017;
    8: op2_01_in00 = reg_0017;
    14: op2_01_in00 = reg_0017;
    19: op2_01_in00 = reg_0017;
    24: op2_01_in00 = reg_0017;
    36: op2_01_in00 = reg_0017;
    42: op2_01_in00 = reg_0017;
    46: op2_01_in00 = reg_0017;
    49: op2_01_in00 = reg_0017;
    50: op2_01_in00 = reg_0017;
    56: op2_01_in00 = reg_0017;
    59: op2_01_in00 = reg_0017;
    65: op2_01_in00 = reg_0017;
    66: op2_01_in00 = reg_0017;
    67: op2_01_in00 = reg_0017;
    68: op2_01_in00 = reg_0017;
    73: op2_01_in00 = reg_0017;
    74: op2_01_in00 = reg_0017;
    79: op2_01_in00 = reg_0017;
    80: op2_01_in00 = reg_0017;
    85: op2_01_in00 = reg_0017;
    90: op2_01_in00 = reg_0017;
    91: op2_01_in00 = reg_0017;
    92: op2_01_in00 = reg_0017;
    7: op2_01_in00 = reg_0487;
    13: op2_01_in00 = reg_0487;
    16: op2_01_in00 = reg_0487;
    9: op2_01_in00 = reg_0011;
    12: op2_01_in00 = reg_0011;
    18: op2_01_in00 = reg_0011;
    20: op2_01_in00 = reg_0011;
    22: op2_01_in00 = reg_0011;
    29: op2_01_in00 = reg_0011;
    32: op2_01_in00 = reg_0011;
    35: op2_01_in00 = reg_0011;
    37: op2_01_in00 = reg_0011;
    43: op2_01_in00 = reg_0011;
    57: op2_01_in00 = reg_0011;
    58: op2_01_in00 = reg_0011;
    61: op2_01_in00 = reg_0011;
    89: op2_01_in00 = reg_0011;
    10: op2_01_in00 = reg_0770;
    15: op2_01_in00 = reg_0759;
    17: op2_01_in00 = reg_0018;
    21: op2_01_in00 = reg_0018;
    26: op2_01_in00 = reg_0018;
    28: op2_01_in00 = reg_0018;
    31: op2_01_in00 = reg_0018;
    45: op2_01_in00 = reg_0018;
    51: op2_01_in00 = reg_0018;
    54: op2_01_in00 = reg_0018;
    55: op2_01_in00 = reg_0018;
    63: op2_01_in00 = reg_0018;
    64: op2_01_in00 = reg_0018;
    70: op2_01_in00 = reg_0018;
    72: op2_01_in00 = reg_0018;
    87: op2_01_in00 = reg_0018;
    88: op2_01_in00 = reg_0018;
    23: op2_01_in00 = reg_0561;
    25: op2_01_in00 = reg_0340;
    27: op2_01_in00 = reg_0340;
    34: op2_01_in00 = reg_0340;
    40: op2_01_in00 = reg_0340;
    48: op2_01_in00 = reg_0340;
    53: op2_01_in00 = reg_0340;
    69: op2_01_in00 = reg_0340;
    78: op2_01_in00 = reg_0340;
    83: op2_01_in00 = reg_0340;
    30: op2_01_in00 = reg_0366;
    33: op2_01_in00 = reg_0366;
    39: op2_01_in00 = reg_0366;
    41: op2_01_in00 = reg_0366;
    44: op2_01_in00 = reg_0366;
    47: op2_01_in00 = reg_0366;
    52: op2_01_in00 = reg_0366;
    60: op2_01_in00 = reg_0366;
    62: op2_01_in00 = reg_0366;
    76: op2_01_in00 = reg_0366;
    77: op2_01_in00 = reg_0366;
    84: op2_01_in00 = reg_0366;
    93: op2_01_in00 = reg_0366;
    94: op2_01_in00 = reg_0366;
    95: op2_01_in00 = reg_0366;
    96: op2_01_in00 = reg_0366;
    38: op2_01_in00 = reg_0378;
    97: op2_01_in00 = reg_0378;
    71: op2_01_in00 = reg_0754;
    75: op2_01_in00 = reg_0754;
    81: op2_01_in00 = reg_0754;
    82: op2_01_in00 = reg_0754;
    86: op2_01_in00 = reg_0754;
    default: op2_01_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_01_in01 = reg_0770;
    11: op2_01_in01 = reg_0770;
    6: op2_01_in01 = reg_0018;
    8: op2_01_in01 = reg_0018;
    14: op2_01_in01 = reg_0018;
    19: op2_01_in01 = reg_0018;
    24: op2_01_in01 = reg_0018;
    36: op2_01_in01 = reg_0018;
    42: op2_01_in01 = reg_0018;
    46: op2_01_in01 = reg_0018;
    49: op2_01_in01 = reg_0018;
    50: op2_01_in01 = reg_0018;
    56: op2_01_in01 = reg_0018;
    59: op2_01_in01 = reg_0018;
    65: op2_01_in01 = reg_0018;
    66: op2_01_in01 = reg_0018;
    67: op2_01_in01 = reg_0018;
    68: op2_01_in01 = reg_0018;
    73: op2_01_in01 = reg_0018;
    74: op2_01_in01 = reg_0018;
    79: op2_01_in01 = reg_0018;
    80: op2_01_in01 = reg_0018;
    85: op2_01_in01 = reg_0018;
    90: op2_01_in01 = reg_0018;
    91: op2_01_in01 = reg_0018;
    92: op2_01_in01 = reg_0018;
    7: op2_01_in01 = reg_0769;
    9: op2_01_in01 = reg_0017;
    12: op2_01_in01 = reg_0017;
    18: op2_01_in01 = reg_0017;
    20: op2_01_in01 = reg_0017;
    22: op2_01_in01 = reg_0017;
    29: op2_01_in01 = reg_0017;
    32: op2_01_in01 = reg_0017;
    35: op2_01_in01 = reg_0017;
    37: op2_01_in01 = reg_0017;
    43: op2_01_in01 = reg_0017;
    57: op2_01_in01 = reg_0017;
    58: op2_01_in01 = reg_0017;
    61: op2_01_in01 = reg_0017;
    71: op2_01_in01 = reg_0017;
    75: op2_01_in01 = reg_0017;
    81: op2_01_in01 = reg_0017;
    82: op2_01_in01 = reg_0017;
    86: op2_01_in01 = reg_0017;
    89: op2_01_in01 = reg_0017;
    10: op2_01_in01 = reg_0771;
    13: op2_01_in01 = reg_0758;
    16: op2_01_in01 = reg_0758;
    15: op2_01_in01 = reg_0760;
    17: op2_01_in01 = reg_0487;
    21: op2_01_in01 = reg_0487;
    23: op2_01_in01 = reg_0562;
    25: op2_01_in01 = reg_0366;
    27: op2_01_in01 = reg_0366;
    34: op2_01_in01 = reg_0366;
    40: op2_01_in01 = reg_0366;
    48: op2_01_in01 = reg_0366;
    53: op2_01_in01 = reg_0366;
    69: op2_01_in01 = reg_0366;
    78: op2_01_in01 = reg_0366;
    83: op2_01_in01 = reg_0366;
    26: op2_01_in01 = reg_0340;
    28: op2_01_in01 = reg_0340;
    31: op2_01_in01 = reg_0340;
    45: op2_01_in01 = reg_0340;
    51: op2_01_in01 = reg_0340;
    54: op2_01_in01 = reg_0340;
    55: op2_01_in01 = reg_0340;
    63: op2_01_in01 = reg_0340;
    64: op2_01_in01 = reg_0340;
    70: op2_01_in01 = reg_0340;
    72: op2_01_in01 = reg_0340;
    87: op2_01_in01 = reg_0340;
    88: op2_01_in01 = reg_0340;
    30: op2_01_in01 = reg_0378;
    33: op2_01_in01 = reg_0378;
    39: op2_01_in01 = reg_0378;
    41: op2_01_in01 = reg_0378;
    44: op2_01_in01 = reg_0378;
    47: op2_01_in01 = reg_0378;
    52: op2_01_in01 = reg_0378;
    60: op2_01_in01 = reg_0378;
    62: op2_01_in01 = reg_0378;
    76: op2_01_in01 = reg_0378;
    77: op2_01_in01 = reg_0378;
    84: op2_01_in01 = reg_0378;
    93: op2_01_in01 = reg_0378;
    94: op2_01_in01 = reg_0378;
    95: op2_01_in01 = reg_0378;
    96: op2_01_in01 = reg_0378;
    38: op2_01_in01 = reg_0400;
    97: op2_01_in01 = reg_0400;
    default: op2_01_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_01_in02 = reg_0771;
    11: op2_01_in02 = reg_0771;
    6: op2_01_in02 = reg_0487;
    8: op2_01_in02 = reg_0487;
    14: op2_01_in02 = reg_0487;
    19: op2_01_in02 = reg_0487;
    7: op2_01_in02 = reg_0770;
    13: op2_01_in02 = reg_0770;
    9: op2_01_in02 = reg_0018;
    12: op2_01_in02 = reg_0018;
    18: op2_01_in02 = reg_0018;
    20: op2_01_in02 = reg_0018;
    22: op2_01_in02 = reg_0018;
    29: op2_01_in02 = reg_0018;
    32: op2_01_in02 = reg_0018;
    35: op2_01_in02 = reg_0018;
    37: op2_01_in02 = reg_0018;
    43: op2_01_in02 = reg_0018;
    57: op2_01_in02 = reg_0018;
    58: op2_01_in02 = reg_0018;
    61: op2_01_in02 = reg_0018;
    71: op2_01_in02 = reg_0018;
    75: op2_01_in02 = reg_0018;
    81: op2_01_in02 = reg_0018;
    82: op2_01_in02 = reg_0018;
    86: op2_01_in02 = reg_0018;
    89: op2_01_in02 = reg_0018;
    10: op2_01_in02 = reg_0772;
    15: op2_01_in02 = reg_0772;
    16: op2_01_in02 = reg_0759;
    17: op2_01_in02 = reg_0758;
    21: op2_01_in02 = reg_0561;
    23: op2_01_in02 = reg_0564;
    24: op2_01_in02 = reg_0340;
    36: op2_01_in02 = reg_0340;
    42: op2_01_in02 = reg_0340;
    46: op2_01_in02 = reg_0340;
    49: op2_01_in02 = reg_0340;
    50: op2_01_in02 = reg_0340;
    56: op2_01_in02 = reg_0340;
    59: op2_01_in02 = reg_0340;
    65: op2_01_in02 = reg_0340;
    66: op2_01_in02 = reg_0340;
    67: op2_01_in02 = reg_0340;
    68: op2_01_in02 = reg_0340;
    73: op2_01_in02 = reg_0340;
    74: op2_01_in02 = reg_0340;
    79: op2_01_in02 = reg_0340;
    80: op2_01_in02 = reg_0340;
    85: op2_01_in02 = reg_0340;
    90: op2_01_in02 = reg_0340;
    91: op2_01_in02 = reg_0340;
    92: op2_01_in02 = reg_0340;
    25: op2_01_in02 = reg_0562;
    26: op2_01_in02 = reg_0366;
    28: op2_01_in02 = reg_0366;
    31: op2_01_in02 = reg_0366;
    45: op2_01_in02 = reg_0366;
    51: op2_01_in02 = reg_0366;
    54: op2_01_in02 = reg_0366;
    55: op2_01_in02 = reg_0366;
    63: op2_01_in02 = reg_0366;
    64: op2_01_in02 = reg_0366;
    70: op2_01_in02 = reg_0366;
    72: op2_01_in02 = reg_0366;
    87: op2_01_in02 = reg_0366;
    88: op2_01_in02 = reg_0366;
    27: op2_01_in02 = reg_0378;
    34: op2_01_in02 = reg_0378;
    40: op2_01_in02 = reg_0378;
    48: op2_01_in02 = reg_0378;
    53: op2_01_in02 = reg_0378;
    69: op2_01_in02 = reg_0378;
    78: op2_01_in02 = reg_0378;
    83: op2_01_in02 = reg_0378;
    30: op2_01_in02 = reg_0400;
    33: op2_01_in02 = reg_0400;
    39: op2_01_in02 = reg_0400;
    41: op2_01_in02 = reg_0400;
    44: op2_01_in02 = reg_0400;
    47: op2_01_in02 = reg_0400;
    52: op2_01_in02 = reg_0400;
    60: op2_01_in02 = reg_0400;
    62: op2_01_in02 = reg_0400;
    76: op2_01_in02 = reg_0400;
    77: op2_01_in02 = reg_0400;
    84: op2_01_in02 = reg_0400;
    93: op2_01_in02 = reg_0400;
    94: op2_01_in02 = reg_0400;
    95: op2_01_in02 = reg_0400;
    96: op2_01_in02 = reg_0400;
    38: op2_01_in02 = reg_0410;
    97: op2_01_in02 = reg_0410;
    default: op2_01_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_01_in03 = reg_0772;
    11: op2_01_in03 = reg_0772;
    6: op2_01_in03 = reg_0769;
    8: op2_01_in03 = reg_0769;
    7: op2_01_in03 = reg_0771;
    13: op2_01_in03 = reg_0771;
    9: op2_01_in03 = reg_0487;
    12: op2_01_in03 = reg_0487;
    18: op2_01_in03 = reg_0487;
    20: op2_01_in03 = reg_0487;
    22: op2_01_in03 = reg_0487;
    10: op2_01_in03 = reg_0773;
    15: op2_01_in03 = reg_0773;
    14: op2_01_in03 = reg_0758;
    19: op2_01_in03 = reg_0758;
    16: op2_01_in03 = reg_0760;
    17: op2_01_in03 = reg_0759;
    21: op2_01_in03 = reg_0562;
    23: op2_01_in03 = reg_0565;
    24: op2_01_in03 = reg_0561;
    25: op2_01_in03 = reg_0564;
    26: op2_01_in03 = reg_0378;
    28: op2_01_in03 = reg_0378;
    31: op2_01_in03 = reg_0378;
    45: op2_01_in03 = reg_0378;
    51: op2_01_in03 = reg_0378;
    54: op2_01_in03 = reg_0378;
    55: op2_01_in03 = reg_0378;
    63: op2_01_in03 = reg_0378;
    64: op2_01_in03 = reg_0378;
    70: op2_01_in03 = reg_0378;
    72: op2_01_in03 = reg_0378;
    87: op2_01_in03 = reg_0378;
    88: op2_01_in03 = reg_0378;
    27: op2_01_in03 = reg_0400;
    34: op2_01_in03 = reg_0400;
    40: op2_01_in03 = reg_0400;
    48: op2_01_in03 = reg_0400;
    53: op2_01_in03 = reg_0400;
    69: op2_01_in03 = reg_0400;
    78: op2_01_in03 = reg_0400;
    83: op2_01_in03 = reg_0400;
    29: op2_01_in03 = reg_0340;
    32: op2_01_in03 = reg_0340;
    35: op2_01_in03 = reg_0340;
    37: op2_01_in03 = reg_0340;
    43: op2_01_in03 = reg_0340;
    57: op2_01_in03 = reg_0340;
    58: op2_01_in03 = reg_0340;
    61: op2_01_in03 = reg_0340;
    71: op2_01_in03 = reg_0340;
    75: op2_01_in03 = reg_0340;
    81: op2_01_in03 = reg_0340;
    82: op2_01_in03 = reg_0340;
    86: op2_01_in03 = reg_0340;
    89: op2_01_in03 = reg_0340;
    30: op2_01_in03 = reg_0410;
    33: op2_01_in03 = reg_0410;
    39: op2_01_in03 = reg_0410;
    41: op2_01_in03 = reg_0410;
    44: op2_01_in03 = reg_0410;
    47: op2_01_in03 = reg_0410;
    52: op2_01_in03 = reg_0410;
    60: op2_01_in03 = reg_0410;
    62: op2_01_in03 = reg_0410;
    76: op2_01_in03 = reg_0410;
    77: op2_01_in03 = reg_0410;
    84: op2_01_in03 = reg_0410;
    93: op2_01_in03 = reg_0410;
    94: op2_01_in03 = reg_0410;
    95: op2_01_in03 = reg_0410;
    96: op2_01_in03 = reg_0410;
    36: op2_01_in03 = reg_0366;
    42: op2_01_in03 = reg_0366;
    46: op2_01_in03 = reg_0366;
    49: op2_01_in03 = reg_0366;
    50: op2_01_in03 = reg_0366;
    56: op2_01_in03 = reg_0366;
    59: op2_01_in03 = reg_0366;
    65: op2_01_in03 = reg_0366;
    66: op2_01_in03 = reg_0366;
    67: op2_01_in03 = reg_0366;
    68: op2_01_in03 = reg_0366;
    73: op2_01_in03 = reg_0366;
    74: op2_01_in03 = reg_0366;
    79: op2_01_in03 = reg_0366;
    80: op2_01_in03 = reg_0366;
    85: op2_01_in03 = reg_0366;
    90: op2_01_in03 = reg_0366;
    91: op2_01_in03 = reg_0366;
    92: op2_01_in03 = reg_0366;
    38: op2_01_in03 = reg_0411;
    97: op2_01_in03 = reg_0411;
    default: op2_01_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_01_in04 = reg_0773;
    7: op2_01_in04 = reg_0772;
    16: op2_01_in04 = reg_0772;
    8: op2_01_in04 = reg_0770;
    9: op2_01_in04 = reg_0755;
    10: op2_01_in04 = reg_0774;
    15: op2_01_in04 = reg_0774;
    11: op2_01_in04 = reg_0757;
    12: op2_01_in04 = reg_0769;
    14: op2_01_in04 = reg_0759;
    19: op2_01_in04 = reg_0759;
    17: op2_01_in04 = reg_0760;
    21: op2_01_in04 = reg_0760;
    20: op2_01_in04 = reg_0562;
    22: op2_01_in04 = reg_0565;
    25: op2_01_in04 = reg_0565;
    27: op2_01_in04 = reg_0565;
    23: op2_01_in04 = reg_0762;
    26: op2_01_in04 = reg_0765;
    28: op2_01_in04 = reg_0400;
    31: op2_01_in04 = reg_0400;
    45: op2_01_in04 = reg_0400;
    51: op2_01_in04 = reg_0400;
    54: op2_01_in04 = reg_0400;
    55: op2_01_in04 = reg_0400;
    63: op2_01_in04 = reg_0400;
    64: op2_01_in04 = reg_0400;
    72: op2_01_in04 = reg_0400;
    87: op2_01_in04 = reg_0400;
    88: op2_01_in04 = reg_0400;
    29: op2_01_in04 = reg_0411;
    33: op2_01_in04 = reg_0411;
    39: op2_01_in04 = reg_0411;
    44: op2_01_in04 = reg_0411;
    47: op2_01_in04 = reg_0411;
    52: op2_01_in04 = reg_0411;
    60: op2_01_in04 = reg_0411;
    62: op2_01_in04 = reg_0411;
    76: op2_01_in04 = reg_0411;
    84: op2_01_in04 = reg_0411;
    93: op2_01_in04 = reg_0411;
    94: op2_01_in04 = reg_0411;
    95: op2_01_in04 = reg_0411;
    32: op2_01_in04 = reg_0366;
    35: op2_01_in04 = reg_0366;
    37: op2_01_in04 = reg_0366;
    43: op2_01_in04 = reg_0366;
    57: op2_01_in04 = reg_0366;
    58: op2_01_in04 = reg_0366;
    61: op2_01_in04 = reg_0366;
    71: op2_01_in04 = reg_0366;
    75: op2_01_in04 = reg_0366;
    81: op2_01_in04 = reg_0366;
    82: op2_01_in04 = reg_0366;
    86: op2_01_in04 = reg_0366;
    34: op2_01_in04 = reg_0410;
    40: op2_01_in04 = reg_0410;
    53: op2_01_in04 = reg_0410;
    69: op2_01_in04 = reg_0410;
    78: op2_01_in04 = reg_0410;
    36: op2_01_in04 = reg_0378;
    42: op2_01_in04 = reg_0378;
    46: op2_01_in04 = reg_0378;
    49: op2_01_in04 = reg_0378;
    50: op2_01_in04 = reg_0378;
    56: op2_01_in04 = reg_0378;
    59: op2_01_in04 = reg_0378;
    65: op2_01_in04 = reg_0378;
    66: op2_01_in04 = reg_0378;
    67: op2_01_in04 = reg_0378;
    73: op2_01_in04 = reg_0378;
    74: op2_01_in04 = reg_0378;
    79: op2_01_in04 = reg_0378;
    80: op2_01_in04 = reg_0378;
    85: op2_01_in04 = reg_0378;
    90: op2_01_in04 = reg_0378;
    91: op2_01_in04 = reg_0378;
    92: op2_01_in04 = reg_0378;
    38: op2_01_in04 = reg_0412;
    97: op2_01_in04 = reg_0412;
    default: op2_01_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の5番目の入力
  always @ ( * ) begin
    case ( state )
    10: op2_01_in05 = reg_0526;
    15: op2_01_in05 = reg_0287;
    17: op2_01_in05 = reg_0762;
    19: op2_01_in05 = reg_0760;
    25: op2_01_in05 = reg_0378;
    57: op2_01_in05 = reg_0378;
    82: op2_01_in05 = reg_0378;
    28: op2_01_in05 = reg_0410;
    51: op2_01_in05 = reg_0410;
    54: op2_01_in05 = reg_0410;
    87: op2_01_in05 = reg_0410;
    32: op2_01_in05 = reg_0413;
    38: op2_01_in05 = reg_0413;
    33: op2_01_in05 = reg_0412;
    60: op2_01_in05 = reg_0412;
    50: op2_01_in05 = reg_0400;
    56: op2_01_in05 = reg_0400;
    79: op2_01_in05 = reg_0400;
    default: op2_01_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の6番目の入力
  always @ ( * ) begin
    case ( state )
    60: op2_01_in06 = reg_0413;
    default: op2_01_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#1のバイアス入力
  always @ ( * ) begin
    case ( state )
    5: op2_01_bias = 67;
    6: op2_01_bias = 55;
    7: op2_01_bias = 63;
    8: op2_01_bias = 83;
    9: op2_01_bias = 62;
    10: op2_01_bias = 67;
    11: op2_01_bias = 74;
    12: op2_01_bias = 64;
    13: op2_01_bias = 60;
    14: op2_01_bias = 74;
    15: op2_01_bias = 89;
    16: op2_01_bias = 71;
    17: op2_01_bias = 79;
    18: op2_01_bias = 58;
    19: op2_01_bias = 86;
    20: op2_01_bias = 53;
    21: op2_01_bias = 79;
    22: op2_01_bias = 65;
    23: op2_01_bias = 70;
    24: op2_01_bias = 63;
    25: op2_01_bias = 90;
    26: op2_01_bias = 72;
    27: op2_01_bias = 74;
    28: op2_01_bias = 70;
    29: op2_01_bias = 62;
    30: op2_01_bias = 55;
    31: op2_01_bias = 82;
    32: op2_01_bias = 70;
    33: op2_01_bias = 82;
    34: op2_01_bias = 67;
    35: op2_01_bias = 69;
    36: op2_01_bias = 62;
    37: op2_01_bias = 71;
    38: op2_01_bias = 84;
    39: op2_01_bias = 71;
    40: op2_01_bias = 69;
    41: op2_01_bias = 64;
    42: op2_01_bias = 73;
    43: op2_01_bias = 66;
    44: op2_01_bias = 65;
    45: op2_01_bias = 56;
    46: op2_01_bias = 64;
    47: op2_01_bias = 76;
    48: op2_01_bias = 65;
    49: op2_01_bias = 58;
    50: op2_01_bias = 80;
    51: op2_01_bias = 90;
    52: op2_01_bias = 72;
    53: op2_01_bias = 77;
    54: op2_01_bias = 86;
    55: op2_01_bias = 64;
    56: op2_01_bias = 81;
    57: op2_01_bias = 79;
    58: op2_01_bias = 77;
    59: op2_01_bias = 84;
    60: op2_01_bias = 118;
    61: op2_01_bias = 69;
    62: op2_01_bias = 68;
    63: op2_01_bias = 73;
    64: op2_01_bias = 69;
    65: op2_01_bias = 71;
    66: op2_01_bias = 64;
    67: op2_01_bias = 64;
    68: op2_01_bias = 64;
    69: op2_01_bias = 72;
    70: op2_01_bias = 51;
    71: op2_01_bias = 78;
    72: op2_01_bias = 68;
    73: op2_01_bias = 74;
    74: op2_01_bias = 61;
    75: op2_01_bias = 82;
    76: op2_01_bias = 57;
    77: op2_01_bias = 61;
    78: op2_01_bias = 58;
    79: op2_01_bias = 81;
    80: op2_01_bias = 56;
    81: op2_01_bias = 72;
    82: op2_01_bias = 84;
    83: op2_01_bias = 57;
    84: op2_01_bias = 61;
    85: op2_01_bias = 74;
    86: op2_01_bias = 71;
    87: op2_01_bias = 86;
    88: op2_01_bias = 61;
    89: op2_01_bias = 64;
    90: op2_01_bias = 87;
    91: op2_01_bias = 63;
    92: op2_01_bias = 72;
    93: op2_01_bias = 72;
    94: op2_01_bias = 84;
    95: op2_01_bias = 83;
    96: op2_01_bias = 50;
    97: op2_01_bias = 64;
    default: op2_01_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#2の0番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_02_in00 = reg_0774;
    6: op2_02_in00 = reg_0770;
    12: op2_02_in00 = reg_0770;
    7: op2_02_in00 = reg_0773;
    11: op2_02_in00 = reg_0773;
    16: op2_02_in00 = reg_0773;
    8: op2_02_in00 = reg_0771;
    14: op2_02_in00 = reg_0771;
    9: op2_02_in00 = reg_0769;
    10: op2_02_in00 = reg_0775;
    15: op2_02_in00 = reg_0775;
    13: op2_02_in00 = reg_0772;
    17: op2_02_in00 = reg_0761;
    19: op2_02_in00 = reg_0761;
    21: op2_02_in00 = reg_0761;
    18: op2_02_in00 = reg_0758;
    20: op2_02_in00 = reg_0758;
    22: op2_02_in00 = reg_0561;
    23: op2_02_in00 = reg_0763;
    24: op2_02_in00 = reg_0562;
    25: op2_02_in00 = reg_0762;
    26: op2_02_in00 = reg_0564;
    27: op2_02_in00 = reg_0566;
    28: op2_02_in00 = reg_0565;
    29: op2_02_in00 = reg_0366;
    89: op2_02_in00 = reg_0366;
    30: op2_02_in00 = reg_0411;
    34: op2_02_in00 = reg_0411;
    40: op2_02_in00 = reg_0411;
    41: op2_02_in00 = reg_0411;
    51: op2_02_in00 = reg_0411;
    53: op2_02_in00 = reg_0411;
    54: op2_02_in00 = reg_0411;
    69: op2_02_in00 = reg_0411;
    77: op2_02_in00 = reg_0411;
    78: op2_02_in00 = reg_0411;
    87: op2_02_in00 = reg_0411;
    96: op2_02_in00 = reg_0411;
    31: op2_02_in00 = reg_0410;
    45: op2_02_in00 = reg_0410;
    48: op2_02_in00 = reg_0410;
    50: op2_02_in00 = reg_0410;
    55: op2_02_in00 = reg_0410;
    56: op2_02_in00 = reg_0410;
    63: op2_02_in00 = reg_0410;
    64: op2_02_in00 = reg_0410;
    72: op2_02_in00 = reg_0410;
    79: op2_02_in00 = reg_0410;
    83: op2_02_in00 = reg_0410;
    88: op2_02_in00 = reg_0410;
    32: op2_02_in00 = reg_0378;
    35: op2_02_in00 = reg_0378;
    37: op2_02_in00 = reg_0378;
    43: op2_02_in00 = reg_0378;
    58: op2_02_in00 = reg_0378;
    61: op2_02_in00 = reg_0378;
    68: op2_02_in00 = reg_0378;
    71: op2_02_in00 = reg_0378;
    75: op2_02_in00 = reg_0378;
    81: op2_02_in00 = reg_0378;
    86: op2_02_in00 = reg_0378;
    33: op2_02_in00 = reg_0413;
    36: op2_02_in00 = reg_0400;
    42: op2_02_in00 = reg_0400;
    46: op2_02_in00 = reg_0400;
    49: op2_02_in00 = reg_0400;
    57: op2_02_in00 = reg_0400;
    59: op2_02_in00 = reg_0400;
    65: op2_02_in00 = reg_0400;
    66: op2_02_in00 = reg_0400;
    67: op2_02_in00 = reg_0400;
    70: op2_02_in00 = reg_0400;
    73: op2_02_in00 = reg_0400;
    74: op2_02_in00 = reg_0400;
    80: op2_02_in00 = reg_0400;
    82: op2_02_in00 = reg_0400;
    85: op2_02_in00 = reg_0400;
    90: op2_02_in00 = reg_0400;
    91: op2_02_in00 = reg_0400;
    92: op2_02_in00 = reg_0400;
    38: op2_02_in00 = reg_0414;
    39: op2_02_in00 = reg_0412;
    44: op2_02_in00 = reg_0412;
    47: op2_02_in00 = reg_0412;
    52: op2_02_in00 = reg_0412;
    62: op2_02_in00 = reg_0412;
    76: op2_02_in00 = reg_0412;
    84: op2_02_in00 = reg_0412;
    93: op2_02_in00 = reg_0412;
    94: op2_02_in00 = reg_0412;
    95: op2_02_in00 = reg_0412;
    default: op2_02_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の1番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_02_in01 = reg_0775;
    6: op2_02_in01 = reg_0771;
    12: op2_02_in01 = reg_0771;
    7: op2_02_in01 = reg_0774;
    11: op2_02_in01 = reg_0774;
    16: op2_02_in01 = reg_0774;
    8: op2_02_in01 = reg_0772;
    14: op2_02_in01 = reg_0772;
    9: op2_02_in01 = reg_0770;
    10: op2_02_in01 = reg_0025;
    15: op2_02_in01 = reg_0025;
    13: op2_02_in01 = reg_0773;
    17: op2_02_in01 = reg_0773;
    18: op2_02_in01 = reg_0759;
    20: op2_02_in01 = reg_0759;
    19: op2_02_in01 = reg_0762;
    21: op2_02_in01 = reg_0762;
    22: op2_02_in01 = reg_0562;
    23: op2_02_in01 = reg_0764;
    24: op2_02_in01 = reg_0564;
    25: op2_02_in01 = reg_0763;
    26: op2_02_in01 = reg_0565;
    27: op2_02_in01 = reg_0567;
    30: op2_02_in01 = reg_0567;
    28: op2_02_in01 = reg_0566;
    29: op2_02_in01 = reg_0378;
    89: op2_02_in01 = reg_0378;
    31: op2_02_in01 = reg_0411;
    45: op2_02_in01 = reg_0411;
    48: op2_02_in01 = reg_0411;
    50: op2_02_in01 = reg_0411;
    55: op2_02_in01 = reg_0411;
    56: op2_02_in01 = reg_0411;
    63: op2_02_in01 = reg_0411;
    64: op2_02_in01 = reg_0411;
    72: op2_02_in01 = reg_0411;
    79: op2_02_in01 = reg_0411;
    83: op2_02_in01 = reg_0411;
    88: op2_02_in01 = reg_0411;
    32: op2_02_in01 = reg_0400;
    35: op2_02_in01 = reg_0400;
    37: op2_02_in01 = reg_0400;
    43: op2_02_in01 = reg_0400;
    58: op2_02_in01 = reg_0400;
    61: op2_02_in01 = reg_0400;
    68: op2_02_in01 = reg_0400;
    71: op2_02_in01 = reg_0400;
    75: op2_02_in01 = reg_0400;
    81: op2_02_in01 = reg_0400;
    86: op2_02_in01 = reg_0400;
    33: op2_02_in01 = reg_0029;
    34: op2_02_in01 = reg_0412;
    40: op2_02_in01 = reg_0412;
    41: op2_02_in01 = reg_0412;
    51: op2_02_in01 = reg_0412;
    53: op2_02_in01 = reg_0412;
    54: op2_02_in01 = reg_0412;
    69: op2_02_in01 = reg_0412;
    77: op2_02_in01 = reg_0412;
    78: op2_02_in01 = reg_0412;
    87: op2_02_in01 = reg_0412;
    96: op2_02_in01 = reg_0412;
    36: op2_02_in01 = reg_0410;
    42: op2_02_in01 = reg_0410;
    46: op2_02_in01 = reg_0410;
    49: op2_02_in01 = reg_0410;
    57: op2_02_in01 = reg_0410;
    59: op2_02_in01 = reg_0410;
    65: op2_02_in01 = reg_0410;
    66: op2_02_in01 = reg_0410;
    67: op2_02_in01 = reg_0410;
    70: op2_02_in01 = reg_0410;
    73: op2_02_in01 = reg_0410;
    74: op2_02_in01 = reg_0410;
    80: op2_02_in01 = reg_0410;
    82: op2_02_in01 = reg_0410;
    85: op2_02_in01 = reg_0410;
    90: op2_02_in01 = reg_0410;
    91: op2_02_in01 = reg_0410;
    92: op2_02_in01 = reg_0410;
    38: op2_02_in01 = reg_0032;
    39: op2_02_in01 = reg_0413;
    44: op2_02_in01 = reg_0413;
    47: op2_02_in01 = reg_0413;
    52: op2_02_in01 = reg_0413;
    62: op2_02_in01 = reg_0413;
    76: op2_02_in01 = reg_0413;
    84: op2_02_in01 = reg_0413;
    93: op2_02_in01 = reg_0413;
    94: op2_02_in01 = reg_0413;
    95: op2_02_in01 = reg_0413;
    default: op2_02_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の2番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_02_in02 = reg_0776;
    6: op2_02_in02 = reg_0772;
    12: op2_02_in02 = reg_0772;
    7: op2_02_in02 = reg_0775;
    11: op2_02_in02 = reg_0775;
    16: op2_02_in02 = reg_0775;
    8: op2_02_in02 = reg_0773;
    14: op2_02_in02 = reg_0773;
    9: op2_02_in02 = reg_0771;
    10: op2_02_in02 = reg_0777;
    13: op2_02_in02 = reg_0774;
    17: op2_02_in02 = reg_0774;
    15: op2_02_in02 = reg_0043;
    18: op2_02_in02 = reg_0760;
    20: op2_02_in02 = reg_0760;
    22: op2_02_in02 = reg_0760;
    19: op2_02_in02 = reg_0763;
    21: op2_02_in02 = reg_0763;
    23: op2_02_in02 = reg_0025;
    62: op2_02_in02 = reg_0025;
    93: op2_02_in02 = reg_0025;
    94: op2_02_in02 = reg_0025;
    95: op2_02_in02 = reg_0025;
    24: op2_02_in02 = reg_0565;
    25: op2_02_in02 = reg_0764;
    87: op2_02_in02 = reg_0764;
    26: op2_02_in02 = reg_0566;
    27: op2_02_in02 = reg_0574;
    30: op2_02_in02 = reg_0574;
    28: op2_02_in02 = reg_0567;
    31: op2_02_in02 = reg_0567;
    29: op2_02_in02 = reg_0400;
    89: op2_02_in02 = reg_0400;
    32: op2_02_in02 = reg_0410;
    35: op2_02_in02 = reg_0410;
    37: op2_02_in02 = reg_0410;
    43: op2_02_in02 = reg_0410;
    58: op2_02_in02 = reg_0410;
    61: op2_02_in02 = reg_0410;
    68: op2_02_in02 = reg_0410;
    71: op2_02_in02 = reg_0410;
    75: op2_02_in02 = reg_0410;
    81: op2_02_in02 = reg_0410;
    86: op2_02_in02 = reg_0410;
    33: op2_02_in02 = reg_0032;
    34: op2_02_in02 = reg_0413;
    40: op2_02_in02 = reg_0413;
    41: op2_02_in02 = reg_0413;
    51: op2_02_in02 = reg_0413;
    53: op2_02_in02 = reg_0413;
    54: op2_02_in02 = reg_0413;
    69: op2_02_in02 = reg_0413;
    77: op2_02_in02 = reg_0413;
    78: op2_02_in02 = reg_0413;
    96: op2_02_in02 = reg_0413;
    36: op2_02_in02 = reg_0411;
    42: op2_02_in02 = reg_0411;
    46: op2_02_in02 = reg_0411;
    49: op2_02_in02 = reg_0411;
    57: op2_02_in02 = reg_0411;
    59: op2_02_in02 = reg_0411;
    65: op2_02_in02 = reg_0411;
    66: op2_02_in02 = reg_0411;
    67: op2_02_in02 = reg_0411;
    70: op2_02_in02 = reg_0411;
    73: op2_02_in02 = reg_0411;
    74: op2_02_in02 = reg_0411;
    80: op2_02_in02 = reg_0411;
    82: op2_02_in02 = reg_0411;
    85: op2_02_in02 = reg_0411;
    90: op2_02_in02 = reg_0411;
    91: op2_02_in02 = reg_0411;
    92: op2_02_in02 = reg_0411;
    38: op2_02_in02 = reg_0634;
    39: op2_02_in02 = reg_0414;
    44: op2_02_in02 = reg_0414;
    47: op2_02_in02 = reg_0414;
    45: op2_02_in02 = reg_0412;
    48: op2_02_in02 = reg_0412;
    50: op2_02_in02 = reg_0412;
    55: op2_02_in02 = reg_0412;
    56: op2_02_in02 = reg_0412;
    63: op2_02_in02 = reg_0412;
    64: op2_02_in02 = reg_0412;
    72: op2_02_in02 = reg_0412;
    79: op2_02_in02 = reg_0412;
    83: op2_02_in02 = reg_0412;
    88: op2_02_in02 = reg_0412;
    52: op2_02_in02 = reg_0039;
    76: op2_02_in02 = reg_0037;
    84: op2_02_in02 = reg_0037;
    default: op2_02_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の3番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_02_in03 = reg_0777;
    6: op2_02_in03 = reg_0773;
    12: op2_02_in03 = reg_0773;
    7: op2_02_in03 = reg_0776;
    8: op2_02_in03 = reg_0774;
    14: op2_02_in03 = reg_0774;
    9: op2_02_in03 = reg_0772;
    10: op2_02_in03 = reg_0732;
    11: op2_02_in03 = reg_0025;
    16: op2_02_in03 = reg_0025;
    25: op2_02_in03 = reg_0025;
    27: op2_02_in03 = reg_0025;
    69: op2_02_in03 = reg_0025;
    96: op2_02_in03 = reg_0025;
    13: op2_02_in03 = reg_0775;
    17: op2_02_in03 = reg_0775;
    19: op2_02_in03 = reg_0775;
    21: op2_02_in03 = reg_0775;
    15: op2_02_in03 = reg_0020;
    33: op2_02_in03 = reg_0020;
    18: op2_02_in03 = reg_0761;
    20: op2_02_in03 = reg_0761;
    22: op2_02_in03 = reg_0761;
    23: op2_02_in03 = reg_0501;
    24: op2_02_in03 = reg_0762;
    26: op2_02_in03 = reg_0567;
    28: op2_02_in03 = reg_0574;
    31: op2_02_in03 = reg_0574;
    29: op2_02_in03 = reg_0410;
    89: op2_02_in03 = reg_0410;
    30: op2_02_in03 = reg_0765;
    32: op2_02_in03 = reg_0411;
    35: op2_02_in03 = reg_0411;
    37: op2_02_in03 = reg_0411;
    43: op2_02_in03 = reg_0411;
    58: op2_02_in03 = reg_0411;
    61: op2_02_in03 = reg_0411;
    68: op2_02_in03 = reg_0411;
    71: op2_02_in03 = reg_0411;
    75: op2_02_in03 = reg_0411;
    81: op2_02_in03 = reg_0411;
    86: op2_02_in03 = reg_0411;
    34: op2_02_in03 = reg_0414;
    40: op2_02_in03 = reg_0414;
    41: op2_02_in03 = reg_0414;
    36: op2_02_in03 = reg_0412;
    42: op2_02_in03 = reg_0412;
    46: op2_02_in03 = reg_0412;
    49: op2_02_in03 = reg_0412;
    57: op2_02_in03 = reg_0412;
    59: op2_02_in03 = reg_0412;
    65: op2_02_in03 = reg_0412;
    66: op2_02_in03 = reg_0412;
    67: op2_02_in03 = reg_0412;
    70: op2_02_in03 = reg_0412;
    73: op2_02_in03 = reg_0412;
    74: op2_02_in03 = reg_0412;
    80: op2_02_in03 = reg_0412;
    82: op2_02_in03 = reg_0412;
    85: op2_02_in03 = reg_0412;
    90: op2_02_in03 = reg_0412;
    91: op2_02_in03 = reg_0412;
    92: op2_02_in03 = reg_0412;
    38: op2_02_in03 = reg_0021;
    39: op2_02_in03 = reg_0032;
    44: op2_02_in03 = reg_0032;
    47: op2_02_in03 = reg_0032;
    52: op2_02_in03 = reg_0032;
    76: op2_02_in03 = reg_0032;
    84: op2_02_in03 = reg_0032;
    45: op2_02_in03 = reg_0413;
    48: op2_02_in03 = reg_0413;
    50: op2_02_in03 = reg_0413;
    55: op2_02_in03 = reg_0413;
    56: op2_02_in03 = reg_0413;
    63: op2_02_in03 = reg_0413;
    64: op2_02_in03 = reg_0413;
    72: op2_02_in03 = reg_0413;
    79: op2_02_in03 = reg_0413;
    83: op2_02_in03 = reg_0413;
    88: op2_02_in03 = reg_0413;
    51: op2_02_in03 = reg_0039;
    53: op2_02_in03 = reg_0039;
    54: op2_02_in03 = reg_0039;
    62: op2_02_in03 = reg_0037;
    77: op2_02_in03 = reg_0037;
    78: op2_02_in03 = reg_0037;
    87: op2_02_in03 = reg_0037;
    93: op2_02_in03 = reg_0014;
    94: op2_02_in03 = reg_0014;
    95: op2_02_in03 = reg_0014;
    default: op2_02_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の4番目の入力
  always @ ( * ) begin
    case ( state )
    5: op2_02_in04 = reg_0497;
    6: op2_02_in04 = reg_0753;
    8: op2_02_in04 = reg_0775;
    14: op2_02_in04 = reg_0775;
    82: op2_02_in04 = reg_0775;
    9: op2_02_in04 = reg_0773;
    10: op2_02_in04 = reg_0527;
    12: op2_02_in04 = reg_0774;
    13: op2_02_in04 = reg_0025;
    17: op2_02_in04 = reg_0025;
    19: op2_02_in04 = reg_0025;
    63: op2_02_in04 = reg_0025;
    64: op2_02_in04 = reg_0025;
    15: op2_02_in04 = reg_0021;
    33: op2_02_in04 = reg_0021;
    16: op2_02_in04 = reg_0777;
    25: op2_02_in04 = reg_0777;
    18: op2_02_in04 = reg_0763;
    20: op2_02_in04 = reg_0316;
    22: op2_02_in04 = reg_0762;
    23: op2_02_in04 = reg_0340;
    26: op2_02_in04 = reg_0574;
    28: op2_02_in04 = reg_0765;
    29: op2_02_in04 = reg_0603;
    30: op2_02_in04 = reg_0603;
    31: op2_02_in04 = reg_0412;
    32: op2_02_in04 = reg_0412;
    35: op2_02_in04 = reg_0412;
    37: op2_02_in04 = reg_0412;
    43: op2_02_in04 = reg_0412;
    58: op2_02_in04 = reg_0412;
    61: op2_02_in04 = reg_0412;
    71: op2_02_in04 = reg_0412;
    75: op2_02_in04 = reg_0412;
    81: op2_02_in04 = reg_0412;
    86: op2_02_in04 = reg_0412;
    34: op2_02_in04 = reg_0634;
    39: op2_02_in04 = reg_0634;
    44: op2_02_in04 = reg_0634;
    47: op2_02_in04 = reg_0634;
    52: op2_02_in04 = reg_0634;
    36: op2_02_in04 = reg_0413;
    42: op2_02_in04 = reg_0413;
    46: op2_02_in04 = reg_0413;
    49: op2_02_in04 = reg_0413;
    57: op2_02_in04 = reg_0413;
    59: op2_02_in04 = reg_0413;
    65: op2_02_in04 = reg_0413;
    66: op2_02_in04 = reg_0413;
    67: op2_02_in04 = reg_0413;
    70: op2_02_in04 = reg_0413;
    73: op2_02_in04 = reg_0413;
    74: op2_02_in04 = reg_0413;
    80: op2_02_in04 = reg_0413;
    85: op2_02_in04 = reg_0413;
    90: op2_02_in04 = reg_0413;
    91: op2_02_in04 = reg_0413;
    40: op2_02_in04 = reg_0032;
    41: op2_02_in04 = reg_0032;
    53: op2_02_in04 = reg_0032;
    54: op2_02_in04 = reg_0032;
    77: op2_02_in04 = reg_0032;
    45: op2_02_in04 = reg_0414;
    48: op2_02_in04 = reg_0414;
    50: op2_02_in04 = reg_0039;
    55: op2_02_in04 = reg_0039;
    51: op2_02_in04 = reg_0063;
    62: op2_02_in04 = reg_0020;
    76: op2_02_in04 = reg_0020;
    93: op2_02_in04 = reg_0020;
    94: op2_02_in04 = reg_0020;
    95: op2_02_in04 = reg_0020;
    69: op2_02_in04 = reg_0113;
    72: op2_02_in04 = reg_0037;
    83: op2_02_in04 = reg_0037;
    79: op2_02_in04 = reg_0136;
    84: op2_02_in04 = reg_0044;
    87: op2_02_in04 = reg_0501;
    96: op2_02_in04 = reg_0014;
    default: op2_02_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の5番目の入力
  always @ ( * ) begin
    case ( state )
    13: op2_02_in05 = reg_0280;
    25: op2_02_in05 = reg_0567;
    28: op2_02_in05 = reg_0767;
    30: op2_02_in05 = reg_0768;
    32: op2_02_in05 = reg_0414;
    35: op2_02_in05 = reg_0413;
    58: op2_02_in05 = reg_0413;
    40: op2_02_in05 = reg_0634;
    65: op2_02_in05 = reg_0025;
    90: op2_02_in05 = reg_0025;
    91: op2_02_in05 = reg_0025;
    67: op2_02_in05 = reg_0039;
    76: op2_02_in05 = reg_0021;
    95: op2_02_in05 = reg_0021;
    83: op2_02_in05 = reg_0043;
    96: op2_02_in05 = reg_0020;
    default: op2_02_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の6番目の入力
  always @ ( * ) begin
    case ( state )
    58: op2_02_in06 = reg_0039;
    96: op2_02_in06 = reg_0021;
    default: op2_02_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#2のバイアス入力
  always @ ( * ) begin
    case ( state )
    5: op2_02_bias = 64;
    6: op2_02_bias = 66;
    7: op2_02_bias = 55;
    8: op2_02_bias = 68;
    9: op2_02_bias = 84;
    10: op2_02_bias = 57;
    11: op2_02_bias = 59;
    12: op2_02_bias = 85;
    13: op2_02_bias = 84;
    14: op2_02_bias = 79;
    15: op2_02_bias = 70;
    16: op2_02_bias = 84;
    17: op2_02_bias = 83;
    18: op2_02_bias = 79;
    19: op2_02_bias = 78;
    20: op2_02_bias = 61;
    21: op2_02_bias = 62;
    22: op2_02_bias = 71;
    23: op2_02_bias = 48;
    24: op2_02_bias = 73;
    25: op2_02_bias = 93;
    26: op2_02_bias = 65;
    27: op2_02_bias = 61;
    28: op2_02_bias = 84;
    29: op2_02_bias = 70;
    30: op2_02_bias = 69;
    31: op2_02_bias = 63;
    32: op2_02_bias = 76;
    33: op2_02_bias = 68;
    34: op2_02_bias = 69;
    35: op2_02_bias = 83;
    36: op2_02_bias = 69;
    37: op2_02_bias = 71;
    38: op2_02_bias = 63;
    39: op2_02_bias = 56;
    40: op2_02_bias = 87;
    41: op2_02_bias = 73;
    42: op2_02_bias = 62;
    43: op2_02_bias = 70;
    44: op2_02_bias = 69;
    45: op2_02_bias = 75;
    46: op2_02_bias = 70;
    47: op2_02_bias = 78;
    48: op2_02_bias = 56;
    49: op2_02_bias = 63;
    50: op2_02_bias = 79;
    51: op2_02_bias = 71;
    52: op2_02_bias = 66;
    53: op2_02_bias = 70;
    54: op2_02_bias = 78;
    55: op2_02_bias = 67;
    56: op2_02_bias = 45;
    57: op2_02_bias = 70;
    58: op2_02_bias = 85;
    59: op2_02_bias = 64;
    61: op2_02_bias = 66;
    62: op2_02_bias = 71;
    63: op2_02_bias = 70;
    64: op2_02_bias = 64;
    65: op2_02_bias = 80;
    66: op2_02_bias = 72;
    67: op2_02_bias = 86;
    68: op2_02_bias = 50;
    69: op2_02_bias = 74;
    70: op2_02_bias = 61;
    71: op2_02_bias = 65;
    72: op2_02_bias = 67;
    73: op2_02_bias = 63;
    74: op2_02_bias = 62;
    75: op2_02_bias = 63;
    76: op2_02_bias = 64;
    77: op2_02_bias = 72;
    78: op2_02_bias = 69;
    79: op2_02_bias = 73;
    80: op2_02_bias = 67;
    81: op2_02_bias = 80;
    82: op2_02_bias = 69;
    83: op2_02_bias = 97;
    84: op2_02_bias = 60;
    85: op2_02_bias = 78;
    86: op2_02_bias = 56;
    87: op2_02_bias = 61;
    88: op2_02_bias = 66;
    89: op2_02_bias = 51;
    90: op2_02_bias = 86;
    91: op2_02_bias = 69;
    92: op2_02_bias = 54;
    93: op2_02_bias = 68;
    94: op2_02_bias = 68;
    95: op2_02_bias = 83;
    96: op2_02_bias = 76;
    default: op2_02_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#3の0番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_03_in00 = reg_0774;
    9: op2_03_in00 = reg_0774;
    12: op2_03_in00 = reg_0775;
    14: op2_03_in00 = reg_0025;
    59: op2_03_in00 = reg_0025;
    18: op2_03_in00 = reg_0762;
    20: op2_03_in00 = reg_0762;
    22: op2_03_in00 = reg_0763;
    24: op2_03_in00 = reg_0763;
    26: op2_03_in00 = reg_0764;
    29: op2_03_in00 = reg_0566;
    32: op2_03_in00 = reg_0574;
    37: op2_03_in00 = reg_0413;
    43: op2_03_in00 = reg_0413;
    61: op2_03_in00 = reg_0413;
    71: op2_03_in00 = reg_0413;
    75: op2_03_in00 = reg_0413;
    92: op2_03_in00 = reg_0413;
    46: op2_03_in00 = reg_0414;
    68: op2_03_in00 = reg_0412;
    89: op2_03_in00 = reg_0411;
    default: op2_03_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の1番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_03_in01 = reg_0775;
    9: op2_03_in01 = reg_0775;
    12: op2_03_in01 = reg_0025;
    26: op2_03_in01 = reg_0025;
    92: op2_03_in01 = reg_0025;
    14: op2_03_in01 = reg_0777;
    18: op2_03_in01 = reg_0774;
    20: op2_03_in01 = reg_0763;
    22: op2_03_in01 = reg_0764;
    24: op2_03_in01 = reg_0764;
    29: op2_03_in01 = reg_0567;
    32: op2_03_in01 = reg_0029;
    37: op2_03_in01 = reg_0414;
    43: op2_03_in01 = reg_0765;
    46: op2_03_in01 = reg_0063;
    59: op2_03_in01 = reg_0032;
    61: op2_03_in01 = reg_0039;
    68: op2_03_in01 = reg_0413;
    71: op2_03_in01 = reg_0037;
    75: op2_03_in01 = reg_0037;
    89: op2_03_in01 = reg_0412;
    default: op2_03_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の2番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_03_in02 = reg_0776;
    9: op2_03_in02 = reg_0025;
    24: op2_03_in02 = reg_0025;
    68: op2_03_in02 = reg_0025;
    12: op2_03_in02 = reg_0043;
    14: op2_03_in02 = reg_0042;
    18: op2_03_in02 = reg_0775;
    20: op2_03_in02 = reg_0775;
    22: op2_03_in02 = reg_0262;
    26: op2_03_in02 = reg_0777;
    29: op2_03_in02 = reg_0574;
    32: op2_03_in02 = reg_0032;
    37: op2_03_in02 = reg_0032;
    71: op2_03_in02 = reg_0032;
    43: op2_03_in02 = reg_0063;
    46: op2_03_in02 = reg_0767;
    59: op2_03_in02 = reg_0767;
    61: op2_03_in02 = reg_0037;
    75: op2_03_in02 = reg_0415;
    89: op2_03_in02 = reg_0413;
    92: op2_03_in02 = reg_0014;
    default: op2_03_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の3番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_03_in03 = reg_0777;
    9: op2_03_in03 = reg_0777;
    22: op2_03_in03 = reg_0777;
    24: op2_03_in03 = reg_0777;
    12: op2_03_in03 = reg_0044;
    14: op2_03_in03 = reg_0779;
    18: op2_03_in03 = reg_0025;
    20: op2_03_in03 = reg_0025;
    26: op2_03_in03 = reg_0778;
    29: op2_03_in03 = reg_0765;
    32: op2_03_in03 = reg_0020;
    71: op2_03_in03 = reg_0020;
    37: op2_03_in03 = reg_0416;
    43: op2_03_in03 = reg_0634;
    46: op2_03_in03 = reg_0021;
    59: op2_03_in03 = reg_0021;
    61: op2_03_in03 = reg_0034;
    68: op2_03_in03 = reg_0113;
    75: op2_03_in03 = reg_0715;
    89: op2_03_in03 = reg_0029;
    92: op2_03_in03 = reg_0357;
    default: op2_03_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の4番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_03_in04 = reg_0020;
    22: op2_03_in04 = reg_0020;
    9: op2_03_in04 = reg_0525;
    12: op2_03_in04 = reg_0779;
    26: op2_03_in04 = reg_0779;
    14: op2_03_in04 = reg_0760;
    18: op2_03_in04 = reg_0043;
    20: op2_03_in04 = reg_0777;
    29: op2_03_in04 = reg_0777;
    24: op2_03_in04 = reg_0034;
    68: op2_03_in04 = reg_0034;
    32: op2_03_in04 = reg_0021;
    43: op2_03_in04 = reg_0021;
    75: op2_03_in04 = reg_0021;
    37: op2_03_in04 = reg_0417;
    61: op2_03_in04 = reg_0417;
    89: op2_03_in04 = reg_0014;
    default: op2_03_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の5番目の入力
  always @ ( * ) begin
    case ( state )
    6: op2_03_in05 = reg_0021;
    22: op2_03_in05 = reg_0021;
    12: op2_03_in05 = reg_0758;
    24: op2_03_in05 = reg_0366;
    26: op2_03_in05 = reg_0575;
    29: op2_03_in05 = reg_0020;
    32: op2_03_in05 = reg_0415;
    default: op2_03_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の6番目の入力
  always @ ( * ) begin
    case ( state )
    29: op2_03_in06 = reg_0021;
    default: op2_03_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#3のバイアス入力
  always @ ( * ) begin
    case ( state )
    6: op2_03_bias = 86;
    9: op2_03_bias = 73;
    12: op2_03_bias = 94;
    14: op2_03_bias = 65;
    18: op2_03_bias = 83;
    20: op2_03_bias = 70;
    22: op2_03_bias = 92;
    24: op2_03_bias = 85;
    26: op2_03_bias = 87;
    29: op2_03_bias = 107;
    32: op2_03_bias = 78;
    37: op2_03_bias = 72;
    43: op2_03_bias = 60;
    46: op2_03_bias = 64;
    59: op2_03_bias = 54;
    61: op2_03_bias = 70;
    68: op2_03_bias = 84;
    71: op2_03_bias = 51;
    75: op2_03_bias = 72;
    89: op2_03_bias = 65;
    92: op2_03_bias = 53;
    default: op2_03_bias = 0;
    endcase
  end // always @ ( * )

  // REG#0の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0000 <= imem03_in[3:0];
    5: reg_0000 <= imem03_in[3:0];
    88: reg_0000 <= imem03_in[3:0];
    90: reg_0000 <= imem00_in[55:52];
    94: reg_0000 <= imem01_in[107:104];
    endcase
  end

  // REG#1の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0001 <= imem03_in[23:20];
    5: reg_0001 <= imem03_in[23:20];
    89: reg_0001 <= imem03_in[23:20];
    endcase
  end

  // REG#2の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0002 <= imem03_in[27:24];
    5: reg_0002 <= imem03_in[27:24];
    89: reg_0002 <= imem03_in[27:24];
    endcase
  end

  // REG#3の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0003 <= imem03_in[35:32];
    5: reg_0003 <= imem03_in[35:32];
    87: reg_0003 <= imem03_in[35:32];
    endcase
  end

  // REG#4の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0004 <= imem03_in[115:112];
    5: reg_0004 <= imem03_in[115:112];
    89: reg_0004 <= imem03_in[115:112];
    endcase
  end

  // REG#5の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0005 <= imem06_in[103:100];
    4: reg_0005 <= op1_00_out;
    5: reg_0005 <= op1_00_out;
    6: reg_0005 <= op1_00_out;
    8: reg_0005 <= imem06_in[103:100];
    30: reg_0005 <= imem06_in[103:100];
    31: reg_0005 <= op1_00_out;
    32: reg_0005 <= op1_00_out;
    33: reg_0005 <= op1_00_out;
    34: reg_0005 <= op1_00_out;
    35: reg_0005 <= op1_00_out;
    36: reg_0005 <= op1_00_out;
    37: reg_0005 <= op1_00_out;
    38: reg_0005 <= op1_00_out;
    39: reg_0005 <= op1_00_out;
    40: reg_0005 <= op1_00_out;
    41: reg_0005 <= op1_00_out;
    42: reg_0005 <= op1_00_out;
    43: reg_0005 <= op1_00_out;
    44: reg_0005 <= op1_00_out;
    45: reg_0005 <= op1_00_out;
    46: reg_0005 <= op1_00_out;
    47: reg_0005 <= op1_00_out;
    48: reg_0005 <= op1_00_out;
    49: reg_0005 <= op1_00_out;
    50: reg_0005 <= op1_00_out;
    51: reg_0005 <= op1_00_out;
    52: reg_0005 <= op1_00_out;
    53: reg_0005 <= op1_00_out;
    54: reg_0005 <= op1_00_out;
    55: reg_0005 <= op1_00_out;
    56: reg_0005 <= op1_00_out;
    57: reg_0005 <= op1_00_out;
    59: reg_0005 <= imem06_in[103:100];
    60: reg_0005 <= op1_00_out;
    61: reg_0005 <= op1_00_out;
    62: reg_0005 <= op1_00_out;
    63: reg_0005 <= op1_00_out;
    64: reg_0005 <= op1_00_out;
    65: reg_0005 <= op1_00_out;
    66: reg_0005 <= op1_00_out;
    67: reg_0005 <= op1_00_out;
    68: reg_0005 <= op1_00_out;
    69: reg_0005 <= op1_00_out;
    70: reg_0005 <= op1_00_out;
    71: reg_0005 <= op1_00_out;
    72: reg_0005 <= op1_00_out;
    73: reg_0005 <= op1_00_out;
    74: reg_0005 <= op1_00_out;
    75: reg_0005 <= op1_00_out;
    76: reg_0005 <= op1_00_out;
    77: reg_0005 <= op1_00_out;
    78: reg_0005 <= op1_00_out;
    79: reg_0005 <= op1_00_out;
    80: reg_0005 <= op1_00_out;
    81: reg_0005 <= op1_00_out;
    82: reg_0005 <= op1_00_out;
    83: reg_0005 <= op1_00_out;
    84: reg_0005 <= op1_00_out;
    85: reg_0005 <= op1_00_out;
    86: reg_0005 <= op1_00_out;
    87: reg_0005 <= op1_00_out;
    88: reg_0005 <= op1_00_out;
    89: reg_0005 <= op1_00_out;
    90: reg_0005 <= op1_00_out;
    91: reg_0005 <= op1_00_out;
    92: reg_0005 <= op1_00_out;
    93: reg_0005 <= op1_00_out;
    94: reg_0005 <= op1_00_out;
    95: reg_0005 <= op1_00_out;
    96: reg_0005 <= op1_00_out;
    endcase
  end

  // REG#6の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0006 <= imem03_in[7:4];
    5: reg_0006 <= imem03_in[7:4];
    88: reg_0006 <= imem03_in[119:116];
    90: reg_0006 <= imem00_in[7:4];
    endcase
  end

  // REG#7の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0007 <= imem03_in[47:44];
    5: reg_0007 <= imem03_in[47:44];
    89: reg_0007 <= imem03_in[47:44];
    92: reg_0007 <= imem01_in[63:60];
    94: reg_0007 <= imem01_in[63:60];
    endcase
  end

  // REG#8の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0008 <= imem03_in[75:72];
    5: reg_0008 <= imem03_in[75:72];
    85: reg_0008 <= imem05_in[99:96];
    87: reg_0008 <= imem03_in[75:72];
    endcase
  end

  // REG#9の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0009 <= imem03_in[103:100];
    5: reg_0009 <= imem03_in[103:100];
    87: reg_0009 <= imem03_in[103:100];
    endcase
  end

  // REG#10の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0010 <= imem03_in[107:104];
    5: reg_0010 <= imem03_in[107:104];
    85: reg_0010 <= imem05_in[7:4];
    87: reg_0010 <= imem03_in[107:104];
    endcase
  end

  // REG#11の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0011 <= imem06_in[107:104];
    4: reg_0011 <= op1_01_out;
    5: reg_0011 <= op1_01_out;
    6: reg_0011 <= op1_01_out;
    7: reg_0011 <= op1_01_out;
    8: reg_0011 <= op1_01_out;
    9: reg_0011 <= op1_01_out;
    10: reg_0011 <= op1_01_out;
    11: reg_0011 <= op1_01_out;
    12: reg_0011 <= op1_01_out;
    13: reg_0011 <= op1_01_out;
    14: reg_0011 <= op1_01_out;
    15: reg_0011 <= op1_01_out;
    16: reg_0011 <= op1_01_out;
    17: reg_0011 <= op1_01_out;
    18: reg_0011 <= op1_01_out;
    19: reg_0011 <= op1_01_out;
    20: reg_0011 <= op1_01_out;
    21: reg_0011 <= op1_01_out;
    22: reg_0011 <= op1_01_out;
    23: reg_0011 <= op1_01_out;
    24: reg_0011 <= op1_01_out;
    25: reg_0011 <= op1_01_out;
    26: reg_0011 <= op1_01_out;
    27: reg_0011 <= op1_01_out;
    28: reg_0011 <= op1_01_out;
    29: reg_0011 <= op1_01_out;
    30: reg_0011 <= op1_01_out;
    31: reg_0011 <= op1_01_out;
    32: reg_0011 <= op1_01_out;
    33: reg_0011 <= op1_01_out;
    34: reg_0011 <= op1_01_out;
    35: reg_0011 <= op1_01_out;
    36: reg_0011 <= op1_01_out;
    37: reg_0011 <= op1_01_out;
    38: reg_0011 <= op1_01_out;
    39: reg_0011 <= op1_01_out;
    40: reg_0011 <= op1_01_out;
    41: reg_0011 <= op1_01_out;
    42: reg_0011 <= op1_01_out;
    43: reg_0011 <= op1_01_out;
    44: reg_0011 <= op1_01_out;
    45: reg_0011 <= op1_01_out;
    46: reg_0011 <= op1_01_out;
    47: reg_0011 <= op1_01_out;
    48: reg_0011 <= op1_01_out;
    49: reg_0011 <= op1_01_out;
    50: reg_0011 <= op1_01_out;
    51: reg_0011 <= op1_01_out;
    52: reg_0011 <= op1_01_out;
    53: reg_0011 <= op1_01_out;
    54: reg_0011 <= op1_01_out;
    55: reg_0011 <= op1_01_out;
    56: reg_0011 <= op1_01_out;
    57: reg_0011 <= op1_01_out;
    58: reg_0011 <= op1_01_out;
    59: reg_0011 <= op1_01_out;
    60: reg_0011 <= op1_01_out;
    61: reg_0011 <= op1_01_out;
    62: reg_0011 <= op1_01_out;
    63: reg_0011 <= op1_01_out;
    64: reg_0011 <= op1_01_out;
    65: reg_0011 <= op1_01_out;
    66: reg_0011 <= op1_01_out;
    67: reg_0011 <= op1_01_out;
    68: reg_0011 <= op1_01_out;
    70: reg_0011 <= imem06_in[107:104];
    87: reg_0011 <= imem06_in[107:104];
    88: reg_0011 <= op1_01_out;
    89: reg_0011 <= op1_01_out;
    90: reg_0011 <= op1_01_out;
    91: reg_0011 <= op1_01_out;
    92: reg_0011 <= op1_01_out;
    93: reg_0011 <= op1_01_out;
    94: reg_0011 <= op1_01_out;
    95: reg_0011 <= op1_01_out;
    96: reg_0011 <= op1_01_out;
    endcase
  end

  // REG#12の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0012 <= imem03_in[19:16];
    5: reg_0012 <= imem03_in[19:16];
    87: reg_0012 <= imem03_in[19:16];
    endcase
  end

  // REG#13の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0013 <= imem03_in[43:40];
    5: reg_0013 <= imem03_in[43:40];
    89: reg_0013 <= imem03_in[43:40];
    93: reg_0013 <= imem01_in[11:8];
    95: reg_0013 <= imem01_in[11:8];
    endcase
  end

  // REG#14の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0014 <= imem03_in[67:64];
    5: reg_0014 <= imem03_in[67:64];
    88: reg_0014 <= op1_13_out;
    89: reg_0014 <= op1_13_out;
    91: reg_0014 <= op1_13_out;
    92: reg_0014 <= op1_13_out;
    93: reg_0014 <= op1_13_out;
    94: reg_0014 <= op1_13_out;
    95: reg_0014 <= op1_13_out;
    endcase
  end

  // REG#15の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0015 <= imem03_in[83:80];
    5: reg_0015 <= imem03_in[83:80];
    85: reg_0015 <= imem05_in[23:20];
    87: reg_0015 <= imem03_in[83:80];
    endcase
  end

  // REG#16の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0016 <= imem03_in[91:88];
    5: reg_0016 <= imem03_in[91:88];
    88: reg_0016 <= imem03_in[91:88];
    90: reg_0016 <= imem00_in[99:96];
    endcase
  end

  // REG#17の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0017 <= imem06_in[55:52];
    4: reg_0017 <= op1_02_out;
    5: reg_0017 <= op1_02_out;
    6: reg_0017 <= op1_02_out;
    7: reg_0017 <= op1_02_out;
    8: reg_0017 <= op1_02_out;
    9: reg_0017 <= op1_02_out;
    10: reg_0017 <= op1_02_out;
    11: reg_0017 <= op1_02_out;
    12: reg_0017 <= op1_02_out;
    13: reg_0017 <= op1_02_out;
    14: reg_0017 <= op1_02_out;
    15: reg_0017 <= op1_02_out;
    16: reg_0017 <= op1_02_out;
    17: reg_0017 <= op1_02_out;
    18: reg_0017 <= op1_02_out;
    19: reg_0017 <= op1_02_out;
    20: reg_0017 <= op1_02_out;
    21: reg_0017 <= op1_02_out;
    22: reg_0017 <= op1_02_out;
    23: reg_0017 <= op1_02_out;
    24: reg_0017 <= op1_02_out;
    25: reg_0017 <= op1_02_out;
    26: reg_0017 <= op1_02_out;
    27: reg_0017 <= op1_02_out;
    28: reg_0017 <= op1_02_out;
    29: reg_0017 <= op1_02_out;
    30: reg_0017 <= op1_02_out;
    31: reg_0017 <= op1_02_out;
    32: reg_0017 <= op1_02_out;
    33: reg_0017 <= op1_02_out;
    34: reg_0017 <= op1_02_out;
    35: reg_0017 <= op1_02_out;
    36: reg_0017 <= op1_02_out;
    37: reg_0017 <= op1_02_out;
    38: reg_0017 <= op1_02_out;
    39: reg_0017 <= op1_02_out;
    40: reg_0017 <= op1_02_out;
    41: reg_0017 <= op1_02_out;
    42: reg_0017 <= op1_02_out;
    43: reg_0017 <= op1_02_out;
    44: reg_0017 <= op1_02_out;
    45: reg_0017 <= op1_02_out;
    46: reg_0017 <= op1_02_out;
    47: reg_0017 <= op1_02_out;
    48: reg_0017 <= op1_02_out;
    49: reg_0017 <= op1_02_out;
    50: reg_0017 <= op1_02_out;
    51: reg_0017 <= op1_02_out;
    52: reg_0017 <= op1_02_out;
    53: reg_0017 <= op1_02_out;
    54: reg_0017 <= op1_02_out;
    55: reg_0017 <= op1_02_out;
    56: reg_0017 <= op1_02_out;
    57: reg_0017 <= op1_02_out;
    58: reg_0017 <= op1_02_out;
    59: reg_0017 <= op1_02_out;
    60: reg_0017 <= op1_02_out;
    61: reg_0017 <= op1_02_out;
    62: reg_0017 <= op1_02_out;
    63: reg_0017 <= op1_02_out;
    64: reg_0017 <= op1_02_out;
    65: reg_0017 <= op1_02_out;
    66: reg_0017 <= op1_02_out;
    67: reg_0017 <= op1_02_out;
    68: reg_0017 <= op1_02_out;
    69: reg_0017 <= op1_02_out;
    70: reg_0017 <= op1_02_out;
    71: reg_0017 <= op1_02_out;
    72: reg_0017 <= op1_02_out;
    73: reg_0017 <= op1_02_out;
    74: reg_0017 <= op1_02_out;
    75: reg_0017 <= op1_02_out;
    76: reg_0017 <= op1_02_out;
    77: reg_0017 <= op1_02_out;
    78: reg_0017 <= op1_02_out;
    79: reg_0017 <= op1_02_out;
    80: reg_0017 <= op1_02_out;
    81: reg_0017 <= op1_02_out;
    82: reg_0017 <= op1_02_out;
    83: reg_0017 <= op1_02_out;
    84: reg_0017 <= op1_02_out;
    85: reg_0017 <= op1_02_out;
    86: reg_0017 <= op1_02_out;
    87: reg_0017 <= op1_02_out;
    88: reg_0017 <= op1_02_out;
    89: reg_0017 <= op1_02_out;
    90: reg_0017 <= op1_02_out;
    91: reg_0017 <= op1_02_out;
    92: reg_0017 <= op1_02_out;
    93: reg_0017 <= op1_02_out;
    94: reg_0017 <= op1_02_out;
    95: reg_0017 <= op1_02_out;
    96: reg_0017 <= op1_02_out;
    endcase
  end

  // REG#18の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0018 <= imem06_in[75:72];
    4: reg_0018 <= op1_03_out;
    5: reg_0018 <= op1_03_out;
    6: reg_0018 <= op1_03_out;
    7: reg_0018 <= op1_03_out;
    8: reg_0018 <= op1_03_out;
    9: reg_0018 <= op1_03_out;
    10: reg_0018 <= op1_03_out;
    11: reg_0018 <= op1_03_out;
    12: reg_0018 <= op1_03_out;
    13: reg_0018 <= op1_03_out;
    14: reg_0018 <= op1_03_out;
    15: reg_0018 <= op1_03_out;
    16: reg_0018 <= op1_03_out;
    17: reg_0018 <= op1_03_out;
    18: reg_0018 <= op1_03_out;
    19: reg_0018 <= op1_03_out;
    20: reg_0018 <= op1_03_out;
    21: reg_0018 <= op1_03_out;
    22: reg_0018 <= op1_03_out;
    23: reg_0018 <= op1_03_out;
    24: reg_0018 <= op1_03_out;
    25: reg_0018 <= op1_03_out;
    26: reg_0018 <= op1_03_out;
    27: reg_0018 <= op1_03_out;
    28: reg_0018 <= op1_03_out;
    29: reg_0018 <= op1_03_out;
    30: reg_0018 <= op1_03_out;
    31: reg_0018 <= op1_03_out;
    32: reg_0018 <= op1_03_out;
    33: reg_0018 <= op1_03_out;
    34: reg_0018 <= op1_03_out;
    35: reg_0018 <= op1_03_out;
    36: reg_0018 <= op1_03_out;
    37: reg_0018 <= op1_03_out;
    38: reg_0018 <= op1_03_out;
    39: reg_0018 <= op1_03_out;
    40: reg_0018 <= op1_03_out;
    41: reg_0018 <= op1_03_out;
    42: reg_0018 <= op1_03_out;
    43: reg_0018 <= op1_03_out;
    44: reg_0018 <= op1_03_out;
    45: reg_0018 <= op1_03_out;
    46: reg_0018 <= op1_03_out;
    47: reg_0018 <= op1_03_out;
    48: reg_0018 <= op1_03_out;
    49: reg_0018 <= op1_03_out;
    50: reg_0018 <= op1_03_out;
    51: reg_0018 <= op1_03_out;
    52: reg_0018 <= op1_03_out;
    53: reg_0018 <= op1_03_out;
    54: reg_0018 <= op1_03_out;
    55: reg_0018 <= op1_03_out;
    56: reg_0018 <= op1_03_out;
    57: reg_0018 <= op1_03_out;
    58: reg_0018 <= op1_03_out;
    59: reg_0018 <= op1_03_out;
    60: reg_0018 <= op1_03_out;
    61: reg_0018 <= op1_03_out;
    62: reg_0018 <= op1_03_out;
    63: reg_0018 <= op1_03_out;
    64: reg_0018 <= op1_03_out;
    65: reg_0018 <= op1_03_out;
    66: reg_0018 <= op1_03_out;
    67: reg_0018 <= op1_03_out;
    68: reg_0018 <= op1_03_out;
    69: reg_0018 <= op1_03_out;
    70: reg_0018 <= op1_03_out;
    71: reg_0018 <= op1_03_out;
    72: reg_0018 <= op1_03_out;
    73: reg_0018 <= op1_03_out;
    74: reg_0018 <= op1_03_out;
    75: reg_0018 <= op1_03_out;
    76: reg_0018 <= op1_03_out;
    77: reg_0018 <= op1_03_out;
    78: reg_0018 <= op1_03_out;
    79: reg_0018 <= op1_03_out;
    80: reg_0018 <= op1_03_out;
    81: reg_0018 <= op1_03_out;
    82: reg_0018 <= op1_03_out;
    83: reg_0018 <= op1_03_out;
    84: reg_0018 <= op1_03_out;
    85: reg_0018 <= op1_03_out;
    86: reg_0018 <= op1_03_out;
    87: reg_0018 <= op1_03_out;
    88: reg_0018 <= op1_03_out;
    89: reg_0018 <= op1_03_out;
    90: reg_0018 <= op1_03_out;
    91: reg_0018 <= op1_03_out;
    92: reg_0018 <= op1_03_out;
    93: reg_0018 <= op1_03_out;
    94: reg_0018 <= op1_03_out;
    95: reg_0018 <= op1_03_out;
    96: reg_0018 <= op1_03_out;
    endcase
  end

  // REG#19の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0019 <= imem03_in[11:8];
    5: reg_0019 <= imem03_in[11:8];
    89: reg_0019 <= imem00_in[15:12];
    91: reg_0019 <= imem01_in[99:96];
    93: reg_0019 <= imem01_in[35:32];
    95: reg_0019 <= imem01_in[35:32];
    endcase
  end

  // REG#20の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0020 <= imem06_in[59:56];
    5: reg_0020 <= op1_14_out;
    7: reg_0020 <= imem06_in[59:56];
    8: reg_0020 <= op1_14_out;
    10: reg_0020 <= op1_14_out;
    12: reg_0020 <= op1_14_out;
    14: reg_0020 <= op1_14_out;
    15: reg_0020 <= op1_14_out;
    17: reg_0020 <= op1_14_out;
    19: reg_0020 <= op1_14_out;
    21: reg_0020 <= op1_14_out;
    22: reg_0020 <= op1_14_out;
    24: reg_0020 <= op1_14_out;
    27: reg_0020 <= imem06_in[59:56];
    28: reg_0020 <= op1_14_out;
    29: reg_0020 <= op1_14_out;
    31: reg_0020 <= op1_14_out;
    32: reg_0020 <= op1_14_out;
    33: reg_0020 <= op1_14_out;
    35: reg_0020 <= op1_14_out;
    38: reg_0020 <= imem06_in[59:56];
    55: reg_0020 <= imem06_in[59:56];
    57: reg_0020 <= op1_14_out;
    59: reg_0020 <= op1_14_out;
    61: reg_0020 <= op1_14_out;
    62: reg_0020 <= op1_14_out;
    64: reg_0020 <= op1_14_out;
    66: reg_0020 <= op1_14_out;
    68: reg_0020 <= op1_14_out;
    70: reg_0020 <= op1_14_out;
    71: reg_0020 <= op1_14_out;
    73: reg_0020 <= op1_14_out;
    75: reg_0020 <= op1_14_out;
    76: reg_0020 <= op1_14_out;
    78: reg_0020 <= op1_14_out;
    80: reg_0020 <= op1_14_out;
    82: reg_0020 <= op1_14_out;
    84: reg_0020 <= op1_14_out;
    86: reg_0020 <= op1_14_out;
    88: reg_0020 <= op1_14_out;
    90: reg_0020 <= op1_14_out;
    92: reg_0020 <= op1_14_out;
    93: reg_0020 <= op1_14_out;
    94: reg_0020 <= op1_14_out;
    95: reg_0020 <= op1_14_out;
    endcase
  end

  // REG#21の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0021 <= imem06_in[83:80];
    5: reg_0021 <= op1_15_out;
    6: reg_0021 <= op1_15_out;
    8: reg_0021 <= op1_15_out;
    10: reg_0021 <= op1_15_out;
    12: reg_0021 <= op1_15_out;
    14: reg_0021 <= op1_15_out;
    15: reg_0021 <= op1_15_out;
    17: reg_0021 <= op1_15_out;
    19: reg_0021 <= op1_15_out;
    21: reg_0021 <= op1_15_out;
    22: reg_0021 <= op1_15_out;
    24: reg_0021 <= op1_15_out;
    26: reg_0021 <= op1_15_out;
    28: reg_0021 <= op1_15_out;
    29: reg_0021 <= op1_15_out;
    31: reg_0021 <= op1_15_out;
    32: reg_0021 <= op1_15_out;
    33: reg_0021 <= op1_15_out;
    35: reg_0021 <= op1_15_out;
    37: reg_0021 <= op1_15_out;
    38: reg_0021 <= op1_15_out;
    40: reg_0021 <= op1_15_out;
    42: reg_0021 <= op1_15_out;
    43: reg_0021 <= op1_15_out;
    45: reg_0021 <= op1_15_out;
    46: reg_0021 <= op1_15_out;
    48: reg_0021 <= op1_15_out;
    50: reg_0021 <= op1_15_out;
    52: reg_0021 <= op1_15_out;
    54: reg_0021 <= op1_15_out;
    56: reg_0021 <= op1_15_out;
    58: reg_0021 <= op1_15_out;
    60: reg_0021 <= imem06_in[83:80];
    66: reg_0021 <= op1_15_out;
    69: reg_0021 <= imem06_in[83:80];
    70: reg_0021 <= op1_15_out;
    72: reg_0021 <= op1_15_out;
    74: reg_0021 <= op1_15_out;
    75: reg_0021 <= op1_15_out;
    76: reg_0021 <= op1_15_out;
    78: reg_0021 <= op1_15_out;
    80: reg_0021 <= op1_15_out;
    82: reg_0021 <= op1_15_out;
    84: reg_0021 <= op1_15_out;
    86: reg_0021 <= op1_15_out;
    88: reg_0021 <= op1_15_out;
    90: reg_0021 <= op1_15_out;
    92: reg_0021 <= op1_15_out;
    94: reg_0021 <= op1_15_out;
    95: reg_0021 <= op1_15_out;
    endcase
  end

  // REG#22の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0022 <= imem06_in[99:96];
    5: reg_0022 <= op2_00_out;
    6: reg_0022 <= op2_00_out;
    9: reg_0022 <= op2_00_out;
    19: reg_0022 <= op2_00_out;
    53: reg_0022 <= op2_00_out;
    80: reg_0022 <= op2_00_out;
    83: reg_0022 <= op2_00_out;
    92: reg_0022 <= op2_00_out;
    endcase
  end

  // REG#23の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0023 <= imem06_in[115:112];
    5: reg_0023 <= op2_01_out;
    7: reg_0023 <= op2_01_out;
    14: reg_0023 <= op2_01_out;
    37: reg_0023 <= op2_01_out;
    71: reg_0023 <= op2_01_out;
    96: reg_0023 <= op2_01_out;
    endcase
  end

  // REG#24の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0024 <= imem06_in[87:84];
    5: reg_0024 <= op2_02_out;
    8: reg_0024 <= op2_02_out;
    18: reg_0024 <= op2_02_out;
    51: reg_0024 <= op2_02_out;
    76: reg_0024 <= op2_02_out;
    endcase
  end

  // REG#25の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0025 <= imem06_in[67:64];
    7: reg_0025 <= imem06_in[15:12];
    8: reg_0025 <= op1_12_out;
    9: reg_0025 <= op1_12_out;
    10: reg_0025 <= op1_12_out;
    11: reg_0025 <= op1_12_out;
    12: reg_0025 <= op1_12_out;
    13: reg_0025 <= op1_12_out;
    14: reg_0025 <= op1_12_out;
    15: reg_0025 <= op1_12_out;
    16: reg_0025 <= op1_12_out;
    17: reg_0025 <= op1_12_out;
    18: reg_0025 <= op1_12_out;
    19: reg_0025 <= op1_12_out;
    20: reg_0025 <= op1_12_out;
    22: reg_0025 <= op1_12_out;
    23: reg_0025 <= op1_12_out;
    24: reg_0025 <= op1_12_out;
    25: reg_0025 <= op1_12_out;
    26: reg_0025 <= op1_12_out;
    28: reg_0025 <= imem06_in[15:12];
    56: reg_0025 <= op1_12_out;
    58: reg_0025 <= op1_12_out;
    59: reg_0025 <= op1_12_out;
    61: reg_0025 <= op1_12_out;
    62: reg_0025 <= op1_12_out;
    63: reg_0025 <= op1_12_out;
    64: reg_0025 <= op1_12_out;
    65: reg_0025 <= op1_12_out;
    67: reg_0025 <= op1_12_out;
    68: reg_0025 <= op1_12_out;
    70: reg_0025 <= imem06_in[15:12];
    87: reg_0025 <= op1_12_out;
    89: reg_0025 <= op1_12_out;
    90: reg_0025 <= op1_12_out;
    91: reg_0025 <= op1_12_out;
    92: reg_0025 <= op1_12_out;
    93: reg_0025 <= op1_12_out;
    94: reg_0025 <= op1_12_out;
    95: reg_0025 <= op1_12_out;
    endcase
  end

  // REG#26の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0026 <= imem06_in[23:20];
    7: reg_0026 <= imem06_in[23:20];
    8: reg_0026 <= op2_00_out;
    16: reg_0026 <= op2_00_out;
    43: reg_0026 <= op2_00_out;
    48: reg_0026 <= op2_00_out;
    65: reg_0026 <= op2_00_out;
    76: reg_0026 <= op2_00_out;
    endcase
  end

  // REG#27の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0027 <= imem06_in[19:16];
    7: reg_0027 <= imem06_in[27:24];
    8: reg_0027 <= op2_01_out;
    17: reg_0027 <= op2_01_out;
    47: reg_0027 <= op2_01_out;
    63: reg_0027 <= op2_01_out;
    72: reg_0027 <= imem05_in[95:92];
    92: reg_0027 <= op2_01_out;
    endcase
  end

  // REG#28の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0028 <= imem06_in[7:4];
    8: reg_0028 <= imem06_in[7:4];
    29: reg_0028 <= imem03_in[15:12];
    31: reg_0028 <= imem06_in[7:4];
    36: reg_0028 <= imem06_in[7:4];
    60: reg_0028 <= imem06_in[7:4];
    67: reg_0028 <= imem01_in[15:12];
    69: reg_0028 <= imem03_in[15:12];
    endcase
  end

  // REG#29の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0029 <= imem06_in[95:92];
    8: reg_0029 <= imem06_in[95:92];
    30: reg_0029 <= imem06_in[7:4];
    31: reg_0029 <= op1_12_out;
    32: reg_0029 <= op1_12_out;
    34: reg_0029 <= imem06_in[7:4];
    36: reg_0029 <= imem06_in[95:92];
    60: reg_0029 <= imem06_in[95:92];
    70: reg_0029 <= imem06_in[7:4];
    87: reg_0029 <= imem06_in[7:4];
    88: reg_0029 <= op1_12_out;
    90: reg_0029 <= imem00_in[123:120];
    endcase
  end

  // REG#30の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0030 <= imem06_in[91:88];
    8: reg_0030 <= imem06_in[91:88];
    31: reg_0030 <= imem06_in[91:88];
    32: reg_0030 <= op2_00_out;
    54: reg_0030 <= op2_00_out;
    84: reg_0030 <= imem02_in[3:0];
    94: reg_0030 <= op2_00_out;
    endcase
  end

  // REG#31の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0031 <= imem06_in[15:12];
    8: reg_0031 <= imem06_in[15:12];
    31: reg_0031 <= imem06_in[15:12];
    34: reg_0031 <= imem06_in[15:12];
    36: reg_0031 <= imem06_in[15:12];
    55: reg_0031 <= imem06_in[115:112];
    57: reg_0031 <= imem06_in[15:12];
    83: reg_0031 <= imem02_in[43:40];
    endcase
  end

  // REG#32の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0032 <= imem06_in[35:32];
    8: reg_0032 <= imem06_in[35:32];
    30: reg_0032 <= imem06_in[15:12];
    31: reg_0032 <= op1_13_out;
    32: reg_0032 <= op1_13_out;
    34: reg_0032 <= imem06_in[35:32];
    36: reg_0032 <= op1_13_out;
    37: reg_0032 <= op1_13_out;
    38: reg_0032 <= op1_13_out;
    39: reg_0032 <= op1_13_out;
    40: reg_0032 <= op1_13_out;
    41: reg_0032 <= op1_13_out;
    43: reg_0032 <= op1_13_out;
    44: reg_0032 <= op1_13_out;
    46: reg_0032 <= op1_13_out;
    47: reg_0032 <= op1_13_out;
    49: reg_0032 <= op1_13_out;
    51: reg_0032 <= op1_13_out;
    52: reg_0032 <= op1_13_out;
    53: reg_0032 <= op1_13_out;
    54: reg_0032 <= op1_13_out;
    56: reg_0032 <= op1_13_out;
    58: reg_0032 <= op1_13_out;
    60: reg_0032 <= imem06_in[35:32];
    66: reg_0032 <= op1_13_out;
    69: reg_0032 <= imem06_in[35:32];
    70: reg_0032 <= op1_13_out;
    71: reg_0032 <= op1_13_out;
    73: reg_0032 <= op1_13_out;
    75: reg_0032 <= op1_13_out;
    76: reg_0032 <= op1_13_out;
    77: reg_0032 <= op1_13_out;
    79: reg_0032 <= op1_13_out;
    81: reg_0032 <= op1_13_out;
    83: reg_0032 <= op1_13_out;
    85: reg_0032 <= imem06_in[15:12];
    endcase
  end

  // REG#33の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0033 <= imem06_in[3:0];
    8: reg_0033 <= imem06_in[3:0];
    30: reg_0033 <= imem06_in[75:72];
    31: reg_0033 <= op2_01_out;
    52: reg_0033 <= op2_01_out;
    78: reg_0033 <= op2_01_out;
    endcase
  end

  // REG#34の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0034 <= imem06_in[39:36];
    8: reg_0034 <= imem06_in[39:36];
    23: reg_0034 <= op1_14_out;
    24: reg_0034 <= op2_02_out;
    29: reg_0034 <= op2_02_out;
    46: reg_0034 <= op2_02_out;
    60: reg_0034 <= op1_14_out;
    61: reg_0034 <= op2_02_out;
    65: reg_0034 <= op1_14_out;
    67: reg_0034 <= op1_14_out;
    69: reg_0034 <= imem06_in[39:36];
    70: reg_0034 <= op2_02_out;
    94: reg_0034 <= op2_02_out;
    endcase
  end

  // REG#35の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0035 <= imem06_in[43:40];
    8: reg_0035 <= imem06_in[43:40];
    30: reg_0035 <= imem06_in[111:108];
    32: reg_0035 <= op2_02_out;
    57: reg_0035 <= imem06_in[111:108];
    82: reg_0035 <= op2_02_out;
    91: reg_0035 <= op2_02_out;
    endcase
  end

  // REG#36の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0036 <= imem06_in[71:68];
    8: reg_0036 <= imem06_in[71:68];
    29: reg_0036 <= op2_01_out;
    45: reg_0036 <= op2_01_out;
    56: reg_0036 <= op2_01_out;
    90: reg_0036 <= op2_01_out;
    endcase
  end

  // REG#37の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0037 <= imem06_in[79:76];
    8: reg_0037 <= imem06_in[79:76];
    30: reg_0037 <= imem06_in[79:76];
    34: reg_0037 <= imem06_in[79:76];
    36: reg_0037 <= imem06_in[79:76];
    59: reg_0037 <= imem06_in[79:76];
    60: reg_0037 <= op1_13_out;
    61: reg_0037 <= op1_13_out;
    62: reg_0037 <= op1_13_out;
    64: reg_0037 <= op1_13_out;
    67: reg_0037 <= imem01_in[55:52];
    69: reg_0037 <= imem06_in[79:76];
    70: reg_0037 <= op1_12_out;
    71: reg_0037 <= op1_12_out;
    72: reg_0037 <= op1_12_out;
    74: reg_0037 <= op1_12_out;
    75: reg_0037 <= op1_12_out;
    76: reg_0037 <= op1_12_out;
    77: reg_0037 <= op1_12_out;
    78: reg_0037 <= op1_13_out;
    80: reg_0037 <= op1_12_out;
    82: reg_0037 <= op1_12_out;
    83: reg_0037 <= op1_12_out;
    84: reg_0037 <= op1_12_out;
    86: reg_0037 <= op1_12_out;
    88: reg_0037 <= imem06_in[79:76];
    endcase
  end

  // REG#38の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0038 <= imem06_in[111:108];
    8: reg_0038 <= imem06_in[111:108];
    26: reg_0038 <= imem03_in[23:20];
    28: reg_0038 <= imem06_in[111:108];
    56: reg_0038 <= imem06_in[111:108];
    endcase
  end

  // REG#39の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0039 <= imem06_in[11:8];
    8: reg_0039 <= imem06_in[11:8];
    30: reg_0039 <= imem03_in[47:44];
    48: reg_0039 <= imem05_in[87:84];
    49: reg_0039 <= op1_12_out;
    50: reg_0039 <= op1_12_out;
    51: reg_0039 <= op1_12_out;
    52: reg_0039 <= op1_12_out;
    53: reg_0039 <= op1_12_out;
    54: reg_0039 <= op1_12_out;
    55: reg_0039 <= op1_12_out;
    57: reg_0039 <= op1_12_out;
    59: reg_0039 <= imem06_in[11:8];
    60: reg_0039 <= op1_12_out;
    62: reg_0039 <= imem02_in[79:76];
    64: reg_0039 <= imem05_in[87:84];
    66: reg_0039 <= op1_12_out;
    68: reg_0039 <= imem03_in[47:44];
    70: reg_0039 <= imem06_in[11:8];
    85: reg_0039 <= imem06_in[11:8];
    endcase
  end

  // REG#40の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0040 <= imem06_in[51:48];
    8: reg_0040 <= imem06_in[51:48];
    29: reg_0040 <= imem03_in[27:24];
    31: reg_0040 <= imem06_in[43:40];
    34: reg_0040 <= imem06_in[51:48];
    36: reg_0040 <= imem06_in[51:48];
    59: reg_0040 <= imem05_in[63:60];
    61: reg_0040 <= imem02_in[19:16];
    63: reg_0040 <= imem05_in[83:80];
    65: reg_0040 <= imem05_in[63:60];
    75: reg_0040 <= op2_03_out;
    endcase
  end

  // REG#41の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0041 <= imem04_in[31:28];
    9: reg_0041 <= imem01_in[107:104];
    37: reg_0041 <= imem06_in[67:64];
    38: reg_0041 <= op2_01_out;
    75: reg_0041 <= op2_01_out;
    endcase
  end

  // REG#42の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0042 <= imem02_in[15:12];
    11: reg_0042 <= imem05_in[39:36];
    13: reg_0042 <= op1_14_out;
    14: reg_0042 <= op2_00_out;
    36: reg_0042 <= op2_00_out;
    67: reg_0042 <= op2_00_out;
    83: reg_0042 <= imem02_in[15:12];
    93: reg_0042 <= op2_00_out;
    endcase
  end

  // REG#43の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0043 <= imem04_in[59:56];
    11: reg_0043 <= op1_13_out;
    12: reg_0043 <= op1_13_out;
    14: reg_0043 <= op1_13_out;
    16: reg_0043 <= imem04_in[59:56];
    17: reg_0043 <= op1_13_out;
    18: reg_0043 <= op1_13_out;
    20: reg_0043 <= op1_13_out;
    23: reg_0043 <= imem04_in[59:56];
    81: reg_0043 <= imem04_in[59:56];
    82: reg_0043 <= op1_13_out;
    84: reg_0043 <= imem02_in[11:8];
    endcase
  end

  // REG#44の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0044 <= imem04_in[111:108];
    11: reg_0044 <= op1_14_out;
    12: reg_0044 <= op2_00_out;
    29: reg_0044 <= op2_00_out;
    44: reg_0044 <= op2_00_out;
    52: reg_0044 <= op2_00_out;
    77: reg_0044 <= op1_14_out;
    79: reg_0044 <= op1_14_out;
    81: reg_0044 <= op1_14_out;
    83: reg_0044 <= op1_14_out;
    84: reg_0044 <= op2_00_out;
    95: reg_0044 <= op2_00_out;
    endcase
  end

  // REG#45の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0045 <= imem02_in[11:8];
    11: reg_0045 <= op2_00_out;
    26: reg_0045 <= op2_00_out;
    34: reg_0045 <= op2_00_out;
    62: reg_0045 <= imem02_in[11:8];
    71: reg_0045 <= imem02_in[11:8];
    81: reg_0045 <= op2_00_out;
    86: reg_0045 <= op2_00_out;
    endcase
  end

  // REG#46の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0046 <= imem04_in[11:8];
    12: reg_0046 <= op2_01_out;
    30: reg_0046 <= op2_01_out;
    49: reg_0046 <= op2_01_out;
    69: reg_0046 <= op2_01_out;
    90: reg_0046 <= op1_13_out;
    93: reg_0046 <= op2_01_out;
    endcase
  end

  // REG#47の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0047 <= imem04_in[19:16];
    13: reg_0047 <= op2_01_out;
    34: reg_0047 <= op2_01_out;
    62: reg_0047 <= op2_01_out;
    68: reg_0047 <= op2_01_out;
    86: reg_0047 <= op2_01_out;
    endcase
  end

  // REG#48の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0048 <= imem04_in[71:68];
    14: reg_0048 <= op2_02_out;
    38: reg_0048 <= op2_02_out;
    77: reg_0048 <= imem05_in[87:84];
    78: reg_0048 <= op2_02_out;
    endcase
  end

  // REG#49の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0049 <= imem02_in[75:72];
    14: reg_0049 <= op2_03_out;
    40: reg_0049 <= imem04_in[71:68];
    41: reg_0049 <= op2_02_out;
    44: reg_0049 <= op2_02_out;
    54: reg_0049 <= op2_02_out;
    85: reg_0049 <= op2_02_out;
    endcase
  end

  // REG#50の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0050 <= imem04_in[115:112];
    16: reg_0050 <= imem04_in[115:112];
    18: reg_0050 <= imem04_in[115:112];
    41: reg_0050 <= imem04_in[115:112];
    endcase
  end

  // REG#51の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0051 <= imem02_in[63:60];
    16: reg_0051 <= imem04_in[119:116];
    18: reg_0051 <= imem04_in[119:116];
    37: reg_0051 <= imem06_in[19:16];
    40: reg_0051 <= imem04_in[119:116];
    42: reg_0051 <= imem07_in[43:40];
    92: reg_0051 <= imem01_in[67:64];
    94: reg_0051 <= imem01_in[67:64];
    endcase
  end

  // REG#52の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0052 <= imem02_in[51:48];
    16: reg_0052 <= imem04_in[35:32];
    18: reg_0052 <= imem04_in[35:32];
    41: reg_0052 <= imem04_in[35:32];
    endcase
  end

  // REG#53の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0053 <= imem04_in[63:60];
    16: reg_0053 <= imem04_in[11:8];
    18: reg_0053 <= imem04_in[11:8];
    40: reg_0053 <= imem04_in[91:88];
    42: reg_0053 <= imem07_in[39:36];
    endcase
  end

  // REG#54の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0054 <= imem04_in[15:12];
    16: reg_0054 <= imem04_in[15:12];
    18: reg_0054 <= imem04_in[15:12];
    38: reg_0054 <= imem01_in[43:40];
    40: reg_0054 <= imem01_in[43:40];
    92: reg_0054 <= imem01_in[103:100];
    94: reg_0054 <= imem01_in[43:40];
    endcase
  end

  // REG#55の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0055 <= imem02_in[87:84];
    16: reg_0055 <= imem04_in[67:64];
    19: reg_0055 <= imem02_in[43:40];
    21: reg_0055 <= imem04_in[51:48];
    23: reg_0055 <= imem04_in[67:64];
    82: reg_0055 <= imem02_in[43:40];
    84: reg_0055 <= imem02_in[87:84];
    endcase
  end

  // REG#56の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0056 <= imem04_in[55:52];
    16: reg_0056 <= imem04_in[55:52];
    19: reg_0056 <= imem02_in[47:44];
    21: reg_0056 <= imem04_in[55:52];
    23: reg_0056 <= imem04_in[55:52];
    81: reg_0056 <= imem04_in[55:52];
    83: reg_0056 <= imem02_in[47:44];
    endcase
  end

  // REG#57の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0057 <= imem04_in[87:84];
    16: reg_0057 <= imem04_in[87:84];
    19: reg_0057 <= imem02_in[7:4];
    21: reg_0057 <= imem04_in[91:88];
    23: reg_0057 <= imem04_in[87:84];
    79: reg_0057 <= imem07_in[23:20];
    81: reg_0057 <= imem04_in[87:84];
    83: reg_0057 <= imem02_in[7:4];
    endcase
  end

  // REG#58の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0058 <= imem04_in[39:36];
    16: reg_0058 <= imem04_in[107:104];
    19: reg_0058 <= imem02_in[107:104];
    21: reg_0058 <= imem04_in[107:104];
    23: reg_0058 <= imem04_in[107:104];
    78: reg_0058 <= imem05_in[123:120];
    82: reg_0058 <= imem04_in[39:36];
    endcase
  end

  // REG#59の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0059 <= imem04_in[3:0];
    16: reg_0059 <= imem04_in[95:92];
    19: reg_0059 <= imem02_in[123:120];
    21: reg_0059 <= imem04_in[3:0];
    23: reg_0059 <= imem04_in[3:0];
    81: reg_0059 <= imem04_in[95:92];
    83: reg_0059 <= imem02_in[123:120];
    endcase
  end

  // REG#60の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0060 <= imem02_in[91:88];
    16: reg_0060 <= imem04_in[79:76];
    19: reg_0060 <= imem02_in[51:48];
    21: reg_0060 <= imem04_in[79:76];
    23: reg_0060 <= imem04_in[79:76];
    82: reg_0060 <= imem04_in[79:76];
    endcase
  end

  // REG#61の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0061 <= imem04_in[7:4];
    17: reg_0061 <= imem04_in[7:4];
    42: reg_0061 <= imem07_in[55:52];
    endcase
  end

  // REG#62の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0062 <= imem04_in[27:24];
    17: reg_0062 <= imem04_in[27:24];
    44: reg_0062 <= imem04_in[27:24];
    46: reg_0062 <= imem01_in[7:4];
    48: reg_0062 <= imem04_in[27:24];
    55: reg_0062 <= imem06_in[11:8];
    58: reg_0062 <= imem04_in[27:24];
    94: reg_0062 <= imem01_in[7:4];
    endcase
  end

  // REG#63の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0063 <= imem04_in[79:76];
    17: reg_0063 <= imem04_in[79:76];
    42: reg_0063 <= op1_13_out;
    44: reg_0063 <= imem04_in[35:32];
    45: reg_0063 <= op1_13_out;
    47: reg_0063 <= imem04_in[35:32];
    48: reg_0063 <= op1_13_out;
    50: reg_0063 <= op1_13_out;
    52: reg_0063 <= imem03_in[3:0];
    54: reg_0063 <= imem03_in[3:0];
    86: reg_0063 <= imem03_in[3:0];
    87: reg_0063 <= op1_13_out;
    90: reg_0063 <= imem00_in[103:100];
    endcase
  end

  // REG#64の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0064 <= imem04_in[103:100];
    17: reg_0064 <= imem04_in[103:100];
    42: reg_0064 <= imem07_in[11:8];
    endcase
  end

  // REG#65の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0065 <= imem04_in[35:32];
    17: reg_0065 <= imem04_in[35:32];
    43: reg_0065 <= imem02_in[127:124];
    45: reg_0065 <= imem04_in[35:32];
    48: reg_0065 <= imem04_in[35:32];
    58: reg_0065 <= imem04_in[35:32];
    endcase
  end

  // REG#66の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0066 <= imem04_in[43:40];
    17: reg_0066 <= imem04_in[43:40];
    45: reg_0066 <= imem04_in[27:24];
    47: reg_0066 <= imem04_in[59:56];
    49: reg_0066 <= imem05_in[95:92];
    63: reg_0066 <= imem05_in[119:116];
    65: reg_0066 <= imem05_in[95:92];
    77: reg_0066 <= imem05_in[119:116];
    79: reg_0066 <= imem07_in[55:52];
    81: reg_0066 <= imem07_in[55:52];
    endcase
  end

  // REG#67の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0067 <= imem04_in[51:48];
    17: reg_0067 <= imem04_in[51:48];
    42: reg_0067 <= imem07_in[35:32];
    endcase
  end

  // REG#68の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0068 <= imem04_in[67:64];
    17: reg_0068 <= imem04_in[67:64];
    44: reg_0068 <= imem04_in[55:52];
    46: reg_0068 <= imem01_in[31:28];
    48: reg_0068 <= imem04_in[67:64];
    55: reg_0068 <= imem06_in[103:100];
    58: reg_0068 <= imem04_in[55:52];
    94: reg_0068 <= imem01_in[31:28];
    endcase
  end

  // REG#69の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0069 <= imem04_in[83:80];
    17: reg_0069 <= imem04_in[83:80];
    44: reg_0069 <= imem04_in[51:48];
    46: reg_0069 <= imem01_in[39:36];
    48: reg_0069 <= imem04_in[83:80];
    55: reg_0069 <= imem06_in[79:76];
    58: reg_0069 <= imem04_in[51:48];
    endcase
  end

  // REG#70の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0070 <= imem04_in[95:92];
    17: reg_0070 <= imem04_in[95:92];
    45: reg_0070 <= imem04_in[95:92];
    47: reg_0070 <= imem04_in[95:92];
    49: reg_0070 <= imem05_in[51:48];
    63: reg_0070 <= imem05_in[51:48];
    66: reg_0070 <= imem05_in[51:48];
    68: reg_0070 <= imem03_in[11:8];
    70: reg_0070 <= imem02_in[31:28];
    72: reg_0070 <= imem05_in[51:48];
    90: reg_0070 <= imem00_in[115:112];
    endcase
  end

  // REG#71の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0071 <= imem04_in[75:72];
    17: reg_0071 <= imem04_in[75:72];
    41: reg_0071 <= imem04_in[75:72];
    endcase
  end

  // REG#72の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0072 <= imem04_in[107:104];
    17: reg_0072 <= imem04_in[107:104];
    36: reg_0072 <= op2_01_out;
    69: reg_0072 <= imem06_in[107:104];
    70: reg_0072 <= op2_01_out;
    94: reg_0072 <= op2_01_out;
    endcase
  end

  // REG#73の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0073 <= imem02_in[111:108];
    16: reg_0073 <= op1_14_out;
    18: reg_0073 <= op1_14_out;
    20: reg_0073 <= op1_14_out;
    23: reg_0073 <= imem01_in[23:20];
    25: reg_0073 <= imem02_in[111:108];
    49: reg_0073 <= op1_14_out;
    52: reg_0073 <= imem01_in[23:20];
    endcase
  end

  // REG#74の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0074 <= imem04_in[99:96];
    17: reg_0074 <= imem04_in[99:96];
    41: reg_0074 <= imem04_in[99:96];
    endcase
  end

  // REG#75の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0075 <= imem04_in[91:88];
    17: reg_0075 <= imem04_in[91:88];
    44: reg_0075 <= imem04_in[47:44];
    46: reg_0075 <= imem01_in[71:68];
    48: reg_0075 <= imem04_in[47:44];
    57: reg_0075 <= imem04_in[91:88];
    59: reg_0075 <= imem06_in[7:4];
    61: reg_0075 <= imem02_in[79:76];
    63: reg_0075 <= imem05_in[15:12];
    65: reg_0075 <= imem05_in[15:12];
    78: reg_0075 <= imem05_in[15:12];
    81: reg_0075 <= imem04_in[91:88];
    83: reg_0075 <= imem02_in[79:76];
    endcase
  end

  // REG#76の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0076 <= imem04_in[47:44];
    17: reg_0076 <= imem04_in[47:44];
    41: reg_0076 <= imem04_in[47:44];
    endcase
  end

  // REG#77の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0077 <= imem02_in[99:96];
    17: reg_0077 <= imem04_in[71:68];
    41: reg_0077 <= imem04_in[71:68];
    90: reg_0077 <= imem00_in[43:40];
    endcase
  end

  // REG#78の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0078 <= imem04_in[23:20];
    17: reg_0078 <= imem04_in[23:20];
    45: reg_0078 <= imem04_in[23:20];
    48: reg_0078 <= imem04_in[23:20];
    58: reg_0078 <= imem04_in[23:20];
    endcase
  end

  // REG#79の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0079 <= imem02_in[115:112];
    17: reg_0079 <= imem04_in[19:16];
    41: reg_0079 <= imem04_in[19:16];
    endcase
  end

  // REG#80の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0080 <= imem02_in[31:28];
    18: reg_0080 <= imem05_in[47:44];
    20: reg_0080 <= imem02_in[31:28];
    81: reg_0080 <= imem04_in[35:32];
    83: reg_0080 <= imem02_in[31:28];
    endcase
  end

  // REG#81の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0081 <= imem02_in[27:24];
    18: reg_0081 <= imem05_in[99:96];
    20: reg_0081 <= imem02_in[27:24];
    83: reg_0081 <= imem02_in[27:24];
    endcase
  end

  // REG#82の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0082 <= imem02_in[67:64];
    18: reg_0082 <= imem05_in[111:108];
    20: reg_0082 <= imem02_in[67:64];
    74: reg_0082 <= op2_02_out;
    endcase
  end

  // REG#83の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0083 <= imem02_in[3:0];
    19: reg_0083 <= imem02_in[83:80];
    21: reg_0083 <= imem04_in[71:68];
    23: reg_0083 <= imem04_in[71:68];
    81: reg_0083 <= imem04_in[71:68];
    83: reg_0083 <= imem02_in[83:80];
    endcase
  end

  // REG#84の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0084 <= imem02_in[79:76];
    19: reg_0084 <= imem05_in[95:92];
    40: reg_0084 <= imem04_in[115:112];
    42: reg_0084 <= imem07_in[103:100];
    endcase
  end

  // REG#85の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0085 <= imem02_in[39:36];
    19: reg_0085 <= imem05_in[59:56];
    46: reg_0085 <= imem01_in[11:8];
    48: reg_0085 <= imem01_in[11:8];
    64: reg_0085 <= imem05_in[67:64];
    66: reg_0085 <= imem05_in[59:56];
    68: reg_0085 <= imem01_in[11:8];
    92: reg_0085 <= imem01_in[11:8];
    endcase
  end

  // REG#86の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0086 <= imem02_in[55:52];
    19: reg_0086 <= imem05_in[123:120];
    46: reg_0086 <= imem01_in[51:48];
    49: reg_0086 <= imem05_in[123:120];
    65: reg_0086 <= imem05_in[123:120];
    77: reg_0086 <= imem05_in[55:52];
    79: reg_0086 <= imem07_in[119:116];
    81: reg_0086 <= imem04_in[79:76];
    83: reg_0086 <= imem02_in[55:52];
    endcase
  end

  // REG#87の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0087 <= imem02_in[95:92];
    19: reg_0087 <= imem02_in[95:92];
    21: reg_0087 <= imem04_in[43:40];
    23: reg_0087 <= imem04_in[43:40];
    81: reg_0087 <= imem04_in[75:72];
    83: reg_0087 <= imem02_in[95:92];
    endcase
  end

  // REG#88の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0088 <= imem02_in[19:16];
    19: reg_0088 <= imem02_in[19:16];
    21: reg_0088 <= imem04_in[63:60];
    23: reg_0088 <= imem04_in[63:60];
    80: reg_0088 <= op1_13_out;
    83: reg_0088 <= imem02_in[19:16];
    endcase
  end

  // REG#89の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0089 <= imem02_in[23:20];
    19: reg_0089 <= imem05_in[127:124];
    46: reg_0089 <= imem01_in[23:20];
    49: reg_0089 <= imem05_in[127:124];
    62: reg_0089 <= imem02_in[23:20];
    71: reg_0089 <= imem05_in[127:124];
    73: reg_0089 <= imem07_in[15:12];
    77: reg_0089 <= imem07_in[15:12];
    79: reg_0089 <= imem07_in[15:12];
    81: reg_0089 <= imem07_in[15:12];
    endcase
  end

  // REG#90の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0090 <= imem02_in[59:56];
    19: reg_0090 <= imem05_in[7:4];
    47: reg_0090 <= imem04_in[51:48];
    49: reg_0090 <= imem05_in[7:4];
    63: reg_0090 <= imem05_in[7:4];
    66: reg_0090 <= imem05_in[83:80];
    68: reg_0090 <= imem03_in[71:68];
    70: reg_0090 <= imem02_in[59:56];
    72: reg_0090 <= imem05_in[83:80];
    endcase
  end

  // REG#91の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0091 <= imem02_in[71:68];
    19: reg_0091 <= imem05_in[3:0];
    47: reg_0091 <= imem04_in[127:124];
    49: reg_0091 <= imem05_in[3:0];
    61: reg_0091 <= imem02_in[23:20];
    62: reg_0091 <= op1_15_out;
    64: reg_0091 <= op1_15_out;
    67: reg_0091 <= imem05_in[3:0];
    68: reg_0091 <= op1_15_out;
    71: reg_0091 <= imem05_in[3:0];
    73: reg_0091 <= op1_15_out;
    77: reg_0091 <= imem05_in[3:0];
    79: reg_0091 <= imem07_in[95:92];
    81: reg_0091 <= imem07_in[95:92];
    endcase
  end

  // REG#92の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0092 <= imem02_in[7:4];
    20: reg_0092 <= imem02_in[7:4];
    84: reg_0092 <= imem02_in[7:4];
    endcase
  end

  // REG#93の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0093 <= imem02_in[107:104];
    20: reg_0093 <= imem02_in[107:104];
    84: reg_0093 <= imem02_in[107:104];
    endcase
  end

  // REG#94の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0094 <= imem02_in[103:100];
    20: reg_0094 <= imem02_in[103:100];
    84: reg_0094 <= imem02_in[103:100];
    endcase
  end

  // REG#95の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0095 <= imem02_in[35:32];
    20: reg_0095 <= imem02_in[35:32];
    84: reg_0095 <= imem02_in[35:32];
    endcase
  end

  // REG#96の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0096 <= imem02_in[43:40];
    20: reg_0096 <= imem02_in[43:40];
    84: reg_0096 <= imem02_in[43:40];
    endcase
  end

  // REG#97の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0097 <= imem02_in[47:44];
    20: reg_0097 <= imem02_in[47:44];
    84: reg_0097 <= imem02_in[47:44];
    endcase
  end

  // REG#98の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0098 <= imem02_in[83:80];
    20: reg_0098 <= imem02_in[83:80];
    84: reg_0098 <= imem02_in[83:80];
    91: reg_0098 <= imem01_in[27:24];
    94: reg_0098 <= imem01_in[27:24];
    endcase
  end

  // REG#99の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0099 <= imem01_in[43:40];
    46: reg_0099 <= imem01_in[55:52];
    49: reg_0099 <= imem05_in[23:20];
    63: reg_0099 <= imem05_in[23:20];
    65: reg_0099 <= imem05_in[23:20];
    77: reg_0099 <= imem05_in[23:20];
    79: reg_0099 <= imem07_in[123:120];
    81: reg_0099 <= imem07_in[59:56];
    endcase
  end

  // REG#100の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0100 <= imem01_in[71:68];
    48: reg_0100 <= imem01_in[71:68];
    67: reg_0100 <= imem01_in[71:68];
    69: reg_0100 <= imem06_in[103:100];
    71: reg_0100 <= imem05_in[119:116];
    73: reg_0100 <= imem07_in[75:72];
    77: reg_0100 <= imem07_in[75:72];
    79: reg_0100 <= imem07_in[75:72];
    81: reg_0100 <= imem07_in[75:72];
    endcase
  end

  // REG#101の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0101 <= imem01_in[79:76];
    49: reg_0101 <= imem05_in[115:112];
    64: reg_0101 <= imem05_in[95:92];
    66: reg_0101 <= imem05_in[115:112];
    68: reg_0101 <= imem01_in[79:76];
    92: reg_0101 <= imem01_in[79:76];
    94: reg_0101 <= imem01_in[79:76];
    endcase
  end

  // REG#102の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0102 <= imem01_in[63:60];
    49: reg_0102 <= imem05_in[55:52];
    64: reg_0102 <= imem05_in[55:52];
    66: reg_0102 <= imem05_in[55:52];
    68: reg_0102 <= imem01_in[63:60];
    endcase
  end

  // REG#103の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0103 <= imem01_in[19:16];
    49: reg_0103 <= imem05_in[47:44];
    65: reg_0103 <= imem05_in[47:44];
    74: reg_0103 <= imem07_in[123:120];
    78: reg_0103 <= imem07_in[123:120];
    91: reg_0103 <= op2_00_out;
    endcase
  end

  // REG#104の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0104 <= imem01_in[39:36];
    50: reg_0104 <= imem02_in[99:96];
    52: reg_0104 <= imem01_in[39:36];
    95: reg_0104 <= imem01_in[39:36];
    endcase
  end

  // REG#105の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0105 <= imem01_in[7:4];
    50: reg_0105 <= imem02_in[63:60];
    52: reg_0105 <= imem01_in[7:4];
    endcase
  end

  // REG#106の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0106 <= imem01_in[75:72];
    50: reg_0106 <= imem02_in[15:12];
    52: reg_0106 <= imem01_in[75:72];
    endcase
  end

  // REG#107の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0107 <= imem01_in[91:88];
    50: reg_0107 <= imem02_in[35:32];
    52: reg_0107 <= imem01_in[91:88];
    91: reg_0107 <= imem01_in[91:88];
    endcase
  end

  // REG#108の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0108 <= imem01_in[59:56];
    50: reg_0108 <= imem02_in[59:56];
    52: reg_0108 <= imem01_in[59:56];
    endcase
  end

  // REG#109の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0109 <= imem01_in[87:84];
    51: reg_0109 <= imem01_in[87:84];
    53: reg_0109 <= imem00_in[83:80];
    55: reg_0109 <= imem06_in[43:40];
    58: reg_0109 <= imem04_in[115:112];
    84: reg_0109 <= imem02_in[27:24];
    endcase
  end

  // REG#110の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0110 <= imem01_in[115:112];
    51: reg_0110 <= imem01_in[7:4];
    53: reg_0110 <= imem00_in[99:96];
    55: reg_0110 <= imem05_in[39:36];
    59: reg_0110 <= imem06_in[71:68];
    61: reg_0110 <= imem02_in[39:36];
    63: reg_0110 <= imem05_in[11:8];
    66: reg_0110 <= imem05_in[11:8];
    68: reg_0110 <= imem01_in[115:112];
    81: reg_0110 <= imem07_in[31:28];
    endcase
  end

  // REG#111の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0111 <= imem01_in[23:20];
    51: reg_0111 <= imem01_in[23:20];
    53: reg_0111 <= imem00_in[119:116];
    55: reg_0111 <= imem05_in[59:56];
    59: reg_0111 <= imem06_in[99:96];
    61: reg_0111 <= imem02_in[83:80];
    63: reg_0111 <= imem05_in[59:56];
    66: reg_0111 <= imem05_in[23:20];
    68: reg_0111 <= imem01_in[23:20];
    92: reg_0111 <= imem01_in[23:20];
    94: reg_0111 <= imem01_in[23:20];
    endcase
  end

  // REG#112の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0112 <= imem01_in[55:52];
    51: reg_0112 <= imem01_in[111:108];
    53: reg_0112 <= imem00_in[27:24];
    55: reg_0112 <= imem05_in[55:52];
    59: reg_0112 <= imem06_in[111:108];
    61: reg_0112 <= imem02_in[87:84];
    63: reg_0112 <= imem05_in[107:104];
    66: reg_0112 <= imem05_in[107:104];
    68: reg_0112 <= imem01_in[55:52];
    90: reg_0112 <= imem00_in[27:24];
    endcase
  end

  // REG#113の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0113 <= imem01_in[103:100];
    51: reg_0113 <= imem01_in[103:100];
    53: reg_0113 <= imem00_in[3:0];
    55: reg_0113 <= imem05_in[75:72];
    60: reg_0113 <= imem05_in[75:72];
    63: reg_0113 <= op1_13_out;
    65: reg_0113 <= op1_13_out;
    67: reg_0113 <= op1_13_out;
    68: reg_0113 <= op1_13_out;
    69: reg_0113 <= op1_13_out;
    72: reg_0113 <= imem05_in[75:72];
    endcase
  end

  // REG#114の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0114 <= imem01_in[67:64];
    51: reg_0114 <= imem01_in[15:12];
    53: reg_0114 <= imem00_in[51:48];
    55: reg_0114 <= imem05_in[119:116];
    60: reg_0114 <= imem05_in[39:36];
    62: reg_0114 <= imem02_in[107:104];
    68: reg_0114 <= imem01_in[67:64];
    91: reg_0114 <= imem01_in[67:64];
    endcase
  end

  // REG#115の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0115 <= imem01_in[83:80];
    51: reg_0115 <= imem01_in[83:80];
    54: reg_0115 <= imem05_in[43:40];
    56: reg_0115 <= imem06_in[23:20];
    89: reg_0115 <= imem00_in[111:108];
    91: reg_0115 <= imem01_in[87:84];
    95: reg_0115 <= imem01_in[87:84];
    endcase
  end

  // REG#116の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0116 <= imem01_in[35:32];
    51: reg_0116 <= imem01_in[79:76];
    54: reg_0116 <= imem03_in[75:72];
    81: reg_0116 <= imem07_in[19:16];
    endcase
  end

  // REG#117の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0117 <= imem01_in[99:96];
    51: reg_0117 <= imem01_in[119:116];
    54: reg_0117 <= imem00_in[91:88];
    82: reg_0117 <= imem02_in[67:64];
    84: reg_0117 <= imem02_in[67:64];
    endcase
  end

  // REG#118の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0118 <= imem01_in[27:24];
    52: reg_0118 <= imem01_in[27:24];
    endcase
  end

  // REG#119の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0119 <= imem01_in[47:44];
    52: reg_0119 <= imem01_in[47:44];
    95: reg_0119 <= imem01_in[47:44];
    endcase
  end

  // REG#120の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0120 <= imem01_in[51:48];
    52: reg_0120 <= imem01_in[51:48];
    endcase
  end

  // REG#121の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0121 <= imem01_in[107:104];
    52: reg_0121 <= imem01_in[107:104];
    endcase
  end

  // REG#122の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0122 <= imem01_in[11:8];
    52: reg_0122 <= imem01_in[11:8];
    endcase
  end

  // REG#123の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0123 <= imem01_in[3:0];
    52: reg_0123 <= imem01_in[3:0];
    endcase
  end

  // REG#124の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0124 <= imem01_in[15:12];
    52: reg_0124 <= imem01_in[15:12];
    94: reg_0124 <= imem01_in[15:12];
    endcase
  end

  // REG#125の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0125 <= imem01_in[31:28];
    52: reg_0125 <= imem01_in[31:28];
    endcase
  end

  // REG#126の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0126 <= imem01_in[111:108];
    52: reg_0126 <= imem01_in[111:108];
    endcase
  end

  // REG#127の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0127 <= imem01_in[95:92];
    52: reg_0127 <= imem01_in[95:92];
    endcase
  end

  // REG#128の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0128 <= imem05_in[43:40];
    65: reg_0128 <= imem05_in[43:40];
    70: reg_0128 <= imem02_in[95:92];
    72: reg_0128 <= imem05_in[43:40];
    endcase
  end

  // REG#129の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0129 <= imem05_in[79:76];
    67: reg_0129 <= op2_01_out;
    83: reg_0129 <= op2_01_out;
    95: reg_0129 <= op2_01_out;
    endcase
  end

  // REG#130の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0130 <= imem05_in[91:88];
    68: reg_0130 <= imem01_in[99:96];
    88: reg_0130 <= imem03_in[103:100];
    90: reg_0130 <= imem00_in[91:88];
    endcase
  end

  // REG#131の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0131 <= imem05_in[107:104];
    68: reg_0131 <= imem01_in[71:68];
    90: reg_0131 <= imem00_in[95:92];
    endcase
  end

  // REG#132の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0132 <= imem05_in[3:0];
    69: reg_0132 <= imem06_in[119:116];
    71: reg_0132 <= imem05_in[91:88];
    74: reg_0132 <= imem07_in[67:64];
    77: reg_0132 <= imem05_in[91:88];
    79: reg_0132 <= imem07_in[115:112];
    82: reg_0132 <= imem02_in[31:28];
    84: reg_0132 <= imem02_in[31:28];
    endcase
  end

  // REG#133の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0133 <= imem05_in[31:28];
    70: reg_0133 <= imem02_in[27:24];
    72: reg_0133 <= imem05_in[31:28];
    endcase
  end

  // REG#134の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0134 <= imem05_in[111:108];
    70: reg_0134 <= imem02_in[63:60];
    72: reg_0134 <= imem05_in[111:108];
    endcase
  end

  // REG#135の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0135 <= imem05_in[23:20];
    70: reg_0135 <= imem02_in[115:112];
    72: reg_0135 <= imem05_in[23:20];
    endcase
  end

  // REG#136の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0136 <= imem05_in[27:24];
    71: reg_0136 <= imem05_in[19:16];
    73: reg_0136 <= op1_12_out;
    77: reg_0136 <= imem05_in[19:16];
    78: reg_0136 <= op1_12_out;
    79: reg_0136 <= op1_12_out;
    81: reg_0136 <= op1_12_out;
    84: reg_0136 <= imem02_in[59:56];
    endcase
  end

  // REG#137の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0137 <= imem05_in[103:100];
    71: reg_0137 <= imem05_in[103:100];
    73: reg_0137 <= imem05_in[103:100];
    endcase
  end

  // REG#138の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0138 <= imem05_in[75:72];
    71: reg_0138 <= imem02_in[123:120];
    78: reg_0138 <= imem05_in[75:72];
    86: reg_0138 <= imem05_in[75:72];
    endcase
  end

  // REG#139の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0139 <= imem05_in[71:68];
    71: reg_0139 <= imem02_in[55:52];
    78: reg_0139 <= imem05_in[71:68];
    81: reg_0139 <= imem07_in[3:0];
    endcase
  end

  // REG#140の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0140 <= imem05_in[95:92];
    71: reg_0140 <= imem02_in[87:84];
    81: reg_0140 <= imem07_in[111:108];
    endcase
  end

  // REG#141の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0141 <= imem05_in[87:84];
    71: reg_0141 <= imem02_in[43:40];
    81: reg_0141 <= imem07_in[71:68];
    endcase
  end

  // REG#142の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0142 <= imem05_in[51:48];
    71: reg_0142 <= imem02_in[19:16];
    81: reg_0142 <= imem07_in[39:36];
    endcase
  end

  // REG#143の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0143 <= imem05_in[67:64];
    71: reg_0143 <= imem05_in[67:64];
    73: reg_0143 <= imem05_in[67:64];
    endcase
  end

  // REG#144の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0144 <= imem05_in[115:112];
    72: reg_0144 <= imem05_in[115:112];
    endcase
  end

  // REG#145の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0145 <= imem05_in[19:16];
    72: reg_0145 <= imem05_in[19:16];
    88: reg_0145 <= imem03_in[67:64];
    90: reg_0145 <= imem00_in[87:84];
    endcase
  end

  // REG#146の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0146 <= imem05_in[55:52];
    72: reg_0146 <= imem05_in[55:52];
    endcase
  end

  // REG#147の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0147 <= imem05_in[7:4];
    73: reg_0147 <= imem05_in[7:4];
    endcase
  end

  // REG#148の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0148 <= imem05_in[11:8];
    73: reg_0148 <= imem05_in[11:8];
    endcase
  end

  // REG#149の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0149 <= imem05_in[15:12];
    73: reg_0149 <= imem05_in[15:12];
    endcase
  end

  // REG#150の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0150 <= imem05_in[35:32];
    73: reg_0150 <= imem05_in[35:32];
    endcase
  end

  // REG#151の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0151 <= imem05_in[39:36];
    73: reg_0151 <= imem05_in[39:36];
    endcase
  end

  // REG#152の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0152 <= imem05_in[47:44];
    73: reg_0152 <= imem05_in[47:44];
    91: reg_0152 <= imem01_in[75:72];
    endcase
  end

  // REG#153の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0153 <= imem05_in[83:80];
    73: reg_0153 <= imem05_in[83:80];
    endcase
  end

  // REG#154の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0154 <= imem05_in[63:60];
    73: reg_0154 <= imem05_in[63:60];
    endcase
  end

  // REG#155の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0155 <= imem05_in[99:96];
    73: reg_0155 <= imem05_in[99:96];
    endcase
  end

  // REG#156の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0156 <= imem05_in[59:56];
    73: reg_0156 <= imem05_in[59:56];
    endcase
  end

  // REG#157の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0157 <= imem07_in[95:92];
    74: reg_0157 <= imem07_in[111:108];
    78: reg_0157 <= imem07_in[111:108];
    endcase
  end

  // REG#158の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0158 <= imem07_in[103:100];
    74: reg_0158 <= imem07_in[103:100];
    78: reg_0158 <= imem07_in[103:100];
    endcase
  end

  // REG#159の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0159 <= imem07_in[43:40];
    78: reg_0159 <= imem07_in[43:40];
    endcase
  end

  // REG#160の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0160 <= imem07_in[55:52];
    78: reg_0160 <= imem07_in[55:52];
    endcase
  end

  // REG#161の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0161 <= imem07_in[31:28];
    78: reg_0161 <= imem07_in[31:28];
    endcase
  end

  // REG#162の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0162 <= imem07_in[35:32];
    78: reg_0162 <= imem07_in[35:32];
    endcase
  end

  // REG#163の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0163 <= imem07_in[59:56];
    78: reg_0163 <= imem07_in[59:56];
    86: reg_0163 <= imem03_in[123:120];
    88: reg_0163 <= imem06_in[7:4];
    90: reg_0163 <= imem00_in[35:32];
    endcase
  end

  // REG#164の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0164 <= imem07_in[75:72];
    78: reg_0164 <= imem07_in[75:72];
    endcase
  end

  // REG#165の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0165 <= imem07_in[19:16];
    77: reg_0165 <= imem07_in[19:16];
    79: reg_0165 <= imem07_in[35:32];
    82: reg_0165 <= imem02_in[63:60];
    85: reg_0165 <= imem05_in[63:60];
    87: reg_0165 <= imem06_in[39:36];
    89: reg_0165 <= imem00_in[79:76];
    91: reg_0165 <= imem01_in[71:68];
    endcase
  end

  // REG#166の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0166 <= imem07_in[67:64];
    78: reg_0166 <= imem07_in[67:64];
    endcase
  end

  // REG#167の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0167 <= imem07_in[39:36];
    78: reg_0167 <= imem07_in[39:36];
    endcase
  end

  // REG#168の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0168 <= imem07_in[83:80];
    79: reg_0168 <= imem07_in[127:124];
    82: reg_0168 <= imem02_in[119:116];
    85: reg_0168 <= imem06_in[23:20];
    endcase
  end

  // REG#169の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0169 <= imem07_in[47:44];
    79: reg_0169 <= imem07_in[43:40];
    82: reg_0169 <= imem02_in[27:24];
    85: reg_0169 <= imem06_in[111:108];
    endcase
  end

  // REG#170の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0170 <= imem07_in[91:88];
    79: reg_0170 <= imem07_in[91:88];
    81: reg_0170 <= imem07_in[91:88];
    endcase
  end

  // REG#171の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0171 <= imem07_in[111:108];
    79: reg_0171 <= imem07_in[111:108];
    82: reg_0171 <= imem04_in[23:20];
    90: reg_0171 <= imem00_in[111:108];
    endcase
  end

  // REG#172の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0172 <= imem07_in[15:12];
    78: reg_0172 <= op2_00_out;
    endcase
  end

  // REG#173の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0173 <= imem07_in[107:104];
    79: reg_0173 <= imem07_in[107:104];
    82: reg_0173 <= imem04_in[27:24];
    endcase
  end

  // REG#174の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0174 <= imem07_in[3:0];
    79: reg_0174 <= imem07_in[3:0];
    82: reg_0174 <= imem04_in[127:124];
    endcase
  end

  // REG#175の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0175 <= imem07_in[7:4];
    79: reg_0175 <= imem07_in[7:4];
    81: reg_0175 <= imem07_in[7:4];
    endcase
  end

  // REG#176の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0176 <= imem07_in[99:96];
    79: reg_0176 <= imem07_in[99:96];
    81: reg_0176 <= imem07_in[99:96];
    endcase
  end

  // REG#177の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0177 <= imem07_in[71:68];
    79: reg_0177 <= imem07_in[71:68];
    82: reg_0177 <= imem04_in[43:40];
    endcase
  end

  // REG#178の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0178 <= imem07_in[87:84];
    81: reg_0178 <= imem07_in[87:84];
    endcase
  end

  // REG#179の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0179 <= imem07_in[27:24];
    79: reg_0179 <= imem07_in[27:24];
    82: reg_0179 <= imem04_in[55:52];
    endcase
  end

  // REG#180の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0180 <= imem07_in[11:8];
    81: reg_0180 <= imem07_in[11:8];
    endcase
  end

  // REG#181の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0181 <= imem07_in[23:20];
    81: reg_0181 <= imem07_in[23:20];
    endcase
  end

  // REG#182の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0182 <= imem07_in[51:48];
    81: reg_0182 <= imem07_in[51:48];
    endcase
  end

  // REG#183の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0183 <= imem07_in[63:60];
    81: reg_0183 <= imem07_in[63:60];
    endcase
  end

  // REG#184の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0184 <= imem07_in[115:112];
    81: reg_0184 <= imem07_in[115:112];
    endcase
  end

  // REG#185の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0185 <= imem07_in[79:76];
    81: reg_0185 <= imem07_in[79:76];
    endcase
  end

  // REG#186の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0186 <= imem00_in[59:56];
    87: reg_0186 <= imem03_in[3:0];
    89: reg_0186 <= imem03_in[3:0];
    endcase
  end

  // REG#187の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0187 <= imem00_in[27:24];
    88: reg_0187 <= imem03_in[35:32];
    89: reg_0187 <= op2_01_out;
    endcase
  end

  // REG#188の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0188 <= imem00_in[39:36];
    89: reg_0188 <= imem03_in[103:100];
    91: reg_0188 <= imem01_in[111:108];
    endcase
  end

  // REG#189の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0189 <= imem00_in[23:20];
    90: reg_0189 <= imem00_in[23:20];
    endcase
  end

  // REG#190の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0190 <= imem00_in[91:88];
    endcase
  end

  // REG#191の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0191 <= imem00_in[15:12];
    endcase
  end

  // REG#192の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0192 <= imem00_in[111:108];
    endcase
  end

  // REG#193の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0193 <= imem00_in[47:44];
    endcase
  end

  // REG#194の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0194 <= imem00_in[63:60];
    endcase
  end

  // REG#195の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0195 <= imem00_in[99:96];
    endcase
  end

  // REG#196の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0196 <= imem00_in[79:76];
    endcase
  end

  // REG#197の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0197 <= imem00_in[115:112];
    endcase
  end

  // REG#198の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0198 <= imem00_in[67:64];
    endcase
  end

  // REG#199の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0199 <= imem00_in[107:104];
    endcase
  end

  // REG#200の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0200 <= imem00_in[7:4];
    endcase
  end

  // REG#201の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0201 <= imem00_in[71:68];
    endcase
  end

  // REG#202の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0202 <= imem00_in[95:92];
    endcase
  end

  // REG#203の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0203 <= imem00_in[43:40];
    endcase
  end

  // REG#204の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0204 <= imem00_in[35:32];
    endcase
  end

  // REG#205の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0205 <= imem00_in[87:84];
    endcase
  end

  // REG#206の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0206 <= imem00_in[103:100];
    endcase
  end

  // REG#207の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0207 <= imem00_in[51:48];
    endcase
  end

  // REG#208の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0208 <= imem00_in[11:8];
    endcase
  end

  // REG#209の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0209 <= imem00_in[31:28];
    endcase
  end

  // REG#210の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0210 <= imem00_in[19:16];
    endcase
  end

  // REG#211の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0211 <= imem00_in[55:52];
    endcase
  end

  // REG#212の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0212 <= imem00_in[83:80];
    endcase
  end

  // REG#213の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0213 <= imem00_in[75:72];
    endcase
  end

  // REG#214の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0214 <= imem00_in[3:0];
    endcase
  end

  // REG#215の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0215 <= imem05_in[11:8];
    7: reg_0215 <= imem06_in[95:92];
    9: reg_0215 <= imem01_in[23:20];
    38: reg_0215 <= imem06_in[95:92];
    49: reg_0215 <= imem05_in[11:8];
    65: reg_0215 <= imem05_in[11:8];
    78: reg_0215 <= imem05_in[11:8];
    85: reg_0215 <= imem06_in[95:92];
    endcase
  end

  // REG#216の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0216 <= imem01_in[67:64];
    7: reg_0216 <= imem06_in[35:32];
    9: reg_0216 <= imem01_in[67:64];
    40: reg_0216 <= imem01_in[67:64];
    89: reg_0216 <= imem03_in[107:104];
    endcase
  end

  // REG#217の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0217 <= imem05_in[15:12];
    7: reg_0217 <= imem06_in[3:0];
    9: reg_0217 <= imem01_in[47:44];
    38: reg_0217 <= imem01_in[47:44];
    40: reg_0217 <= imem01_in[47:44];
    91: reg_0217 <= imem01_in[47:44];
    93: reg_0217 <= imem01_in[47:44];
    endcase
  end

  // REG#218の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0218 <= imem01_in[35:32];
    7: reg_0218 <= imem06_in[47:44];
    9: reg_0218 <= imem01_in[35:32];
    38: reg_0218 <= imem06_in[47:44];
    55: reg_0218 <= imem05_in[115:112];
    60: reg_0218 <= imem06_in[47:44];
    70: reg_0218 <= imem06_in[47:44];
    88: reg_0218 <= imem06_in[47:44];
    endcase
  end

  // REG#219の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0219 <= imem01_in[119:116];
    7: reg_0219 <= imem06_in[55:52];
    9: reg_0219 <= imem01_in[119:116];
    37: reg_0219 <= imem06_in[55:52];
    40: reg_0219 <= imem01_in[119:116];
    94: reg_0219 <= imem01_in[119:116];
    endcase
  end

  // REG#220の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0220 <= imem01_in[71:68];
    7: reg_0220 <= imem06_in[127:124];
    9: reg_0220 <= imem01_in[71:68];
    40: reg_0220 <= imem01_in[71:68];
    92: reg_0220 <= imem01_in[71:68];
    endcase
  end

  // REG#221の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0221 <= imem01_in[115:112];
    6: reg_0221 <= op2_01_out;
    10: reg_0221 <= op2_01_out;
    24: reg_0221 <= op2_01_out;
    28: reg_0221 <= op2_01_out;
    42: reg_0221 <= op2_01_out;
    46: reg_0221 <= op2_01_out;
    59: reg_0221 <= op2_01_out;
    endcase
  end

  // REG#222の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0222 <= imem01_in[23:20];
    6: reg_0222 <= op2_02_out;
    11: reg_0222 <= op2_02_out;
    28: reg_0222 <= op2_02_out;
    43: reg_0222 <= op2_02_out;
    50: reg_0222 <= op2_02_out;
    73: reg_0222 <= op2_02_out;
    endcase
  end

  // REG#223の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0223 <= imem05_in[127:124];
    6: reg_0223 <= op2_03_out;
    12: reg_0223 <= op2_03_out;
    32: reg_0223 <= op2_03_out;
    58: reg_0223 <= imem04_in[15:12];
    88: reg_0223 <= imem03_in[87:84];
    89: reg_0223 <= op2_03_out;
    endcase
  end

  // REG#224の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0224 <= imem01_in[59:56];
    8: reg_0224 <= imem01_in[59:56];
    11: reg_0224 <= imem05_in[75:72];
    16: reg_0224 <= imem04_in[91:88];
    19: reg_0224 <= imem05_in[75:72];
    47: reg_0224 <= imem04_in[91:88];
    49: reg_0224 <= imem05_in[75:72];
    61: reg_0224 <= imem02_in[119:116];
    63: reg_0224 <= imem05_in[75:72];
    66: reg_0224 <= imem05_in[75:72];
    68: reg_0224 <= imem01_in[59:56];
    88: reg_0224 <= imem06_in[111:108];
    endcase
  end

  // REG#225の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0225 <= imem01_in[127:124];
    8: reg_0225 <= imem01_in[127:124];
    10: reg_0225 <= imem01_in[127:124];
    19: reg_0225 <= imem05_in[11:8];
    48: reg_0225 <= imem01_in[127:124];
    64: reg_0225 <= imem05_in[11:8];
    66: reg_0225 <= imem05_in[71:68];
    68: reg_0225 <= imem01_in[127:124];
    91: reg_0225 <= imem01_in[127:124];
    93: reg_0225 <= imem01_in[127:124];
    endcase
  end

  // REG#226の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0226 <= imem01_in[11:8];
    8: reg_0226 <= imem01_in[11:8];
    11: reg_0226 <= imem05_in[63:60];
    16: reg_0226 <= imem04_in[75:72];
    19: reg_0226 <= imem05_in[63:60];
    49: reg_0226 <= imem05_in[63:60];
    63: reg_0226 <= imem05_in[123:120];
    67: reg_0226 <= imem05_in[63:60];
    72: reg_0226 <= imem05_in[123:120];
    endcase
  end

  // REG#227の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0227 <= imem01_in[63:60];
    8: reg_0227 <= imem01_in[63:60];
    10: reg_0227 <= imem01_in[63:60];
    24: reg_0227 <= imem01_in[63:60];
    44: reg_0227 <= imem04_in[75:72];
    46: reg_0227 <= imem01_in[63:60];
    48: reg_0227 <= imem04_in[75:72];
    57: reg_0227 <= imem04_in[43:40];
    59: reg_0227 <= imem06_in[95:92];
    61: reg_0227 <= imem02_in[27:24];
    64: reg_0227 <= imem05_in[83:80];
    67: reg_0227 <= imem05_in[83:80];
    72: reg_0227 <= imem05_in[35:32];
    endcase
  end

  // REG#228の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0228 <= imem01_in[107:104];
    8: reg_0228 <= imem01_in[107:104];
    11: reg_0228 <= imem05_in[127:124];
    15: reg_0228 <= op2_00_out;
    40: reg_0228 <= op2_00_out;
    81: reg_0228 <= imem07_in[67:64];
    96: reg_0228 <= op2_00_out;
    endcase
  end

  // REG#229の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0229 <= imem05_in[63:60];
    8: reg_0229 <= imem01_in[43:40];
    10: reg_0229 <= imem01_in[43:40];
    23: reg_0229 <= imem01_in[59:56];
    25: reg_0229 <= imem02_in[35:32];
    45: reg_0229 <= imem04_in[99:96];
    47: reg_0229 <= imem04_in[99:96];
    49: reg_0229 <= imem05_in[59:56];
    65: reg_0229 <= imem05_in[59:56];
    78: reg_0229 <= imem05_in[63:60];
    86: reg_0229 <= imem05_in[63:60];
    endcase
  end

  // REG#230の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0230 <= imem01_in[31:28];
    8: reg_0230 <= imem01_in[31:28];
    11: reg_0230 <= imem05_in[95:92];
    15: reg_0230 <= op2_01_out;
    41: reg_0230 <= op2_01_out;
    43: reg_0230 <= op2_01_out;
    50: reg_0230 <= imem02_in[115:112];
    51: reg_0230 <= op2_01_out;
    76: reg_0230 <= op2_01_out;
    endcase
  end

  // REG#231の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0231 <= op1_00_out;
    7: reg_0231 <= op1_00_out;
    8: reg_0231 <= op1_00_out;
    9: reg_0231 <= op1_00_out;
    10: reg_0231 <= op1_00_out;
    11: reg_0231 <= op1_00_out;
    12: reg_0231 <= op1_00_out;
    13: reg_0231 <= op1_00_out;
    14: reg_0231 <= op1_00_out;
    15: reg_0231 <= op1_00_out;
    16: reg_0231 <= op1_00_out;
    17: reg_0231 <= op1_00_out;
    18: reg_0231 <= op1_00_out;
    19: reg_0231 <= op1_00_out;
    20: reg_0231 <= op1_00_out;
    21: reg_0231 <= op1_00_out;
    22: reg_0231 <= op1_00_out;
    23: reg_0231 <= op1_00_out;
    24: reg_0231 <= op1_00_out;
    25: reg_0231 <= op1_00_out;
    26: reg_0231 <= op1_00_out;
    27: reg_0231 <= op1_00_out;
    28: reg_0231 <= op1_00_out;
    29: reg_0231 <= op1_00_out;
    30: reg_0231 <= op1_00_out;
    34: reg_0231 <= imem06_in[87:84];
    36: reg_0231 <= imem06_in[87:84];
    58: reg_0231 <= op1_00_out;
    59: reg_0231 <= op1_00_out;
    61: reg_0231 <= imem02_in[99:96];
    64: reg_0231 <= imem05_in[23:20];
    67: reg_0231 <= imem05_in[23:20];
    72: reg_0231 <= imem05_in[79:76];
    endcase
  end

  // REG#232の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0232 <= imem01_in[3:0];
    9: reg_0232 <= imem01_in[3:0];
    35: reg_0232 <= imem06_in[119:116];
    38: reg_0232 <= imem01_in[3:0];
    40: reg_0232 <= imem01_in[3:0];
    91: reg_0232 <= imem01_in[3:0];
    94: reg_0232 <= imem01_in[3:0];
    endcase
  end

  // REG#233の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0233 <= imem01_in[19:16];
    9: reg_0233 <= imem01_in[19:16];
    38: reg_0233 <= imem01_in[107:104];
    41: reg_0233 <= imem07_in[59:56];
    44: reg_0233 <= imem04_in[103:100];
    46: reg_0233 <= imem01_in[19:16];
    48: reg_0233 <= imem04_in[103:100];
    58: reg_0233 <= imem04_in[103:100];
    endcase
  end

  // REG#234の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0234 <= imem01_in[95:92];
    9: reg_0234 <= imem01_in[95:92];
    40: reg_0234 <= imem01_in[95:92];
    91: reg_0234 <= imem01_in[95:92];
    endcase
  end

  // REG#235の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0235 <= imem01_in[7:4];
    9: reg_0235 <= imem01_in[7:4];
    40: reg_0235 <= imem01_in[7:4];
    93: reg_0235 <= imem01_in[7:4];
    endcase
  end

  // REG#236の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0236 <= imem01_in[83:80];
    9: reg_0236 <= imem01_in[83:80];
    34: reg_0236 <= imem06_in[107:104];
    36: reg_0236 <= imem06_in[107:104];
    59: reg_0236 <= imem06_in[127:124];
    61: reg_0236 <= imem02_in[123:120];
    65: reg_0236 <= imem05_in[115:112];
    77: reg_0236 <= imem05_in[115:112];
    81: reg_0236 <= imem07_in[35:32];
    endcase
  end

  // REG#237の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0237 <= imem01_in[91:88];
    9: reg_0237 <= imem01_in[91:88];
    34: reg_0237 <= imem06_in[95:92];
    38: reg_0237 <= imem01_in[119:116];
    41: reg_0237 <= imem07_in[79:76];
    44: reg_0237 <= imem04_in[127:124];
    46: reg_0237 <= imem01_in[91:88];
    48: reg_0237 <= imem01_in[91:88];
    62: reg_0237 <= imem02_in[123:120];
    68: reg_0237 <= imem01_in[91:88];
    91: reg_0237 <= imem01_in[119:116];
    endcase
  end

  // REG#238の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0238 <= imem01_in[111:108];
    9: reg_0238 <= imem01_in[111:108];
    36: reg_0238 <= imem06_in[91:88];
    56: reg_0238 <= imem06_in[91:88];
    95: reg_0238 <= imem01_in[111:108];
    endcase
  end

  // REG#239の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0239 <= imem01_in[43:40];
    9: reg_0239 <= imem01_in[43:40];
    40: reg_0239 <= imem04_in[27:24];
    42: reg_0239 <= imem07_in[71:68];
    endcase
  end

  // REG#240の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0240 <= imem01_in[55:52];
    9: reg_0240 <= imem01_in[55:52];
    40: reg_0240 <= imem01_in[55:52];
    92: reg_0240 <= imem01_in[55:52];
    94: reg_0240 <= imem01_in[55:52];
    endcase
  end

  // REG#241の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0241 <= imem05_in[47:44];
    9: reg_0241 <= imem01_in[11:8];
    38: reg_0241 <= imem01_in[11:8];
    40: reg_0241 <= imem01_in[11:8];
    91: reg_0241 <= imem01_in[11:8];
    endcase
  end

  // REG#242の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0242 <= imem01_in[51:48];
    9: reg_0242 <= imem01_in[51:48];
    36: reg_0242 <= imem06_in[11:8];
    57: reg_0242 <= imem06_in[11:8];
    85: reg_0242 <= imem06_in[115:112];
    endcase
  end

  // REG#243の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0243 <= imem05_in[71:68];
    9: reg_0243 <= imem01_in[115:112];
    40: reg_0243 <= imem01_in[115:112];
    91: reg_0243 <= imem01_in[115:112];
    endcase
  end

  // REG#244の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0244 <= imem05_in[95:92];
    9: reg_0244 <= imem01_in[63:60];
    40: reg_0244 <= imem01_in[63:60];
    89: reg_0244 <= imem03_in[91:88];
    endcase
  end

  // REG#245の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0245 <= imem01_in[103:100];
    9: reg_0245 <= imem01_in[103:100];
    38: reg_0245 <= imem01_in[67:64];
    41: reg_0245 <= imem07_in[47:44];
    44: reg_0245 <= imem04_in[7:4];
    46: reg_0245 <= imem01_in[67:64];
    49: reg_0245 <= imem05_in[35:32];
    65: reg_0245 <= imem05_in[35:32];
    78: reg_0245 <= imem05_in[35:32];
    86: reg_0245 <= imem05_in[35:32];
    endcase
  end

  // REG#246の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0246 <= imem01_in[27:24];
    9: reg_0246 <= imem01_in[27:24];
    38: reg_0246 <= imem01_in[27:24];
    41: reg_0246 <= imem07_in[7:4];
    44: reg_0246 <= imem04_in[111:108];
    46: reg_0246 <= imem01_in[27:24];
    49: reg_0246 <= imem05_in[19:16];
    65: reg_0246 <= imem05_in[19:16];
    78: reg_0246 <= imem05_in[19:16];
    85: reg_0246 <= imem06_in[67:64];
    endcase
  end

  // REG#247の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0247 <= imem01_in[75:72];
    9: reg_0247 <= imem01_in[75:72];
    38: reg_0247 <= imem06_in[23:20];
    54: reg_0247 <= imem00_in[115:112];
    82: reg_0247 <= imem04_in[3:0];
    endcase
  end

  // REG#248の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0248 <= imem01_in[87:84];
    9: reg_0248 <= imem01_in[87:84];
    38: reg_0248 <= imem01_in[87:84];
    40: reg_0248 <= imem01_in[87:84];
    89: reg_0248 <= imem03_in[35:32];
    endcase
  end

  // REG#249の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0249 <= imem01_in[123:120];
    9: reg_0249 <= imem01_in[123:120];
    38: reg_0249 <= imem01_in[123:120];
    41: reg_0249 <= imem07_in[39:36];
    44: reg_0249 <= imem04_in[119:116];
    47: reg_0249 <= imem04_in[15:12];
    49: reg_0249 <= imem05_in[83:80];
    65: reg_0249 <= imem05_in[83:80];
    77: reg_0249 <= imem05_in[83:80];
    79: reg_0249 <= imem07_in[39:36];
    82: reg_0249 <= imem04_in[119:116];
    endcase
  end

  // REG#250の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0250 <= imem05_in[35:32];
    10: reg_0250 <= imem05_in[7:4];
    11: reg_0250 <= op2_01_out;
    27: reg_0250 <= op2_01_out;
    39: reg_0250 <= op2_01_out;
    79: reg_0250 <= op2_01_out;
    81: reg_0250 <= op2_01_out;
    87: reg_0250 <= op2_01_out;
    endcase
  end

  // REG#251の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0251 <= imem05_in[67:64];
    10: reg_0251 <= imem05_in[123:120];
    12: reg_0251 <= op2_02_out;
    31: reg_0251 <= op2_02_out;
    53: reg_0251 <= op2_02_out;
    83: reg_0251 <= imem02_in[127:124];
    96: reg_0251 <= op2_02_out;
    endcase
  end

  // REG#252の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0252 <= imem05_in[51:48];
    10: reg_0252 <= imem05_in[11:8];
    13: reg_0252 <= op2_02_out;
    35: reg_0252 <= op2_02_out;
    67: reg_0252 <= imem05_in[51:48];
    71: reg_0252 <= imem05_in[11:8];
    74: reg_0252 <= imem07_in[31:28];
    78: reg_0252 <= imem05_in[51:48];
    86: reg_0252 <= imem05_in[51:48];
    92: reg_0252 <= op2_02_out;
    endcase
  end

  // REG#253の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0253 <= imem05_in[115:112];
    10: reg_0253 <= imem05_in[55:52];
    17: reg_0253 <= imem04_in[31:28];
    42: reg_0253 <= imem07_in[15:12];
    endcase
  end

  // REG#254の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0254 <= imem05_in[103:100];
    10: reg_0254 <= imem05_in[3:0];
    17: reg_0254 <= imem04_in[63:60];
    44: reg_0254 <= imem02_in[27:24];
    49: reg_0254 <= op2_02_out;
    71: reg_0254 <= imem02_in[27:24];
    80: reg_0254 <= op2_02_out;
    86: reg_0254 <= imem05_in[103:100];
    93: reg_0254 <= op2_02_out;
    endcase
  end

  // REG#255の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0255 <= imem05_in[111:108];
    10: reg_0255 <= imem05_in[95:92];
    17: reg_0255 <= imem04_in[59:56];
    45: reg_0255 <= imem04_in[59:56];
    48: reg_0255 <= imem05_in[111:108];
    51: reg_0255 <= imem01_in[27:24];
    54: reg_0255 <= imem00_in[87:84];
    84: reg_0255 <= imem02_in[71:68];
    endcase
  end

  // REG#256の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0256 <= imem05_in[39:36];
    10: reg_0256 <= imem05_in[39:36];
    17: reg_0256 <= imem04_in[111:108];
    45: reg_0256 <= imem04_in[111:108];
    47: reg_0256 <= imem04_in[111:108];
    49: reg_0256 <= imem05_in[39:36];
    64: reg_0256 <= imem05_in[39:36];
    67: reg_0256 <= imem05_in[39:36];
    70: reg_0256 <= imem06_in[115:112];
    81: reg_0256 <= imem04_in[111:108];
    83: reg_0256 <= imem02_in[115:112];
    endcase
  end

  // REG#257の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0257 <= imem05_in[75:72];
    10: reg_0257 <= imem05_in[99:96];
    17: reg_0257 <= imem04_in[3:0];
    45: reg_0257 <= imem04_in[3:0];
    47: reg_0257 <= imem04_in[3:0];
    49: reg_0257 <= imem05_in[99:96];
    65: reg_0257 <= imem05_in[75:72];
    73: reg_0257 <= imem05_in[75:72];
    endcase
  end

  // REG#258の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0258 <= imem05_in[79:76];
    10: reg_0258 <= imem05_in[91:88];
    17: reg_0258 <= imem04_in[11:8];
    45: reg_0258 <= imem04_in[83:80];
    47: reg_0258 <= imem04_in[11:8];
    49: reg_0258 <= imem05_in[79:76];
    64: reg_0258 <= imem05_in[91:88];
    66: reg_0258 <= imem05_in[79:76];
    68: reg_0258 <= imem01_in[107:104];
    91: reg_0258 <= imem01_in[31:28];
    endcase
  end

  // REG#259の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0259 <= imem05_in[27:24];
    11: reg_0259 <= imem05_in[27:24];
    18: reg_0259 <= imem05_in[23:20];
    20: reg_0259 <= imem04_in[87:84];
    22: reg_0259 <= imem04_in[87:84];
    24: reg_0259 <= imem02_in[67:64];
    26: reg_0259 <= imem03_in[27:24];
    27: reg_0259 <= op1_14_out;
    30: reg_0259 <= imem03_in[27:24];
    50: reg_0259 <= op1_14_out;
    52: reg_0259 <= op1_14_out;
    55: reg_0259 <= imem05_in[23:20];
    58: reg_0259 <= imem04_in[87:84];
    endcase
  end

  // REG#260の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0260 <= imem05_in[83:80];
    11: reg_0260 <= imem05_in[83:80];
    19: reg_0260 <= imem05_in[83:80];
    48: reg_0260 <= imem05_in[23:20];
    51: reg_0260 <= imem01_in[75:72];
    54: reg_0260 <= imem05_in[83:80];
    56: reg_0260 <= imem06_in[127:124];
    94: reg_0260 <= imem01_in[75:72];
    endcase
  end

  // REG#261の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0261 <= imem05_in[107:104];
    11: reg_0261 <= imem05_in[107:104];
    16: reg_0261 <= op2_01_out;
    44: reg_0261 <= op2_01_out;
    53: reg_0261 <= op2_01_out;
    82: reg_0261 <= imem04_in[87:84];
    97: reg_0261 <= op2_01_out;
    endcase
  end

  // REG#262の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0262 <= imem05_in[19:16];
    11: reg_0262 <= imem05_in[19:16];
    18: reg_0262 <= imem05_in[115:112];
    20: reg_0262 <= imem04_in[7:4];
    21: reg_0262 <= op1_12_out;
    23: reg_0262 <= imem04_in[7:4];
    82: reg_0262 <= imem04_in[7:4];
    endcase
  end

  // REG#263の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0263 <= imem05_in[119:116];
    11: reg_0263 <= imem05_in[119:116];
    16: reg_0263 <= op2_02_out;
    45: reg_0263 <= op2_02_out;
    57: reg_0263 <= op2_02_out;
    95: reg_0263 <= op2_02_out;
    endcase
  end

  // REG#264の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0264 <= imem05_in[59:56];
    11: reg_0264 <= imem05_in[79:76];
    18: reg_0264 <= imem05_in[127:124];
    20: reg_0264 <= imem04_in[31:28];
    22: reg_0264 <= imem04_in[75:72];
    24: reg_0264 <= imem02_in[51:48];
    26: reg_0264 <= imem03_in[83:80];
    27: reg_0264 <= op2_02_out;
    40: reg_0264 <= op2_02_out;
    83: reg_0264 <= imem02_in[51:48];
    endcase
  end

  // REG#265の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0265 <= imem05_in[91:88];
    11: reg_0265 <= imem05_in[91:88];
    18: reg_0265 <= imem04_in[71:68];
    38: reg_0265 <= imem06_in[119:116];
    54: reg_0265 <= imem05_in[91:88];
    56: reg_0265 <= imem06_in[119:116];
    endcase
  end

  // REG#266の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0266 <= imem05_in[123:120];
    11: reg_0266 <= imem05_in[123:120];
    18: reg_0266 <= imem04_in[111:108];
    40: reg_0266 <= imem04_in[79:76];
    42: reg_0266 <= imem07_in[19:16];
    endcase
  end

  // REG#267の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0267 <= imem05_in[3:0];
    11: reg_0267 <= imem05_in[3:0];
    18: reg_0267 <= imem04_in[83:80];
    40: reg_0267 <= imem04_in[19:16];
    42: reg_0267 <= imem07_in[111:108];
    endcase
  end

  // REG#268の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0268 <= imem05_in[7:4];
    11: reg_0268 <= imem05_in[7:4];
    18: reg_0268 <= imem04_in[87:84];
    40: reg_0268 <= imem04_in[103:100];
    42: reg_0268 <= imem07_in[127:124];
    endcase
  end

  // REG#269の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0269 <= imem05_in[87:84];
    11: reg_0269 <= imem05_in[87:84];
    19: reg_0269 <= imem05_in[87:84];
    49: reg_0269 <= imem05_in[87:84];
    59: reg_0269 <= imem05_in[87:84];
    60: reg_0269 <= op2_01_out;
    63: reg_0269 <= imem05_in[87:84];
    64: reg_0269 <= op2_01_out;
    74: reg_0269 <= op2_01_out;
    endcase
  end

  // REG#270の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0270 <= imem05_in[43:40];
    11: reg_0270 <= imem05_in[43:40];
    18: reg_0270 <= imem05_in[43:40];
    20: reg_0270 <= imem04_in[51:48];
    22: reg_0270 <= imem04_in[51:48];
    24: reg_0270 <= imem02_in[19:16];
    26: reg_0270 <= imem03_in[111:108];
    28: reg_0270 <= imem06_in[83:80];
    52: reg_0270 <= imem03_in[111:108];
    55: reg_0270 <= imem05_in[43:40];
    57: reg_0270 <= imem06_in[83:80];
    85: reg_0270 <= imem06_in[83:80];
    90: reg_0270 <= op2_02_out;
    endcase
  end

  // REG#271の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0271 <= imem05_in[23:20];
    11: reg_0271 <= imem05_in[23:20];
    19: reg_0271 <= imem05_in[23:20];
    46: reg_0271 <= op2_03_out;
    61: reg_0271 <= op2_03_out;
    67: reg_0271 <= imem01_in[87:84];
    68: reg_0271 <= op2_03_out;
    89: reg_0271 <= imem03_in[7:4];
    endcase
  end

  // REG#272の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0272 <= imem05_in[99:96];
    11: reg_0272 <= imem05_in[99:96];
    19: reg_0272 <= imem05_in[99:96];
    48: reg_0272 <= imem05_in[75:72];
    50: reg_0272 <= op2_01_out;
    72: reg_0272 <= op2_01_out;
    endcase
  end

  // REG#273の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0273 <= imem05_in[31:28];
    11: reg_0273 <= imem05_in[31:28];
    18: reg_0273 <= imem04_in[39:36];
    39: reg_0273 <= op2_00_out;
    77: reg_0273 <= op2_00_out;
    endcase
  end

  // REG#274の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0274 <= imem05_in[55:52];
    11: reg_0274 <= imem05_in[55:52];
    18: reg_0274 <= imem04_in[47:44];
    39: reg_0274 <= op2_02_out;
    79: reg_0274 <= op2_02_out;
    83: reg_0274 <= imem02_in[119:116];
    endcase
  end

  // REG#275の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0275 <= imem04_in[111:108];
    16: reg_0275 <= imem04_in[111:108];
    19: reg_0275 <= imem05_in[55:52];
    48: reg_0275 <= imem04_in[111:108];
    57: reg_0275 <= imem04_in[35:32];
    59: reg_0275 <= imem05_in[15:12];
    62: reg_0275 <= imem02_in[127:124];
    69: reg_0275 <= imem06_in[43:40];
    71: reg_0275 <= imem02_in[127:124];
    82: reg_0275 <= imem04_in[35:32];
    endcase
  end

  // REG#276の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0276 <= imem04_in[71:68];
    16: reg_0276 <= imem04_in[71:68];
    19: reg_0276 <= imem05_in[67:64];
    49: reg_0276 <= imem05_in[67:64];
    65: reg_0276 <= imem05_in[67:64];
    74: reg_0276 <= imem07_in[99:96];
    78: reg_0276 <= imem05_in[67:64];
    85: reg_0276 <= imem06_in[51:48];
    endcase
  end

  // REG#277の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0277 <= imem04_in[47:44];
    16: reg_0277 <= imem04_in[47:44];
    19: reg_0277 <= imem05_in[107:104];
    49: reg_0277 <= imem05_in[107:104];
    64: reg_0277 <= imem05_in[107:104];
    67: reg_0277 <= imem05_in[107:104];
    71: reg_0277 <= imem05_in[107:104];
    74: reg_0277 <= imem07_in[71:68];
    78: reg_0277 <= imem05_in[107:104];
    86: reg_0277 <= imem05_in[107:104];
    endcase
  end

  // REG#278の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0278 <= imem04_in[127:124];
    18: reg_0278 <= imem04_in[127:124];
    38: reg_0278 <= imem06_in[123:120];
    55: reg_0278 <= imem05_in[79:76];
    60: reg_0278 <= imem05_in[79:76];
    65: reg_0278 <= imem05_in[79:76];
    74: reg_0278 <= imem07_in[15:12];
    78: reg_0278 <= imem05_in[79:76];
    85: reg_0278 <= imem05_in[79:76];
    87: reg_0278 <= imem06_in[123:120];
    89: reg_0278 <= imem03_in[83:80];
    endcase
  end

  // REG#279の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0279 <= imem04_in[31:28];
    16: reg_0279 <= imem04_in[31:28];
    19: reg_0279 <= imem05_in[39:36];
    49: reg_0279 <= imem05_in[71:68];
    65: reg_0279 <= imem05_in[39:36];
    74: reg_0279 <= imem07_in[107:104];
    77: reg_0279 <= imem05_in[39:36];
    81: reg_0279 <= imem07_in[107:104];
    endcase
  end

  // REG#280の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0280 <= op1_01_out;
    18: reg_0280 <= imem04_in[31:28];
    41: reg_0280 <= imem04_in[31:28];
    endcase
  end

  // REG#281の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0281 <= imem04_in[15:12];
    17: reg_0281 <= imem04_in[15:12];
    43: reg_0281 <= op2_03_out;
    52: reg_0281 <= imem03_in[103:100];
    54: reg_0281 <= imem03_in[103:100];
    84: reg_0281 <= imem02_in[23:20];
    endcase
  end

  // REG#282の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0282 <= imem04_in[51:48];
    16: reg_0282 <= imem04_in[51:48];
    19: reg_0282 <= imem05_in[79:76];
    48: reg_0282 <= op2_01_out;
    67: reg_0282 <= imem05_in[79:76];
    71: reg_0282 <= imem05_in[79:76];
    73: reg_0282 <= op2_01_out;
    endcase
  end

  // REG#283の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0283 <= imem04_in[23:20];
    16: reg_0283 <= imem04_in[23:20];
    18: reg_0283 <= imem04_in[23:20];
    41: reg_0283 <= imem04_in[23:20];
    endcase
  end

  // REG#284の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0284 <= imem04_in[123:120];
    16: reg_0284 <= imem04_in[123:120];
    18: reg_0284 <= imem04_in[123:120];
    35: reg_0284 <= op2_00_out;
    64: reg_0284 <= op2_00_out;
    73: reg_0284 <= op2_00_out;
    endcase
  end

  // REG#285の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0285 <= imem04_in[83:80];
    16: reg_0285 <= imem04_in[83:80];
    19: reg_0285 <= imem05_in[119:116];
    49: reg_0285 <= imem05_in[119:116];
    65: reg_0285 <= imem05_in[119:116];
    78: reg_0285 <= imem05_in[119:116];
    86: reg_0285 <= imem05_in[119:116];
    endcase
  end

  // REG#286の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0286 <= imem04_in[103:100];
    18: reg_0286 <= imem04_in[103:100];
    34: reg_0286 <= imem06_in[63:60];
    38: reg_0286 <= imem06_in[63:60];
    55: reg_0286 <= imem06_in[63:60];
    57: reg_0286 <= op2_00_out;
    97: reg_0286 <= op2_00_out;
    endcase
  end

  // REG#287の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0287 <= op1_02_out;
    17: reg_0287 <= op2_00_out;
    46: reg_0287 <= op2_00_out;
    58: reg_0287 <= op2_00_out;
    endcase
  end

  // REG#288の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0288 <= imem04_in[115:112];
    17: reg_0288 <= imem04_in[115:112];
    41: reg_0288 <= imem07_in[3:0];
    44: reg_0288 <= imem04_in[115:112];
    48: reg_0288 <= imem04_in[115:112];
    55: reg_0288 <= imem05_in[67:64];
    60: reg_0288 <= imem05_in[83:80];
    63: reg_0288 <= imem05_in[67:64];
    65: reg_0288 <= imem05_in[71:68];
    78: reg_0288 <= imem05_in[83:80];
    86: reg_0288 <= imem05_in[83:80];
    endcase
  end

  // REG#289の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0289 <= imem04_in[55:52];
    17: reg_0289 <= imem04_in[55:52];
    38: reg_0289 <= imem06_in[3:0];
    56: reg_0289 <= imem06_in[3:0];
    endcase
  end

  // REG#290の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0290 <= imem04_in[75:72];
    18: reg_0290 <= imem04_in[75:72];
    40: reg_0290 <= imem01_in[75:72];
    87: reg_0290 <= imem06_in[95:92];
    89: reg_0290 <= imem03_in[87:84];
    endcase
  end

  // REG#291の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0291 <= imem04_in[79:76];
    18: reg_0291 <= imem04_in[79:76];
    38: reg_0291 <= imem06_in[27:24];
    56: reg_0291 <= imem06_in[27:24];
    endcase
  end

  // REG#292の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0292 <= imem04_in[95:92];
    18: reg_0292 <= imem04_in[95:92];
    41: reg_0292 <= imem04_in[95:92];
    endcase
  end

  // REG#293の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0293 <= imem04_in[67:64];
    18: reg_0293 <= imem04_in[67:64];
    34: reg_0293 <= imem06_in[115:112];
    38: reg_0293 <= imem06_in[115:112];
    56: reg_0293 <= imem06_in[115:112];
    endcase
  end

  // REG#294の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0294 <= imem04_in[43:40];
    18: reg_0294 <= imem04_in[43:40];
    40: reg_0294 <= imem01_in[79:76];
    89: reg_0294 <= imem03_in[75:72];
    endcase
  end

  // REG#295の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0295 <= imem04_in[99:96];
    18: reg_0295 <= imem04_in[99:96];
    40: reg_0295 <= imem04_in[99:96];
    42: reg_0295 <= imem07_in[23:20];
    endcase
  end

  // REG#296の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0296 <= imem04_in[87:84];
    17: reg_0296 <= imem04_in[87:84];
    44: reg_0296 <= imem04_in[87:84];
    48: reg_0296 <= imem04_in[87:84];
    58: reg_0296 <= imem04_in[95:92];
    endcase
  end

  // REG#297の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0297 <= imem04_in[91:88];
    18: reg_0297 <= imem04_in[91:88];
    41: reg_0297 <= imem04_in[91:88];
    endcase
  end

  // REG#298の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0298 <= imem04_in[107:104];
    18: reg_0298 <= imem04_in[107:104];
    38: reg_0298 <= imem06_in[75:72];
    56: reg_0298 <= imem06_in[75:72];
    endcase
  end

  // REG#299の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0299 <= imem04_in[39:36];
    17: reg_0299 <= imem04_in[39:36];
    38: reg_0299 <= imem06_in[11:8];
    56: reg_0299 <= imem06_in[11:8];
    endcase
  end

  // REG#300の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0300 <= imem04_in[35:32];
    17: reg_0300 <= op2_02_out;
    48: reg_0300 <= op2_02_out;
    67: reg_0300 <= op2_02_out;
    84: reg_0300 <= op2_02_out;
    endcase
  end

  // REG#301の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0301 <= imem04_in[19:16];
    18: reg_0301 <= imem04_in[19:16];
    41: reg_0301 <= imem07_in[67:64];
    44: reg_0301 <= imem02_in[79:76];
    58: reg_0301 <= imem04_in[19:16];
    endcase
  end

  // REG#302の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0302 <= imem04_in[63:60];
    18: reg_0302 <= imem04_in[63:60];
    41: reg_0302 <= imem04_in[63:60];
    endcase
  end

  // REG#303の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0303 <= imem04_in[3:0];
    18: reg_0303 <= imem04_in[3:0];
    41: reg_0303 <= imem04_in[3:0];
    endcase
  end

  // REG#304の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0304 <= imem04_in[11:8];
    19: reg_0304 <= imem05_in[27:24];
    49: reg_0304 <= imem05_in[27:24];
    64: reg_0304 <= imem05_in[27:24];
    67: reg_0304 <= imem01_in[91:88];
    69: reg_0304 <= imem06_in[91:88];
    71: reg_0304 <= imem02_in[91:88];
    81: reg_0304 <= imem04_in[11:8];
    83: reg_0304 <= imem02_in[91:88];
    94: reg_0304 <= imem01_in[91:88];
    endcase
  end

  // REG#305の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0305 <= imem04_in[27:24];
    18: reg_0305 <= imem04_in[27:24];
    41: reg_0305 <= imem04_in[27:24];
    endcase
  end

  // REG#306の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0306 <= imem04_in[59:56];
    18: reg_0306 <= imem04_in[59:56];
    40: reg_0306 <= imem01_in[27:24];
    89: reg_0306 <= imem03_in[71:68];
    endcase
  end

  // REG#307の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0307 <= imem04_in[119:116];
    19: reg_0307 <= imem05_in[91:88];
    49: reg_0307 <= imem05_in[91:88];
    65: reg_0307 <= imem05_in[91:88];
    78: reg_0307 <= imem05_in[91:88];
    85: reg_0307 <= imem06_in[63:60];
    endcase
  end

  // REG#308の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0308 <= imem04_in[7:4];
    18: reg_0308 <= imem04_in[7:4];
    41: reg_0308 <= imem04_in[7:4];
    endcase
  end

  // REG#309の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0309 <= imem03_in[115:112];
    19: reg_0309 <= imem05_in[31:28];
    49: reg_0309 <= imem05_in[31:28];
    65: reg_0309 <= imem05_in[31:28];
    78: reg_0309 <= imem05_in[31:28];
    86: reg_0309 <= imem05_in[31:28];
    endcase
  end

  // REG#310の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0310 <= imem02_in[87:84];
    18: reg_0310 <= op2_00_out;
    49: reg_0310 <= op2_00_out;
    68: reg_0310 <= op2_00_out;
    85: reg_0310 <= op2_00_out;
    endcase
  end

  // REG#311の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0311 <= imem03_in[35:32];
    20: reg_0311 <= imem04_in[123:120];
    22: reg_0311 <= imem04_in[123:120];
    24: reg_0311 <= imem02_in[115:112];
    26: reg_0311 <= imem03_in[123:120];
    28: reg_0311 <= imem06_in[127:124];
    52: reg_0311 <= imem03_in[123:120];
    55: reg_0311 <= imem06_in[127:124];
    58: reg_0311 <= imem04_in[67:64];
    endcase
  end

  // REG#312の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0312 <= imem03_in[95:92];
    19: reg_0312 <= op2_01_out;
    54: reg_0312 <= op2_01_out;
    84: reg_0312 <= op2_01_out;
    endcase
  end

  // REG#313の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0313 <= imem06_in[71:68];
    19: reg_0313 <= op2_02_out;
    55: reg_0313 <= op2_02_out;
    88: reg_0313 <= op2_02_out;
    endcase
  end

  // REG#314の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0314 <= imem02_in[119:116];
    20: reg_0314 <= imem02_in[15:12];
    78: reg_0314 <= imem05_in[95:92];
    84: reg_0314 <= imem02_in[15:12];
    endcase
  end

  // REG#315の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0315 <= imem06_in[99:96];
    21: reg_0315 <= imem04_in[23:20];
    23: reg_0315 <= imem04_in[23:20];
    78: reg_0315 <= imem05_in[23:20];
    84: reg_0315 <= imem02_in[99:96];
    endcase
  end

  // REG#316の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0316 <= op1_03_out;
    21: reg_0316 <= imem04_in[15:12];
    23: reg_0316 <= imem04_in[15:12];
    82: reg_0316 <= imem04_in[15:12];
    endcase
  end

  // REG#317の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0317 <= imem03_in[39:36];
    22: reg_0317 <= imem04_in[115:112];
    24: reg_0317 <= imem02_in[31:28];
    26: reg_0317 <= imem03_in[19:16];
    28: reg_0317 <= imem06_in[19:16];
    54: reg_0317 <= imem03_in[19:16];
    86: reg_0317 <= imem03_in[23:20];
    88: reg_0317 <= imem03_in[23:20];
    endcase
  end

  // REG#318の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0318 <= imem02_in[59:56];
    22: reg_0318 <= imem04_in[83:80];
    24: reg_0318 <= imem02_in[59:56];
    26: reg_0318 <= imem03_in[71:68];
    28: reg_0318 <= imem06_in[11:8];
    54: reg_0318 <= imem03_in[71:68];
    87: reg_0318 <= imem03_in[71:68];
    endcase
  end

  // REG#319の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0319 <= imem03_in[59:56];
    22: reg_0319 <= imem04_in[3:0];
    24: reg_0319 <= imem02_in[43:40];
    26: reg_0319 <= imem03_in[59:56];
    28: reg_0319 <= imem06_in[103:100];
    54: reg_0319 <= imem03_in[59:56];
    87: reg_0319 <= imem06_in[103:100];
    89: reg_0319 <= imem03_in[59:56];
    endcase
  end

  // REG#320の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0320 <= imem02_in[31:28];
    23: reg_0320 <= imem01_in[63:60];
    25: reg_0320 <= imem02_in[31:28];
    51: reg_0320 <= imem02_in[31:28];
    endcase
  end

  // REG#321の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0321 <= imem03_in[23:20];
    23: reg_0321 <= imem01_in[119:116];
    25: reg_0321 <= imem02_in[119:116];
    48: reg_0321 <= imem01_in[119:116];
    67: reg_0321 <= imem01_in[119:116];
    69: reg_0321 <= imem03_in[23:20];
    endcase
  end

  // REG#322の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0322 <= imem03_in[79:76];
    23: reg_0322 <= imem01_in[67:64];
    25: reg_0322 <= imem02_in[99:96];
    48: reg_0322 <= imem01_in[67:64];
    67: reg_0322 <= imem05_in[119:116];
    70: reg_0322 <= imem06_in[27:24];
    83: reg_0322 <= imem02_in[99:96];
    endcase
  end

  // REG#323の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0323 <= imem03_in[83:80];
    23: reg_0323 <= imem01_in[71:68];
    25: reg_0323 <= imem02_in[127:124];
    48: reg_0323 <= imem05_in[107:104];
    51: reg_0323 <= imem02_in[127:124];
    endcase
  end

  // REG#324の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0324 <= imem02_in[79:76];
    23: reg_0324 <= imem01_in[103:100];
    25: reg_0324 <= imem02_in[79:76];
    51: reg_0324 <= imem02_in[79:76];
    93: reg_0324 <= imem01_in[103:100];
    endcase
  end

  // REG#325の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0325 <= imem02_in[23:20];
    22: reg_0325 <= op2_00_out;
    63: reg_0325 <= op2_00_out;
    71: reg_0325 <= imem02_in[23:20];
    81: reg_0325 <= imem07_in[83:80];
    endcase
  end

  // REG#326の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0326 <= imem02_in[35:32];
    22: reg_0326 <= op2_01_out;
    65: reg_0326 <= imem05_in[7:4];
    78: reg_0326 <= imem05_in[7:4];
    86: reg_0326 <= imem05_in[7:4];
    endcase
  end

  // REG#327の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0327 <= imem03_in[71:68];
    22: reg_0327 <= op2_02_out;
    65: reg_0327 <= op2_02_out;
    81: reg_0327 <= imem07_in[47:44];
    endcase
  end

  // REG#328の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0328 <= imem02_in[115:112];
    23: reg_0328 <= imem04_in[35:32];
    73: reg_0328 <= imem07_in[55:52];
    78: reg_0328 <= imem05_in[39:36];
    85: reg_0328 <= imem06_in[107:104];
    endcase
  end

  // REG#329の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0329 <= imem02_in[55:52];
    24: reg_0329 <= imem02_in[79:76];
    26: reg_0329 <= imem03_in[87:84];
    28: reg_0329 <= imem06_in[99:96];
    54: reg_0329 <= imem03_in[87:84];
    86: reg_0329 <= imem03_in[51:48];
    88: reg_0329 <= imem03_in[51:48];
    endcase
  end

  // REG#330の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0330 <= imem02_in[63:60];
    24: reg_0330 <= imem02_in[123:120];
    25: reg_0330 <= op2_00_out;
    31: reg_0330 <= op2_00_out;
    51: reg_0330 <= op2_00_out;
    74: reg_0330 <= op2_00_out;
    endcase
  end

  // REG#331の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0331 <= imem03_in[127:124];
    23: reg_0331 <= op2_01_out;
    26: reg_0331 <= imem03_in[127:124];
    28: reg_0331 <= imem06_in[27:24];
    54: reg_0331 <= imem03_in[127:124];
    82: reg_0331 <= imem04_in[107:104];
    endcase
  end

  // REG#332の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0332 <= imem06_in[11:8];
    23: reg_0332 <= op2_02_out;
    26: reg_0332 <= op2_02_out;
    36: reg_0332 <= op2_02_out;
    69: reg_0332 <= op2_02_out;
    endcase
  end

  // REG#333の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0333 <= imem02_in[11:8];
    24: reg_0333 <= imem01_in[87:84];
    42: reg_0333 <= imem07_in[59:56];
    endcase
  end

  // REG#334の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0334 <= imem02_in[7:4];
    24: reg_0334 <= imem01_in[55:52];
    42: reg_0334 <= imem07_in[3:0];
    endcase
  end

  // REG#335の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0335 <= imem02_in[111:108];
    24: reg_0335 <= imem02_in[111:108];
    25: reg_0335 <= op2_01_out;
    32: reg_0335 <= op2_01_out;
    55: reg_0335 <= op2_01_out;
    88: reg_0335 <= imem06_in[27:24];
    endcase
  end

  // REG#336の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0336 <= imem02_in[127:124];
    24: reg_0336 <= imem01_in[7:4];
    44: reg_0336 <= imem02_in[127:124];
    59: reg_0336 <= imem05_in[35:32];
    61: reg_0336 <= imem02_in[127:124];
    63: reg_0336 <= imem05_in[35:32];
    66: reg_0336 <= imem05_in[35:32];
    68: reg_0336 <= imem01_in[7:4];
    endcase
  end

  // REG#337の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0337 <= imem06_in[119:116];
    24: reg_0337 <= imem01_in[43:40];
    44: reg_0337 <= imem02_in[11:8];
    60: reg_0337 <= imem05_in[19:16];
    64: reg_0337 <= imem05_in[19:16];
    67: reg_0337 <= imem05_in[19:16];
    72: reg_0337 <= imem05_in[11:8];
    endcase
  end

  // REG#338の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0338 <= imem02_in[99:96];
    24: reg_0338 <= imem02_in[99:96];
    27: reg_0338 <= imem06_in[63:60];
    29: reg_0338 <= imem03_in[43:40];
    31: reg_0338 <= imem06_in[63:60];
    36: reg_0338 <= imem06_in[63:60];
    54: reg_0338 <= imem03_in[43:40];
    87: reg_0338 <= imem03_in[43:40];
    endcase
  end

  // REG#339の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0339 <= imem02_in[71:68];
    24: reg_0339 <= imem02_in[71:68];
    27: reg_0339 <= imem06_in[107:104];
    29: reg_0339 <= imem03_in[71:68];
    31: reg_0339 <= imem06_in[107:104];
    38: reg_0339 <= imem06_in[107:104];
    56: reg_0339 <= imem06_in[107:104];
    endcase
  end

  // REG#340の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0340 <= op1_04_out;
    23: reg_0340 <= op1_04_out;
    24: reg_0340 <= op1_04_out;
    25: reg_0340 <= op1_04_out;
    26: reg_0340 <= op1_04_out;
    27: reg_0340 <= op1_04_out;
    28: reg_0340 <= op1_04_out;
    29: reg_0340 <= op1_04_out;
    30: reg_0340 <= op1_04_out;
    31: reg_0340 <= op1_04_out;
    32: reg_0340 <= op1_04_out;
    33: reg_0340 <= op1_04_out;
    34: reg_0340 <= op1_04_out;
    35: reg_0340 <= op1_04_out;
    36: reg_0340 <= op1_04_out;
    37: reg_0340 <= op1_04_out;
    38: reg_0340 <= op1_04_out;
    39: reg_0340 <= op1_04_out;
    40: reg_0340 <= op1_04_out;
    41: reg_0340 <= op1_04_out;
    42: reg_0340 <= op1_04_out;
    43: reg_0340 <= op1_04_out;
    44: reg_0340 <= op1_04_out;
    45: reg_0340 <= op1_04_out;
    46: reg_0340 <= op1_04_out;
    47: reg_0340 <= op1_04_out;
    48: reg_0340 <= op1_04_out;
    49: reg_0340 <= op1_04_out;
    50: reg_0340 <= op1_04_out;
    51: reg_0340 <= op1_04_out;
    52: reg_0340 <= op1_04_out;
    53: reg_0340 <= op1_04_out;
    54: reg_0340 <= op1_04_out;
    55: reg_0340 <= op1_04_out;
    56: reg_0340 <= op1_04_out;
    57: reg_0340 <= op1_04_out;
    58: reg_0340 <= op1_04_out;
    59: reg_0340 <= op1_04_out;
    60: reg_0340 <= op1_04_out;
    61: reg_0340 <= op1_04_out;
    62: reg_0340 <= op1_04_out;
    63: reg_0340 <= op1_04_out;
    64: reg_0340 <= op1_04_out;
    65: reg_0340 <= op1_04_out;
    66: reg_0340 <= op1_04_out;
    67: reg_0340 <= op1_04_out;
    68: reg_0340 <= op1_04_out;
    69: reg_0340 <= op1_04_out;
    70: reg_0340 <= op1_04_out;
    71: reg_0340 <= op1_04_out;
    72: reg_0340 <= op1_04_out;
    73: reg_0340 <= op1_04_out;
    74: reg_0340 <= op1_04_out;
    75: reg_0340 <= op1_04_out;
    76: reg_0340 <= op1_04_out;
    77: reg_0340 <= op1_04_out;
    78: reg_0340 <= op1_04_out;
    79: reg_0340 <= op1_04_out;
    80: reg_0340 <= op1_04_out;
    81: reg_0340 <= op1_04_out;
    82: reg_0340 <= op1_04_out;
    83: reg_0340 <= op1_04_out;
    84: reg_0340 <= op1_04_out;
    85: reg_0340 <= op1_04_out;
    86: reg_0340 <= op1_04_out;
    87: reg_0340 <= op1_04_out;
    88: reg_0340 <= op1_04_out;
    89: reg_0340 <= op1_04_out;
    90: reg_0340 <= op1_04_out;
    91: reg_0340 <= op1_04_out;
    92: reg_0340 <= op1_04_out;
    93: reg_0340 <= op1_04_out;
    94: reg_0340 <= op1_04_out;
    95: reg_0340 <= op1_04_out;
    96: reg_0340 <= op1_04_out;
    endcase
  end

  // REG#341の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0341 <= imem02_in[43:40];
    25: reg_0341 <= imem02_in[43:40];
    51: reg_0341 <= imem02_in[43:40];
    endcase
  end

  // REG#342の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0342 <= imem02_in[95:92];
    25: reg_0342 <= imem02_in[95:92];
    51: reg_0342 <= imem02_in[95:92];
    endcase
  end

  // REG#343の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0343 <= imem03_in[43:40];
    25: reg_0343 <= imem02_in[115:112];
    48: reg_0343 <= imem04_in[11:8];
    51: reg_0343 <= imem02_in[115:112];
    endcase
  end

  // REG#344の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0344 <= imem06_in[23:20];
    25: reg_0344 <= imem02_in[11:8];
    51: reg_0344 <= imem02_in[11:8];
    endcase
  end

  // REG#345の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0345 <= imem02_in[51:48];
    25: reg_0345 <= imem02_in[51:48];
    51: reg_0345 <= imem02_in[51:48];
    endcase
  end

  // REG#346の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0346 <= imem02_in[75:72];
    25: reg_0346 <= imem02_in[75:72];
    44: reg_0346 <= imem02_in[75:72];
    56: reg_0346 <= imem06_in[19:16];
    endcase
  end

  // REG#347の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0347 <= imem02_in[123:120];
    25: reg_0347 <= imem02_in[123:120];
    50: reg_0347 <= imem02_in[123:120];
    52: reg_0347 <= imem03_in[43:40];
    54: reg_0347 <= imem03_in[11:8];
    86: reg_0347 <= imem03_in[127:124];
    88: reg_0347 <= imem03_in[43:40];
    endcase
  end

  // REG#348の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0348 <= imem06_in[7:4];
    25: reg_0348 <= imem02_in[55:52];
    50: reg_0348 <= imem02_in[55:52];
    52: reg_0348 <= imem03_in[7:4];
    56: reg_0348 <= imem06_in[7:4];
    endcase
  end

  // REG#349の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0349 <= imem06_in[39:36];
    25: reg_0349 <= imem02_in[7:4];
    50: reg_0349 <= imem02_in[7:4];
    52: reg_0349 <= imem03_in[47:44];
    56: reg_0349 <= imem06_in[39:36];
    endcase
  end

  // REG#350の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0350 <= imem02_in[107:104];
    25: reg_0350 <= imem02_in[107:104];
    48: reg_0350 <= imem04_in[95:92];
    54: reg_0350 <= imem03_in[83:80];
    85: reg_0350 <= op1_12_out;
    88: reg_0350 <= imem03_in[83:80];
    endcase
  end

  // REG#351の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0351 <= imem06_in[51:48];
    25: reg_0351 <= imem02_in[87:84];
    51: reg_0351 <= imem02_in[87:84];
    85: reg_0351 <= op1_13_out;
    88: reg_0351 <= imem06_in[51:48];
    endcase
  end

  // REG#352の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0352 <= imem02_in[3:0];
    25: reg_0352 <= imem02_in[3:0];
    51: reg_0352 <= imem02_in[3:0];
    endcase
  end

  // REG#353の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0353 <= imem02_in[83:80];
    25: reg_0353 <= imem02_in[83:80];
    45: reg_0353 <= imem04_in[107:104];
    47: reg_0353 <= imem04_in[107:104];
    51: reg_0353 <= imem02_in[83:80];
    endcase
  end

  // REG#354の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0354 <= imem02_in[39:36];
    25: reg_0354 <= imem02_in[39:36];
    50: reg_0354 <= imem02_in[39:36];
    52: reg_0354 <= imem03_in[71:68];
    56: reg_0354 <= imem06_in[87:84];
    endcase
  end

  // REG#355の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0355 <= imem02_in[103:100];
    25: reg_0355 <= imem02_in[103:100];
    41: reg_0355 <= imem07_in[111:108];
    44: reg_0355 <= imem02_in[103:100];
    62: reg_0355 <= imem02_in[103:100];
    70: reg_0355 <= imem02_in[103:100];
    72: reg_0355 <= imem05_in[99:96];
    endcase
  end

  // REG#356の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0356 <= imem06_in[19:16];
    25: reg_0356 <= imem02_in[63:60];
    51: reg_0356 <= imem02_in[63:60];
    endcase
  end

  // REG#357の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0357 <= imem02_in[15:12];
    25: reg_0357 <= imem02_in[15:12];
    48: reg_0357 <= imem04_in[3:0];
    54: reg_0357 <= imem03_in[107:104];
    85: reg_0357 <= op1_14_out;
    88: reg_0357 <= imem03_in[107:104];
    89: reg_0357 <= op1_14_out;
    91: reg_0357 <= op1_14_out;
    endcase
  end

  // REG#358の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0358 <= imem02_in[19:16];
    25: reg_0358 <= imem02_in[19:16];
    51: reg_0358 <= imem02_in[19:16];
    endcase
  end

  // REG#359の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0359 <= imem02_in[47:44];
    25: reg_0359 <= imem02_in[47:44];
    51: reg_0359 <= imem02_in[47:44];
    endcase
  end

  // REG#360の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0360 <= imem03_in[27:24];
    25: reg_0360 <= imem02_in[71:68];
    51: reg_0360 <= imem02_in[71:68];
    endcase
  end

  // REG#361の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0361 <= imem03_in[107:104];
    25: reg_0361 <= imem02_in[59:56];
    51: reg_0361 <= imem02_in[59:56];
    endcase
  end

  // REG#362の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0362 <= imem03_in[51:48];
    25: reg_0362 <= imem02_in[23:20];
    51: reg_0362 <= imem02_in[23:20];
    endcase
  end

  // REG#363の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0363 <= imem02_in[67:64];
    25: reg_0363 <= imem02_in[67:64];
    51: reg_0363 <= imem02_in[67:64];
    endcase
  end

  // REG#364の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0364 <= imem02_in[27:24];
    25: reg_0364 <= imem02_in[27:24];
    51: reg_0364 <= imem02_in[27:24];
    endcase
  end

  // REG#365の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0365 <= imem02_in[91:88];
    25: reg_0365 <= imem02_in[91:88];
    51: reg_0365 <= imem02_in[91:88];
    endcase
  end

  // REG#366の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0366 <= op1_05_out;
    24: reg_0366 <= op1_05_out;
    25: reg_0366 <= op1_05_out;
    26: reg_0366 <= op1_05_out;
    27: reg_0366 <= op1_05_out;
    28: reg_0366 <= op1_05_out;
    29: reg_0366 <= op1_05_out;
    30: reg_0366 <= op1_05_out;
    31: reg_0366 <= op1_05_out;
    32: reg_0366 <= op1_05_out;
    33: reg_0366 <= op1_05_out;
    34: reg_0366 <= op1_05_out;
    35: reg_0366 <= op1_05_out;
    36: reg_0366 <= op1_05_out;
    37: reg_0366 <= op1_05_out;
    38: reg_0366 <= op1_05_out;
    39: reg_0366 <= op1_05_out;
    40: reg_0366 <= op1_05_out;
    41: reg_0366 <= op1_05_out;
    42: reg_0366 <= op1_05_out;
    43: reg_0366 <= op1_05_out;
    44: reg_0366 <= op1_05_out;
    45: reg_0366 <= op1_05_out;
    46: reg_0366 <= op1_05_out;
    47: reg_0366 <= op1_05_out;
    48: reg_0366 <= op1_05_out;
    49: reg_0366 <= op1_05_out;
    50: reg_0366 <= op1_05_out;
    51: reg_0366 <= op1_05_out;
    52: reg_0366 <= op1_05_out;
    53: reg_0366 <= op1_05_out;
    54: reg_0366 <= op1_05_out;
    55: reg_0366 <= op1_05_out;
    56: reg_0366 <= op1_05_out;
    57: reg_0366 <= op1_05_out;
    58: reg_0366 <= op1_05_out;
    59: reg_0366 <= op1_05_out;
    60: reg_0366 <= op1_05_out;
    61: reg_0366 <= op1_05_out;
    62: reg_0366 <= op1_05_out;
    63: reg_0366 <= op1_05_out;
    64: reg_0366 <= op1_05_out;
    65: reg_0366 <= op1_05_out;
    66: reg_0366 <= op1_05_out;
    67: reg_0366 <= op1_05_out;
    68: reg_0366 <= op1_05_out;
    69: reg_0366 <= op1_05_out;
    70: reg_0366 <= op1_05_out;
    71: reg_0366 <= op1_05_out;
    72: reg_0366 <= op1_05_out;
    73: reg_0366 <= op1_05_out;
    74: reg_0366 <= op1_05_out;
    75: reg_0366 <= op1_05_out;
    76: reg_0366 <= op1_05_out;
    77: reg_0366 <= op1_05_out;
    78: reg_0366 <= op1_05_out;
    79: reg_0366 <= op1_05_out;
    80: reg_0366 <= op1_05_out;
    81: reg_0366 <= op1_05_out;
    82: reg_0366 <= op1_05_out;
    83: reg_0366 <= op1_05_out;
    84: reg_0366 <= op1_05_out;
    85: reg_0366 <= op1_05_out;
    86: reg_0366 <= op1_05_out;
    87: reg_0366 <= op1_05_out;
    88: reg_0366 <= op1_05_out;
    89: reg_0366 <= op1_05_out;
    90: reg_0366 <= op1_05_out;
    91: reg_0366 <= op1_05_out;
    92: reg_0366 <= op1_05_out;
    93: reg_0366 <= op1_05_out;
    94: reg_0366 <= op1_05_out;
    95: reg_0366 <= op1_05_out;
    96: reg_0366 <= op1_05_out;
    endcase
  end

  // REG#367の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0367 <= imem06_in[111:108];
    27: reg_0367 <= imem06_in[123:120];
    29: reg_0367 <= imem03_in[31:28];
    31: reg_0367 <= imem06_in[111:108];
    36: reg_0367 <= imem06_in[111:108];
    60: reg_0367 <= imem06_in[111:108];
    70: reg_0367 <= imem06_in[111:108];
    87: reg_0367 <= imem03_in[31:28];
    endcase
  end

  // REG#368の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0368 <= imem06_in[127:124];
    27: reg_0368 <= imem06_in[71:68];
    29: reg_0368 <= imem03_in[55:52];
    31: reg_0368 <= imem06_in[71:68];
    36: reg_0368 <= imem06_in[71:68];
    60: reg_0368 <= imem06_in[71:68];
    69: reg_0368 <= imem03_in[55:52];
    89: reg_0368 <= imem03_in[55:52];
    endcase
  end

  // REG#369の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0369 <= imem03_in[63:60];
    26: reg_0369 <= imem03_in[63:60];
    28: reg_0369 <= imem06_in[23:20];
    55: reg_0369 <= imem06_in[23:20];
    57: reg_0369 <= imem06_in[23:20];
    84: reg_0369 <= imem06_in[23:20];
    86: reg_0369 <= imem05_in[111:108];
    endcase
  end

  // REG#370の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0370 <= imem03_in[31:28];
    26: reg_0370 <= imem03_in[31:28];
    28: reg_0370 <= imem06_in[39:36];
    56: reg_0370 <= imem06_in[59:56];
    endcase
  end

  // REG#371の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0371 <= imem06_in[67:64];
    27: reg_0371 <= imem06_in[67:64];
    29: reg_0371 <= imem03_in[23:20];
    31: reg_0371 <= imem06_in[67:64];
    35: reg_0371 <= imem06_in[67:64];
    38: reg_0371 <= imem06_in[67:64];
    55: reg_0371 <= imem06_in[67:64];
    58: reg_0371 <= imem04_in[75:72];
    endcase
  end

  // REG#372の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0372 <= imem06_in[31:28];
    27: reg_0372 <= imem06_in[31:28];
    29: reg_0372 <= imem03_in[59:56];
    31: reg_0372 <= imem06_in[31:28];
    36: reg_0372 <= imem06_in[31:28];
    59: reg_0372 <= imem06_in[31:28];
    62: reg_0372 <= imem02_in[111:108];
    69: reg_0372 <= imem03_in[59:56];
    endcase
  end

  // REG#373の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0373 <= imem03_in[55:52];
    27: reg_0373 <= imem03_in[55:52];
    68: reg_0373 <= op2_02_out;
    87: reg_0373 <= op2_02_out;
    endcase
  end

  // REG#374の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0374 <= imem03_in[119:116];
    27: reg_0374 <= imem03_in[119:116];
    67: reg_0374 <= imem05_in[95:92];
    71: reg_0374 <= imem02_in[107:104];
    83: reg_0374 <= imem02_in[107:104];
    endcase
  end

  // REG#375の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0375 <= imem06_in[75:72];
    27: reg_0375 <= imem06_in[87:84];
    29: reg_0375 <= imem03_in[111:108];
    31: reg_0375 <= imem06_in[75:72];
    36: reg_0375 <= imem06_in[75:72];
    55: reg_0375 <= imem06_in[75:72];
    57: reg_0375 <= imem06_in[87:84];
    84: reg_0375 <= imem06_in[75:72];
    86: reg_0375 <= imem03_in[111:108];
    88: reg_0375 <= imem03_in[111:108];
    endcase
  end

  // REG#376の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0376 <= imem03_in[91:88];
    27: reg_0376 <= imem03_in[91:88];
    68: reg_0376 <= imem01_in[3:0];
    92: reg_0376 <= imem01_in[3:0];
    endcase
  end

  // REG#377の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0377 <= imem03_in[75:72];
    26: reg_0377 <= imem03_in[75:72];
    28: reg_0377 <= imem06_in[51:48];
    55: reg_0377 <= imem06_in[51:48];
    57: reg_0377 <= imem06_in[51:48];
    84: reg_0377 <= imem06_in[51:48];
    86: reg_0377 <= imem03_in[75:72];
    88: reg_0377 <= imem03_in[75:72];
    endcase
  end

  // REG#378の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0378 <= op1_06_out;
    25: reg_0378 <= op1_06_out;
    26: reg_0378 <= op1_06_out;
    27: reg_0378 <= op1_06_out;
    28: reg_0378 <= op1_06_out;
    29: reg_0378 <= op1_06_out;
    30: reg_0378 <= op1_06_out;
    31: reg_0378 <= op1_06_out;
    32: reg_0378 <= op1_06_out;
    33: reg_0378 <= op1_06_out;
    34: reg_0378 <= op1_06_out;
    35: reg_0378 <= op1_06_out;
    36: reg_0378 <= op1_06_out;
    37: reg_0378 <= op1_06_out;
    38: reg_0378 <= op1_06_out;
    39: reg_0378 <= op1_06_out;
    40: reg_0378 <= op1_06_out;
    41: reg_0378 <= op1_06_out;
    42: reg_0378 <= op1_06_out;
    43: reg_0378 <= op1_06_out;
    44: reg_0378 <= op1_06_out;
    45: reg_0378 <= op1_06_out;
    46: reg_0378 <= op1_06_out;
    47: reg_0378 <= op1_06_out;
    48: reg_0378 <= op1_06_out;
    49: reg_0378 <= op1_06_out;
    50: reg_0378 <= op1_06_out;
    51: reg_0378 <= op1_06_out;
    52: reg_0378 <= op1_06_out;
    53: reg_0378 <= op1_06_out;
    54: reg_0378 <= op1_06_out;
    55: reg_0378 <= op1_06_out;
    56: reg_0378 <= op1_06_out;
    57: reg_0378 <= op1_06_out;
    58: reg_0378 <= op1_06_out;
    59: reg_0378 <= op1_06_out;
    60: reg_0378 <= op1_06_out;
    61: reg_0378 <= op1_06_out;
    62: reg_0378 <= op1_06_out;
    63: reg_0378 <= op1_06_out;
    64: reg_0378 <= op1_06_out;
    65: reg_0378 <= op1_06_out;
    66: reg_0378 <= op1_06_out;
    67: reg_0378 <= op1_06_out;
    68: reg_0378 <= op1_06_out;
    69: reg_0378 <= op1_06_out;
    70: reg_0378 <= op1_06_out;
    71: reg_0378 <= op1_06_out;
    72: reg_0378 <= op1_06_out;
    73: reg_0378 <= op1_06_out;
    74: reg_0378 <= op1_06_out;
    75: reg_0378 <= op1_06_out;
    76: reg_0378 <= op1_06_out;
    77: reg_0378 <= op1_06_out;
    78: reg_0378 <= op1_06_out;
    79: reg_0378 <= op1_06_out;
    80: reg_0378 <= op1_06_out;
    81: reg_0378 <= op1_06_out;
    82: reg_0378 <= op1_06_out;
    83: reg_0378 <= op1_06_out;
    84: reg_0378 <= op1_06_out;
    85: reg_0378 <= op1_06_out;
    86: reg_0378 <= op1_06_out;
    87: reg_0378 <= op1_06_out;
    88: reg_0378 <= op1_06_out;
    89: reg_0378 <= op1_06_out;
    90: reg_0378 <= op1_06_out;
    91: reg_0378 <= op1_06_out;
    92: reg_0378 <= op1_06_out;
    93: reg_0378 <= op1_06_out;
    94: reg_0378 <= op1_06_out;
    95: reg_0378 <= op1_06_out;
    96: reg_0378 <= op1_06_out;
    endcase
  end

  // REG#379の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0379 <= imem06_in[15:12];
    26: reg_0379 <= op2_01_out;
    35: reg_0379 <= op2_01_out;
    65: reg_0379 <= op2_01_out;
    77: reg_0379 <= op2_01_out;
    endcase
  end

  // REG#380の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0380 <= imem06_in[115:112];
    27: reg_0380 <= imem06_in[115:112];
    29: reg_0380 <= imem03_in[7:4];
    31: reg_0380 <= imem06_in[115:112];
    35: reg_0380 <= imem06_in[115:112];
    37: reg_0380 <= op2_00_out;
    70: reg_0380 <= op2_00_out;
    endcase
  end

  // REG#381の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0381 <= imem06_in[27:24];
    27: reg_0381 <= imem06_in[27:24];
    29: reg_0381 <= imem03_in[103:100];
    31: reg_0381 <= imem06_in[27:24];
    34: reg_0381 <= op2_02_out;
    63: reg_0381 <= op2_02_out;
    72: reg_0381 <= op2_02_out;
    endcase
  end

  // REG#382の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0382 <= imem06_in[79:76];
    26: reg_0382 <= op2_03_out;
    37: reg_0382 <= op2_03_out;
    74: reg_0382 <= imem07_in[63:60];
    78: reg_0382 <= imem07_in[63:60];
    endcase
  end

  // REG#383の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0383 <= imem06_in[83:80];
    27: reg_0383 <= imem03_in[51:48];
    65: reg_0383 <= imem05_in[111:108];
    78: reg_0383 <= imem05_in[111:108];
    85: reg_0383 <= imem05_in[111:108];
    87: reg_0383 <= imem03_in[51:48];
    endcase
  end

  // REG#384の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0384 <= imem03_in[11:8];
    27: reg_0384 <= imem03_in[11:8];
    69: reg_0384 <= imem03_in[11:8];
    endcase
  end

  // REG#385の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0385 <= imem03_in[67:64];
    27: reg_0385 <= imem03_in[67:64];
    68: reg_0385 <= imem01_in[47:44];
    endcase
  end

  // REG#386の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0386 <= imem06_in[59:56];
    27: reg_0386 <= imem03_in[115:112];
    65: reg_0386 <= imem05_in[3:0];
    78: reg_0386 <= imem05_in[3:0];
    84: reg_0386 <= imem06_in[59:56];
    86: reg_0386 <= imem05_in[3:0];
    endcase
  end

  // REG#387の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0387 <= imem03_in[15:12];
    27: reg_0387 <= imem03_in[15:12];
    69: reg_0387 <= imem03_in[99:96];
    endcase
  end

  // REG#388の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0388 <= imem03_in[47:44];
    27: reg_0388 <= imem03_in[47:44];
    68: reg_0388 <= imem01_in[95:92];
    92: reg_0388 <= imem01_in[95:92];
    endcase
  end

  // REG#389の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0389 <= imem03_in[123:120];
    27: reg_0389 <= imem03_in[123:120];
    67: reg_0389 <= imem05_in[115:112];
    71: reg_0389 <= imem05_in[115:112];
    74: reg_0389 <= imem07_in[87:84];
    78: reg_0389 <= imem05_in[115:112];
    85: reg_0389 <= imem05_in[115:112];
    87: reg_0389 <= imem03_in[123:120];
    endcase
  end

  // REG#390の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0390 <= imem06_in[103:100];
    27: reg_0390 <= imem06_in[103:100];
    28: reg_0390 <= op2_00_out;
    41: reg_0390 <= op2_00_out;
    42: reg_0390 <= op2_00_out;
    45: reg_0390 <= op2_00_out;
    55: reg_0390 <= op2_00_out;
    87: reg_0390 <= imem06_in[127:124];
    88: reg_0390 <= op2_00_out;
    endcase
  end

  // REG#391の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0391 <= imem03_in[19:16];
    27: reg_0391 <= imem03_in[19:16];
    67: reg_0391 <= imem05_in[35:32];
    71: reg_0391 <= imem05_in[35:32];
    73: reg_0391 <= imem07_in[23:20];
    78: reg_0391 <= imem07_in[23:20];
    endcase
  end

  // REG#392の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0392 <= imem06_in[43:40];
    27: reg_0392 <= imem03_in[71:68];
    67: reg_0392 <= imem05_in[59:56];
    71: reg_0392 <= imem02_in[35:32];
    83: reg_0392 <= imem02_in[35:32];
    endcase
  end

  // REG#393の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0393 <= imem03_in[103:100];
    27: reg_0393 <= imem03_in[103:100];
    67: reg_0393 <= imem05_in[99:96];
    71: reg_0393 <= imem05_in[99:96];
    74: reg_0393 <= imem07_in[119:116];
    78: reg_0393 <= imem05_in[99:96];
    86: reg_0393 <= imem05_in[99:96];
    endcase
  end

  // REG#394の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0394 <= imem03_in[3:0];
    27: reg_0394 <= imem03_in[3:0];
    68: reg_0394 <= imem01_in[75:72];
    endcase
  end

  // REG#395の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0395 <= imem03_in[7:4];
    27: reg_0395 <= imem03_in[7:4];
    69: reg_0395 <= imem03_in[7:4];
    endcase
  end

  // REG#396の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0396 <= imem03_in[111:108];
    27: reg_0396 <= imem03_in[111:108];
    69: reg_0396 <= imem03_in[111:108];
    endcase
  end

  // REG#397の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0397 <= imem03_in[99:96];
    27: reg_0397 <= imem03_in[99:96];
    68: reg_0397 <= imem01_in[103:100];
    endcase
  end

  // REG#398の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0398 <= imem03_in[87:84];
    27: reg_0398 <= imem03_in[87:84];
    69: reg_0398 <= imem03_in[87:84];
    endcase
  end

  // REG#399の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0399 <= imem06_in[91:88];
    27: reg_0399 <= imem06_in[91:88];
    29: reg_0399 <= op2_03_out;
    48: reg_0399 <= imem04_in[59:56];
    54: reg_0399 <= imem03_in[99:96];
    86: reg_0399 <= imem05_in[79:76];
    92: reg_0399 <= op2_03_out;
    endcase
  end

  // REG#400の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0400 <= op1_07_out;
    26: reg_0400 <= op1_07_out;
    27: reg_0400 <= op1_07_out;
    28: reg_0400 <= op1_07_out;
    29: reg_0400 <= op1_07_out;
    30: reg_0400 <= op1_07_out;
    31: reg_0400 <= op1_07_out;
    32: reg_0400 <= op1_07_out;
    33: reg_0400 <= op1_07_out;
    34: reg_0400 <= op1_07_out;
    35: reg_0400 <= op1_07_out;
    36: reg_0400 <= op1_07_out;
    37: reg_0400 <= op1_07_out;
    38: reg_0400 <= op1_07_out;
    39: reg_0400 <= op1_07_out;
    40: reg_0400 <= op1_07_out;
    41: reg_0400 <= op1_07_out;
    42: reg_0400 <= op1_07_out;
    43: reg_0400 <= op1_07_out;
    44: reg_0400 <= op1_07_out;
    45: reg_0400 <= op1_07_out;
    46: reg_0400 <= op1_07_out;
    47: reg_0400 <= op1_07_out;
    48: reg_0400 <= op1_07_out;
    49: reg_0400 <= op1_07_out;
    50: reg_0400 <= op1_07_out;
    51: reg_0400 <= op1_07_out;
    52: reg_0400 <= op1_07_out;
    53: reg_0400 <= op1_07_out;
    54: reg_0400 <= op1_07_out;
    55: reg_0400 <= op1_07_out;
    56: reg_0400 <= op1_07_out;
    57: reg_0400 <= op1_07_out;
    58: reg_0400 <= op1_07_out;
    59: reg_0400 <= op1_07_out;
    60: reg_0400 <= op1_07_out;
    61: reg_0400 <= op1_07_out;
    62: reg_0400 <= op1_07_out;
    63: reg_0400 <= op1_07_out;
    64: reg_0400 <= op1_07_out;
    65: reg_0400 <= op1_07_out;
    66: reg_0400 <= op1_07_out;
    67: reg_0400 <= op1_07_out;
    68: reg_0400 <= op1_07_out;
    69: reg_0400 <= op1_07_out;
    70: reg_0400 <= op1_07_out;
    71: reg_0400 <= op1_07_out;
    72: reg_0400 <= op1_07_out;
    73: reg_0400 <= op1_07_out;
    74: reg_0400 <= op1_07_out;
    75: reg_0400 <= op1_07_out;
    76: reg_0400 <= op1_07_out;
    77: reg_0400 <= op1_07_out;
    78: reg_0400 <= op1_07_out;
    79: reg_0400 <= op1_07_out;
    80: reg_0400 <= op1_07_out;
    81: reg_0400 <= op1_07_out;
    82: reg_0400 <= op1_07_out;
    83: reg_0400 <= op1_07_out;
    84: reg_0400 <= op1_07_out;
    85: reg_0400 <= op1_07_out;
    86: reg_0400 <= op1_07_out;
    87: reg_0400 <= op1_07_out;
    88: reg_0400 <= op1_07_out;
    89: reg_0400 <= op1_07_out;
    90: reg_0400 <= op1_07_out;
    91: reg_0400 <= op1_07_out;
    92: reg_0400 <= op1_07_out;
    93: reg_0400 <= op1_07_out;
    94: reg_0400 <= op1_07_out;
    95: reg_0400 <= op1_07_out;
    96: reg_0400 <= op1_07_out;
    endcase
  end

  // REG#401の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0401 <= imem06_in[123:120];
    28: reg_0401 <= imem06_in[123:120];
    52: reg_0401 <= imem03_in[119:116];
    56: reg_0401 <= imem06_in[123:120];
    endcase
  end

  // REG#402の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0402 <= imem06_in[3:0];
    28: reg_0402 <= imem06_in[3:0];
    52: reg_0402 <= imem03_in[11:8];
    55: reg_0402 <= imem06_in[3:0];
    57: reg_0402 <= imem06_in[3:0];
    85: reg_0402 <= imem06_in[3:0];
    endcase
  end

  // REG#403の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0403 <= imem06_in[87:84];
    28: reg_0403 <= imem06_in[87:84];
    57: reg_0403 <= imem04_in[127:124];
    59: reg_0403 <= imem05_in[115:112];
    62: reg_0403 <= imem02_in[15:12];
    69: reg_0403 <= imem03_in[67:64];
    endcase
  end

  // REG#404の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0404 <= imem06_in[95:92];
    28: reg_0404 <= imem06_in[95:92];
    56: reg_0404 <= imem06_in[95:92];
    endcase
  end

  // REG#405の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0405 <= imem06_in[55:52];
    28: reg_0405 <= imem06_in[55:52];
    55: reg_0405 <= imem06_in[55:52];
    57: reg_0405 <= imem06_in[55:52];
    85: reg_0405 <= imem06_in[55:52];
    endcase
  end

  // REG#406の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0406 <= imem06_in[107:104];
    28: reg_0406 <= imem06_in[107:104];
    51: reg_0406 <= imem02_in[107:104];
    endcase
  end

  // REG#407の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0407 <= imem06_in[47:44];
    28: reg_0407 <= imem06_in[47:44];
    54: reg_0407 <= imem00_in[95:92];
    86: reg_0407 <= imem05_in[91:88];
    endcase
  end

  // REG#408の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0408 <= imem06_in[35:32];
    28: reg_0408 <= imem06_in[35:32];
    57: reg_0408 <= imem06_in[35:32];
    85: reg_0408 <= imem06_in[35:32];
    endcase
  end

  // REG#409の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0409 <= imem06_in[63:60];
    28: reg_0409 <= imem06_in[63:60];
    56: reg_0409 <= imem06_in[63:60];
    endcase
  end

  // REG#410の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0410 <= op1_08_out;
    28: reg_0410 <= op1_08_out;
    29: reg_0410 <= op1_08_out;
    30: reg_0410 <= op1_08_out;
    31: reg_0410 <= op1_08_out;
    32: reg_0410 <= op1_08_out;
    33: reg_0410 <= op1_08_out;
    34: reg_0410 <= op1_08_out;
    35: reg_0410 <= op1_08_out;
    36: reg_0410 <= op1_08_out;
    37: reg_0410 <= op1_08_out;
    38: reg_0410 <= op1_08_out;
    39: reg_0410 <= op1_08_out;
    40: reg_0410 <= op1_08_out;
    41: reg_0410 <= op1_08_out;
    42: reg_0410 <= op1_08_out;
    43: reg_0410 <= op1_08_out;
    44: reg_0410 <= op1_08_out;
    45: reg_0410 <= op1_08_out;
    46: reg_0410 <= op1_08_out;
    47: reg_0410 <= op1_08_out;
    48: reg_0410 <= op1_08_out;
    49: reg_0410 <= op1_08_out;
    50: reg_0410 <= op1_08_out;
    51: reg_0410 <= op1_08_out;
    52: reg_0410 <= op1_08_out;
    53: reg_0410 <= op1_08_out;
    54: reg_0410 <= op1_08_out;
    55: reg_0410 <= op1_08_out;
    56: reg_0410 <= op1_08_out;
    57: reg_0410 <= op1_08_out;
    58: reg_0410 <= op1_08_out;
    59: reg_0410 <= op1_08_out;
    60: reg_0410 <= op1_08_out;
    61: reg_0410 <= op1_08_out;
    62: reg_0410 <= op1_08_out;
    63: reg_0410 <= op1_08_out;
    64: reg_0410 <= op1_08_out;
    65: reg_0410 <= op1_08_out;
    66: reg_0410 <= op1_08_out;
    67: reg_0410 <= op1_08_out;
    68: reg_0410 <= op1_08_out;
    69: reg_0410 <= op1_08_out;
    70: reg_0410 <= op1_08_out;
    71: reg_0410 <= op1_08_out;
    72: reg_0410 <= op1_08_out;
    73: reg_0410 <= op1_08_out;
    74: reg_0410 <= op1_08_out;
    75: reg_0410 <= op1_08_out;
    76: reg_0410 <= op1_08_out;
    77: reg_0410 <= op1_08_out;
    78: reg_0410 <= op1_08_out;
    79: reg_0410 <= op1_08_out;
    80: reg_0410 <= op1_08_out;
    81: reg_0410 <= op1_08_out;
    82: reg_0410 <= op1_08_out;
    83: reg_0410 <= op1_08_out;
    84: reg_0410 <= op1_08_out;
    85: reg_0410 <= op1_08_out;
    86: reg_0410 <= op1_08_out;
    87: reg_0410 <= op1_08_out;
    88: reg_0410 <= op1_08_out;
    89: reg_0410 <= op1_08_out;
    90: reg_0410 <= op1_08_out;
    91: reg_0410 <= op1_08_out;
    92: reg_0410 <= op1_08_out;
    93: reg_0410 <= op1_08_out;
    94: reg_0410 <= op1_08_out;
    95: reg_0410 <= op1_08_out;
    96: reg_0410 <= op1_08_out;
    endcase
  end

  // REG#411の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0411 <= op1_09_out;
    29: reg_0411 <= op1_09_out;
    30: reg_0411 <= op1_09_out;
    31: reg_0411 <= op1_09_out;
    32: reg_0411 <= op1_09_out;
    33: reg_0411 <= op1_09_out;
    34: reg_0411 <= op1_09_out;
    35: reg_0411 <= op1_09_out;
    36: reg_0411 <= op1_09_out;
    37: reg_0411 <= op1_09_out;
    38: reg_0411 <= op1_09_out;
    39: reg_0411 <= op1_09_out;
    40: reg_0411 <= op1_09_out;
    41: reg_0411 <= op1_09_out;
    42: reg_0411 <= op1_09_out;
    43: reg_0411 <= op1_09_out;
    44: reg_0411 <= op1_09_out;
    45: reg_0411 <= op1_09_out;
    46: reg_0411 <= op1_09_out;
    47: reg_0411 <= op1_09_out;
    48: reg_0411 <= op1_09_out;
    49: reg_0411 <= op1_09_out;
    50: reg_0411 <= op1_09_out;
    51: reg_0411 <= op1_09_out;
    52: reg_0411 <= op1_09_out;
    53: reg_0411 <= op1_09_out;
    54: reg_0411 <= op1_09_out;
    55: reg_0411 <= op1_09_out;
    56: reg_0411 <= op1_09_out;
    57: reg_0411 <= op1_09_out;
    58: reg_0411 <= op1_09_out;
    59: reg_0411 <= op1_09_out;
    60: reg_0411 <= op1_09_out;
    61: reg_0411 <= op1_09_out;
    62: reg_0411 <= op1_09_out;
    63: reg_0411 <= op1_09_out;
    64: reg_0411 <= op1_09_out;
    65: reg_0411 <= op1_09_out;
    66: reg_0411 <= op1_09_out;
    67: reg_0411 <= op1_09_out;
    68: reg_0411 <= op1_09_out;
    69: reg_0411 <= op1_09_out;
    70: reg_0411 <= op1_09_out;
    71: reg_0411 <= op1_09_out;
    72: reg_0411 <= op1_09_out;
    73: reg_0411 <= op1_09_out;
    74: reg_0411 <= op1_09_out;
    75: reg_0411 <= op1_09_out;
    76: reg_0411 <= op1_09_out;
    77: reg_0411 <= op1_09_out;
    78: reg_0411 <= op1_09_out;
    79: reg_0411 <= op1_09_out;
    80: reg_0411 <= op1_09_out;
    81: reg_0411 <= op1_09_out;
    82: reg_0411 <= op1_09_out;
    83: reg_0411 <= op1_09_out;
    84: reg_0411 <= op1_09_out;
    85: reg_0411 <= op1_09_out;
    86: reg_0411 <= op1_09_out;
    87: reg_0411 <= op1_09_out;
    88: reg_0411 <= op1_09_out;
    89: reg_0411 <= op1_09_out;
    90: reg_0411 <= op1_09_out;
    91: reg_0411 <= op1_09_out;
    92: reg_0411 <= op1_09_out;
    93: reg_0411 <= op1_09_out;
    94: reg_0411 <= op1_09_out;
    95: reg_0411 <= op1_09_out;
    96: reg_0411 <= op1_09_out;
    endcase
  end

  // REG#412の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0412 <= op1_10_out;
    31: reg_0412 <= op1_10_out;
    32: reg_0412 <= op1_10_out;
    33: reg_0412 <= op1_10_out;
    34: reg_0412 <= op1_10_out;
    35: reg_0412 <= op1_10_out;
    36: reg_0412 <= op1_10_out;
    37: reg_0412 <= op1_10_out;
    38: reg_0412 <= op1_10_out;
    39: reg_0412 <= op1_10_out;
    40: reg_0412 <= op1_10_out;
    41: reg_0412 <= op1_10_out;
    42: reg_0412 <= op1_10_out;
    43: reg_0412 <= op1_10_out;
    44: reg_0412 <= op1_10_out;
    45: reg_0412 <= op1_10_out;
    46: reg_0412 <= op1_10_out;
    47: reg_0412 <= op1_10_out;
    48: reg_0412 <= op1_10_out;
    49: reg_0412 <= op1_10_out;
    50: reg_0412 <= op1_10_out;
    51: reg_0412 <= op1_10_out;
    52: reg_0412 <= op1_10_out;
    53: reg_0412 <= op1_10_out;
    54: reg_0412 <= op1_10_out;
    55: reg_0412 <= op1_10_out;
    56: reg_0412 <= op1_10_out;
    57: reg_0412 <= op1_10_out;
    58: reg_0412 <= op1_10_out;
    59: reg_0412 <= op1_10_out;
    60: reg_0412 <= op1_10_out;
    61: reg_0412 <= op1_10_out;
    62: reg_0412 <= op1_10_out;
    63: reg_0412 <= op1_10_out;
    64: reg_0412 <= op1_10_out;
    65: reg_0412 <= op1_10_out;
    66: reg_0412 <= op1_10_out;
    67: reg_0412 <= op1_10_out;
    68: reg_0412 <= op1_10_out;
    69: reg_0412 <= op1_10_out;
    70: reg_0412 <= op1_10_out;
    71: reg_0412 <= op1_10_out;
    72: reg_0412 <= op1_10_out;
    73: reg_0412 <= op1_10_out;
    74: reg_0412 <= op1_10_out;
    75: reg_0412 <= op1_10_out;
    76: reg_0412 <= op1_10_out;
    77: reg_0412 <= op1_10_out;
    78: reg_0412 <= op1_10_out;
    79: reg_0412 <= op1_10_out;
    80: reg_0412 <= op1_10_out;
    81: reg_0412 <= op1_10_out;
    82: reg_0412 <= op1_10_out;
    83: reg_0412 <= op1_10_out;
    84: reg_0412 <= op1_10_out;
    85: reg_0412 <= op1_10_out;
    86: reg_0412 <= op1_10_out;
    87: reg_0412 <= op1_10_out;
    88: reg_0412 <= op1_10_out;
    89: reg_0412 <= op1_10_out;
    90: reg_0412 <= op1_10_out;
    91: reg_0412 <= op1_10_out;
    92: reg_0412 <= op1_10_out;
    93: reg_0412 <= op1_10_out;
    94: reg_0412 <= op1_10_out;
    95: reg_0412 <= op1_10_out;
    96: reg_0412 <= op1_10_out;
    endcase
  end

  // REG#413の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0413 <= op1_11_out;
    32: reg_0413 <= op1_11_out;
    33: reg_0413 <= op1_11_out;
    34: reg_0413 <= op1_11_out;
    35: reg_0413 <= op1_11_out;
    36: reg_0413 <= op1_11_out;
    37: reg_0413 <= op1_11_out;
    38: reg_0413 <= op1_11_out;
    39: reg_0413 <= op1_11_out;
    40: reg_0413 <= op1_11_out;
    41: reg_0413 <= op1_11_out;
    42: reg_0413 <= op1_11_out;
    43: reg_0413 <= op1_11_out;
    44: reg_0413 <= op1_11_out;
    45: reg_0413 <= op1_11_out;
    46: reg_0413 <= op1_11_out;
    47: reg_0413 <= op1_11_out;
    48: reg_0413 <= op1_11_out;
    49: reg_0413 <= op1_11_out;
    50: reg_0413 <= op1_11_out;
    51: reg_0413 <= op1_11_out;
    52: reg_0413 <= op1_11_out;
    53: reg_0413 <= op1_11_out;
    54: reg_0413 <= op1_11_out;
    55: reg_0413 <= op1_11_out;
    56: reg_0413 <= op1_11_out;
    57: reg_0413 <= op1_11_out;
    58: reg_0413 <= op1_11_out;
    59: reg_0413 <= op1_11_out;
    60: reg_0413 <= op1_11_out;
    61: reg_0413 <= op1_11_out;
    62: reg_0413 <= op1_11_out;
    63: reg_0413 <= op1_11_out;
    64: reg_0413 <= op1_11_out;
    65: reg_0413 <= op1_11_out;
    66: reg_0413 <= op1_11_out;
    67: reg_0413 <= op1_11_out;
    68: reg_0413 <= op1_11_out;
    69: reg_0413 <= op1_11_out;
    70: reg_0413 <= op1_11_out;
    71: reg_0413 <= op1_11_out;
    72: reg_0413 <= op1_11_out;
    73: reg_0413 <= op1_11_out;
    74: reg_0413 <= op1_11_out;
    75: reg_0413 <= op1_11_out;
    76: reg_0413 <= op1_11_out;
    77: reg_0413 <= op1_11_out;
    78: reg_0413 <= op1_11_out;
    79: reg_0413 <= op1_11_out;
    80: reg_0413 <= op1_11_out;
    82: reg_0413 <= op1_11_out;
    83: reg_0413 <= op1_11_out;
    84: reg_0413 <= op1_11_out;
    85: reg_0413 <= op1_11_out;
    87: reg_0413 <= op1_11_out;
    88: reg_0413 <= op1_11_out;
    89: reg_0413 <= op1_11_out;
    90: reg_0413 <= op1_11_out;
    91: reg_0413 <= op1_11_out;
    92: reg_0413 <= op1_11_out;
    93: reg_0413 <= op1_11_out;
    94: reg_0413 <= op1_11_out;
    95: reg_0413 <= op1_11_out;
    endcase
  end

  // REG#414の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0414 <= op1_12_out;
    33: reg_0414 <= op1_12_out;
    34: reg_0414 <= op1_12_out;
    36: reg_0414 <= op1_12_out;
    37: reg_0414 <= op1_12_out;
    38: reg_0414 <= op1_12_out;
    39: reg_0414 <= op1_12_out;
    40: reg_0414 <= op1_12_out;
    41: reg_0414 <= op1_12_out;
    43: reg_0414 <= op1_12_out;
    44: reg_0414 <= op1_12_out;
    45: reg_0414 <= op1_12_out;
    46: reg_0414 <= op1_12_out;
    47: reg_0414 <= op1_12_out;
    48: reg_0414 <= op1_12_out;
    51: reg_0414 <= imem02_in[99:96];
    endcase
  end

  // REG#415の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0415 <= op1_13_out;
    33: reg_0415 <= op1_13_out;
    35: reg_0415 <= op1_13_out;
    37: reg_0415 <= op2_02_out;
    72: reg_0415 <= op1_13_out;
    74: reg_0415 <= op1_13_out;
    75: reg_0415 <= op2_02_out;
    endcase
  end

  // REG#416の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0416 <= op1_14_out;
    34: reg_0416 <= imem06_in[43:40];
    36: reg_0416 <= op1_14_out;
    38: reg_0416 <= imem06_in[43:40];
    53: reg_0416 <= op1_14_out;
    55: reg_0416 <= op1_14_out;
    58: reg_0416 <= imem04_in[111:108];
    endcase
  end

  // REG#417の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0417 <= op1_15_out;
    34: reg_0417 <= op1_15_out;
    36: reg_0417 <= op1_15_out;
    39: reg_0417 <= op1_15_out;
    41: reg_0417 <= op1_15_out;
    44: reg_0417 <= imem02_in[87:84];
    60: reg_0417 <= op1_15_out;
    62: reg_0417 <= imem02_in[87:84];
    69: reg_0417 <= imem03_in[31:28];
    endcase
  end

  // REG#418の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0418 <= imem07_in[51:48];
    40: reg_0418 <= imem01_in[23:20];
    89: reg_0418 <= imem03_in[39:36];
    endcase
  end

  // REG#419の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0419 <= imem07_in[55:52];
    40: reg_0419 <= imem01_in[107:104];
    93: reg_0419 <= imem01_in[107:104];
    endcase
  end

  // REG#420の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0420 <= imem07_in[111:108];
    40: reg_0420 <= imem01_in[127:124];
    94: reg_0420 <= imem01_in[127:124];
    endcase
  end

  // REG#421の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0421 <= imem07_in[39:36];
    40: reg_0421 <= imem01_in[19:16];
    91: reg_0421 <= imem01_in[19:16];
    endcase
  end

  // REG#422の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0422 <= imem07_in[31:28];
    40: reg_0422 <= imem01_in[35:32];
    91: reg_0422 <= imem01_in[35:32];
    endcase
  end

  // REG#423の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0423 <= imem07_in[59:56];
    40: reg_0423 <= imem01_in[15:12];
    endcase
  end

  // REG#424の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0424 <= imem07_in[11:8];
    40: reg_0424 <= imem01_in[111:108];
    92: reg_0424 <= imem01_in[111:108];
    94: reg_0424 <= imem01_in[111:108];
    endcase
  end

  // REG#425の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0425 <= imem07_in[3:0];
    40: reg_0425 <= imem01_in[83:80];
    92: reg_0425 <= imem01_in[83:80];
    94: reg_0425 <= imem01_in[83:80];
    endcase
  end

  // REG#426の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0426 <= imem07_in[43:40];
    41: reg_0426 <= imem07_in[63:60];
    44: reg_0426 <= imem02_in[115:112];
    62: reg_0426 <= imem02_in[115:112];
    71: reg_0426 <= imem02_in[115:112];
    81: reg_0426 <= imem07_in[43:40];
    endcase
  end

  // REG#427の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0427 <= imem07_in[103:100];
    41: reg_0427 <= imem07_in[103:100];
    44: reg_0427 <= imem02_in[119:116];
    62: reg_0427 <= imem02_in[119:116];
    71: reg_0427 <= imem02_in[119:116];
    81: reg_0427 <= imem07_in[103:100];
    endcase
  end

  // REG#428の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0428 <= imem07_in[71:68];
    40: reg_0428 <= op2_01_out;
    82: reg_0428 <= op2_01_out;
    91: reg_0428 <= op2_01_out;
    endcase
  end

  // REG#429の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0429 <= imem07_in[19:16];
    41: reg_0429 <= imem04_in[11:8];
    endcase
  end

  // REG#430の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0430 <= imem07_in[15:12];
    41: reg_0430 <= imem04_in[67:64];
    endcase
  end

  // REG#431の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0431 <= imem07_in[127:124];
    41: reg_0431 <= imem04_in[103:100];
    endcase
  end

  // REG#432の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0432 <= imem07_in[23:20];
    41: reg_0432 <= imem04_in[15:12];
    endcase
  end

  // REG#433の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0433 <= imem07_in[35:32];
    41: reg_0433 <= imem04_in[39:36];
    endcase
  end

  // REG#434の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0434 <= imem07_in[75:72];
    42: reg_0434 <= imem07_in[75:72];
    endcase
  end

  // REG#435の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0435 <= imem07_in[123:120];
    42: reg_0435 <= imem07_in[123:120];
    endcase
  end

  // REG#436の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0436 <= imem07_in[27:24];
    42: reg_0436 <= imem07_in[27:24];
    endcase
  end

  // REG#437の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0437 <= imem07_in[107:104];
    42: reg_0437 <= imem07_in[107:104];
    endcase
  end

  // REG#438の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0438 <= imem07_in[115:112];
    42: reg_0438 <= imem07_in[115:112];
    endcase
  end

  // REG#439の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0439 <= imem07_in[67:64];
    42: reg_0439 <= imem07_in[67:64];
    endcase
  end

  // REG#440の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0440 <= imem07_in[87:84];
    42: reg_0440 <= imem07_in[87:84];
    endcase
  end

  // REG#441の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0441 <= imem07_in[7:4];
    42: reg_0441 <= imem07_in[7:4];
    endcase
  end

  // REG#442の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0442 <= imem07_in[95:92];
    42: reg_0442 <= imem07_in[95:92];
    endcase
  end

  // REG#443の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0443 <= imem07_in[99:96];
    42: reg_0443 <= imem07_in[99:96];
    endcase
  end

  // REG#444の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0444 <= imem07_in[91:88];
    42: reg_0444 <= imem07_in[91:88];
    endcase
  end

  // REG#445の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0445 <= imem07_in[63:60];
    42: reg_0445 <= imem07_in[63:60];
    endcase
  end

  // REG#446の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0446 <= imem07_in[79:76];
    42: reg_0446 <= imem07_in[79:76];
    endcase
  end

  // REG#447の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0447 <= imem07_in[47:44];
    42: reg_0447 <= imem07_in[47:44];
    endcase
  end

  // REG#448の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0448 <= imem07_in[119:116];
    42: reg_0448 <= imem07_in[119:116];
    endcase
  end

  // REG#449の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0449 <= imem07_in[83:80];
    42: reg_0449 <= imem07_in[83:80];
    endcase
  end

  // REG#450の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0450 <= imem00_in[19:16];
    endcase
  end

  // REG#451の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0451 <= imem00_in[23:20];
    endcase
  end

  // REG#452の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0452 <= imem00_in[115:112];
    endcase
  end

  // REG#453の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0453 <= imem00_in[11:8];
    endcase
  end

  // REG#454の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0454 <= imem00_in[15:12];
    endcase
  end

  // REG#455の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0455 <= imem00_in[27:24];
    endcase
  end

  // REG#456の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0456 <= imem00_in[119:116];
    endcase
  end

  // REG#457の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0457 <= imem00_in[31:28];
    endcase
  end

  // REG#458の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0458 <= imem00_in[127:124];
    endcase
  end

  // REG#459の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0459 <= imem00_in[111:108];
    endcase
  end

  // REG#460の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0460 <= imem00_in[63:60];
    endcase
  end

  // REG#461の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0461 <= imem00_in[39:36];
    endcase
  end

  // REG#462の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0462 <= imem00_in[67:64];
    endcase
  end

  // REG#463の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0463 <= imem00_in[3:0];
    endcase
  end

  // REG#464の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0464 <= imem00_in[35:32];
    endcase
  end

  // REG#465の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0465 <= imem00_in[7:4];
    endcase
  end

  // REG#466の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0466 <= imem00_in[55:52];
    endcase
  end

  // REG#467の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0467 <= imem00_in[87:84];
    endcase
  end

  // REG#468の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0468 <= imem00_in[103:100];
    endcase
  end

  // REG#469の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0469 <= imem00_in[47:44];
    endcase
  end

  // REG#470の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0470 <= imem00_in[91:88];
    endcase
  end

  // REG#471の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0471 <= imem00_in[99:96];
    endcase
  end

  // REG#472の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0472 <= imem00_in[75:72];
    endcase
  end

  // REG#473の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0473 <= imem00_in[83:80];
    endcase
  end

  // REG#474の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0474 <= imem00_in[95:92];
    endcase
  end

  // REG#475の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0475 <= imem00_in[59:56];
    endcase
  end

  // REG#476の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0476 <= imem00_in[51:48];
    endcase
  end

  // REG#477の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0477 <= imem00_in[43:40];
    endcase
  end

  // REG#478の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0478 <= imem00_in[123:120];
    endcase
  end

  // REG#479の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0479 <= imem00_in[107:104];
    endcase
  end

  // REG#480の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0480 <= imem00_in[79:76];
    endcase
  end

  // REG#481の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0481 <= imem00_in[71:68];
    endcase
  end

  // REG#482の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0482 <= imem05_in[19:16];
    5: reg_0482 <= imem05_in[19:16];
    57: reg_0482 <= imem04_in[71:68];
    58: reg_0482 <= op2_01_out;
    endcase
  end

  // REG#483の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0483 <= imem05_in[23:20];
    5: reg_0483 <= imem05_in[23:20];
    57: reg_0483 <= imem04_in[119:116];
    59: reg_0483 <= imem05_in[23:20];
    62: reg_0483 <= imem02_in[59:56];
    69: reg_0483 <= imem03_in[51:48];
    endcase
  end

  // REG#484の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0484 <= imem05_in[43:40];
    5: reg_0484 <= imem05_in[43:40];
    57: reg_0484 <= imem04_in[3:0];
    59: reg_0484 <= imem05_in[43:40];
    62: reg_0484 <= imem02_in[83:80];
    70: reg_0484 <= imem06_in[71:68];
    85: reg_0484 <= imem06_in[71:68];
    endcase
  end

  // REG#485の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0485 <= imem05_in[115:112];
    5: reg_0485 <= imem05_in[115:112];
    51: reg_0485 <= imem02_in[7:4];
    endcase
  end

  // REG#486の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0486 <= imem05_in[127:124];
    5: reg_0486 <= imem05_in[127:124];
    55: reg_0486 <= imem05_in[127:124];
    60: reg_0486 <= imem05_in[127:124];
    63: reg_0486 <= imem05_in[127:124];
    65: reg_0486 <= imem05_in[127:124];
    78: reg_0486 <= imem05_in[27:24];
    85: reg_0486 <= imem05_in[27:24];
    87: reg_0486 <= imem03_in[119:116];
    endcase
  end

  // REG#487の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0487 <= imem01_in[99:96];
    4: reg_0487 <= op1_04_out;
    5: reg_0487 <= op1_04_out;
    6: reg_0487 <= op1_04_out;
    7: reg_0487 <= op1_04_out;
    8: reg_0487 <= op1_04_out;
    9: reg_0487 <= op1_04_out;
    10: reg_0487 <= op1_04_out;
    11: reg_0487 <= op1_04_out;
    12: reg_0487 <= op1_04_out;
    13: reg_0487 <= op1_04_out;
    14: reg_0487 <= op1_04_out;
    15: reg_0487 <= op1_04_out;
    16: reg_0487 <= op1_04_out;
    17: reg_0487 <= op1_04_out;
    18: reg_0487 <= op1_04_out;
    19: reg_0487 <= op1_04_out;
    20: reg_0487 <= op1_04_out;
    21: reg_0487 <= op1_04_out;
    22: reg_0487 <= op1_04_out;
    24: reg_0487 <= imem01_in[99:96];
    45: reg_0487 <= imem04_in[103:100];
    48: reg_0487 <= imem01_in[99:96];
    67: reg_0487 <= imem05_in[75:72];
    71: reg_0487 <= imem02_in[51:48];
    82: reg_0487 <= imem02_in[51:48];
    84: reg_0487 <= imem02_in[51:48];
    endcase
  end

  // REG#488の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0488 <= imem05_in[39:36];
    5: reg_0488 <= imem05_in[39:36];
    54: reg_0488 <= imem03_in[95:92];
    86: reg_0488 <= imem05_in[39:36];
    endcase
  end

  // REG#489の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0489 <= imem05_in[123:120];
    5: reg_0489 <= imem05_in[123:120];
    57: reg_0489 <= imem04_in[23:20];
    60: reg_0489 <= imem05_in[123:120];
    64: reg_0489 <= imem05_in[123:120];
    67: reg_0489 <= imem05_in[123:120];
    72: reg_0489 <= imem05_in[119:116];
    endcase
  end

  // REG#490の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0490 <= imem05_in[35:32];
    5: reg_0490 <= imem05_in[35:32];
    55: reg_0490 <= imem05_in[35:32];
    60: reg_0490 <= imem05_in[43:40];
    64: reg_0490 <= imem05_in[35:32];
    66: reg_0490 <= imem05_in[43:40];
    69: reg_0490 <= imem03_in[71:68];
    endcase
  end

  // REG#491の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0491 <= imem05_in[55:52];
    5: reg_0491 <= imem05_in[55:52];
    54: reg_0491 <= imem05_in[55:52];
    57: reg_0491 <= imem04_in[95:92];
    60: reg_0491 <= imem05_in[55:52];
    65: reg_0491 <= imem05_in[55:52];
    78: reg_0491 <= imem05_in[55:52];
    86: reg_0491 <= imem05_in[55:52];
    endcase
  end

  // REG#492の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0492 <= imem05_in[59:56];
    5: reg_0492 <= imem05_in[59:56];
    54: reg_0492 <= imem00_in[35:32];
    86: reg_0492 <= imem05_in[59:56];
    endcase
  end

  // REG#493の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0493 <= imem05_in[67:64];
    5: reg_0493 <= imem05_in[67:64];
    54: reg_0493 <= imem03_in[51:48];
    87: reg_0493 <= imem03_in[99:96];
    endcase
  end

  // REG#494の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0494 <= imem05_in[75:72];
    5: reg_0494 <= imem05_in[75:72];
    54: reg_0494 <= imem00_in[99:96];
    87: reg_0494 <= imem03_in[67:64];
    endcase
  end

  // REG#495の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0495 <= imem05_in[87:84];
    5: reg_0495 <= imem05_in[87:84];
    55: reg_0495 <= imem05_in[87:84];
    60: reg_0495 <= imem06_in[107:104];
    65: reg_0495 <= imem05_in[87:84];
    78: reg_0495 <= imem05_in[87:84];
    86: reg_0495 <= imem05_in[87:84];
    endcase
  end

  // REG#496の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0496 <= imem01_in[19:16];
    8: reg_0496 <= imem01_in[47:44];
    10: reg_0496 <= imem01_in[19:16];
    24: reg_0496 <= imem01_in[19:16];
    48: reg_0496 <= imem01_in[47:44];
    60: reg_0496 <= imem06_in[75:72];
    67: reg_0496 <= imem01_in[19:16];
    69: reg_0496 <= imem03_in[91:88];
    endcase
  end

  // REG#497の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0497 <= op1_00_out;
    8: reg_0497 <= imem01_in[15:12];
    10: reg_0497 <= imem01_in[15:12];
    24: reg_0497 <= imem01_in[15:12];
    48: reg_0497 <= imem01_in[15:12];
    68: reg_0497 <= imem01_in[15:12];
    endcase
  end

  // REG#498の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0498 <= imem01_in[115:112];
    8: reg_0498 <= imem01_in[115:112];
    11: reg_0498 <= imem05_in[11:8];
    18: reg_0498 <= imem05_in[11:8];
    20: reg_0498 <= imem02_in[87:84];
    83: reg_0498 <= imem02_in[87:84];
    94: reg_0498 <= imem01_in[115:112];
    endcase
  end

  // REG#499の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0499 <= imem01_in[75:72];
    8: reg_0499 <= imem01_in[27:24];
    10: reg_0499 <= imem01_in[75:72];
    23: reg_0499 <= imem01_in[27:24];
    27: reg_0499 <= imem03_in[95:92];
    67: reg_0499 <= imem05_in[87:84];
    72: reg_0499 <= imem05_in[87:84];
    95: reg_0499 <= imem01_in[27:24];
    endcase
  end

  // REG#500の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0500 <= imem01_in[55:52];
    8: reg_0500 <= imem01_in[55:52];
    10: reg_0500 <= imem01_in[55:52];
    23: reg_0500 <= imem04_in[119:116];
    78: reg_0500 <= imem05_in[43:40];
    86: reg_0500 <= imem05_in[43:40];
    endcase
  end

  // REG#501の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0501 <= imem01_in[11:8];
    7: reg_0501 <= op1_13_out;
    10: reg_0501 <= imem01_in[11:8];
    22: reg_0501 <= op1_13_out;
    24: reg_0501 <= imem01_in[11:8];
    48: reg_0501 <= imem04_in[39:36];
    55: reg_0501 <= op1_13_out;
    57: reg_0501 <= op1_13_out;
    59: reg_0501 <= op1_13_out;
    62: reg_0501 <= imem02_in[3:0];
    70: reg_0501 <= imem06_in[75:72];
    84: reg_0501 <= op1_13_out;
    86: reg_0501 <= op1_13_out;
    88: reg_0501 <= imem06_in[75:72];
    endcase
  end

  // REG#502の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0502 <= imem01_in[59:56];
    9: reg_0502 <= imem01_in[59:56];
    38: reg_0502 <= imem01_in[59:56];
    40: reg_0502 <= imem01_in[59:56];
    endcase
  end

  // REG#503の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0503 <= imem01_in[79:76];
    9: reg_0503 <= imem01_in[79:76];
    38: reg_0503 <= imem01_in[79:76];
    41: reg_0503 <= imem04_in[83:80];
    endcase
  end

  // REG#504の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0504 <= imem01_in[7:4];
    9: reg_0504 <= imem01_in[99:96];
    40: reg_0504 <= imem01_in[99:96];
    94: reg_0504 <= imem01_in[99:96];
    endcase
  end

  // REG#505の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0505 <= imem01_in[123:120];
    9: reg_0505 <= imem01_in[15:12];
    40: reg_0505 <= imem01_in[123:120];
    91: reg_0505 <= imem01_in[123:120];
    endcase
  end

  // REG#506の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0506 <= imem01_in[103:100];
    9: reg_0506 <= imem01_in[39:36];
    40: reg_0506 <= imem01_in[103:100];
    91: reg_0506 <= imem01_in[103:100];
    endcase
  end

  // REG#507の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0507 <= imem01_in[119:116];
    10: reg_0507 <= imem01_in[119:116];
    24: reg_0507 <= imem01_in[119:116];
    48: reg_0507 <= imem04_in[51:48];
    57: reg_0507 <= imem04_in[67:64];
    60: reg_0507 <= imem06_in[63:60];
    68: reg_0507 <= imem01_in[119:116];
    87: reg_0507 <= imem03_in[115:112];
    endcase
  end

  // REG#508の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0508 <= imem01_in[127:124];
    9: reg_0508 <= imem01_in[127:124];
    38: reg_0508 <= imem01_in[127:124];
    41: reg_0508 <= imem04_in[111:108];
    endcase
  end

  // REG#509の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0509 <= imem01_in[43:40];
    10: reg_0509 <= imem01_in[31:28];
    18: reg_0509 <= op2_01_out;
    51: reg_0509 <= imem01_in[43:40];
    54: reg_0509 <= imem03_in[123:120];
    87: reg_0509 <= imem03_in[11:8];
    endcase
  end

  // REG#510の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0510 <= imem01_in[111:108];
    10: reg_0510 <= imem01_in[111:108];
    23: reg_0510 <= imem04_in[111:108];
    82: reg_0510 <= imem04_in[111:108];
    93: reg_0510 <= imem01_in[111:108];
    endcase
  end

  // REG#511の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0511 <= imem01_in[31:28];
    9: reg_0511 <= imem01_in[31:28];
    40: reg_0511 <= imem01_in[31:28];
    92: reg_0511 <= imem01_in[31:28];
    endcase
  end

  // REG#512の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0512 <= imem01_in[27:24];
    10: reg_0512 <= imem01_in[27:24];
    24: reg_0512 <= imem01_in[27:24];
    45: reg_0512 <= imem04_in[7:4];
    48: reg_0512 <= imem04_in[7:4];
    57: reg_0512 <= imem06_in[127:124];
    85: reg_0512 <= imem06_in[127:124];
    endcase
  end

  // REG#513の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0513 <= imem01_in[23:20];
    10: reg_0513 <= imem01_in[23:20];
    24: reg_0513 <= imem01_in[23:20];
    45: reg_0513 <= imem04_in[19:16];
    48: reg_0513 <= imem04_in[19:16];
    58: reg_0513 <= imem04_in[71:68];
    95: reg_0513 <= imem01_in[23:20];
    endcase
  end

  // REG#514の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0514 <= imem01_in[47:44];
    10: reg_0514 <= imem01_in[47:44];
    24: reg_0514 <= imem01_in[47:44];
    46: reg_0514 <= imem01_in[47:44];
    51: reg_0514 <= imem02_in[123:120];
    endcase
  end

  // REG#515の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0515 <= imem01_in[95:92];
    10: reg_0515 <= imem01_in[95:92];
    22: reg_0515 <= imem04_in[55:52];
    24: reg_0515 <= imem01_in[95:92];
    48: reg_0515 <= imem04_in[55:52];
    57: reg_0515 <= imem06_in[123:120];
    85: reg_0515 <= imem06_in[123:120];
    endcase
  end

  // REG#516の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0516 <= imem01_in[107:104];
    10: reg_0516 <= imem01_in[107:104];
    23: reg_0516 <= imem04_in[115:112];
    82: reg_0516 <= imem04_in[115:112];
    endcase
  end

  // REG#517の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0517 <= imem01_in[83:80];
    10: reg_0517 <= imem01_in[83:80];
    23: reg_0517 <= imem01_in[83:80];
    27: reg_0517 <= imem03_in[59:56];
    67: reg_0517 <= imem05_in[127:124];
    72: reg_0517 <= imem05_in[127:124];
    endcase
  end

  // REG#518の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0518 <= imem01_in[91:88];
    10: reg_0518 <= imem01_in[91:88];
    20: reg_0518 <= imem02_in[3:0];
    82: reg_0518 <= imem02_in[3:0];
    86: reg_0518 <= imem05_in[11:8];
    93: reg_0518 <= imem01_in[91:88];
    endcase
  end

  // REG#519の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0519 <= imem01_in[67:64];
    10: reg_0519 <= imem01_in[67:64];
    24: reg_0519 <= imem01_in[67:64];
    45: reg_0519 <= imem04_in[87:84];
    48: reg_0519 <= imem04_in[99:96];
    57: reg_0519 <= imem06_in[19:16];
    85: reg_0519 <= imem06_in[19:16];
    endcase
  end

  // REG#520の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0520 <= imem01_in[35:32];
    10: reg_0520 <= imem01_in[35:32];
    22: reg_0520 <= imem04_in[91:88];
    24: reg_0520 <= imem01_in[35:32];
    45: reg_0520 <= imem04_in[15:12];
    48: reg_0520 <= imem04_in[15:12];
    57: reg_0520 <= imem04_in[15:12];
    60: reg_0520 <= imem06_in[15:12];
    68: reg_0520 <= imem01_in[35:32];
    92: reg_0520 <= imem01_in[35:32];
    94: reg_0520 <= imem01_in[35:32];
    endcase
  end

  // REG#521の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0521 <= imem01_in[71:68];
    10: reg_0521 <= imem01_in[71:68];
    21: reg_0521 <= op2_00_out;
    60: reg_0521 <= op2_00_out;
    61: reg_0521 <= op2_00_out;
    66: reg_0521 <= op2_00_out;
    79: reg_0521 <= op2_00_out;
    82: reg_0521 <= op2_00_out;
    89: reg_0521 <= op2_00_out;
    endcase
  end

  // REG#522の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0522 <= imem01_in[15:12];
    10: reg_0522 <= imem01_in[7:4];
    20: reg_0522 <= op2_00_out;
    56: reg_0522 <= op2_00_out;
    91: reg_0522 <= imem01_in[7:4];
    endcase
  end

  // REG#523の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0523 <= imem01_in[3:0];
    10: reg_0523 <= imem01_in[3:0];
    23: reg_0523 <= imem04_in[95:92];
    82: reg_0523 <= imem04_in[95:92];
    endcase
  end

  // REG#524の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0524 <= imem01_in[63:60];
    9: reg_0524 <= op2_01_out;
    20: reg_0524 <= op2_01_out;
    57: reg_0524 <= op2_01_out;
    endcase
  end

  // REG#525の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0525 <= op1_01_out;
    10: reg_0525 <= imem01_in[103:100];
    21: reg_0525 <= op2_01_out;
    61: reg_0525 <= op2_01_out;
    66: reg_0525 <= op2_01_out;
    80: reg_0525 <= op2_01_out;
    84: reg_0525 <= op1_01_out;
    85: reg_0525 <= op2_01_out;
    endcase
  end

  // REG#526の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0526 <= op1_02_out;
    11: reg_0526 <= imem05_in[67:64];
    18: reg_0526 <= imem05_in[67:64];
    20: reg_0526 <= imem02_in[95:92];
    84: reg_0526 <= imem02_in[95:92];
    endcase
  end

  // REG#527の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0527 <= op1_03_out;
    11: reg_0527 <= imem05_in[51:48];
    19: reg_0527 <= imem05_in[51:48];
    48: reg_0527 <= imem05_in[51:48];
    51: reg_0527 <= imem02_in[103:100];
    endcase
  end

  // REG#528の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0528 <= imem04_in[43:40];
    18: reg_0528 <= op2_03_out;
    54: reg_0528 <= imem03_in[79:76];
    87: reg_0528 <= imem03_in[79:76];
    endcase
  end

  // REG#529の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0529 <= imem04_in[55:52];
    18: reg_0529 <= imem04_in[55:52];
    41: reg_0529 <= imem04_in[55:52];
    endcase
  end

  // REG#530の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0530 <= imem04_in[23:20];
    20: reg_0530 <= imem02_in[39:36];
    81: reg_0530 <= imem04_in[23:20];
    83: reg_0530 <= imem02_in[39:36];
    endcase
  end

  // REG#531の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0531 <= imem04_in[115:112];
    20: reg_0531 <= imem02_in[79:76];
    82: reg_0531 <= imem02_in[79:76];
    86: reg_0531 <= imem05_in[95:92];
    endcase
  end

  // REG#532の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0532 <= imem04_in[95:92];
    20: reg_0532 <= imem02_in[115:112];
    82: reg_0532 <= imem02_in[115:112];
    84: reg_0532 <= imem02_in[115:112];
    endcase
  end

  // REG#533の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0533 <= imem04_in[107:104];
    20: reg_0533 <= imem02_in[23:20];
    81: reg_0533 <= imem04_in[107:104];
    83: reg_0533 <= imem02_in[23:20];
    endcase
  end

  // REG#534の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0534 <= imem04_in[51:48];
    18: reg_0534 <= imem04_in[51:48];
    33: reg_0534 <= op2_01_out;
    60: reg_0534 <= imem06_in[11:8];
    69: reg_0534 <= imem06_in[11:8];
    71: reg_0534 <= imem02_in[15:12];
    82: reg_0534 <= imem04_in[51:48];
    endcase
  end

  // REG#535の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0535 <= imem04_in[59:56];
    20: reg_0535 <= imem02_in[59:56];
    82: reg_0535 <= imem04_in[59:56];
    endcase
  end

  // REG#536の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0536 <= imem04_in[15:12];
    20: reg_0536 <= imem04_in[15:12];
    23: reg_0536 <= imem04_in[91:88];
    82: reg_0536 <= imem04_in[91:88];
    endcase
  end

  // REG#537の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0537 <= imem04_in[71:68];
    20: reg_0537 <= imem04_in[71:68];
    23: reg_0537 <= imem04_in[51:48];
    82: reg_0537 <= imem04_in[71:68];
    endcase
  end

  // REG#538の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0538 <= op1_04_out;
    20: reg_0538 <= imem02_in[99:96];
    82: reg_0538 <= imem02_in[99:96];
    86: reg_0538 <= imem05_in[15:12];
    endcase
  end

  // REG#539の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0539 <= imem04_in[63:60];
    20: reg_0539 <= imem02_in[71:68];
    82: reg_0539 <= imem04_in[63:60];
    endcase
  end

  // REG#540の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0540 <= imem04_in[91:88];
    20: reg_0540 <= imem02_in[55:52];
    84: reg_0540 <= imem02_in[55:52];
    endcase
  end

  // REG#541の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0541 <= imem04_in[119:116];
    20: reg_0541 <= imem02_in[11:8];
    83: reg_0541 <= imem02_in[11:8];
    endcase
  end

  // REG#542の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0542 <= imem04_in[47:44];
    20: reg_0542 <= imem04_in[47:44];
    23: reg_0542 <= imem04_in[47:44];
    82: reg_0542 <= imem04_in[47:44];
    endcase
  end

  // REG#543の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0543 <= imem04_in[3:0];
    20: reg_0543 <= op2_02_out;
    58: reg_0543 <= op2_02_out;
    endcase
  end

  // REG#544の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0544 <= imem04_in[7:4];
    21: reg_0544 <= imem04_in[7:4];
    23: reg_0544 <= imem04_in[19:16];
    82: reg_0544 <= imem04_in[19:16];
    endcase
  end

  // REG#545の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0545 <= imem04_in[11:8];
    21: reg_0545 <= imem04_in[11:8];
    23: reg_0545 <= imem04_in[11:8];
    82: reg_0545 <= imem04_in[11:8];
    endcase
  end

  // REG#546の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0546 <= imem04_in[87:84];
    20: reg_0546 <= op2_03_out;
    59: reg_0546 <= op2_03_out;
    endcase
  end

  // REG#547の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0547 <= imem04_in[127:124];
    23: reg_0547 <= imem04_in[127:124];
    81: reg_0547 <= imem04_in[127:124];
    86: reg_0547 <= imem05_in[123:120];
    endcase
  end

  // REG#548の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0548 <= imem04_in[67:64];
    22: reg_0548 <= imem04_in[67:64];
    24: reg_0548 <= imem01_in[107:104];
    44: reg_0548 <= imem02_in[99:96];
    62: reg_0548 <= imem02_in[99:96];
    71: reg_0548 <= imem02_in[99:96];
    82: reg_0548 <= imem04_in[67:64];
    endcase
  end

  // REG#549の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0549 <= imem04_in[79:76];
    24: reg_0549 <= imem01_in[71:68];
    45: reg_0549 <= imem04_in[115:112];
    48: reg_0549 <= imem04_in[79:76];
    57: reg_0549 <= imem04_in[115:112];
    60: reg_0549 <= imem06_in[79:76];
    69: reg_0549 <= imem03_in[83:80];
    endcase
  end

  // REG#550の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0550 <= imem04_in[35:32];
    22: reg_0550 <= imem04_in[35:32];
    24: reg_0550 <= imem01_in[115:112];
    48: reg_0550 <= imem01_in[115:112];
    67: reg_0550 <= imem05_in[67:64];
    72: reg_0550 <= imem05_in[67:64];
    endcase
  end

  // REG#551の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0551 <= imem04_in[103:100];
    21: reg_0551 <= imem04_in[103:100];
    23: reg_0551 <= imem04_in[103:100];
    82: reg_0551 <= imem04_in[103:100];
    endcase
  end

  // REG#552の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0552 <= imem04_in[39:36];
    23: reg_0552 <= imem04_in[39:36];
    81: reg_0552 <= imem04_in[39:36];
    86: reg_0552 <= imem05_in[23:20];
    endcase
  end

  // REG#553の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0553 <= imem04_in[31:28];
    23: reg_0553 <= imem04_in[31:28];
    82: reg_0553 <= imem04_in[31:28];
    endcase
  end

  // REG#554の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0554 <= imem04_in[83:80];
    21: reg_0554 <= imem04_in[83:80];
    23: reg_0554 <= imem04_in[83:80];
    82: reg_0554 <= imem04_in[83:80];
    endcase
  end

  // REG#555の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0555 <= imem04_in[75:72];
    21: reg_0555 <= imem04_in[75:72];
    23: reg_0555 <= imem04_in[75:72];
    82: reg_0555 <= imem04_in[75:72];
    endcase
  end

  // REG#556の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0556 <= imem04_in[123:120];
    23: reg_0556 <= imem04_in[123:120];
    82: reg_0556 <= imem04_in[123:120];
    endcase
  end

  // REG#557の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0557 <= imem04_in[19:16];
    22: reg_0557 <= imem04_in[19:16];
    24: reg_0557 <= imem01_in[103:100];
    48: reg_0557 <= imem01_in[103:100];
    67: reg_0557 <= imem01_in[103:100];
    69: reg_0557 <= imem03_in[115:112];
    endcase
  end

  // REG#558の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0558 <= imem04_in[99:96];
    23: reg_0558 <= imem04_in[99:96];
    82: reg_0558 <= imem04_in[99:96];
    endcase
  end

  // REG#559の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0559 <= imem04_in[111:108];
    22: reg_0559 <= imem04_in[111:108];
    24: reg_0559 <= imem01_in[127:124];
    46: reg_0559 <= imem01_in[127:124];
    51: reg_0559 <= imem01_in[127:124];
    54: reg_0559 <= imem03_in[47:44];
    87: reg_0559 <= imem03_in[47:44];
    endcase
  end

  // REG#560の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0560 <= imem04_in[27:24];
    21: reg_0560 <= imem04_in[27:24];
    23: reg_0560 <= imem04_in[27:24];
    81: reg_0560 <= imem04_in[27:24];
    86: reg_0560 <= imem05_in[127:124];
    endcase
  end

  // REG#561の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0561 <= op1_05_out;
    20: reg_0561 <= op1_05_out;
    21: reg_0561 <= op1_05_out;
    22: reg_0561 <= op1_05_out;
    23: reg_0561 <= op1_05_out;
    27: reg_0561 <= imem03_in[31:28];
    66: reg_0561 <= op2_02_out;
    81: reg_0561 <= op2_02_out;
    89: reg_0561 <= imem03_in[31:28];
    endcase
  end

  // REG#562の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0562 <= op1_06_out;
    20: reg_0562 <= op1_06_out;
    21: reg_0562 <= op1_06_out;
    22: reg_0562 <= op1_06_out;
    23: reg_0562 <= op1_06_out;
    24: reg_0562 <= op1_06_out;
    27: reg_0562 <= imem03_in[79:76];
    69: reg_0562 <= imem03_in[79:76];
    endcase
  end

  // REG#563の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0563 <= imem03_in[67:64];
    24: reg_0563 <= imem01_in[75:72];
    48: reg_0563 <= imem01_in[75:72];
    62: reg_0563 <= imem02_in[43:40];
    70: reg_0563 <= imem06_in[35:32];
    86: reg_0563 <= imem05_in[19:16];
    endcase
  end

  // REG#564の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0564 <= op1_07_out;
    22: reg_0564 <= op1_07_out;
    23: reg_0564 <= op1_07_out;
    24: reg_0564 <= op1_07_out;
    25: reg_0564 <= op1_07_out;
    27: reg_0564 <= imem03_in[39:36];
    69: reg_0564 <= imem03_in[39:36];
    endcase
  end

  // REG#565の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0565 <= op1_08_out;
    22: reg_0565 <= op1_08_out;
    23: reg_0565 <= op1_08_out;
    24: reg_0565 <= op1_08_out;
    25: reg_0565 <= op1_08_out;
    26: reg_0565 <= op1_08_out;
    27: reg_0565 <= op1_08_out;
    30: reg_0565 <= imem03_in[43:40];
    51: reg_0565 <= imem02_in[55:52];
    endcase
  end

  // REG#566の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0566 <= op1_09_out;
    25: reg_0566 <= op1_09_out;
    26: reg_0566 <= op1_09_out;
    27: reg_0566 <= op1_09_out;
    28: reg_0566 <= op1_09_out;
    30: reg_0566 <= imem03_in[23:20];
    51: reg_0566 <= imem02_in[119:116];
    endcase
  end

  // REG#567の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0567 <= op1_10_out;
    25: reg_0567 <= op1_10_out;
    26: reg_0567 <= op1_10_out;
    27: reg_0567 <= op1_10_out;
    28: reg_0567 <= op1_10_out;
    29: reg_0567 <= op1_10_out;
    30: reg_0567 <= op1_10_out;
    40: reg_0567 <= imem01_in[51:48];
    92: reg_0567 <= imem01_in[51:48];
    94: reg_0567 <= imem01_in[51:48];
    endcase
  end

  // REG#568の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0568 <= imem03_in[43:40];
    27: reg_0568 <= imem03_in[43:40];
    69: reg_0568 <= imem03_in[43:40];
    endcase
  end

  // REG#569の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0569 <= imem03_in[55:52];
    27: reg_0569 <= imem03_in[75:72];
    69: reg_0569 <= imem03_in[75:72];
    endcase
  end

  // REG#570の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0570 <= imem03_in[119:116];
    27: reg_0570 <= imem03_in[127:124];
    69: reg_0570 <= imem03_in[127:124];
    endcase
  end

  // REG#571の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0571 <= imem03_in[19:16];
    27: reg_0571 <= imem03_in[63:60];
    69: reg_0571 <= imem03_in[19:16];
    endcase
  end

  // REG#572の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0572 <= imem03_in[47:44];
    27: reg_0572 <= imem03_in[83:80];
    69: reg_0572 <= imem03_in[47:44];
    87: reg_0572 <= imem03_in[127:124];
    endcase
  end

  // REG#573の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0573 <= imem03_in[23:20];
    27: reg_0573 <= imem03_in[23:20];
    68: reg_0573 <= imem03_in[23:20];
    70: reg_0573 <= imem06_in[3:0];
    87: reg_0573 <= imem03_in[23:20];
    endcase
  end

  // REG#574の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0574 <= op1_11_out;
    26: reg_0574 <= op1_11_out;
    27: reg_0574 <= op1_11_out;
    28: reg_0574 <= op1_11_out;
    29: reg_0574 <= op1_11_out;
    30: reg_0574 <= op1_11_out;
    31: reg_0574 <= op1_11_out;
    40: reg_0574 <= imem01_in[39:36];
    92: reg_0574 <= imem01_in[39:36];
    94: reg_0574 <= imem01_in[39:36];
    endcase
  end

  // REG#575の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0575 <= op1_12_out;
    27: reg_0575 <= imem03_in[27:24];
    69: reg_0575 <= imem03_in[27:24];
    endcase
  end

  // REG#576の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0576 <= imem03_in[127:124];
    28: reg_0576 <= imem06_in[119:116];
    57: reg_0576 <= imem06_in[119:116];
    85: reg_0576 <= imem06_in[119:116];
    endcase
  end

  // REG#577の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0577 <= imem06_in[95:92];
    28: reg_0577 <= imem06_in[31:28];
    56: reg_0577 <= imem06_in[31:28];
    endcase
  end

  // REG#578の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0578 <= imem03_in[99:96];
    30: reg_0578 <= imem03_in[99:96];
    52: reg_0578 <= imem03_in[75:72];
    57: reg_0578 <= imem06_in[27:24];
    85: reg_0578 <= imem06_in[27:24];
    endcase
  end

  // REG#579の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0579 <= imem03_in[35:32];
    30: reg_0579 <= imem03_in[35:32];
    54: reg_0579 <= imem03_in[35:32];
    86: reg_0579 <= imem05_in[115:112];
    endcase
  end

  // REG#580の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0580 <= imem03_in[95:92];
    30: reg_0580 <= imem03_in[95:92];
    52: reg_0580 <= imem03_in[95:92];
    57: reg_0580 <= imem06_in[107:104];
    84: reg_0580 <= imem06_in[107:104];
    86: reg_0580 <= imem05_in[67:64];
    endcase
  end

  // REG#581の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0581 <= imem03_in[107:104];
    30: reg_0581 <= imem03_in[107:104];
    51: reg_0581 <= imem02_in[39:36];
    endcase
  end

  // REG#582の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0582 <= imem03_in[15:12];
    30: reg_0582 <= imem03_in[15:12];
    54: reg_0582 <= imem03_in[15:12];
    87: reg_0582 <= imem03_in[15:12];
    endcase
  end

  // REG#583の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0583 <= imem03_in[39:36];
    30: reg_0583 <= imem03_in[39:36];
    52: reg_0583 <= imem03_in[39:36];
    57: reg_0583 <= imem06_in[95:92];
    86: reg_0583 <= imem05_in[47:44];
    endcase
  end

  // REG#584の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0584 <= imem03_in[79:76];
    30: reg_0584 <= imem03_in[79:76];
    44: reg_0584 <= imem02_in[39:36];
    62: reg_0584 <= imem02_in[39:36];
    71: reg_0584 <= imem02_in[39:36];
    84: reg_0584 <= imem02_in[39:36];
    endcase
  end

  // REG#585の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0585 <= imem03_in[83:80];
    30: reg_0585 <= imem03_in[83:80];
    45: reg_0585 <= imem04_in[31:28];
    48: reg_0585 <= imem04_in[31:28];
    58: reg_0585 <= imem04_in[31:28];
    endcase
  end

  // REG#586の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0586 <= imem03_in[11:8];
    30: reg_0586 <= imem03_in[11:8];
    51: reg_0586 <= imem02_in[35:32];
    endcase
  end

  // REG#587の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0587 <= imem03_in[51:48];
    30: reg_0587 <= imem03_in[51:48];
    51: reg_0587 <= imem02_in[15:12];
    endcase
  end

  // REG#588の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0588 <= imem03_in[115:112];
    30: reg_0588 <= imem03_in[115:112];
    52: reg_0588 <= imem03_in[115:112];
    54: reg_0588 <= imem03_in[115:112];
    86: reg_0588 <= imem03_in[115:112];
    88: reg_0588 <= imem03_in[115:112];
    endcase
  end

  // REG#589の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0589 <= imem03_in[71:68];
    30: reg_0589 <= imem03_in[71:68];
    54: reg_0589 <= imem03_in[23:20];
    87: reg_0589 <= imem03_in[95:92];
    endcase
  end

  // REG#590の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0590 <= imem03_in[123:120];
    30: reg_0590 <= imem03_in[123:120];
    51: reg_0590 <= imem02_in[111:108];
    endcase
  end

  // REG#591の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0591 <= imem03_in[63:60];
    30: reg_0591 <= imem03_in[63:60];
    54: reg_0591 <= imem03_in[63:60];
    87: reg_0591 <= imem03_in[63:60];
    endcase
  end

  // REG#592の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0592 <= imem03_in[59:56];
    30: reg_0592 <= imem03_in[59:56];
    52: reg_0592 <= imem01_in[43:40];
    endcase
  end

  // REG#593の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0593 <= imem03_in[87:84];
    30: reg_0593 <= imem03_in[87:84];
    52: reg_0593 <= imem03_in[87:84];
    57: reg_0593 <= imem06_in[103:100];
    85: reg_0593 <= imem06_in[103:100];
    endcase
  end

  // REG#594の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0594 <= imem03_in[75:72];
    30: reg_0594 <= imem03_in[75:72];
    51: reg_0594 <= imem02_in[75:72];
    endcase
  end

  // REG#595の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0595 <= imem03_in[111:108];
    30: reg_0595 <= imem03_in[111:108];
    54: reg_0595 <= imem03_in[111:108];
    87: reg_0595 <= imem03_in[111:108];
    endcase
  end

  // REG#596の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0596 <= imem03_in[27:24];
    30: reg_0596 <= imem03_in[55:52];
    52: reg_0596 <= imem03_in[55:52];
    54: reg_0596 <= imem03_in[55:52];
    86: reg_0596 <= imem03_in[27:24];
    88: reg_0596 <= imem03_in[27:24];
    endcase
  end

  // REG#597の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0597 <= imem03_in[103:100];
    30: reg_0597 <= imem03_in[103:100];
    54: reg_0597 <= imem03_in[27:24];
    87: reg_0597 <= imem03_in[27:24];
    endcase
  end

  // REG#598の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0598 <= imem03_in[3:0];
    30: reg_0598 <= imem03_in[3:0];
    48: reg_0598 <= imem04_in[43:40];
    58: reg_0598 <= imem04_in[43:40];
    endcase
  end

  // REG#599の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0599 <= imem03_in[31:28];
    30: reg_0599 <= imem03_in[31:28];
    54: reg_0599 <= imem03_in[31:28];
    87: reg_0599 <= imem03_in[55:52];
    endcase
  end

  // REG#600の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0600 <= imem03_in[91:88];
    30: reg_0600 <= imem03_in[91:88];
    54: reg_0600 <= imem03_in[91:88];
    87: reg_0600 <= imem03_in[91:88];
    endcase
  end

  // REG#601の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0601 <= imem06_in[123:120];
    30: reg_0601 <= imem03_in[19:16];
    52: reg_0601 <= imem01_in[83:80];
    endcase
  end

  // REG#602の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0602 <= imem03_in[7:4];
    30: reg_0602 <= imem03_in[7:4];
    54: reg_0602 <= imem03_in[7:4];
    87: reg_0602 <= imem03_in[7:4];
    endcase
  end

  // REG#603の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0603 <= op1_13_out;
    29: reg_0603 <= op1_13_out;
    30: reg_0603 <= op1_13_out;
    34: reg_0603 <= op1_13_out;
    40: reg_0603 <= imem01_in[91:88];
    endcase
  end

  // REG#604の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0604 <= imem06_in[19:16];
    31: reg_0604 <= imem06_in[11:8];
    35: reg_0604 <= imem06_in[19:16];
    38: reg_0604 <= imem06_in[19:16];
    54: reg_0604 <= imem03_in[39:36];
    87: reg_0604 <= imem03_in[39:36];
    endcase
  end

  // REG#605の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0605 <= imem06_in[51:48];
    31: reg_0605 <= imem06_in[95:92];
    35: reg_0605 <= imem06_in[51:48];
    38: reg_0605 <= imem06_in[51:48];
    56: reg_0605 <= imem06_in[51:48];
    endcase
  end

  // REG#606の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0606 <= imem06_in[67:64];
    31: reg_0606 <= imem06_in[79:76];
    35: reg_0606 <= imem06_in[79:76];
    38: reg_0606 <= imem06_in[79:76];
    56: reg_0606 <= imem06_in[79:76];
    endcase
  end

  // REG#607の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0607 <= imem06_in[27:24];
    36: reg_0607 <= imem06_in[27:24];
    60: reg_0607 <= imem06_in[27:24];
    69: reg_0607 <= imem06_in[27:24];
    71: reg_0607 <= imem02_in[83:80];
    82: reg_0607 <= imem02_in[83:80];
    87: reg_0607 <= imem06_in[27:24];
    89: reg_0607 <= imem03_in[19:16];
    endcase
  end

  // REG#608の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0608 <= imem06_in[91:88];
    34: reg_0608 <= imem06_in[91:88];
    38: reg_0608 <= imem06_in[91:88];
    57: reg_0608 <= imem06_in[91:88];
    85: reg_0608 <= imem06_in[91:88];
    endcase
  end

  // REG#609の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0609 <= imem06_in[71:68];
    34: reg_0609 <= imem06_in[71:68];
    38: reg_0609 <= imem06_in[71:68];
    56: reg_0609 <= imem06_in[71:68];
    88: reg_0609 <= imem06_in[71:68];
    endcase
  end

  // REG#610の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0610 <= imem06_in[11:8];
    35: reg_0610 <= imem06_in[11:8];
    37: reg_0610 <= imem06_in[11:8];
    41: reg_0610 <= imem04_in[127:124];
    endcase
  end

  // REG#611の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0611 <= imem06_in[79:76];
    41: reg_0611 <= imem04_in[59:56];
    endcase
  end

  // REG#612の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0612 <= imem06_in[127:124];
    35: reg_0612 <= imem06_in[127:124];
    38: reg_0612 <= imem06_in[127:124];
    54: reg_0612 <= imem00_in[43:40];
    88: reg_0612 <= imem06_in[35:32];
    endcase
  end

  // REG#613の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0613 <= imem06_in[39:36];
    35: reg_0613 <= imem06_in[39:36];
    38: reg_0613 <= imem06_in[39:36];
    57: reg_0613 <= imem06_in[39:36];
    85: reg_0613 <= imem06_in[39:36];
    endcase
  end

  // REG#614の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0614 <= imem06_in[3:0];
    34: reg_0614 <= imem06_in[3:0];
    36: reg_0614 <= imem06_in[3:0];
    58: reg_0614 <= imem04_in[3:0];
    endcase
  end

  // REG#615の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0615 <= imem06_in[119:116];
    34: reg_0615 <= imem06_in[119:116];
    37: reg_0615 <= imem06_in[119:116];
    41: reg_0615 <= imem04_in[43:40];
    endcase
  end

  // REG#616の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0616 <= imem06_in[59:56];
    34: reg_0616 <= imem06_in[59:56];
    37: reg_0616 <= imem06_in[59:56];
    41: reg_0616 <= imem04_in[79:76];
    endcase
  end

  // REG#617の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0617 <= imem06_in[47:44];
    35: reg_0617 <= imem06_in[47:44];
    37: reg_0617 <= imem06_in[47:44];
    41: reg_0617 <= imem04_in[119:116];
    endcase
  end

  // REG#618の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0618 <= imem06_in[99:96];
    35: reg_0618 <= imem06_in[99:96];
    38: reg_0618 <= imem06_in[99:96];
    56: reg_0618 <= imem06_in[99:96];
    endcase
  end

  // REG#619の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0619 <= imem06_in[83:80];
    34: reg_0619 <= imem06_in[83:80];
    38: reg_0619 <= imem06_in[83:80];
    56: reg_0619 <= imem06_in[83:80];
    endcase
  end

  // REG#620の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0620 <= imem06_in[43:40];
    36: reg_0620 <= imem06_in[43:40];
    60: reg_0620 <= imem06_in[43:40];
    70: reg_0620 <= imem06_in[43:40];
    88: reg_0620 <= imem06_in[43:40];
    endcase
  end

  // REG#621の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0621 <= imem06_in[55:52];
    36: reg_0621 <= imem06_in[55:52];
    59: reg_0621 <= imem06_in[55:52];
    62: reg_0621 <= imem02_in[47:44];
    71: reg_0621 <= imem02_in[47:44];
    88: reg_0621 <= imem06_in[55:52];
    endcase
  end

  // REG#622の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0622 <= imem06_in[111:108];
    35: reg_0622 <= imem06_in[111:108];
    38: reg_0622 <= imem06_in[111:108];
    55: reg_0622 <= imem06_in[111:108];
    58: reg_0622 <= imem04_in[47:44];
    endcase
  end

  // REG#623の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0623 <= imem06_in[115:112];
    36: reg_0623 <= imem06_in[115:112];
    60: reg_0623 <= imem06_in[115:112];
    69: reg_0623 <= imem03_in[119:116];
    endcase
  end

  // REG#624の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0624 <= imem06_in[35:32];
    35: reg_0624 <= imem06_in[35:32];
    38: reg_0624 <= imem06_in[35:32];
    56: reg_0624 <= imem06_in[35:32];
    endcase
  end

  // REG#625の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0625 <= imem06_in[15:12];
    35: reg_0625 <= imem06_in[15:12];
    38: reg_0625 <= imem06_in[15:12];
    56: reg_0625 <= imem06_in[15:12];
    endcase
  end

  // REG#626の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0626 <= imem06_in[75:72];
    35: reg_0626 <= imem06_in[75:72];
    37: reg_0626 <= imem06_in[75:72];
    41: reg_0626 <= imem04_in[123:120];
    endcase
  end

  // REG#627の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0627 <= imem06_in[107:104];
    35: reg_0627 <= imem06_in[107:104];
    41: reg_0627 <= imem04_in[107:104];
    endcase
  end

  // REG#628の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0628 <= imem06_in[7:4];
    35: reg_0628 <= imem06_in[7:4];
    38: reg_0628 <= imem06_in[7:4];
    57: reg_0628 <= imem06_in[7:4];
    85: reg_0628 <= imem06_in[7:4];
    endcase
  end

  // REG#629の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0629 <= imem06_in[23:20];
    35: reg_0629 <= imem06_in[23:20];
    37: reg_0629 <= imem06_in[23:20];
    41: reg_0629 <= imem04_in[87:84];
    endcase
  end

  // REG#630の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0630 <= imem06_in[31:28];
    35: reg_0630 <= imem06_in[31:28];
    38: reg_0630 <= imem06_in[31:28];
    57: reg_0630 <= imem06_in[31:28];
    85: reg_0630 <= imem06_in[31:28];
    endcase
  end

  // REG#631の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0631 <= imem06_in[63:60];
    35: reg_0631 <= imem06_in[63:60];
    41: reg_0631 <= imem04_in[51:48];
    endcase
  end

  // REG#632の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0632 <= imem06_in[103:100];
    36: reg_0632 <= imem06_in[103:100];
    60: reg_0632 <= imem06_in[103:100];
    70: reg_0632 <= imem06_in[103:100];
    84: reg_0632 <= imem06_in[103:100];
    88: reg_0632 <= imem06_in[103:100];
    endcase
  end

  // REG#633の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0633 <= imem06_in[87:84];
    35: reg_0633 <= imem06_in[87:84];
    38: reg_0633 <= imem06_in[87:84];
    54: reg_0633 <= imem00_in[111:108];
    88: reg_0633 <= imem06_in[87:84];
    endcase
  end

  // REG#634の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0634 <= op1_14_out;
    34: reg_0634 <= op1_14_out;
    37: reg_0634 <= op1_14_out;
    38: reg_0634 <= op1_14_out;
    39: reg_0634 <= op1_14_out;
    40: reg_0634 <= op1_14_out;
    42: reg_0634 <= op1_14_out;
    43: reg_0634 <= op1_14_out;
    44: reg_0634 <= op1_14_out;
    46: reg_0634 <= op1_14_out;
    47: reg_0634 <= op1_14_out;
    51: reg_0634 <= op1_14_out;
    54: reg_0634 <= imem00_in[123:120];
    89: reg_0634 <= imem00_in[123:120];
    endcase
  end

  // REG#635の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0635 <= op1_15_out;
    42: reg_0635 <= imem07_in[51:48];
    endcase
  end

  // REG#636の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0636 <= imem02_in[115:112];
    42: reg_0636 <= imem07_in[31:28];
    endcase
  end

  // REG#637の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0637 <= imem02_in[35:32];
    44: reg_0637 <= imem02_in[35:32];
    62: reg_0637 <= imem02_in[35:32];
    69: reg_0637 <= imem03_in[103:100];
    endcase
  end

  // REG#638の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0638 <= imem02_in[83:80];
    44: reg_0638 <= imem02_in[83:80];
    57: reg_0638 <= imem06_in[99:96];
    85: reg_0638 <= imem06_in[99:96];
    endcase
  end

  // REG#639の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0639 <= imem02_in[63:60];
    44: reg_0639 <= imem02_in[63:60];
    62: reg_0639 <= imem02_in[63:60];
    71: reg_0639 <= imem02_in[63:60];
    83: reg_0639 <= imem02_in[63:60];
    endcase
  end

  // REG#640の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0640 <= imem02_in[75:72];
    45: reg_0640 <= imem04_in[55:52];
    48: reg_0640 <= imem04_in[91:88];
    58: reg_0640 <= imem04_in[91:88];
    endcase
  end

  // REG#641の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0641 <= imem02_in[91:88];
    44: reg_0641 <= imem02_in[91:88];
    62: reg_0641 <= imem02_in[91:88];
    70: reg_0641 <= imem02_in[91:88];
    72: reg_0641 <= imem05_in[59:56];
    endcase
  end

  // REG#642の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0642 <= imem02_in[3:0];
    44: reg_0642 <= imem02_in[3:0];
    60: reg_0642 <= imem06_in[67:64];
    69: reg_0642 <= imem06_in[67:64];
    71: reg_0642 <= imem02_in[3:0];
    83: reg_0642 <= imem02_in[3:0];
    endcase
  end

  // REG#643の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0643 <= imem02_in[103:100];
    45: reg_0643 <= imem04_in[63:60];
    48: reg_0643 <= imem04_in[63:60];
    58: reg_0643 <= imem04_in[63:60];
    endcase
  end

  // REG#644の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0644 <= imem02_in[99:96];
    43: reg_0644 <= imem02_in[99:96];
    48: reg_0644 <= imem04_in[107:104];
    58: reg_0644 <= imem04_in[107:104];
    endcase
  end

  // REG#645の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0645 <= imem02_in[11:8];
    43: reg_0645 <= imem02_in[11:8];
    48: reg_0645 <= imem01_in[43:40];
    61: reg_0645 <= imem02_in[11:8];
    68: reg_0645 <= imem01_in[43:40];
    93: reg_0645 <= imem01_in[43:40];
    endcase
  end

  // REG#646の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0646 <= imem02_in[39:36];
    43: reg_0646 <= imem02_in[39:36];
    48: reg_0646 <= imem01_in[3:0];
    67: reg_0646 <= imem01_in[3:0];
    69: reg_0646 <= imem03_in[63:60];
    endcase
  end

  // REG#647の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0647 <= imem02_in[71:68];
    44: reg_0647 <= imem02_in[71:68];
    62: reg_0647 <= imem02_in[71:68];
    71: reg_0647 <= imem02_in[71:68];
    83: reg_0647 <= imem02_in[71:68];
    endcase
  end

  // REG#648の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0648 <= imem02_in[79:76];
    43: reg_0648 <= imem02_in[79:76];
    47: reg_0648 <= op2_00_out;
    62: reg_0648 <= op2_00_out;
    69: reg_0648 <= imem03_in[3:0];
    endcase
  end

  // REG#649の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0649 <= imem02_in[87:84];
    43: reg_0649 <= imem02_in[87:84];
    48: reg_0649 <= imem01_in[63:60];
    69: reg_0649 <= imem03_in[123:120];
    endcase
  end

  // REG#650の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0650 <= imem02_in[7:4];
    44: reg_0650 <= imem02_in[7:4];
    62: reg_0650 <= imem02_in[7:4];
    71: reg_0650 <= imem02_in[7:4];
    88: reg_0650 <= imem06_in[107:104];
    endcase
  end

  // REG#651の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0651 <= imem02_in[67:64];
    44: reg_0651 <= imem02_in[67:64];
    62: reg_0651 <= imem02_in[67:64];
    70: reg_0651 <= imem06_in[55:52];
    88: reg_0651 <= imem06_in[11:8];
    endcase
  end

  // REG#652の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0652 <= imem02_in[119:116];
    43: reg_0652 <= imem02_in[119:116];
    48: reg_0652 <= imem01_in[107:104];
    67: reg_0652 <= imem01_in[107:104];
    70: reg_0652 <= imem06_in[79:76];
    87: reg_0652 <= imem06_in[79:76];
    88: reg_0652 <= op2_01_out;
    endcase
  end

  // REG#653の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0653 <= imem02_in[27:24];
    43: reg_0653 <= imem02_in[27:24];
    48: reg_0653 <= imem01_in[19:16];
    68: reg_0653 <= imem01_in[19:16];
    endcase
  end

  // REG#654の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0654 <= imem02_in[31:28];
    44: reg_0654 <= imem02_in[31:28];
    57: reg_0654 <= imem06_in[47:44];
    85: reg_0654 <= imem06_in[47:44];
    endcase
  end

  // REG#655の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0655 <= imem02_in[23:20];
    44: reg_0655 <= imem02_in[23:20];
    62: reg_0655 <= imem02_in[95:92];
    71: reg_0655 <= imem02_in[95:92];
    82: reg_0655 <= imem02_in[23:20];
    88: reg_0655 <= imem06_in[3:0];
    endcase
  end

  // REG#656の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0656 <= imem02_in[59:56];
    44: reg_0656 <= imem02_in[59:56];
    60: reg_0656 <= imem06_in[55:52];
    69: reg_0656 <= imem06_in[55:52];
    71: reg_0656 <= imem02_in[59:56];
    83: reg_0656 <= imem02_in[59:56];
    endcase
  end

  // REG#657の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0657 <= imem02_in[51:48];
    44: reg_0657 <= imem02_in[51:48];
    62: reg_0657 <= imem02_in[51:48];
    70: reg_0657 <= imem06_in[63:60];
    88: reg_0657 <= imem06_in[63:60];
    endcase
  end

  // REG#658の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0658 <= imem02_in[15:12];
    44: reg_0658 <= imem02_in[15:12];
    54: reg_0658 <= imem00_in[75:72];
    90: reg_0658 <= imem00_in[75:72];
    endcase
  end

  // REG#659の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0659 <= imem02_in[111:108];
    44: reg_0659 <= imem02_in[111:108];
    57: reg_0659 <= imem06_in[43:40];
    85: reg_0659 <= imem06_in[43:40];
    endcase
  end

  // REG#660の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0660 <= imem02_in[47:44];
    44: reg_0660 <= imem02_in[47:44];
    52: reg_0660 <= imem01_in[63:60];
    endcase
  end

  // REG#661の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0661 <= imem02_in[55:52];
    44: reg_0661 <= imem02_in[55:52];
    62: reg_0661 <= imem02_in[55:52];
    70: reg_0661 <= imem06_in[95:92];
    88: reg_0661 <= imem06_in[95:92];
    endcase
  end

  // REG#662の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0662 <= imem02_in[95:92];
    44: reg_0662 <= imem02_in[95:92];
    56: reg_0662 <= op2_02_out;
    endcase
  end

  // REG#663の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0663 <= imem02_in[127:124];
    48: reg_0663 <= imem01_in[35:32];
    67: reg_0663 <= imem01_in[35:32];
    70: reg_0663 <= imem06_in[23:20];
    88: reg_0663 <= imem06_in[23:20];
    endcase
  end

  // REG#664の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0664 <= imem02_in[43:40];
    44: reg_0664 <= imem02_in[43:40];
    61: reg_0664 <= imem02_in[43:40];
    70: reg_0664 <= imem06_in[67:64];
    88: reg_0664 <= imem06_in[67:64];
    endcase
  end

  // REG#665の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0665 <= imem02_in[107:104];
    44: reg_0665 <= imem02_in[107:104];
    61: reg_0665 <= imem02_in[107:104];
    70: reg_0665 <= imem02_in[107:104];
    72: reg_0665 <= imem05_in[107:104];
    endcase
  end

  // REG#666の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0666 <= imem02_in[19:16];
    44: reg_0666 <= imem02_in[19:16];
    62: reg_0666 <= imem02_in[19:16];
    70: reg_0666 <= imem02_in[19:16];
    72: reg_0666 <= imem05_in[39:36];
    endcase
  end

  // REG#667の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0667 <= imem02_in[123:120];
    44: reg_0667 <= imem02_in[123:120];
    60: reg_0667 <= imem06_in[3:0];
    70: reg_0667 <= imem02_in[123:120];
    72: reg_0667 <= imem05_in[27:24];
    endcase
  end

  // REG#668の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0668 <= imem00_in[95:92];
    48: reg_0668 <= imem01_in[27:24];
    68: reg_0668 <= imem01_in[27:24];
    endcase
  end

  // REG#669の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0669 <= imem00_in[123:120];
    52: reg_0669 <= imem01_in[79:76];
    endcase
  end

  // REG#670の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0670 <= imem00_in[63:60];
    52: reg_0670 <= imem01_in[35:32];
    endcase
  end

  // REG#671の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0671 <= imem00_in[87:84];
    52: reg_0671 <= imem01_in[87:84];
    endcase
  end

  // REG#672の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0672 <= imem00_in[35:32];
    52: reg_0672 <= imem01_in[55:52];
    endcase
  end

  // REG#673の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0673 <= imem00_in[111:108];
    52: reg_0673 <= imem01_in[19:16];
    endcase
  end

  // REG#674の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0674 <= imem00_in[83:80];
    52: reg_0674 <= imem01_in[103:100];
    endcase
  end

  // REG#675の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0675 <= imem00_in[99:96];
    52: reg_0675 <= imem01_in[71:68];
    endcase
  end

  // REG#676の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0676 <= imem00_in[43:40];
    52: reg_0676 <= imem01_in[99:96];
    endcase
  end

  // REG#677の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0677 <= imem00_in[75:72];
    52: reg_0677 <= imem01_in[67:64];
    endcase
  end

  // REG#678の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0678 <= imem00_in[91:88];
    52: reg_0678 <= imem01_in[115:112];
    endcase
  end

  // REG#679の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0679 <= imem00_in[67:64];
    53: reg_0679 <= imem00_in[67:64];
    58: reg_0679 <= imem04_in[11:8];
    endcase
  end

  // REG#680の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0680 <= imem00_in[103:100];
    54: reg_0680 <= imem00_in[103:100];
    88: reg_0680 <= imem06_in[91:88];
    endcase
  end

  // REG#681の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0681 <= imem00_in[23:20];
    54: reg_0681 <= imem00_in[23:20];
    88: reg_0681 <= imem06_in[15:12];
    endcase
  end

  // REG#682の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0682 <= imem00_in[7:4];
    54: reg_0682 <= imem00_in[7:4];
    87: reg_0682 <= op2_00_out;
    endcase
  end

  // REG#683の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0683 <= imem00_in[19:16];
    54: reg_0683 <= imem00_in[19:16];
    90: reg_0683 <= imem00_in[19:16];
    endcase
  end

  // REG#684の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0684 <= imem00_in[55:52];
    54: reg_0684 <= imem00_in[55:52];
    89: reg_0684 <= imem00_in[55:52];
    endcase
  end

  // REG#685の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0685 <= imem00_in[31:28];
    54: reg_0685 <= imem00_in[31:28];
    90: reg_0685 <= imem00_in[31:28];
    endcase
  end

  // REG#686の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0686 <= imem00_in[59:56];
    54: reg_0686 <= imem00_in[59:56];
    90: reg_0686 <= imem00_in[59:56];
    endcase
  end

  // REG#687の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0687 <= imem00_in[115:112];
    53: reg_0687 <= imem00_in[115:112];
    58: reg_0687 <= imem04_in[39:36];
    endcase
  end

  // REG#688の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0688 <= imem00_in[107:104];
    54: reg_0688 <= imem00_in[107:104];
    90: reg_0688 <= imem00_in[107:104];
    endcase
  end

  // REG#689の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0689 <= imem00_in[51:48];
    54: reg_0689 <= imem00_in[51:48];
    90: reg_0689 <= imem00_in[51:48];
    endcase
  end

  // REG#690の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0690 <= imem00_in[71:68];
    54: reg_0690 <= imem00_in[71:68];
    90: reg_0690 <= imem00_in[71:68];
    endcase
  end

  // REG#691の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0691 <= imem00_in[79:76];
    54: reg_0691 <= imem00_in[79:76];
    90: reg_0691 <= imem00_in[79:76];
    endcase
  end

  // REG#692の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0692 <= imem00_in[119:116];
    54: reg_0692 <= imem00_in[119:116];
    90: reg_0692 <= imem00_in[119:116];
    endcase
  end

  // REG#693の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0693 <= imem00_in[11:8];
    54: reg_0693 <= imem00_in[11:8];
    90: reg_0693 <= imem00_in[11:8];
    endcase
  end

  // REG#694の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0694 <= imem00_in[39:36];
    54: reg_0694 <= imem00_in[39:36];
    endcase
  end

  // REG#695の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0695 <= imem00_in[3:0];
    54: reg_0695 <= imem00_in[3:0];
    90: reg_0695 <= imem00_in[3:0];
    endcase
  end

  // REG#696の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0696 <= imem00_in[27:24];
    54: reg_0696 <= imem00_in[27:24];
    89: reg_0696 <= imem00_in[27:24];
    endcase
  end

  // REG#697の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0697 <= imem00_in[15:12];
    54: reg_0697 <= imem00_in[15:12];
    90: reg_0697 <= imem00_in[15:12];
    endcase
  end

  // REG#698の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0698 <= imem00_in[47:44];
    54: reg_0698 <= imem00_in[47:44];
    90: reg_0698 <= imem00_in[47:44];
    endcase
  end

  // REG#699の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0699 <= imem00_in[127:124];
    54: reg_0699 <= imem00_in[127:124];
    90: reg_0699 <= imem00_in[127:124];
    endcase
  end

  // REG#700の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0700 <= imem07_in[123:120];
    60: reg_0700 <= imem06_in[19:16];
    70: reg_0700 <= imem06_in[19:16];
    88: reg_0700 <= imem06_in[19:16];
    endcase
  end

  // REG#701の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0701 <= imem07_in[115:112];
    69: reg_0701 <= op2_00_out;
    90: reg_0701 <= op2_00_out;
    endcase
  end

  // REG#702の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0702 <= imem07_in[63:60];
    71: reg_0702 <= imem02_in[103:100];
    83: reg_0702 <= imem02_in[103:100];
    endcase
  end

  // REG#703の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0703 <= imem07_in[67:64];
    71: reg_0703 <= imem02_in[79:76];
    84: reg_0703 <= imem02_in[79:76];
    endcase
  end

  // REG#704の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0704 <= imem07_in[15:12];
    71: reg_0704 <= imem02_in[67:64];
    83: reg_0704 <= imem02_in[67:64];
    endcase
  end

  // REG#705の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0705 <= imem07_in[91:88];
    71: reg_0705 <= imem02_in[111:108];
    83: reg_0705 <= imem02_in[111:108];
    endcase
  end

  // REG#706の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0706 <= imem07_in[119:116];
    71: reg_0706 <= op2_02_out;
    endcase
  end

  // REG#707の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0707 <= imem07_in[111:108];
    71: reg_0707 <= op2_03_out;
    endcase
  end

  // REG#708の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0708 <= imem07_in[83:80];
    73: reg_0708 <= imem07_in[83:80];
    78: reg_0708 <= imem07_in[83:80];
    endcase
  end

  // REG#709の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0709 <= imem07_in[87:84];
    73: reg_0709 <= imem07_in[91:88];
    78: reg_0709 <= imem07_in[87:84];
    endcase
  end

  // REG#710の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0710 <= imem07_in[31:28];
    73: reg_0710 <= imem07_in[19:16];
    78: reg_0710 <= imem07_in[19:16];
    endcase
  end

  // REG#711の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0711 <= imem07_in[107:104];
    73: reg_0711 <= imem07_in[107:104];
    78: reg_0711 <= imem07_in[107:104];
    endcase
  end

  // REG#712の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0712 <= imem07_in[71:68];
    73: reg_0712 <= imem07_in[35:32];
    78: reg_0712 <= imem07_in[71:68];
    endcase
  end

  // REG#713の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0713 <= imem07_in[95:92];
    73: reg_0713 <= imem07_in[39:36];
    78: reg_0713 <= imem07_in[95:92];
    endcase
  end

  // REG#714の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0714 <= imem07_in[59:56];
    73: reg_0714 <= imem07_in[127:124];
    77: reg_0714 <= imem07_in[127:124];
    79: reg_0714 <= imem07_in[59:56];
    endcase
  end

  // REG#715の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0715 <= imem07_in[99:96];
    72: reg_0715 <= op1_14_out;
    74: reg_0715 <= op1_14_out;
    78: reg_0715 <= imem07_in[99:96];
    endcase
  end

  // REG#716の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0716 <= imem07_in[11:8];
    73: reg_0716 <= imem07_in[11:8];
    78: reg_0716 <= imem07_in[11:8];
    endcase
  end

  // REG#717の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0717 <= imem07_in[51:48];
    74: reg_0717 <= imem07_in[51:48];
    77: reg_0717 <= imem07_in[51:48];
    79: reg_0717 <= imem07_in[51:48];
    endcase
  end

  // REG#718の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0718 <= imem07_in[103:100];
    77: reg_0718 <= imem07_in[103:100];
    endcase
  end

  // REG#719の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0719 <= imem07_in[19:16];
    74: reg_0719 <= imem07_in[19:16];
    78: reg_0719 <= imem05_in[103:100];
    endcase
  end

  // REG#720の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0720 <= imem07_in[23:20];
    74: reg_0720 <= imem07_in[23:20];
    78: reg_0720 <= imem05_in[59:56];
    endcase
  end

  // REG#721の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0721 <= imem07_in[39:36];
    74: reg_0721 <= imem07_in[39:36];
    78: reg_0721 <= imem07_in[15:12];
    endcase
  end

  // REG#722の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0722 <= imem07_in[3:0];
    74: reg_0722 <= imem07_in[3:0];
    78: reg_0722 <= imem07_in[3:0];
    endcase
  end

  // REG#723の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0723 <= imem07_in[43:40];
    74: reg_0723 <= imem07_in[43:40];
    78: reg_0723 <= imem07_in[27:24];
    endcase
  end

  // REG#724の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0724 <= imem07_in[75:72];
    78: reg_0724 <= imem07_in[115:112];
    endcase
  end

  // REG#725の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0725 <= imem07_in[55:52];
    74: reg_0725 <= imem07_in[55:52];
    78: reg_0725 <= imem07_in[79:76];
    endcase
  end

  // REG#726の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0726 <= imem07_in[47:44];
    74: reg_0726 <= imem07_in[47:44];
    78: reg_0726 <= imem07_in[47:44];
    endcase
  end

  // REG#727の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0727 <= imem07_in[127:124];
    74: reg_0727 <= imem07_in[127:124];
    78: reg_0727 <= imem07_in[127:124];
    endcase
  end

  // REG#728の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0728 <= imem07_in[7:4];
    74: reg_0728 <= imem07_in[7:4];
    78: reg_0728 <= imem07_in[7:4];
    endcase
  end

  // REG#729の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0729 <= imem07_in[79:76];
    74: reg_0729 <= imem07_in[79:76];
    77: reg_0729 <= imem07_in[79:76];
    79: reg_0729 <= imem07_in[79:76];
    endcase
  end

  // REG#730の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0730 <= imem07_in[27:24];
    77: reg_0730 <= imem07_in[27:24];
    81: reg_0730 <= imem07_in[27:24];
    endcase
  end

  // REG#731の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0731 <= imem07_in[35:32];
    74: reg_0731 <= imem07_in[35:32];
    78: reg_0731 <= imem07_in[119:116];
    endcase
  end

  // REG#732の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0732 <= imem03_in[7:4];
    7: reg_0732 <= op1_14_out;
    9: reg_0732 <= op1_14_out;
    11: reg_0732 <= imem05_in[103:100];
    19: reg_0732 <= imem05_in[103:100];
    49: reg_0732 <= imem05_in[103:100];
    63: reg_0732 <= op1_14_out;
    67: reg_0732 <= imem05_in[103:100];
    69: reg_0732 <= op1_14_out;
    72: reg_0732 <= imem05_in[103:100];
    endcase
  end

  // REG#733の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0733 <= imem03_in[95:92];
    8: reg_0733 <= imem01_in[23:20];
    11: reg_0733 <= imem05_in[71:68];
    19: reg_0733 <= imem05_in[71:68];
    48: reg_0733 <= imem01_in[23:20];
    69: reg_0733 <= imem03_in[95:92];
    endcase
  end

  // REG#734の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0734 <= imem05_in[115:112];
    8: reg_0734 <= imem01_in[95:92];
    11: reg_0734 <= imem05_in[115:112];
    19: reg_0734 <= imem05_in[115:112];
    48: reg_0734 <= imem01_in[95:92];
    67: reg_0734 <= imem01_in[95:92];
    73: reg_0734 <= imem05_in[115:112];
    endcase
  end

  // REG#735の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0735 <= imem03_in[27:24];
    8: reg_0735 <= imem01_in[119:116];
    11: reg_0735 <= imem05_in[47:44];
    19: reg_0735 <= imem05_in[47:44];
    48: reg_0735 <= imem01_in[7:4];
    68: reg_0735 <= imem03_in[27:24];
    71: reg_0735 <= imem05_in[47:44];
    78: reg_0735 <= imem05_in[47:44];
    85: reg_0735 <= imem05_in[47:44];
    endcase
  end

  // REG#736の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0736 <= imem05_in[15:12];
    8: reg_0736 <= imem01_in[35:32];
    11: reg_0736 <= imem05_in[15:12];
    19: reg_0736 <= imem05_in[15:12];
    46: reg_0736 <= imem01_in[35:32];
    49: reg_0736 <= imem05_in[15:12];
    67: reg_0736 <= imem05_in[15:12];
    72: reg_0736 <= imem05_in[15:12];
    endcase
  end

  // REG#737の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0737 <= imem05_in[55:52];
    8: reg_0737 <= imem01_in[111:108];
    11: reg_0737 <= imem05_in[35:32];
    19: reg_0737 <= imem05_in[35:32];
    48: reg_0737 <= imem01_in[111:108];
    68: reg_0737 <= imem01_in[111:108];
    endcase
  end

  // REG#738の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0738 <= imem03_in[3:0];
    8: reg_0738 <= imem01_in[3:0];
    10: reg_0738 <= op2_00_out;
    23: reg_0738 <= op2_00_out;
    24: reg_0738 <= op2_00_out;
    27: reg_0738 <= op2_00_out;
    38: reg_0738 <= op2_00_out;
    75: reg_0738 <= op2_00_out;
    endcase
  end

  // REG#739の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0739 <= imem03_in[119:116];
    8: reg_0739 <= imem01_in[7:4];
    10: reg_0739 <= op2_02_out;
    25: reg_0739 <= op2_02_out;
    33: reg_0739 <= op2_02_out;
    62: reg_0739 <= imem02_in[31:28];
    71: reg_0739 <= imem02_in[31:28];
    83: reg_0739 <= op2_02_out;
    endcase
  end

  // REG#740の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0740 <= imem03_in[83:80];
    8: reg_0740 <= imem01_in[123:120];
    20: reg_0740 <= imem02_in[111:108];
    84: reg_0740 <= imem02_in[111:108];
    endcase
  end

  // REG#741の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0741 <= imem05_in[19:16];
    8: reg_0741 <= imem01_in[39:36];
    19: reg_0741 <= imem05_in[19:16];
    48: reg_0741 <= imem01_in[39:36];
    68: reg_0741 <= imem01_in[39:36];
    91: reg_0741 <= imem01_in[39:36];
    endcase
  end

  // REG#742の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0742 <= imem05_in[43:40];
    8: reg_0742 <= imem01_in[51:48];
    19: reg_0742 <= imem05_in[43:40];
    49: reg_0742 <= imem05_in[43:40];
    64: reg_0742 <= imem05_in[43:40];
    67: reg_0742 <= imem05_in[43:40];
    73: reg_0742 <= imem05_in[43:40];
    endcase
  end

  // REG#743の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0743 <= imem05_in[87:84];
    8: reg_0743 <= imem01_in[67:64];
    20: reg_0743 <= imem02_in[19:16];
    84: reg_0743 <= imem02_in[19:16];
    endcase
  end

  // REG#744の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0744 <= imem05_in[111:108];
    8: reg_0744 <= imem01_in[83:80];
    11: reg_0744 <= imem05_in[111:108];
    19: reg_0744 <= imem05_in[111:108];
    49: reg_0744 <= imem05_in[111:108];
    54: reg_0744 <= imem00_in[63:60];
    90: reg_0744 <= imem00_in[63:60];
    endcase
  end

  // REG#745の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0745 <= imem03_in[11:8];
    7: reg_0745 <= op2_00_out;
    13: reg_0745 <= op2_00_out;
    33: reg_0745 <= op2_00_out;
    59: reg_0745 <= op2_00_out;
    endcase
  end

  // REG#746の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0746 <= imem03_in[103:100];
    7: reg_0746 <= op2_02_out;
    15: reg_0746 <= op2_02_out;
    42: reg_0746 <= op2_02_out;
    47: reg_0746 <= op2_02_out;
    64: reg_0746 <= op2_02_out;
    77: reg_0746 <= op2_02_out;
    endcase
  end

  // REG#747の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0747 <= imem05_in[123:120];
    8: reg_0747 <= imem06_in[27:24];
    27: reg_0747 <= imem03_in[107:104];
    69: reg_0747 <= imem03_in[107:104];
    endcase
  end

  // REG#748の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0748 <= imem03_in[35:32];
    8: reg_0748 <= imem06_in[75:72];
    28: reg_0748 <= imem06_in[75:72];
    57: reg_0748 <= imem06_in[75:72];
    85: reg_0748 <= imem06_in[75:72];
    endcase
  end

  // REG#749の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0749 <= imem05_in[7:4];
    8: reg_0749 <= imem06_in[115:112];
    30: reg_0749 <= imem03_in[127:124];
    54: reg_0749 <= imem00_in[67:64];
    90: reg_0749 <= imem00_in[67:64];
    endcase
  end

  // REG#750の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0750 <= imem05_in[27:24];
    8: reg_0750 <= imem06_in[87:84];
    30: reg_0750 <= imem03_in[67:64];
    54: reg_0750 <= imem03_in[67:64];
    85: reg_0750 <= imem06_in[87:84];
    endcase
  end

  // REG#751の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0751 <= imem05_in[71:68];
    8: reg_0751 <= imem06_in[107:104];
    30: reg_0751 <= imem03_in[119:116];
    54: reg_0751 <= imem03_in[119:116];
    86: reg_0751 <= imem05_in[71:68];
    endcase
  end

  // REG#752の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0752 <= imem05_in[103:100];
    8: reg_0752 <= imem06_in[99:96];
    30: reg_0752 <= imem06_in[99:96];
    36: reg_0752 <= imem06_in[99:96];
    55: reg_0752 <= imem05_in[103:100];
    60: reg_0752 <= imem06_in[99:96];
    70: reg_0752 <= imem06_in[99:96];
    endcase
  end

  // REG#753の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0753 <= op1_00_out;
    8: reg_0753 <= imem06_in[19:16];
    30: reg_0753 <= imem06_in[19:16];
    34: reg_0753 <= imem06_in[19:16];
    36: reg_0753 <= imem06_in[19:16];
    59: reg_0753 <= imem06_in[19:16];
    62: reg_0753 <= imem02_in[75:72];
    71: reg_0753 <= imem02_in[75:72];
    83: reg_0753 <= imem02_in[75:72];
    endcase
  end

  // REG#754の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0754 <= op1_01_out;
    9: reg_0754 <= op2_02_out;
    21: reg_0754 <= op2_02_out;
    62: reg_0754 <= op2_02_out;
    69: reg_0754 <= op1_01_out;
    70: reg_0754 <= op1_01_out;
    71: reg_0754 <= op1_01_out;
    72: reg_0754 <= op1_01_out;
    73: reg_0754 <= op1_01_out;
    74: reg_0754 <= op1_01_out;
    75: reg_0754 <= op1_01_out;
    76: reg_0754 <= op1_01_out;
    77: reg_0754 <= op1_01_out;
    78: reg_0754 <= op1_01_out;
    79: reg_0754 <= op1_01_out;
    80: reg_0754 <= op1_01_out;
    81: reg_0754 <= op1_01_out;
    82: reg_0754 <= op1_01_out;
    83: reg_0754 <= op1_01_out;
    85: reg_0754 <= op1_01_out;
    86: reg_0754 <= op1_01_out;
    87: reg_0754 <= op1_01_out;
    89: reg_0754 <= op2_02_out;
    endcase
  end

  // REG#755の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0755 <= op1_02_out;
    10: reg_0755 <= imem01_in[115:112];
    23: reg_0755 <= imem01_in[115:112];
    27: reg_0755 <= imem03_in[35:32];
    69: reg_0755 <= imem03_in[35:32];
    92: reg_0755 <= imem01_in[115:112];
    endcase
  end

  // REG#756の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0756 <= op1_03_out;
    20: reg_0756 <= imem02_in[75:72];
    84: reg_0756 <= imem02_in[75:72];
    endcase
  end

  // REG#757の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0757 <= op1_04_out;
    20: reg_0757 <= imem02_in[91:88];
    84: reg_0757 <= imem02_in[91:88];
    endcase
  end

  // REG#758の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0758 <= op1_05_out;
    12: reg_0758 <= op1_05_out;
    13: reg_0758 <= op1_05_out;
    14: reg_0758 <= op1_05_out;
    15: reg_0758 <= op1_05_out;
    16: reg_0758 <= op1_05_out;
    17: reg_0758 <= op1_05_out;
    18: reg_0758 <= op1_05_out;
    19: reg_0758 <= op1_05_out;
    24: reg_0758 <= imem01_in[3:0];
    46: reg_0758 <= imem01_in[3:0];
    54: reg_0758 <= imem00_in[83:80];
    90: reg_0758 <= imem00_in[83:80];
    endcase
  end

  // REG#759の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0759 <= op1_06_out;
    13: reg_0759 <= op1_06_out;
    14: reg_0759 <= op1_06_out;
    15: reg_0759 <= op1_06_out;
    16: reg_0759 <= op1_06_out;
    17: reg_0759 <= op1_06_out;
    18: reg_0759 <= op1_06_out;
    19: reg_0759 <= op1_06_out;
    24: reg_0759 <= imem01_in[83:80];
    48: reg_0759 <= imem01_in[83:80];
    68: reg_0759 <= imem01_in[83:80];
    endcase
  end

  // REG#760の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0760 <= op1_07_out;
    14: reg_0760 <= op1_07_out;
    15: reg_0760 <= op1_07_out;
    16: reg_0760 <= op1_07_out;
    17: reg_0760 <= op1_07_out;
    18: reg_0760 <= op1_07_out;
    19: reg_0760 <= op1_07_out;
    20: reg_0760 <= op1_07_out;
    21: reg_0760 <= op1_07_out;
    24: reg_0760 <= imem01_in[123:120];
    48: reg_0760 <= imem01_in[123:120];
    68: reg_0760 <= imem01_in[123:120];
    94: reg_0760 <= imem01_in[123:120];
    endcase
  end

  // REG#761の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0761 <= op1_08_out;
    16: reg_0761 <= op1_08_out;
    17: reg_0761 <= op1_08_out;
    18: reg_0761 <= op1_08_out;
    19: reg_0761 <= op1_08_out;
    20: reg_0761 <= op1_08_out;
    21: reg_0761 <= op1_08_out;
    24: reg_0761 <= imem01_in[111:108];
    48: reg_0761 <= imem01_in[55:52];
    73: reg_0761 <= imem05_in[91:88];
    91: reg_0761 <= imem01_in[55:52];
    endcase
  end

  // REG#762の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0762 <= op1_09_out;
    17: reg_0762 <= op1_09_out;
    18: reg_0762 <= op1_09_out;
    19: reg_0762 <= op1_09_out;
    20: reg_0762 <= op1_09_out;
    21: reg_0762 <= op1_09_out;
    22: reg_0762 <= op1_09_out;
    23: reg_0762 <= op1_09_out;
    24: reg_0762 <= op1_09_out;
    28: reg_0762 <= imem06_in[43:40];
    56: reg_0762 <= imem06_in[43:40];
    endcase
  end

  // REG#763の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0763 <= op1_10_out;
    18: reg_0763 <= op1_10_out;
    19: reg_0763 <= op1_10_out;
    20: reg_0763 <= op1_10_out;
    21: reg_0763 <= op1_10_out;
    22: reg_0763 <= op1_10_out;
    23: reg_0763 <= op1_10_out;
    24: reg_0763 <= op1_10_out;
    28: reg_0763 <= imem06_in[79:76];
    57: reg_0763 <= imem06_in[79:76];
    85: reg_0763 <= imem06_in[79:76];
    endcase
  end

  // REG#764の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0764 <= op1_11_out;
    21: reg_0764 <= op1_11_out;
    22: reg_0764 <= op1_11_out;
    23: reg_0764 <= op1_11_out;
    24: reg_0764 <= op1_11_out;
    25: reg_0764 <= op1_11_out;
    28: reg_0764 <= imem06_in[115:112];
    57: reg_0764 <= imem06_in[115:112];
    84: reg_0764 <= imem06_in[115:112];
    86: reg_0764 <= op1_11_out;
    88: reg_0764 <= imem06_in[115:112];
    endcase
  end

  // REG#765の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0765 <= op1_12_out;
    27: reg_0765 <= op1_12_out;
    28: reg_0765 <= op1_12_out;
    29: reg_0765 <= op1_12_out;
    30: reg_0765 <= op1_12_out;
    35: reg_0765 <= op1_12_out;
    42: reg_0765 <= op1_12_out;
    48: reg_0765 <= imem01_in[59:56];
    69: reg_0765 <= op1_12_out;
    73: reg_0765 <= imem05_in[95:92];
    endcase
  end

  // REG#766の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0766 <= op1_13_out;
    27: reg_0766 <= op1_13_out;
    31: reg_0766 <= imem06_in[103:100];
    38: reg_0766 <= imem06_in[103:100];
    56: reg_0766 <= imem06_in[103:100];
    endcase
  end

  // REG#767の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0767 <= op1_14_out;
    30: reg_0767 <= op1_14_out;
    41: reg_0767 <= op1_14_out;
    45: reg_0767 <= op1_14_out;
    48: reg_0767 <= op1_14_out;
    54: reg_0767 <= op1_14_out;
    56: reg_0767 <= op1_14_out;
    58: reg_0767 <= op1_14_out;
    60: reg_0767 <= imem06_in[91:88];
    70: reg_0767 <= imem06_in[91:88];
    87: reg_0767 <= op1_14_out;
    endcase
  end

  // REG#768の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0768 <= op1_15_out;
    30: reg_0768 <= op1_15_out;
    44: reg_0768 <= op1_15_out;
    47: reg_0768 <= op1_15_out;
    49: reg_0768 <= op1_15_out;
    51: reg_0768 <= op1_15_out;
    53: reg_0768 <= op1_15_out;
    55: reg_0768 <= op1_15_out;
    57: reg_0768 <= op1_15_out;
    59: reg_0768 <= op1_15_out;
    61: reg_0768 <= op1_15_out;
    63: reg_0768 <= op1_15_out;
    65: reg_0768 <= op1_15_out;
    67: reg_0768 <= op1_15_out;
    69: reg_0768 <= op1_15_out;
    71: reg_0768 <= op1_15_out;
    77: reg_0768 <= op1_15_out;
    79: reg_0768 <= op1_15_out;
    81: reg_0768 <= op1_15_out;
    83: reg_0768 <= op1_15_out;
    85: reg_0768 <= op1_15_out;
    87: reg_0768 <= op1_15_out;
    89: reg_0768 <= op1_15_out;
    91: reg_0768 <= op1_15_out;
    93: reg_0768 <= op1_15_out;
    endcase
  end

  // REG#769の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0769 <= op1_05_out;
    5: reg_0769 <= op1_05_out;
    6: reg_0769 <= op1_05_out;
    7: reg_0769 <= op1_05_out;
    8: reg_0769 <= op1_05_out;
    9: reg_0769 <= op1_05_out;
    10: reg_0769 <= op1_05_out;
    11: reg_0769 <= op1_05_out;
    20: reg_0769 <= imem02_in[51:48];
    endcase
  end

  // REG#770の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0770 <= op1_06_out;
    5: reg_0770 <= op1_06_out;
    6: reg_0770 <= op1_06_out;
    7: reg_0770 <= op1_06_out;
    8: reg_0770 <= op1_06_out;
    9: reg_0770 <= op1_06_out;
    10: reg_0770 <= op1_06_out;
    11: reg_0770 <= op1_06_out;
    12: reg_0770 <= op1_06_out;
    20: reg_0770 <= imem02_in[63:60];
    84: reg_0770 <= imem02_in[63:60];
    endcase
  end

  // REG#771の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0771 <= op1_07_out;
    5: reg_0771 <= op1_07_out;
    6: reg_0771 <= op1_07_out;
    7: reg_0771 <= op1_07_out;
    8: reg_0771 <= op1_07_out;
    9: reg_0771 <= op1_07_out;
    10: reg_0771 <= op1_07_out;
    11: reg_0771 <= op1_07_out;
    12: reg_0771 <= op1_07_out;
    13: reg_0771 <= op1_07_out;
    24: reg_0771 <= imem01_in[91:88];
    51: reg_0771 <= imem01_in[91:88];
    58: reg_0771 <= imem04_in[83:80];
    endcase
  end

  // REG#772の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0772 <= op1_08_out;
    5: reg_0772 <= op1_08_out;
    6: reg_0772 <= op1_08_out;
    7: reg_0772 <= op1_08_out;
    8: reg_0772 <= op1_08_out;
    9: reg_0772 <= op1_08_out;
    10: reg_0772 <= op1_08_out;
    11: reg_0772 <= op1_08_out;
    12: reg_0772 <= op1_08_out;
    13: reg_0772 <= op1_08_out;
    14: reg_0772 <= op1_08_out;
    15: reg_0772 <= op1_08_out;
    24: reg_0772 <= imem01_in[31:28];
    48: reg_0772 <= imem01_in[31:28];
    68: reg_0772 <= imem01_in[31:28];
    endcase
  end

  // REG#773の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0773 <= op1_09_out;
    5: reg_0773 <= op1_09_out;
    6: reg_0773 <= op1_09_out;
    7: reg_0773 <= op1_09_out;
    8: reg_0773 <= op1_09_out;
    9: reg_0773 <= op1_09_out;
    10: reg_0773 <= op1_09_out;
    11: reg_0773 <= op1_09_out;
    12: reg_0773 <= op1_09_out;
    13: reg_0773 <= op1_09_out;
    14: reg_0773 <= op1_09_out;
    15: reg_0773 <= op1_09_out;
    16: reg_0773 <= op1_09_out;
    28: reg_0773 <= imem06_in[67:64];
    57: reg_0773 <= imem06_in[67:64];
    84: reg_0773 <= imem06_in[67:64];
    endcase
  end

  // REG#774の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0774 <= op1_10_out;
    5: reg_0774 <= op1_10_out;
    6: reg_0774 <= op1_10_out;
    7: reg_0774 <= op1_10_out;
    8: reg_0774 <= op1_10_out;
    9: reg_0774 <= op1_10_out;
    10: reg_0774 <= op1_10_out;
    11: reg_0774 <= op1_10_out;
    12: reg_0774 <= op1_10_out;
    13: reg_0774 <= op1_10_out;
    14: reg_0774 <= op1_10_out;
    15: reg_0774 <= op1_10_out;
    16: reg_0774 <= op1_10_out;
    17: reg_0774 <= op1_10_out;
    28: reg_0774 <= imem06_in[7:4];
    58: reg_0774 <= imem04_in[79:76];
    endcase
  end

  // REG#775の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0775 <= op1_11_out;
    5: reg_0775 <= op1_11_out;
    6: reg_0775 <= op1_11_out;
    7: reg_0775 <= op1_11_out;
    8: reg_0775 <= op1_11_out;
    9: reg_0775 <= op1_11_out;
    10: reg_0775 <= op1_11_out;
    11: reg_0775 <= op1_11_out;
    12: reg_0775 <= op1_11_out;
    13: reg_0775 <= op1_11_out;
    14: reg_0775 <= op1_11_out;
    15: reg_0775 <= op1_11_out;
    16: reg_0775 <= op1_11_out;
    17: reg_0775 <= op1_11_out;
    18: reg_0775 <= op1_11_out;
    19: reg_0775 <= op1_11_out;
    20: reg_0775 <= op1_11_out;
    28: reg_0775 <= imem06_in[59:56];
    57: reg_0775 <= imem06_in[59:56];
    81: reg_0775 <= op1_11_out;
    85: reg_0775 <= imem06_in[59:56];
    endcase
  end

  // REG#776の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0776 <= op1_12_out;
    5: reg_0776 <= op1_12_out;
    6: reg_0776 <= op1_12_out;
    7: reg_0776 <= op1_12_out;
    10: reg_0776 <= imem01_in[99:96];
    28: reg_0776 <= imem06_in[91:88];
    58: reg_0776 <= imem04_in[99:96];
    endcase
  end

  // REG#777の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0777 <= op1_13_out;
    5: reg_0777 <= op1_13_out;
    6: reg_0777 <= op1_13_out;
    8: reg_0777 <= op1_13_out;
    9: reg_0777 <= op1_13_out;
    10: reg_0777 <= op1_13_out;
    13: reg_0777 <= op1_13_out;
    15: reg_0777 <= op1_13_out;
    16: reg_0777 <= op1_13_out;
    19: reg_0777 <= op1_13_out;
    21: reg_0777 <= op1_13_out;
    23: reg_0777 <= op1_13_out;
    24: reg_0777 <= op1_13_out;
    25: reg_0777 <= op1_13_out;
    26: reg_0777 <= op1_13_out;
    28: reg_0777 <= op1_13_out;
    31: reg_0777 <= imem06_in[39:36];
    36: reg_0777 <= imem06_in[39:36];
    60: reg_0777 <= imem06_in[39:36];
    70: reg_0777 <= imem06_in[39:36];
    88: reg_0777 <= imem06_in[39:36];
    endcase
  end

  // REG#778の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0778 <= op1_14_out;
    6: reg_0778 <= op1_14_out;
    10: reg_0778 <= imem01_in[87:84];
    23: reg_0778 <= imem01_in[87:84];
    25: reg_0778 <= op1_14_out;
    26: reg_0778 <= op1_14_out;
    31: reg_0778 <= imem06_in[35:32];
    36: reg_0778 <= imem06_in[35:32];
    48: reg_0778 <= imem01_in[87:84];
    68: reg_0778 <= imem01_in[87:84];
    93: reg_0778 <= imem01_in[87:84];
    endcase
  end

  // REG#779の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0779 <= op1_15_out;
    7: reg_0779 <= op1_15_out;
    9: reg_0779 <= op1_15_out;
    11: reg_0779 <= op1_15_out;
    13: reg_0779 <= op1_15_out;
    16: reg_0779 <= op1_15_out;
    18: reg_0779 <= op1_15_out;
    20: reg_0779 <= op1_15_out;
    23: reg_0779 <= op1_15_out;
    25: reg_0779 <= op1_15_out;
    27: reg_0779 <= op1_15_out;
    31: reg_0779 <= imem06_in[87:84];
    55: reg_0779 <= imem06_in[87:84];
    58: reg_0779 <= imem04_in[7:4];
    endcase
  end

  // REG#780の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0780 <= imem05_in[79:76];
    54: reg_0780 <= imem05_in[79:76];
    58: reg_0780 <= imem04_in[59:56];
    endcase
  end

  // REG#781の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0781 <= imem05_in[31:28];
    55: reg_0781 <= imem05_in[31:28];
    60: reg_0781 <= imem05_in[31:28];
    67: reg_0781 <= imem05_in[31:28];
    71: reg_0781 <= imem05_in[31:28];
    73: reg_0781 <= imem05_in[31:28];
    endcase
  end

  // REG#782の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0782 <= imem05_in[91:88];
    55: reg_0782 <= imem05_in[91:88];
    60: reg_0782 <= imem05_in[91:88];
    67: reg_0782 <= imem05_in[91:88];
    72: reg_0782 <= imem05_in[91:88];
    endcase
  end

  // REG#783の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0783 <= imem05_in[99:96];
    60: reg_0783 <= imem05_in[99:96];
    65: reg_0783 <= imem05_in[99:96];
    73: reg_0783 <= imem05_in[87:84];
    endcase
  end

  // REG#784の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0784 <= imem05_in[111:108];
    60: reg_0784 <= imem05_in[111:108];
    64: reg_0784 <= imem05_in[111:108];
    66: reg_0784 <= imem05_in[111:108];
    71: reg_0784 <= imem05_in[111:108];
    78: reg_0784 <= imem07_in[51:48];
    endcase
  end

  // REG#785の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0785 <= imem05_in[83:80];
    55: reg_0785 <= imem05_in[83:80];
    59: reg_0785 <= imem05_in[83:80];
    62: reg_0785 <= imem02_in[27:24];
    73: reg_0785 <= imem05_in[23:20];
    endcase
  end

  // REG#786の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0786 <= imem05_in[103:100];
    60: reg_0786 <= imem05_in[103:100];
    65: reg_0786 <= imem05_in[103:100];
    77: reg_0786 <= imem05_in[103:100];
    endcase
  end

  // REG#787の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0787 <= imem05_in[119:116];
    54: reg_0787 <= imem05_in[119:116];
    60: reg_0787 <= imem06_in[87:84];
    70: reg_0787 <= imem06_in[87:84];
    endcase
  end

  // REG#788の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0788 <= imem05_in[47:44];
    55: reg_0788 <= imem05_in[47:44];
    59: reg_0788 <= imem05_in[47:44];
    64: reg_0788 <= imem05_in[47:44];
    67: reg_0788 <= imem05_in[47:44];
    72: reg_0788 <= imem05_in[47:44];
    endcase
  end

  // REG#789の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0789 <= imem05_in[51:48];
    54: reg_0789 <= imem05_in[51:48];
    60: reg_0789 <= imem05_in[51:48];
    65: reg_0789 <= imem05_in[51:48];
    78: reg_0789 <= imem07_in[91:88];
    endcase
  end

  // REG#790の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0790 <= imem05_in[107:104];
    55: reg_0790 <= imem05_in[107:104];
    60: reg_0790 <= imem05_in[107:104];
    65: reg_0790 <= imem05_in[107:104];
    endcase
  end

  // REG#791の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0791 <= imem05_in[3:0];
    55: reg_0791 <= imem05_in[3:0];
    60: reg_0791 <= imem05_in[3:0];
    64: reg_0791 <= imem05_in[3:0];
    72: reg_0791 <= imem05_in[3:0];
    endcase
  end

  // REG#792の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0792 <= imem05_in[7:4];
    55: reg_0792 <= imem05_in[7:4];
    60: reg_0792 <= imem05_in[7:4];
    64: reg_0792 <= imem05_in[7:4];
    67: reg_0792 <= imem05_in[7:4];
    72: reg_0792 <= imem05_in[7:4];
    endcase
  end

  // REG#793の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0793 <= imem05_in[71:68];
    55: reg_0793 <= imem05_in[71:68];
    60: reg_0793 <= imem05_in[71:68];
    64: reg_0793 <= imem05_in[71:68];
    67: reg_0793 <= imem05_in[71:68];
    72: reg_0793 <= imem05_in[71:68];
    endcase
  end

  // REG#794の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0794 <= imem05_in[95:92];
    60: reg_0794 <= imem06_in[51:48];
    70: reg_0794 <= imem06_in[51:48];
    87: reg_0794 <= imem06_in[51:48];
    endcase
  end

  // REG#795の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0795 <= imem05_in[63:60];
    55: reg_0795 <= imem05_in[63:60];
    60: reg_0795 <= imem05_in[63:60];
    64: reg_0795 <= imem05_in[63:60];
    72: reg_0795 <= imem05_in[63:60];
    endcase
  end

  // REG#796の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0796 <= imem05_in[15:12];
    55: reg_0796 <= imem05_in[15:12];
    60: reg_0796 <= imem05_in[15:12];
    73: reg_0796 <= imem05_in[79:76];
    endcase
  end

  // REG#797の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0797 <= imem05_in[27:24];
    55: reg_0797 <= imem05_in[27:24];
    60: reg_0797 <= imem05_in[27:24];
    63: reg_0797 <= imem05_in[27:24];
    65: reg_0797 <= imem05_in[27:24];
    77: reg_0797 <= imem05_in[27:24];
    86: reg_0797 <= imem05_in[27:24];
    endcase
  end

  // REG#798の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0798 <= imem05_in[11:8];
    55: reg_0798 <= imem05_in[11:8];
    59: reg_0798 <= op2_02_out;
    endcase
  end

  // REG#799の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0799 <= imem03_in[87:84];
    87: reg_0799 <= imem03_in[87:84];
    endcase
  end

  // REG#800の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0800 <= imem03_in[63:60];
    89: reg_0800 <= imem03_in[63:60];
    endcase
  end

  // REG#801の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0801 <= imem03_in[59:56];
    87: reg_0801 <= imem03_in[59:56];
    endcase
  end

  // REG#802の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0802 <= imem03_in[79:76];
    89: reg_0802 <= imem03_in[79:76];
    endcase
  end

  // REG#803の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0803 <= imem03_in[39:36];
    88: reg_0803 <= imem03_in[39:36];
    endcase
  end

  // REG#804の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0804 <= imem03_in[55:52];
    endcase
  end

  // REG#805の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0805 <= imem03_in[71:68];
    88: reg_0805 <= imem03_in[71:68];
    endcase
  end

  // REG#806の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0806 <= imem03_in[95:92];
    89: reg_0806 <= imem03_in[95:92];
    endcase
  end

  // REG#807の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0807 <= imem03_in[51:48];
    89: reg_0807 <= imem03_in[51:48];
    endcase
  end

  // REG#808の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0808 <= imem03_in[31:28];
    endcase
  end

  // REG#809の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0809 <= imem03_in[111:108];
    89: reg_0809 <= imem03_in[111:108];
    endcase
  end

  // REG#810の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0810 <= imem03_in[99:96];
    endcase
  end

  // REG#811の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0811 <= imem03_in[15:12];
    89: reg_0811 <= imem03_in[15:12];
    endcase
  end

  // REG#812の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0812 <= imem06_in[23:20];
    31: reg_0812 <= imem06_in[23:20];
    34: reg_0812 <= imem06_in[23:20];
    36: reg_0812 <= imem06_in[23:20];
    60: reg_0812 <= imem06_in[23:20];
    69: reg_0812 <= imem06_in[23:20];
    73: reg_0812 <= imem05_in[3:0];
    endcase
  end

  // REG#813の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0813 <= imem06_in[31:28];
    30: reg_0813 <= imem06_in[31:28];
    34: reg_0813 <= imem06_in[31:28];
    60: reg_0813 <= imem06_in[31:28];
    70: reg_0813 <= imem06_in[31:28];
    88: reg_0813 <= imem06_in[31:28];
    endcase
  end

  // REG#814の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0814 <= imem06_in[67:64];
    31: reg_0814 <= imem06_in[3:0];
    36: reg_0814 <= imem06_in[67:64];
    56: reg_0814 <= imem06_in[67:64];
    endcase
  end

  // REG#815の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0815 <= imem06_in[47:44];
    30: reg_0815 <= imem06_in[47:44];
    36: reg_0815 <= imem06_in[47:44];
    56: reg_0815 <= imem06_in[47:44];
    endcase
  end

  // REG#816の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0816 <= imem06_in[63:60];
    31: reg_0816 <= imem06_in[47:44];
    57: reg_0816 <= imem06_in[63:60];
    84: reg_0816 <= imem06_in[63:60];
    87: reg_0816 <= imem06_in[47:44];
    endcase
  end

  // REG#817の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0817 <= imem06_in[55:52];
    31: reg_0817 <= imem06_in[55:52];
    38: reg_0817 <= imem06_in[55:52];
    56: reg_0817 <= imem06_in[55:52];
    endcase
  end

  // REG#818の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0818 <= imem06_in[83:80];
    31: reg_0818 <= imem06_in[83:80];
    36: reg_0818 <= imem06_in[83:80];
    59: reg_0818 <= imem06_in[83:80];
    70: reg_0818 <= imem06_in[83:80];
    endcase
  end

  // REG#819の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0819 <= imem06_in[59:56];
    31: reg_0819 <= imem06_in[59:56];
    36: reg_0819 <= imem06_in[59:56];
    60: reg_0819 <= imem06_in[59:56];
    70: reg_0819 <= imem06_in[59:56];
    88: reg_0819 <= imem06_in[59:56];
    endcase
  end

  // REG#820の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0820 <= imem01_in[51:48];
    24: reg_0820 <= imem01_in[51:48];
    48: reg_0820 <= imem01_in[51:48];
    68: reg_0820 <= imem01_in[51:48];
    91: reg_0820 <= imem01_in[51:48];
    endcase
  end

  // REG#821の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0821 <= imem01_in[123:120];
    23: reg_0821 <= imem01_in[123:120];
    28: reg_0821 <= imem06_in[71:68];
    57: reg_0821 <= imem06_in[71:68];
    endcase
  end

  // REG#822の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0822 <= imem01_in[39:36];
    24: reg_0822 <= imem01_in[39:36];
    73: reg_0822 <= imem05_in[27:24];
    endcase
  end

  // REG#823の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0823 <= op2_03_out;
    22: reg_0823 <= op2_03_out;
    24: reg_0823 <= op2_03_out;
    30: reg_0823 <= op2_00_out;
    50: reg_0823 <= op2_00_out;
    71: reg_0823 <= op2_00_out;
    endcase
  end

  // REG#824の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0824 <= imem01_in[59:56];
    24: reg_0824 <= imem01_in[59:56];
    46: reg_0824 <= imem01_in[59:56];
    51: reg_0824 <= imem01_in[59:56];
    73: reg_0824 <= imem05_in[111:108];
    endcase
  end

  // REG#825の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0825 <= imem01_in[79:76];
    24: reg_0825 <= imem01_in[79:76];
    48: reg_0825 <= imem01_in[79:76];
    67: reg_0825 <= imem01_in[79:76];
    73: reg_0825 <= imem05_in[51:48];
    endcase
  end

  // REG#826の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0826 <= op2_02_out;
    52: reg_0826 <= op2_02_out;
    86: reg_0826 <= op2_02_out;
    endcase
  end

  // REG#827の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_0827 <= imem05_in[19:16];
    endcase
  end

  // REG#828の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_0828 <= imem05_in[107:104];
    endcase
  end

  // REG#829の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_0829 <= imem05_in[71:68];
    endcase
  end

  // REG#830の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_0830 <= imem05_in[55:52];
    endcase
  end

  // REG#831の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_0831 <= op2_00_out;
    endcase
  end
endmodule
