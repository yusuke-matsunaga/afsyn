module affine2(
  input clock,
  input reset,
  input start,
  output busy,
  output [4:0] imem00_bank,
  output imem00_rd,
  input [15:0] imem00_in,
  output [4:0] imem01_bank,
  output imem01_rd,
  input [15:0] imem01_in,
  output [4:0] imem02_bank,
  output imem02_rd,
  input [15:0] imem02_in,
  output [4:0] imem03_bank,
  output imem03_rd,
  input [15:0] imem03_in,
  output [4:0] imem04_bank,
  output imem04_rd,
  input [15:0] imem04_in,
  output [4:0] imem05_bank,
  output imem05_rd,
  input [15:0] imem05_in,
  output [4:0] imem06_bank,
  output imem06_rd,
  input [15:0] imem06_in,
  output [4:0] imem07_bank,
  output imem07_rd,
  input [15:0] imem07_in,
  output [5:0] omem00_bank,
  output omem00_wr,
  output [8:0] omem00_out,
  output [5:0] omem01_bank,
  output omem01_wr,
  output [8:0] omem01_out,
  output [5:0] omem02_bank,
  output omem02_wr,
  output [8:0] omem02_out,
  output [5:0] omem03_bank,
  output omem03_wr,
  output [8:0] omem03_out,
  output [5:0] omem04_bank,
  output omem04_wr,
  output [8:0] omem04_out);


  // 0 番目の OP1
  reg [3:0] op1_00_in00;
  reg       op1_00_inv00;
  reg [3:0] op1_00_in01;
  reg       op1_00_inv01;
  reg [3:0] op1_00_in02;
  reg       op1_00_inv02;
  reg [3:0] op1_00_in03;
  reg       op1_00_inv03;
  reg [3:0] op1_00_in04;
  reg       op1_00_inv04;
  reg [3:0] op1_00_in05;
  reg       op1_00_inv05;
  reg [3:0] op1_00_in06;
  reg       op1_00_inv06;
  reg [3:0] op1_00_in07;
  reg       op1_00_inv07;
  reg [3:0] op1_00_in08;
  reg       op1_00_inv08;
  reg [3:0] op1_00_in09;
  reg       op1_00_inv09;
  reg [3:0] op1_00_in10;
  reg       op1_00_inv10;
  reg [3:0] op1_00_in11;
  reg       op1_00_inv11;
  reg [3:0] op1_00_in12;
  reg       op1_00_inv12;
  reg [3:0] op1_00_in13;
  reg       op1_00_inv13;
  reg [3:0] op1_00_in14;
  reg       op1_00_inv14;
  reg [3:0] op1_00_in15;
  reg       op1_00_inv15;
  reg [3:0] op1_00_in16;
  reg       op1_00_inv16;
  reg [3:0] op1_00_in17;
  reg       op1_00_inv17;
  reg [3:0] op1_00_in18;
  reg       op1_00_inv18;
  reg [3:0] op1_00_in19;
  reg       op1_00_inv19;
  reg [3:0] op1_00_in20;
  reg       op1_00_inv20;
  reg [3:0] op1_00_in21;
  reg       op1_00_inv21;
  reg [3:0] op1_00_in22;
  reg       op1_00_inv22;
  reg [3:0] op1_00_in23;
  reg       op1_00_inv23;
  reg [3:0] op1_00_in24;
  reg       op1_00_inv24;
  reg [3:0] op1_00_in25;
  reg       op1_00_inv25;
  reg [3:0] op1_00_in26;
  reg       op1_00_inv26;
  reg [3:0] op1_00_in27;
  reg       op1_00_inv27;
  reg [3:0] op1_00_in28;
  reg       op1_00_inv28;
  reg [3:0] op1_00_in29;
  reg       op1_00_inv29;
  reg [3:0] op1_00_in30;
  reg       op1_00_inv30;
  reg [3:0] op1_00_in31;
  reg       op1_00_inv31;
  wire [8:0] op1_00_out;
  affine2_op1 op1_00(
    .data0_in(op1_00_in00),
    .inv0_in(op1_00_inv00),
    .data1_in(op1_00_in01),
    .inv1_in(op1_00_inv01),
    .data2_in(op1_00_in02),
    .inv2_in(op1_00_inv02),
    .data3_in(op1_00_in03),
    .inv3_in(op1_00_inv03),
    .data4_in(op1_00_in04),
    .inv4_in(op1_00_inv04),
    .data5_in(op1_00_in05),
    .inv5_in(op1_00_inv05),
    .data6_in(op1_00_in06),
    .inv6_in(op1_00_inv06),
    .data7_in(op1_00_in07),
    .inv7_in(op1_00_inv07),
    .data8_in(op1_00_in08),
    .inv8_in(op1_00_inv08),
    .data9_in(op1_00_in09),
    .inv9_in(op1_00_inv09),
    .data10_in(op1_00_in10),
    .inv10_in(op1_00_inv10),
    .data11_in(op1_00_in11),
    .inv11_in(op1_00_inv11),
    .data12_in(op1_00_in12),
    .inv12_in(op1_00_inv12),
    .data13_in(op1_00_in13),
    .inv13_in(op1_00_inv13),
    .data14_in(op1_00_in14),
    .inv14_in(op1_00_inv14),
    .data15_in(op1_00_in15),
    .inv15_in(op1_00_inv15),
    .data16_in(op1_00_in16),
    .inv16_in(op1_00_inv16),
    .data17_in(op1_00_in17),
    .inv17_in(op1_00_inv17),
    .data18_in(op1_00_in18),
    .inv18_in(op1_00_inv18),
    .data19_in(op1_00_in19),
    .inv19_in(op1_00_inv19),
    .data20_in(op1_00_in20),
    .inv20_in(op1_00_inv20),
    .data21_in(op1_00_in21),
    .inv21_in(op1_00_inv21),
    .data22_in(op1_00_in22),
    .inv22_in(op1_00_inv22),
    .data23_in(op1_00_in23),
    .inv23_in(op1_00_inv23),
    .data24_in(op1_00_in24),
    .inv24_in(op1_00_inv24),
    .data25_in(op1_00_in25),
    .inv25_in(op1_00_inv25),
    .data26_in(op1_00_in26),
    .inv26_in(op1_00_inv26),
    .data27_in(op1_00_in27),
    .inv27_in(op1_00_inv27),
    .data28_in(op1_00_in28),
    .inv28_in(op1_00_inv28),
    .data29_in(op1_00_in29),
    .inv29_in(op1_00_inv29),
    .data30_in(op1_00_in30),
    .inv30_in(op1_00_inv30),
    .data31_in(op1_00_in31),
    .inv31_in(op1_00_inv31),
    .data_out(op1_00_out));

  // 1 番目の OP1
  reg [3:0] op1_01_in00;
  reg       op1_01_inv00;
  reg [3:0] op1_01_in01;
  reg       op1_01_inv01;
  reg [3:0] op1_01_in02;
  reg       op1_01_inv02;
  reg [3:0] op1_01_in03;
  reg       op1_01_inv03;
  reg [3:0] op1_01_in04;
  reg       op1_01_inv04;
  reg [3:0] op1_01_in05;
  reg       op1_01_inv05;
  reg [3:0] op1_01_in06;
  reg       op1_01_inv06;
  reg [3:0] op1_01_in07;
  reg       op1_01_inv07;
  reg [3:0] op1_01_in08;
  reg       op1_01_inv08;
  reg [3:0] op1_01_in09;
  reg       op1_01_inv09;
  reg [3:0] op1_01_in10;
  reg       op1_01_inv10;
  reg [3:0] op1_01_in11;
  reg       op1_01_inv11;
  reg [3:0] op1_01_in12;
  reg       op1_01_inv12;
  reg [3:0] op1_01_in13;
  reg       op1_01_inv13;
  reg [3:0] op1_01_in14;
  reg       op1_01_inv14;
  reg [3:0] op1_01_in15;
  reg       op1_01_inv15;
  reg [3:0] op1_01_in16;
  reg       op1_01_inv16;
  reg [3:0] op1_01_in17;
  reg       op1_01_inv17;
  reg [3:0] op1_01_in18;
  reg       op1_01_inv18;
  reg [3:0] op1_01_in19;
  reg       op1_01_inv19;
  reg [3:0] op1_01_in20;
  reg       op1_01_inv20;
  reg [3:0] op1_01_in21;
  reg       op1_01_inv21;
  reg [3:0] op1_01_in22;
  reg       op1_01_inv22;
  reg [3:0] op1_01_in23;
  reg       op1_01_inv23;
  reg [3:0] op1_01_in24;
  reg       op1_01_inv24;
  reg [3:0] op1_01_in25;
  reg       op1_01_inv25;
  reg [3:0] op1_01_in26;
  reg       op1_01_inv26;
  reg [3:0] op1_01_in27;
  reg       op1_01_inv27;
  reg [3:0] op1_01_in28;
  reg       op1_01_inv28;
  reg [3:0] op1_01_in29;
  reg       op1_01_inv29;
  reg [3:0] op1_01_in30;
  reg       op1_01_inv30;
  reg [3:0] op1_01_in31;
  reg       op1_01_inv31;
  wire [8:0] op1_01_out;
  affine2_op1 op1_01(
    .data0_in(op1_01_in00),
    .inv0_in(op1_01_inv00),
    .data1_in(op1_01_in01),
    .inv1_in(op1_01_inv01),
    .data2_in(op1_01_in02),
    .inv2_in(op1_01_inv02),
    .data3_in(op1_01_in03),
    .inv3_in(op1_01_inv03),
    .data4_in(op1_01_in04),
    .inv4_in(op1_01_inv04),
    .data5_in(op1_01_in05),
    .inv5_in(op1_01_inv05),
    .data6_in(op1_01_in06),
    .inv6_in(op1_01_inv06),
    .data7_in(op1_01_in07),
    .inv7_in(op1_01_inv07),
    .data8_in(op1_01_in08),
    .inv8_in(op1_01_inv08),
    .data9_in(op1_01_in09),
    .inv9_in(op1_01_inv09),
    .data10_in(op1_01_in10),
    .inv10_in(op1_01_inv10),
    .data11_in(op1_01_in11),
    .inv11_in(op1_01_inv11),
    .data12_in(op1_01_in12),
    .inv12_in(op1_01_inv12),
    .data13_in(op1_01_in13),
    .inv13_in(op1_01_inv13),
    .data14_in(op1_01_in14),
    .inv14_in(op1_01_inv14),
    .data15_in(op1_01_in15),
    .inv15_in(op1_01_inv15),
    .data16_in(op1_01_in16),
    .inv16_in(op1_01_inv16),
    .data17_in(op1_01_in17),
    .inv17_in(op1_01_inv17),
    .data18_in(op1_01_in18),
    .inv18_in(op1_01_inv18),
    .data19_in(op1_01_in19),
    .inv19_in(op1_01_inv19),
    .data20_in(op1_01_in20),
    .inv20_in(op1_01_inv20),
    .data21_in(op1_01_in21),
    .inv21_in(op1_01_inv21),
    .data22_in(op1_01_in22),
    .inv22_in(op1_01_inv22),
    .data23_in(op1_01_in23),
    .inv23_in(op1_01_inv23),
    .data24_in(op1_01_in24),
    .inv24_in(op1_01_inv24),
    .data25_in(op1_01_in25),
    .inv25_in(op1_01_inv25),
    .data26_in(op1_01_in26),
    .inv26_in(op1_01_inv26),
    .data27_in(op1_01_in27),
    .inv27_in(op1_01_inv27),
    .data28_in(op1_01_in28),
    .inv28_in(op1_01_inv28),
    .data29_in(op1_01_in29),
    .inv29_in(op1_01_inv29),
    .data30_in(op1_01_in30),
    .inv30_in(op1_01_inv30),
    .data31_in(op1_01_in31),
    .inv31_in(op1_01_inv31),
    .data_out(op1_01_out));

  // 2 番目の OP1
  reg [3:0] op1_02_in00;
  reg       op1_02_inv00;
  reg [3:0] op1_02_in01;
  reg       op1_02_inv01;
  reg [3:0] op1_02_in02;
  reg       op1_02_inv02;
  reg [3:0] op1_02_in03;
  reg       op1_02_inv03;
  reg [3:0] op1_02_in04;
  reg       op1_02_inv04;
  reg [3:0] op1_02_in05;
  reg       op1_02_inv05;
  reg [3:0] op1_02_in06;
  reg       op1_02_inv06;
  reg [3:0] op1_02_in07;
  reg       op1_02_inv07;
  reg [3:0] op1_02_in08;
  reg       op1_02_inv08;
  reg [3:0] op1_02_in09;
  reg       op1_02_inv09;
  reg [3:0] op1_02_in10;
  reg       op1_02_inv10;
  reg [3:0] op1_02_in11;
  reg       op1_02_inv11;
  reg [3:0] op1_02_in12;
  reg       op1_02_inv12;
  reg [3:0] op1_02_in13;
  reg       op1_02_inv13;
  reg [3:0] op1_02_in14;
  reg       op1_02_inv14;
  reg [3:0] op1_02_in15;
  reg       op1_02_inv15;
  reg [3:0] op1_02_in16;
  reg       op1_02_inv16;
  reg [3:0] op1_02_in17;
  reg       op1_02_inv17;
  reg [3:0] op1_02_in18;
  reg       op1_02_inv18;
  reg [3:0] op1_02_in19;
  reg       op1_02_inv19;
  reg [3:0] op1_02_in20;
  reg       op1_02_inv20;
  reg [3:0] op1_02_in21;
  reg       op1_02_inv21;
  reg [3:0] op1_02_in22;
  reg       op1_02_inv22;
  reg [3:0] op1_02_in23;
  reg       op1_02_inv23;
  reg [3:0] op1_02_in24;
  reg       op1_02_inv24;
  reg [3:0] op1_02_in25;
  reg       op1_02_inv25;
  reg [3:0] op1_02_in26;
  reg       op1_02_inv26;
  reg [3:0] op1_02_in27;
  reg       op1_02_inv27;
  reg [3:0] op1_02_in28;
  reg       op1_02_inv28;
  reg [3:0] op1_02_in29;
  reg       op1_02_inv29;
  reg [3:0] op1_02_in30;
  reg       op1_02_inv30;
  reg [3:0] op1_02_in31;
  reg       op1_02_inv31;
  wire [8:0] op1_02_out;
  affine2_op1 op1_02(
    .data0_in(op1_02_in00),
    .inv0_in(op1_02_inv00),
    .data1_in(op1_02_in01),
    .inv1_in(op1_02_inv01),
    .data2_in(op1_02_in02),
    .inv2_in(op1_02_inv02),
    .data3_in(op1_02_in03),
    .inv3_in(op1_02_inv03),
    .data4_in(op1_02_in04),
    .inv4_in(op1_02_inv04),
    .data5_in(op1_02_in05),
    .inv5_in(op1_02_inv05),
    .data6_in(op1_02_in06),
    .inv6_in(op1_02_inv06),
    .data7_in(op1_02_in07),
    .inv7_in(op1_02_inv07),
    .data8_in(op1_02_in08),
    .inv8_in(op1_02_inv08),
    .data9_in(op1_02_in09),
    .inv9_in(op1_02_inv09),
    .data10_in(op1_02_in10),
    .inv10_in(op1_02_inv10),
    .data11_in(op1_02_in11),
    .inv11_in(op1_02_inv11),
    .data12_in(op1_02_in12),
    .inv12_in(op1_02_inv12),
    .data13_in(op1_02_in13),
    .inv13_in(op1_02_inv13),
    .data14_in(op1_02_in14),
    .inv14_in(op1_02_inv14),
    .data15_in(op1_02_in15),
    .inv15_in(op1_02_inv15),
    .data16_in(op1_02_in16),
    .inv16_in(op1_02_inv16),
    .data17_in(op1_02_in17),
    .inv17_in(op1_02_inv17),
    .data18_in(op1_02_in18),
    .inv18_in(op1_02_inv18),
    .data19_in(op1_02_in19),
    .inv19_in(op1_02_inv19),
    .data20_in(op1_02_in20),
    .inv20_in(op1_02_inv20),
    .data21_in(op1_02_in21),
    .inv21_in(op1_02_inv21),
    .data22_in(op1_02_in22),
    .inv22_in(op1_02_inv22),
    .data23_in(op1_02_in23),
    .inv23_in(op1_02_inv23),
    .data24_in(op1_02_in24),
    .inv24_in(op1_02_inv24),
    .data25_in(op1_02_in25),
    .inv25_in(op1_02_inv25),
    .data26_in(op1_02_in26),
    .inv26_in(op1_02_inv26),
    .data27_in(op1_02_in27),
    .inv27_in(op1_02_inv27),
    .data28_in(op1_02_in28),
    .inv28_in(op1_02_inv28),
    .data29_in(op1_02_in29),
    .inv29_in(op1_02_inv29),
    .data30_in(op1_02_in30),
    .inv30_in(op1_02_inv30),
    .data31_in(op1_02_in31),
    .inv31_in(op1_02_inv31),
    .data_out(op1_02_out));

  // 3 番目の OP1
  reg [3:0] op1_03_in00;
  reg       op1_03_inv00;
  reg [3:0] op1_03_in01;
  reg       op1_03_inv01;
  reg [3:0] op1_03_in02;
  reg       op1_03_inv02;
  reg [3:0] op1_03_in03;
  reg       op1_03_inv03;
  reg [3:0] op1_03_in04;
  reg       op1_03_inv04;
  reg [3:0] op1_03_in05;
  reg       op1_03_inv05;
  reg [3:0] op1_03_in06;
  reg       op1_03_inv06;
  reg [3:0] op1_03_in07;
  reg       op1_03_inv07;
  reg [3:0] op1_03_in08;
  reg       op1_03_inv08;
  reg [3:0] op1_03_in09;
  reg       op1_03_inv09;
  reg [3:0] op1_03_in10;
  reg       op1_03_inv10;
  reg [3:0] op1_03_in11;
  reg       op1_03_inv11;
  reg [3:0] op1_03_in12;
  reg       op1_03_inv12;
  reg [3:0] op1_03_in13;
  reg       op1_03_inv13;
  reg [3:0] op1_03_in14;
  reg       op1_03_inv14;
  reg [3:0] op1_03_in15;
  reg       op1_03_inv15;
  reg [3:0] op1_03_in16;
  reg       op1_03_inv16;
  reg [3:0] op1_03_in17;
  reg       op1_03_inv17;
  reg [3:0] op1_03_in18;
  reg       op1_03_inv18;
  reg [3:0] op1_03_in19;
  reg       op1_03_inv19;
  reg [3:0] op1_03_in20;
  reg       op1_03_inv20;
  reg [3:0] op1_03_in21;
  reg       op1_03_inv21;
  reg [3:0] op1_03_in22;
  reg       op1_03_inv22;
  reg [3:0] op1_03_in23;
  reg       op1_03_inv23;
  reg [3:0] op1_03_in24;
  reg       op1_03_inv24;
  reg [3:0] op1_03_in25;
  reg       op1_03_inv25;
  reg [3:0] op1_03_in26;
  reg       op1_03_inv26;
  reg [3:0] op1_03_in27;
  reg       op1_03_inv27;
  reg [3:0] op1_03_in28;
  reg       op1_03_inv28;
  reg [3:0] op1_03_in29;
  reg       op1_03_inv29;
  reg [3:0] op1_03_in30;
  reg       op1_03_inv30;
  reg [3:0] op1_03_in31;
  reg       op1_03_inv31;
  wire [8:0] op1_03_out;
  affine2_op1 op1_03(
    .data0_in(op1_03_in00),
    .inv0_in(op1_03_inv00),
    .data1_in(op1_03_in01),
    .inv1_in(op1_03_inv01),
    .data2_in(op1_03_in02),
    .inv2_in(op1_03_inv02),
    .data3_in(op1_03_in03),
    .inv3_in(op1_03_inv03),
    .data4_in(op1_03_in04),
    .inv4_in(op1_03_inv04),
    .data5_in(op1_03_in05),
    .inv5_in(op1_03_inv05),
    .data6_in(op1_03_in06),
    .inv6_in(op1_03_inv06),
    .data7_in(op1_03_in07),
    .inv7_in(op1_03_inv07),
    .data8_in(op1_03_in08),
    .inv8_in(op1_03_inv08),
    .data9_in(op1_03_in09),
    .inv9_in(op1_03_inv09),
    .data10_in(op1_03_in10),
    .inv10_in(op1_03_inv10),
    .data11_in(op1_03_in11),
    .inv11_in(op1_03_inv11),
    .data12_in(op1_03_in12),
    .inv12_in(op1_03_inv12),
    .data13_in(op1_03_in13),
    .inv13_in(op1_03_inv13),
    .data14_in(op1_03_in14),
    .inv14_in(op1_03_inv14),
    .data15_in(op1_03_in15),
    .inv15_in(op1_03_inv15),
    .data16_in(op1_03_in16),
    .inv16_in(op1_03_inv16),
    .data17_in(op1_03_in17),
    .inv17_in(op1_03_inv17),
    .data18_in(op1_03_in18),
    .inv18_in(op1_03_inv18),
    .data19_in(op1_03_in19),
    .inv19_in(op1_03_inv19),
    .data20_in(op1_03_in20),
    .inv20_in(op1_03_inv20),
    .data21_in(op1_03_in21),
    .inv21_in(op1_03_inv21),
    .data22_in(op1_03_in22),
    .inv22_in(op1_03_inv22),
    .data23_in(op1_03_in23),
    .inv23_in(op1_03_inv23),
    .data24_in(op1_03_in24),
    .inv24_in(op1_03_inv24),
    .data25_in(op1_03_in25),
    .inv25_in(op1_03_inv25),
    .data26_in(op1_03_in26),
    .inv26_in(op1_03_inv26),
    .data27_in(op1_03_in27),
    .inv27_in(op1_03_inv27),
    .data28_in(op1_03_in28),
    .inv28_in(op1_03_inv28),
    .data29_in(op1_03_in29),
    .inv29_in(op1_03_inv29),
    .data30_in(op1_03_in30),
    .inv30_in(op1_03_inv30),
    .data31_in(op1_03_in31),
    .inv31_in(op1_03_inv31),
    .data_out(op1_03_out));

  // 4 番目の OP1
  reg [3:0] op1_04_in00;
  reg       op1_04_inv00;
  reg [3:0] op1_04_in01;
  reg       op1_04_inv01;
  reg [3:0] op1_04_in02;
  reg       op1_04_inv02;
  reg [3:0] op1_04_in03;
  reg       op1_04_inv03;
  reg [3:0] op1_04_in04;
  reg       op1_04_inv04;
  reg [3:0] op1_04_in05;
  reg       op1_04_inv05;
  reg [3:0] op1_04_in06;
  reg       op1_04_inv06;
  reg [3:0] op1_04_in07;
  reg       op1_04_inv07;
  reg [3:0] op1_04_in08;
  reg       op1_04_inv08;
  reg [3:0] op1_04_in09;
  reg       op1_04_inv09;
  reg [3:0] op1_04_in10;
  reg       op1_04_inv10;
  reg [3:0] op1_04_in11;
  reg       op1_04_inv11;
  reg [3:0] op1_04_in12;
  reg       op1_04_inv12;
  reg [3:0] op1_04_in13;
  reg       op1_04_inv13;
  reg [3:0] op1_04_in14;
  reg       op1_04_inv14;
  reg [3:0] op1_04_in15;
  reg       op1_04_inv15;
  reg [3:0] op1_04_in16;
  reg       op1_04_inv16;
  reg [3:0] op1_04_in17;
  reg       op1_04_inv17;
  reg [3:0] op1_04_in18;
  reg       op1_04_inv18;
  reg [3:0] op1_04_in19;
  reg       op1_04_inv19;
  reg [3:0] op1_04_in20;
  reg       op1_04_inv20;
  reg [3:0] op1_04_in21;
  reg       op1_04_inv21;
  reg [3:0] op1_04_in22;
  reg       op1_04_inv22;
  reg [3:0] op1_04_in23;
  reg       op1_04_inv23;
  reg [3:0] op1_04_in24;
  reg       op1_04_inv24;
  reg [3:0] op1_04_in25;
  reg       op1_04_inv25;
  reg [3:0] op1_04_in26;
  reg       op1_04_inv26;
  reg [3:0] op1_04_in27;
  reg       op1_04_inv27;
  reg [3:0] op1_04_in28;
  reg       op1_04_inv28;
  reg [3:0] op1_04_in29;
  reg       op1_04_inv29;
  reg [3:0] op1_04_in30;
  reg       op1_04_inv30;
  reg [3:0] op1_04_in31;
  reg       op1_04_inv31;
  wire [8:0] op1_04_out;
  affine2_op1 op1_04(
    .data0_in(op1_04_in00),
    .inv0_in(op1_04_inv00),
    .data1_in(op1_04_in01),
    .inv1_in(op1_04_inv01),
    .data2_in(op1_04_in02),
    .inv2_in(op1_04_inv02),
    .data3_in(op1_04_in03),
    .inv3_in(op1_04_inv03),
    .data4_in(op1_04_in04),
    .inv4_in(op1_04_inv04),
    .data5_in(op1_04_in05),
    .inv5_in(op1_04_inv05),
    .data6_in(op1_04_in06),
    .inv6_in(op1_04_inv06),
    .data7_in(op1_04_in07),
    .inv7_in(op1_04_inv07),
    .data8_in(op1_04_in08),
    .inv8_in(op1_04_inv08),
    .data9_in(op1_04_in09),
    .inv9_in(op1_04_inv09),
    .data10_in(op1_04_in10),
    .inv10_in(op1_04_inv10),
    .data11_in(op1_04_in11),
    .inv11_in(op1_04_inv11),
    .data12_in(op1_04_in12),
    .inv12_in(op1_04_inv12),
    .data13_in(op1_04_in13),
    .inv13_in(op1_04_inv13),
    .data14_in(op1_04_in14),
    .inv14_in(op1_04_inv14),
    .data15_in(op1_04_in15),
    .inv15_in(op1_04_inv15),
    .data16_in(op1_04_in16),
    .inv16_in(op1_04_inv16),
    .data17_in(op1_04_in17),
    .inv17_in(op1_04_inv17),
    .data18_in(op1_04_in18),
    .inv18_in(op1_04_inv18),
    .data19_in(op1_04_in19),
    .inv19_in(op1_04_inv19),
    .data20_in(op1_04_in20),
    .inv20_in(op1_04_inv20),
    .data21_in(op1_04_in21),
    .inv21_in(op1_04_inv21),
    .data22_in(op1_04_in22),
    .inv22_in(op1_04_inv22),
    .data23_in(op1_04_in23),
    .inv23_in(op1_04_inv23),
    .data24_in(op1_04_in24),
    .inv24_in(op1_04_inv24),
    .data25_in(op1_04_in25),
    .inv25_in(op1_04_inv25),
    .data26_in(op1_04_in26),
    .inv26_in(op1_04_inv26),
    .data27_in(op1_04_in27),
    .inv27_in(op1_04_inv27),
    .data28_in(op1_04_in28),
    .inv28_in(op1_04_inv28),
    .data29_in(op1_04_in29),
    .inv29_in(op1_04_inv29),
    .data30_in(op1_04_in30),
    .inv30_in(op1_04_inv30),
    .data31_in(op1_04_in31),
    .inv31_in(op1_04_inv31),
    .data_out(op1_04_out));

  // 5 番目の OP1
  reg [3:0] op1_05_in00;
  reg       op1_05_inv00;
  reg [3:0] op1_05_in01;
  reg       op1_05_inv01;
  reg [3:0] op1_05_in02;
  reg       op1_05_inv02;
  reg [3:0] op1_05_in03;
  reg       op1_05_inv03;
  reg [3:0] op1_05_in04;
  reg       op1_05_inv04;
  reg [3:0] op1_05_in05;
  reg       op1_05_inv05;
  reg [3:0] op1_05_in06;
  reg       op1_05_inv06;
  reg [3:0] op1_05_in07;
  reg       op1_05_inv07;
  reg [3:0] op1_05_in08;
  reg       op1_05_inv08;
  reg [3:0] op1_05_in09;
  reg       op1_05_inv09;
  reg [3:0] op1_05_in10;
  reg       op1_05_inv10;
  reg [3:0] op1_05_in11;
  reg       op1_05_inv11;
  reg [3:0] op1_05_in12;
  reg       op1_05_inv12;
  reg [3:0] op1_05_in13;
  reg       op1_05_inv13;
  reg [3:0] op1_05_in14;
  reg       op1_05_inv14;
  reg [3:0] op1_05_in15;
  reg       op1_05_inv15;
  reg [3:0] op1_05_in16;
  reg       op1_05_inv16;
  reg [3:0] op1_05_in17;
  reg       op1_05_inv17;
  reg [3:0] op1_05_in18;
  reg       op1_05_inv18;
  reg [3:0] op1_05_in19;
  reg       op1_05_inv19;
  reg [3:0] op1_05_in20;
  reg       op1_05_inv20;
  reg [3:0] op1_05_in21;
  reg       op1_05_inv21;
  reg [3:0] op1_05_in22;
  reg       op1_05_inv22;
  reg [3:0] op1_05_in23;
  reg       op1_05_inv23;
  reg [3:0] op1_05_in24;
  reg       op1_05_inv24;
  reg [3:0] op1_05_in25;
  reg       op1_05_inv25;
  reg [3:0] op1_05_in26;
  reg       op1_05_inv26;
  reg [3:0] op1_05_in27;
  reg       op1_05_inv27;
  reg [3:0] op1_05_in28;
  reg       op1_05_inv28;
  reg [3:0] op1_05_in29;
  reg       op1_05_inv29;
  reg [3:0] op1_05_in30;
  reg       op1_05_inv30;
  reg [3:0] op1_05_in31;
  reg       op1_05_inv31;
  wire [8:0] op1_05_out;
  affine2_op1 op1_05(
    .data0_in(op1_05_in00),
    .inv0_in(op1_05_inv00),
    .data1_in(op1_05_in01),
    .inv1_in(op1_05_inv01),
    .data2_in(op1_05_in02),
    .inv2_in(op1_05_inv02),
    .data3_in(op1_05_in03),
    .inv3_in(op1_05_inv03),
    .data4_in(op1_05_in04),
    .inv4_in(op1_05_inv04),
    .data5_in(op1_05_in05),
    .inv5_in(op1_05_inv05),
    .data6_in(op1_05_in06),
    .inv6_in(op1_05_inv06),
    .data7_in(op1_05_in07),
    .inv7_in(op1_05_inv07),
    .data8_in(op1_05_in08),
    .inv8_in(op1_05_inv08),
    .data9_in(op1_05_in09),
    .inv9_in(op1_05_inv09),
    .data10_in(op1_05_in10),
    .inv10_in(op1_05_inv10),
    .data11_in(op1_05_in11),
    .inv11_in(op1_05_inv11),
    .data12_in(op1_05_in12),
    .inv12_in(op1_05_inv12),
    .data13_in(op1_05_in13),
    .inv13_in(op1_05_inv13),
    .data14_in(op1_05_in14),
    .inv14_in(op1_05_inv14),
    .data15_in(op1_05_in15),
    .inv15_in(op1_05_inv15),
    .data16_in(op1_05_in16),
    .inv16_in(op1_05_inv16),
    .data17_in(op1_05_in17),
    .inv17_in(op1_05_inv17),
    .data18_in(op1_05_in18),
    .inv18_in(op1_05_inv18),
    .data19_in(op1_05_in19),
    .inv19_in(op1_05_inv19),
    .data20_in(op1_05_in20),
    .inv20_in(op1_05_inv20),
    .data21_in(op1_05_in21),
    .inv21_in(op1_05_inv21),
    .data22_in(op1_05_in22),
    .inv22_in(op1_05_inv22),
    .data23_in(op1_05_in23),
    .inv23_in(op1_05_inv23),
    .data24_in(op1_05_in24),
    .inv24_in(op1_05_inv24),
    .data25_in(op1_05_in25),
    .inv25_in(op1_05_inv25),
    .data26_in(op1_05_in26),
    .inv26_in(op1_05_inv26),
    .data27_in(op1_05_in27),
    .inv27_in(op1_05_inv27),
    .data28_in(op1_05_in28),
    .inv28_in(op1_05_inv28),
    .data29_in(op1_05_in29),
    .inv29_in(op1_05_inv29),
    .data30_in(op1_05_in30),
    .inv30_in(op1_05_inv30),
    .data31_in(op1_05_in31),
    .inv31_in(op1_05_inv31),
    .data_out(op1_05_out));

  // 6 番目の OP1
  reg [3:0] op1_06_in00;
  reg       op1_06_inv00;
  reg [3:0] op1_06_in01;
  reg       op1_06_inv01;
  reg [3:0] op1_06_in02;
  reg       op1_06_inv02;
  reg [3:0] op1_06_in03;
  reg       op1_06_inv03;
  reg [3:0] op1_06_in04;
  reg       op1_06_inv04;
  reg [3:0] op1_06_in05;
  reg       op1_06_inv05;
  reg [3:0] op1_06_in06;
  reg       op1_06_inv06;
  reg [3:0] op1_06_in07;
  reg       op1_06_inv07;
  reg [3:0] op1_06_in08;
  reg       op1_06_inv08;
  reg [3:0] op1_06_in09;
  reg       op1_06_inv09;
  reg [3:0] op1_06_in10;
  reg       op1_06_inv10;
  reg [3:0] op1_06_in11;
  reg       op1_06_inv11;
  reg [3:0] op1_06_in12;
  reg       op1_06_inv12;
  reg [3:0] op1_06_in13;
  reg       op1_06_inv13;
  reg [3:0] op1_06_in14;
  reg       op1_06_inv14;
  reg [3:0] op1_06_in15;
  reg       op1_06_inv15;
  reg [3:0] op1_06_in16;
  reg       op1_06_inv16;
  reg [3:0] op1_06_in17;
  reg       op1_06_inv17;
  reg [3:0] op1_06_in18;
  reg       op1_06_inv18;
  reg [3:0] op1_06_in19;
  reg       op1_06_inv19;
  reg [3:0] op1_06_in20;
  reg       op1_06_inv20;
  reg [3:0] op1_06_in21;
  reg       op1_06_inv21;
  reg [3:0] op1_06_in22;
  reg       op1_06_inv22;
  reg [3:0] op1_06_in23;
  reg       op1_06_inv23;
  reg [3:0] op1_06_in24;
  reg       op1_06_inv24;
  reg [3:0] op1_06_in25;
  reg       op1_06_inv25;
  reg [3:0] op1_06_in26;
  reg       op1_06_inv26;
  reg [3:0] op1_06_in27;
  reg       op1_06_inv27;
  reg [3:0] op1_06_in28;
  reg       op1_06_inv28;
  reg [3:0] op1_06_in29;
  reg       op1_06_inv29;
  reg [3:0] op1_06_in30;
  reg       op1_06_inv30;
  reg [3:0] op1_06_in31;
  reg       op1_06_inv31;
  wire [8:0] op1_06_out;
  affine2_op1 op1_06(
    .data0_in(op1_06_in00),
    .inv0_in(op1_06_inv00),
    .data1_in(op1_06_in01),
    .inv1_in(op1_06_inv01),
    .data2_in(op1_06_in02),
    .inv2_in(op1_06_inv02),
    .data3_in(op1_06_in03),
    .inv3_in(op1_06_inv03),
    .data4_in(op1_06_in04),
    .inv4_in(op1_06_inv04),
    .data5_in(op1_06_in05),
    .inv5_in(op1_06_inv05),
    .data6_in(op1_06_in06),
    .inv6_in(op1_06_inv06),
    .data7_in(op1_06_in07),
    .inv7_in(op1_06_inv07),
    .data8_in(op1_06_in08),
    .inv8_in(op1_06_inv08),
    .data9_in(op1_06_in09),
    .inv9_in(op1_06_inv09),
    .data10_in(op1_06_in10),
    .inv10_in(op1_06_inv10),
    .data11_in(op1_06_in11),
    .inv11_in(op1_06_inv11),
    .data12_in(op1_06_in12),
    .inv12_in(op1_06_inv12),
    .data13_in(op1_06_in13),
    .inv13_in(op1_06_inv13),
    .data14_in(op1_06_in14),
    .inv14_in(op1_06_inv14),
    .data15_in(op1_06_in15),
    .inv15_in(op1_06_inv15),
    .data16_in(op1_06_in16),
    .inv16_in(op1_06_inv16),
    .data17_in(op1_06_in17),
    .inv17_in(op1_06_inv17),
    .data18_in(op1_06_in18),
    .inv18_in(op1_06_inv18),
    .data19_in(op1_06_in19),
    .inv19_in(op1_06_inv19),
    .data20_in(op1_06_in20),
    .inv20_in(op1_06_inv20),
    .data21_in(op1_06_in21),
    .inv21_in(op1_06_inv21),
    .data22_in(op1_06_in22),
    .inv22_in(op1_06_inv22),
    .data23_in(op1_06_in23),
    .inv23_in(op1_06_inv23),
    .data24_in(op1_06_in24),
    .inv24_in(op1_06_inv24),
    .data25_in(op1_06_in25),
    .inv25_in(op1_06_inv25),
    .data26_in(op1_06_in26),
    .inv26_in(op1_06_inv26),
    .data27_in(op1_06_in27),
    .inv27_in(op1_06_inv27),
    .data28_in(op1_06_in28),
    .inv28_in(op1_06_inv28),
    .data29_in(op1_06_in29),
    .inv29_in(op1_06_inv29),
    .data30_in(op1_06_in30),
    .inv30_in(op1_06_inv30),
    .data31_in(op1_06_in31),
    .inv31_in(op1_06_inv31),
    .data_out(op1_06_out));

  // 7 番目の OP1
  reg [3:0] op1_07_in00;
  reg       op1_07_inv00;
  reg [3:0] op1_07_in01;
  reg       op1_07_inv01;
  reg [3:0] op1_07_in02;
  reg       op1_07_inv02;
  reg [3:0] op1_07_in03;
  reg       op1_07_inv03;
  reg [3:0] op1_07_in04;
  reg       op1_07_inv04;
  reg [3:0] op1_07_in05;
  reg       op1_07_inv05;
  reg [3:0] op1_07_in06;
  reg       op1_07_inv06;
  reg [3:0] op1_07_in07;
  reg       op1_07_inv07;
  reg [3:0] op1_07_in08;
  reg       op1_07_inv08;
  reg [3:0] op1_07_in09;
  reg       op1_07_inv09;
  reg [3:0] op1_07_in10;
  reg       op1_07_inv10;
  reg [3:0] op1_07_in11;
  reg       op1_07_inv11;
  reg [3:0] op1_07_in12;
  reg       op1_07_inv12;
  reg [3:0] op1_07_in13;
  reg       op1_07_inv13;
  reg [3:0] op1_07_in14;
  reg       op1_07_inv14;
  reg [3:0] op1_07_in15;
  reg       op1_07_inv15;
  reg [3:0] op1_07_in16;
  reg       op1_07_inv16;
  reg [3:0] op1_07_in17;
  reg       op1_07_inv17;
  reg [3:0] op1_07_in18;
  reg       op1_07_inv18;
  reg [3:0] op1_07_in19;
  reg       op1_07_inv19;
  reg [3:0] op1_07_in20;
  reg       op1_07_inv20;
  reg [3:0] op1_07_in21;
  reg       op1_07_inv21;
  reg [3:0] op1_07_in22;
  reg       op1_07_inv22;
  reg [3:0] op1_07_in23;
  reg       op1_07_inv23;
  reg [3:0] op1_07_in24;
  reg       op1_07_inv24;
  reg [3:0] op1_07_in25;
  reg       op1_07_inv25;
  reg [3:0] op1_07_in26;
  reg       op1_07_inv26;
  reg [3:0] op1_07_in27;
  reg       op1_07_inv27;
  reg [3:0] op1_07_in28;
  reg       op1_07_inv28;
  reg [3:0] op1_07_in29;
  reg       op1_07_inv29;
  reg [3:0] op1_07_in30;
  reg       op1_07_inv30;
  reg [3:0] op1_07_in31;
  reg       op1_07_inv31;
  wire [8:0] op1_07_out;
  affine2_op1 op1_07(
    .data0_in(op1_07_in00),
    .inv0_in(op1_07_inv00),
    .data1_in(op1_07_in01),
    .inv1_in(op1_07_inv01),
    .data2_in(op1_07_in02),
    .inv2_in(op1_07_inv02),
    .data3_in(op1_07_in03),
    .inv3_in(op1_07_inv03),
    .data4_in(op1_07_in04),
    .inv4_in(op1_07_inv04),
    .data5_in(op1_07_in05),
    .inv5_in(op1_07_inv05),
    .data6_in(op1_07_in06),
    .inv6_in(op1_07_inv06),
    .data7_in(op1_07_in07),
    .inv7_in(op1_07_inv07),
    .data8_in(op1_07_in08),
    .inv8_in(op1_07_inv08),
    .data9_in(op1_07_in09),
    .inv9_in(op1_07_inv09),
    .data10_in(op1_07_in10),
    .inv10_in(op1_07_inv10),
    .data11_in(op1_07_in11),
    .inv11_in(op1_07_inv11),
    .data12_in(op1_07_in12),
    .inv12_in(op1_07_inv12),
    .data13_in(op1_07_in13),
    .inv13_in(op1_07_inv13),
    .data14_in(op1_07_in14),
    .inv14_in(op1_07_inv14),
    .data15_in(op1_07_in15),
    .inv15_in(op1_07_inv15),
    .data16_in(op1_07_in16),
    .inv16_in(op1_07_inv16),
    .data17_in(op1_07_in17),
    .inv17_in(op1_07_inv17),
    .data18_in(op1_07_in18),
    .inv18_in(op1_07_inv18),
    .data19_in(op1_07_in19),
    .inv19_in(op1_07_inv19),
    .data20_in(op1_07_in20),
    .inv20_in(op1_07_inv20),
    .data21_in(op1_07_in21),
    .inv21_in(op1_07_inv21),
    .data22_in(op1_07_in22),
    .inv22_in(op1_07_inv22),
    .data23_in(op1_07_in23),
    .inv23_in(op1_07_inv23),
    .data24_in(op1_07_in24),
    .inv24_in(op1_07_inv24),
    .data25_in(op1_07_in25),
    .inv25_in(op1_07_inv25),
    .data26_in(op1_07_in26),
    .inv26_in(op1_07_inv26),
    .data27_in(op1_07_in27),
    .inv27_in(op1_07_inv27),
    .data28_in(op1_07_in28),
    .inv28_in(op1_07_inv28),
    .data29_in(op1_07_in29),
    .inv29_in(op1_07_inv29),
    .data30_in(op1_07_in30),
    .inv30_in(op1_07_inv30),
    .data31_in(op1_07_in31),
    .inv31_in(op1_07_inv31),
    .data_out(op1_07_out));

  // 8 番目の OP1
  reg [3:0] op1_08_in00;
  reg       op1_08_inv00;
  reg [3:0] op1_08_in01;
  reg       op1_08_inv01;
  reg [3:0] op1_08_in02;
  reg       op1_08_inv02;
  reg [3:0] op1_08_in03;
  reg       op1_08_inv03;
  reg [3:0] op1_08_in04;
  reg       op1_08_inv04;
  reg [3:0] op1_08_in05;
  reg       op1_08_inv05;
  reg [3:0] op1_08_in06;
  reg       op1_08_inv06;
  reg [3:0] op1_08_in07;
  reg       op1_08_inv07;
  reg [3:0] op1_08_in08;
  reg       op1_08_inv08;
  reg [3:0] op1_08_in09;
  reg       op1_08_inv09;
  reg [3:0] op1_08_in10;
  reg       op1_08_inv10;
  reg [3:0] op1_08_in11;
  reg       op1_08_inv11;
  reg [3:0] op1_08_in12;
  reg       op1_08_inv12;
  reg [3:0] op1_08_in13;
  reg       op1_08_inv13;
  reg [3:0] op1_08_in14;
  reg       op1_08_inv14;
  reg [3:0] op1_08_in15;
  reg       op1_08_inv15;
  reg [3:0] op1_08_in16;
  reg       op1_08_inv16;
  reg [3:0] op1_08_in17;
  reg       op1_08_inv17;
  reg [3:0] op1_08_in18;
  reg       op1_08_inv18;
  reg [3:0] op1_08_in19;
  reg       op1_08_inv19;
  reg [3:0] op1_08_in20;
  reg       op1_08_inv20;
  reg [3:0] op1_08_in21;
  reg       op1_08_inv21;
  reg [3:0] op1_08_in22;
  reg       op1_08_inv22;
  reg [3:0] op1_08_in23;
  reg       op1_08_inv23;
  reg [3:0] op1_08_in24;
  reg       op1_08_inv24;
  reg [3:0] op1_08_in25;
  reg       op1_08_inv25;
  reg [3:0] op1_08_in26;
  reg       op1_08_inv26;
  reg [3:0] op1_08_in27;
  reg       op1_08_inv27;
  reg [3:0] op1_08_in28;
  reg       op1_08_inv28;
  reg [3:0] op1_08_in29;
  reg       op1_08_inv29;
  reg [3:0] op1_08_in30;
  reg       op1_08_inv30;
  reg [3:0] op1_08_in31;
  reg       op1_08_inv31;
  wire [8:0] op1_08_out;
  affine2_op1 op1_08(
    .data0_in(op1_08_in00),
    .inv0_in(op1_08_inv00),
    .data1_in(op1_08_in01),
    .inv1_in(op1_08_inv01),
    .data2_in(op1_08_in02),
    .inv2_in(op1_08_inv02),
    .data3_in(op1_08_in03),
    .inv3_in(op1_08_inv03),
    .data4_in(op1_08_in04),
    .inv4_in(op1_08_inv04),
    .data5_in(op1_08_in05),
    .inv5_in(op1_08_inv05),
    .data6_in(op1_08_in06),
    .inv6_in(op1_08_inv06),
    .data7_in(op1_08_in07),
    .inv7_in(op1_08_inv07),
    .data8_in(op1_08_in08),
    .inv8_in(op1_08_inv08),
    .data9_in(op1_08_in09),
    .inv9_in(op1_08_inv09),
    .data10_in(op1_08_in10),
    .inv10_in(op1_08_inv10),
    .data11_in(op1_08_in11),
    .inv11_in(op1_08_inv11),
    .data12_in(op1_08_in12),
    .inv12_in(op1_08_inv12),
    .data13_in(op1_08_in13),
    .inv13_in(op1_08_inv13),
    .data14_in(op1_08_in14),
    .inv14_in(op1_08_inv14),
    .data15_in(op1_08_in15),
    .inv15_in(op1_08_inv15),
    .data16_in(op1_08_in16),
    .inv16_in(op1_08_inv16),
    .data17_in(op1_08_in17),
    .inv17_in(op1_08_inv17),
    .data18_in(op1_08_in18),
    .inv18_in(op1_08_inv18),
    .data19_in(op1_08_in19),
    .inv19_in(op1_08_inv19),
    .data20_in(op1_08_in20),
    .inv20_in(op1_08_inv20),
    .data21_in(op1_08_in21),
    .inv21_in(op1_08_inv21),
    .data22_in(op1_08_in22),
    .inv22_in(op1_08_inv22),
    .data23_in(op1_08_in23),
    .inv23_in(op1_08_inv23),
    .data24_in(op1_08_in24),
    .inv24_in(op1_08_inv24),
    .data25_in(op1_08_in25),
    .inv25_in(op1_08_inv25),
    .data26_in(op1_08_in26),
    .inv26_in(op1_08_inv26),
    .data27_in(op1_08_in27),
    .inv27_in(op1_08_inv27),
    .data28_in(op1_08_in28),
    .inv28_in(op1_08_inv28),
    .data29_in(op1_08_in29),
    .inv29_in(op1_08_inv29),
    .data30_in(op1_08_in30),
    .inv30_in(op1_08_inv30),
    .data31_in(op1_08_in31),
    .inv31_in(op1_08_inv31),
    .data_out(op1_08_out));

  // 9 番目の OP1
  reg [3:0] op1_09_in00;
  reg       op1_09_inv00;
  reg [3:0] op1_09_in01;
  reg       op1_09_inv01;
  reg [3:0] op1_09_in02;
  reg       op1_09_inv02;
  reg [3:0] op1_09_in03;
  reg       op1_09_inv03;
  reg [3:0] op1_09_in04;
  reg       op1_09_inv04;
  reg [3:0] op1_09_in05;
  reg       op1_09_inv05;
  reg [3:0] op1_09_in06;
  reg       op1_09_inv06;
  reg [3:0] op1_09_in07;
  reg       op1_09_inv07;
  reg [3:0] op1_09_in08;
  reg       op1_09_inv08;
  reg [3:0] op1_09_in09;
  reg       op1_09_inv09;
  reg [3:0] op1_09_in10;
  reg       op1_09_inv10;
  reg [3:0] op1_09_in11;
  reg       op1_09_inv11;
  reg [3:0] op1_09_in12;
  reg       op1_09_inv12;
  reg [3:0] op1_09_in13;
  reg       op1_09_inv13;
  reg [3:0] op1_09_in14;
  reg       op1_09_inv14;
  reg [3:0] op1_09_in15;
  reg       op1_09_inv15;
  reg [3:0] op1_09_in16;
  reg       op1_09_inv16;
  reg [3:0] op1_09_in17;
  reg       op1_09_inv17;
  reg [3:0] op1_09_in18;
  reg       op1_09_inv18;
  reg [3:0] op1_09_in19;
  reg       op1_09_inv19;
  reg [3:0] op1_09_in20;
  reg       op1_09_inv20;
  reg [3:0] op1_09_in21;
  reg       op1_09_inv21;
  reg [3:0] op1_09_in22;
  reg       op1_09_inv22;
  reg [3:0] op1_09_in23;
  reg       op1_09_inv23;
  reg [3:0] op1_09_in24;
  reg       op1_09_inv24;
  reg [3:0] op1_09_in25;
  reg       op1_09_inv25;
  reg [3:0] op1_09_in26;
  reg       op1_09_inv26;
  reg [3:0] op1_09_in27;
  reg       op1_09_inv27;
  reg [3:0] op1_09_in28;
  reg       op1_09_inv28;
  reg [3:0] op1_09_in29;
  reg       op1_09_inv29;
  reg [3:0] op1_09_in30;
  reg       op1_09_inv30;
  reg [3:0] op1_09_in31;
  reg       op1_09_inv31;
  wire [8:0] op1_09_out;
  affine2_op1 op1_09(
    .data0_in(op1_09_in00),
    .inv0_in(op1_09_inv00),
    .data1_in(op1_09_in01),
    .inv1_in(op1_09_inv01),
    .data2_in(op1_09_in02),
    .inv2_in(op1_09_inv02),
    .data3_in(op1_09_in03),
    .inv3_in(op1_09_inv03),
    .data4_in(op1_09_in04),
    .inv4_in(op1_09_inv04),
    .data5_in(op1_09_in05),
    .inv5_in(op1_09_inv05),
    .data6_in(op1_09_in06),
    .inv6_in(op1_09_inv06),
    .data7_in(op1_09_in07),
    .inv7_in(op1_09_inv07),
    .data8_in(op1_09_in08),
    .inv8_in(op1_09_inv08),
    .data9_in(op1_09_in09),
    .inv9_in(op1_09_inv09),
    .data10_in(op1_09_in10),
    .inv10_in(op1_09_inv10),
    .data11_in(op1_09_in11),
    .inv11_in(op1_09_inv11),
    .data12_in(op1_09_in12),
    .inv12_in(op1_09_inv12),
    .data13_in(op1_09_in13),
    .inv13_in(op1_09_inv13),
    .data14_in(op1_09_in14),
    .inv14_in(op1_09_inv14),
    .data15_in(op1_09_in15),
    .inv15_in(op1_09_inv15),
    .data16_in(op1_09_in16),
    .inv16_in(op1_09_inv16),
    .data17_in(op1_09_in17),
    .inv17_in(op1_09_inv17),
    .data18_in(op1_09_in18),
    .inv18_in(op1_09_inv18),
    .data19_in(op1_09_in19),
    .inv19_in(op1_09_inv19),
    .data20_in(op1_09_in20),
    .inv20_in(op1_09_inv20),
    .data21_in(op1_09_in21),
    .inv21_in(op1_09_inv21),
    .data22_in(op1_09_in22),
    .inv22_in(op1_09_inv22),
    .data23_in(op1_09_in23),
    .inv23_in(op1_09_inv23),
    .data24_in(op1_09_in24),
    .inv24_in(op1_09_inv24),
    .data25_in(op1_09_in25),
    .inv25_in(op1_09_inv25),
    .data26_in(op1_09_in26),
    .inv26_in(op1_09_inv26),
    .data27_in(op1_09_in27),
    .inv27_in(op1_09_inv27),
    .data28_in(op1_09_in28),
    .inv28_in(op1_09_inv28),
    .data29_in(op1_09_in29),
    .inv29_in(op1_09_inv29),
    .data30_in(op1_09_in30),
    .inv30_in(op1_09_inv30),
    .data31_in(op1_09_in31),
    .inv31_in(op1_09_inv31),
    .data_out(op1_09_out));

  // 10 番目の OP1
  reg [3:0] op1_10_in00;
  reg       op1_10_inv00;
  reg [3:0] op1_10_in01;
  reg       op1_10_inv01;
  reg [3:0] op1_10_in02;
  reg       op1_10_inv02;
  reg [3:0] op1_10_in03;
  reg       op1_10_inv03;
  reg [3:0] op1_10_in04;
  reg       op1_10_inv04;
  reg [3:0] op1_10_in05;
  reg       op1_10_inv05;
  reg [3:0] op1_10_in06;
  reg       op1_10_inv06;
  reg [3:0] op1_10_in07;
  reg       op1_10_inv07;
  reg [3:0] op1_10_in08;
  reg       op1_10_inv08;
  reg [3:0] op1_10_in09;
  reg       op1_10_inv09;
  reg [3:0] op1_10_in10;
  reg       op1_10_inv10;
  reg [3:0] op1_10_in11;
  reg       op1_10_inv11;
  reg [3:0] op1_10_in12;
  reg       op1_10_inv12;
  reg [3:0] op1_10_in13;
  reg       op1_10_inv13;
  reg [3:0] op1_10_in14;
  reg       op1_10_inv14;
  reg [3:0] op1_10_in15;
  reg       op1_10_inv15;
  reg [3:0] op1_10_in16;
  reg       op1_10_inv16;
  reg [3:0] op1_10_in17;
  reg       op1_10_inv17;
  reg [3:0] op1_10_in18;
  reg       op1_10_inv18;
  reg [3:0] op1_10_in19;
  reg       op1_10_inv19;
  reg [3:0] op1_10_in20;
  reg       op1_10_inv20;
  reg [3:0] op1_10_in21;
  reg       op1_10_inv21;
  reg [3:0] op1_10_in22;
  reg       op1_10_inv22;
  reg [3:0] op1_10_in23;
  reg       op1_10_inv23;
  reg [3:0] op1_10_in24;
  reg       op1_10_inv24;
  reg [3:0] op1_10_in25;
  reg       op1_10_inv25;
  reg [3:0] op1_10_in26;
  reg       op1_10_inv26;
  reg [3:0] op1_10_in27;
  reg       op1_10_inv27;
  reg [3:0] op1_10_in28;
  reg       op1_10_inv28;
  reg [3:0] op1_10_in29;
  reg       op1_10_inv29;
  reg [3:0] op1_10_in30;
  reg       op1_10_inv30;
  reg [3:0] op1_10_in31;
  reg       op1_10_inv31;
  wire [8:0] op1_10_out;
  affine2_op1 op1_10(
    .data0_in(op1_10_in00),
    .inv0_in(op1_10_inv00),
    .data1_in(op1_10_in01),
    .inv1_in(op1_10_inv01),
    .data2_in(op1_10_in02),
    .inv2_in(op1_10_inv02),
    .data3_in(op1_10_in03),
    .inv3_in(op1_10_inv03),
    .data4_in(op1_10_in04),
    .inv4_in(op1_10_inv04),
    .data5_in(op1_10_in05),
    .inv5_in(op1_10_inv05),
    .data6_in(op1_10_in06),
    .inv6_in(op1_10_inv06),
    .data7_in(op1_10_in07),
    .inv7_in(op1_10_inv07),
    .data8_in(op1_10_in08),
    .inv8_in(op1_10_inv08),
    .data9_in(op1_10_in09),
    .inv9_in(op1_10_inv09),
    .data10_in(op1_10_in10),
    .inv10_in(op1_10_inv10),
    .data11_in(op1_10_in11),
    .inv11_in(op1_10_inv11),
    .data12_in(op1_10_in12),
    .inv12_in(op1_10_inv12),
    .data13_in(op1_10_in13),
    .inv13_in(op1_10_inv13),
    .data14_in(op1_10_in14),
    .inv14_in(op1_10_inv14),
    .data15_in(op1_10_in15),
    .inv15_in(op1_10_inv15),
    .data16_in(op1_10_in16),
    .inv16_in(op1_10_inv16),
    .data17_in(op1_10_in17),
    .inv17_in(op1_10_inv17),
    .data18_in(op1_10_in18),
    .inv18_in(op1_10_inv18),
    .data19_in(op1_10_in19),
    .inv19_in(op1_10_inv19),
    .data20_in(op1_10_in20),
    .inv20_in(op1_10_inv20),
    .data21_in(op1_10_in21),
    .inv21_in(op1_10_inv21),
    .data22_in(op1_10_in22),
    .inv22_in(op1_10_inv22),
    .data23_in(op1_10_in23),
    .inv23_in(op1_10_inv23),
    .data24_in(op1_10_in24),
    .inv24_in(op1_10_inv24),
    .data25_in(op1_10_in25),
    .inv25_in(op1_10_inv25),
    .data26_in(op1_10_in26),
    .inv26_in(op1_10_inv26),
    .data27_in(op1_10_in27),
    .inv27_in(op1_10_inv27),
    .data28_in(op1_10_in28),
    .inv28_in(op1_10_inv28),
    .data29_in(op1_10_in29),
    .inv29_in(op1_10_inv29),
    .data30_in(op1_10_in30),
    .inv30_in(op1_10_inv30),
    .data31_in(op1_10_in31),
    .inv31_in(op1_10_inv31),
    .data_out(op1_10_out));

  // 11 番目の OP1
  reg [3:0] op1_11_in00;
  reg       op1_11_inv00;
  reg [3:0] op1_11_in01;
  reg       op1_11_inv01;
  reg [3:0] op1_11_in02;
  reg       op1_11_inv02;
  reg [3:0] op1_11_in03;
  reg       op1_11_inv03;
  reg [3:0] op1_11_in04;
  reg       op1_11_inv04;
  reg [3:0] op1_11_in05;
  reg       op1_11_inv05;
  reg [3:0] op1_11_in06;
  reg       op1_11_inv06;
  reg [3:0] op1_11_in07;
  reg       op1_11_inv07;
  reg [3:0] op1_11_in08;
  reg       op1_11_inv08;
  reg [3:0] op1_11_in09;
  reg       op1_11_inv09;
  reg [3:0] op1_11_in10;
  reg       op1_11_inv10;
  reg [3:0] op1_11_in11;
  reg       op1_11_inv11;
  reg [3:0] op1_11_in12;
  reg       op1_11_inv12;
  reg [3:0] op1_11_in13;
  reg       op1_11_inv13;
  reg [3:0] op1_11_in14;
  reg       op1_11_inv14;
  reg [3:0] op1_11_in15;
  reg       op1_11_inv15;
  reg [3:0] op1_11_in16;
  reg       op1_11_inv16;
  reg [3:0] op1_11_in17;
  reg       op1_11_inv17;
  reg [3:0] op1_11_in18;
  reg       op1_11_inv18;
  reg [3:0] op1_11_in19;
  reg       op1_11_inv19;
  reg [3:0] op1_11_in20;
  reg       op1_11_inv20;
  reg [3:0] op1_11_in21;
  reg       op1_11_inv21;
  reg [3:0] op1_11_in22;
  reg       op1_11_inv22;
  reg [3:0] op1_11_in23;
  reg       op1_11_inv23;
  reg [3:0] op1_11_in24;
  reg       op1_11_inv24;
  reg [3:0] op1_11_in25;
  reg       op1_11_inv25;
  reg [3:0] op1_11_in26;
  reg       op1_11_inv26;
  reg [3:0] op1_11_in27;
  reg       op1_11_inv27;
  reg [3:0] op1_11_in28;
  reg       op1_11_inv28;
  reg [3:0] op1_11_in29;
  reg       op1_11_inv29;
  reg [3:0] op1_11_in30;
  reg       op1_11_inv30;
  reg [3:0] op1_11_in31;
  reg       op1_11_inv31;
  wire [8:0] op1_11_out;
  affine2_op1 op1_11(
    .data0_in(op1_11_in00),
    .inv0_in(op1_11_inv00),
    .data1_in(op1_11_in01),
    .inv1_in(op1_11_inv01),
    .data2_in(op1_11_in02),
    .inv2_in(op1_11_inv02),
    .data3_in(op1_11_in03),
    .inv3_in(op1_11_inv03),
    .data4_in(op1_11_in04),
    .inv4_in(op1_11_inv04),
    .data5_in(op1_11_in05),
    .inv5_in(op1_11_inv05),
    .data6_in(op1_11_in06),
    .inv6_in(op1_11_inv06),
    .data7_in(op1_11_in07),
    .inv7_in(op1_11_inv07),
    .data8_in(op1_11_in08),
    .inv8_in(op1_11_inv08),
    .data9_in(op1_11_in09),
    .inv9_in(op1_11_inv09),
    .data10_in(op1_11_in10),
    .inv10_in(op1_11_inv10),
    .data11_in(op1_11_in11),
    .inv11_in(op1_11_inv11),
    .data12_in(op1_11_in12),
    .inv12_in(op1_11_inv12),
    .data13_in(op1_11_in13),
    .inv13_in(op1_11_inv13),
    .data14_in(op1_11_in14),
    .inv14_in(op1_11_inv14),
    .data15_in(op1_11_in15),
    .inv15_in(op1_11_inv15),
    .data16_in(op1_11_in16),
    .inv16_in(op1_11_inv16),
    .data17_in(op1_11_in17),
    .inv17_in(op1_11_inv17),
    .data18_in(op1_11_in18),
    .inv18_in(op1_11_inv18),
    .data19_in(op1_11_in19),
    .inv19_in(op1_11_inv19),
    .data20_in(op1_11_in20),
    .inv20_in(op1_11_inv20),
    .data21_in(op1_11_in21),
    .inv21_in(op1_11_inv21),
    .data22_in(op1_11_in22),
    .inv22_in(op1_11_inv22),
    .data23_in(op1_11_in23),
    .inv23_in(op1_11_inv23),
    .data24_in(op1_11_in24),
    .inv24_in(op1_11_inv24),
    .data25_in(op1_11_in25),
    .inv25_in(op1_11_inv25),
    .data26_in(op1_11_in26),
    .inv26_in(op1_11_inv26),
    .data27_in(op1_11_in27),
    .inv27_in(op1_11_inv27),
    .data28_in(op1_11_in28),
    .inv28_in(op1_11_inv28),
    .data29_in(op1_11_in29),
    .inv29_in(op1_11_inv29),
    .data30_in(op1_11_in30),
    .inv30_in(op1_11_inv30),
    .data31_in(op1_11_in31),
    .inv31_in(op1_11_inv31),
    .data_out(op1_11_out));

  // 12 番目の OP1
  reg [3:0] op1_12_in00;
  reg       op1_12_inv00;
  reg [3:0] op1_12_in01;
  reg       op1_12_inv01;
  reg [3:0] op1_12_in02;
  reg       op1_12_inv02;
  reg [3:0] op1_12_in03;
  reg       op1_12_inv03;
  reg [3:0] op1_12_in04;
  reg       op1_12_inv04;
  reg [3:0] op1_12_in05;
  reg       op1_12_inv05;
  reg [3:0] op1_12_in06;
  reg       op1_12_inv06;
  reg [3:0] op1_12_in07;
  reg       op1_12_inv07;
  reg [3:0] op1_12_in08;
  reg       op1_12_inv08;
  reg [3:0] op1_12_in09;
  reg       op1_12_inv09;
  reg [3:0] op1_12_in10;
  reg       op1_12_inv10;
  reg [3:0] op1_12_in11;
  reg       op1_12_inv11;
  reg [3:0] op1_12_in12;
  reg       op1_12_inv12;
  reg [3:0] op1_12_in13;
  reg       op1_12_inv13;
  reg [3:0] op1_12_in14;
  reg       op1_12_inv14;
  reg [3:0] op1_12_in15;
  reg       op1_12_inv15;
  reg [3:0] op1_12_in16;
  reg       op1_12_inv16;
  reg [3:0] op1_12_in17;
  reg       op1_12_inv17;
  reg [3:0] op1_12_in18;
  reg       op1_12_inv18;
  reg [3:0] op1_12_in19;
  reg       op1_12_inv19;
  reg [3:0] op1_12_in20;
  reg       op1_12_inv20;
  reg [3:0] op1_12_in21;
  reg       op1_12_inv21;
  reg [3:0] op1_12_in22;
  reg       op1_12_inv22;
  reg [3:0] op1_12_in23;
  reg       op1_12_inv23;
  reg [3:0] op1_12_in24;
  reg       op1_12_inv24;
  reg [3:0] op1_12_in25;
  reg       op1_12_inv25;
  reg [3:0] op1_12_in26;
  reg       op1_12_inv26;
  reg [3:0] op1_12_in27;
  reg       op1_12_inv27;
  reg [3:0] op1_12_in28;
  reg       op1_12_inv28;
  reg [3:0] op1_12_in29;
  reg       op1_12_inv29;
  reg [3:0] op1_12_in30;
  reg       op1_12_inv30;
  reg [3:0] op1_12_in31;
  reg       op1_12_inv31;
  wire [8:0] op1_12_out;
  affine2_op1 op1_12(
    .data0_in(op1_12_in00),
    .inv0_in(op1_12_inv00),
    .data1_in(op1_12_in01),
    .inv1_in(op1_12_inv01),
    .data2_in(op1_12_in02),
    .inv2_in(op1_12_inv02),
    .data3_in(op1_12_in03),
    .inv3_in(op1_12_inv03),
    .data4_in(op1_12_in04),
    .inv4_in(op1_12_inv04),
    .data5_in(op1_12_in05),
    .inv5_in(op1_12_inv05),
    .data6_in(op1_12_in06),
    .inv6_in(op1_12_inv06),
    .data7_in(op1_12_in07),
    .inv7_in(op1_12_inv07),
    .data8_in(op1_12_in08),
    .inv8_in(op1_12_inv08),
    .data9_in(op1_12_in09),
    .inv9_in(op1_12_inv09),
    .data10_in(op1_12_in10),
    .inv10_in(op1_12_inv10),
    .data11_in(op1_12_in11),
    .inv11_in(op1_12_inv11),
    .data12_in(op1_12_in12),
    .inv12_in(op1_12_inv12),
    .data13_in(op1_12_in13),
    .inv13_in(op1_12_inv13),
    .data14_in(op1_12_in14),
    .inv14_in(op1_12_inv14),
    .data15_in(op1_12_in15),
    .inv15_in(op1_12_inv15),
    .data16_in(op1_12_in16),
    .inv16_in(op1_12_inv16),
    .data17_in(op1_12_in17),
    .inv17_in(op1_12_inv17),
    .data18_in(op1_12_in18),
    .inv18_in(op1_12_inv18),
    .data19_in(op1_12_in19),
    .inv19_in(op1_12_inv19),
    .data20_in(op1_12_in20),
    .inv20_in(op1_12_inv20),
    .data21_in(op1_12_in21),
    .inv21_in(op1_12_inv21),
    .data22_in(op1_12_in22),
    .inv22_in(op1_12_inv22),
    .data23_in(op1_12_in23),
    .inv23_in(op1_12_inv23),
    .data24_in(op1_12_in24),
    .inv24_in(op1_12_inv24),
    .data25_in(op1_12_in25),
    .inv25_in(op1_12_inv25),
    .data26_in(op1_12_in26),
    .inv26_in(op1_12_inv26),
    .data27_in(op1_12_in27),
    .inv27_in(op1_12_inv27),
    .data28_in(op1_12_in28),
    .inv28_in(op1_12_inv28),
    .data29_in(op1_12_in29),
    .inv29_in(op1_12_inv29),
    .data30_in(op1_12_in30),
    .inv30_in(op1_12_inv30),
    .data31_in(op1_12_in31),
    .inv31_in(op1_12_inv31),
    .data_out(op1_12_out));

  // 13 番目の OP1
  reg [3:0] op1_13_in00;
  reg       op1_13_inv00;
  reg [3:0] op1_13_in01;
  reg       op1_13_inv01;
  reg [3:0] op1_13_in02;
  reg       op1_13_inv02;
  reg [3:0] op1_13_in03;
  reg       op1_13_inv03;
  reg [3:0] op1_13_in04;
  reg       op1_13_inv04;
  reg [3:0] op1_13_in05;
  reg       op1_13_inv05;
  reg [3:0] op1_13_in06;
  reg       op1_13_inv06;
  reg [3:0] op1_13_in07;
  reg       op1_13_inv07;
  reg [3:0] op1_13_in08;
  reg       op1_13_inv08;
  reg [3:0] op1_13_in09;
  reg       op1_13_inv09;
  reg [3:0] op1_13_in10;
  reg       op1_13_inv10;
  reg [3:0] op1_13_in11;
  reg       op1_13_inv11;
  reg [3:0] op1_13_in12;
  reg       op1_13_inv12;
  reg [3:0] op1_13_in13;
  reg       op1_13_inv13;
  reg [3:0] op1_13_in14;
  reg       op1_13_inv14;
  reg [3:0] op1_13_in15;
  reg       op1_13_inv15;
  reg [3:0] op1_13_in16;
  reg       op1_13_inv16;
  reg [3:0] op1_13_in17;
  reg       op1_13_inv17;
  reg [3:0] op1_13_in18;
  reg       op1_13_inv18;
  reg [3:0] op1_13_in19;
  reg       op1_13_inv19;
  reg [3:0] op1_13_in20;
  reg       op1_13_inv20;
  reg [3:0] op1_13_in21;
  reg       op1_13_inv21;
  reg [3:0] op1_13_in22;
  reg       op1_13_inv22;
  reg [3:0] op1_13_in23;
  reg       op1_13_inv23;
  reg [3:0] op1_13_in24;
  reg       op1_13_inv24;
  reg [3:0] op1_13_in25;
  reg       op1_13_inv25;
  reg [3:0] op1_13_in26;
  reg       op1_13_inv26;
  reg [3:0] op1_13_in27;
  reg       op1_13_inv27;
  reg [3:0] op1_13_in28;
  reg       op1_13_inv28;
  reg [3:0] op1_13_in29;
  reg       op1_13_inv29;
  reg [3:0] op1_13_in30;
  reg       op1_13_inv30;
  reg [3:0] op1_13_in31;
  reg       op1_13_inv31;
  wire [8:0] op1_13_out;
  affine2_op1 op1_13(
    .data0_in(op1_13_in00),
    .inv0_in(op1_13_inv00),
    .data1_in(op1_13_in01),
    .inv1_in(op1_13_inv01),
    .data2_in(op1_13_in02),
    .inv2_in(op1_13_inv02),
    .data3_in(op1_13_in03),
    .inv3_in(op1_13_inv03),
    .data4_in(op1_13_in04),
    .inv4_in(op1_13_inv04),
    .data5_in(op1_13_in05),
    .inv5_in(op1_13_inv05),
    .data6_in(op1_13_in06),
    .inv6_in(op1_13_inv06),
    .data7_in(op1_13_in07),
    .inv7_in(op1_13_inv07),
    .data8_in(op1_13_in08),
    .inv8_in(op1_13_inv08),
    .data9_in(op1_13_in09),
    .inv9_in(op1_13_inv09),
    .data10_in(op1_13_in10),
    .inv10_in(op1_13_inv10),
    .data11_in(op1_13_in11),
    .inv11_in(op1_13_inv11),
    .data12_in(op1_13_in12),
    .inv12_in(op1_13_inv12),
    .data13_in(op1_13_in13),
    .inv13_in(op1_13_inv13),
    .data14_in(op1_13_in14),
    .inv14_in(op1_13_inv14),
    .data15_in(op1_13_in15),
    .inv15_in(op1_13_inv15),
    .data16_in(op1_13_in16),
    .inv16_in(op1_13_inv16),
    .data17_in(op1_13_in17),
    .inv17_in(op1_13_inv17),
    .data18_in(op1_13_in18),
    .inv18_in(op1_13_inv18),
    .data19_in(op1_13_in19),
    .inv19_in(op1_13_inv19),
    .data20_in(op1_13_in20),
    .inv20_in(op1_13_inv20),
    .data21_in(op1_13_in21),
    .inv21_in(op1_13_inv21),
    .data22_in(op1_13_in22),
    .inv22_in(op1_13_inv22),
    .data23_in(op1_13_in23),
    .inv23_in(op1_13_inv23),
    .data24_in(op1_13_in24),
    .inv24_in(op1_13_inv24),
    .data25_in(op1_13_in25),
    .inv25_in(op1_13_inv25),
    .data26_in(op1_13_in26),
    .inv26_in(op1_13_inv26),
    .data27_in(op1_13_in27),
    .inv27_in(op1_13_inv27),
    .data28_in(op1_13_in28),
    .inv28_in(op1_13_inv28),
    .data29_in(op1_13_in29),
    .inv29_in(op1_13_inv29),
    .data30_in(op1_13_in30),
    .inv30_in(op1_13_inv30),
    .data31_in(op1_13_in31),
    .inv31_in(op1_13_inv31),
    .data_out(op1_13_out));

  // 14 番目の OP1
  reg [3:0] op1_14_in00;
  reg       op1_14_inv00;
  reg [3:0] op1_14_in01;
  reg       op1_14_inv01;
  reg [3:0] op1_14_in02;
  reg       op1_14_inv02;
  reg [3:0] op1_14_in03;
  reg       op1_14_inv03;
  reg [3:0] op1_14_in04;
  reg       op1_14_inv04;
  reg [3:0] op1_14_in05;
  reg       op1_14_inv05;
  reg [3:0] op1_14_in06;
  reg       op1_14_inv06;
  reg [3:0] op1_14_in07;
  reg       op1_14_inv07;
  reg [3:0] op1_14_in08;
  reg       op1_14_inv08;
  reg [3:0] op1_14_in09;
  reg       op1_14_inv09;
  reg [3:0] op1_14_in10;
  reg       op1_14_inv10;
  reg [3:0] op1_14_in11;
  reg       op1_14_inv11;
  reg [3:0] op1_14_in12;
  reg       op1_14_inv12;
  reg [3:0] op1_14_in13;
  reg       op1_14_inv13;
  reg [3:0] op1_14_in14;
  reg       op1_14_inv14;
  reg [3:0] op1_14_in15;
  reg       op1_14_inv15;
  reg [3:0] op1_14_in16;
  reg       op1_14_inv16;
  reg [3:0] op1_14_in17;
  reg       op1_14_inv17;
  reg [3:0] op1_14_in18;
  reg       op1_14_inv18;
  reg [3:0] op1_14_in19;
  reg       op1_14_inv19;
  reg [3:0] op1_14_in20;
  reg       op1_14_inv20;
  reg [3:0] op1_14_in21;
  reg       op1_14_inv21;
  reg [3:0] op1_14_in22;
  reg       op1_14_inv22;
  reg [3:0] op1_14_in23;
  reg       op1_14_inv23;
  reg [3:0] op1_14_in24;
  reg       op1_14_inv24;
  reg [3:0] op1_14_in25;
  reg       op1_14_inv25;
  reg [3:0] op1_14_in26;
  reg       op1_14_inv26;
  reg [3:0] op1_14_in27;
  reg       op1_14_inv27;
  reg [3:0] op1_14_in28;
  reg       op1_14_inv28;
  reg [3:0] op1_14_in29;
  reg       op1_14_inv29;
  reg [3:0] op1_14_in30;
  reg       op1_14_inv30;
  reg [3:0] op1_14_in31;
  reg       op1_14_inv31;
  wire [8:0] op1_14_out;
  affine2_op1 op1_14(
    .data0_in(op1_14_in00),
    .inv0_in(op1_14_inv00),
    .data1_in(op1_14_in01),
    .inv1_in(op1_14_inv01),
    .data2_in(op1_14_in02),
    .inv2_in(op1_14_inv02),
    .data3_in(op1_14_in03),
    .inv3_in(op1_14_inv03),
    .data4_in(op1_14_in04),
    .inv4_in(op1_14_inv04),
    .data5_in(op1_14_in05),
    .inv5_in(op1_14_inv05),
    .data6_in(op1_14_in06),
    .inv6_in(op1_14_inv06),
    .data7_in(op1_14_in07),
    .inv7_in(op1_14_inv07),
    .data8_in(op1_14_in08),
    .inv8_in(op1_14_inv08),
    .data9_in(op1_14_in09),
    .inv9_in(op1_14_inv09),
    .data10_in(op1_14_in10),
    .inv10_in(op1_14_inv10),
    .data11_in(op1_14_in11),
    .inv11_in(op1_14_inv11),
    .data12_in(op1_14_in12),
    .inv12_in(op1_14_inv12),
    .data13_in(op1_14_in13),
    .inv13_in(op1_14_inv13),
    .data14_in(op1_14_in14),
    .inv14_in(op1_14_inv14),
    .data15_in(op1_14_in15),
    .inv15_in(op1_14_inv15),
    .data16_in(op1_14_in16),
    .inv16_in(op1_14_inv16),
    .data17_in(op1_14_in17),
    .inv17_in(op1_14_inv17),
    .data18_in(op1_14_in18),
    .inv18_in(op1_14_inv18),
    .data19_in(op1_14_in19),
    .inv19_in(op1_14_inv19),
    .data20_in(op1_14_in20),
    .inv20_in(op1_14_inv20),
    .data21_in(op1_14_in21),
    .inv21_in(op1_14_inv21),
    .data22_in(op1_14_in22),
    .inv22_in(op1_14_inv22),
    .data23_in(op1_14_in23),
    .inv23_in(op1_14_inv23),
    .data24_in(op1_14_in24),
    .inv24_in(op1_14_inv24),
    .data25_in(op1_14_in25),
    .inv25_in(op1_14_inv25),
    .data26_in(op1_14_in26),
    .inv26_in(op1_14_inv26),
    .data27_in(op1_14_in27),
    .inv27_in(op1_14_inv27),
    .data28_in(op1_14_in28),
    .inv28_in(op1_14_inv28),
    .data29_in(op1_14_in29),
    .inv29_in(op1_14_inv29),
    .data30_in(op1_14_in30),
    .inv30_in(op1_14_inv30),
    .data31_in(op1_14_in31),
    .inv31_in(op1_14_inv31),
    .data_out(op1_14_out));

  // 15 番目の OP1
  reg [3:0] op1_15_in00;
  reg       op1_15_inv00;
  reg [3:0] op1_15_in01;
  reg       op1_15_inv01;
  reg [3:0] op1_15_in02;
  reg       op1_15_inv02;
  reg [3:0] op1_15_in03;
  reg       op1_15_inv03;
  reg [3:0] op1_15_in04;
  reg       op1_15_inv04;
  reg [3:0] op1_15_in05;
  reg       op1_15_inv05;
  reg [3:0] op1_15_in06;
  reg       op1_15_inv06;
  reg [3:0] op1_15_in07;
  reg       op1_15_inv07;
  reg [3:0] op1_15_in08;
  reg       op1_15_inv08;
  reg [3:0] op1_15_in09;
  reg       op1_15_inv09;
  reg [3:0] op1_15_in10;
  reg       op1_15_inv10;
  reg [3:0] op1_15_in11;
  reg       op1_15_inv11;
  reg [3:0] op1_15_in12;
  reg       op1_15_inv12;
  reg [3:0] op1_15_in13;
  reg       op1_15_inv13;
  reg [3:0] op1_15_in14;
  reg       op1_15_inv14;
  reg [3:0] op1_15_in15;
  reg       op1_15_inv15;
  reg [3:0] op1_15_in16;
  reg       op1_15_inv16;
  reg [3:0] op1_15_in17;
  reg       op1_15_inv17;
  reg [3:0] op1_15_in18;
  reg       op1_15_inv18;
  reg [3:0] op1_15_in19;
  reg       op1_15_inv19;
  reg [3:0] op1_15_in20;
  reg       op1_15_inv20;
  reg [3:0] op1_15_in21;
  reg       op1_15_inv21;
  reg [3:0] op1_15_in22;
  reg       op1_15_inv22;
  reg [3:0] op1_15_in23;
  reg       op1_15_inv23;
  reg [3:0] op1_15_in24;
  reg       op1_15_inv24;
  reg [3:0] op1_15_in25;
  reg       op1_15_inv25;
  reg [3:0] op1_15_in26;
  reg       op1_15_inv26;
  reg [3:0] op1_15_in27;
  reg       op1_15_inv27;
  reg [3:0] op1_15_in28;
  reg       op1_15_inv28;
  reg [3:0] op1_15_in29;
  reg       op1_15_inv29;
  reg [3:0] op1_15_in30;
  reg       op1_15_inv30;
  reg [3:0] op1_15_in31;
  reg       op1_15_inv31;
  wire [8:0] op1_15_out;
  affine2_op1 op1_15(
    .data0_in(op1_15_in00),
    .inv0_in(op1_15_inv00),
    .data1_in(op1_15_in01),
    .inv1_in(op1_15_inv01),
    .data2_in(op1_15_in02),
    .inv2_in(op1_15_inv02),
    .data3_in(op1_15_in03),
    .inv3_in(op1_15_inv03),
    .data4_in(op1_15_in04),
    .inv4_in(op1_15_inv04),
    .data5_in(op1_15_in05),
    .inv5_in(op1_15_inv05),
    .data6_in(op1_15_in06),
    .inv6_in(op1_15_inv06),
    .data7_in(op1_15_in07),
    .inv7_in(op1_15_inv07),
    .data8_in(op1_15_in08),
    .inv8_in(op1_15_inv08),
    .data9_in(op1_15_in09),
    .inv9_in(op1_15_inv09),
    .data10_in(op1_15_in10),
    .inv10_in(op1_15_inv10),
    .data11_in(op1_15_in11),
    .inv11_in(op1_15_inv11),
    .data12_in(op1_15_in12),
    .inv12_in(op1_15_inv12),
    .data13_in(op1_15_in13),
    .inv13_in(op1_15_inv13),
    .data14_in(op1_15_in14),
    .inv14_in(op1_15_inv14),
    .data15_in(op1_15_in15),
    .inv15_in(op1_15_inv15),
    .data16_in(op1_15_in16),
    .inv16_in(op1_15_inv16),
    .data17_in(op1_15_in17),
    .inv17_in(op1_15_inv17),
    .data18_in(op1_15_in18),
    .inv18_in(op1_15_inv18),
    .data19_in(op1_15_in19),
    .inv19_in(op1_15_inv19),
    .data20_in(op1_15_in20),
    .inv20_in(op1_15_inv20),
    .data21_in(op1_15_in21),
    .inv21_in(op1_15_inv21),
    .data22_in(op1_15_in22),
    .inv22_in(op1_15_inv22),
    .data23_in(op1_15_in23),
    .inv23_in(op1_15_inv23),
    .data24_in(op1_15_in24),
    .inv24_in(op1_15_inv24),
    .data25_in(op1_15_in25),
    .inv25_in(op1_15_inv25),
    .data26_in(op1_15_in26),
    .inv26_in(op1_15_inv26),
    .data27_in(op1_15_in27),
    .inv27_in(op1_15_inv27),
    .data28_in(op1_15_in28),
    .inv28_in(op1_15_inv28),
    .data29_in(op1_15_in29),
    .inv29_in(op1_15_inv29),
    .data30_in(op1_15_in30),
    .inv30_in(op1_15_inv30),
    .data31_in(op1_15_in31),
    .inv31_in(op1_15_inv31),
    .data_out(op1_15_out));

  // 0 番目の OP2
  reg [8:0] op2_00_in00;
  reg [8:0] op2_00_in01;
  reg [8:0] op2_00_in02;
  reg [8:0] op2_00_in03;
  reg [8:0] op2_00_in04;
  reg [8:0] op2_00_in05;
  reg [8:0] op2_00_in06;
  reg [8:0] op2_00_in07;
  reg [8:0] op2_00_in08;
  reg [8:0] op2_00_in09;
  reg [8:0] op2_00_in10;
  reg [8:0] op2_00_in11;
  reg [8:0] op2_00_in12;
  reg [8:0] op2_00_in13;
  reg [8:0] op2_00_in14;
  reg [8:0] op2_00_in15;
  reg [8:0] op2_00_in16;
  reg [8:0] op2_00_in17;
  reg [8:0] op2_00_in18;
  reg [8:0] op2_00_in19;
  reg [8:0] op2_00_in20;
  reg [8:0] op2_00_in21;
  reg [8:0] op2_00_in22;
  reg [8:0] op2_00_in23;
  reg [8:0] op2_00_in24;
  reg [8:0] op2_00_in25;
  reg [8:0] op2_00_in26;
  reg [8:0] op2_00_in27;
  reg [8:0] op2_00_in28;
  reg [8:0] op2_00_in29;
  reg [8:0] op2_00_in30;
  reg [8:0] op2_00_bias;
  wire [8:0] op2_00_out;
  affine2_op2 op2_00(
    .data0_in(op2_00_in00),
    .data1_in(op2_00_in01),
    .data2_in(op2_00_in02),
    .data3_in(op2_00_in03),
    .data4_in(op2_00_in04),
    .data5_in(op2_00_in05),
    .data6_in(op2_00_in06),
    .data7_in(op2_00_in07),
    .data8_in(op2_00_in08),
    .data9_in(op2_00_in09),
    .data10_in(op2_00_in10),
    .data11_in(op2_00_in11),
    .data12_in(op2_00_in12),
    .data13_in(op2_00_in13),
    .data14_in(op2_00_in14),
    .data15_in(op2_00_in15),
    .data16_in(op2_00_in16),
    .data17_in(op2_00_in17),
    .data18_in(op2_00_in18),
    .data19_in(op2_00_in19),
    .data20_in(op2_00_in20),
    .data21_in(op2_00_in21),
    .data22_in(op2_00_in22),
    .data23_in(op2_00_in23),
    .data24_in(op2_00_in24),
    .data25_in(op2_00_in25),
    .data26_in(op2_00_in26),
    .data27_in(op2_00_in27),
    .data28_in(op2_00_in28),
    .data29_in(op2_00_in29),
    .data30_in(op2_00_in30),
    .data31_in(op2_00_bias),
    .data_out(op2_00_out));

  // 1 番目の OP2
  reg [8:0] op2_01_in00;
  reg [8:0] op2_01_in01;
  reg [8:0] op2_01_in02;
  reg [8:0] op2_01_in03;
  reg [8:0] op2_01_in04;
  reg [8:0] op2_01_in05;
  reg [8:0] op2_01_in06;
  reg [8:0] op2_01_in07;
  reg [8:0] op2_01_in08;
  reg [8:0] op2_01_in09;
  reg [8:0] op2_01_in10;
  reg [8:0] op2_01_in11;
  reg [8:0] op2_01_in12;
  reg [8:0] op2_01_in13;
  reg [8:0] op2_01_in14;
  reg [8:0] op2_01_in15;
  reg [8:0] op2_01_in16;
  reg [8:0] op2_01_in17;
  reg [8:0] op2_01_in18;
  reg [8:0] op2_01_in19;
  reg [8:0] op2_01_in20;
  reg [8:0] op2_01_in21;
  reg [8:0] op2_01_in22;
  reg [8:0] op2_01_in23;
  reg [8:0] op2_01_in24;
  reg [8:0] op2_01_in25;
  reg [8:0] op2_01_in26;
  reg [8:0] op2_01_in27;
  reg [8:0] op2_01_in28;
  reg [8:0] op2_01_in29;
  reg [8:0] op2_01_in30;
  reg [8:0] op2_01_bias;
  wire [8:0] op2_01_out;
  affine2_op2 op2_01(
    .data0_in(op2_01_in00),
    .data1_in(op2_01_in01),
    .data2_in(op2_01_in02),
    .data3_in(op2_01_in03),
    .data4_in(op2_01_in04),
    .data5_in(op2_01_in05),
    .data6_in(op2_01_in06),
    .data7_in(op2_01_in07),
    .data8_in(op2_01_in08),
    .data9_in(op2_01_in09),
    .data10_in(op2_01_in10),
    .data11_in(op2_01_in11),
    .data12_in(op2_01_in12),
    .data13_in(op2_01_in13),
    .data14_in(op2_01_in14),
    .data15_in(op2_01_in15),
    .data16_in(op2_01_in16),
    .data17_in(op2_01_in17),
    .data18_in(op2_01_in18),
    .data19_in(op2_01_in19),
    .data20_in(op2_01_in20),
    .data21_in(op2_01_in21),
    .data22_in(op2_01_in22),
    .data23_in(op2_01_in23),
    .data24_in(op2_01_in24),
    .data25_in(op2_01_in25),
    .data26_in(op2_01_in26),
    .data27_in(op2_01_in27),
    .data28_in(op2_01_in28),
    .data29_in(op2_01_in29),
    .data30_in(op2_01_in30),
    .data31_in(op2_01_bias),
    .data_out(op2_01_out));

  // 2 番目の OP2
  reg [8:0] op2_02_in00;
  reg [8:0] op2_02_in01;
  reg [8:0] op2_02_in02;
  reg [8:0] op2_02_in03;
  reg [8:0] op2_02_in04;
  reg [8:0] op2_02_in05;
  reg [8:0] op2_02_in06;
  reg [8:0] op2_02_in07;
  reg [8:0] op2_02_in08;
  reg [8:0] op2_02_in09;
  reg [8:0] op2_02_in10;
  reg [8:0] op2_02_in11;
  reg [8:0] op2_02_in12;
  reg [8:0] op2_02_in13;
  reg [8:0] op2_02_in14;
  reg [8:0] op2_02_in15;
  reg [8:0] op2_02_in16;
  reg [8:0] op2_02_in17;
  reg [8:0] op2_02_in18;
  reg [8:0] op2_02_in19;
  reg [8:0] op2_02_in20;
  reg [8:0] op2_02_in21;
  reg [8:0] op2_02_in22;
  reg [8:0] op2_02_in23;
  reg [8:0] op2_02_in24;
  reg [8:0] op2_02_in25;
  reg [8:0] op2_02_in26;
  reg [8:0] op2_02_in27;
  reg [8:0] op2_02_in28;
  reg [8:0] op2_02_in29;
  reg [8:0] op2_02_in30;
  reg [8:0] op2_02_bias;
  wire [8:0] op2_02_out;
  affine2_op2 op2_02(
    .data0_in(op2_02_in00),
    .data1_in(op2_02_in01),
    .data2_in(op2_02_in02),
    .data3_in(op2_02_in03),
    .data4_in(op2_02_in04),
    .data5_in(op2_02_in05),
    .data6_in(op2_02_in06),
    .data7_in(op2_02_in07),
    .data8_in(op2_02_in08),
    .data9_in(op2_02_in09),
    .data10_in(op2_02_in10),
    .data11_in(op2_02_in11),
    .data12_in(op2_02_in12),
    .data13_in(op2_02_in13),
    .data14_in(op2_02_in14),
    .data15_in(op2_02_in15),
    .data16_in(op2_02_in16),
    .data17_in(op2_02_in17),
    .data18_in(op2_02_in18),
    .data19_in(op2_02_in19),
    .data20_in(op2_02_in20),
    .data21_in(op2_02_in21),
    .data22_in(op2_02_in22),
    .data23_in(op2_02_in23),
    .data24_in(op2_02_in24),
    .data25_in(op2_02_in25),
    .data26_in(op2_02_in26),
    .data27_in(op2_02_in27),
    .data28_in(op2_02_in28),
    .data29_in(op2_02_in29),
    .data30_in(op2_02_in30),
    .data31_in(op2_02_bias),
    .data_out(op2_02_out));

  // 3 番目の OP2
  reg [8:0] op2_03_in00;
  reg [8:0] op2_03_in01;
  reg [8:0] op2_03_in02;
  reg [8:0] op2_03_in03;
  reg [8:0] op2_03_in04;
  reg [8:0] op2_03_in05;
  reg [8:0] op2_03_in06;
  reg [8:0] op2_03_in07;
  reg [8:0] op2_03_in08;
  reg [8:0] op2_03_in09;
  reg [8:0] op2_03_in10;
  reg [8:0] op2_03_in11;
  reg [8:0] op2_03_in12;
  reg [8:0] op2_03_in13;
  reg [8:0] op2_03_in14;
  reg [8:0] op2_03_in15;
  reg [8:0] op2_03_in16;
  reg [8:0] op2_03_in17;
  reg [8:0] op2_03_in18;
  reg [8:0] op2_03_in19;
  reg [8:0] op2_03_in20;
  reg [8:0] op2_03_in21;
  reg [8:0] op2_03_in22;
  reg [8:0] op2_03_in23;
  reg [8:0] op2_03_in24;
  reg [8:0] op2_03_in25;
  reg [8:0] op2_03_in26;
  reg [8:0] op2_03_in27;
  reg [8:0] op2_03_in28;
  reg [8:0] op2_03_in29;
  reg [8:0] op2_03_in30;
  reg [8:0] op2_03_bias;
  wire [8:0] op2_03_out;
  affine2_op2 op2_03(
    .data0_in(op2_03_in00),
    .data1_in(op2_03_in01),
    .data2_in(op2_03_in02),
    .data3_in(op2_03_in03),
    .data4_in(op2_03_in04),
    .data5_in(op2_03_in05),
    .data6_in(op2_03_in06),
    .data7_in(op2_03_in07),
    .data8_in(op2_03_in08),
    .data9_in(op2_03_in09),
    .data10_in(op2_03_in10),
    .data11_in(op2_03_in11),
    .data12_in(op2_03_in12),
    .data13_in(op2_03_in13),
    .data14_in(op2_03_in14),
    .data15_in(op2_03_in15),
    .data16_in(op2_03_in16),
    .data17_in(op2_03_in17),
    .data18_in(op2_03_in18),
    .data19_in(op2_03_in19),
    .data20_in(op2_03_in20),
    .data21_in(op2_03_in21),
    .data22_in(op2_03_in22),
    .data23_in(op2_03_in23),
    .data24_in(op2_03_in24),
    .data25_in(op2_03_in25),
    .data26_in(op2_03_in26),
    .data27_in(op2_03_in27),
    .data28_in(op2_03_in28),
    .data29_in(op2_03_in29),
    .data30_in(op2_03_in30),
    .data31_in(op2_03_bias),
    .data_out(op2_03_out));

  // 4 番目の OP2
  reg [8:0] op2_04_in00;
  reg [8:0] op2_04_in01;
  reg [8:0] op2_04_in02;
  reg [8:0] op2_04_in03;
  reg [8:0] op2_04_in04;
  reg [8:0] op2_04_in05;
  reg [8:0] op2_04_in06;
  reg [8:0] op2_04_in07;
  reg [8:0] op2_04_in08;
  reg [8:0] op2_04_in09;
  reg [8:0] op2_04_in10;
  reg [8:0] op2_04_in11;
  reg [8:0] op2_04_in12;
  reg [8:0] op2_04_in13;
  reg [8:0] op2_04_in14;
  reg [8:0] op2_04_in15;
  reg [8:0] op2_04_in16;
  reg [8:0] op2_04_in17;
  reg [8:0] op2_04_in18;
  reg [8:0] op2_04_in19;
  reg [8:0] op2_04_in20;
  reg [8:0] op2_04_in21;
  reg [8:0] op2_04_in22;
  reg [8:0] op2_04_in23;
  reg [8:0] op2_04_in24;
  reg [8:0] op2_04_in25;
  reg [8:0] op2_04_in26;
  reg [8:0] op2_04_in27;
  reg [8:0] op2_04_in28;
  reg [8:0] op2_04_in29;
  reg [8:0] op2_04_in30;
  reg [8:0] op2_04_bias;
  wire [8:0] op2_04_out;
  affine2_op2 op2_04(
    .data0_in(op2_04_in00),
    .data1_in(op2_04_in01),
    .data2_in(op2_04_in02),
    .data3_in(op2_04_in03),
    .data4_in(op2_04_in04),
    .data5_in(op2_04_in05),
    .data6_in(op2_04_in06),
    .data7_in(op2_04_in07),
    .data8_in(op2_04_in08),
    .data9_in(op2_04_in09),
    .data10_in(op2_04_in10),
    .data11_in(op2_04_in11),
    .data12_in(op2_04_in12),
    .data13_in(op2_04_in13),
    .data14_in(op2_04_in14),
    .data15_in(op2_04_in15),
    .data16_in(op2_04_in16),
    .data17_in(op2_04_in17),
    .data18_in(op2_04_in18),
    .data19_in(op2_04_in19),
    .data20_in(op2_04_in20),
    .data21_in(op2_04_in21),
    .data22_in(op2_04_in22),
    .data23_in(op2_04_in23),
    .data24_in(op2_04_in24),
    .data25_in(op2_04_in25),
    .data26_in(op2_04_in26),
    .data27_in(op2_04_in27),
    .data28_in(op2_04_in28),
    .data29_in(op2_04_in29),
    .data30_in(op2_04_in30),
    .data31_in(op2_04_bias),
    .data_out(op2_04_out));

  // 5 番目の OP2
  reg [8:0] op2_05_in00;
  reg [8:0] op2_05_in01;
  reg [8:0] op2_05_in02;
  reg [8:0] op2_05_in03;
  reg [8:0] op2_05_in04;
  reg [8:0] op2_05_in05;
  reg [8:0] op2_05_in06;
  reg [8:0] op2_05_in07;
  reg [8:0] op2_05_in08;
  reg [8:0] op2_05_in09;
  reg [8:0] op2_05_in10;
  reg [8:0] op2_05_in11;
  reg [8:0] op2_05_in12;
  reg [8:0] op2_05_in13;
  reg [8:0] op2_05_in14;
  reg [8:0] op2_05_in15;
  reg [8:0] op2_05_in16;
  reg [8:0] op2_05_in17;
  reg [8:0] op2_05_in18;
  reg [8:0] op2_05_in19;
  reg [8:0] op2_05_in20;
  reg [8:0] op2_05_in21;
  reg [8:0] op2_05_in22;
  reg [8:0] op2_05_in23;
  reg [8:0] op2_05_in24;
  reg [8:0] op2_05_in25;
  reg [8:0] op2_05_in26;
  reg [8:0] op2_05_in27;
  reg [8:0] op2_05_in28;
  reg [8:0] op2_05_in29;
  reg [8:0] op2_05_in30;
  reg [8:0] op2_05_bias;
  wire [8:0] op2_05_out;
  affine2_op2 op2_05(
    .data0_in(op2_05_in00),
    .data1_in(op2_05_in01),
    .data2_in(op2_05_in02),
    .data3_in(op2_05_in03),
    .data4_in(op2_05_in04),
    .data5_in(op2_05_in05),
    .data6_in(op2_05_in06),
    .data7_in(op2_05_in07),
    .data8_in(op2_05_in08),
    .data9_in(op2_05_in09),
    .data10_in(op2_05_in10),
    .data11_in(op2_05_in11),
    .data12_in(op2_05_in12),
    .data13_in(op2_05_in13),
    .data14_in(op2_05_in14),
    .data15_in(op2_05_in15),
    .data16_in(op2_05_in16),
    .data17_in(op2_05_in17),
    .data18_in(op2_05_in18),
    .data19_in(op2_05_in19),
    .data20_in(op2_05_in20),
    .data21_in(op2_05_in21),
    .data22_in(op2_05_in22),
    .data23_in(op2_05_in23),
    .data24_in(op2_05_in24),
    .data25_in(op2_05_in25),
    .data26_in(op2_05_in26),
    .data27_in(op2_05_in27),
    .data28_in(op2_05_in28),
    .data29_in(op2_05_in29),
    .data30_in(op2_05_in30),
    .data31_in(op2_05_bias),
    .data_out(op2_05_out));

  // 6 番目の OP2
  reg [8:0] op2_06_in00;
  reg [8:0] op2_06_in01;
  reg [8:0] op2_06_in02;
  reg [8:0] op2_06_in03;
  reg [8:0] op2_06_in04;
  reg [8:0] op2_06_in05;
  reg [8:0] op2_06_in06;
  reg [8:0] op2_06_in07;
  reg [8:0] op2_06_in08;
  reg [8:0] op2_06_in09;
  reg [8:0] op2_06_in10;
  reg [8:0] op2_06_in11;
  reg [8:0] op2_06_in12;
  reg [8:0] op2_06_in13;
  reg [8:0] op2_06_in14;
  reg [8:0] op2_06_in15;
  reg [8:0] op2_06_in16;
  reg [8:0] op2_06_in17;
  reg [8:0] op2_06_in18;
  reg [8:0] op2_06_in19;
  reg [8:0] op2_06_in20;
  reg [8:0] op2_06_in21;
  reg [8:0] op2_06_in22;
  reg [8:0] op2_06_in23;
  reg [8:0] op2_06_in24;
  reg [8:0] op2_06_in25;
  reg [8:0] op2_06_in26;
  reg [8:0] op2_06_in27;
  reg [8:0] op2_06_in28;
  reg [8:0] op2_06_in29;
  reg [8:0] op2_06_in30;
  reg [8:0] op2_06_bias;
  wire [8:0] op2_06_out;
  affine2_op2 op2_06(
    .data0_in(op2_06_in00),
    .data1_in(op2_06_in01),
    .data2_in(op2_06_in02),
    .data3_in(op2_06_in03),
    .data4_in(op2_06_in04),
    .data5_in(op2_06_in05),
    .data6_in(op2_06_in06),
    .data7_in(op2_06_in07),
    .data8_in(op2_06_in08),
    .data9_in(op2_06_in09),
    .data10_in(op2_06_in10),
    .data11_in(op2_06_in11),
    .data12_in(op2_06_in12),
    .data13_in(op2_06_in13),
    .data14_in(op2_06_in14),
    .data15_in(op2_06_in15),
    .data16_in(op2_06_in16),
    .data17_in(op2_06_in17),
    .data18_in(op2_06_in18),
    .data19_in(op2_06_in19),
    .data20_in(op2_06_in20),
    .data21_in(op2_06_in21),
    .data22_in(op2_06_in22),
    .data23_in(op2_06_in23),
    .data24_in(op2_06_in24),
    .data25_in(op2_06_in25),
    .data26_in(op2_06_in26),
    .data27_in(op2_06_in27),
    .data28_in(op2_06_in28),
    .data29_in(op2_06_in29),
    .data30_in(op2_06_in30),
    .data31_in(op2_06_bias),
    .data_out(op2_06_out));

  // 7 番目の OP2
  reg [8:0] op2_07_in00;
  reg [8:0] op2_07_in01;
  reg [8:0] op2_07_in02;
  reg [8:0] op2_07_in03;
  reg [8:0] op2_07_in04;
  reg [8:0] op2_07_in05;
  reg [8:0] op2_07_in06;
  reg [8:0] op2_07_in07;
  reg [8:0] op2_07_in08;
  reg [8:0] op2_07_in09;
  reg [8:0] op2_07_in10;
  reg [8:0] op2_07_in11;
  reg [8:0] op2_07_in12;
  reg [8:0] op2_07_in13;
  reg [8:0] op2_07_in14;
  reg [8:0] op2_07_in15;
  reg [8:0] op2_07_in16;
  reg [8:0] op2_07_in17;
  reg [8:0] op2_07_in18;
  reg [8:0] op2_07_in19;
  reg [8:0] op2_07_in20;
  reg [8:0] op2_07_in21;
  reg [8:0] op2_07_in22;
  reg [8:0] op2_07_in23;
  reg [8:0] op2_07_in24;
  reg [8:0] op2_07_in25;
  reg [8:0] op2_07_in26;
  reg [8:0] op2_07_in27;
  reg [8:0] op2_07_in28;
  reg [8:0] op2_07_in29;
  reg [8:0] op2_07_in30;
  reg [8:0] op2_07_bias;
  wire [8:0] op2_07_out;
  affine2_op2 op2_07(
    .data0_in(op2_07_in00),
    .data1_in(op2_07_in01),
    .data2_in(op2_07_in02),
    .data3_in(op2_07_in03),
    .data4_in(op2_07_in04),
    .data5_in(op2_07_in05),
    .data6_in(op2_07_in06),
    .data7_in(op2_07_in07),
    .data8_in(op2_07_in08),
    .data9_in(op2_07_in09),
    .data10_in(op2_07_in10),
    .data11_in(op2_07_in11),
    .data12_in(op2_07_in12),
    .data13_in(op2_07_in13),
    .data14_in(op2_07_in14),
    .data15_in(op2_07_in15),
    .data16_in(op2_07_in16),
    .data17_in(op2_07_in17),
    .data18_in(op2_07_in18),
    .data19_in(op2_07_in19),
    .data20_in(op2_07_in20),
    .data21_in(op2_07_in21),
    .data22_in(op2_07_in22),
    .data23_in(op2_07_in23),
    .data24_in(op2_07_in24),
    .data25_in(op2_07_in25),
    .data26_in(op2_07_in26),
    .data27_in(op2_07_in27),
    .data28_in(op2_07_in28),
    .data29_in(op2_07_in29),
    .data30_in(op2_07_in30),
    .data31_in(op2_07_bias),
    .data_out(op2_07_out));

  // 8 番目の OP2
  reg [8:0] op2_08_in00;
  reg [8:0] op2_08_in01;
  reg [8:0] op2_08_in02;
  reg [8:0] op2_08_in03;
  reg [8:0] op2_08_in04;
  reg [8:0] op2_08_in05;
  reg [8:0] op2_08_in06;
  reg [8:0] op2_08_in07;
  reg [8:0] op2_08_in08;
  reg [8:0] op2_08_in09;
  reg [8:0] op2_08_in10;
  reg [8:0] op2_08_in11;
  reg [8:0] op2_08_in12;
  reg [8:0] op2_08_in13;
  reg [8:0] op2_08_in14;
  reg [8:0] op2_08_in15;
  reg [8:0] op2_08_in16;
  reg [8:0] op2_08_in17;
  reg [8:0] op2_08_in18;
  reg [8:0] op2_08_in19;
  reg [8:0] op2_08_in20;
  reg [8:0] op2_08_in21;
  reg [8:0] op2_08_in22;
  reg [8:0] op2_08_in23;
  reg [8:0] op2_08_in24;
  reg [8:0] op2_08_in25;
  reg [8:0] op2_08_in26;
  reg [8:0] op2_08_in27;
  reg [8:0] op2_08_in28;
  reg [8:0] op2_08_in29;
  reg [8:0] op2_08_in30;
  reg [8:0] op2_08_bias;
  wire [8:0] op2_08_out;
  affine2_op2 op2_08(
    .data0_in(op2_08_in00),
    .data1_in(op2_08_in01),
    .data2_in(op2_08_in02),
    .data3_in(op2_08_in03),
    .data4_in(op2_08_in04),
    .data5_in(op2_08_in05),
    .data6_in(op2_08_in06),
    .data7_in(op2_08_in07),
    .data8_in(op2_08_in08),
    .data9_in(op2_08_in09),
    .data10_in(op2_08_in10),
    .data11_in(op2_08_in11),
    .data12_in(op2_08_in12),
    .data13_in(op2_08_in13),
    .data14_in(op2_08_in14),
    .data15_in(op2_08_in15),
    .data16_in(op2_08_in16),
    .data17_in(op2_08_in17),
    .data18_in(op2_08_in18),
    .data19_in(op2_08_in19),
    .data20_in(op2_08_in20),
    .data21_in(op2_08_in21),
    .data22_in(op2_08_in22),
    .data23_in(op2_08_in23),
    .data24_in(op2_08_in24),
    .data25_in(op2_08_in25),
    .data26_in(op2_08_in26),
    .data27_in(op2_08_in27),
    .data28_in(op2_08_in28),
    .data29_in(op2_08_in29),
    .data30_in(op2_08_in30),
    .data31_in(op2_08_bias),
    .data_out(op2_08_out));

  // 9 番目の OP2
  reg [8:0] op2_09_in00;
  reg [8:0] op2_09_in01;
  reg [8:0] op2_09_in02;
  reg [8:0] op2_09_in03;
  reg [8:0] op2_09_in04;
  reg [8:0] op2_09_in05;
  reg [8:0] op2_09_in06;
  reg [8:0] op2_09_in07;
  reg [8:0] op2_09_in08;
  reg [8:0] op2_09_in09;
  reg [8:0] op2_09_in10;
  reg [8:0] op2_09_in11;
  reg [8:0] op2_09_in12;
  reg [8:0] op2_09_in13;
  reg [8:0] op2_09_in14;
  reg [8:0] op2_09_in15;
  reg [8:0] op2_09_in16;
  reg [8:0] op2_09_in17;
  reg [8:0] op2_09_in18;
  reg [8:0] op2_09_in19;
  reg [8:0] op2_09_in20;
  reg [8:0] op2_09_in21;
  reg [8:0] op2_09_in22;
  reg [8:0] op2_09_in23;
  reg [8:0] op2_09_in24;
  reg [8:0] op2_09_in25;
  reg [8:0] op2_09_in26;
  reg [8:0] op2_09_in27;
  reg [8:0] op2_09_in28;
  reg [8:0] op2_09_in29;
  reg [8:0] op2_09_in30;
  reg [8:0] op2_09_bias;
  wire [8:0] op2_09_out;
  affine2_op2 op2_09(
    .data0_in(op2_09_in00),
    .data1_in(op2_09_in01),
    .data2_in(op2_09_in02),
    .data3_in(op2_09_in03),
    .data4_in(op2_09_in04),
    .data5_in(op2_09_in05),
    .data6_in(op2_09_in06),
    .data7_in(op2_09_in07),
    .data8_in(op2_09_in08),
    .data9_in(op2_09_in09),
    .data10_in(op2_09_in10),
    .data11_in(op2_09_in11),
    .data12_in(op2_09_in12),
    .data13_in(op2_09_in13),
    .data14_in(op2_09_in14),
    .data15_in(op2_09_in15),
    .data16_in(op2_09_in16),
    .data17_in(op2_09_in17),
    .data18_in(op2_09_in18),
    .data19_in(op2_09_in19),
    .data20_in(op2_09_in20),
    .data21_in(op2_09_in21),
    .data22_in(op2_09_in22),
    .data23_in(op2_09_in23),
    .data24_in(op2_09_in24),
    .data25_in(op2_09_in25),
    .data26_in(op2_09_in26),
    .data27_in(op2_09_in27),
    .data28_in(op2_09_in28),
    .data29_in(op2_09_in29),
    .data30_in(op2_09_in30),
    .data31_in(op2_09_bias),
    .data_out(op2_09_out));

  // 10 番目の OP2
  reg [8:0] op2_10_in00;
  reg [8:0] op2_10_in01;
  reg [8:0] op2_10_in02;
  reg [8:0] op2_10_in03;
  reg [8:0] op2_10_in04;
  reg [8:0] op2_10_in05;
  reg [8:0] op2_10_in06;
  reg [8:0] op2_10_in07;
  reg [8:0] op2_10_in08;
  reg [8:0] op2_10_in09;
  reg [8:0] op2_10_in10;
  reg [8:0] op2_10_in11;
  reg [8:0] op2_10_in12;
  reg [8:0] op2_10_in13;
  reg [8:0] op2_10_in14;
  reg [8:0] op2_10_in15;
  reg [8:0] op2_10_in16;
  reg [8:0] op2_10_in17;
  reg [8:0] op2_10_in18;
  reg [8:0] op2_10_in19;
  reg [8:0] op2_10_in20;
  reg [8:0] op2_10_in21;
  reg [8:0] op2_10_in22;
  reg [8:0] op2_10_in23;
  reg [8:0] op2_10_in24;
  reg [8:0] op2_10_in25;
  reg [8:0] op2_10_in26;
  reg [8:0] op2_10_in27;
  reg [8:0] op2_10_in28;
  reg [8:0] op2_10_in29;
  reg [8:0] op2_10_in30;
  reg [8:0] op2_10_bias;
  wire [8:0] op2_10_out;
  affine2_op2 op2_10(
    .data0_in(op2_10_in00),
    .data1_in(op2_10_in01),
    .data2_in(op2_10_in02),
    .data3_in(op2_10_in03),
    .data4_in(op2_10_in04),
    .data5_in(op2_10_in05),
    .data6_in(op2_10_in06),
    .data7_in(op2_10_in07),
    .data8_in(op2_10_in08),
    .data9_in(op2_10_in09),
    .data10_in(op2_10_in10),
    .data11_in(op2_10_in11),
    .data12_in(op2_10_in12),
    .data13_in(op2_10_in13),
    .data14_in(op2_10_in14),
    .data15_in(op2_10_in15),
    .data16_in(op2_10_in16),
    .data17_in(op2_10_in17),
    .data18_in(op2_10_in18),
    .data19_in(op2_10_in19),
    .data20_in(op2_10_in20),
    .data21_in(op2_10_in21),
    .data22_in(op2_10_in22),
    .data23_in(op2_10_in23),
    .data24_in(op2_10_in24),
    .data25_in(op2_10_in25),
    .data26_in(op2_10_in26),
    .data27_in(op2_10_in27),
    .data28_in(op2_10_in28),
    .data29_in(op2_10_in29),
    .data30_in(op2_10_in30),
    .data31_in(op2_10_bias),
    .data_out(op2_10_out));

  // 11 番目の OP2
  reg [8:0] op2_11_in00;
  reg [8:0] op2_11_in01;
  reg [8:0] op2_11_in02;
  reg [8:0] op2_11_in03;
  reg [8:0] op2_11_in04;
  reg [8:0] op2_11_in05;
  reg [8:0] op2_11_in06;
  reg [8:0] op2_11_in07;
  reg [8:0] op2_11_in08;
  reg [8:0] op2_11_in09;
  reg [8:0] op2_11_in10;
  reg [8:0] op2_11_in11;
  reg [8:0] op2_11_in12;
  reg [8:0] op2_11_in13;
  reg [8:0] op2_11_in14;
  reg [8:0] op2_11_in15;
  reg [8:0] op2_11_in16;
  reg [8:0] op2_11_in17;
  reg [8:0] op2_11_in18;
  reg [8:0] op2_11_in19;
  reg [8:0] op2_11_in20;
  reg [8:0] op2_11_in21;
  reg [8:0] op2_11_in22;
  reg [8:0] op2_11_in23;
  reg [8:0] op2_11_in24;
  reg [8:0] op2_11_in25;
  reg [8:0] op2_11_in26;
  reg [8:0] op2_11_in27;
  reg [8:0] op2_11_in28;
  reg [8:0] op2_11_in29;
  reg [8:0] op2_11_in30;
  reg [8:0] op2_11_bias;
  wire [8:0] op2_11_out;
  affine2_op2 op2_11(
    .data0_in(op2_11_in00),
    .data1_in(op2_11_in01),
    .data2_in(op2_11_in02),
    .data3_in(op2_11_in03),
    .data4_in(op2_11_in04),
    .data5_in(op2_11_in05),
    .data6_in(op2_11_in06),
    .data7_in(op2_11_in07),
    .data8_in(op2_11_in08),
    .data9_in(op2_11_in09),
    .data10_in(op2_11_in10),
    .data11_in(op2_11_in11),
    .data12_in(op2_11_in12),
    .data13_in(op2_11_in13),
    .data14_in(op2_11_in14),
    .data15_in(op2_11_in15),
    .data16_in(op2_11_in16),
    .data17_in(op2_11_in17),
    .data18_in(op2_11_in18),
    .data19_in(op2_11_in19),
    .data20_in(op2_11_in20),
    .data21_in(op2_11_in21),
    .data22_in(op2_11_in22),
    .data23_in(op2_11_in23),
    .data24_in(op2_11_in24),
    .data25_in(op2_11_in25),
    .data26_in(op2_11_in26),
    .data27_in(op2_11_in27),
    .data28_in(op2_11_in28),
    .data29_in(op2_11_in29),
    .data30_in(op2_11_in30),
    .data31_in(op2_11_bias),
    .data_out(op2_11_out));

  // 12 番目の OP2
  reg [8:0] op2_12_in00;
  reg [8:0] op2_12_in01;
  reg [8:0] op2_12_in02;
  reg [8:0] op2_12_in03;
  reg [8:0] op2_12_in04;
  reg [8:0] op2_12_in05;
  reg [8:0] op2_12_in06;
  reg [8:0] op2_12_in07;
  reg [8:0] op2_12_in08;
  reg [8:0] op2_12_in09;
  reg [8:0] op2_12_in10;
  reg [8:0] op2_12_in11;
  reg [8:0] op2_12_in12;
  reg [8:0] op2_12_in13;
  reg [8:0] op2_12_in14;
  reg [8:0] op2_12_in15;
  reg [8:0] op2_12_in16;
  reg [8:0] op2_12_in17;
  reg [8:0] op2_12_in18;
  reg [8:0] op2_12_in19;
  reg [8:0] op2_12_in20;
  reg [8:0] op2_12_in21;
  reg [8:0] op2_12_in22;
  reg [8:0] op2_12_in23;
  reg [8:0] op2_12_in24;
  reg [8:0] op2_12_in25;
  reg [8:0] op2_12_in26;
  reg [8:0] op2_12_in27;
  reg [8:0] op2_12_in28;
  reg [8:0] op2_12_in29;
  reg [8:0] op2_12_in30;
  reg [8:0] op2_12_bias;
  wire [8:0] op2_12_out;
  affine2_op2 op2_12(
    .data0_in(op2_12_in00),
    .data1_in(op2_12_in01),
    .data2_in(op2_12_in02),
    .data3_in(op2_12_in03),
    .data4_in(op2_12_in04),
    .data5_in(op2_12_in05),
    .data6_in(op2_12_in06),
    .data7_in(op2_12_in07),
    .data8_in(op2_12_in08),
    .data9_in(op2_12_in09),
    .data10_in(op2_12_in10),
    .data11_in(op2_12_in11),
    .data12_in(op2_12_in12),
    .data13_in(op2_12_in13),
    .data14_in(op2_12_in14),
    .data15_in(op2_12_in15),
    .data16_in(op2_12_in16),
    .data17_in(op2_12_in17),
    .data18_in(op2_12_in18),
    .data19_in(op2_12_in19),
    .data20_in(op2_12_in20),
    .data21_in(op2_12_in21),
    .data22_in(op2_12_in22),
    .data23_in(op2_12_in23),
    .data24_in(op2_12_in24),
    .data25_in(op2_12_in25),
    .data26_in(op2_12_in26),
    .data27_in(op2_12_in27),
    .data28_in(op2_12_in28),
    .data29_in(op2_12_in29),
    .data30_in(op2_12_in30),
    .data31_in(op2_12_bias),
    .data_out(op2_12_out));

  // 13 番目の OP2
  reg [8:0] op2_13_in00;
  reg [8:0] op2_13_in01;
  reg [8:0] op2_13_in02;
  reg [8:0] op2_13_in03;
  reg [8:0] op2_13_in04;
  reg [8:0] op2_13_in05;
  reg [8:0] op2_13_in06;
  reg [8:0] op2_13_in07;
  reg [8:0] op2_13_in08;
  reg [8:0] op2_13_in09;
  reg [8:0] op2_13_in10;
  reg [8:0] op2_13_in11;
  reg [8:0] op2_13_in12;
  reg [8:0] op2_13_in13;
  reg [8:0] op2_13_in14;
  reg [8:0] op2_13_in15;
  reg [8:0] op2_13_in16;
  reg [8:0] op2_13_in17;
  reg [8:0] op2_13_in18;
  reg [8:0] op2_13_in19;
  reg [8:0] op2_13_in20;
  reg [8:0] op2_13_in21;
  reg [8:0] op2_13_in22;
  reg [8:0] op2_13_in23;
  reg [8:0] op2_13_in24;
  reg [8:0] op2_13_in25;
  reg [8:0] op2_13_in26;
  reg [8:0] op2_13_in27;
  reg [8:0] op2_13_in28;
  reg [8:0] op2_13_in29;
  reg [8:0] op2_13_in30;
  reg [8:0] op2_13_bias;
  wire [8:0] op2_13_out;
  affine2_op2 op2_13(
    .data0_in(op2_13_in00),
    .data1_in(op2_13_in01),
    .data2_in(op2_13_in02),
    .data3_in(op2_13_in03),
    .data4_in(op2_13_in04),
    .data5_in(op2_13_in05),
    .data6_in(op2_13_in06),
    .data7_in(op2_13_in07),
    .data8_in(op2_13_in08),
    .data9_in(op2_13_in09),
    .data10_in(op2_13_in10),
    .data11_in(op2_13_in11),
    .data12_in(op2_13_in12),
    .data13_in(op2_13_in13),
    .data14_in(op2_13_in14),
    .data15_in(op2_13_in15),
    .data16_in(op2_13_in16),
    .data17_in(op2_13_in17),
    .data18_in(op2_13_in18),
    .data19_in(op2_13_in19),
    .data20_in(op2_13_in20),
    .data21_in(op2_13_in21),
    .data22_in(op2_13_in22),
    .data23_in(op2_13_in23),
    .data24_in(op2_13_in24),
    .data25_in(op2_13_in25),
    .data26_in(op2_13_in26),
    .data27_in(op2_13_in27),
    .data28_in(op2_13_in28),
    .data29_in(op2_13_in29),
    .data30_in(op2_13_in30),
    .data31_in(op2_13_bias),
    .data_out(op2_13_out));

  // 14 番目の OP2
  reg [8:0] op2_14_in00;
  reg [8:0] op2_14_in01;
  reg [8:0] op2_14_in02;
  reg [8:0] op2_14_in03;
  reg [8:0] op2_14_in04;
  reg [8:0] op2_14_in05;
  reg [8:0] op2_14_in06;
  reg [8:0] op2_14_in07;
  reg [8:0] op2_14_in08;
  reg [8:0] op2_14_in09;
  reg [8:0] op2_14_in10;
  reg [8:0] op2_14_in11;
  reg [8:0] op2_14_in12;
  reg [8:0] op2_14_in13;
  reg [8:0] op2_14_in14;
  reg [8:0] op2_14_in15;
  reg [8:0] op2_14_in16;
  reg [8:0] op2_14_in17;
  reg [8:0] op2_14_in18;
  reg [8:0] op2_14_in19;
  reg [8:0] op2_14_in20;
  reg [8:0] op2_14_in21;
  reg [8:0] op2_14_in22;
  reg [8:0] op2_14_in23;
  reg [8:0] op2_14_in24;
  reg [8:0] op2_14_in25;
  reg [8:0] op2_14_in26;
  reg [8:0] op2_14_in27;
  reg [8:0] op2_14_in28;
  reg [8:0] op2_14_in29;
  reg [8:0] op2_14_in30;
  reg [8:0] op2_14_bias;
  wire [8:0] op2_14_out;
  affine2_op2 op2_14(
    .data0_in(op2_14_in00),
    .data1_in(op2_14_in01),
    .data2_in(op2_14_in02),
    .data3_in(op2_14_in03),
    .data4_in(op2_14_in04),
    .data5_in(op2_14_in05),
    .data6_in(op2_14_in06),
    .data7_in(op2_14_in07),
    .data8_in(op2_14_in08),
    .data9_in(op2_14_in09),
    .data10_in(op2_14_in10),
    .data11_in(op2_14_in11),
    .data12_in(op2_14_in12),
    .data13_in(op2_14_in13),
    .data14_in(op2_14_in14),
    .data15_in(op2_14_in15),
    .data16_in(op2_14_in16),
    .data17_in(op2_14_in17),
    .data18_in(op2_14_in18),
    .data19_in(op2_14_in19),
    .data20_in(op2_14_in20),
    .data21_in(op2_14_in21),
    .data22_in(op2_14_in22),
    .data23_in(op2_14_in23),
    .data24_in(op2_14_in24),
    .data25_in(op2_14_in25),
    .data26_in(op2_14_in26),
    .data27_in(op2_14_in27),
    .data28_in(op2_14_in28),
    .data29_in(op2_14_in29),
    .data30_in(op2_14_in30),
    .data31_in(op2_14_bias),
    .data_out(op2_14_out));

  // 15 番目の OP2
  reg [8:0] op2_15_in00;
  reg [8:0] op2_15_in01;
  reg [8:0] op2_15_in02;
  reg [8:0] op2_15_in03;
  reg [8:0] op2_15_in04;
  reg [8:0] op2_15_in05;
  reg [8:0] op2_15_in06;
  reg [8:0] op2_15_in07;
  reg [8:0] op2_15_in08;
  reg [8:0] op2_15_in09;
  reg [8:0] op2_15_in10;
  reg [8:0] op2_15_in11;
  reg [8:0] op2_15_in12;
  reg [8:0] op2_15_in13;
  reg [8:0] op2_15_in14;
  reg [8:0] op2_15_in15;
  reg [8:0] op2_15_in16;
  reg [8:0] op2_15_in17;
  reg [8:0] op2_15_in18;
  reg [8:0] op2_15_in19;
  reg [8:0] op2_15_in20;
  reg [8:0] op2_15_in21;
  reg [8:0] op2_15_in22;
  reg [8:0] op2_15_in23;
  reg [8:0] op2_15_in24;
  reg [8:0] op2_15_in25;
  reg [8:0] op2_15_in26;
  reg [8:0] op2_15_in27;
  reg [8:0] op2_15_in28;
  reg [8:0] op2_15_in29;
  reg [8:0] op2_15_in30;
  reg [8:0] op2_15_bias;
  wire [8:0] op2_15_out;
  affine2_op2 op2_15(
    .data0_in(op2_15_in00),
    .data1_in(op2_15_in01),
    .data2_in(op2_15_in02),
    .data3_in(op2_15_in03),
    .data4_in(op2_15_in04),
    .data5_in(op2_15_in05),
    .data6_in(op2_15_in06),
    .data7_in(op2_15_in07),
    .data8_in(op2_15_in08),
    .data9_in(op2_15_in09),
    .data10_in(op2_15_in10),
    .data11_in(op2_15_in11),
    .data12_in(op2_15_in12),
    .data13_in(op2_15_in13),
    .data14_in(op2_15_in14),
    .data15_in(op2_15_in15),
    .data16_in(op2_15_in16),
    .data17_in(op2_15_in17),
    .data18_in(op2_15_in18),
    .data19_in(op2_15_in19),
    .data20_in(op2_15_in20),
    .data21_in(op2_15_in21),
    .data22_in(op2_15_in22),
    .data23_in(op2_15_in23),
    .data24_in(op2_15_in24),
    .data25_in(op2_15_in25),
    .data26_in(op2_15_in26),
    .data27_in(op2_15_in27),
    .data28_in(op2_15_in28),
    .data29_in(op2_15_in29),
    .data30_in(op2_15_in30),
    .data31_in(op2_15_bias),
    .data_out(op2_15_out));

  // 中間レジスタ
  reg [8:0] reg_0000;
  reg [8:0] reg_0001;
  reg [8:0] reg_0002;
  reg [8:0] reg_0003;
  reg [8:0] reg_0004;
  reg [8:0] reg_0005;
  reg [8:0] reg_0006;
  reg [8:0] reg_0007;
  reg [8:0] reg_0008;
  reg [8:0] reg_0009;
  reg [8:0] reg_0010;
  reg [8:0] reg_0011;
  reg [8:0] reg_0012;
  reg [8:0] reg_0013;
  reg [8:0] reg_0014;
  reg [8:0] reg_0015;
  reg [8:0] reg_0016;
  reg [8:0] reg_0017;
  reg [8:0] reg_0018;
  reg [8:0] reg_0019;
  reg [8:0] reg_0020;
  reg [8:0] reg_0021;
  reg [8:0] reg_0022;
  reg [8:0] reg_0023;
  reg [8:0] reg_0024;
  reg [8:0] reg_0025;
  reg [8:0] reg_0026;
  reg [8:0] reg_0027;
  reg [8:0] reg_0028;
  reg [8:0] reg_0029;
  reg [8:0] reg_0030;
  reg [8:0] reg_0031;
  reg [8:0] reg_0032;
  reg [8:0] reg_0033;
  reg [8:0] reg_0034;
  reg [8:0] reg_0035;
  reg [8:0] reg_0036;
  reg [8:0] reg_0037;
  reg [8:0] reg_0038;
  reg [8:0] reg_0039;
  reg [8:0] reg_0040;
  reg [8:0] reg_0041;
  reg [8:0] reg_0042;
  reg [8:0] reg_0043;
  reg [8:0] reg_0044;
  reg [8:0] reg_0045;
  reg [8:0] reg_0046;
  reg [8:0] reg_0047;
  reg [8:0] reg_0048;
  reg [8:0] reg_0049;
  reg [8:0] reg_0050;
  reg [8:0] reg_0051;
  reg [8:0] reg_0052;
  reg [8:0] reg_0053;
  reg [8:0] reg_0054;
  reg [8:0] reg_0055;
  reg [8:0] reg_0056;
  reg [8:0] reg_0057;
  reg [8:0] reg_0058;
  reg [8:0] reg_0059;
  reg [8:0] reg_0060;
  reg [8:0] reg_0061;
  reg [8:0] reg_0062;
  reg [8:0] reg_0063;
  reg [8:0] reg_0064;
  reg [8:0] reg_0065;
  reg [8:0] reg_0066;
  reg [8:0] reg_0067;
  reg [8:0] reg_0068;
  reg [8:0] reg_0069;
  reg [8:0] reg_0070;
  reg [8:0] reg_0071;
  reg [8:0] reg_0072;
  reg [8:0] reg_0073;
  reg [8:0] reg_0074;
  reg [8:0] reg_0075;
  reg [8:0] reg_0076;
  reg [8:0] reg_0077;
  reg [8:0] reg_0078;
  reg [8:0] reg_0079;
  reg [8:0] reg_0080;
  reg [8:0] reg_0081;
  reg [8:0] reg_0082;
  reg [8:0] reg_0083;
  reg [8:0] reg_0084;
  reg [8:0] reg_0085;
  reg [8:0] reg_0086;
  reg [8:0] reg_0087;
  reg [8:0] reg_0088;
  reg [8:0] reg_0089;
  reg [8:0] reg_0090;
  reg [8:0] reg_0091;
  reg [8:0] reg_0092;
  reg [8:0] reg_0093;
  reg [8:0] reg_0094;
  reg [8:0] reg_0095;
  reg [8:0] reg_0096;
  reg [8:0] reg_0097;
  reg [8:0] reg_0098;
  reg [8:0] reg_0099;
  reg [8:0] reg_0100;
  reg [8:0] reg_0101;
  reg [8:0] reg_0102;
  reg [8:0] reg_0103;
  reg [8:0] reg_0104;
  reg [8:0] reg_0105;
  reg [8:0] reg_0106;
  reg [8:0] reg_0107;
  reg [8:0] reg_0108;
  reg [8:0] reg_0109;
  reg [8:0] reg_0110;
  reg [8:0] reg_0111;
  reg [8:0] reg_0112;
  reg [8:0] reg_0113;
  reg [8:0] reg_0114;
  reg [8:0] reg_0115;
  reg [8:0] reg_0116;
  reg [8:0] reg_0117;
  reg [8:0] reg_0118;
  reg [8:0] reg_0119;
  reg [8:0] reg_0120;
  reg [8:0] reg_0121;
  reg [8:0] reg_0122;
  reg [8:0] reg_0123;
  reg [8:0] reg_0124;
  reg [8:0] reg_0125;
  reg [8:0] reg_0126;
  reg [8:0] reg_0127;
  reg [8:0] reg_0128;
  reg [8:0] reg_0129;
  reg [8:0] reg_0130;
  reg [8:0] reg_0131;
  reg [8:0] reg_0132;
  reg [8:0] reg_0133;
  reg [8:0] reg_0134;
  reg [8:0] reg_0135;
  reg [8:0] reg_0136;
  reg [8:0] reg_0137;
  reg [8:0] reg_0138;
  reg [8:0] reg_0139;
  reg [8:0] reg_0140;
  reg [8:0] reg_0141;
  reg [8:0] reg_0142;
  reg [8:0] reg_0143;
  reg [8:0] reg_0144;
  reg [8:0] reg_0145;
  reg [8:0] reg_0146;
  reg [8:0] reg_0147;
  reg [8:0] reg_0148;
  reg [8:0] reg_0149;
  reg [8:0] reg_0150;
  reg [8:0] reg_0151;
  reg [8:0] reg_0152;
  reg [8:0] reg_0153;
  reg [8:0] reg_0154;
  reg [8:0] reg_0155;
  reg [8:0] reg_0156;
  reg [8:0] reg_0157;
  reg [8:0] reg_0158;
  reg [8:0] reg_0159;
  reg [8:0] reg_0160;
  reg [8:0] reg_0161;
  reg [8:0] reg_0162;
  reg [8:0] reg_0163;
  reg [8:0] reg_0164;
  reg [8:0] reg_0165;
  reg [8:0] reg_0166;
  reg [8:0] reg_0167;
  reg [8:0] reg_0168;
  reg [8:0] reg_0169;
  reg [8:0] reg_0170;
  reg [8:0] reg_0171;
  reg [8:0] reg_0172;
  reg [8:0] reg_0173;
  reg [8:0] reg_0174;
  reg [8:0] reg_0175;
  reg [8:0] reg_0176;
  reg [8:0] reg_0177;
  reg [8:0] reg_0178;
  reg [8:0] reg_0179;
  reg [8:0] reg_0180;
  reg [8:0] reg_0181;
  reg [8:0] reg_0182;
  reg [8:0] reg_0183;
  reg [8:0] reg_0184;
  reg [8:0] reg_0185;
  reg [8:0] reg_0186;
  reg [8:0] reg_0187;
  reg [8:0] reg_0188;
  reg [8:0] reg_0189;
  reg [8:0] reg_0190;
  reg [8:0] reg_0191;
  reg [8:0] reg_0192;
  reg [8:0] reg_0193;
  reg [8:0] reg_0194;
  reg [8:0] reg_0195;
  reg [8:0] reg_0196;
  reg [8:0] reg_0197;
  reg [8:0] reg_0198;
  reg [8:0] reg_0199;
  reg [8:0] reg_0200;
  reg [8:0] reg_0201;
  reg [8:0] reg_0202;
  reg [8:0] reg_0203;
  reg [8:0] reg_0204;
  reg [8:0] reg_0205;
  reg [8:0] reg_0206;
  reg [8:0] reg_0207;
  reg [8:0] reg_0208;
  reg [8:0] reg_0209;
  reg [8:0] reg_0210;
  reg [8:0] reg_0211;
  reg [8:0] reg_0212;
  reg [8:0] reg_0213;
  reg [8:0] reg_0214;
  reg [8:0] reg_0215;
  reg [8:0] reg_0216;
  reg [8:0] reg_0217;
  reg [8:0] reg_0218;
  reg [8:0] reg_0219;
  reg [8:0] reg_0220;
  reg [8:0] reg_0221;
  reg [8:0] reg_0222;
  reg [8:0] reg_0223;
  reg [8:0] reg_0224;
  reg [8:0] reg_0225;
  reg [8:0] reg_0226;
  reg [8:0] reg_0227;
  reg [8:0] reg_0228;
  reg [8:0] reg_0229;
  reg [8:0] reg_0230;
  reg [8:0] reg_0231;
  reg [8:0] reg_0232;
  reg [8:0] reg_0233;
  reg [8:0] reg_0234;
  reg [8:0] reg_0235;
  reg [8:0] reg_0236;
  reg [8:0] reg_0237;
  reg [8:0] reg_0238;
  reg [8:0] reg_0239;
  reg [8:0] reg_0240;
  reg [8:0] reg_0241;
  reg [8:0] reg_0242;
  reg [8:0] reg_0243;
  reg [8:0] reg_0244;
  reg [8:0] reg_0245;
  reg [8:0] reg_0246;
  reg [8:0] reg_0247;
  reg [8:0] reg_0248;
  reg [8:0] reg_0249;
  reg [8:0] reg_0250;
  reg [8:0] reg_0251;
  reg [8:0] reg_0252;
  reg [8:0] reg_0253;
  reg [8:0] reg_0254;
  reg [8:0] reg_0255;
  reg [8:0] reg_0256;
  reg [8:0] reg_0257;
  reg [8:0] reg_0258;
  reg [8:0] reg_0259;
  reg [8:0] reg_0260;
  reg [8:0] reg_0261;
  reg [8:0] reg_0262;
  reg [8:0] reg_0263;
  reg [8:0] reg_0264;
  reg [8:0] reg_0265;
  reg [8:0] reg_0266;
  reg [8:0] reg_0267;
  reg [8:0] reg_0268;
  reg [8:0] reg_0269;
  reg [8:0] reg_0270;
  reg [8:0] reg_0271;
  reg [8:0] reg_0272;
  reg [8:0] reg_0273;
  reg [8:0] reg_0274;
  reg [8:0] reg_0275;
  reg [8:0] reg_0276;
  reg [8:0] reg_0277;
  reg [8:0] reg_0278;
  reg [8:0] reg_0279;
  reg [8:0] reg_0280;
  reg [8:0] reg_0281;
  reg [8:0] reg_0282;
  reg [8:0] reg_0283;
  reg [8:0] reg_0284;
  reg [8:0] reg_0285;
  reg [8:0] reg_0286;
  reg [8:0] reg_0287;
  reg [8:0] reg_0288;
  reg [8:0] reg_0289;
  reg [8:0] reg_0290;
  reg [8:0] reg_0291;
  reg [8:0] reg_0292;
  reg [8:0] reg_0293;
  reg [8:0] reg_0294;
  reg [8:0] reg_0295;
  reg [8:0] reg_0296;
  reg [8:0] reg_0297;
  reg [8:0] reg_0298;
  reg [8:0] reg_0299;
  reg [8:0] reg_0300;
  reg [8:0] reg_0301;
  reg [8:0] reg_0302;
  reg [8:0] reg_0303;
  reg [8:0] reg_0304;
  reg [8:0] reg_0305;
  reg [8:0] reg_0306;
  reg [8:0] reg_0307;
  reg [8:0] reg_0308;
  reg [8:0] reg_0309;
  reg [8:0] reg_0310;
  reg [8:0] reg_0311;
  reg [8:0] reg_0312;
  reg [8:0] reg_0313;
  reg [8:0] reg_0314;
  reg [8:0] reg_0315;
  reg [8:0] reg_0316;
  reg [8:0] reg_0317;
  reg [8:0] reg_0318;
  reg [8:0] reg_0319;
  reg [8:0] reg_0320;
  reg [8:0] reg_0321;
  reg [8:0] reg_0322;
  reg [8:0] reg_0323;
  reg [8:0] reg_0324;
  reg [8:0] reg_0325;
  reg [8:0] reg_0326;
  reg [8:0] reg_0327;
  reg [8:0] reg_0328;
  reg [8:0] reg_0329;
  reg [8:0] reg_0330;
  reg [8:0] reg_0331;
  reg [8:0] reg_0332;
  reg [8:0] reg_0333;
  reg [8:0] reg_0334;
  reg [8:0] reg_0335;
  reg [8:0] reg_0336;
  reg [8:0] reg_0337;
  reg [8:0] reg_0338;
  reg [8:0] reg_0339;
  reg [8:0] reg_0340;
  reg [8:0] reg_0341;
  reg [8:0] reg_0342;
  reg [8:0] reg_0343;
  reg [8:0] reg_0344;
  reg [8:0] reg_0345;
  reg [8:0] reg_0346;
  reg [8:0] reg_0347;
  reg [8:0] reg_0348;
  reg [8:0] reg_0349;
  reg [8:0] reg_0350;
  reg [8:0] reg_0351;
  reg [8:0] reg_0352;
  reg [8:0] reg_0353;
  reg [8:0] reg_0354;
  reg [8:0] reg_0355;
  reg [8:0] reg_0356;
  reg [8:0] reg_0357;
  reg [8:0] reg_0358;
  reg [8:0] reg_0359;
  reg [8:0] reg_0360;
  reg [8:0] reg_0361;
  reg [8:0] reg_0362;
  reg [8:0] reg_0363;
  reg [8:0] reg_0364;
  reg [8:0] reg_0365;
  reg [8:0] reg_0366;
  reg [8:0] reg_0367;
  reg [8:0] reg_0368;
  reg [8:0] reg_0369;
  reg [8:0] reg_0370;
  reg [8:0] reg_0371;
  reg [8:0] reg_0372;
  reg [8:0] reg_0373;
  reg [8:0] reg_0374;
  reg [8:0] reg_0375;
  reg [8:0] reg_0376;
  reg [8:0] reg_0377;
  reg [8:0] reg_0378;
  reg [8:0] reg_0379;
  reg [8:0] reg_0380;
  reg [8:0] reg_0381;
  reg [8:0] reg_0382;
  reg [8:0] reg_0383;
  reg [8:0] reg_0384;
  reg [8:0] reg_0385;
  reg [8:0] reg_0386;
  reg [8:0] reg_0387;
  reg [8:0] reg_0388;
  reg [8:0] reg_0389;
  reg [8:0] reg_0390;
  reg [8:0] reg_0391;
  reg [8:0] reg_0392;
  reg [8:0] reg_0393;
  reg [8:0] reg_0394;
  reg [8:0] reg_0395;
  reg [8:0] reg_0396;
  reg [8:0] reg_0397;
  reg [8:0] reg_0398;
  reg [8:0] reg_0399;
  reg [8:0] reg_0400;
  reg [8:0] reg_0401;
  reg [8:0] reg_0402;
  reg [8:0] reg_0403;
  reg [8:0] reg_0404;
  reg [8:0] reg_0405;
  reg [8:0] reg_0406;
  reg [8:0] reg_0407;
  reg [8:0] reg_0408;
  reg [8:0] reg_0409;
  reg [8:0] reg_0410;
  reg [8:0] reg_0411;
  reg [8:0] reg_0412;
  reg [8:0] reg_0413;
  reg [8:0] reg_0414;
  reg [8:0] reg_0415;
  reg [8:0] reg_0416;
  reg [8:0] reg_0417;
  reg [8:0] reg_0418;
  reg [8:0] reg_0419;
  reg [8:0] reg_0420;
  reg [8:0] reg_0421;
  reg [8:0] reg_0422;
  reg [8:0] reg_0423;
  reg [8:0] reg_0424;
  reg [8:0] reg_0425;
  reg [8:0] reg_0426;
  reg [8:0] reg_0427;
  reg [8:0] reg_0428;
  reg [8:0] reg_0429;
  reg [8:0] reg_0430;
  reg [8:0] reg_0431;
  reg [8:0] reg_0432;
  reg [8:0] reg_0433;
  reg [8:0] reg_0434;
  reg [8:0] reg_0435;
  reg [8:0] reg_0436;
  reg [8:0] reg_0437;
  reg [8:0] reg_0438;
  reg [8:0] reg_0439;
  reg [8:0] reg_0440;
  reg [8:0] reg_0441;
  reg [8:0] reg_0442;
  reg [8:0] reg_0443;
  reg [8:0] reg_0444;
  reg [8:0] reg_0445;
  reg [8:0] reg_0446;
  reg [8:0] reg_0447;
  reg [8:0] reg_0448;
  reg [8:0] reg_0449;
  reg [8:0] reg_0450;
  reg [8:0] reg_0451;
  reg [8:0] reg_0452;
  reg [8:0] reg_0453;
  reg [8:0] reg_0454;
  reg [8:0] reg_0455;
  reg [8:0] reg_0456;
  reg [8:0] reg_0457;
  reg [8:0] reg_0458;
  reg [8:0] reg_0459;
  reg [8:0] reg_0460;
  reg [8:0] reg_0461;
  reg [8:0] reg_0462;
  reg [8:0] reg_0463;
  reg [8:0] reg_0464;
  reg [8:0] reg_0465;
  reg [8:0] reg_0466;
  reg [8:0] reg_0467;
  reg [8:0] reg_0468;
  reg [8:0] reg_0469;
  reg [8:0] reg_0470;
  reg [8:0] reg_0471;
  reg [8:0] reg_0472;
  reg [8:0] reg_0473;
  reg [8:0] reg_0474;
  reg [8:0] reg_0475;
  reg [8:0] reg_0476;
  reg [8:0] reg_0477;
  reg [8:0] reg_0478;
  reg [8:0] reg_0479;
  reg [8:0] reg_0480;
  reg [8:0] reg_0481;
  reg [8:0] reg_0482;
  reg [8:0] reg_0483;
  reg [8:0] reg_0484;
  reg [8:0] reg_0485;
  reg [8:0] reg_0486;
  reg [8:0] reg_0487;
  reg [8:0] reg_0488;
  reg [8:0] reg_0489;
  reg [8:0] reg_0490;
  reg [8:0] reg_0491;
  reg [8:0] reg_0492;
  reg [8:0] reg_0493;
  reg [8:0] reg_0494;
  reg [8:0] reg_0495;
  reg [8:0] reg_0496;
  reg [8:0] reg_0497;
  reg [8:0] reg_0498;
  reg [8:0] reg_0499;
  reg [8:0] reg_0500;
  reg [8:0] reg_0501;
  reg [8:0] reg_0502;
  reg [8:0] reg_0503;
  reg [8:0] reg_0504;
  reg [8:0] reg_0505;
  reg [8:0] reg_0506;
  reg [8:0] reg_0507;
  reg [8:0] reg_0508;
  reg [8:0] reg_0509;
  reg [8:0] reg_0510;
  reg [8:0] reg_0511;
  reg [8:0] reg_0512;
  reg [8:0] reg_0513;
  reg [8:0] reg_0514;
  reg [8:0] reg_0515;
  reg [8:0] reg_0516;
  reg [8:0] reg_0517;
  reg [8:0] reg_0518;
  reg [8:0] reg_0519;
  reg [8:0] reg_0520;
  reg [8:0] reg_0521;
  reg [8:0] reg_0522;
  reg [8:0] reg_0523;
  reg [8:0] reg_0524;
  reg [8:0] reg_0525;
  reg [8:0] reg_0526;
  reg [8:0] reg_0527;
  reg [8:0] reg_0528;
  reg [8:0] reg_0529;
  reg [8:0] reg_0530;
  reg [8:0] reg_0531;
  reg [8:0] reg_0532;
  reg [8:0] reg_0533;
  reg [8:0] reg_0534;
  reg [8:0] reg_0535;
  reg [8:0] reg_0536;
  reg [8:0] reg_0537;
  reg [8:0] reg_0538;
  reg [8:0] reg_0539;
  reg [8:0] reg_0540;
  reg [8:0] reg_0541;
  reg [8:0] reg_0542;
  reg [8:0] reg_0543;
  reg [8:0] reg_0544;
  reg [8:0] reg_0545;
  reg [8:0] reg_0546;
  reg [8:0] reg_0547;
  reg [8:0] reg_0548;
  reg [8:0] reg_0549;
  reg [8:0] reg_0550;
  reg [8:0] reg_0551;
  reg [8:0] reg_0552;
  reg [8:0] reg_0553;
  reg [8:0] reg_0554;
  reg [8:0] reg_0555;
  reg [8:0] reg_0556;
  reg [8:0] reg_0557;
  reg [8:0] reg_0558;
  reg [8:0] reg_0559;
  reg [8:0] reg_0560;
  reg [8:0] reg_0561;
  reg [8:0] reg_0562;
  reg [8:0] reg_0563;
  reg [8:0] reg_0564;
  reg [8:0] reg_0565;
  reg [8:0] reg_0566;
  reg [8:0] reg_0567;
  reg [8:0] reg_0568;
  reg [8:0] reg_0569;
  reg [8:0] reg_0570;
  reg [8:0] reg_0571;
  reg [8:0] reg_0572;
  reg [8:0] reg_0573;
  reg [8:0] reg_0574;
  reg [8:0] reg_0575;
  reg [8:0] reg_0576;
  reg [8:0] reg_0577;
  reg [8:0] reg_0578;
  reg [8:0] reg_0579;
  reg [8:0] reg_0580;
  reg [8:0] reg_0581;
  reg [8:0] reg_0582;
  reg [8:0] reg_0583;
  reg [8:0] reg_0584;
  reg [8:0] reg_0585;
  reg [8:0] reg_0586;
  reg [8:0] reg_0587;
  reg [8:0] reg_0588;
  reg [8:0] reg_0589;
  reg [8:0] reg_0590;
  reg [8:0] reg_0591;
  reg [8:0] reg_0592;
  reg [8:0] reg_0593;
  reg [8:0] reg_0594;
  reg [8:0] reg_0595;
  reg [8:0] reg_0596;
  reg [8:0] reg_0597;
  reg [8:0] reg_0598;
  reg [8:0] reg_0599;
  reg [8:0] reg_0600;
  reg [8:0] reg_0601;
  reg [8:0] reg_0602;
  reg [8:0] reg_0603;
  reg [8:0] reg_0604;
  reg [8:0] reg_0605;
  reg [8:0] reg_0606;
  reg [8:0] reg_0607;
  reg [8:0] reg_0608;
  reg [8:0] reg_0609;
  reg [8:0] reg_0610;
  reg [8:0] reg_0611;
  reg [8:0] reg_0612;
  reg [8:0] reg_0613;
  reg [8:0] reg_0614;
  reg [8:0] reg_0615;
  reg [8:0] reg_0616;
  reg [8:0] reg_0617;
  reg [8:0] reg_0618;
  reg [8:0] reg_0619;
  reg [8:0] reg_0620;
  reg [8:0] reg_0621;
  reg [8:0] reg_0622;
  reg [8:0] reg_0623;
  reg [8:0] reg_0624;
  reg [8:0] reg_0625;
  reg [8:0] reg_0626;
  reg [8:0] reg_0627;
  reg [8:0] reg_0628;
  reg [8:0] reg_0629;
  reg [8:0] reg_0630;
  reg [8:0] reg_0631;
  reg [8:0] reg_0632;
  reg [8:0] reg_0633;
  reg [8:0] reg_0634;
  reg [8:0] reg_0635;
  reg [8:0] reg_0636;
  reg [8:0] reg_0637;
  reg [8:0] reg_0638;
  reg [8:0] reg_0639;
  reg [8:0] reg_0640;
  reg [8:0] reg_0641;
  reg [8:0] reg_0642;
  reg [8:0] reg_0643;
  reg [8:0] reg_0644;
  reg [8:0] reg_0645;
  reg [8:0] reg_0646;
  reg [8:0] reg_0647;
  reg [8:0] reg_0648;
  reg [8:0] reg_0649;
  reg [8:0] reg_0650;
  reg [8:0] reg_0651;
  reg [8:0] reg_0652;
  reg [8:0] reg_0653;
  reg [8:0] reg_0654;
  reg [8:0] reg_0655;
  reg [8:0] reg_0656;
  reg [8:0] reg_0657;
  reg [8:0] reg_0658;
  reg [8:0] reg_0659;
  reg [8:0] reg_0660;
  reg [8:0] reg_0661;
  reg [8:0] reg_0662;
  reg [8:0] reg_0663;
  reg [8:0] reg_0664;
  reg [8:0] reg_0665;
  reg [8:0] reg_0666;
  reg [8:0] reg_0667;
  reg [8:0] reg_0668;
  reg [8:0] reg_0669;
  reg [8:0] reg_0670;
  reg [8:0] reg_0671;
  reg [8:0] reg_0672;
  reg [8:0] reg_0673;
  reg [8:0] reg_0674;
  reg [8:0] reg_0675;
  reg [8:0] reg_0676;
  reg [8:0] reg_0677;
  reg [8:0] reg_0678;
  reg [8:0] reg_0679;
  reg [8:0] reg_0680;
  reg [8:0] reg_0681;
  reg [8:0] reg_0682;
  reg [8:0] reg_0683;
  reg [8:0] reg_0684;
  reg [8:0] reg_0685;
  reg [8:0] reg_0686;
  reg [8:0] reg_0687;
  reg [8:0] reg_0688;
  reg [8:0] reg_0689;
  reg [8:0] reg_0690;
  reg [8:0] reg_0691;
  reg [8:0] reg_0692;
  reg [8:0] reg_0693;
  reg [8:0] reg_0694;
  reg [8:0] reg_0695;
  reg [8:0] reg_0696;
  reg [8:0] reg_0697;
  reg [8:0] reg_0698;
  reg [8:0] reg_0699;
  reg [8:0] reg_0700;
  reg [8:0] reg_0701;
  reg [8:0] reg_0702;
  reg [8:0] reg_0703;
  reg [8:0] reg_0704;
  reg [8:0] reg_0705;
  reg [8:0] reg_0706;
  reg [8:0] reg_0707;
  reg [8:0] reg_0708;
  reg [8:0] reg_0709;
  reg [8:0] reg_0710;
  reg [8:0] reg_0711;
  reg [8:0] reg_0712;
  reg [8:0] reg_0713;
  reg [8:0] reg_0714;
  reg [8:0] reg_0715;
  reg [8:0] reg_0716;
  reg [8:0] reg_0717;
  reg [8:0] reg_0718;
  reg [8:0] reg_0719;
  reg [8:0] reg_0720;
  reg [8:0] reg_0721;
  reg [8:0] reg_0722;
  reg [8:0] reg_0723;
  reg [8:0] reg_0724;
  reg [8:0] reg_0725;
  reg [8:0] reg_0726;
  reg [8:0] reg_0727;
  reg [8:0] reg_0728;
  reg [8:0] reg_0729;
  reg [8:0] reg_0730;
  reg [8:0] reg_0731;
  reg [8:0] reg_0732;
  reg [8:0] reg_0733;
  reg [8:0] reg_0734;
  reg [8:0] reg_0735;
  reg [8:0] reg_0736;
  reg [8:0] reg_0737;
  reg [8:0] reg_0738;
  reg [8:0] reg_0739;
  reg [8:0] reg_0740;
  reg [8:0] reg_0741;
  reg [8:0] reg_0742;
  reg [8:0] reg_0743;
  reg [8:0] reg_0744;
  reg [8:0] reg_0745;
  reg [8:0] reg_0746;
  reg [8:0] reg_0747;
  reg [8:0] reg_0748;
  reg [8:0] reg_0749;
  reg [8:0] reg_0750;
  reg [8:0] reg_0751;
  reg [8:0] reg_0752;
  reg [8:0] reg_0753;
  reg [8:0] reg_0754;
  reg [8:0] reg_0755;
  reg [8:0] reg_0756;
  reg [8:0] reg_0757;
  reg [8:0] reg_0758;
  reg [8:0] reg_0759;
  reg [8:0] reg_0760;
  reg [8:0] reg_0761;
  reg [8:0] reg_0762;
  reg [8:0] reg_0763;
  reg [8:0] reg_0764;
  reg [8:0] reg_0765;
  reg [8:0] reg_0766;
  reg [8:0] reg_0767;
  reg [8:0] reg_0768;
  reg [8:0] reg_0769;
  reg [8:0] reg_0770;
  reg [8:0] reg_0771;
  reg [8:0] reg_0772;
  reg [8:0] reg_0773;
  reg [8:0] reg_0774;
  reg [8:0] reg_0775;
  reg [8:0] reg_0776;
  reg [8:0] reg_0777;
  reg [8:0] reg_0778;
  reg [8:0] reg_0779;
  reg [8:0] reg_0780;
  reg [8:0] reg_0781;
  reg [8:0] reg_0782;
  reg [8:0] reg_0783;
  reg [8:0] reg_0784;
  reg [8:0] reg_0785;
  reg [8:0] reg_0786;
  reg [8:0] reg_0787;
  reg [8:0] reg_0788;
  reg [8:0] reg_0789;
  reg [8:0] reg_0790;
  reg [8:0] reg_0791;
  reg [8:0] reg_0792;
  reg [8:0] reg_0793;
  reg [8:0] reg_0794;
  reg [8:0] reg_0795;
  reg [8:0] reg_0796;
  reg [8:0] reg_0797;
  reg [8:0] reg_0798;
  reg [8:0] reg_0799;
  reg [8:0] reg_0800;
  reg [8:0] reg_0801;
  reg [8:0] reg_0802;
  reg [8:0] reg_0803;
  reg [8:0] reg_0804;
  reg [8:0] reg_0805;
  reg [8:0] reg_0806;
  reg [8:0] reg_0807;
  reg [8:0] reg_0808;
  reg [8:0] reg_0809;
  reg [8:0] reg_0810;
  reg [8:0] reg_0811;
  reg [8:0] reg_0812;
  reg [8:0] reg_0813;
  reg [8:0] reg_0814;
  reg [8:0] reg_0815;
  reg [8:0] reg_0816;
  reg [8:0] reg_0817;
  reg [8:0] reg_0818;
  reg [8:0] reg_0819;
  reg [8:0] reg_0820;
  reg [8:0] reg_0821;
  reg [8:0] reg_0822;
  reg [8:0] reg_0823;
  reg [8:0] reg_0824;
  reg [8:0] reg_0825;
  reg [8:0] reg_0826;
  reg [8:0] reg_0827;
  reg [8:0] reg_0828;
  reg [8:0] reg_0829;
  reg [8:0] reg_0830;
  reg [8:0] reg_0831;
  reg [8:0] reg_0832;
  reg [8:0] reg_0833;
  reg [8:0] reg_0834;
  reg [8:0] reg_0835;
  reg [8:0] reg_0836;
  reg [8:0] reg_0837;
  reg [8:0] reg_0838;
  reg [8:0] reg_0839;
  reg [8:0] reg_0840;
  reg [8:0] reg_0841;
  reg [8:0] reg_0842;
  reg [8:0] reg_0843;
  reg [8:0] reg_0844;
  reg [8:0] reg_0845;
  reg [8:0] reg_0846;
  reg [8:0] reg_0847;
  reg [8:0] reg_0848;
  reg [8:0] reg_0849;
  reg [8:0] reg_0850;
  reg [8:0] reg_0851;
  reg [8:0] reg_0852;
  reg [8:0] reg_0853;
  reg [8:0] reg_0854;
  reg [8:0] reg_0855;
  reg [8:0] reg_0856;
  reg [8:0] reg_0857;
  reg [8:0] reg_0858;
  reg [8:0] reg_0859;
  reg [8:0] reg_0860;
  reg [8:0] reg_0861;
  reg [8:0] reg_0862;
  reg [8:0] reg_0863;
  reg [8:0] reg_0864;
  reg [8:0] reg_0865;
  reg [8:0] reg_0866;
  reg [8:0] reg_0867;
  reg [8:0] reg_0868;
  reg [8:0] reg_0869;
  reg [8:0] reg_0870;
  reg [8:0] reg_0871;
  reg [8:0] reg_0872;
  reg [8:0] reg_0873;
  reg [8:0] reg_0874;
  reg [8:0] reg_0875;
  reg [8:0] reg_0876;
  reg [8:0] reg_0877;
  reg [8:0] reg_0878;
  reg [8:0] reg_0879;
  reg [8:0] reg_0880;
  reg [8:0] reg_0881;
  reg [8:0] reg_0882;
  reg [8:0] reg_0883;
  reg [8:0] reg_0884;
  reg [8:0] reg_0885;
  reg [8:0] reg_0886;
  reg [8:0] reg_0887;
  reg [8:0] reg_0888;
  reg [8:0] reg_0889;
  reg [8:0] reg_0890;
  reg [8:0] reg_0891;
  reg [8:0] reg_0892;
  reg [8:0] reg_0893;
  reg [8:0] reg_0894;
  reg [8:0] reg_0895;
  reg [8:0] reg_0896;
  reg [8:0] reg_0897;
  reg [8:0] reg_0898;
  reg [8:0] reg_0899;
  reg [8:0] reg_0900;
  reg [8:0] reg_0901;
  reg [8:0] reg_0902;
  reg [8:0] reg_0903;
  reg [8:0] reg_0904;
  reg [8:0] reg_0905;
  reg [8:0] reg_0906;
  reg [8:0] reg_0907;
  reg [8:0] reg_0908;
  reg [8:0] reg_0909;
  reg [8:0] reg_0910;
  reg [8:0] reg_0911;
  reg [8:0] reg_0912;
  reg [8:0] reg_0913;
  reg [8:0] reg_0914;
  reg [8:0] reg_0915;
  reg [8:0] reg_0916;
  reg [8:0] reg_0917;
  reg [8:0] reg_0918;
  reg [8:0] reg_0919;
  reg [8:0] reg_0920;
  reg [8:0] reg_0921;
  reg [8:0] reg_0922;
  reg [8:0] reg_0923;
  reg [8:0] reg_0924;
  reg [8:0] reg_0925;
  reg [8:0] reg_0926;
  reg [8:0] reg_0927;
  reg [8:0] reg_0928;
  reg [8:0] reg_0929;
  reg [8:0] reg_0930;
  reg [8:0] reg_0931;
  reg [8:0] reg_0932;
  reg [8:0] reg_0933;
  reg [8:0] reg_0934;
  reg [8:0] reg_0935;
  reg [8:0] reg_0936;
  reg [8:0] reg_0937;
  reg [8:0] reg_0938;
  reg [8:0] reg_0939;
  reg [8:0] reg_0940;
  reg [8:0] reg_0941;
  reg [8:0] reg_0942;
  reg [8:0] reg_0943;
  reg [8:0] reg_0944;
  reg [8:0] reg_0945;
  reg [8:0] reg_0946;
  reg [8:0] reg_0947;
  reg [8:0] reg_0948;
  reg [8:0] reg_0949;
  reg [8:0] reg_0950;
  reg [8:0] reg_0951;
  reg [8:0] reg_0952;
  reg [8:0] reg_0953;
  reg [8:0] reg_0954;
  reg [8:0] reg_0955;
  reg [8:0] reg_0956;
  reg [8:0] reg_0957;
  reg [8:0] reg_0958;
  reg [8:0] reg_0959;
  reg [8:0] reg_0960;
  reg [8:0] reg_0961;
  reg [8:0] reg_0962;
  reg [8:0] reg_0963;
  reg [8:0] reg_0964;
  reg [8:0] reg_0965;
  reg [8:0] reg_0966;
  reg [8:0] reg_0967;
  reg [8:0] reg_0968;
  reg [8:0] reg_0969;
  reg [8:0] reg_0970;
  reg [8:0] reg_0971;
  reg [8:0] reg_0972;
  reg [8:0] reg_0973;
  reg [8:0] reg_0974;
  reg [8:0] reg_0975;
  reg [8:0] reg_0976;
  reg [8:0] reg_0977;
  reg [8:0] reg_0978;
  reg [8:0] reg_0979;
  reg [8:0] reg_0980;
  reg [8:0] reg_0981;
  reg [8:0] reg_0982;
  reg [8:0] reg_0983;
  reg [8:0] reg_0984;
  reg [8:0] reg_0985;
  reg [8:0] reg_0986;
  reg [8:0] reg_0987;
  reg [8:0] reg_0988;
  reg [8:0] reg_0989;
  reg [8:0] reg_0990;
  reg [8:0] reg_0991;
  reg [8:0] reg_0992;
  reg [8:0] reg_0993;
  reg [8:0] reg_0994;
  reg [8:0] reg_0995;
  reg [8:0] reg_0996;
  reg [8:0] reg_0997;
  reg [8:0] reg_0998;
  reg [8:0] reg_0999;
  reg [8:0] reg_1000;
  reg [8:0] reg_1001;
  reg [8:0] reg_1002;
  reg [8:0] reg_1003;
  reg [8:0] reg_1004;
  reg [8:0] reg_1005;
  reg [8:0] reg_1006;
  reg [8:0] reg_1007;
  reg [8:0] reg_1008;
  reg [8:0] reg_1009;
  reg [8:0] reg_1010;
  reg [8:0] reg_1011;
  reg [8:0] reg_1012;
  reg [8:0] reg_1013;
  reg [8:0] reg_1014;
  reg [8:0] reg_1015;
  reg [8:0] reg_1016;
  reg [8:0] reg_1017;
  reg [8:0] reg_1018;
  reg [8:0] reg_1019;
  reg [8:0] reg_1020;
  reg [8:0] reg_1021;
  reg [8:0] reg_1022;
  reg [8:0] reg_1023;
  reg [8:0] reg_1024;
  reg [8:0] reg_1025;
  reg [8:0] reg_1026;
  reg [8:0] reg_1027;
  reg [8:0] reg_1028;
  reg [8:0] reg_1029;
  reg [8:0] reg_1030;
  reg [8:0] reg_1031;
  reg [8:0] reg_1032;
  reg [8:0] reg_1033;
  reg [8:0] reg_1034;
  reg [8:0] reg_1035;
  reg [8:0] reg_1036;
  reg [8:0] reg_1037;
  reg [8:0] reg_1038;
  reg [8:0] reg_1039;
  reg [8:0] reg_1040;
  reg [8:0] reg_1041;
  reg [8:0] reg_1042;
  reg [8:0] reg_1043;
  reg [8:0] reg_1044;
  reg [8:0] reg_1045;
  reg [8:0] reg_1046;
  reg [8:0] reg_1047;
  reg [8:0] reg_1048;
  reg [8:0] reg_1049;
  reg [8:0] reg_1050;
  reg [8:0] reg_1051;
  reg [8:0] reg_1052;
  reg [8:0] reg_1053;
  reg [8:0] reg_1054;
  reg [8:0] reg_1055;
  reg [8:0] reg_1056;
  reg [8:0] reg_1057;
  reg [8:0] reg_1058;
  reg [8:0] reg_1059;
  reg [8:0] reg_1060;
  reg [8:0] reg_1061;
  reg [8:0] reg_1062;
  reg [8:0] reg_1063;
  reg [8:0] reg_1064;
  reg [8:0] reg_1065;
  reg [8:0] reg_1066;
  reg [8:0] reg_1067;
  reg [8:0] reg_1068;
  reg [8:0] reg_1069;
  reg [8:0] reg_1070;
  reg [8:0] reg_1071;
  reg [8:0] reg_1072;
  reg [8:0] reg_1073;
  reg [8:0] reg_1074;
  reg [8:0] reg_1075;
  reg [8:0] reg_1076;
  reg [8:0] reg_1077;
  reg [8:0] reg_1078;
  reg [8:0] reg_1079;
  reg [8:0] reg_1080;
  reg [8:0] reg_1081;
  reg [8:0] reg_1082;
  reg [8:0] reg_1083;
  reg [8:0] reg_1084;
  reg [8:0] reg_1085;
  reg [8:0] reg_1086;
  reg [8:0] reg_1087;
  reg [8:0] reg_1088;
  reg [8:0] reg_1089;
  reg [8:0] reg_1090;
  reg [8:0] reg_1091;
  reg [8:0] reg_1092;
  reg [8:0] reg_1093;
  reg [8:0] reg_1094;
  reg [8:0] reg_1095;
  reg [8:0] reg_1096;
  reg [8:0] reg_1097;
  reg [8:0] reg_1098;
  reg [8:0] reg_1099;
  reg [8:0] reg_1100;
  reg [8:0] reg_1101;
  reg [8:0] reg_1102;
  reg [8:0] reg_1103;
  reg [8:0] reg_1104;
  reg [8:0] reg_1105;
  reg [8:0] reg_1106;
  reg [8:0] reg_1107;
  reg [8:0] reg_1108;
  reg [8:0] reg_1109;
  reg [8:0] reg_1110;
  reg [8:0] reg_1111;
  reg [8:0] reg_1112;
  reg [8:0] reg_1113;
  reg [8:0] reg_1114;
  reg [8:0] reg_1115;
  reg [8:0] reg_1116;
  reg [8:0] reg_1117;
  reg [8:0] reg_1118;
  reg [8:0] reg_1119;
  reg [8:0] reg_1120;
  reg [8:0] reg_1121;
  reg [8:0] reg_1122;
  reg [8:0] reg_1123;
  reg [8:0] reg_1124;
  reg [8:0] reg_1125;
  reg [8:0] reg_1126;
  reg [8:0] reg_1127;
  reg [8:0] reg_1128;
  reg [8:0] reg_1129;
  reg [8:0] reg_1130;
  reg [8:0] reg_1131;
  reg [8:0] reg_1132;
  reg [8:0] reg_1133;
  reg [8:0] reg_1134;
  reg [8:0] reg_1135;
  reg [8:0] reg_1136;
  reg [8:0] reg_1137;
  reg [8:0] reg_1138;
  reg [8:0] reg_1139;
  reg [8:0] reg_1140;
  reg [8:0] reg_1141;
  reg [8:0] reg_1142;
  reg [8:0] reg_1143;
  reg [8:0] reg_1144;
  reg [8:0] reg_1145;
  reg [8:0] reg_1146;
  reg [8:0] reg_1147;
  reg [8:0] reg_1148;
  reg [8:0] reg_1149;
  reg [8:0] reg_1150;
  reg [8:0] reg_1151;
  reg [8:0] reg_1152;
  reg [8:0] reg_1153;
  reg [8:0] reg_1154;
  reg [8:0] reg_1155;
  reg [8:0] reg_1156;
  reg [8:0] reg_1157;
  reg [8:0] reg_1158;
  reg [8:0] reg_1159;
  reg [8:0] reg_1160;
  reg [8:0] reg_1161;
  reg [8:0] reg_1162;
  reg [8:0] reg_1163;
  reg [8:0] reg_1164;
  reg [8:0] reg_1165;
  reg [8:0] reg_1166;
  reg [8:0] reg_1167;
  reg [8:0] reg_1168;
  reg [8:0] reg_1169;
  reg [8:0] reg_1170;
  reg [8:0] reg_1171;
  reg [8:0] reg_1172;
  reg [8:0] reg_1173;
  reg [8:0] reg_1174;
  reg [8:0] reg_1175;
  reg [8:0] reg_1176;
  reg [8:0] reg_1177;
  reg [8:0] reg_1178;
  reg [8:0] reg_1179;
  reg [8:0] reg_1180;
  reg [8:0] reg_1181;
  reg [8:0] reg_1182;
  reg [8:0] reg_1183;
  reg [8:0] reg_1184;
  reg [8:0] reg_1185;
  reg [8:0] reg_1186;
  reg [8:0] reg_1187;
  reg [8:0] reg_1188;
  reg [8:0] reg_1189;
  reg [8:0] reg_1190;
  reg [8:0] reg_1191;
  reg [8:0] reg_1192;
  reg [8:0] reg_1193;
  reg [8:0] reg_1194;
  reg [8:0] reg_1195;
  reg [8:0] reg_1196;
  reg [8:0] reg_1197;
  reg [8:0] reg_1198;
  reg [8:0] reg_1199;
  reg [8:0] reg_1200;
  reg [8:0] reg_1201;
  reg [8:0] reg_1202;
  reg [8:0] reg_1203;
  reg [8:0] reg_1204;
  reg [8:0] reg_1205;
  reg [8:0] reg_1206;
  reg [8:0] reg_1207;
  reg [8:0] reg_1208;
  reg [8:0] reg_1209;
  reg [8:0] reg_1210;
  reg [8:0] reg_1211;
  reg [8:0] reg_1212;
  reg [8:0] reg_1213;
  reg [8:0] reg_1214;
  reg [8:0] reg_1215;
  reg [8:0] reg_1216;
  reg [8:0] reg_1217;
  reg [8:0] reg_1218;
  reg [8:0] reg_1219;
  reg [8:0] reg_1220;
  reg [8:0] reg_1221;
  reg [8:0] reg_1222;
  reg [8:0] reg_1223;
  reg [8:0] reg_1224;
  reg [8:0] reg_1225;
  reg [8:0] reg_1226;
  reg [8:0] reg_1227;
  reg [8:0] reg_1228;
  reg [8:0] reg_1229;
  reg [8:0] reg_1230;
  reg [8:0] reg_1231;
  reg [8:0] reg_1232;
  reg [8:0] reg_1233;
  reg [8:0] reg_1234;
  reg [8:0] reg_1235;
  reg [8:0] reg_1236;
  reg [8:0] reg_1237;
  reg [8:0] reg_1238;
  reg [8:0] reg_1239;
  reg [8:0] reg_1240;
  reg [8:0] reg_1241;
  reg [8:0] reg_1242;
  reg [8:0] reg_1243;
  reg [8:0] reg_1244;
  reg [8:0] reg_1245;
  reg [8:0] reg_1246;
  reg [8:0] reg_1247;
  reg [8:0] reg_1248;
  reg [8:0] reg_1249;
  reg [8:0] reg_1250;
  reg [8:0] reg_1251;
  reg [8:0] reg_1252;
  reg [8:0] reg_1253;
  reg [8:0] reg_1254;
  reg [8:0] reg_1255;
  reg [8:0] reg_1256;
  reg [8:0] reg_1257;
  reg [8:0] reg_1258;
  reg [8:0] reg_1259;
  reg [8:0] reg_1260;
  reg [8:0] reg_1261;
  reg [8:0] reg_1262;
  reg [8:0] reg_1263;
  reg [8:0] reg_1264;
  reg [8:0] reg_1265;
  reg [8:0] reg_1266;
  reg [8:0] reg_1267;
  reg [8:0] reg_1268;
  reg [8:0] reg_1269;
  reg [8:0] reg_1270;
  reg [8:0] reg_1271;
  reg [8:0] reg_1272;
  reg [8:0] reg_1273;
  reg [8:0] reg_1274;
  reg [8:0] reg_1275;
  reg [8:0] reg_1276;
  reg [8:0] reg_1277;
  reg [8:0] reg_1278;
  reg [8:0] reg_1279;
  reg [8:0] reg_1280;
  reg [8:0] reg_1281;
  reg [8:0] reg_1282;
  reg [8:0] reg_1283;
  reg [8:0] reg_1284;
  reg [8:0] reg_1285;
  reg [8:0] reg_1286;
  reg [8:0] reg_1287;
  reg [8:0] reg_1288;
  reg [8:0] reg_1289;
  reg [8:0] reg_1290;
  reg [8:0] reg_1291;
  reg [8:0] reg_1292;
  reg [8:0] reg_1293;
  reg [8:0] reg_1294;
  reg [8:0] reg_1295;
  reg [8:0] reg_1296;
  reg [8:0] reg_1297;
  reg [8:0] reg_1298;
  reg [8:0] reg_1299;
  reg [8:0] reg_1300;
  reg [8:0] reg_1301;
  reg [8:0] reg_1302;
  reg [8:0] reg_1303;
  reg [8:0] reg_1304;
  reg [8:0] reg_1305;
  reg [8:0] reg_1306;
  reg [8:0] reg_1307;
  reg [8:0] reg_1308;
  reg [8:0] reg_1309;
  reg [8:0] reg_1310;
  reg [8:0] reg_1311;
  reg [8:0] reg_1312;
  reg [8:0] reg_1313;
  reg [8:0] reg_1314;
  reg [8:0] reg_1315;
  reg [8:0] reg_1316;
  reg [8:0] reg_1317;
  reg [8:0] reg_1318;
  reg [8:0] reg_1319;
  reg [8:0] reg_1320;
  reg [8:0] reg_1321;
  reg [8:0] reg_1322;
  reg [8:0] reg_1323;
  reg [8:0] reg_1324;
  reg [8:0] reg_1325;
  reg [8:0] reg_1326;
  reg [8:0] reg_1327;
  reg [8:0] reg_1328;
  reg [8:0] reg_1329;
  reg [8:0] reg_1330;
  reg [8:0] reg_1331;
  reg [8:0] reg_1332;
  reg [8:0] reg_1333;
  reg [8:0] reg_1334;
  reg [8:0] reg_1335;
  reg [8:0] reg_1336;
  reg [8:0] reg_1337;
  reg [8:0] reg_1338;
  reg [8:0] reg_1339;
  reg [8:0] reg_1340;
  reg [8:0] reg_1341;
  reg [8:0] reg_1342;
  reg [8:0] reg_1343;
  reg [8:0] reg_1344;
  reg [8:0] reg_1345;
  reg [8:0] reg_1346;
  reg [8:0] reg_1347;
  reg [8:0] reg_1348;
  reg [8:0] reg_1349;
  reg [8:0] reg_1350;
  reg [8:0] reg_1351;
  reg [8:0] reg_1352;
  reg [8:0] reg_1353;
  reg [8:0] reg_1354;
  reg [8:0] reg_1355;
  reg [8:0] reg_1356;
  reg [8:0] reg_1357;
  reg [8:0] reg_1358;
  reg [8:0] reg_1359;
  reg [8:0] reg_1360;
  reg [8:0] reg_1361;
  reg [8:0] reg_1362;
  reg [8:0] reg_1363;
  reg [8:0] reg_1364;
  reg [8:0] reg_1365;
  reg [8:0] reg_1366;
  reg [8:0] reg_1367;
  reg [8:0] reg_1368;
  reg [8:0] reg_1369;
  reg [8:0] reg_1370;
  reg [8:0] reg_1371;
  reg [8:0] reg_1372;
  reg [8:0] reg_1373;
  reg [8:0] reg_1374;
  reg [8:0] reg_1375;
  reg [8:0] reg_1376;
  reg [8:0] reg_1377;
  reg [8:0] reg_1378;
  reg [8:0] reg_1379;
  reg [8:0] reg_1380;
  reg [8:0] reg_1381;
  reg [8:0] reg_1382;
  reg [8:0] reg_1383;
  reg [8:0] reg_1384;
  reg [8:0] reg_1385;
  reg [8:0] reg_1386;
  reg [8:0] reg_1387;
  reg [8:0] reg_1388;
  reg [8:0] reg_1389;
  reg [8:0] reg_1390;
  reg [8:0] reg_1391;
  reg [8:0] reg_1392;
  reg [8:0] reg_1393;
  reg [8:0] reg_1394;
  reg [8:0] reg_1395;
  reg [8:0] reg_1396;
  reg [8:0] reg_1397;
  reg [8:0] reg_1398;
  reg [8:0] reg_1399;
  reg [8:0] reg_1400;
  reg [8:0] reg_1401;
  reg [8:0] reg_1402;
  reg [8:0] reg_1403;
  reg [8:0] reg_1404;
  reg [8:0] reg_1405;
  reg [8:0] reg_1406;
  reg [8:0] reg_1407;
  reg [8:0] reg_1408;
  reg [8:0] reg_1409;
  reg [8:0] reg_1410;
  reg [8:0] reg_1411;
  reg [8:0] reg_1412;
  reg [8:0] reg_1413;
  reg [8:0] reg_1414;
  reg [8:0] reg_1415;
  reg [8:0] reg_1416;
  reg [8:0] reg_1417;
  reg [8:0] reg_1418;
  reg [8:0] reg_1419;
  reg [8:0] reg_1420;
  reg [8:0] reg_1421;
  reg [8:0] reg_1422;
  reg [8:0] reg_1423;
  reg [8:0] reg_1424;
  reg [8:0] reg_1425;
  reg [8:0] reg_1426;
  reg [8:0] reg_1427;
  reg [8:0] reg_1428;
  reg [8:0] reg_1429;
  reg [8:0] reg_1430;
  reg [8:0] reg_1431;
  reg [8:0] reg_1432;
  reg [8:0] reg_1433;
  reg [8:0] reg_1434;
  reg [8:0] reg_1435;
  reg [8:0] reg_1436;
  reg [8:0] reg_1437;
  reg [8:0] reg_1438;
  reg [8:0] reg_1439;
  reg [8:0] reg_1440;
  reg [8:0] reg_1441;
  reg [8:0] reg_1442;
  reg [8:0] reg_1443;
  reg [8:0] reg_1444;
  reg [8:0] reg_1445;
  reg [8:0] reg_1446;
  reg [8:0] reg_1447;
  reg [8:0] reg_1448;
  reg [8:0] reg_1449;
  reg [8:0] reg_1450;
  reg [8:0] reg_1451;
  reg [8:0] reg_1452;
  reg [8:0] reg_1453;
  reg [8:0] reg_1454;
  reg [8:0] reg_1455;
  reg [8:0] reg_1456;
  reg [8:0] reg_1457;
  reg [8:0] reg_1458;
  reg [8:0] reg_1459;
  reg [8:0] reg_1460;
  reg [8:0] reg_1461;
  reg [8:0] reg_1462;
  reg [8:0] reg_1463;
  reg [8:0] reg_1464;
  reg [8:0] reg_1465;
  reg [8:0] reg_1466;
  reg [8:0] reg_1467;
  reg [8:0] reg_1468;
  reg [8:0] reg_1469;
  reg [8:0] reg_1470;
  reg [8:0] reg_1471;
  reg [8:0] reg_1472;
  reg [8:0] reg_1473;
  reg [8:0] reg_1474;
  reg [8:0] reg_1475;
  reg [8:0] reg_1476;
  reg [8:0] reg_1477;
  reg [8:0] reg_1478;
  reg [8:0] reg_1479;
  reg [8:0] reg_1480;
  reg [8:0] reg_1481;
  reg [8:0] reg_1482;
  reg [8:0] reg_1483;
  reg [8:0] reg_1484;
  reg [8:0] reg_1485;
  reg [8:0] reg_1486;
  reg [8:0] reg_1487;
  reg [8:0] reg_1488;
  reg [8:0] reg_1489;
  reg [8:0] reg_1490;
  reg [8:0] reg_1491;
  reg [8:0] reg_1492;
  reg [8:0] reg_1493;
  reg [8:0] reg_1494;
  reg [8:0] reg_1495;
  reg [8:0] reg_1496;
  reg [8:0] reg_1497;
  reg [8:0] reg_1498;
  reg [8:0] reg_1499;
  reg [8:0] reg_1500;
  reg [8:0] reg_1501;
  reg [8:0] reg_1502;
  reg [8:0] reg_1503;
  reg [8:0] reg_1504;
  reg [8:0] reg_1505;
  reg [8:0] reg_1506;
  reg [8:0] reg_1507;
  reg [8:0] reg_1508;
  reg [8:0] reg_1509;
  reg [8:0] reg_1510;
  reg [8:0] reg_1511;
  reg [8:0] reg_1512;
  reg [8:0] reg_1513;
  reg [8:0] reg_1514;
  reg [8:0] reg_1515;
  reg [8:0] reg_1516;
  reg [8:0] reg_1517;
  reg [8:0] reg_1518;

  // 制御マシンの状態
  reg [7:0] state;
  reg _busy;
  assign busy = _busy;
  // 制御マシンの動作
  always @ ( posedge clock or negedge reset ) begin
    if ( !reset ) begin
      _busy <= 0;
      state <= 0;
    end
    else if ( _busy ) begin
      if ( state < 174 ) begin
        state <= state + 1;
      end
      else begin
        _busy <= 0;
        state <= 0;
      end
    end
    else if ( start ) begin
      _busy <= 1;
    end
  end

  // 0番目の入力用メモリブロックの制御
  reg [4:0] _imem00_bank;
  always @ ( * ) begin
    case ( state )
    18: _imem00_bank = 3;
    17: _imem00_bank = 6;
    16: _imem00_bank = 7;
    15: _imem00_bank = 9;
    14: _imem00_bank = 11;
    13: _imem00_bank = 12;
    12: _imem00_bank = 13;
    11: _imem00_bank = 14;
    10: _imem00_bank = 15;
    9: _imem00_bank = 16;
    8: _imem00_bank = 17;
    7: _imem00_bank = 19;
    6: _imem00_bank = 21;
    5: _imem00_bank = 23;
    4: _imem00_bank = 25;
    3: _imem00_bank = 27;
    2: _imem00_bank = 28;
    1: _imem00_bank = 29;
    0: _imem00_bank = 30;
    31: _imem00_bank = 1;
    30: _imem00_bank = 2;
    29: _imem00_bank = 3;
    28: _imem00_bank = 6;
    27: _imem00_bank = 7;
    26: _imem00_bank = 13;
    25: _imem00_bank = 19;
    24: _imem00_bank = 23;
    23: _imem00_bank = 24;
    22: _imem00_bank = 25;
    21: _imem00_bank = 26;
    20: _imem00_bank = 29;
    39: _imem00_bank = 6;
    38: _imem00_bank = 7;
    37: _imem00_bank = 9;
    36: _imem00_bank = 11;
    35: _imem00_bank = 12;
    34: _imem00_bank = 14;
    33: _imem00_bank = 17;
    32: _imem00_bank = 21;
    19: _imem00_bank = 22;
    50: _imem00_bank = 0;
    49: _imem00_bank = 3;
    48: _imem00_bank = 5;
    47: _imem00_bank = 11;
    46: _imem00_bank = 12;
    45: _imem00_bank = 16;
    44: _imem00_bank = 17;
    43: _imem00_bank = 19;
    42: _imem00_bank = 22;
    41: _imem00_bank = 30;
    56: _imem00_bank = 2;
    55: _imem00_bank = 7;
    54: _imem00_bank = 14;
    53: _imem00_bank = 15;
    52: _imem00_bank = 16;
    51: _imem00_bank = 18;
    40: _imem00_bank = 20;
    58: _imem00_bank = 3;
    57: _imem00_bank = 4;
    74: _imem00_bank = 1;
    73: _imem00_bank = 2;
    72: _imem00_bank = 3;
    71: _imem00_bank = 6;
    70: _imem00_bank = 8;
    69: _imem00_bank = 10;
    68: _imem00_bank = 13;
    67: _imem00_bank = 16;
    66: _imem00_bank = 17;
    65: _imem00_bank = 18;
    64: _imem00_bank = 19;
    63: _imem00_bank = 21;
    62: _imem00_bank = 26;
    61: _imem00_bank = 27;
    60: _imem00_bank = 28;
    59: _imem00_bank = 31;
    75: _imem00_bank = 3;
    76: _imem00_bank = 8;
    77: _imem00_bank = 1;
    78: _imem00_bank = 0;
    79: _imem00_bank = 0;
    80: _imem00_bank = 5;
    81: _imem00_bank = 1;
    82: _imem00_bank = 1;
    83: _imem00_bank = 1;
    88: _imem00_bank = 1;
    87: _imem00_bank = 3;
    86: _imem00_bank = 7;
    85: _imem00_bank = 9;
    84: _imem00_bank = 10;
    89: _imem00_bank = 0;
    90: _imem00_bank = 0;
    91: _imem00_bank = 2;
    92: _imem00_bank = 0;
    93: _imem00_bank = 3;
    94: _imem00_bank = 0;
    95: _imem00_bank = 2;
    96: _imem00_bank = 1;
    97: _imem00_bank = 0;
    98: _imem00_bank = 5;
    99: _imem00_bank = 0;
    100: _imem00_bank = 3;
    101: _imem00_bank = 1;
    102: _imem00_bank = 2;
    103: _imem00_bank = 0;
    104: _imem00_bank = 0;
    105: _imem00_bank = 1;
    106: _imem00_bank = 0;
    107: _imem00_bank = 0;
    108: _imem00_bank = 0;
    109: _imem00_bank = 1;
    110: _imem00_bank = 2;
    111: _imem00_bank = 0;
    112: _imem00_bank = 0;
    113: _imem00_bank = 2;
    114: _imem00_bank = 0;
    115: _imem00_bank = 1;
    116: _imem00_bank = 0;
    117: _imem00_bank = 0;
    118: _imem00_bank = 0;
    119: _imem00_bank = 1;
    120: _imem00_bank = 0;
    121: _imem00_bank = 2;
    122: _imem00_bank = 3;
    123: _imem00_bank = 3;
    124: _imem00_bank = 8;
    125: _imem00_bank = 0;
    126: _imem00_bank = 0;
    127: _imem00_bank = 0;
    128: _imem00_bank = 4;
    129: _imem00_bank = 0;
    default: _imem00_bank = 0;
    endcase
  end // always @ ( * )
  assign imem00_bank = _imem00_bank;
  reg _imem00_rd;
  always @ ( * ) begin
    case ( state )
    18: _imem00_rd = 1;
    17: _imem00_rd = 1;
    16: _imem00_rd = 1;
    15: _imem00_rd = 1;
    14: _imem00_rd = 1;
    13: _imem00_rd = 1;
    12: _imem00_rd = 1;
    11: _imem00_rd = 1;
    10: _imem00_rd = 1;
    9: _imem00_rd = 1;
    8: _imem00_rd = 1;
    7: _imem00_rd = 1;
    6: _imem00_rd = 1;
    5: _imem00_rd = 1;
    4: _imem00_rd = 1;
    3: _imem00_rd = 1;
    2: _imem00_rd = 1;
    1: _imem00_rd = 1;
    0: _imem00_rd = 1;
    31: _imem00_rd = 1;
    30: _imem00_rd = 1;
    29: _imem00_rd = 1;
    28: _imem00_rd = 1;
    27: _imem00_rd = 1;
    26: _imem00_rd = 1;
    25: _imem00_rd = 1;
    24: _imem00_rd = 1;
    23: _imem00_rd = 1;
    22: _imem00_rd = 1;
    21: _imem00_rd = 1;
    20: _imem00_rd = 1;
    39: _imem00_rd = 1;
    38: _imem00_rd = 1;
    37: _imem00_rd = 1;
    36: _imem00_rd = 1;
    35: _imem00_rd = 1;
    34: _imem00_rd = 1;
    33: _imem00_rd = 1;
    32: _imem00_rd = 1;
    19: _imem00_rd = 1;
    50: _imem00_rd = 1;
    49: _imem00_rd = 1;
    48: _imem00_rd = 1;
    47: _imem00_rd = 1;
    46: _imem00_rd = 1;
    45: _imem00_rd = 1;
    44: _imem00_rd = 1;
    43: _imem00_rd = 1;
    42: _imem00_rd = 1;
    41: _imem00_rd = 1;
    56: _imem00_rd = 1;
    55: _imem00_rd = 1;
    54: _imem00_rd = 1;
    53: _imem00_rd = 1;
    52: _imem00_rd = 1;
    51: _imem00_rd = 1;
    40: _imem00_rd = 1;
    58: _imem00_rd = 1;
    57: _imem00_rd = 1;
    74: _imem00_rd = 1;
    73: _imem00_rd = 1;
    72: _imem00_rd = 1;
    71: _imem00_rd = 1;
    70: _imem00_rd = 1;
    69: _imem00_rd = 1;
    68: _imem00_rd = 1;
    67: _imem00_rd = 1;
    66: _imem00_rd = 1;
    65: _imem00_rd = 1;
    64: _imem00_rd = 1;
    63: _imem00_rd = 1;
    62: _imem00_rd = 1;
    61: _imem00_rd = 1;
    60: _imem00_rd = 1;
    59: _imem00_rd = 1;
    75: _imem00_rd = 1;
    76: _imem00_rd = 1;
    77: _imem00_rd = 1;
    78: _imem00_rd = 1;
    79: _imem00_rd = 1;
    80: _imem00_rd = 1;
    81: _imem00_rd = 1;
    82: _imem00_rd = 1;
    83: _imem00_rd = 1;
    88: _imem00_rd = 1;
    87: _imem00_rd = 1;
    86: _imem00_rd = 1;
    85: _imem00_rd = 1;
    84: _imem00_rd = 1;
    89: _imem00_rd = 1;
    90: _imem00_rd = 1;
    91: _imem00_rd = 1;
    92: _imem00_rd = 1;
    93: _imem00_rd = 1;
    94: _imem00_rd = 1;
    95: _imem00_rd = 1;
    96: _imem00_rd = 1;
    97: _imem00_rd = 1;
    98: _imem00_rd = 1;
    99: _imem00_rd = 1;
    100: _imem00_rd = 1;
    101: _imem00_rd = 1;
    102: _imem00_rd = 1;
    103: _imem00_rd = 1;
    104: _imem00_rd = 1;
    105: _imem00_rd = 1;
    106: _imem00_rd = 1;
    107: _imem00_rd = 1;
    108: _imem00_rd = 1;
    109: _imem00_rd = 1;
    110: _imem00_rd = 1;
    111: _imem00_rd = 1;
    112: _imem00_rd = 1;
    113: _imem00_rd = 1;
    114: _imem00_rd = 1;
    115: _imem00_rd = 1;
    116: _imem00_rd = 1;
    117: _imem00_rd = 1;
    118: _imem00_rd = 1;
    119: _imem00_rd = 1;
    120: _imem00_rd = 1;
    121: _imem00_rd = 1;
    122: _imem00_rd = 1;
    123: _imem00_rd = 1;
    124: _imem00_rd = 1;
    125: _imem00_rd = 1;
    126: _imem00_rd = 1;
    127: _imem00_rd = 1;
    128: _imem00_rd = 1;
    129: _imem00_rd = 1;
    default: _imem00_rd = 0;
    endcase
  end // always @ ( * )
  assign imem00_rd = _imem00_rd;

  // 1番目の入力用メモリブロックの制御
  reg [4:0] _imem01_bank;
  always @ ( * ) begin
    case ( state )
    18: _imem01_bank = 2;
    17: _imem01_bank = 3;
    16: _imem01_bank = 5;
    15: _imem01_bank = 9;
    13: _imem01_bank = 10;
    12: _imem01_bank = 11;
    11: _imem01_bank = 12;
    10: _imem01_bank = 13;
    9: _imem01_bank = 15;
    8: _imem01_bank = 16;
    7: _imem01_bank = 17;
    6: _imem01_bank = 18;
    5: _imem01_bank = 21;
    4: _imem01_bank = 23;
    3: _imem01_bank = 25;
    2: _imem01_bank = 26;
    1: _imem01_bank = 28;
    0: _imem01_bank = 29;
    31: _imem01_bank = 1;
    30: _imem01_bank = 3;
    29: _imem01_bank = 5;
    28: _imem01_bank = 8;
    27: _imem01_bank = 13;
    26: _imem01_bank = 14;
    25: _imem01_bank = 15;
    24: _imem01_bank = 16;
    23: _imem01_bank = 19;
    22: _imem01_bank = 20;
    21: _imem01_bank = 21;
    20: _imem01_bank = 22;
    19: _imem01_bank = 26;
    14: _imem01_bank = 27;
    33: _imem01_bank = 30;
    32: _imem01_bank = 31;
    39: _imem01_bank = 3;
    38: _imem01_bank = 5;
    37: _imem01_bank = 6;
    36: _imem01_bank = 12;
    35: _imem01_bank = 13;
    34: _imem01_bank = 14;
    50: _imem01_bank = 2;
    49: _imem01_bank = 3;
    48: _imem01_bank = 4;
    47: _imem01_bank = 5;
    46: _imem01_bank = 7;
    45: _imem01_bank = 13;
    44: _imem01_bank = 15;
    43: _imem01_bank = 17;
    42: _imem01_bank = 22;
    41: _imem01_bank = 23;
    40: _imem01_bank = 24;
    56: _imem01_bank = 1;
    55: _imem01_bank = 3;
    54: _imem01_bank = 6;
    53: _imem01_bank = 9;
    52: _imem01_bank = 12;
    51: _imem01_bank = 13;
    58: _imem01_bank = 2;
    57: _imem01_bank = 6;
    74: _imem01_bank = 4;
    73: _imem01_bank = 5;
    72: _imem01_bank = 7;
    71: _imem01_bank = 10;
    70: _imem01_bank = 12;
    69: _imem01_bank = 13;
    68: _imem01_bank = 17;
    59: _imem01_bank = 0;
    67: _imem01_bank = 6;
    66: _imem01_bank = 22;
    65: _imem01_bank = 23;
    64: _imem01_bank = 24;
    63: _imem01_bank = 1;
    62: _imem01_bank = 5;
    61: _imem01_bank = 7;
    60: _imem01_bank = 10;
    86: _imem01_bank = 23;
    85: _imem01_bank = 24;
    84: _imem01_bank = 25;
    83: _imem01_bank = 26;
    82: _imem01_bank = 27;
    75: _imem01_bank = 0;
    76: _imem01_bank = 4;
    77: _imem01_bank = 1;
    78: _imem01_bank = 1;
    81: _imem01_bank = 30;
    79: _imem01_bank = 1;
    80: _imem01_bank = 0;
    88: _imem01_bank = 1;
    87: _imem01_bank = 2;
    89: _imem01_bank = 0;
    90: _imem01_bank = 2;
    91: _imem01_bank = 0;
    92: _imem01_bank = 0;
    93: _imem01_bank = 5;
    94: _imem01_bank = 19;
    95: _imem01_bank = 27;
    96: _imem01_bank = 0;
    97: _imem01_bank = 0;
    98: _imem01_bank = 4;
    99: _imem01_bank = 1;
    100: _imem01_bank = 0;
    101: _imem01_bank = 4;
    102: _imem01_bank = 2;
    103: _imem01_bank = 29;
    104: _imem01_bank = 29;
    105: _imem01_bank = 0;
    106: _imem01_bank = 0;
    107: _imem01_bank = 3;
    108: _imem01_bank = 1;
    109: _imem01_bank = 0;
    110: _imem01_bank = 2;
    111: _imem01_bank = 2;
    112: _imem01_bank = 29;
    113: _imem01_bank = 1;
    114: _imem01_bank = 0;
    115: _imem01_bank = 0;
    116: _imem01_bank = 3;
    117: _imem01_bank = 2;
    118: _imem01_bank = 19;
    119: _imem01_bank = 1;
    120: _imem01_bank = 0;
    121: _imem01_bank = 1;
    122: _imem01_bank = 20;
    123: _imem01_bank = 0;
    124: _imem01_bank = 6;
    125: _imem01_bank = 1;
    126: _imem01_bank = 2;
    127: _imem01_bank = 1;
    128: _imem01_bank = 4;
    129: _imem01_bank = 2;
    default: _imem01_bank = 0;
    endcase
  end // always @ ( * )
  assign imem01_bank = _imem01_bank;
  reg _imem01_rd;
  always @ ( * ) begin
    case ( state )
    18: _imem01_rd = 1;
    17: _imem01_rd = 1;
    16: _imem01_rd = 1;
    15: _imem01_rd = 1;
    13: _imem01_rd = 1;
    12: _imem01_rd = 1;
    11: _imem01_rd = 1;
    10: _imem01_rd = 1;
    9: _imem01_rd = 1;
    8: _imem01_rd = 1;
    7: _imem01_rd = 1;
    6: _imem01_rd = 1;
    5: _imem01_rd = 1;
    4: _imem01_rd = 1;
    3: _imem01_rd = 1;
    2: _imem01_rd = 1;
    1: _imem01_rd = 1;
    0: _imem01_rd = 1;
    31: _imem01_rd = 1;
    30: _imem01_rd = 1;
    29: _imem01_rd = 1;
    28: _imem01_rd = 1;
    27: _imem01_rd = 1;
    26: _imem01_rd = 1;
    25: _imem01_rd = 1;
    24: _imem01_rd = 1;
    23: _imem01_rd = 1;
    22: _imem01_rd = 1;
    21: _imem01_rd = 1;
    20: _imem01_rd = 1;
    19: _imem01_rd = 1;
    14: _imem01_rd = 1;
    33: _imem01_rd = 1;
    32: _imem01_rd = 1;
    39: _imem01_rd = 1;
    38: _imem01_rd = 1;
    37: _imem01_rd = 1;
    36: _imem01_rd = 1;
    35: _imem01_rd = 1;
    34: _imem01_rd = 1;
    50: _imem01_rd = 1;
    49: _imem01_rd = 1;
    48: _imem01_rd = 1;
    47: _imem01_rd = 1;
    46: _imem01_rd = 1;
    45: _imem01_rd = 1;
    44: _imem01_rd = 1;
    43: _imem01_rd = 1;
    42: _imem01_rd = 1;
    41: _imem01_rd = 1;
    40: _imem01_rd = 1;
    56: _imem01_rd = 1;
    55: _imem01_rd = 1;
    54: _imem01_rd = 1;
    53: _imem01_rd = 1;
    52: _imem01_rd = 1;
    51: _imem01_rd = 1;
    58: _imem01_rd = 1;
    57: _imem01_rd = 1;
    74: _imem01_rd = 1;
    73: _imem01_rd = 1;
    72: _imem01_rd = 1;
    71: _imem01_rd = 1;
    70: _imem01_rd = 1;
    69: _imem01_rd = 1;
    68: _imem01_rd = 1;
    59: _imem01_rd = 1;
    67: _imem01_rd = 1;
    66: _imem01_rd = 1;
    65: _imem01_rd = 1;
    64: _imem01_rd = 1;
    63: _imem01_rd = 1;
    62: _imem01_rd = 1;
    61: _imem01_rd = 1;
    60: _imem01_rd = 1;
    86: _imem01_rd = 1;
    85: _imem01_rd = 1;
    84: _imem01_rd = 1;
    83: _imem01_rd = 1;
    82: _imem01_rd = 1;
    75: _imem01_rd = 1;
    76: _imem01_rd = 1;
    77: _imem01_rd = 1;
    78: _imem01_rd = 1;
    81: _imem01_rd = 1;
    79: _imem01_rd = 1;
    80: _imem01_rd = 1;
    88: _imem01_rd = 1;
    87: _imem01_rd = 1;
    89: _imem01_rd = 1;
    90: _imem01_rd = 1;
    91: _imem01_rd = 1;
    92: _imem01_rd = 1;
    93: _imem01_rd = 1;
    94: _imem01_rd = 1;
    95: _imem01_rd = 1;
    96: _imem01_rd = 1;
    97: _imem01_rd = 1;
    98: _imem01_rd = 1;
    99: _imem01_rd = 1;
    100: _imem01_rd = 1;
    101: _imem01_rd = 1;
    102: _imem01_rd = 1;
    103: _imem01_rd = 1;
    104: _imem01_rd = 1;
    105: _imem01_rd = 1;
    106: _imem01_rd = 1;
    107: _imem01_rd = 1;
    108: _imem01_rd = 1;
    109: _imem01_rd = 1;
    110: _imem01_rd = 1;
    111: _imem01_rd = 1;
    112: _imem01_rd = 1;
    113: _imem01_rd = 1;
    114: _imem01_rd = 1;
    115: _imem01_rd = 1;
    116: _imem01_rd = 1;
    117: _imem01_rd = 1;
    118: _imem01_rd = 1;
    119: _imem01_rd = 1;
    120: _imem01_rd = 1;
    121: _imem01_rd = 1;
    122: _imem01_rd = 1;
    123: _imem01_rd = 1;
    124: _imem01_rd = 1;
    125: _imem01_rd = 1;
    126: _imem01_rd = 1;
    127: _imem01_rd = 1;
    128: _imem01_rd = 1;
    129: _imem01_rd = 1;
    default: _imem01_rd = 0;
    endcase
  end // always @ ( * )
  assign imem01_rd = _imem01_rd;

  // 2番目の入力用メモリブロックの制御
  reg [4:0] _imem02_bank;
  always @ ( * ) begin
    case ( state )
    13: _imem02_bank = 1;
    12: _imem02_bank = 2;
    11: _imem02_bank = 4;
    10: _imem02_bank = 8;
    9: _imem02_bank = 10;
    8: _imem02_bank = 12;
    7: _imem02_bank = 13;
    6: _imem02_bank = 14;
    5: _imem02_bank = 17;
    4: _imem02_bank = 18;
    3: _imem02_bank = 19;
    2: _imem02_bank = 21;
    1: _imem02_bank = 24;
    17: _imem02_bank = 24;
    16: _imem02_bank = 25;
    33: _imem02_bank = 0;
    32: _imem02_bank = 2;
    31: _imem02_bank = 4;
    30: _imem02_bank = 6;
    29: _imem02_bank = 7;
    28: _imem02_bank = 8;
    27: _imem02_bank = 10;
    26: _imem02_bank = 11;
    25: _imem02_bank = 12;
    24: _imem02_bank = 13;
    23: _imem02_bank = 16;
    22: _imem02_bank = 19;
    21: _imem02_bank = 20;
    20: _imem02_bank = 23;
    19: _imem02_bank = 24;
    18: _imem02_bank = 27;
    15: _imem02_bank = 28;
    14: _imem02_bank = 30;
    36: _imem02_bank = 14;
    35: _imem02_bank = 16;
    34: _imem02_bank = 22;
    0: _imem02_bank = 26;
    50: _imem02_bank = 1;
    49: _imem02_bank = 2;
    48: _imem02_bank = 3;
    47: _imem02_bank = 4;
    46: _imem02_bank = 5;
    45: _imem02_bank = 12;
    44: _imem02_bank = 15;
    43: _imem02_bank = 16;
    42: _imem02_bank = 20;
    41: _imem02_bank = 21;
    40: _imem02_bank = 24;
    39: _imem02_bank = 25;
    38: _imem02_bank = 27;
    37: _imem02_bank = 29;
    52: _imem02_bank = 0;
    51: _imem02_bank = 9;
    59: _imem02_bank = 2;
    58: _imem02_bank = 4;
    57: _imem02_bank = 8;
    56: _imem02_bank = 9;
    55: _imem02_bank = 10;
    54: _imem02_bank = 11;
    53: _imem02_bank = 12;
    72: _imem02_bank = 0;
    71: _imem02_bank = 1;
    70: _imem02_bank = 6;
    69: _imem02_bank = 7;
    68: _imem02_bank = 16;
    67: _imem02_bank = 19;
    66: _imem02_bank = 21;
    65: _imem02_bank = 24;
    64: _imem02_bank = 26;
    63: _imem02_bank = 27;
    62: _imem02_bank = 1;
    61: _imem02_bank = 8;
    60: _imem02_bank = 10;
    84: _imem02_bank = 22;
    83: _imem02_bank = 23;
    82: _imem02_bank = 24;
    81: _imem02_bank = 29;
    80: _imem02_bank = 30;
    79: _imem02_bank = 27;
    78: _imem02_bank = 25;
    86: _imem02_bank = 0;
    85: _imem02_bank = 1;
    77: _imem02_bank = 3;
    76: _imem02_bank = 4;
    75: _imem02_bank = 10;
    74: _imem02_bank = 20;
    73: _imem02_bank = 31;
    87: _imem02_bank = 11;
    88: _imem02_bank = 9;
    89: _imem02_bank = 20;
    90: _imem02_bank = 2;
    91: _imem02_bank = 0;
    92: _imem02_bank = 0;
    93: _imem02_bank = 1;
    94: _imem02_bank = 1;
    95: _imem02_bank = 0;
    96: _imem02_bank = 1;
    97: _imem02_bank = 1;
    98: _imem02_bank = 1;
    99: _imem02_bank = 5;
    100: _imem02_bank = 8;
    101: _imem02_bank = 2;
    102: _imem02_bank = 0;
    103: _imem02_bank = 0;
    104: _imem02_bank = 0;
    105: _imem02_bank = 26;
    106: _imem02_bank = 1;
    107: _imem02_bank = 11;
    108: _imem02_bank = 1;
    109: _imem02_bank = 3;
    110: _imem02_bank = 0;
    111: _imem02_bank = 1;
    112: _imem02_bank = 0;
    113: _imem02_bank = 1;
    114: _imem02_bank = 1;
    115: _imem02_bank = 3;
    116: _imem02_bank = 3;
    117: _imem02_bank = 0;
    118: _imem02_bank = 0;
    119: _imem02_bank = 1;
    120: _imem02_bank = 0;
    121: _imem02_bank = 0;
    122: _imem02_bank = 1;
    123: _imem02_bank = 1;
    124: _imem02_bank = 2;
    125: _imem02_bank = 1;
    126: _imem02_bank = 0;
    127: _imem02_bank = 0;
    128: _imem02_bank = 1;
    129: _imem02_bank = 0;
    default: _imem02_bank = 0;
    endcase
  end // always @ ( * )
  assign imem02_bank = _imem02_bank;
  reg _imem02_rd;
  always @ ( * ) begin
    case ( state )
    13: _imem02_rd = 1;
    12: _imem02_rd = 1;
    11: _imem02_rd = 1;
    10: _imem02_rd = 1;
    9: _imem02_rd = 1;
    8: _imem02_rd = 1;
    7: _imem02_rd = 1;
    6: _imem02_rd = 1;
    5: _imem02_rd = 1;
    4: _imem02_rd = 1;
    3: _imem02_rd = 1;
    2: _imem02_rd = 1;
    1: _imem02_rd = 1;
    17: _imem02_rd = 1;
    16: _imem02_rd = 1;
    33: _imem02_rd = 1;
    32: _imem02_rd = 1;
    31: _imem02_rd = 1;
    30: _imem02_rd = 1;
    29: _imem02_rd = 1;
    28: _imem02_rd = 1;
    27: _imem02_rd = 1;
    26: _imem02_rd = 1;
    25: _imem02_rd = 1;
    24: _imem02_rd = 1;
    23: _imem02_rd = 1;
    22: _imem02_rd = 1;
    21: _imem02_rd = 1;
    20: _imem02_rd = 1;
    19: _imem02_rd = 1;
    18: _imem02_rd = 1;
    15: _imem02_rd = 1;
    14: _imem02_rd = 1;
    36: _imem02_rd = 1;
    35: _imem02_rd = 1;
    34: _imem02_rd = 1;
    0: _imem02_rd = 1;
    50: _imem02_rd = 1;
    49: _imem02_rd = 1;
    48: _imem02_rd = 1;
    47: _imem02_rd = 1;
    46: _imem02_rd = 1;
    45: _imem02_rd = 1;
    44: _imem02_rd = 1;
    43: _imem02_rd = 1;
    42: _imem02_rd = 1;
    41: _imem02_rd = 1;
    40: _imem02_rd = 1;
    39: _imem02_rd = 1;
    38: _imem02_rd = 1;
    37: _imem02_rd = 1;
    52: _imem02_rd = 1;
    51: _imem02_rd = 1;
    59: _imem02_rd = 1;
    58: _imem02_rd = 1;
    57: _imem02_rd = 1;
    56: _imem02_rd = 1;
    55: _imem02_rd = 1;
    54: _imem02_rd = 1;
    53: _imem02_rd = 1;
    72: _imem02_rd = 1;
    71: _imem02_rd = 1;
    70: _imem02_rd = 1;
    69: _imem02_rd = 1;
    68: _imem02_rd = 1;
    67: _imem02_rd = 1;
    66: _imem02_rd = 1;
    65: _imem02_rd = 1;
    64: _imem02_rd = 1;
    63: _imem02_rd = 1;
    62: _imem02_rd = 1;
    61: _imem02_rd = 1;
    60: _imem02_rd = 1;
    84: _imem02_rd = 1;
    83: _imem02_rd = 1;
    82: _imem02_rd = 1;
    81: _imem02_rd = 1;
    80: _imem02_rd = 1;
    79: _imem02_rd = 1;
    78: _imem02_rd = 1;
    86: _imem02_rd = 1;
    85: _imem02_rd = 1;
    77: _imem02_rd = 1;
    76: _imem02_rd = 1;
    75: _imem02_rd = 1;
    74: _imem02_rd = 1;
    73: _imem02_rd = 1;
    87: _imem02_rd = 1;
    88: _imem02_rd = 1;
    89: _imem02_rd = 1;
    90: _imem02_rd = 1;
    91: _imem02_rd = 1;
    92: _imem02_rd = 1;
    93: _imem02_rd = 1;
    94: _imem02_rd = 1;
    95: _imem02_rd = 1;
    96: _imem02_rd = 1;
    97: _imem02_rd = 1;
    98: _imem02_rd = 1;
    99: _imem02_rd = 1;
    100: _imem02_rd = 1;
    101: _imem02_rd = 1;
    102: _imem02_rd = 1;
    103: _imem02_rd = 1;
    104: _imem02_rd = 1;
    105: _imem02_rd = 1;
    106: _imem02_rd = 1;
    107: _imem02_rd = 1;
    108: _imem02_rd = 1;
    109: _imem02_rd = 1;
    110: _imem02_rd = 1;
    111: _imem02_rd = 1;
    112: _imem02_rd = 1;
    113: _imem02_rd = 1;
    114: _imem02_rd = 1;
    115: _imem02_rd = 1;
    116: _imem02_rd = 1;
    117: _imem02_rd = 1;
    118: _imem02_rd = 1;
    119: _imem02_rd = 1;
    120: _imem02_rd = 1;
    121: _imem02_rd = 1;
    122: _imem02_rd = 1;
    123: _imem02_rd = 1;
    124: _imem02_rd = 1;
    125: _imem02_rd = 1;
    126: _imem02_rd = 1;
    127: _imem02_rd = 1;
    128: _imem02_rd = 1;
    129: _imem02_rd = 1;
    default: _imem02_rd = 0;
    endcase
  end // always @ ( * )
  assign imem02_rd = _imem02_rd;

  // 3番目の入力用メモリブロックの制御
  reg [4:0] _imem03_bank;
  always @ ( * ) begin
    case ( state )
    17: _imem03_bank = 0;
    16: _imem03_bank = 2;
    15: _imem03_bank = 4;
    14: _imem03_bank = 6;
    13: _imem03_bank = 8;
    12: _imem03_bank = 10;
    11: _imem03_bank = 11;
    10: _imem03_bank = 12;
    9: _imem03_bank = 13;
    8: _imem03_bank = 14;
    7: _imem03_bank = 15;
    6: _imem03_bank = 17;
    5: _imem03_bank = 18;
    4: _imem03_bank = 23;
    3: _imem03_bank = 24;
    2: _imem03_bank = 25;
    1: _imem03_bank = 26;
    0: _imem03_bank = 31;
    33: _imem03_bank = 3;
    32: _imem03_bank = 5;
    31: _imem03_bank = 12;
    30: _imem03_bank = 20;
    29: _imem03_bank = 21;
    28: _imem03_bank = 24;
    27: _imem03_bank = 25;
    26: _imem03_bank = 26;
    25: _imem03_bank = 28;
    24: _imem03_bank = 30;
    23: _imem03_bank = 31;
    36: _imem03_bank = 1;
    35: _imem03_bank = 2;
    34: _imem03_bank = 6;
    22: _imem03_bank = 8;
    21: _imem03_bank = 11;
    20: _imem03_bank = 15;
    19: _imem03_bank = 18;
    18: _imem03_bank = 29;
    50: _imem03_bank = 0;
    49: _imem03_bank = 5;
    48: _imem03_bank = 7;
    47: _imem03_bank = 10;
    46: _imem03_bank = 12;
    45: _imem03_bank = 15;
    44: _imem03_bank = 16;
    43: _imem03_bank = 18;
    42: _imem03_bank = 19;
    41: _imem03_bank = 20;
    40: _imem03_bank = 24;
    39: _imem03_bank = 28;
    38: _imem03_bank = 29;
    52: _imem03_bank = 5;
    51: _imem03_bank = 10;
    37: _imem03_bank = 13;
    59: _imem03_bank = 17;
    58: _imem03_bank = 20;
    57: _imem03_bank = 29;
    65: _imem03_bank = 2;
    64: _imem03_bank = 5;
    63: _imem03_bank = 8;
    62: _imem03_bank = 10;
    61: _imem03_bank = 11;
    60: _imem03_bank = 12;
    56: _imem03_bank = 13;
    55: _imem03_bank = 14;
    54: _imem03_bank = 21;
    53: _imem03_bank = 22;
    66: _imem03_bank = 27;
    72: _imem03_bank = 1;
    71: _imem03_bank = 2;
    70: _imem03_bank = 3;
    69: _imem03_bank = 5;
    68: _imem03_bank = 7;
    67: _imem03_bank = 9;
    85: _imem03_bank = 25;
    84: _imem03_bank = 27;
    83: _imem03_bank = 28;
    82: _imem03_bank = 4;
    81: _imem03_bank = 5;
    80: _imem03_bank = 6;
    79: _imem03_bank = 8;
    78: _imem03_bank = 9;
    77: _imem03_bank = 10;
    76: _imem03_bank = 11;
    75: _imem03_bank = 14;
    74: _imem03_bank = 15;
    73: _imem03_bank = 16;
    86: _imem03_bank = 1;
    87: _imem03_bank = 11;
    88: _imem03_bank = 26;
    89: _imem03_bank = 0;
    90: _imem03_bank = 0;
    91: _imem03_bank = 14;
    92: _imem03_bank = 0;
    93: _imem03_bank = 0;
    94: _imem03_bank = 0;
    95: _imem03_bank = 0;
    96: _imem03_bank = 0;
    97: _imem03_bank = 0;
    98: _imem03_bank = 1;
    99: _imem03_bank = 0;
    100: _imem03_bank = 4;
    101: _imem03_bank = 2;
    102: _imem03_bank = 7;
    103: _imem03_bank = 2;
    104: _imem03_bank = 0;
    105: _imem03_bank = 0;
    106: _imem03_bank = 2;
    107: _imem03_bank = 2;
    108: _imem03_bank = 1;
    109: _imem03_bank = 19;
    110: _imem03_bank = 7;
    111: _imem03_bank = 1;
    112: _imem03_bank = 1;
    113: _imem03_bank = 0;
    114: _imem03_bank = 1;
    115: _imem03_bank = 0;
    116: _imem03_bank = 3;
    117: _imem03_bank = 2;
    118: _imem03_bank = 2;
    119: _imem03_bank = 20;
    120: _imem03_bank = 0;
    121: _imem03_bank = 26;
    122: _imem03_bank = 0;
    123: _imem03_bank = 2;
    124: _imem03_bank = 1;
    125: _imem03_bank = 3;
    126: _imem03_bank = 1;
    127: _imem03_bank = 2;
    128: _imem03_bank = 0;
    129: _imem03_bank = 1;
    default: _imem03_bank = 0;
    endcase
  end // always @ ( * )
  assign imem03_bank = _imem03_bank;
  reg _imem03_rd;
  always @ ( * ) begin
    case ( state )
    17: _imem03_rd = 1;
    16: _imem03_rd = 1;
    15: _imem03_rd = 1;
    14: _imem03_rd = 1;
    13: _imem03_rd = 1;
    12: _imem03_rd = 1;
    11: _imem03_rd = 1;
    10: _imem03_rd = 1;
    9: _imem03_rd = 1;
    8: _imem03_rd = 1;
    7: _imem03_rd = 1;
    6: _imem03_rd = 1;
    5: _imem03_rd = 1;
    4: _imem03_rd = 1;
    3: _imem03_rd = 1;
    2: _imem03_rd = 1;
    1: _imem03_rd = 1;
    0: _imem03_rd = 1;
    33: _imem03_rd = 1;
    32: _imem03_rd = 1;
    31: _imem03_rd = 1;
    30: _imem03_rd = 1;
    29: _imem03_rd = 1;
    28: _imem03_rd = 1;
    27: _imem03_rd = 1;
    26: _imem03_rd = 1;
    25: _imem03_rd = 1;
    24: _imem03_rd = 1;
    23: _imem03_rd = 1;
    36: _imem03_rd = 1;
    35: _imem03_rd = 1;
    34: _imem03_rd = 1;
    22: _imem03_rd = 1;
    21: _imem03_rd = 1;
    20: _imem03_rd = 1;
    19: _imem03_rd = 1;
    18: _imem03_rd = 1;
    50: _imem03_rd = 1;
    49: _imem03_rd = 1;
    48: _imem03_rd = 1;
    47: _imem03_rd = 1;
    46: _imem03_rd = 1;
    45: _imem03_rd = 1;
    44: _imem03_rd = 1;
    43: _imem03_rd = 1;
    42: _imem03_rd = 1;
    41: _imem03_rd = 1;
    40: _imem03_rd = 1;
    39: _imem03_rd = 1;
    38: _imem03_rd = 1;
    52: _imem03_rd = 1;
    51: _imem03_rd = 1;
    37: _imem03_rd = 1;
    59: _imem03_rd = 1;
    58: _imem03_rd = 1;
    57: _imem03_rd = 1;
    65: _imem03_rd = 1;
    64: _imem03_rd = 1;
    63: _imem03_rd = 1;
    62: _imem03_rd = 1;
    61: _imem03_rd = 1;
    60: _imem03_rd = 1;
    56: _imem03_rd = 1;
    55: _imem03_rd = 1;
    54: _imem03_rd = 1;
    53: _imem03_rd = 1;
    66: _imem03_rd = 1;
    72: _imem03_rd = 1;
    71: _imem03_rd = 1;
    70: _imem03_rd = 1;
    69: _imem03_rd = 1;
    68: _imem03_rd = 1;
    67: _imem03_rd = 1;
    85: _imem03_rd = 1;
    84: _imem03_rd = 1;
    83: _imem03_rd = 1;
    82: _imem03_rd = 1;
    81: _imem03_rd = 1;
    80: _imem03_rd = 1;
    79: _imem03_rd = 1;
    78: _imem03_rd = 1;
    77: _imem03_rd = 1;
    76: _imem03_rd = 1;
    75: _imem03_rd = 1;
    74: _imem03_rd = 1;
    73: _imem03_rd = 1;
    86: _imem03_rd = 1;
    87: _imem03_rd = 1;
    88: _imem03_rd = 1;
    89: _imem03_rd = 1;
    90: _imem03_rd = 1;
    91: _imem03_rd = 1;
    92: _imem03_rd = 1;
    93: _imem03_rd = 1;
    94: _imem03_rd = 1;
    95: _imem03_rd = 1;
    96: _imem03_rd = 1;
    97: _imem03_rd = 1;
    98: _imem03_rd = 1;
    99: _imem03_rd = 1;
    100: _imem03_rd = 1;
    101: _imem03_rd = 1;
    102: _imem03_rd = 1;
    103: _imem03_rd = 1;
    104: _imem03_rd = 1;
    105: _imem03_rd = 1;
    106: _imem03_rd = 1;
    107: _imem03_rd = 1;
    108: _imem03_rd = 1;
    109: _imem03_rd = 1;
    110: _imem03_rd = 1;
    111: _imem03_rd = 1;
    112: _imem03_rd = 1;
    113: _imem03_rd = 1;
    114: _imem03_rd = 1;
    115: _imem03_rd = 1;
    116: _imem03_rd = 1;
    117: _imem03_rd = 1;
    118: _imem03_rd = 1;
    119: _imem03_rd = 1;
    120: _imem03_rd = 1;
    121: _imem03_rd = 1;
    122: _imem03_rd = 1;
    123: _imem03_rd = 1;
    124: _imem03_rd = 1;
    125: _imem03_rd = 1;
    126: _imem03_rd = 1;
    127: _imem03_rd = 1;
    128: _imem03_rd = 1;
    129: _imem03_rd = 1;
    default: _imem03_rd = 0;
    endcase
  end // always @ ( * )
  assign imem03_rd = _imem03_rd;

  // 4番目の入力用メモリブロックの制御
  reg [4:0] _imem04_bank;
  always @ ( * ) begin
    case ( state )
    17: _imem04_bank = 0;
    16: _imem04_bank = 1;
    15: _imem04_bank = 4;
    14: _imem04_bank = 8;
    13: _imem04_bank = 13;
    9: _imem04_bank = 15;
    8: _imem04_bank = 17;
    7: _imem04_bank = 19;
    6: _imem04_bank = 20;
    5: _imem04_bank = 23;
    4: _imem04_bank = 24;
    3: _imem04_bank = 25;
    2: _imem04_bank = 28;
    1: _imem04_bank = 30;
    30: _imem04_bank = 0;
    29: _imem04_bank = 1;
    28: _imem04_bank = 3;
    27: _imem04_bank = 4;
    26: _imem04_bank = 6;
    25: _imem04_bank = 7;
    24: _imem04_bank = 12;
    23: _imem04_bank = 13;
    22: _imem04_bank = 17;
    21: _imem04_bank = 19;
    20: _imem04_bank = 20;
    19: _imem04_bank = 21;
    18: _imem04_bank = 23;
    12: _imem04_bank = 25;
    11: _imem04_bank = 26;
    10: _imem04_bank = 27;
    0: _imem04_bank = 29;
    36: _imem04_bank = 1;
    35: _imem04_bank = 8;
    34: _imem04_bank = 10;
    33: _imem04_bank = 11;
    32: _imem04_bank = 12;
    37: _imem04_bank = 15;
    31: _imem04_bank = 16;
    47: _imem04_bank = 4;
    46: _imem04_bank = 6;
    45: _imem04_bank = 8;
    44: _imem04_bank = 14;
    43: _imem04_bank = 16;
    42: _imem04_bank = 17;
    41: _imem04_bank = 18;
    40: _imem04_bank = 19;
    39: _imem04_bank = 21;
    38: _imem04_bank = 22;
    52: _imem04_bank = 0;
    51: _imem04_bank = 1;
    50: _imem04_bank = 4;
    49: _imem04_bank = 8;
    48: _imem04_bank = 10;
    59: _imem04_bank = 1;
    58: _imem04_bank = 2;
    57: _imem04_bank = 4;
    56: _imem04_bank = 6;
    55: _imem04_bank = 7;
    54: _imem04_bank = 8;
    53: _imem04_bank = 9;
    65: _imem04_bank = 0;
    64: _imem04_bank = 2;
    63: _imem04_bank = 3;
    62: _imem04_bank = 4;
    61: _imem04_bank = 6;
    60: _imem04_bank = 12;
    69: _imem04_bank = 15;
    68: _imem04_bank = 16;
    67: _imem04_bank = 18;
    66: _imem04_bank = 19;
    85: _imem04_bank = 0;
    84: _imem04_bank = 5;
    83: _imem04_bank = 8;
    82: _imem04_bank = 10;
    81: _imem04_bank = 11;
    80: _imem04_bank = 12;
    79: _imem04_bank = 15;
    78: _imem04_bank = 16;
    77: _imem04_bank = 18;
    76: _imem04_bank = 24;
    75: _imem04_bank = 25;
    74: _imem04_bank = 26;
    73: _imem04_bank = 27;
    72: _imem04_bank = 28;
    71: _imem04_bank = 30;
    70: _imem04_bank = 31;
    86: _imem04_bank = 0;
    87: _imem04_bank = 0;
    88: _imem04_bank = 2;
    89: _imem04_bank = 1;
    90: _imem04_bank = 6;
    91: _imem04_bank = 0;
    92: _imem04_bank = 2;
    93: _imem04_bank = 20;
    94: _imem04_bank = 1;
    95: _imem04_bank = 1;
    96: _imem04_bank = 0;
    97: _imem04_bank = 1;
    98: _imem04_bank = 0;
    99: _imem04_bank = 1;
    100: _imem04_bank = 0;
    101: _imem04_bank = 0;
    102: _imem04_bank = 0;
    103: _imem04_bank = 0;
    104: _imem04_bank = 0;
    105: _imem04_bank = 1;
    106: _imem04_bank = 23;
    107: _imem04_bank = 0;
    108: _imem04_bank = 0;
    109: _imem04_bank = 6;
    110: _imem04_bank = 3;
    111: _imem04_bank = 3;
    112: _imem04_bank = 1;
    113: _imem04_bank = 0;
    114: _imem04_bank = 0;
    115: _imem04_bank = 0;
    116: _imem04_bank = 2;
    117: _imem04_bank = 0;
    118: _imem04_bank = 2;
    119: _imem04_bank = 1;
    120: _imem04_bank = 1;
    121: _imem04_bank = 5;
    122: _imem04_bank = 1;
    123: _imem04_bank = 4;
    124: _imem04_bank = 0;
    125: _imem04_bank = 3;
    126: _imem04_bank = 0;
    127: _imem04_bank = 25;
    128: _imem04_bank = 2;
    129: _imem04_bank = 29;
    default: _imem04_bank = 0;
    endcase
  end // always @ ( * )
  assign imem04_bank = _imem04_bank;
  reg _imem04_rd;
  always @ ( * ) begin
    case ( state )
    17: _imem04_rd = 1;
    16: _imem04_rd = 1;
    15: _imem04_rd = 1;
    14: _imem04_rd = 1;
    13: _imem04_rd = 1;
    9: _imem04_rd = 1;
    8: _imem04_rd = 1;
    7: _imem04_rd = 1;
    6: _imem04_rd = 1;
    5: _imem04_rd = 1;
    4: _imem04_rd = 1;
    3: _imem04_rd = 1;
    2: _imem04_rd = 1;
    1: _imem04_rd = 1;
    30: _imem04_rd = 1;
    29: _imem04_rd = 1;
    28: _imem04_rd = 1;
    27: _imem04_rd = 1;
    26: _imem04_rd = 1;
    25: _imem04_rd = 1;
    24: _imem04_rd = 1;
    23: _imem04_rd = 1;
    22: _imem04_rd = 1;
    21: _imem04_rd = 1;
    20: _imem04_rd = 1;
    19: _imem04_rd = 1;
    18: _imem04_rd = 1;
    12: _imem04_rd = 1;
    11: _imem04_rd = 1;
    10: _imem04_rd = 1;
    0: _imem04_rd = 1;
    36: _imem04_rd = 1;
    35: _imem04_rd = 1;
    34: _imem04_rd = 1;
    33: _imem04_rd = 1;
    32: _imem04_rd = 1;
    37: _imem04_rd = 1;
    31: _imem04_rd = 1;
    47: _imem04_rd = 1;
    46: _imem04_rd = 1;
    45: _imem04_rd = 1;
    44: _imem04_rd = 1;
    43: _imem04_rd = 1;
    42: _imem04_rd = 1;
    41: _imem04_rd = 1;
    40: _imem04_rd = 1;
    39: _imem04_rd = 1;
    38: _imem04_rd = 1;
    52: _imem04_rd = 1;
    51: _imem04_rd = 1;
    50: _imem04_rd = 1;
    49: _imem04_rd = 1;
    48: _imem04_rd = 1;
    59: _imem04_rd = 1;
    58: _imem04_rd = 1;
    57: _imem04_rd = 1;
    56: _imem04_rd = 1;
    55: _imem04_rd = 1;
    54: _imem04_rd = 1;
    53: _imem04_rd = 1;
    65: _imem04_rd = 1;
    64: _imem04_rd = 1;
    63: _imem04_rd = 1;
    62: _imem04_rd = 1;
    61: _imem04_rd = 1;
    60: _imem04_rd = 1;
    69: _imem04_rd = 1;
    68: _imem04_rd = 1;
    67: _imem04_rd = 1;
    66: _imem04_rd = 1;
    85: _imem04_rd = 1;
    84: _imem04_rd = 1;
    83: _imem04_rd = 1;
    82: _imem04_rd = 1;
    81: _imem04_rd = 1;
    80: _imem04_rd = 1;
    79: _imem04_rd = 1;
    78: _imem04_rd = 1;
    77: _imem04_rd = 1;
    76: _imem04_rd = 1;
    75: _imem04_rd = 1;
    74: _imem04_rd = 1;
    73: _imem04_rd = 1;
    72: _imem04_rd = 1;
    71: _imem04_rd = 1;
    70: _imem04_rd = 1;
    86: _imem04_rd = 1;
    87: _imem04_rd = 1;
    88: _imem04_rd = 1;
    89: _imem04_rd = 1;
    90: _imem04_rd = 1;
    91: _imem04_rd = 1;
    92: _imem04_rd = 1;
    93: _imem04_rd = 1;
    94: _imem04_rd = 1;
    95: _imem04_rd = 1;
    96: _imem04_rd = 1;
    97: _imem04_rd = 1;
    98: _imem04_rd = 1;
    99: _imem04_rd = 1;
    100: _imem04_rd = 1;
    101: _imem04_rd = 1;
    102: _imem04_rd = 1;
    103: _imem04_rd = 1;
    104: _imem04_rd = 1;
    105: _imem04_rd = 1;
    106: _imem04_rd = 1;
    107: _imem04_rd = 1;
    108: _imem04_rd = 1;
    109: _imem04_rd = 1;
    110: _imem04_rd = 1;
    111: _imem04_rd = 1;
    112: _imem04_rd = 1;
    113: _imem04_rd = 1;
    114: _imem04_rd = 1;
    115: _imem04_rd = 1;
    116: _imem04_rd = 1;
    117: _imem04_rd = 1;
    118: _imem04_rd = 1;
    119: _imem04_rd = 1;
    120: _imem04_rd = 1;
    121: _imem04_rd = 1;
    122: _imem04_rd = 1;
    123: _imem04_rd = 1;
    124: _imem04_rd = 1;
    125: _imem04_rd = 1;
    126: _imem04_rd = 1;
    127: _imem04_rd = 1;
    128: _imem04_rd = 1;
    129: _imem04_rd = 1;
    default: _imem04_rd = 0;
    endcase
  end // always @ ( * )
  assign imem04_rd = _imem04_rd;

  // 5番目の入力用メモリブロックの制御
  reg [4:0] _imem05_bank;
  always @ ( * ) begin
    case ( state )
    9: _imem05_bank = 1;
    8: _imem05_bank = 9;
    7: _imem05_bank = 10;
    6: _imem05_bank = 15;
    5: _imem05_bank = 17;
    4: _imem05_bank = 21;
    3: _imem05_bank = 24;
    2: _imem05_bank = 25;
    1: _imem05_bank = 30;
    0: _imem05_bank = 31;
    30: _imem05_bank = 1;
    24: _imem05_bank = 1;
    23: _imem05_bank = 2;
    22: _imem05_bank = 4;
    21: _imem05_bank = 5;
    20: _imem05_bank = 7;
    19: _imem05_bank = 10;
    18: _imem05_bank = 15;
    17: _imem05_bank = 16;
    16: _imem05_bank = 22;
    15: _imem05_bank = 24;
    14: _imem05_bank = 26;
    13: _imem05_bank = 28;
    37: _imem05_bank = 0;
    36: _imem05_bank = 3;
    35: _imem05_bank = 4;
    34: _imem05_bank = 7;
    33: _imem05_bank = 10;
    32: _imem05_bank = 11;
    31: _imem05_bank = 12;
    29: _imem05_bank = 13;
    28: _imem05_bank = 17;
    27: _imem05_bank = 18;
    26: _imem05_bank = 20;
    25: _imem05_bank = 23;
    12: _imem05_bank = 25;
    47: _imem05_bank = 9;
    46: _imem05_bank = 10;
    45: _imem05_bank = 12;
    44: _imem05_bank = 15;
    43: _imem05_bank = 18;
    42: _imem05_bank = 19;
    41: _imem05_bank = 21;
    40: _imem05_bank = 23;
    39: _imem05_bank = 28;
    50: _imem05_bank = 1;
    49: _imem05_bank = 2;
    48: _imem05_bank = 5;
    38: _imem05_bank = 6;
    11: _imem05_bank = 14;
    10: _imem05_bank = 29;
    59: _imem05_bank = 2;
    58: _imem05_bank = 3;
    57: _imem05_bank = 5;
    56: _imem05_bank = 7;
    55: _imem05_bank = 9;
    54: _imem05_bank = 12;
    53: _imem05_bank = 14;
    52: _imem05_bank = 15;
    65: _imem05_bank = 16;
    64: _imem05_bank = 21;
    63: _imem05_bank = 23;
    62: _imem05_bank = 24;
    61: _imem05_bank = 26;
    60: _imem05_bank = 29;
    69: _imem05_bank = 0;
    68: _imem05_bank = 1;
    67: _imem05_bank = 4;
    66: _imem05_bank = 6;
    51: _imem05_bank = 8;
    70: _imem05_bank = 27;
    85: _imem05_bank = 5;
    84: _imem05_bank = 6;
    83: _imem05_bank = 7;
    82: _imem05_bank = 10;
    81: _imem05_bank = 11;
    80: _imem05_bank = 12;
    79: _imem05_bank = 13;
    78: _imem05_bank = 14;
    76: _imem05_bank = 14;
    75: _imem05_bank = 17;
    74: _imem05_bank = 18;
    73: _imem05_bank = 19;
    72: _imem05_bank = 20;
    71: _imem05_bank = 22;
    77: _imem05_bank = 0;
    86: _imem05_bank = 0;
    87: _imem05_bank = 0;
    88: _imem05_bank = 0;
    89: _imem05_bank = 27;
    90: _imem05_bank = 8;
    91: _imem05_bank = 1;
    92: _imem05_bank = 0;
    93: _imem05_bank = 3;
    94: _imem05_bank = 2;
    95: _imem05_bank = 0;
    96: _imem05_bank = 0;
    97: _imem05_bank = 0;
    98: _imem05_bank = 1;
    99: _imem05_bank = 0;
    100: _imem05_bank = 22;
    101: _imem05_bank = 18;
    102: _imem05_bank = 0;
    103: _imem05_bank = 1;
    104: _imem05_bank = 3;
    105: _imem05_bank = 1;
    106: _imem05_bank = 3;
    107: _imem05_bank = 3;
    108: _imem05_bank = 1;
    109: _imem05_bank = 0;
    110: _imem05_bank = 0;
    111: _imem05_bank = 0;
    112: _imem05_bank = 4;
    113: _imem05_bank = 30;
    114: _imem05_bank = 1;
    115: _imem05_bank = 3;
    116: _imem05_bank = 31;
    117: _imem05_bank = 6;
    118: _imem05_bank = 1;
    119: _imem05_bank = 2;
    120: _imem05_bank = 10;
    121: _imem05_bank = 1;
    122: _imem05_bank = 0;
    123: _imem05_bank = 2;
    124: _imem05_bank = 0;
    125: _imem05_bank = 23;
    126: _imem05_bank = 0;
    127: _imem05_bank = 0;
    128: _imem05_bank = 1;
    129: _imem05_bank = 0;
    default: _imem05_bank = 0;
    endcase
  end // always @ ( * )
  assign imem05_bank = _imem05_bank;
  reg _imem05_rd;
  always @ ( * ) begin
    case ( state )
    9: _imem05_rd = 1;
    8: _imem05_rd = 1;
    7: _imem05_rd = 1;
    6: _imem05_rd = 1;
    5: _imem05_rd = 1;
    4: _imem05_rd = 1;
    3: _imem05_rd = 1;
    2: _imem05_rd = 1;
    1: _imem05_rd = 1;
    0: _imem05_rd = 1;
    30: _imem05_rd = 1;
    24: _imem05_rd = 1;
    23: _imem05_rd = 1;
    22: _imem05_rd = 1;
    21: _imem05_rd = 1;
    20: _imem05_rd = 1;
    19: _imem05_rd = 1;
    18: _imem05_rd = 1;
    17: _imem05_rd = 1;
    16: _imem05_rd = 1;
    15: _imem05_rd = 1;
    14: _imem05_rd = 1;
    13: _imem05_rd = 1;
    37: _imem05_rd = 1;
    36: _imem05_rd = 1;
    35: _imem05_rd = 1;
    34: _imem05_rd = 1;
    33: _imem05_rd = 1;
    32: _imem05_rd = 1;
    31: _imem05_rd = 1;
    29: _imem05_rd = 1;
    28: _imem05_rd = 1;
    27: _imem05_rd = 1;
    26: _imem05_rd = 1;
    25: _imem05_rd = 1;
    12: _imem05_rd = 1;
    47: _imem05_rd = 1;
    46: _imem05_rd = 1;
    45: _imem05_rd = 1;
    44: _imem05_rd = 1;
    43: _imem05_rd = 1;
    42: _imem05_rd = 1;
    41: _imem05_rd = 1;
    40: _imem05_rd = 1;
    39: _imem05_rd = 1;
    50: _imem05_rd = 1;
    49: _imem05_rd = 1;
    48: _imem05_rd = 1;
    38: _imem05_rd = 1;
    11: _imem05_rd = 1;
    10: _imem05_rd = 1;
    59: _imem05_rd = 1;
    58: _imem05_rd = 1;
    57: _imem05_rd = 1;
    56: _imem05_rd = 1;
    55: _imem05_rd = 1;
    54: _imem05_rd = 1;
    53: _imem05_rd = 1;
    52: _imem05_rd = 1;
    65: _imem05_rd = 1;
    64: _imem05_rd = 1;
    63: _imem05_rd = 1;
    62: _imem05_rd = 1;
    61: _imem05_rd = 1;
    60: _imem05_rd = 1;
    69: _imem05_rd = 1;
    68: _imem05_rd = 1;
    67: _imem05_rd = 1;
    66: _imem05_rd = 1;
    51: _imem05_rd = 1;
    70: _imem05_rd = 1;
    85: _imem05_rd = 1;
    84: _imem05_rd = 1;
    83: _imem05_rd = 1;
    82: _imem05_rd = 1;
    81: _imem05_rd = 1;
    80: _imem05_rd = 1;
    79: _imem05_rd = 1;
    78: _imem05_rd = 1;
    76: _imem05_rd = 1;
    75: _imem05_rd = 1;
    74: _imem05_rd = 1;
    73: _imem05_rd = 1;
    72: _imem05_rd = 1;
    71: _imem05_rd = 1;
    77: _imem05_rd = 1;
    86: _imem05_rd = 1;
    87: _imem05_rd = 1;
    88: _imem05_rd = 1;
    89: _imem05_rd = 1;
    90: _imem05_rd = 1;
    91: _imem05_rd = 1;
    92: _imem05_rd = 1;
    93: _imem05_rd = 1;
    94: _imem05_rd = 1;
    95: _imem05_rd = 1;
    96: _imem05_rd = 1;
    97: _imem05_rd = 1;
    98: _imem05_rd = 1;
    99: _imem05_rd = 1;
    100: _imem05_rd = 1;
    101: _imem05_rd = 1;
    102: _imem05_rd = 1;
    103: _imem05_rd = 1;
    104: _imem05_rd = 1;
    105: _imem05_rd = 1;
    106: _imem05_rd = 1;
    107: _imem05_rd = 1;
    108: _imem05_rd = 1;
    109: _imem05_rd = 1;
    110: _imem05_rd = 1;
    111: _imem05_rd = 1;
    112: _imem05_rd = 1;
    113: _imem05_rd = 1;
    114: _imem05_rd = 1;
    115: _imem05_rd = 1;
    116: _imem05_rd = 1;
    117: _imem05_rd = 1;
    118: _imem05_rd = 1;
    119: _imem05_rd = 1;
    120: _imem05_rd = 1;
    121: _imem05_rd = 1;
    122: _imem05_rd = 1;
    123: _imem05_rd = 1;
    124: _imem05_rd = 1;
    125: _imem05_rd = 1;
    126: _imem05_rd = 1;
    127: _imem05_rd = 1;
    128: _imem05_rd = 1;
    129: _imem05_rd = 1;
    default: _imem05_rd = 0;
    endcase
  end // always @ ( * )
  assign imem05_rd = _imem05_rd;

  // 6番目の入力用メモリブロックの制御
  reg [4:0] _imem06_bank;
  always @ ( * ) begin
    case ( state )
    9: _imem06_bank = 2;
    8: _imem06_bank = 3;
    7: _imem06_bank = 6;
    6: _imem06_bank = 10;
    5: _imem06_bank = 11;
    4: _imem06_bank = 14;
    3: _imem06_bank = 15;
    2: _imem06_bank = 16;
    1: _imem06_bank = 17;
    13: _imem06_bank = 23;
    12: _imem06_bank = 24;
    11: _imem06_bank = 28;
    10: _imem06_bank = 29;
    0: _imem06_bank = 30;
    24: _imem06_bank = 0;
    23: _imem06_bank = 9;
    22: _imem06_bank = 11;
    21: _imem06_bank = 12;
    20: _imem06_bank = 16;
    19: _imem06_bank = 18;
    18: _imem06_bank = 21;
    17: _imem06_bank = 22;
    16: _imem06_bank = 23;
    15: _imem06_bank = 25;
    14: _imem06_bank = 27;
    37: _imem06_bank = 0;
    36: _imem06_bank = 1;
    35: _imem06_bank = 3;
    43: _imem06_bank = 3;
    42: _imem06_bank = 5;
    41: _imem06_bank = 6;
    40: _imem06_bank = 8;
    39: _imem06_bank = 10;
    38: _imem06_bank = 12;
    34: _imem06_bank = 15;
    33: _imem06_bank = 16;
    32: _imem06_bank = 17;
    31: _imem06_bank = 19;
    30: _imem06_bank = 20;
    29: _imem06_bank = 21;
    28: _imem06_bank = 22;
    27: _imem06_bank = 23;
    26: _imem06_bank = 24;
    25: _imem06_bank = 26;
    47: _imem06_bank = 0;
    46: _imem06_bank = 4;
    45: _imem06_bank = 5;
    44: _imem06_bank = 7;
    50: _imem06_bank = 2;
    49: _imem06_bank = 4;
    48: _imem06_bank = 5;
    65: _imem06_bank = 0;
    64: _imem06_bank = 1;
    63: _imem06_bank = 4;
    62: _imem06_bank = 8;
    61: _imem06_bank = 9;
    60: _imem06_bank = 11;
    59: _imem06_bank = 12;
    58: _imem06_bank = 16;
    57: _imem06_bank = 17;
    56: _imem06_bank = 18;
    55: _imem06_bank = 20;
    54: _imem06_bank = 22;
    53: _imem06_bank = 26;
    52: _imem06_bank = 27;
    51: _imem06_bank = 31;
    70: _imem06_bank = 2;
    69: _imem06_bank = 3;
    68: _imem06_bank = 4;
    67: _imem06_bank = 5;
    66: _imem06_bank = 7;
    76: _imem06_bank = 2;
    75: _imem06_bank = 4;
    74: _imem06_bank = 6;
    73: _imem06_bank = 8;
    72: _imem06_bank = 12;
    71: _imem06_bank = 13;
    77: _imem06_bank = 0;
    78: _imem06_bank = 13;
    87: _imem06_bank = 2;
    86: _imem06_bank = 3;
    85: _imem06_bank = 5;
    79: _imem06_bank = 1;
    80: _imem06_bank = 1;
    81: _imem06_bank = 3;
    82: _imem06_bank = 0;
    84: _imem06_bank = 0;
    83: _imem06_bank = 9;
    88: _imem06_bank = 3;
    89: _imem06_bank = 0;
    90: _imem06_bank = 0;
    91: _imem06_bank = 8;
    92: _imem06_bank = 0;
    93: _imem06_bank = 8;
    94: _imem06_bank = 0;
    95: _imem06_bank = 1;
    96: _imem06_bank = 27;
    97: _imem06_bank = 3;
    98: _imem06_bank = 0;
    99: _imem06_bank = 13;
    100: _imem06_bank = 0;
    101: _imem06_bank = 0;
    102: _imem06_bank = 0;
    103: _imem06_bank = 0;
    104: _imem06_bank = 0;
    105: _imem06_bank = 0;
    106: _imem06_bank = 2;
    107: _imem06_bank = 0;
    108: _imem06_bank = 2;
    109: _imem06_bank = 0;
    110: _imem06_bank = 3;
    111: _imem06_bank = 0;
    112: _imem06_bank = 4;
    113: _imem06_bank = 3;
    114: _imem06_bank = 1;
    115: _imem06_bank = 0;
    116: _imem06_bank = 0;
    117: _imem06_bank = 1;
    118: _imem06_bank = 3;
    119: _imem06_bank = 0;
    120: _imem06_bank = 1;
    121: _imem06_bank = 2;
    122: _imem06_bank = 0;
    123: _imem06_bank = 0;
    124: _imem06_bank = 4;
    125: _imem06_bank = 0;
    126: _imem06_bank = 1;
    127: _imem06_bank = 2;
    128: _imem06_bank = 5;
    129: _imem06_bank = 0;
    default: _imem06_bank = 0;
    endcase
  end // always @ ( * )
  assign imem06_bank = _imem06_bank;
  reg _imem06_rd;
  always @ ( * ) begin
    case ( state )
    9: _imem06_rd = 1;
    8: _imem06_rd = 1;
    7: _imem06_rd = 1;
    6: _imem06_rd = 1;
    5: _imem06_rd = 1;
    4: _imem06_rd = 1;
    3: _imem06_rd = 1;
    2: _imem06_rd = 1;
    1: _imem06_rd = 1;
    13: _imem06_rd = 1;
    12: _imem06_rd = 1;
    11: _imem06_rd = 1;
    10: _imem06_rd = 1;
    0: _imem06_rd = 1;
    24: _imem06_rd = 1;
    23: _imem06_rd = 1;
    22: _imem06_rd = 1;
    21: _imem06_rd = 1;
    20: _imem06_rd = 1;
    19: _imem06_rd = 1;
    18: _imem06_rd = 1;
    17: _imem06_rd = 1;
    16: _imem06_rd = 1;
    15: _imem06_rd = 1;
    14: _imem06_rd = 1;
    37: _imem06_rd = 1;
    36: _imem06_rd = 1;
    35: _imem06_rd = 1;
    43: _imem06_rd = 1;
    42: _imem06_rd = 1;
    41: _imem06_rd = 1;
    40: _imem06_rd = 1;
    39: _imem06_rd = 1;
    38: _imem06_rd = 1;
    34: _imem06_rd = 1;
    33: _imem06_rd = 1;
    32: _imem06_rd = 1;
    31: _imem06_rd = 1;
    30: _imem06_rd = 1;
    29: _imem06_rd = 1;
    28: _imem06_rd = 1;
    27: _imem06_rd = 1;
    26: _imem06_rd = 1;
    25: _imem06_rd = 1;
    47: _imem06_rd = 1;
    46: _imem06_rd = 1;
    45: _imem06_rd = 1;
    44: _imem06_rd = 1;
    50: _imem06_rd = 1;
    49: _imem06_rd = 1;
    48: _imem06_rd = 1;
    65: _imem06_rd = 1;
    64: _imem06_rd = 1;
    63: _imem06_rd = 1;
    62: _imem06_rd = 1;
    61: _imem06_rd = 1;
    60: _imem06_rd = 1;
    59: _imem06_rd = 1;
    58: _imem06_rd = 1;
    57: _imem06_rd = 1;
    56: _imem06_rd = 1;
    55: _imem06_rd = 1;
    54: _imem06_rd = 1;
    53: _imem06_rd = 1;
    52: _imem06_rd = 1;
    51: _imem06_rd = 1;
    70: _imem06_rd = 1;
    69: _imem06_rd = 1;
    68: _imem06_rd = 1;
    67: _imem06_rd = 1;
    66: _imem06_rd = 1;
    76: _imem06_rd = 1;
    75: _imem06_rd = 1;
    74: _imem06_rd = 1;
    73: _imem06_rd = 1;
    72: _imem06_rd = 1;
    71: _imem06_rd = 1;
    77: _imem06_rd = 1;
    78: _imem06_rd = 1;
    87: _imem06_rd = 1;
    86: _imem06_rd = 1;
    85: _imem06_rd = 1;
    79: _imem06_rd = 1;
    80: _imem06_rd = 1;
    81: _imem06_rd = 1;
    82: _imem06_rd = 1;
    84: _imem06_rd = 1;
    83: _imem06_rd = 1;
    88: _imem06_rd = 1;
    89: _imem06_rd = 1;
    90: _imem06_rd = 1;
    91: _imem06_rd = 1;
    92: _imem06_rd = 1;
    93: _imem06_rd = 1;
    94: _imem06_rd = 1;
    95: _imem06_rd = 1;
    96: _imem06_rd = 1;
    97: _imem06_rd = 1;
    98: _imem06_rd = 1;
    99: _imem06_rd = 1;
    100: _imem06_rd = 1;
    101: _imem06_rd = 1;
    102: _imem06_rd = 1;
    103: _imem06_rd = 1;
    104: _imem06_rd = 1;
    105: _imem06_rd = 1;
    106: _imem06_rd = 1;
    107: _imem06_rd = 1;
    108: _imem06_rd = 1;
    109: _imem06_rd = 1;
    110: _imem06_rd = 1;
    111: _imem06_rd = 1;
    112: _imem06_rd = 1;
    113: _imem06_rd = 1;
    114: _imem06_rd = 1;
    115: _imem06_rd = 1;
    116: _imem06_rd = 1;
    117: _imem06_rd = 1;
    118: _imem06_rd = 1;
    119: _imem06_rd = 1;
    120: _imem06_rd = 1;
    121: _imem06_rd = 1;
    122: _imem06_rd = 1;
    123: _imem06_rd = 1;
    124: _imem06_rd = 1;
    125: _imem06_rd = 1;
    126: _imem06_rd = 1;
    127: _imem06_rd = 1;
    128: _imem06_rd = 1;
    129: _imem06_rd = 1;
    default: _imem06_rd = 0;
    endcase
  end // always @ ( * )
  assign imem06_rd = _imem06_rd;

  // 7番目の入力用メモリブロックの制御
  reg [4:0] _imem07_bank;
  always @ ( * ) begin
    case ( state )
    13: _imem07_bank = 0;
    12: _imem07_bank = 1;
    11: _imem07_bank = 6;
    10: _imem07_bank = 7;
    9: _imem07_bank = 8;
    8: _imem07_bank = 11;
    7: _imem07_bank = 14;
    6: _imem07_bank = 15;
    5: _imem07_bank = 19;
    4: _imem07_bank = 24;
    3: _imem07_bank = 28;
    2: _imem07_bank = 29;
    19: _imem07_bank = 2;
    18: _imem07_bank = 7;
    17: _imem07_bank = 9;
    16: _imem07_bank = 10;
    15: _imem07_bank = 11;
    14: _imem07_bank = 18;
    1: _imem07_bank = 25;
    0: _imem07_bank = 27;
    43: _imem07_bank = 0;
    42: _imem07_bank = 1;
    41: _imem07_bank = 8;
    40: _imem07_bank = 9;
    39: _imem07_bank = 10;
    38: _imem07_bank = 12;
    37: _imem07_bank = 14;
    36: _imem07_bank = 15;
    35: _imem07_bank = 20;
    22: _imem07_bank = 23;
    21: _imem07_bank = 25;
    20: _imem07_bank = 26;
    44: _imem07_bank = 2;
    34: _imem07_bank = 7;
    33: _imem07_bank = 11;
    32: _imem07_bank = 17;
    31: _imem07_bank = 22;
    30: _imem07_bank = 23;
    29: _imem07_bank = 26;
    28: _imem07_bank = 27;
    27: _imem07_bank = 29;
    26: _imem07_bank = 30;
    46: _imem07_bank = 0;
    45: _imem07_bank = 4;
    25: _imem07_bank = 16;
    24: _imem07_bank = 19;
    23: _imem07_bank = 21;
    65: _imem07_bank = 0;
    64: _imem07_bank = 3;
    63: _imem07_bank = 7;
    62: _imem07_bank = 8;
    61: _imem07_bank = 11;
    47: _imem07_bank = 13;
    70: _imem07_bank = 0;
    69: _imem07_bank = 1;
    68: _imem07_bank = 2;
    67: _imem07_bank = 3;
    66: _imem07_bank = 4;
    60: _imem07_bank = 5;
    59: _imem07_bank = 6;
    51: _imem07_bank = 0;
    50: _imem07_bank = 1;
    49: _imem07_bank = 2;
    48: _imem07_bank = 3;
    52: _imem07_bank = 31;
    76: _imem07_bank = 0;
    75: _imem07_bank = 1;
    56: _imem07_bank = 2;
    55: _imem07_bank = 3;
    54: _imem07_bank = 4;
    53: _imem07_bank = 5;
    71: _imem07_bank = 0;
    58: _imem07_bank = 9;
    57: _imem07_bank = 14;
    72: _imem07_bank = 1;
    73: _imem07_bank = 3;
    74: _imem07_bank = 3;
    77: _imem07_bank = 1;
    78: _imem07_bank = 1;
    79: _imem07_bank = 1;
    80: _imem07_bank = 2;
    81: _imem07_bank = 3;
    82: _imem07_bank = 2;
    83: _imem07_bank = 0;
    88: _imem07_bank = 0;
    87: _imem07_bank = 3;
    86: _imem07_bank = 5;
    85: _imem07_bank = 8;
    84: _imem07_bank = 10;
    89: _imem07_bank = 0;
    90: _imem07_bank = 1;
    91: _imem07_bank = 1;
    92: _imem07_bank = 0;
    93: _imem07_bank = 5;
    94: _imem07_bank = 0;
    95: _imem07_bank = 0;
    96: _imem07_bank = 0;
    97: _imem07_bank = 1;
    98: _imem07_bank = 0;
    99: _imem07_bank = 0;
    100: _imem07_bank = 0;
    101: _imem07_bank = 2;
    102: _imem07_bank = 1;
    103: _imem07_bank = 1;
    104: _imem07_bank = 0;
    105: _imem07_bank = 0;
    106: _imem07_bank = 0;
    107: _imem07_bank = 0;
    108: _imem07_bank = 0;
    109: _imem07_bank = 3;
    110: _imem07_bank = 0;
    111: _imem07_bank = 4;
    112: _imem07_bank = 0;
    113: _imem07_bank = 1;
    114: _imem07_bank = 2;
    115: _imem07_bank = 0;
    116: _imem07_bank = 26;
    117: _imem07_bank = 28;
    118: _imem07_bank = 1;
    119: _imem07_bank = 0;
    120: _imem07_bank = 2;
    121: _imem07_bank = 2;
    122: _imem07_bank = 0;
    123: _imem07_bank = 7;
    124: _imem07_bank = 0;
    125: _imem07_bank = 29;
    126: _imem07_bank = 1;
    127: _imem07_bank = 2;
    128: _imem07_bank = 0;
    129: _imem07_bank = 1;
    default: _imem07_bank = 0;
    endcase
  end // always @ ( * )
  assign imem07_bank = _imem07_bank;
  reg _imem07_rd;
  always @ ( * ) begin
    case ( state )
    13: _imem07_rd = 1;
    12: _imem07_rd = 1;
    11: _imem07_rd = 1;
    10: _imem07_rd = 1;
    9: _imem07_rd = 1;
    8: _imem07_rd = 1;
    7: _imem07_rd = 1;
    6: _imem07_rd = 1;
    5: _imem07_rd = 1;
    4: _imem07_rd = 1;
    3: _imem07_rd = 1;
    2: _imem07_rd = 1;
    19: _imem07_rd = 1;
    18: _imem07_rd = 1;
    17: _imem07_rd = 1;
    16: _imem07_rd = 1;
    15: _imem07_rd = 1;
    14: _imem07_rd = 1;
    1: _imem07_rd = 1;
    0: _imem07_rd = 1;
    43: _imem07_rd = 1;
    42: _imem07_rd = 1;
    41: _imem07_rd = 1;
    40: _imem07_rd = 1;
    39: _imem07_rd = 1;
    38: _imem07_rd = 1;
    37: _imem07_rd = 1;
    36: _imem07_rd = 1;
    35: _imem07_rd = 1;
    22: _imem07_rd = 1;
    21: _imem07_rd = 1;
    20: _imem07_rd = 1;
    44: _imem07_rd = 1;
    34: _imem07_rd = 1;
    33: _imem07_rd = 1;
    32: _imem07_rd = 1;
    31: _imem07_rd = 1;
    30: _imem07_rd = 1;
    29: _imem07_rd = 1;
    28: _imem07_rd = 1;
    27: _imem07_rd = 1;
    26: _imem07_rd = 1;
    46: _imem07_rd = 1;
    45: _imem07_rd = 1;
    25: _imem07_rd = 1;
    24: _imem07_rd = 1;
    23: _imem07_rd = 1;
    65: _imem07_rd = 1;
    64: _imem07_rd = 1;
    63: _imem07_rd = 1;
    62: _imem07_rd = 1;
    61: _imem07_rd = 1;
    47: _imem07_rd = 1;
    70: _imem07_rd = 1;
    69: _imem07_rd = 1;
    68: _imem07_rd = 1;
    67: _imem07_rd = 1;
    66: _imem07_rd = 1;
    60: _imem07_rd = 1;
    59: _imem07_rd = 1;
    51: _imem07_rd = 1;
    50: _imem07_rd = 1;
    49: _imem07_rd = 1;
    48: _imem07_rd = 1;
    52: _imem07_rd = 1;
    76: _imem07_rd = 1;
    75: _imem07_rd = 1;
    56: _imem07_rd = 1;
    55: _imem07_rd = 1;
    54: _imem07_rd = 1;
    53: _imem07_rd = 1;
    71: _imem07_rd = 1;
    58: _imem07_rd = 1;
    57: _imem07_rd = 1;
    72: _imem07_rd = 1;
    73: _imem07_rd = 1;
    74: _imem07_rd = 1;
    77: _imem07_rd = 1;
    78: _imem07_rd = 1;
    79: _imem07_rd = 1;
    80: _imem07_rd = 1;
    81: _imem07_rd = 1;
    82: _imem07_rd = 1;
    83: _imem07_rd = 1;
    88: _imem07_rd = 1;
    87: _imem07_rd = 1;
    86: _imem07_rd = 1;
    85: _imem07_rd = 1;
    84: _imem07_rd = 1;
    89: _imem07_rd = 1;
    90: _imem07_rd = 1;
    91: _imem07_rd = 1;
    92: _imem07_rd = 1;
    93: _imem07_rd = 1;
    94: _imem07_rd = 1;
    95: _imem07_rd = 1;
    96: _imem07_rd = 1;
    97: _imem07_rd = 1;
    98: _imem07_rd = 1;
    99: _imem07_rd = 1;
    100: _imem07_rd = 1;
    101: _imem07_rd = 1;
    102: _imem07_rd = 1;
    103: _imem07_rd = 1;
    104: _imem07_rd = 1;
    105: _imem07_rd = 1;
    106: _imem07_rd = 1;
    107: _imem07_rd = 1;
    108: _imem07_rd = 1;
    109: _imem07_rd = 1;
    110: _imem07_rd = 1;
    111: _imem07_rd = 1;
    112: _imem07_rd = 1;
    113: _imem07_rd = 1;
    114: _imem07_rd = 1;
    115: _imem07_rd = 1;
    116: _imem07_rd = 1;
    117: _imem07_rd = 1;
    118: _imem07_rd = 1;
    119: _imem07_rd = 1;
    120: _imem07_rd = 1;
    121: _imem07_rd = 1;
    122: _imem07_rd = 1;
    123: _imem07_rd = 1;
    124: _imem07_rd = 1;
    125: _imem07_rd = 1;
    126: _imem07_rd = 1;
    127: _imem07_rd = 1;
    128: _imem07_rd = 1;
    129: _imem07_rd = 1;
    default: _imem07_rd = 0;
    endcase
  end // always @ ( * )
  assign imem07_rd = _imem07_rd;

  // 0番目の出力用メモリブロックの制御
  reg [5:0] _omem00_bank;
  always @ ( * ) begin
    case ( state )
    22: _omem00_bank = 0;
    37: _omem00_bank = 1;
    47: _omem00_bank = 2;
    54: _omem00_bank = 3;
    60: _omem00_bank = 4;
    69: _omem00_bank = 5;
    78: _omem00_bank = 6;
    70: _omem00_bank = 7;
    89: _omem00_bank = 8;
    75: _omem00_bank = 9;
    88: _omem00_bank = 10;
    74: _omem00_bank = 11;
    90: _omem00_bank = 12;
    76: _omem00_bank = 13;
    91: _omem00_bank = 14;
    92: _omem00_bank = 15;
    93: _omem00_bank = 16;
    94: _omem00_bank = 17;
    95: _omem00_bank = 18;
    71: _omem00_bank = 19;
    96: _omem00_bank = 20;
    77: _omem00_bank = 21;
    97: _omem00_bank = 22;
    79: _omem00_bank = 23;
    80: _omem00_bank = 24;
    98: _omem00_bank = 25;
    99: _omem00_bank = 26;
    81: _omem00_bank = 27;
    82: _omem00_bank = 28;
    100: _omem00_bank = 29;
    101: _omem00_bank = 30;
    83: _omem00_bank = 31;
    102: _omem00_bank = 32;
    84: _omem00_bank = 33;
    103: _omem00_bank = 34;
    85: _omem00_bank = 35;
    104: _omem00_bank = 36;
    86: _omem00_bank = 37;
    87: _omem00_bank = 38;
    105: _omem00_bank = 39;
    106: _omem00_bank = 40;
    107: _omem00_bank = 41;
    108: _omem00_bank = 42;
    109: _omem00_bank = 43;
    110: _omem00_bank = 44;
    111: _omem00_bank = 45;
    112: _omem00_bank = 46;
    113: _omem00_bank = 47;
    114: _omem00_bank = 48;
    115: _omem00_bank = 49;
    116: _omem00_bank = 50;
    117: _omem00_bank = 51;
    62: _omem00_bank = 52;
    118: _omem00_bank = 53;
    119: _omem00_bank = 54;
    73: _omem00_bank = 55;
    120: _omem00_bank = 56;
    121: _omem00_bank = 57;
    122: _omem00_bank = 58;
    123: _omem00_bank = 59;
    default: _omem00_bank = 0;
    endcase
  end // always @ ( * )
  assign omem00_bank = _omem00_bank;
  reg _omem00_wr;
  always @ ( * ) begin
    case ( state )
    22: _omem00_wr = 1;
    37: _omem00_wr = 1;
    47: _omem00_wr = 1;
    54: _omem00_wr = 1;
    60: _omem00_wr = 1;
    69: _omem00_wr = 1;
    78: _omem00_wr = 1;
    70: _omem00_wr = 1;
    89: _omem00_wr = 1;
    75: _omem00_wr = 1;
    88: _omem00_wr = 1;
    74: _omem00_wr = 1;
    90: _omem00_wr = 1;
    76: _omem00_wr = 1;
    91: _omem00_wr = 1;
    92: _omem00_wr = 1;
    93: _omem00_wr = 1;
    94: _omem00_wr = 1;
    95: _omem00_wr = 1;
    71: _omem00_wr = 1;
    96: _omem00_wr = 1;
    77: _omem00_wr = 1;
    97: _omem00_wr = 1;
    79: _omem00_wr = 1;
    80: _omem00_wr = 1;
    98: _omem00_wr = 1;
    99: _omem00_wr = 1;
    81: _omem00_wr = 1;
    82: _omem00_wr = 1;
    100: _omem00_wr = 1;
    101: _omem00_wr = 1;
    83: _omem00_wr = 1;
    102: _omem00_wr = 1;
    84: _omem00_wr = 1;
    103: _omem00_wr = 1;
    85: _omem00_wr = 1;
    104: _omem00_wr = 1;
    86: _omem00_wr = 1;
    87: _omem00_wr = 1;
    105: _omem00_wr = 1;
    106: _omem00_wr = 1;
    107: _omem00_wr = 1;
    108: _omem00_wr = 1;
    109: _omem00_wr = 1;
    110: _omem00_wr = 1;
    111: _omem00_wr = 1;
    112: _omem00_wr = 1;
    113: _omem00_wr = 1;
    114: _omem00_wr = 1;
    115: _omem00_wr = 1;
    116: _omem00_wr = 1;
    117: _omem00_wr = 1;
    62: _omem00_wr = 1;
    118: _omem00_wr = 1;
    119: _omem00_wr = 1;
    73: _omem00_wr = 1;
    120: _omem00_wr = 1;
    121: _omem00_wr = 1;
    122: _omem00_wr = 1;
    123: _omem00_wr = 1;
    default: _omem00_wr = 0;
    endcase
  end // always @ ( * )
  assign omem00_wr = _omem00_wr;

  // 1番目の出力用メモリブロックの制御
  reg [5:0] _omem01_bank;
  always @ ( * ) begin
    case ( state )
    89: _omem01_bank = 0;
    78: _omem01_bank = 1;
    73: _omem01_bank = 2;
    90: _omem01_bank = 3;
    79: _omem01_bank = 4;
    91: _omem01_bank = 5;
    80: _omem01_bank = 6;
    92: _omem01_bank = 7;
    93: _omem01_bank = 8;
    81: _omem01_bank = 9;
    94: _omem01_bank = 10;
    82: _omem01_bank = 11;
    95: _omem01_bank = 12;
    83: _omem01_bank = 13;
    96: _omem01_bank = 14;
    84: _omem01_bank = 15;
    85: _omem01_bank = 16;
    86: _omem01_bank = 17;
    97: _omem01_bank = 18;
    98: _omem01_bank = 19;
    99: _omem01_bank = 20;
    87: _omem01_bank = 21;
    88: _omem01_bank = 22;
    100: _omem01_bank = 23;
    101: _omem01_bank = 24;
    102: _omem01_bank = 25;
    103: _omem01_bank = 26;
    104: _omem01_bank = 27;
    105: _omem01_bank = 28;
    106: _omem01_bank = 29;
    107: _omem01_bank = 30;
    108: _omem01_bank = 31;
    109: _omem01_bank = 32;
    110: _omem01_bank = 33;
    111: _omem01_bank = 34;
    112: _omem01_bank = 35;
    113: _omem01_bank = 36;
    114: _omem01_bank = 37;
    115: _omem01_bank = 38;
    116: _omem01_bank = 39;
    117: _omem01_bank = 40;
    118: _omem01_bank = 41;
    119: _omem01_bank = 42;
    120: _omem01_bank = 43;
    121: _omem01_bank = 44;
    122: _omem01_bank = 45;
    123: _omem01_bank = 46;
    124: _omem01_bank = 47;
    125: _omem01_bank = 48;
    126: _omem01_bank = 49;
    127: _omem01_bank = 50;
    128: _omem01_bank = 51;
    129: _omem01_bank = 52;
    130: _omem01_bank = 53;
    131: _omem01_bank = 54;
    132: _omem01_bank = 55;
    133: _omem01_bank = 56;
    134: _omem01_bank = 57;
    135: _omem01_bank = 58;
    136: _omem01_bank = 59;
    default: _omem01_bank = 0;
    endcase
  end // always @ ( * )
  assign omem01_bank = _omem01_bank;
  reg _omem01_wr;
  always @ ( * ) begin
    case ( state )
    89: _omem01_wr = 1;
    78: _omem01_wr = 1;
    73: _omem01_wr = 1;
    90: _omem01_wr = 1;
    79: _omem01_wr = 1;
    91: _omem01_wr = 1;
    80: _omem01_wr = 1;
    92: _omem01_wr = 1;
    93: _omem01_wr = 1;
    81: _omem01_wr = 1;
    94: _omem01_wr = 1;
    82: _omem01_wr = 1;
    95: _omem01_wr = 1;
    83: _omem01_wr = 1;
    96: _omem01_wr = 1;
    84: _omem01_wr = 1;
    85: _omem01_wr = 1;
    86: _omem01_wr = 1;
    97: _omem01_wr = 1;
    98: _omem01_wr = 1;
    99: _omem01_wr = 1;
    87: _omem01_wr = 1;
    88: _omem01_wr = 1;
    100: _omem01_wr = 1;
    101: _omem01_wr = 1;
    102: _omem01_wr = 1;
    103: _omem01_wr = 1;
    104: _omem01_wr = 1;
    105: _omem01_wr = 1;
    106: _omem01_wr = 1;
    107: _omem01_wr = 1;
    108: _omem01_wr = 1;
    109: _omem01_wr = 1;
    110: _omem01_wr = 1;
    111: _omem01_wr = 1;
    112: _omem01_wr = 1;
    113: _omem01_wr = 1;
    114: _omem01_wr = 1;
    115: _omem01_wr = 1;
    116: _omem01_wr = 1;
    117: _omem01_wr = 1;
    118: _omem01_wr = 1;
    119: _omem01_wr = 1;
    120: _omem01_wr = 1;
    121: _omem01_wr = 1;
    122: _omem01_wr = 1;
    123: _omem01_wr = 1;
    124: _omem01_wr = 1;
    125: _omem01_wr = 1;
    126: _omem01_wr = 1;
    127: _omem01_wr = 1;
    128: _omem01_wr = 1;
    129: _omem01_wr = 1;
    130: _omem01_wr = 1;
    131: _omem01_wr = 1;
    132: _omem01_wr = 1;
    133: _omem01_wr = 1;
    134: _omem01_wr = 1;
    135: _omem01_wr = 1;
    136: _omem01_wr = 1;
    default: _omem01_wr = 0;
    endcase
  end // always @ ( * )
  assign omem01_wr = _omem01_wr;

  // 2番目の出力用メモリブロックの制御
  reg [5:0] _omem02_bank;
  always @ ( * ) begin
    case ( state )
    91: _omem02_bank = 0;
    84: _omem02_bank = 1;
    92: _omem02_bank = 2;
    93: _omem02_bank = 3;
    94: _omem02_bank = 4;
    85: _omem02_bank = 5;
    86: _omem02_bank = 6;
    95: _omem02_bank = 7;
    87: _omem02_bank = 8;
    88: _omem02_bank = 9;
    66: _omem02_bank = 10;
    96: _omem02_bank = 11;
    97: _omem02_bank = 12;
    98: _omem02_bank = 13;
    89: _omem02_bank = 14;
    99: _omem02_bank = 15;
    90: _omem02_bank = 16;
    100: _omem02_bank = 17;
    101: _omem02_bank = 18;
    102: _omem02_bank = 19;
    103: _omem02_bank = 20;
    104: _omem02_bank = 21;
    105: _omem02_bank = 22;
    106: _omem02_bank = 23;
    107: _omem02_bank = 24;
    108: _omem02_bank = 25;
    109: _omem02_bank = 26;
    110: _omem02_bank = 27;
    111: _omem02_bank = 28;
    112: _omem02_bank = 29;
    113: _omem02_bank = 30;
    114: _omem02_bank = 31;
    115: _omem02_bank = 32;
    116: _omem02_bank = 33;
    117: _omem02_bank = 34;
    118: _omem02_bank = 35;
    119: _omem02_bank = 36;
    120: _omem02_bank = 37;
    121: _omem02_bank = 38;
    122: _omem02_bank = 39;
    123: _omem02_bank = 40;
    124: _omem02_bank = 41;
    125: _omem02_bank = 42;
    126: _omem02_bank = 43;
    127: _omem02_bank = 44;
    128: _omem02_bank = 45;
    129: _omem02_bank = 46;
    130: _omem02_bank = 47;
    131: _omem02_bank = 48;
    132: _omem02_bank = 49;
    133: _omem02_bank = 50;
    134: _omem02_bank = 51;
    135: _omem02_bank = 52;
    136: _omem02_bank = 53;
    137: _omem02_bank = 54;
    138: _omem02_bank = 55;
    139: _omem02_bank = 56;
    140: _omem02_bank = 57;
    141: _omem02_bank = 58;
    142: _omem02_bank = 59;
    default: _omem02_bank = 0;
    endcase
  end // always @ ( * )
  assign omem02_bank = _omem02_bank;
  reg _omem02_wr;
  always @ ( * ) begin
    case ( state )
    91: _omem02_wr = 1;
    84: _omem02_wr = 1;
    92: _omem02_wr = 1;
    93: _omem02_wr = 1;
    94: _omem02_wr = 1;
    85: _omem02_wr = 1;
    86: _omem02_wr = 1;
    95: _omem02_wr = 1;
    87: _omem02_wr = 1;
    88: _omem02_wr = 1;
    66: _omem02_wr = 1;
    96: _omem02_wr = 1;
    97: _omem02_wr = 1;
    98: _omem02_wr = 1;
    89: _omem02_wr = 1;
    99: _omem02_wr = 1;
    90: _omem02_wr = 1;
    100: _omem02_wr = 1;
    101: _omem02_wr = 1;
    102: _omem02_wr = 1;
    103: _omem02_wr = 1;
    104: _omem02_wr = 1;
    105: _omem02_wr = 1;
    106: _omem02_wr = 1;
    107: _omem02_wr = 1;
    108: _omem02_wr = 1;
    109: _omem02_wr = 1;
    110: _omem02_wr = 1;
    111: _omem02_wr = 1;
    112: _omem02_wr = 1;
    113: _omem02_wr = 1;
    114: _omem02_wr = 1;
    115: _omem02_wr = 1;
    116: _omem02_wr = 1;
    117: _omem02_wr = 1;
    118: _omem02_wr = 1;
    119: _omem02_wr = 1;
    120: _omem02_wr = 1;
    121: _omem02_wr = 1;
    122: _omem02_wr = 1;
    123: _omem02_wr = 1;
    124: _omem02_wr = 1;
    125: _omem02_wr = 1;
    126: _omem02_wr = 1;
    127: _omem02_wr = 1;
    128: _omem02_wr = 1;
    129: _omem02_wr = 1;
    130: _omem02_wr = 1;
    131: _omem02_wr = 1;
    132: _omem02_wr = 1;
    133: _omem02_wr = 1;
    134: _omem02_wr = 1;
    135: _omem02_wr = 1;
    136: _omem02_wr = 1;
    137: _omem02_wr = 1;
    138: _omem02_wr = 1;
    139: _omem02_wr = 1;
    140: _omem02_wr = 1;
    141: _omem02_wr = 1;
    142: _omem02_wr = 1;
    default: _omem02_wr = 0;
    endcase
  end // always @ ( * )
  assign omem02_wr = _omem02_wr;

  // 3番目の出力用メモリブロックの制御
  reg [5:0] _omem03_bank;
  always @ ( * ) begin
    case ( state )
    100: _omem03_bank = 0;
    101: _omem03_bank = 1;
    102: _omem03_bank = 2;
    103: _omem03_bank = 3;
    104: _omem03_bank = 4;
    105: _omem03_bank = 5;
    106: _omem03_bank = 6;
    107: _omem03_bank = 7;
    108: _omem03_bank = 8;
    109: _omem03_bank = 9;
    110: _omem03_bank = 10;
    111: _omem03_bank = 11;
    112: _omem03_bank = 12;
    113: _omem03_bank = 13;
    114: _omem03_bank = 14;
    115: _omem03_bank = 15;
    116: _omem03_bank = 16;
    117: _omem03_bank = 17;
    118: _omem03_bank = 18;
    119: _omem03_bank = 19;
    120: _omem03_bank = 20;
    121: _omem03_bank = 21;
    122: _omem03_bank = 22;
    123: _omem03_bank = 23;
    124: _omem03_bank = 24;
    125: _omem03_bank = 25;
    126: _omem03_bank = 26;
    127: _omem03_bank = 27;
    128: _omem03_bank = 28;
    129: _omem03_bank = 29;
    130: _omem03_bank = 30;
    131: _omem03_bank = 31;
    132: _omem03_bank = 32;
    133: _omem03_bank = 33;
    134: _omem03_bank = 34;
    135: _omem03_bank = 35;
    136: _omem03_bank = 36;
    137: _omem03_bank = 37;
    138: _omem03_bank = 38;
    139: _omem03_bank = 39;
    140: _omem03_bank = 40;
    141: _omem03_bank = 41;
    142: _omem03_bank = 42;
    143: _omem03_bank = 43;
    144: _omem03_bank = 44;
    145: _omem03_bank = 45;
    146: _omem03_bank = 46;
    147: _omem03_bank = 47;
    148: _omem03_bank = 48;
    149: _omem03_bank = 49;
    150: _omem03_bank = 50;
    151: _omem03_bank = 51;
    152: _omem03_bank = 52;
    153: _omem03_bank = 53;
    154: _omem03_bank = 54;
    155: _omem03_bank = 55;
    156: _omem03_bank = 56;
    157: _omem03_bank = 57;
    158: _omem03_bank = 58;
    159: _omem03_bank = 59;
    default: _omem03_bank = 0;
    endcase
  end // always @ ( * )
  assign omem03_bank = _omem03_bank;
  reg _omem03_wr;
  always @ ( * ) begin
    case ( state )
    100: _omem03_wr = 1;
    101: _omem03_wr = 1;
    102: _omem03_wr = 1;
    103: _omem03_wr = 1;
    104: _omem03_wr = 1;
    105: _omem03_wr = 1;
    106: _omem03_wr = 1;
    107: _omem03_wr = 1;
    108: _omem03_wr = 1;
    109: _omem03_wr = 1;
    110: _omem03_wr = 1;
    111: _omem03_wr = 1;
    112: _omem03_wr = 1;
    113: _omem03_wr = 1;
    114: _omem03_wr = 1;
    115: _omem03_wr = 1;
    116: _omem03_wr = 1;
    117: _omem03_wr = 1;
    118: _omem03_wr = 1;
    119: _omem03_wr = 1;
    120: _omem03_wr = 1;
    121: _omem03_wr = 1;
    122: _omem03_wr = 1;
    123: _omem03_wr = 1;
    124: _omem03_wr = 1;
    125: _omem03_wr = 1;
    126: _omem03_wr = 1;
    127: _omem03_wr = 1;
    128: _omem03_wr = 1;
    129: _omem03_wr = 1;
    130: _omem03_wr = 1;
    131: _omem03_wr = 1;
    132: _omem03_wr = 1;
    133: _omem03_wr = 1;
    134: _omem03_wr = 1;
    135: _omem03_wr = 1;
    136: _omem03_wr = 1;
    137: _omem03_wr = 1;
    138: _omem03_wr = 1;
    139: _omem03_wr = 1;
    140: _omem03_wr = 1;
    141: _omem03_wr = 1;
    142: _omem03_wr = 1;
    143: _omem03_wr = 1;
    144: _omem03_wr = 1;
    145: _omem03_wr = 1;
    146: _omem03_wr = 1;
    147: _omem03_wr = 1;
    148: _omem03_wr = 1;
    149: _omem03_wr = 1;
    150: _omem03_wr = 1;
    151: _omem03_wr = 1;
    152: _omem03_wr = 1;
    153: _omem03_wr = 1;
    154: _omem03_wr = 1;
    155: _omem03_wr = 1;
    156: _omem03_wr = 1;
    157: _omem03_wr = 1;
    158: _omem03_wr = 1;
    159: _omem03_wr = 1;
    default: _omem03_wr = 0;
    endcase
  end // always @ ( * )
  assign omem03_wr = _omem03_wr;

  // 4番目の出力用メモリブロックの制御
  reg [5:0] _omem04_bank;
  always @ ( * ) begin
    case ( state )
    117: _omem04_bank = 0;
    118: _omem04_bank = 1;
    119: _omem04_bank = 2;
    120: _omem04_bank = 3;
    121: _omem04_bank = 4;
    122: _omem04_bank = 5;
    123: _omem04_bank = 6;
    124: _omem04_bank = 7;
    125: _omem04_bank = 8;
    126: _omem04_bank = 9;
    127: _omem04_bank = 10;
    128: _omem04_bank = 11;
    129: _omem04_bank = 12;
    130: _omem04_bank = 13;
    131: _omem04_bank = 14;
    132: _omem04_bank = 15;
    133: _omem04_bank = 16;
    134: _omem04_bank = 17;
    135: _omem04_bank = 18;
    136: _omem04_bank = 19;
    137: _omem04_bank = 20;
    138: _omem04_bank = 21;
    139: _omem04_bank = 22;
    140: _omem04_bank = 23;
    141: _omem04_bank = 24;
    142: _omem04_bank = 25;
    143: _omem04_bank = 26;
    144: _omem04_bank = 27;
    145: _omem04_bank = 28;
    146: _omem04_bank = 29;
    147: _omem04_bank = 30;
    148: _omem04_bank = 31;
    149: _omem04_bank = 32;
    150: _omem04_bank = 33;
    151: _omem04_bank = 34;
    152: _omem04_bank = 35;
    153: _omem04_bank = 36;
    154: _omem04_bank = 37;
    155: _omem04_bank = 38;
    156: _omem04_bank = 39;
    157: _omem04_bank = 40;
    158: _omem04_bank = 41;
    159: _omem04_bank = 42;
    160: _omem04_bank = 43;
    161: _omem04_bank = 44;
    162: _omem04_bank = 45;
    163: _omem04_bank = 46;
    164: _omem04_bank = 47;
    165: _omem04_bank = 48;
    166: _omem04_bank = 49;
    167: _omem04_bank = 50;
    168: _omem04_bank = 51;
    169: _omem04_bank = 52;
    170: _omem04_bank = 53;
    171: _omem04_bank = 54;
    172: _omem04_bank = 55;
    173: _omem04_bank = 56;
    174: _omem04_bank = 57;
    default: _omem04_bank = 0;
    endcase
  end // always @ ( * )
  assign omem04_bank = _omem04_bank;
  reg _omem04_wr;
  always @ ( * ) begin
    case ( state )
    117: _omem04_wr = 1;
    118: _omem04_wr = 1;
    119: _omem04_wr = 1;
    120: _omem04_wr = 1;
    121: _omem04_wr = 1;
    122: _omem04_wr = 1;
    123: _omem04_wr = 1;
    124: _omem04_wr = 1;
    125: _omem04_wr = 1;
    126: _omem04_wr = 1;
    127: _omem04_wr = 1;
    128: _omem04_wr = 1;
    129: _omem04_wr = 1;
    130: _omem04_wr = 1;
    131: _omem04_wr = 1;
    132: _omem04_wr = 1;
    133: _omem04_wr = 1;
    134: _omem04_wr = 1;
    135: _omem04_wr = 1;
    136: _omem04_wr = 1;
    137: _omem04_wr = 1;
    138: _omem04_wr = 1;
    139: _omem04_wr = 1;
    140: _omem04_wr = 1;
    141: _omem04_wr = 1;
    142: _omem04_wr = 1;
    143: _omem04_wr = 1;
    144: _omem04_wr = 1;
    145: _omem04_wr = 1;
    146: _omem04_wr = 1;
    147: _omem04_wr = 1;
    148: _omem04_wr = 1;
    149: _omem04_wr = 1;
    150: _omem04_wr = 1;
    151: _omem04_wr = 1;
    152: _omem04_wr = 1;
    153: _omem04_wr = 1;
    154: _omem04_wr = 1;
    155: _omem04_wr = 1;
    156: _omem04_wr = 1;
    157: _omem04_wr = 1;
    158: _omem04_wr = 1;
    159: _omem04_wr = 1;
    160: _omem04_wr = 1;
    161: _omem04_wr = 1;
    162: _omem04_wr = 1;
    163: _omem04_wr = 1;
    164: _omem04_wr = 1;
    165: _omem04_wr = 1;
    166: _omem04_wr = 1;
    167: _omem04_wr = 1;
    168: _omem04_wr = 1;
    169: _omem04_wr = 1;
    170: _omem04_wr = 1;
    171: _omem04_wr = 1;
    172: _omem04_wr = 1;
    173: _omem04_wr = 1;
    174: _omem04_wr = 1;
    default: _omem04_wr = 0;
    endcase
  end // always @ ( * )
  assign omem04_wr = _omem04_wr;
  reg [8:0] _omem00_out;
  always @ ( * ) begin
    case ( state )
    22: _omem00_out = reg_0134;
    37: _omem00_out = reg_0325;
    47: _omem00_out = reg_0976;
    54: _omem00_out = reg_0249;
    60: _omem00_out = reg_0187;
    69: _omem00_out = reg_0600;
    78: _omem00_out = reg_0237;
    70: _omem00_out = reg_0370;
    89: _omem00_out = reg_0237;
    75: _omem00_out = reg_0600;
    88: _omem00_out = reg_0525;
    74: _omem00_out = reg_0844;
    90: _omem00_out = reg_0282;
    76: _omem00_out = reg_0605;
    91: _omem00_out = reg_0959;
    92: _omem00_out = reg_0679;
    93: _omem00_out = reg_1506;
    94: _omem00_out = reg_1507;
    95: _omem00_out = reg_0708;
    71: _omem00_out = reg_0600;
    96: _omem00_out = reg_0788;
    77: _omem00_out = reg_0991;
    97: _omem00_out = reg_0852;
    79: _omem00_out = reg_1106;
    80: _omem00_out = reg_1234;
    98: _omem00_out = reg_0874;
    99: _omem00_out = reg_0877;
    81: _omem00_out = reg_1037;
    82: _omem00_out = reg_1506;
    100: _omem00_out = reg_0898;
    101: _omem00_out = reg_0525;
    83: _omem00_out = reg_1507;
    102: _omem00_out = reg_0982;
    84: _omem00_out = reg_0844;
    103: _omem00_out = reg_1034;
    85: _omem00_out = reg_0842;
    104: _omem00_out = reg_1042;
    86: _omem00_out = reg_0959;
    87: _omem00_out = reg_0600;
    105: _omem00_out = reg_1080;
    106: _omem00_out = reg_1038;
    107: _omem00_out = reg_1062;
    108: _omem00_out = reg_0990;
    109: _omem00_out = reg_1066;
    110: _omem00_out = reg_1039;
    111: _omem00_out = reg_0283;
    112: _omem00_out = reg_1069;
    113: _omem00_out = reg_1045;
    114: _omem00_out = reg_1084;
    115: _omem00_out = reg_1085;
    116: _omem00_out = reg_1086;
    117: _omem00_out = reg_1087;
    62: _omem00_out = reg_0187;
    118: _omem00_out = reg_0605;
    119: _omem00_out = reg_1103;
    73: _omem00_out = reg_0600;
    120: _omem00_out = reg_0997;
    121: _omem00_out = reg_1110;
    122: _omem00_out = reg_1186;
    123: _omem00_out = reg_1212;
    default: _omem00_out = 0;
    endcase
  end // always @ ( * )
  assign omem00_out = _omem00_out[8:0];
  reg [8:0] _omem01_out;
  always @ ( * ) begin
    case ( state )
    89: _omem01_out = reg_0322;
    78: _omem01_out = reg_0422;
    73: _omem01_out = reg_0605;
    90: _omem01_out = reg_0475;
    79: _omem01_out = reg_0540;
    91: _omem01_out = reg_0834;
    80: _omem01_out = reg_0587;
    92: _omem01_out = reg_0893;
    93: _omem01_out = reg_0942;
    81: _omem01_out = reg_0594;
    94: _omem01_out = reg_0943;
    82: _omem01_out = reg_0991;
    95: _omem01_out = reg_0652;
    83: _omem01_out = reg_0596;
    96: _omem01_out = reg_0678;
    84: _omem01_out = reg_0644;
    85: _omem01_out = reg_0237;
    86: _omem01_out = reg_0675;
    97: _omem01_out = reg_0596;
    98: _omem01_out = reg_0683;
    99: _omem01_out = reg_0756;
    87: _omem01_out = reg_0755;
    88: _omem01_out = reg_0933;
    100: _omem01_out = reg_0980;
    101: _omem01_out = reg_0761;
    102: _omem01_out = reg_0565;
    103: _omem01_out = reg_1106;
    104: _omem01_out = reg_0853;
    105: _omem01_out = reg_0680;
    106: _omem01_out = reg_0910;
    107: _omem01_out = reg_0704;
    108: _omem01_out = reg_0936;
    109: _omem01_out = reg_0941;
    110: _omem01_out = reg_0540;
    111: _omem01_out = reg_1005;
    112: _omem01_out = reg_0933;
    113: _omem01_out = reg_0587;
    114: _omem01_out = reg_0944;
    115: _omem01_out = reg_0981;
    116: _omem01_out = reg_0567;
    117: _omem01_out = reg_1234;
    118: _omem01_out = reg_0646;
    119: _omem01_out = reg_0674;
    120: _omem01_out = reg_0988;
    121: _omem01_out = reg_0422;
    122: _omem01_out = reg_1011;
    123: _omem01_out = reg_1088;
    124: _omem01_out = reg_0844;
    125: _omem01_out = reg_0671;
    126: _omem01_out = reg_0976;
    127: _omem01_out = reg_0594;
    128: _omem01_out = reg_0676;
    129: _omem01_out = reg_0280;
    130: _omem01_out = reg_0685;
    131: _omem01_out = reg_0325;
    132: _omem01_out = reg_0849;
    133: _omem01_out = reg_0713;
    134: _omem01_out = reg_0991;
    135: _omem01_out = reg_0749;
    136: _omem01_out = reg_0757;
    default: _omem01_out = 0;
    endcase
  end // always @ ( * )
  assign omem01_out = _omem01_out[8:0];
  reg [8:0] _omem02_out;
  always @ ( * ) begin
    case ( state )
    91: _omem02_out = reg_0200;
    84: _omem02_out = reg_1037;
    92: _omem02_out = reg_0265;
    93: _omem02_out = reg_0479;
    94: _omem02_out = reg_0322;
    85: _omem02_out = reg_0187;
    86: _omem02_out = reg_0282;
    95: _omem02_out = reg_0481;
    87: _omem02_out = reg_0283;
    88: _omem02_out = reg_0596;
    66: _omem02_out = reg_0369;
    96: _omem02_out = reg_0508;
    97: _omem02_out = reg_0534;
    98: _omem02_out = reg_0614;
    89: _omem02_out = reg_0844;
    99: _omem02_out = reg_0656;
    90: _omem02_out = reg_0160;
    100: _omem02_out = reg_0357;
    101: _omem02_out = reg_0187;
    102: _omem02_out = reg_0160;
    103: _omem02_out = reg_0502;
    104: _omem02_out = reg_0539;
    105: _omem02_out = reg_0842;
    106: _omem02_out = reg_0245;
    107: _omem02_out = reg_0273;
    108: _omem02_out = reg_0581;
    109: _omem02_out = reg_0639;
    110: _omem02_out = reg_0647;
    111: _omem02_out = reg_0650;
    112: _omem02_out = reg_0651;
    113: _omem02_out = reg_0200;
    114: _omem02_out = reg_0480;
    115: _omem02_out = reg_0959;
    116: _omem02_out = reg_1037;
    117: _omem02_out = reg_0644;
    118: _omem02_out = reg_0578;
    119: _omem02_out = reg_0675;
    120: _omem02_out = reg_0611;
    121: _omem02_out = reg_0679;
    122: _omem02_out = reg_0641;
    123: _omem02_out = reg_0643;
    124: _omem02_out = reg_0653;
    125: _omem02_out = reg_0655;
    126: _omem02_out = reg_0682;
    127: _omem02_out = reg_0686;
    128: _omem02_out = reg_0737;
    129: _omem02_out = reg_0237;
    130: _omem02_out = reg_0247;
    131: _omem02_out = reg_0304;
    132: _omem02_out = reg_0230;
    133: _omem02_out = reg_0652;
    134: _omem02_out = reg_0341;
    135: _omem02_out = reg_0506;
    136: _omem02_out = reg_0305;
    137: _omem02_out = reg_0508;
    138: _omem02_out = reg_0678;
    139: _omem02_out = reg_0474;
    140: _omem02_out = reg_0481;
    141: _omem02_out = reg_0504;
    142: _omem02_out = reg_0596;
    default: _omem02_out = 0;
    endcase
  end // always @ ( * )
  assign omem02_out = _omem02_out[8:0];
  reg [8:0] _omem03_out;
  always @ ( * ) begin
    case ( state )
    100: _omem03_out = reg_0509;
    101: _omem03_out = reg_0534;
    102: _omem03_out = reg_0672;
    103: _omem03_out = reg_0677;
    104: _omem03_out = reg_0683;
    105: _omem03_out = reg_0710;
    106: _omem03_out = reg_0357;
    107: _omem03_out = reg_0509;
    108: _omem03_out = reg_0657;
    109: _omem03_out = reg_0187;
    110: _omem03_out = reg_0642;
    111: _omem03_out = reg_0534;
    112: _omem03_out = reg_0656;
    113: _omem03_out = reg_0565;
    114: _omem03_out = reg_0160;
    115: _omem03_out = reg_0499;
    116: _omem03_out = reg_0753;
    117: _omem03_out = reg_1106;
    118: _omem03_out = reg_0502;
    119: _omem03_out = reg_0525;
    120: _omem03_out = reg_0490;
    121: _omem03_out = reg_0683;
    122: _omem03_out = reg_0539;
    123: _omem03_out = reg_0514;
    124: _omem03_out = reg_0842;
    125: _omem03_out = reg_0680;
    126: _omem03_out = reg_0590;
    127: _omem03_out = reg_0357;
    128: _omem03_out = reg_0121;
    129: _omem03_out = reg_0245;
    130: _omem03_out = reg_0339;
    131: _omem03_out = reg_0509;
    132: _omem03_out = reg_0755;
    133: _omem03_out = reg_0273;
    134: _omem03_out = reg_0482;
    135: _omem03_out = reg_0990;
    136: _omem03_out = reg_0657;
    137: _omem03_out = reg_1038;
    138: _omem03_out = reg_0187;
    139: _omem03_out = reg_0639;
    140: _omem03_out = reg_1066;
    141: _omem03_out = reg_0704;
    142: _omem03_out = reg_0037;
    143: _omem03_out = reg_0642;
    144: _omem03_out = reg_0098;
    145: _omem03_out = reg_0672;
    146: _omem03_out = reg_1039;
    147: _omem03_out = reg_0283;
    148: _omem03_out = reg_0710;
    149: _omem03_out = reg_0530;
    150: _omem03_out = reg_0607;
    151: _omem03_out = reg_0614;
    152: _omem03_out = reg_0200;
    153: _omem03_out = reg_0336;
    154: _omem03_out = reg_0654;
    155: _omem03_out = reg_1045;
    156: _omem03_out = reg_0277;
    157: _omem03_out = reg_0160;
    158: _omem03_out = reg_0467;
    159: _omem03_out = reg_0587;
    default: _omem03_out = 0;
    endcase
  end // always @ ( * )
  assign omem03_out = _omem03_out[8:0];
  reg [8:0] _omem04_out;
  always @ ( * ) begin
    case ( state )
    117: _omem04_out = reg_0013;
    118: _omem04_out = reg_0959;
    119: _omem04_out = reg_1069;
    120: _omem04_out = reg_0753;
    121: _omem04_out = reg_0567;
    122: _omem04_out = reg_0204;
    123: _omem04_out = reg_0100;
    124: _omem04_out = reg_0013;
    125: _omem04_out = reg_1234;
    126: _omem04_out = reg_0578;
    127: _omem04_out = reg_0282;
    128: _omem04_out = reg_0502;
    129: _omem04_out = reg_0525;
    130: _omem04_out = reg_0605;
    131: _omem04_out = reg_0499;
    132: _omem04_out = reg_0656;
    133: _omem04_out = reg_0370;
    134: _omem04_out = reg_1106;
    135: _omem04_out = reg_0611;
    136: _omem04_out = reg_0933;
    137: _omem04_out = reg_0093;
    138: _omem04_out = reg_0480;
    139: _omem04_out = reg_0683;
    140: _omem04_out = reg_0015;
    141: _omem04_out = reg_0490;
    142: _omem04_out = reg_0204;
    143: _omem04_out = reg_0514;
    144: _omem04_out = reg_0102;
    145: _omem04_out = reg_0997;
    146: _omem04_out = reg_1037;
    147: _omem04_out = reg_0844;
    148: _omem04_out = reg_0842;
    149: _omem04_out = reg_0208;
    150: _omem04_out = reg_0655;
    151: _omem04_out = reg_0671;
    152: _omem04_out = reg_0680;
    153: _omem04_out = reg_0646;
    154: _omem04_out = reg_0578;
    155: _omem04_out = reg_0675;
    156: _omem04_out = reg_0534;
    157: _omem04_out = reg_0357;
    158: _omem04_out = reg_0282;
    159: _omem04_out = reg_0686;
    160: _omem04_out = reg_0590;
    161: _omem04_out = reg_0644;
    162: _omem04_out = reg_0753;
    163: _omem04_out = reg_0567;
    164: _omem04_out = reg_0502;
    165: _omem04_out = reg_0237;
    166: _omem04_out = reg_0677;
    167: _omem04_out = reg_0245;
    168: _omem04_out = reg_0249;
    169: _omem04_out = reg_0121;
    170: _omem04_out = reg_0280;
    171: _omem04_out = reg_0679;
    172: _omem04_out = reg_0100;
    173: _omem04_out = reg_0013;
    174: _omem04_out = reg_0304;
    default: _omem04_out = 0;
    endcase
  end // always @ ( * )
  assign omem04_out = _omem04_out[8:0];

  // OP1#0の0番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in00 = imem00_in[11:8];
    58: op1_00_in00 = imem00_in[11:8];
    79: op1_00_in00 = imem00_in[11:8];
    100: op1_00_in00 = imem00_in[11:8];
    112: op1_00_in00 = imem00_in[11:8];
    15: op1_00_in00 = imem01_in[15:12];
    106: op1_00_in00 = imem01_in[15:12];
    19: op1_00_in00 = imem02_in[15:12];
    102: op1_00_in00 = imem02_in[15:12];
    109: op1_00_in00 = imem02_in[15:12];
    11: op1_00_in00 = imem04_in[15:12];
    33: op1_00_in00 = imem00_in[15:12];
    76: op1_00_in00 = imem00_in[15:12];
    83: op1_00_in00 = imem00_in[15:12];
    110: op1_00_in00 = imem00_in[15:12];
    35: op1_00_in00 = imem01_in[11:8];
    96: op1_00_in00 = imem01_in[11:8];
    120: op1_00_in00 = imem01_in[11:8];
    32: op1_00_in00 = reg_0478;
    26: op1_00_in00 = imem05_in[15:12];
    67: op1_00_in00 = imem05_in[15:12];
    78: op1_00_in00 = imem05_in[15:12];
    103: op1_00_in00 = imem05_in[15:12];
    21: op1_00_in00 = imem07_in[11:8];
    24: op1_00_in00 = imem07_in[11:8];
    4: op1_00_in00 = imem07_in[11:8];
    127: op1_00_in00 = imem07_in[11:8];
    41: op1_00_in00 = imem00_in[7:4];
    60: op1_00_in00 = imem00_in[7:4];
    81: op1_00_in00 = imem00_in[7:4];
    91: op1_00_in00 = imem00_in[7:4];
    116: op1_00_in00 = imem00_in[7:4];
    38: op1_00_in00 = reg_0400;
    39: op1_00_in00 = imem04_in[3:0];
    95: op1_00_in00 = imem04_in[3:0];
    113: op1_00_in00 = imem04_in[3:0];
    129: op1_00_in00 = imem04_in[3:0];
    45: op1_00_in00 = imem06_in[11:8];
    117: op1_00_in00 = imem06_in[11:8];
    130: op1_00_in00 = imem06_in[11:8];
    52: op1_00_in00 = imem00_in[3:0];
    94: op1_00_in00 = imem00_in[3:0];
    128: op1_00_in00 = imem00_in[3:0];
    49: op1_00_in00 = reg_0823;
    46: op1_00_in00 = imem06_in[15:12];
    63: op1_00_in00 = imem06_in[15:12];
    54: op1_00_in00 = reg_0875;
    48: op1_00_in00 = reg_0526;
    53: op1_00_in00 = reg_0283;
    61: op1_00_in00 = imem03_in[3:0];
    68: op1_00_in00 = imem03_in[3:0];
    90: op1_00_in00 = imem03_in[3:0];
    93: op1_00_in00 = imem03_in[3:0];
    121: op1_00_in00 = imem03_in[3:0];
    123: op1_00_in00 = imem03_in[3:0];
    71: op1_00_in00 = imem04_in[7:4];
    108: op1_00_in00 = imem04_in[7:4];
    72: op1_00_in00 = imem05_in[3:0];
    92: op1_00_in00 = imem05_in[3:0];
    40: op1_00_in00 = reg_0704;
    55: op1_00_in00 = imem02_in[11:8];
    107: op1_00_in00 = imem02_in[11:8];
    74: op1_00_in00 = reg_0896;
    87: op1_00_in00 = imem03_in[7:4];
    111: op1_00_in00 = imem03_in[7:4];
    73: op1_00_in00 = reg_0905;
    59: op1_00_in00 = reg_0580;
    50: op1_00_in00 = reg_0282;
    86: op1_00_in00 = reg_0121;
    69: op1_00_in00 = reg_0079;
    36: op1_00_in00 = reg_0365;
    42: op1_00_in00 = reg_0365;
    37: op1_00_in00 = reg_0286;
    44: op1_00_in00 = reg_0603;
    22: op1_00_in00 = reg_0114;
    88: op1_00_in00 = imem01_in[3:0];
    105: op1_00_in00 = imem01_in[3:0];
    114: op1_00_in00 = imem01_in[3:0];
    47: op1_00_in00 = reg_0522;
    28: op1_00_in00 = reg_0028;
    56: op1_00_in00 = reg_0330;
    75: op1_00_in00 = reg_0874;
    25: op1_00_in00 = reg_0284;
    34: op1_00_in00 = reg_0245;
    70: op1_00_in00 = reg_0363;
    57: op1_00_in00 = reg_0842;
    77: op1_00_in00 = reg_0396;
    51: op1_00_in00 = reg_0866;
    43: op1_00_in00 = reg_0798;
    62: op1_00_in00 = reg_0555;
    80: op1_00_in00 = reg_0381;
    2: op1_00_in00 = imem07_in[3:0];
    118: op1_00_in00 = imem07_in[3:0];
    125: op1_00_in00 = imem07_in[3:0];
    27: op1_00_in00 = imem07_in[15:12];
    89: op1_00_in00 = imem03_in[11:8];
    82: op1_00_in00 = reg_1449;
    64: op1_00_in00 = reg_0401;
    84: op1_00_in00 = reg_1484;
    65: op1_00_in00 = reg_0554;
    85: op1_00_in00 = reg_0434;
    66: op1_00_in00 = reg_0540;
    97: op1_00_in00 = imem01_in[7:4];
    124: op1_00_in00 = imem01_in[7:4];
    98: op1_00_in00 = imem06_in[7:4];
    99: op1_00_in00 = imem05_in[11:8];
    122: op1_00_in00 = imem05_in[11:8];
    101: op1_00_in00 = imem06_in[3:0];
    104: op1_00_in00 = imem07_in[7:4];
    119: op1_00_in00 = imem07_in[7:4];
    5: op1_00_in00 = reg_0004;
    29: op1_00_in00 = reg_0321;
    115: op1_00_in00 = imem05_in[7:4];
    126: op1_00_in00 = imem02_in[3:0];
    131: op1_00_in00 = imem04_in[11:8];
    default: op1_00_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv00 = 1;
    15: op1_00_inv00 = 1;
    19: op1_00_inv00 = 1;
    11: op1_00_inv00 = 1;
    33: op1_00_inv00 = 1;
    35: op1_00_inv00 = 1;
    21: op1_00_inv00 = 1;
    41: op1_00_inv00 = 1;
    39: op1_00_inv00 = 1;
    52: op1_00_inv00 = 1;
    46: op1_00_inv00 = 1;
    58: op1_00_inv00 = 1;
    48: op1_00_inv00 = 1;
    60: op1_00_inv00 = 1;
    61: op1_00_inv00 = 1;
    76: op1_00_inv00 = 1;
    71: op1_00_inv00 = 1;
    40: op1_00_inv00 = 1;
    55: op1_00_inv00 = 1;
    68: op1_00_inv00 = 1;
    74: op1_00_inv00 = 1;
    87: op1_00_inv00 = 1;
    73: op1_00_inv00 = 1;
    88: op1_00_inv00 = 1;
    56: op1_00_inv00 = 1;
    25: op1_00_inv00 = 1;
    42: op1_00_inv00 = 1;
    4: op1_00_inv00 = 1;
    34: op1_00_inv00 = 1;
    77: op1_00_inv00 = 1;
    51: op1_00_inv00 = 1;
    62: op1_00_inv00 = 1;
    2: op1_00_inv00 = 1;
    27: op1_00_inv00 = 1;
    81: op1_00_inv00 = 1;
    63: op1_00_inv00 = 1;
    83: op1_00_inv00 = 1;
    65: op1_00_inv00 = 1;
    66: op1_00_inv00 = 1;
    91: op1_00_inv00 = 1;
    94: op1_00_inv00 = 1;
    96: op1_00_inv00 = 1;
    97: op1_00_inv00 = 1;
    98: op1_00_inv00 = 1;
    100: op1_00_inv00 = 1;
    101: op1_00_inv00 = 1;
    102: op1_00_inv00 = 1;
    106: op1_00_inv00 = 1;
    107: op1_00_inv00 = 1;
    108: op1_00_inv00 = 1;
    111: op1_00_inv00 = 1;
    112: op1_00_inv00 = 1;
    29: op1_00_inv00 = 1;
    115: op1_00_inv00 = 1;
    117: op1_00_inv00 = 1;
    122: op1_00_inv00 = 1;
    125: op1_00_inv00 = 1;
    126: op1_00_inv00 = 1;
    129: op1_00_inv00 = 1;
    130: op1_00_inv00 = 1;
    131: op1_00_inv00 = 1;
    default: op1_00_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の1番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in01 = reg_0306;
    15: op1_00_in01 = reg_0238;
    19: op1_00_in01 = reg_0133;
    45: op1_00_in01 = reg_0133;
    11: op1_00_in01 = reg_0164;
    33: op1_00_in01 = reg_0581;
    35: op1_00_in01 = reg_0662;
    32: op1_00_in01 = reg_0444;
    26: op1_00_in01 = reg_0395;
    21: op1_00_in01 = reg_0321;
    41: op1_00_in01 = reg_0820;
    38: op1_00_in01 = reg_0363;
    39: op1_00_in01 = reg_0598;
    24: op1_00_in01 = reg_0028;
    52: op1_00_in01 = reg_1099;
    59: op1_00_in01 = reg_1099;
    110: op1_00_in01 = reg_1099;
    49: op1_00_in01 = imem04_in[3:0];
    46: op1_00_in01 = reg_0141;
    51: op1_00_in01 = reg_0141;
    58: op1_00_in01 = reg_1241;
    54: op1_00_in01 = reg_0043;
    48: op1_00_in01 = reg_0528;
    60: op1_00_in01 = reg_1277;
    53: op1_00_in01 = reg_0012;
    61: op1_00_in01 = imem03_in[7:4];
    121: op1_00_in01 = imem03_in[7:4];
    123: op1_00_in01 = imem03_in[7:4];
    67: op1_00_in01 = reg_0873;
    76: op1_00_in01 = reg_0791;
    71: op1_00_in01 = reg_0061;
    72: op1_00_in01 = reg_0317;
    40: op1_00_in01 = reg_0187;
    55: op1_00_in01 = reg_0433;
    68: op1_00_in01 = imem03_in[11:8];
    93: op1_00_in01 = imem03_in[11:8];
    74: op1_00_in01 = imem02_in[3:0];
    87: op1_00_in01 = imem03_in[15:12];
    78: op1_00_in01 = reg_0939;
    73: op1_00_in01 = reg_0827;
    50: op1_00_in01 = reg_0011;
    86: op1_00_in01 = reg_0154;
    69: op1_00_in01 = reg_0290;
    36: op1_00_in01 = reg_0320;
    37: op1_00_in01 = reg_0437;
    44: op1_00_in01 = reg_0538;
    22: op1_00_in01 = reg_0029;
    88: op1_00_in01 = reg_0400;
    85: op1_00_in01 = reg_0400;
    47: op1_00_in01 = reg_0171;
    28: op1_00_in01 = reg_0361;
    56: op1_00_in01 = reg_0247;
    75: op1_00_in01 = reg_0079;
    25: op1_00_in01 = reg_0124;
    42: op1_00_in01 = reg_0047;
    34: op1_00_in01 = reg_0465;
    70: op1_00_in01 = reg_0091;
    57: op1_00_in01 = reg_0843;
    77: op1_00_in01 = reg_0414;
    79: op1_00_in01 = reg_0983;
    43: op1_00_in01 = reg_0370;
    62: op1_00_in01 = reg_0748;
    80: op1_00_in01 = reg_0632;
    2: op1_00_in01 = imem07_in[7:4];
    27: op1_00_in01 = reg_0287;
    81: op1_00_in01 = reg_0907;
    112: op1_00_in01 = reg_0907;
    89: op1_00_in01 = reg_0145;
    63: op1_00_in01 = reg_0720;
    82: op1_00_in01 = reg_0049;
    83: op1_00_in01 = reg_1510;
    64: op1_00_in01 = reg_0384;
    84: op1_00_in01 = reg_0601;
    65: op1_00_in01 = reg_0580;
    90: op1_00_in01 = reg_0288;
    66: op1_00_in01 = reg_0477;
    91: op1_00_in01 = reg_1244;
    92: op1_00_in01 = imem05_in[15:12];
    94: op1_00_in01 = reg_1141;
    95: op1_00_in01 = reg_0835;
    96: op1_00_in01 = reg_0360;
    97: op1_00_in01 = reg_0042;
    98: op1_00_in01 = reg_0215;
    99: op1_00_in01 = reg_0750;
    100: op1_00_in01 = reg_1487;
    101: op1_00_in01 = reg_0115;
    102: op1_00_in01 = reg_0390;
    103: op1_00_in01 = reg_0302;
    104: op1_00_in01 = reg_0893;
    105: op1_00_in01 = imem01_in[7:4];
    106: op1_00_in01 = reg_1068;
    107: op1_00_in01 = reg_0279;
    108: op1_00_in01 = imem04_in[11:8];
    129: op1_00_in01 = imem04_in[11:8];
    109: op1_00_in01 = reg_0495;
    5: op1_00_in01 = imem07_in[3:0];
    111: op1_00_in01 = reg_1093;
    113: op1_00_in01 = reg_1369;
    29: op1_00_in01 = reg_0219;
    114: op1_00_in01 = reg_0895;
    115: op1_00_in01 = imem06_in[3:0];
    116: op1_00_in01 = imem00_in[11:8];
    128: op1_00_in01 = imem00_in[11:8];
    117: op1_00_in01 = reg_1030;
    118: op1_00_in01 = reg_0052;
    119: op1_00_in01 = reg_0520;
    120: op1_00_in01 = reg_0383;
    122: op1_00_in01 = reg_1181;
    124: op1_00_in01 = reg_0362;
    125: op1_00_in01 = imem07_in[15:12];
    127: op1_00_in01 = imem07_in[15:12];
    126: op1_00_in01 = reg_0455;
    130: op1_00_in01 = reg_1209;
    131: op1_00_in01 = imem05_in[3:0];
    default: op1_00_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_00_inv01 = 1;
    11: op1_00_inv01 = 1;
    33: op1_00_inv01 = 1;
    35: op1_00_inv01 = 1;
    32: op1_00_inv01 = 1;
    21: op1_00_inv01 = 1;
    41: op1_00_inv01 = 1;
    38: op1_00_inv01 = 1;
    39: op1_00_inv01 = 1;
    52: op1_00_inv01 = 1;
    54: op1_00_inv01 = 1;
    60: op1_00_inv01 = 1;
    53: op1_00_inv01 = 1;
    67: op1_00_inv01 = 1;
    71: op1_00_inv01 = 1;
    55: op1_00_inv01 = 1;
    73: op1_00_inv01 = 1;
    50: op1_00_inv01 = 1;
    69: op1_00_inv01 = 1;
    44: op1_00_inv01 = 1;
    22: op1_00_inv01 = 1;
    88: op1_00_inv01 = 1;
    47: op1_00_inv01 = 1;
    75: op1_00_inv01 = 1;
    42: op1_00_inv01 = 1;
    70: op1_00_inv01 = 1;
    79: op1_00_inv01 = 1;
    2: op1_00_inv01 = 1;
    89: op1_00_inv01 = 1;
    63: op1_00_inv01 = 1;
    82: op1_00_inv01 = 1;
    83: op1_00_inv01 = 1;
    64: op1_00_inv01 = 1;
    90: op1_00_inv01 = 1;
    85: op1_00_inv01 = 1;
    91: op1_00_inv01 = 1;
    93: op1_00_inv01 = 1;
    94: op1_00_inv01 = 1;
    95: op1_00_inv01 = 1;
    98: op1_00_inv01 = 1;
    101: op1_00_inv01 = 1;
    102: op1_00_inv01 = 1;
    103: op1_00_inv01 = 1;
    105: op1_00_inv01 = 1;
    107: op1_00_inv01 = 1;
    109: op1_00_inv01 = 1;
    110: op1_00_inv01 = 1;
    112: op1_00_inv01 = 1;
    113: op1_00_inv01 = 1;
    29: op1_00_inv01 = 1;
    114: op1_00_inv01 = 1;
    115: op1_00_inv01 = 1;
    117: op1_00_inv01 = 1;
    118: op1_00_inv01 = 1;
    120: op1_00_inv01 = 1;
    121: op1_00_inv01 = 1;
    123: op1_00_inv01 = 1;
    125: op1_00_inv01 = 1;
    126: op1_00_inv01 = 1;
    130: op1_00_inv01 = 1;
    131: op1_00_inv01 = 1;
    default: op1_00_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の2番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in02 = reg_0293;
    15: op1_00_in02 = reg_0165;
    19: op1_00_in02 = imem03_in[7:4];
    11: op1_00_in02 = reg_0150;
    33: op1_00_in02 = reg_0554;
    35: op1_00_in02 = imem02_in[3:0];
    32: op1_00_in02 = reg_0426;
    26: op1_00_in02 = reg_0391;
    21: op1_00_in02 = reg_0324;
    41: op1_00_in02 = reg_0803;
    38: op1_00_in02 = reg_0041;
    39: op1_00_in02 = reg_0596;
    71: op1_00_in02 = reg_0596;
    45: op1_00_in02 = reg_0160;
    24: op1_00_in02 = reg_0186;
    52: op1_00_in02 = reg_1078;
    65: op1_00_in02 = reg_1078;
    49: op1_00_in02 = reg_0594;
    46: op1_00_in02 = reg_0397;
    51: op1_00_in02 = reg_0397;
    58: op1_00_in02 = reg_1227;
    54: op1_00_in02 = reg_0679;
    48: op1_00_in02 = reg_0458;
    60: op1_00_in02 = reg_1242;
    53: op1_00_in02 = reg_0011;
    61: op1_00_in02 = imem03_in[15:12];
    68: op1_00_in02 = imem03_in[15:12];
    123: op1_00_in02 = imem03_in[15:12];
    67: op1_00_in02 = reg_0492;
    76: op1_00_in02 = reg_1510;
    72: op1_00_in02 = reg_0038;
    40: op1_00_in02 = reg_0298;
    55: op1_00_in02 = reg_0971;
    74: op1_00_in02 = imem02_in[11:8];
    87: op1_00_in02 = reg_0218;
    78: op1_00_in02 = reg_0183;
    73: op1_00_in02 = imem06_in[15:12];
    59: op1_00_in02 = imem00_in[15:12];
    116: op1_00_in02 = imem00_in[15:12];
    50: op1_00_in02 = reg_0667;
    86: op1_00_in02 = reg_0573;
    69: op1_00_in02 = reg_0222;
    36: op1_00_in02 = reg_0091;
    37: op1_00_in02 = imem07_in[15:12];
    25: op1_00_in02 = imem07_in[15:12];
    44: op1_00_in02 = reg_0539;
    22: op1_00_in02 = reg_0030;
    88: op1_00_in02 = reg_0335;
    47: op1_00_in02 = reg_0308;
    28: op1_00_in02 = reg_0051;
    56: op1_00_in02 = reg_0698;
    75: op1_00_in02 = reg_0012;
    42: op1_00_in02 = imem01_in[7:4];
    34: op1_00_in02 = imem07_in[7:4];
    70: op1_00_in02 = reg_0724;
    57: op1_00_in02 = reg_1052;
    77: op1_00_in02 = reg_0969;
    79: op1_00_in02 = reg_0907;
    43: op1_00_in02 = imem04_in[7:4];
    62: op1_00_in02 = reg_1278;
    80: op1_00_in02 = reg_0006;
    27: op1_00_in02 = reg_0408;
    81: op1_00_in02 = reg_1487;
    89: op1_00_in02 = reg_0143;
    63: op1_00_in02 = reg_0133;
    82: op1_00_in02 = reg_1063;
    83: op1_00_in02 = reg_0616;
    64: op1_00_in02 = reg_0092;
    96: op1_00_in02 = reg_0092;
    84: op1_00_in02 = reg_0196;
    90: op1_00_in02 = reg_0790;
    85: op1_00_in02 = reg_0363;
    124: op1_00_in02 = reg_0363;
    66: op1_00_in02 = imem05_in[7:4];
    91: op1_00_in02 = reg_1241;
    92: op1_00_in02 = reg_0648;
    93: op1_00_in02 = reg_0314;
    94: op1_00_in02 = reg_1243;
    95: op1_00_in02 = reg_0337;
    97: op1_00_in02 = imem02_in[15:12];
    98: op1_00_in02 = reg_0213;
    99: op1_00_in02 = reg_0266;
    100: op1_00_in02 = reg_0804;
    101: op1_00_in02 = reg_0717;
    102: op1_00_in02 = reg_0497;
    103: op1_00_in02 = reg_0090;
    104: op1_00_in02 = reg_0498;
    105: op1_00_in02 = reg_0662;
    106: op1_00_in02 = reg_0447;
    107: op1_00_in02 = imem03_in[3:0];
    108: op1_00_in02 = reg_1503;
    109: op1_00_in02 = reg_1207;
    110: op1_00_in02 = reg_0501;
    111: op1_00_in02 = reg_1199;
    121: op1_00_in02 = reg_1199;
    112: op1_00_in02 = reg_0613;
    113: op1_00_in02 = reg_0264;
    29: op1_00_in02 = reg_0004;
    114: op1_00_in02 = imem02_in[7:4];
    115: op1_00_in02 = reg_0316;
    117: op1_00_in02 = reg_1058;
    118: op1_00_in02 = reg_0053;
    119: op1_00_in02 = reg_0483;
    120: op1_00_in02 = reg_0899;
    122: op1_00_in02 = reg_0697;
    125: op1_00_in02 = reg_0299;
    126: op1_00_in02 = reg_0822;
    127: op1_00_in02 = reg_1182;
    128: op1_00_in02 = reg_1079;
    129: op1_00_in02 = reg_0536;
    130: op1_00_in02 = reg_0782;
    131: op1_00_in02 = reg_0833;
    default: op1_00_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv02 = 1;
    19: op1_00_inv02 = 1;
    35: op1_00_inv02 = 1;
    21: op1_00_inv02 = 1;
    45: op1_00_inv02 = 1;
    49: op1_00_inv02 = 1;
    46: op1_00_inv02 = 1;
    58: op1_00_inv02 = 1;
    48: op1_00_inv02 = 1;
    60: op1_00_inv02 = 1;
    76: op1_00_inv02 = 1;
    40: op1_00_inv02 = 1;
    55: op1_00_inv02 = 1;
    68: op1_00_inv02 = 1;
    87: op1_00_inv02 = 1;
    73: op1_00_inv02 = 1;
    50: op1_00_inv02 = 1;
    69: op1_00_inv02 = 1;
    36: op1_00_inv02 = 1;
    22: op1_00_inv02 = 1;
    88: op1_00_inv02 = 1;
    47: op1_00_inv02 = 1;
    28: op1_00_inv02 = 1;
    56: op1_00_inv02 = 1;
    75: op1_00_inv02 = 1;
    25: op1_00_inv02 = 1;
    42: op1_00_inv02 = 1;
    70: op1_00_inv02 = 1;
    77: op1_00_inv02 = 1;
    51: op1_00_inv02 = 1;
    43: op1_00_inv02 = 1;
    62: op1_00_inv02 = 1;
    89: op1_00_inv02 = 1;
    83: op1_00_inv02 = 1;
    64: op1_00_inv02 = 1;
    90: op1_00_inv02 = 1;
    91: op1_00_inv02 = 1;
    92: op1_00_inv02 = 1;
    93: op1_00_inv02 = 1;
    95: op1_00_inv02 = 1;
    101: op1_00_inv02 = 1;
    105: op1_00_inv02 = 1;
    106: op1_00_inv02 = 1;
    109: op1_00_inv02 = 1;
    110: op1_00_inv02 = 1;
    112: op1_00_inv02 = 1;
    115: op1_00_inv02 = 1;
    117: op1_00_inv02 = 1;
    119: op1_00_inv02 = 1;
    120: op1_00_inv02 = 1;
    125: op1_00_inv02 = 1;
    126: op1_00_inv02 = 1;
    127: op1_00_inv02 = 1;
    128: op1_00_inv02 = 1;
    129: op1_00_inv02 = 1;
    130: op1_00_inv02 = 1;
    131: op1_00_inv02 = 1;
    default: op1_00_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の3番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in03 = reg_0153;
    15: op1_00_in03 = reg_0196;
    19: op1_00_in03 = reg_0290;
    11: op1_00_in03 = reg_0129;
    33: op1_00_in03 = reg_0186;
    35: op1_00_in03 = imem02_in[7:4];
    54: op1_00_in03 = imem02_in[7:4];
    32: op1_00_in03 = reg_0427;
    26: op1_00_in03 = reg_0367;
    21: op1_00_in03 = reg_0170;
    41: op1_00_in03 = reg_0248;
    38: op1_00_in03 = imem02_in[15:12];
    114: op1_00_in03 = imem02_in[15:12];
    39: op1_00_in03 = reg_0340;
    45: op1_00_in03 = reg_0905;
    24: op1_00_in03 = reg_0002;
    52: op1_00_in03 = reg_0250;
    59: op1_00_in03 = reg_0250;
    57: op1_00_in03 = reg_0250;
    49: op1_00_in03 = reg_0574;
    46: op1_00_in03 = reg_0859;
    58: op1_00_in03 = reg_0249;
    48: op1_00_in03 = reg_0459;
    60: op1_00_in03 = reg_0804;
    53: op1_00_in03 = reg_0975;
    61: op1_00_in03 = reg_1301;
    67: op1_00_in03 = reg_0393;
    76: op1_00_in03 = reg_0613;
    71: op1_00_in03 = reg_0470;
    108: op1_00_in03 = reg_0470;
    72: op1_00_in03 = imem06_in[3:0];
    40: op1_00_in03 = imem07_in[11:8];
    55: op1_00_in03 = reg_0934;
    68: op1_00_in03 = reg_0411;
    74: op1_00_in03 = reg_0457;
    87: op1_00_in03 = reg_1325;
    78: op1_00_in03 = reg_1514;
    73: op1_00_in03 = reg_0637;
    50: op1_00_in03 = reg_0553;
    86: op1_00_in03 = reg_0706;
    69: op1_00_in03 = reg_0612;
    36: op1_00_in03 = reg_0092;
    85: op1_00_in03 = reg_0092;
    37: op1_00_in03 = reg_0618;
    44: op1_00_in03 = reg_0896;
    22: op1_00_in03 = imem07_in[7:4];
    98: op1_00_in03 = imem07_in[7:4];
    88: op1_00_in03 = reg_0078;
    120: op1_00_in03 = reg_0078;
    47: op1_00_in03 = reg_0289;
    28: op1_00_in03 = reg_0052;
    56: op1_00_in03 = reg_0535;
    75: op1_00_in03 = reg_0679;
    25: op1_00_in03 = reg_0029;
    42: op1_00_in03 = reg_0010;
    70: op1_00_in03 = reg_0010;
    34: op1_00_in03 = reg_0437;
    77: op1_00_in03 = reg_0599;
    51: op1_00_in03 = reg_0398;
    79: op1_00_in03 = reg_1278;
    116: op1_00_in03 = reg_1278;
    43: op1_00_in03 = reg_0488;
    62: op1_00_in03 = reg_1277;
    80: op1_00_in03 = reg_0069;
    27: op1_00_in03 = reg_0415;
    81: op1_00_in03 = reg_1470;
    89: op1_00_in03 = reg_0000;
    63: op1_00_in03 = reg_0109;
    82: op1_00_in03 = reg_0823;
    83: op1_00_in03 = reg_1079;
    64: op1_00_in03 = reg_0899;
    84: op1_00_in03 = reg_0631;
    65: op1_00_in03 = reg_0523;
    90: op1_00_in03 = reg_1280;
    66: op1_00_in03 = reg_0303;
    91: op1_00_in03 = reg_0791;
    92: op1_00_in03 = reg_0562;
    93: op1_00_in03 = reg_0558;
    94: op1_00_in03 = reg_1281;
    95: op1_00_in03 = reg_1189;
    96: op1_00_in03 = reg_0400;
    124: op1_00_in03 = reg_0400;
    97: op1_00_in03 = reg_0499;
    99: op1_00_in03 = reg_0333;
    100: op1_00_in03 = reg_0803;
    101: op1_00_in03 = reg_0194;
    102: op1_00_in03 = reg_0054;
    103: op1_00_in03 = reg_0872;
    104: op1_00_in03 = reg_1415;
    105: op1_00_in03 = imem02_in[11:8];
    106: op1_00_in03 = reg_0662;
    107: op1_00_in03 = imem03_in[11:8];
    109: op1_00_in03 = reg_0307;
    110: op1_00_in03 = reg_1490;
    111: op1_00_in03 = reg_0178;
    112: op1_00_in03 = reg_0486;
    113: op1_00_in03 = reg_0034;
    29: op1_00_in03 = reg_0087;
    115: op1_00_in03 = reg_1508;
    117: op1_00_in03 = reg_0784;
    118: op1_00_in03 = reg_1182;
    119: op1_00_in03 = reg_0123;
    121: op1_00_in03 = reg_0107;
    122: op1_00_in03 = reg_0477;
    123: op1_00_in03 = reg_0291;
    125: op1_00_in03 = reg_0156;
    126: op1_00_in03 = reg_0533;
    128: op1_00_in03 = reg_0958;
    129: op1_00_in03 = reg_0019;
    130: op1_00_in03 = reg_0752;
    131: op1_00_in03 = reg_0466;
    default: op1_00_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    11: op1_00_inv03 = 1;
    33: op1_00_inv03 = 1;
    32: op1_00_inv03 = 1;
    26: op1_00_inv03 = 1;
    39: op1_00_inv03 = 1;
    45: op1_00_inv03 = 1;
    24: op1_00_inv03 = 1;
    52: op1_00_inv03 = 1;
    49: op1_00_inv03 = 1;
    54: op1_00_inv03 = 1;
    60: op1_00_inv03 = 1;
    67: op1_00_inv03 = 1;
    76: op1_00_inv03 = 1;
    74: op1_00_inv03 = 1;
    87: op1_00_inv03 = 1;
    86: op1_00_inv03 = 1;
    37: op1_00_inv03 = 1;
    88: op1_00_inv03 = 1;
    47: op1_00_inv03 = 1;
    75: op1_00_inv03 = 1;
    25: op1_00_inv03 = 1;
    34: op1_00_inv03 = 1;
    57: op1_00_inv03 = 1;
    62: op1_00_inv03 = 1;
    27: op1_00_inv03 = 1;
    81: op1_00_inv03 = 1;
    89: op1_00_inv03 = 1;
    63: op1_00_inv03 = 1;
    64: op1_00_inv03 = 1;
    84: op1_00_inv03 = 1;
    65: op1_00_inv03 = 1;
    85: op1_00_inv03 = 1;
    66: op1_00_inv03 = 1;
    94: op1_00_inv03 = 1;
    96: op1_00_inv03 = 1;
    100: op1_00_inv03 = 1;
    101: op1_00_inv03 = 1;
    102: op1_00_inv03 = 1;
    103: op1_00_inv03 = 1;
    107: op1_00_inv03 = 1;
    111: op1_00_inv03 = 1;
    112: op1_00_inv03 = 1;
    113: op1_00_inv03 = 1;
    114: op1_00_inv03 = 1;
    115: op1_00_inv03 = 1;
    116: op1_00_inv03 = 1;
    119: op1_00_inv03 = 1;
    120: op1_00_inv03 = 1;
    121: op1_00_inv03 = 1;
    123: op1_00_inv03 = 1;
    128: op1_00_inv03 = 1;
    129: op1_00_inv03 = 1;
    default: op1_00_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の4番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in04 = reg_0267;
    15: op1_00_in04 = reg_0183;
    19: op1_00_in04 = reg_0291;
    11: op1_00_in04 = reg_0117;
    33: op1_00_in04 = reg_0523;
    60: op1_00_in04 = reg_0523;
    35: op1_00_in04 = reg_0631;
    32: op1_00_in04 = reg_0411;
    26: op1_00_in04 = reg_0347;
    21: op1_00_in04 = reg_0309;
    41: op1_00_in04 = reg_0725;
    38: op1_00_in04 = reg_0154;
    39: op1_00_in04 = reg_0305;
    43: op1_00_in04 = reg_0305;
    45: op1_00_in04 = reg_0866;
    52: op1_00_in04 = reg_0293;
    112: op1_00_in04 = reg_0293;
    49: op1_00_in04 = reg_0978;
    68: op1_00_in04 = reg_0978;
    46: op1_00_in04 = reg_0372;
    58: op1_00_in04 = reg_1201;
    54: op1_00_in04 = reg_0256;
    48: op1_00_in04 = reg_0023;
    53: op1_00_in04 = reg_0455;
    61: op1_00_in04 = reg_0348;
    67: op1_00_in04 = reg_0575;
    76: op1_00_in04 = reg_1490;
    94: op1_00_in04 = reg_1490;
    71: op1_00_in04 = reg_1419;
    72: op1_00_in04 = reg_1064;
    40: op1_00_in04 = reg_0779;
    55: op1_00_in04 = reg_0933;
    74: op1_00_in04 = reg_0608;
    87: op1_00_in04 = imem04_in[11:8];
    78: op1_00_in04 = reg_0303;
    44: op1_00_in04 = reg_0303;
    73: op1_00_in04 = reg_0526;
    59: op1_00_in04 = reg_1027;
    50: op1_00_in04 = imem02_in[3:0];
    86: op1_00_in04 = reg_0177;
    69: op1_00_in04 = reg_0606;
    36: op1_00_in04 = reg_0278;
    37: op1_00_in04 = reg_0620;
    22: op1_00_in04 = reg_0003;
    88: op1_00_in04 = reg_0079;
    96: op1_00_in04 = reg_0079;
    47: op1_00_in04 = reg_0459;
    28: op1_00_in04 = imem07_in[7:4];
    56: op1_00_in04 = reg_0695;
    109: op1_00_in04 = reg_0695;
    75: op1_00_in04 = reg_0332;
    25: op1_00_in04 = reg_0114;
    42: op1_00_in04 = reg_0254;
    34: op1_00_in04 = reg_0618;
    70: op1_00_in04 = reg_0222;
    57: op1_00_in04 = reg_0249;
    77: op1_00_in04 = reg_0094;
    51: op1_00_in04 = reg_0396;
    79: op1_00_in04 = reg_1487;
    62: op1_00_in04 = reg_0842;
    80: op1_00_in04 = reg_1132;
    27: op1_00_in04 = reg_0413;
    81: op1_00_in04 = reg_0961;
    89: op1_00_in04 = reg_0180;
    63: op1_00_in04 = reg_0716;
    82: op1_00_in04 = reg_1517;
    83: op1_00_in04 = reg_0501;
    64: op1_00_in04 = reg_0044;
    84: op1_00_in04 = reg_0039;
    65: op1_00_in04 = reg_0221;
    90: op1_00_in04 = reg_0427;
    85: op1_00_in04 = reg_1103;
    66: op1_00_in04 = reg_0393;
    91: op1_00_in04 = reg_1243;
    92: op1_00_in04 = reg_0131;
    93: op1_00_in04 = reg_1226;
    95: op1_00_in04 = reg_0236;
    97: op1_00_in04 = reg_0169;
    98: op1_00_in04 = imem07_in[15:12];
    99: op1_00_in04 = reg_0701;
    100: op1_00_in04 = reg_0805;
    101: op1_00_in04 = reg_0584;
    102: op1_00_in04 = reg_0776;
    103: op1_00_in04 = reg_0275;
    104: op1_00_in04 = reg_1060;
    105: op1_00_in04 = imem02_in[15:12];
    106: op1_00_in04 = imem02_in[7:4];
    107: op1_00_in04 = reg_0699;
    108: op1_00_in04 = imem05_in[11:8];
    110: op1_00_in04 = reg_0250;
    111: op1_00_in04 = reg_0113;
    121: op1_00_in04 = reg_0113;
    113: op1_00_in04 = reg_0731;
    29: op1_00_in04 = reg_0123;
    114: op1_00_in04 = reg_1344;
    115: op1_00_in04 = reg_0115;
    116: op1_00_in04 = reg_1099;
    117: op1_00_in04 = reg_0161;
    119: op1_00_in04 = reg_1182;
    120: op1_00_in04 = reg_0724;
    122: op1_00_in04 = reg_0937;
    123: op1_00_in04 = reg_1139;
    124: op1_00_in04 = reg_0257;
    125: op1_00_in04 = reg_0158;
    126: op1_00_in04 = reg_0900;
    128: op1_00_in04 = reg_1242;
    129: op1_00_in04 = reg_0210;
    130: op1_00_in04 = reg_0110;
    131: op1_00_in04 = reg_0272;
    default: op1_00_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv04 = 1;
    15: op1_00_inv04 = 1;
    19: op1_00_inv04 = 1;
    35: op1_00_inv04 = 1;
    32: op1_00_inv04 = 1;
    26: op1_00_inv04 = 1;
    41: op1_00_inv04 = 1;
    38: op1_00_inv04 = 1;
    39: op1_00_inv04 = 1;
    52: op1_00_inv04 = 1;
    49: op1_00_inv04 = 1;
    53: op1_00_inv04 = 1;
    61: op1_00_inv04 = 1;
    72: op1_00_inv04 = 1;
    40: op1_00_inv04 = 1;
    74: op1_00_inv04 = 1;
    50: op1_00_inv04 = 1;
    86: op1_00_inv04 = 1;
    37: op1_00_inv04 = 1;
    44: op1_00_inv04 = 1;
    22: op1_00_inv04 = 1;
    88: op1_00_inv04 = 1;
    47: op1_00_inv04 = 1;
    28: op1_00_inv04 = 1;
    56: op1_00_inv04 = 1;
    25: op1_00_inv04 = 1;
    42: op1_00_inv04 = 1;
    51: op1_00_inv04 = 1;
    79: op1_00_inv04 = 1;
    43: op1_00_inv04 = 1;
    62: op1_00_inv04 = 1;
    80: op1_00_inv04 = 1;
    64: op1_00_inv04 = 1;
    66: op1_00_inv04 = 1;
    92: op1_00_inv04 = 1;
    94: op1_00_inv04 = 1;
    98: op1_00_inv04 = 1;
    99: op1_00_inv04 = 1;
    100: op1_00_inv04 = 1;
    102: op1_00_inv04 = 1;
    103: op1_00_inv04 = 1;
    107: op1_00_inv04 = 1;
    109: op1_00_inv04 = 1;
    110: op1_00_inv04 = 1;
    111: op1_00_inv04 = 1;
    112: op1_00_inv04 = 1;
    113: op1_00_inv04 = 1;
    114: op1_00_inv04 = 1;
    117: op1_00_inv04 = 1;
    120: op1_00_inv04 = 1;
    121: op1_00_inv04 = 1;
    124: op1_00_inv04 = 1;
    125: op1_00_inv04 = 1;
    128: op1_00_inv04 = 1;
    131: op1_00_inv04 = 1;
    default: op1_00_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の5番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in05 = reg_0248;
    15: op1_00_in05 = reg_0166;
    19: op1_00_in05 = reg_0198;
    11: op1_00_in05 = reg_0094;
    33: op1_00_in05 = reg_0485;
    35: op1_00_in05 = reg_0605;
    69: op1_00_in05 = reg_0605;
    32: op1_00_in05 = imem04_in[11:8];
    26: op1_00_in05 = reg_0345;
    21: op1_00_in05 = reg_0298;
    41: op1_00_in05 = reg_0722;
    38: op1_00_in05 = reg_0705;
    39: op1_00_in05 = reg_0319;
    43: op1_00_in05 = reg_0319;
    45: op1_00_in05 = reg_0860;
    52: op1_00_in05 = reg_0983;
    49: op1_00_in05 = reg_0969;
    46: op1_00_in05 = reg_0822;
    58: op1_00_in05 = reg_0460;
    54: op1_00_in05 = reg_0432;
    48: op1_00_in05 = reg_0212;
    60: op1_00_in05 = reg_0221;
    53: op1_00_in05 = reg_0588;
    74: op1_00_in05 = reg_0588;
    97: op1_00_in05 = reg_0588;
    61: op1_00_in05 = imem04_in[7:4];
    67: op1_00_in05 = reg_1346;
    76: op1_00_in05 = reg_0552;
    71: op1_00_in05 = reg_0698;
    72: op1_00_in05 = reg_0795;
    40: op1_00_in05 = reg_0663;
    55: op1_00_in05 = reg_0390;
    68: op1_00_in05 = reg_0676;
    87: op1_00_in05 = reg_0088;
    78: op1_00_in05 = reg_1485;
    73: op1_00_in05 = reg_0529;
    59: op1_00_in05 = reg_0172;
    62: op1_00_in05 = reg_0172;
    50: op1_00_in05 = reg_0976;
    86: op1_00_in05 = reg_0557;
    36: op1_00_in05 = reg_0012;
    37: op1_00_in05 = reg_0593;
    44: op1_00_in05 = reg_0300;
    88: op1_00_in05 = reg_0724;
    47: op1_00_in05 = reg_0215;
    56: op1_00_in05 = reg_0574;
    75: op1_00_in05 = reg_1103;
    25: op1_00_in05 = reg_0186;
    42: op1_00_in05 = reg_0631;
    34: op1_00_in05 = reg_0620;
    70: op1_00_in05 = reg_0679;
    57: op1_00_in05 = reg_1141;
    77: op1_00_in05 = reg_0369;
    51: op1_00_in05 = reg_0863;
    79: op1_00_in05 = reg_0803;
    80: op1_00_in05 = reg_0311;
    27: op1_00_in05 = reg_0002;
    81: op1_00_in05 = reg_1418;
    89: op1_00_in05 = reg_0789;
    63: op1_00_in05 = reg_0374;
    82: op1_00_in05 = reg_0957;
    83: op1_00_in05 = reg_0580;
    64: op1_00_in05 = reg_1029;
    84: op1_00_in05 = imem06_in[15:12];
    65: op1_00_in05 = reg_0136;
    90: op1_00_in05 = imem04_in[3:0];
    85: op1_00_in05 = reg_0608;
    66: op1_00_in05 = reg_0243;
    91: op1_00_in05 = reg_1081;
    92: op1_00_in05 = reg_1404;
    93: op1_00_in05 = reg_1208;
    94: op1_00_in05 = reg_0804;
    95: op1_00_in05 = imem05_in[3:0];
    96: op1_00_in05 = reg_0257;
    98: op1_00_in05 = reg_0995;
    99: op1_00_in05 = reg_0564;
    100: op1_00_in05 = reg_0523;
    101: op1_00_in05 = reg_0617;
    102: op1_00_in05 = reg_0970;
    103: op1_00_in05 = reg_0575;
    104: op1_00_in05 = reg_0135;
    105: op1_00_in05 = reg_0423;
    106: op1_00_in05 = imem02_in[15:12];
    107: op1_00_in05 = reg_0732;
    108: op1_00_in05 = reg_0832;
    109: op1_00_in05 = reg_0227;
    110: op1_00_in05 = reg_1028;
    111: op1_00_in05 = reg_0411;
    112: op1_00_in05 = reg_1459;
    113: op1_00_in05 = reg_1083;
    114: op1_00_in05 = reg_0846;
    115: op1_00_in05 = reg_0636;
    116: op1_00_in05 = reg_0501;
    117: op1_00_in05 = reg_0925;
    120: op1_00_in05 = reg_0896;
    121: op1_00_in05 = reg_0448;
    122: op1_00_in05 = reg_0450;
    123: op1_00_in05 = reg_1325;
    124: op1_00_in05 = reg_0634;
    125: op1_00_in05 = reg_0924;
    126: op1_00_in05 = reg_0436;
    128: op1_00_in05 = reg_1278;
    129: op1_00_in05 = imem05_in[11:8];
    130: op1_00_in05 = reg_0716;
    131: op1_00_in05 = reg_0205;
    default: op1_00_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    19: op1_00_inv05 = 1;
    11: op1_00_inv05 = 1;
    26: op1_00_inv05 = 1;
    39: op1_00_inv05 = 1;
    52: op1_00_inv05 = 1;
    49: op1_00_inv05 = 1;
    54: op1_00_inv05 = 1;
    60: op1_00_inv05 = 1;
    67: op1_00_inv05 = 1;
    72: op1_00_inv05 = 1;
    74: op1_00_inv05 = 1;
    73: op1_00_inv05 = 1;
    50: op1_00_inv05 = 1;
    86: op1_00_inv05 = 1;
    69: op1_00_inv05 = 1;
    36: op1_00_inv05 = 1;
    44: op1_00_inv05 = 1;
    88: op1_00_inv05 = 1;
    47: op1_00_inv05 = 1;
    56: op1_00_inv05 = 1;
    75: op1_00_inv05 = 1;
    25: op1_00_inv05 = 1;
    42: op1_00_inv05 = 1;
    70: op1_00_inv05 = 1;
    51: op1_00_inv05 = 1;
    43: op1_00_inv05 = 1;
    62: op1_00_inv05 = 1;
    27: op1_00_inv05 = 1;
    89: op1_00_inv05 = 1;
    65: op1_00_inv05 = 1;
    85: op1_00_inv05 = 1;
    66: op1_00_inv05 = 1;
    94: op1_00_inv05 = 1;
    96: op1_00_inv05 = 1;
    97: op1_00_inv05 = 1;
    99: op1_00_inv05 = 1;
    101: op1_00_inv05 = 1;
    102: op1_00_inv05 = 1;
    103: op1_00_inv05 = 1;
    104: op1_00_inv05 = 1;
    106: op1_00_inv05 = 1;
    107: op1_00_inv05 = 1;
    108: op1_00_inv05 = 1;
    112: op1_00_inv05 = 1;
    113: op1_00_inv05 = 1;
    114: op1_00_inv05 = 1;
    116: op1_00_inv05 = 1;
    117: op1_00_inv05 = 1;
    120: op1_00_inv05 = 1;
    121: op1_00_inv05 = 1;
    124: op1_00_inv05 = 1;
    129: op1_00_inv05 = 1;
    default: op1_00_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の6番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in06 = reg_0229;
    15: op1_00_in06 = reg_0167;
    19: op1_00_in06 = reg_0261;
    11: op1_00_in06 = reg_0065;
    33: op1_00_in06 = reg_0476;
    35: op1_00_in06 = reg_0590;
    32: op1_00_in06 = reg_0552;
    68: op1_00_in06 = reg_0552;
    87: op1_00_in06 = reg_0552;
    26: op1_00_in06 = reg_0136;
    21: op1_00_in06 = reg_0228;
    41: op1_00_in06 = reg_0723;
    38: op1_00_in06 = reg_0007;
    39: op1_00_in06 = reg_0237;
    45: op1_00_in06 = reg_0827;
    52: op1_00_in06 = reg_0959;
    49: op1_00_in06 = reg_0932;
    46: op1_00_in06 = reg_0110;
    58: op1_00_in06 = reg_0135;
    54: op1_00_in06 = reg_0776;
    48: op1_00_in06 = reg_0213;
    60: op1_00_in06 = reg_0249;
    53: op1_00_in06 = reg_0562;
    61: op1_00_in06 = imem04_in[11:8];
    67: op1_00_in06 = reg_0317;
    76: op1_00_in06 = reg_1469;
    79: op1_00_in06 = reg_1469;
    71: op1_00_in06 = reg_0835;
    72: op1_00_in06 = reg_0268;
    40: op1_00_in06 = reg_0664;
    55: op1_00_in06 = reg_0055;
    74: op1_00_in06 = reg_0934;
    78: op1_00_in06 = reg_0196;
    73: op1_00_in06 = reg_1225;
    59: op1_00_in06 = reg_0961;
    50: op1_00_in06 = reg_0588;
    42: op1_00_in06 = reg_0588;
    85: op1_00_in06 = reg_0588;
    86: op1_00_in06 = reg_1001;
    69: op1_00_in06 = reg_0587;
    36: op1_00_in06 = reg_0011;
    37: op1_00_in06 = reg_0102;
    44: op1_00_in06 = reg_0873;
    88: op1_00_in06 = reg_0162;
    47: op1_00_in06 = reg_0921;
    56: op1_00_in06 = reg_0681;
    75: op1_00_in06 = reg_1029;
    25: op1_00_in06 = reg_0053;
    34: op1_00_in06 = reg_0361;
    70: op1_00_in06 = reg_0457;
    57: op1_00_in06 = reg_0887;
    77: op1_00_in06 = reg_0698;
    51: op1_00_in06 = reg_0718;
    43: op1_00_in06 = reg_0719;
    62: op1_00_in06 = reg_0202;
    80: op1_00_in06 = reg_1495;
    27: op1_00_in06 = reg_0004;
    81: op1_00_in06 = reg_0524;
    89: op1_00_in06 = reg_0142;
    63: op1_00_in06 = reg_0584;
    82: op1_00_in06 = reg_0190;
    83: op1_00_in06 = reg_1471;
    64: op1_00_in06 = reg_0608;
    84: op1_00_in06 = reg_1437;
    65: op1_00_in06 = reg_1205;
    90: op1_00_in06 = imem04_in[15:12];
    66: op1_00_in06 = reg_0449;
    91: op1_00_in06 = reg_1278;
    92: op1_00_in06 = reg_0939;
    93: op1_00_in06 = reg_0107;
    94: op1_00_in06 = reg_0580;
    116: op1_00_in06 = reg_0580;
    95: op1_00_in06 = reg_0832;
    96: op1_00_in06 = reg_0043;
    97: op1_00_in06 = reg_1343;
    98: op1_00_in06 = reg_1414;
    99: op1_00_in06 = reg_0334;
    100: op1_00_in06 = reg_1230;
    101: op1_00_in06 = reg_0522;
    102: op1_00_in06 = reg_0971;
    103: op1_00_in06 = reg_0589;
    104: op1_00_in06 = reg_0786;
    105: op1_00_in06 = reg_0056;
    106: op1_00_in06 = reg_0456;
    107: op1_00_in06 = reg_0789;
    108: op1_00_in06 = reg_0251;
    109: op1_00_in06 = imem03_in[11:8];
    110: op1_00_in06 = reg_1459;
    111: op1_00_in06 = imem04_in[3:0];
    112: op1_00_in06 = reg_1229;
    113: op1_00_in06 = reg_1200;
    114: op1_00_in06 = reg_0423;
    115: op1_00_in06 = reg_0398;
    117: op1_00_in06 = reg_0960;
    120: op1_00_in06 = reg_0403;
    121: op1_00_in06 = reg_0350;
    122: op1_00_in06 = reg_0393;
    123: op1_00_in06 = reg_0426;
    124: op1_00_in06 = reg_0662;
    125: op1_00_in06 = reg_0489;
    126: op1_00_in06 = reg_0972;
    128: op1_00_in06 = reg_0748;
    129: op1_00_in06 = reg_0338;
    130: op1_00_in06 = reg_1302;
    131: op1_00_in06 = reg_0992;
    default: op1_00_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_00_inv06 = 1;
    19: op1_00_inv06 = 1;
    33: op1_00_inv06 = 1;
    32: op1_00_inv06 = 1;
    26: op1_00_inv06 = 1;
    21: op1_00_inv06 = 1;
    38: op1_00_inv06 = 1;
    45: op1_00_inv06 = 1;
    52: op1_00_inv06 = 1;
    54: op1_00_inv06 = 1;
    48: op1_00_inv06 = 1;
    53: op1_00_inv06 = 1;
    71: op1_00_inv06 = 1;
    72: op1_00_inv06 = 1;
    55: op1_00_inv06 = 1;
    74: op1_00_inv06 = 1;
    87: op1_00_inv06 = 1;
    73: op1_00_inv06 = 1;
    50: op1_00_inv06 = 1;
    86: op1_00_inv06 = 1;
    36: op1_00_inv06 = 1;
    47: op1_00_inv06 = 1;
    75: op1_00_inv06 = 1;
    25: op1_00_inv06 = 1;
    42: op1_00_inv06 = 1;
    34: op1_00_inv06 = 1;
    77: op1_00_inv06 = 1;
    43: op1_00_inv06 = 1;
    62: op1_00_inv06 = 1;
    80: op1_00_inv06 = 1;
    27: op1_00_inv06 = 1;
    81: op1_00_inv06 = 1;
    63: op1_00_inv06 = 1;
    82: op1_00_inv06 = 1;
    64: op1_00_inv06 = 1;
    65: op1_00_inv06 = 1;
    85: op1_00_inv06 = 1;
    92: op1_00_inv06 = 1;
    93: op1_00_inv06 = 1;
    94: op1_00_inv06 = 1;
    95: op1_00_inv06 = 1;
    98: op1_00_inv06 = 1;
    99: op1_00_inv06 = 1;
    104: op1_00_inv06 = 1;
    105: op1_00_inv06 = 1;
    109: op1_00_inv06 = 1;
    110: op1_00_inv06 = 1;
    111: op1_00_inv06 = 1;
    112: op1_00_inv06 = 1;
    115: op1_00_inv06 = 1;
    116: op1_00_inv06 = 1;
    117: op1_00_inv06 = 1;
    121: op1_00_inv06 = 1;
    122: op1_00_inv06 = 1;
    124: op1_00_inv06 = 1;
    126: op1_00_inv06 = 1;
    128: op1_00_inv06 = 1;
    130: op1_00_inv06 = 1;
    default: op1_00_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の7番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in07 = reg_0219;
    15: op1_00_in07 = reg_0160;
    19: op1_00_in07 = reg_0246;
    11: op1_00_in07 = reg_0063;
    33: op1_00_in07 = reg_0445;
    35: op1_00_in07 = reg_0587;
    32: op1_00_in07 = reg_0534;
    26: op1_00_in07 = reg_0070;
    21: op1_00_in07 = reg_0285;
    41: op1_00_in07 = reg_0485;
    38: op1_00_in07 = reg_0327;
    39: op1_00_in07 = reg_0181;
    45: op1_00_in07 = reg_0716;
    52: op1_00_in07 = reg_0927;
    49: op1_00_in07 = reg_0452;
    46: op1_00_in07 = reg_0670;
    58: op1_00_in07 = reg_1148;
    54: op1_00_in07 = reg_0127;
    48: op1_00_in07 = reg_0015;
    60: op1_00_in07 = reg_0987;
    53: op1_00_in07 = reg_0531;
    61: op1_00_in07 = reg_0232;
    67: op1_00_in07 = reg_0207;
    76: op1_00_in07 = reg_1470;
    71: op1_00_in07 = reg_0237;
    72: op1_00_in07 = reg_0316;
    40: op1_00_in07 = reg_0408;
    55: op1_00_in07 = reg_0900;
    68: op1_00_in07 = reg_0464;
    74: op1_00_in07 = reg_1455;
    87: op1_00_in07 = reg_0488;
    78: op1_00_in07 = reg_0130;
    73: op1_00_in07 = imem07_in[3:0];
    59: op1_00_in07 = reg_0641;
    50: op1_00_in07 = reg_0563;
    69: op1_00_in07 = reg_0563;
    42: op1_00_in07 = reg_0563;
    86: op1_00_in07 = reg_0783;
    36: op1_00_in07 = reg_0486;
    37: op1_00_in07 = reg_0484;
    44: op1_00_in07 = reg_0274;
    88: op1_00_in07 = reg_0120;
    47: op1_00_in07 = reg_0922;
    56: op1_00_in07 = reg_0407;
    75: op1_00_in07 = reg_0606;
    70: op1_00_in07 = reg_0742;
    57: op1_00_in07 = reg_0886;
    77: op1_00_in07 = reg_0368;
    51: op1_00_in07 = reg_0524;
    62: op1_00_in07 = reg_0524;
    79: op1_00_in07 = reg_1459;
    43: op1_00_in07 = reg_0129;
    80: op1_00_in07 = reg_1000;
    27: op1_00_in07 = reg_0003;
    81: op1_00_in07 = reg_0476;
    89: op1_00_in07 = reg_1314;
    63: op1_00_in07 = reg_0622;
    115: op1_00_in07 = reg_0622;
    82: op1_00_in07 = reg_0107;
    83: op1_00_in07 = reg_1469;
    64: op1_00_in07 = reg_1260;
    84: op1_00_in07 = reg_0133;
    65: op1_00_in07 = reg_0440;
    90: op1_00_in07 = reg_0263;
    85: op1_00_in07 = reg_1343;
    66: op1_00_in07 = reg_0206;
    91: op1_00_in07 = reg_0672;
    92: op1_00_in07 = reg_0986;
    93: op1_00_in07 = reg_0113;
    94: op1_00_in07 = reg_0221;
    95: op1_00_in07 = reg_0251;
    96: op1_00_in07 = reg_0041;
    97: op1_00_in07 = reg_0712;
    98: op1_00_in07 = reg_0135;
    99: op1_00_in07 = reg_1070;
    100: op1_00_in07 = reg_1418;
    101: op1_00_in07 = reg_0308;
    102: op1_00_in07 = reg_0972;
    103: op1_00_in07 = reg_0449;
    104: op1_00_in07 = reg_0309;
    105: op1_00_in07 = reg_0055;
    106: op1_00_in07 = reg_0889;
    107: op1_00_in07 = reg_0965;
    108: op1_00_in07 = reg_0045;
    109: op1_00_in07 = imem03_in[15:12];
    110: op1_00_in07 = reg_0961;
    111: op1_00_in07 = reg_0297;
    112: op1_00_in07 = reg_1417;
    113: op1_00_in07 = reg_0500;
    114: op1_00_in07 = reg_0934;
    116: op1_00_in07 = reg_0153;
    117: op1_00_in07 = reg_0718;
    120: op1_00_in07 = reg_0447;
    121: op1_00_in07 = reg_0707;
    122: op1_00_in07 = reg_0240;
    123: op1_00_in07 = imem04_in[3:0];
    124: op1_00_in07 = imem02_in[3:0];
    125: op1_00_in07 = reg_0139;
    126: op1_00_in07 = reg_1458;
    128: op1_00_in07 = reg_0806;
    129: op1_00_in07 = reg_0315;
    130: op1_00_in07 = reg_0373;
    131: op1_00_in07 = reg_0340;
    default: op1_00_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv07 = 1;
    15: op1_00_inv07 = 1;
    11: op1_00_inv07 = 1;
    33: op1_00_inv07 = 1;
    32: op1_00_inv07 = 1;
    21: op1_00_inv07 = 1;
    41: op1_00_inv07 = 1;
    45: op1_00_inv07 = 1;
    52: op1_00_inv07 = 1;
    46: op1_00_inv07 = 1;
    58: op1_00_inv07 = 1;
    61: op1_00_inv07 = 1;
    67: op1_00_inv07 = 1;
    76: op1_00_inv07 = 1;
    71: op1_00_inv07 = 1;
    72: op1_00_inv07 = 1;
    74: op1_00_inv07 = 1;
    73: op1_00_inv07 = 1;
    70: op1_00_inv07 = 1;
    77: op1_00_inv07 = 1;
    79: op1_00_inv07 = 1;
    43: op1_00_inv07 = 1;
    62: op1_00_inv07 = 1;
    80: op1_00_inv07 = 1;
    27: op1_00_inv07 = 1;
    82: op1_00_inv07 = 1;
    84: op1_00_inv07 = 1;
    65: op1_00_inv07 = 1;
    92: op1_00_inv07 = 1;
    93: op1_00_inv07 = 1;
    94: op1_00_inv07 = 1;
    96: op1_00_inv07 = 1;
    98: op1_00_inv07 = 1;
    99: op1_00_inv07 = 1;
    100: op1_00_inv07 = 1;
    101: op1_00_inv07 = 1;
    103: op1_00_inv07 = 1;
    104: op1_00_inv07 = 1;
    105: op1_00_inv07 = 1;
    106: op1_00_inv07 = 1;
    107: op1_00_inv07 = 1;
    109: op1_00_inv07 = 1;
    113: op1_00_inv07 = 1;
    114: op1_00_inv07 = 1;
    115: op1_00_inv07 = 1;
    117: op1_00_inv07 = 1;
    121: op1_00_inv07 = 1;
    122: op1_00_inv07 = 1;
    126: op1_00_inv07 = 1;
    131: op1_00_inv07 = 1;
    default: op1_00_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の8番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in08 = reg_0220;
    89: op1_00_in08 = reg_0220;
    15: op1_00_in08 = reg_0147;
    19: op1_00_in08 = reg_0232;
    11: op1_00_in08 = reg_0061;
    33: op1_00_in08 = reg_0428;
    57: op1_00_in08 = reg_0428;
    35: op1_00_in08 = reg_0560;
    73: op1_00_in08 = reg_0560;
    50: op1_00_in08 = reg_0560;
    32: op1_00_in08 = reg_0488;
    26: op1_00_in08 = reg_0331;
    21: op1_00_in08 = reg_0028;
    41: op1_00_in08 = reg_0249;
    38: op1_00_in08 = reg_0069;
    39: op1_00_in08 = imem05_in[3:0];
    45: op1_00_in08 = reg_0714;
    52: op1_00_in08 = reg_0926;
    49: op1_00_in08 = reg_0470;
    46: op1_00_in08 = reg_0617;
    58: op1_00_in08 = reg_0881;
    54: op1_00_in08 = reg_0111;
    48: op1_00_in08 = imem07_in[11:8];
    60: op1_00_in08 = reg_0459;
    53: op1_00_in08 = imem02_in[15:12];
    61: op1_00_in08 = reg_0397;
    67: op1_00_in08 = imem06_in[3:0];
    76: op1_00_in08 = reg_1454;
    71: op1_00_in08 = reg_0211;
    72: op1_00_in08 = reg_0974;
    40: op1_00_in08 = reg_0415;
    55: op1_00_in08 = reg_0712;
    68: op1_00_in08 = reg_0451;
    56: op1_00_in08 = reg_0451;
    74: op1_00_in08 = reg_1433;
    87: op1_00_in08 = reg_0500;
    78: op1_00_in08 = reg_0864;
    122: op1_00_in08 = reg_0864;
    59: op1_00_in08 = reg_0642;
    86: op1_00_in08 = reg_0707;
    69: op1_00_in08 = reg_0631;
    36: op1_00_in08 = reg_0662;
    120: op1_00_in08 = reg_0662;
    37: op1_00_in08 = reg_0124;
    44: op1_00_in08 = reg_0205;
    88: op1_00_in08 = imem02_in[7:4];
    47: op1_00_in08 = reg_0191;
    75: op1_00_in08 = reg_0254;
    42: op1_00_in08 = reg_0532;
    70: op1_00_in08 = reg_0744;
    77: op1_00_in08 = reg_0719;
    51: op1_00_in08 = reg_0619;
    79: op1_00_in08 = reg_1229;
    43: op1_00_in08 = reg_0033;
    62: op1_00_in08 = reg_0883;
    81: op1_00_in08 = reg_0883;
    80: op1_00_in08 = reg_0840;
    27: op1_00_in08 = reg_0050;
    63: op1_00_in08 = reg_0528;
    82: op1_00_in08 = reg_0880;
    83: op1_00_in08 = reg_1053;
    64: op1_00_in08 = reg_0475;
    84: op1_00_in08 = reg_1509;
    65: op1_00_in08 = reg_1322;
    90: op1_00_in08 = reg_1367;
    85: op1_00_in08 = reg_0256;
    66: op1_00_in08 = reg_0040;
    91: op1_00_in08 = reg_1490;
    92: op1_00_in08 = reg_0303;
    93: op1_00_in08 = reg_0104;
    94: op1_00_in08 = reg_1227;
    95: op1_00_in08 = reg_0992;
    96: op1_00_in08 = reg_0010;
    97: op1_00_in08 = reg_0472;
    98: op1_00_in08 = reg_0225;
    99: op1_00_in08 = reg_0183;
    100: op1_00_in08 = reg_0352;
    101: op1_00_in08 = reg_1202;
    102: op1_00_in08 = reg_0382;
    103: op1_00_in08 = reg_0038;
    104: op1_00_in08 = reg_0665;
    105: op1_00_in08 = reg_1493;
    106: op1_00_in08 = reg_0659;
    107: op1_00_in08 = reg_0964;
    108: op1_00_in08 = reg_1180;
    109: op1_00_in08 = reg_0233;
    110: op1_00_in08 = reg_1432;
    111: op1_00_in08 = reg_1203;
    112: op1_00_in08 = reg_0524;
    113: op1_00_in08 = reg_1082;
    114: op1_00_in08 = reg_0561;
    115: op1_00_in08 = reg_1204;
    116: op1_00_in08 = reg_0554;
    117: op1_00_in08 = reg_0586;
    130: op1_00_in08 = reg_0586;
    121: op1_00_in08 = reg_1282;
    123: op1_00_in08 = reg_1233;
    124: op1_00_in08 = reg_0399;
    125: op1_00_in08 = reg_0284;
    126: op1_00_in08 = reg_0128;
    128: op1_00_in08 = reg_1052;
    129: op1_00_in08 = reg_0538;
    131: op1_00_in08 = reg_0562;
    default: op1_00_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv08 = 1;
    15: op1_00_inv08 = 1;
    33: op1_00_inv08 = 1;
    26: op1_00_inv08 = 1;
    39: op1_00_inv08 = 1;
    52: op1_00_inv08 = 1;
    49: op1_00_inv08 = 1;
    60: op1_00_inv08 = 1;
    53: op1_00_inv08 = 1;
    61: op1_00_inv08 = 1;
    67: op1_00_inv08 = 1;
    72: op1_00_inv08 = 1;
    40: op1_00_inv08 = 1;
    68: op1_00_inv08 = 1;
    74: op1_00_inv08 = 1;
    87: op1_00_inv08 = 1;
    73: op1_00_inv08 = 1;
    69: op1_00_inv08 = 1;
    88: op1_00_inv08 = 1;
    56: op1_00_inv08 = 1;
    42: op1_00_inv08 = 1;
    77: op1_00_inv08 = 1;
    79: op1_00_inv08 = 1;
    62: op1_00_inv08 = 1;
    27: op1_00_inv08 = 1;
    81: op1_00_inv08 = 1;
    89: op1_00_inv08 = 1;
    83: op1_00_inv08 = 1;
    64: op1_00_inv08 = 1;
    65: op1_00_inv08 = 1;
    85: op1_00_inv08 = 1;
    91: op1_00_inv08 = 1;
    92: op1_00_inv08 = 1;
    94: op1_00_inv08 = 1;
    98: op1_00_inv08 = 1;
    104: op1_00_inv08 = 1;
    106: op1_00_inv08 = 1;
    107: op1_00_inv08 = 1;
    108: op1_00_inv08 = 1;
    110: op1_00_inv08 = 1;
    113: op1_00_inv08 = 1;
    116: op1_00_inv08 = 1;
    117: op1_00_inv08 = 1;
    125: op1_00_inv08 = 1;
    129: op1_00_inv08 = 1;
    130: op1_00_inv08 = 1;
    default: op1_00_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の9番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in09 = reg_0221;
    15: op1_00_in09 = reg_0120;
    19: op1_00_in09 = reg_0233;
    11: op1_00_in09 = reg_0033;
    33: op1_00_in09 = reg_0410;
    35: op1_00_in09 = reg_0530;
    32: op1_00_in09 = reg_0493;
    26: op1_00_in09 = reg_0315;
    21: op1_00_in09 = reg_0001;
    41: op1_00_in09 = reg_0267;
    38: op1_00_in09 = reg_0279;
    39: op1_00_in09 = imem05_in[15:12];
    45: op1_00_in09 = reg_0524;
    52: op1_00_in09 = reg_0722;
    49: op1_00_in09 = reg_0596;
    46: op1_00_in09 = reg_0295;
    58: op1_00_in09 = reg_0638;
    54: op1_00_in09 = reg_0112;
    48: op1_00_in09 = imem07_in[15:12];
    60: op1_00_in09 = reg_0492;
    53: op1_00_in09 = reg_0497;
    105: op1_00_in09 = reg_0497;
    61: op1_00_in09 = reg_0252;
    67: op1_00_in09 = reg_1105;
    76: op1_00_in09 = reg_1432;
    71: op1_00_in09 = reg_0210;
    72: op1_00_in09 = reg_0925;
    40: op1_00_in09 = reg_0621;
    55: op1_00_in09 = reg_0708;
    68: op1_00_in09 = reg_0862;
    74: op1_00_in09 = reg_0878;
    87: op1_00_in09 = reg_1147;
    78: op1_00_in09 = imem06_in[3:0];
    73: op1_00_in09 = reg_1440;
    59: op1_00_in09 = reg_0201;
    50: op1_00_in09 = reg_0531;
    86: op1_00_in09 = reg_0541;
    69: op1_00_in09 = reg_0876;
    36: op1_00_in09 = reg_0666;
    44: op1_00_in09 = reg_0204;
    88: op1_00_in09 = reg_0474;
    47: op1_00_in09 = reg_0491;
    56: op1_00_in09 = reg_0320;
    75: op1_00_in09 = reg_0475;
    42: op1_00_in09 = reg_0473;
    70: op1_00_in09 = reg_0997;
    57: op1_00_in09 = reg_0416;
    77: op1_00_in09 = reg_0835;
    51: op1_00_in09 = reg_0586;
    79: op1_00_in09 = reg_0821;
    112: op1_00_in09 = reg_0821;
    43: op1_00_in09 = reg_0833;
    62: op1_00_in09 = reg_0642;
    80: op1_00_in09 = reg_0328;
    81: op1_00_in09 = reg_0431;
    89: op1_00_in09 = reg_0107;
    63: op1_00_in09 = reg_0568;
    82: op1_00_in09 = reg_0505;
    83: op1_00_in09 = reg_1459;
    64: op1_00_in09 = reg_0776;
    84: op1_00_in09 = reg_0397;
    65: op1_00_in09 = reg_0122;
    90: op1_00_in09 = reg_0088;
    85: op1_00_in09 = reg_0390;
    66: op1_00_in09 = reg_1036;
    91: op1_00_in09 = reg_0907;
    92: op1_00_in09 = reg_0873;
    93: op1_00_in09 = reg_0880;
    94: op1_00_in09 = reg_0459;
    95: op1_00_in09 = reg_1180;
    96: op1_00_in09 = imem02_in[3:0];
    120: op1_00_in09 = imem02_in[3:0];
    97: op1_00_in09 = reg_0495;
    98: op1_00_in09 = reg_0170;
    99: op1_00_in09 = reg_0302;
    100: op1_00_in09 = reg_0189;
    101: op1_00_in09 = reg_0067;
    102: op1_00_in09 = reg_0629;
    103: op1_00_in09 = imem06_in[11:8];
    104: op1_00_in09 = reg_0441;
    106: op1_00_in09 = reg_0846;
    107: op1_00_in09 = reg_1208;
    108: op1_00_in09 = reg_0939;
    109: op1_00_in09 = reg_0049;
    110: op1_00_in09 = reg_0155;
    111: op1_00_in09 = reg_1200;
    113: op1_00_in09 = reg_0094;
    114: op1_00_in09 = reg_0975;
    115: op1_00_in09 = reg_0212;
    116: op1_00_in09 = reg_0186;
    117: op1_00_in09 = reg_0529;
    121: op1_00_in09 = reg_0348;
    122: op1_00_in09 = imem06_in[7:4];
    123: op1_00_in09 = reg_0281;
    124: op1_00_in09 = reg_0423;
    125: op1_00_in09 = reg_0437;
    126: op1_00_in09 = reg_1140;
    128: op1_00_in09 = reg_0987;
    129: op1_00_in09 = reg_0136;
    130: op1_00_in09 = reg_0522;
    131: op1_00_in09 = reg_0391;
    default: op1_00_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_00_inv09 = 1;
    19: op1_00_inv09 = 1;
    11: op1_00_inv09 = 1;
    33: op1_00_inv09 = 1;
    32: op1_00_inv09 = 1;
    41: op1_00_inv09 = 1;
    38: op1_00_inv09 = 1;
    39: op1_00_inv09 = 1;
    45: op1_00_inv09 = 1;
    52: op1_00_inv09 = 1;
    46: op1_00_inv09 = 1;
    54: op1_00_inv09 = 1;
    71: op1_00_inv09 = 1;
    72: op1_00_inv09 = 1;
    40: op1_00_inv09 = 1;
    55: op1_00_inv09 = 1;
    68: op1_00_inv09 = 1;
    87: op1_00_inv09 = 1;
    59: op1_00_inv09 = 1;
    50: op1_00_inv09 = 1;
    86: op1_00_inv09 = 1;
    44: op1_00_inv09 = 1;
    56: op1_00_inv09 = 1;
    42: op1_00_inv09 = 1;
    70: op1_00_inv09 = 1;
    51: op1_00_inv09 = 1;
    62: op1_00_inv09 = 1;
    64: op1_00_inv09 = 1;
    84: op1_00_inv09 = 1;
    65: op1_00_inv09 = 1;
    85: op1_00_inv09 = 1;
    92: op1_00_inv09 = 1;
    95: op1_00_inv09 = 1;
    98: op1_00_inv09 = 1;
    114: op1_00_inv09 = 1;
    115: op1_00_inv09 = 1;
    116: op1_00_inv09 = 1;
    120: op1_00_inv09 = 1;
    122: op1_00_inv09 = 1;
    123: op1_00_inv09 = 1;
    126: op1_00_inv09 = 1;
    130: op1_00_inv09 = 1;
    default: op1_00_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の10番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in10 = reg_0201;
    15: op1_00_in10 = reg_0088;
    19: op1_00_in10 = reg_0218;
    11: op1_00_in10 = imem05_in[7:4];
    33: op1_00_in10 = reg_0405;
    81: op1_00_in10 = reg_0405;
    100: op1_00_in10 = reg_0405;
    35: op1_00_in10 = reg_0497;
    32: op1_00_in10 = reg_0466;
    26: op1_00_in10 = reg_0300;
    21: op1_00_in10 = reg_0085;
    41: op1_00_in10 = reg_0641;
    38: op1_00_in10 = imem03_in[11:8];
    39: op1_00_in10 = reg_0749;
    45: op1_00_in10 = reg_0636;
    52: op1_00_in10 = reg_0723;
    49: op1_00_in10 = reg_0862;
    46: op1_00_in10 = reg_0171;
    58: op1_00_in10 = reg_0642;
    60: op1_00_in10 = reg_0642;
    54: op1_00_in10 = reg_0708;
    48: op1_00_in10 = reg_0993;
    53: op1_00_in10 = reg_0433;
    75: op1_00_in10 = reg_0433;
    61: op1_00_in10 = reg_0462;
    67: op1_00_in10 = reg_0268;
    76: op1_00_in10 = reg_0459;
    71: op1_00_in10 = reg_0064;
    72: op1_00_in10 = reg_0172;
    40: op1_00_in10 = reg_0620;
    55: op1_00_in10 = reg_0711;
    68: op1_00_in10 = reg_0237;
    74: op1_00_in10 = reg_0009;
    87: op1_00_in10 = reg_1040;
    78: op1_00_in10 = reg_0795;
    73: op1_00_in10 = reg_0162;
    59: op1_00_in10 = reg_0072;
    50: op1_00_in10 = reg_0496;
    86: op1_00_in10 = reg_0962;
    69: op1_00_in10 = reg_0705;
    36: op1_00_in10 = reg_0606;
    44: op1_00_in10 = reg_0206;
    88: op1_00_in10 = reg_0626;
    47: op1_00_in10 = imem07_in[11:8];
    56: op1_00_in10 = reg_0341;
    42: op1_00_in10 = reg_0456;
    70: op1_00_in10 = reg_0608;
    57: op1_00_in10 = reg_0352;
    77: op1_00_in10 = reg_1107;
    51: op1_00_in10 = reg_0569;
    79: op1_00_in10 = reg_0431;
    43: op1_00_in10 = reg_0649;
    62: op1_00_in10 = reg_0640;
    80: op1_00_in10 = reg_0233;
    89: op1_00_in10 = reg_0113;
    63: op1_00_in10 = reg_0571;
    117: op1_00_in10 = reg_0571;
    82: op1_00_in10 = reg_0480;
    83: op1_00_in10 = reg_1432;
    64: op1_00_in10 = reg_0112;
    84: op1_00_in10 = reg_0752;
    65: op1_00_in10 = reg_1254;
    90: op1_00_in10 = reg_1340;
    85: op1_00_in10 = reg_0666;
    66: op1_00_in10 = reg_0974;
    91: op1_00_in10 = reg_0615;
    92: op1_00_in10 = reg_1486;
    93: op1_00_in10 = reg_0884;
    107: op1_00_in10 = reg_0884;
    94: op1_00_in10 = reg_0416;
    95: op1_00_in10 = reg_0938;
    96: op1_00_in10 = reg_0169;
    97: op1_00_in10 = reg_0494;
    98: op1_00_in10 = reg_0309;
    99: op1_00_in10 = reg_1373;
    101: op1_00_in10 = imem07_in[3:0];
    102: op1_00_in10 = reg_0380;
    103: op1_00_in10 = reg_0670;
    104: op1_00_in10 = reg_0740;
    125: op1_00_in10 = reg_0740;
    105: op1_00_in10 = reg_0256;
    106: op1_00_in10 = reg_0423;
    108: op1_00_in10 = reg_0303;
    109: op1_00_in10 = reg_0709;
    110: op1_00_in10 = reg_1418;
    111: op1_00_in10 = reg_1214;
    112: op1_00_in10 = reg_1405;
    113: op1_00_in10 = reg_0451;
    114: op1_00_in10 = reg_0712;
    115: op1_00_in10 = reg_0214;
    116: op1_00_in10 = reg_0555;
    120: op1_00_in10 = reg_0322;
    121: op1_00_in10 = imem04_in[7:4];
    122: op1_00_in10 = reg_0333;
    123: op1_00_in10 = reg_0406;
    124: op1_00_in10 = reg_0588;
    126: op1_00_in10 = reg_0294;
    128: op1_00_in10 = reg_1406;
    129: op1_00_in10 = reg_0890;
    130: op1_00_in10 = reg_0323;
    131: op1_00_in10 = reg_0167;
    default: op1_00_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    11: op1_00_inv10 = 1;
    35: op1_00_inv10 = 1;
    32: op1_00_inv10 = 1;
    21: op1_00_inv10 = 1;
    38: op1_00_inv10 = 1;
    39: op1_00_inv10 = 1;
    52: op1_00_inv10 = 1;
    46: op1_00_inv10 = 1;
    58: op1_00_inv10 = 1;
    60: op1_00_inv10 = 1;
    67: op1_00_inv10 = 1;
    72: op1_00_inv10 = 1;
    40: op1_00_inv10 = 1;
    55: op1_00_inv10 = 1;
    74: op1_00_inv10 = 1;
    73: op1_00_inv10 = 1;
    59: op1_00_inv10 = 1;
    50: op1_00_inv10 = 1;
    69: op1_00_inv10 = 1;
    44: op1_00_inv10 = 1;
    47: op1_00_inv10 = 1;
    56: op1_00_inv10 = 1;
    42: op1_00_inv10 = 1;
    70: op1_00_inv10 = 1;
    57: op1_00_inv10 = 1;
    77: op1_00_inv10 = 1;
    51: op1_00_inv10 = 1;
    43: op1_00_inv10 = 1;
    63: op1_00_inv10 = 1;
    82: op1_00_inv10 = 1;
    64: op1_00_inv10 = 1;
    66: op1_00_inv10 = 1;
    92: op1_00_inv10 = 1;
    93: op1_00_inv10 = 1;
    94: op1_00_inv10 = 1;
    95: op1_00_inv10 = 1;
    96: op1_00_inv10 = 1;
    99: op1_00_inv10 = 1;
    100: op1_00_inv10 = 1;
    102: op1_00_inv10 = 1;
    103: op1_00_inv10 = 1;
    105: op1_00_inv10 = 1;
    106: op1_00_inv10 = 1;
    108: op1_00_inv10 = 1;
    109: op1_00_inv10 = 1;
    111: op1_00_inv10 = 1;
    112: op1_00_inv10 = 1;
    115: op1_00_inv10 = 1;
    117: op1_00_inv10 = 1;
    120: op1_00_inv10 = 1;
    123: op1_00_inv10 = 1;
    125: op1_00_inv10 = 1;
    128: op1_00_inv10 = 1;
    default: op1_00_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の11番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in11 = reg_0186;
    15: op1_00_in11 = reg_0077;
    19: op1_00_in11 = reg_0199;
    11: op1_00_in11 = reg_0173;
    33: op1_00_in11 = reg_0389;
    94: op1_00_in11 = reg_0389;
    35: op1_00_in11 = reg_0494;
    32: op1_00_in11 = reg_0467;
    26: op1_00_in11 = reg_0168;
    41: op1_00_in11 = reg_0218;
    38: op1_00_in11 = reg_0573;
    39: op1_00_in11 = reg_0735;
    45: op1_00_in11 = reg_0622;
    52: op1_00_in11 = imem01_in[11:8];
    49: op1_00_in11 = reg_0835;
    46: op1_00_in11 = reg_0067;
    58: op1_00_in11 = reg_0640;
    54: op1_00_in11 = reg_0711;
    48: op1_00_in11 = reg_0892;
    60: op1_00_in11 = reg_0410;
    53: op1_00_in11 = reg_0776;
    61: op1_00_in11 = reg_1214;
    67: op1_00_in11 = reg_0870;
    76: op1_00_in11 = reg_1405;
    71: op1_00_in11 = reg_0062;
    72: op1_00_in11 = reg_0869;
    40: op1_00_in11 = reg_0102;
    55: op1_00_in11 = reg_0294;
    68: op1_00_in11 = reg_0129;
    74: op1_00_in11 = reg_0531;
    87: op1_00_in11 = reg_0454;
    78: op1_00_in11 = reg_0908;
    73: op1_00_in11 = reg_0922;
    59: op1_00_in11 = reg_0057;
    57: op1_00_in11 = reg_0057;
    50: op1_00_in11 = reg_0473;
    102: op1_00_in11 = reg_0473;
    86: op1_00_in11 = reg_0989;
    69: op1_00_in11 = reg_0009;
    36: op1_00_in11 = reg_0587;
    44: op1_00_in11 = reg_0040;
    129: op1_00_in11 = reg_0040;
    88: op1_00_in11 = reg_0846;
    47: op1_00_in11 = reg_0704;
    56: op1_00_in11 = reg_0305;
    75: op1_00_in11 = reg_0054;
    42: op1_00_in11 = reg_0433;
    70: op1_00_in11 = reg_0631;
    77: op1_00_in11 = reg_0633;
    51: op1_00_in11 = reg_0529;
    79: op1_00_in11 = reg_0435;
    43: op1_00_in11 = reg_0315;
    62: op1_00_in11 = reg_0189;
    80: op1_00_in11 = reg_0709;
    81: op1_00_in11 = reg_0388;
    89: op1_00_in11 = reg_0350;
    63: op1_00_in11 = reg_1228;
    82: op1_00_in11 = reg_0481;
    83: op1_00_in11 = reg_1417;
    64: op1_00_in11 = reg_0106;
    84: op1_00_in11 = reg_0109;
    65: op1_00_in11 = reg_0257;
    90: op1_00_in11 = reg_0462;
    85: op1_00_in11 = reg_0474;
    66: op1_00_in11 = imem06_in[7:4];
    91: op1_00_in11 = reg_0486;
    92: op1_00_in11 = reg_1485;
    93: op1_00_in11 = reg_0348;
    95: op1_00_in11 = reg_0794;
    96: op1_00_in11 = reg_0608;
    97: op1_00_in11 = reg_1451;
    98: op1_00_in11 = reg_0923;
    99: op1_00_in11 = reg_0240;
    100: op1_00_in11 = reg_0134;
    101: op1_00_in11 = imem07_in[11:8];
    103: op1_00_in11 = reg_0270;
    104: op1_00_in11 = reg_0408;
    105: op1_00_in11 = reg_1260;
    106: op1_00_in11 = reg_0879;
    107: op1_00_in11 = reg_0291;
    108: op1_00_in11 = reg_0090;
    109: op1_00_in11 = reg_1063;
    110: op1_00_in11 = reg_0459;
    111: op1_00_in11 = reg_0796;
    112: op1_00_in11 = reg_0722;
    113: op1_00_in11 = reg_0342;
    114: op1_00_in11 = reg_0839;
    115: op1_00_in11 = reg_0213;
    116: op1_00_in11 = reg_1205;
    117: op1_00_in11 = reg_1225;
    120: op1_00_in11 = reg_1235;
    121: op1_00_in11 = reg_0252;
    122: op1_00_in11 = reg_0669;
    123: op1_00_in11 = reg_1041;
    124: op1_00_in11 = reg_0975;
    125: op1_00_in11 = reg_0620;
    126: op1_00_in11 = reg_0217;
    128: op1_00_in11 = reg_0927;
    130: op1_00_in11 = reg_0308;
    131: op1_00_in11 = reg_0334;
    default: op1_00_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv11 = 1;
    15: op1_00_inv11 = 1;
    19: op1_00_inv11 = 1;
    33: op1_00_inv11 = 1;
    38: op1_00_inv11 = 1;
    45: op1_00_inv11 = 1;
    49: op1_00_inv11 = 1;
    58: op1_00_inv11 = 1;
    53: op1_00_inv11 = 1;
    61: op1_00_inv11 = 1;
    76: op1_00_inv11 = 1;
    40: op1_00_inv11 = 1;
    74: op1_00_inv11 = 1;
    87: op1_00_inv11 = 1;
    73: op1_00_inv11 = 1;
    50: op1_00_inv11 = 1;
    86: op1_00_inv11 = 1;
    36: op1_00_inv11 = 1;
    44: op1_00_inv11 = 1;
    88: op1_00_inv11 = 1;
    47: op1_00_inv11 = 1;
    42: op1_00_inv11 = 1;
    70: op1_00_inv11 = 1;
    57: op1_00_inv11 = 1;
    77: op1_00_inv11 = 1;
    51: op1_00_inv11 = 1;
    79: op1_00_inv11 = 1;
    43: op1_00_inv11 = 1;
    62: op1_00_inv11 = 1;
    81: op1_00_inv11 = 1;
    63: op1_00_inv11 = 1;
    82: op1_00_inv11 = 1;
    90: op1_00_inv11 = 1;
    66: op1_00_inv11 = 1;
    92: op1_00_inv11 = 1;
    94: op1_00_inv11 = 1;
    95: op1_00_inv11 = 1;
    102: op1_00_inv11 = 1;
    104: op1_00_inv11 = 1;
    105: op1_00_inv11 = 1;
    109: op1_00_inv11 = 1;
    111: op1_00_inv11 = 1;
    114: op1_00_inv11 = 1;
    116: op1_00_inv11 = 1;
    117: op1_00_inv11 = 1;
    124: op1_00_inv11 = 1;
    125: op1_00_inv11 = 1;
    126: op1_00_inv11 = 1;
    130: op1_00_inv11 = 1;
    default: op1_00_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の12番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in12 = reg_0171;
    15: op1_00_in12 = reg_0047;
    19: op1_00_in12 = reg_0185;
    11: op1_00_in12 = reg_0175;
    33: op1_00_in12 = reg_0351;
    35: op1_00_in12 = reg_0473;
    32: op1_00_in12 = reg_0462;
    26: op1_00_in12 = reg_0196;
    41: op1_00_in12 = reg_0428;
    38: op1_00_in12 = reg_0710;
    80: op1_00_in12 = reg_0710;
    39: op1_00_in12 = reg_0702;
    45: op1_00_in12 = reg_0584;
    52: op1_00_in12 = reg_0161;
    49: op1_00_in12 = reg_0181;
    46: op1_00_in12 = imem07_in[15:12];
    58: op1_00_in12 = reg_0722;
    54: op1_00_in12 = reg_0877;
    48: op1_00_in12 = reg_0297;
    60: op1_00_in12 = reg_0134;
    53: op1_00_in12 = reg_0933;
    61: op1_00_in12 = reg_1216;
    67: op1_00_in12 = reg_0536;
    76: op1_00_in12 = reg_0476;
    71: op1_00_in12 = reg_0016;
    77: op1_00_in12 = reg_0016;
    72: op1_00_in12 = reg_0264;
    40: op1_00_in12 = reg_0028;
    55: op1_00_in12 = reg_0839;
    68: op1_00_in12 = reg_0033;
    74: op1_00_in12 = reg_0327;
    87: op1_00_in12 = reg_0232;
    123: op1_00_in12 = reg_0232;
    78: op1_00_in12 = reg_0905;
    73: op1_00_in12 = reg_0245;
    59: op1_00_in12 = reg_0089;
    50: op1_00_in12 = reg_0475;
    70: op1_00_in12 = reg_0475;
    86: op1_00_in12 = reg_0965;
    69: op1_00_in12 = reg_0531;
    36: op1_00_in12 = reg_0562;
    44: op1_00_in12 = reg_0039;
    88: op1_00_in12 = reg_0822;
    47: op1_00_in12 = reg_0324;
    56: op1_00_in12 = reg_0862;
    75: op1_00_in12 = reg_0128;
    42: op1_00_in12 = reg_0138;
    64: op1_00_in12 = reg_0138;
    57: op1_00_in12 = reg_0027;
    51: op1_00_in12 = reg_0522;
    79: op1_00_in12 = reg_0071;
    81: op1_00_in12 = reg_0071;
    43: op1_00_in12 = reg_0070;
    62: op1_00_in12 = reg_0416;
    89: op1_00_in12 = reg_0291;
    63: op1_00_in12 = reg_0132;
    82: op1_00_in12 = reg_0734;
    83: op1_00_in12 = reg_1405;
    84: op1_00_in12 = reg_0398;
    65: op1_00_in12 = reg_0634;
    90: op1_00_in12 = reg_0574;
    85: op1_00_in12 = reg_0971;
    66: op1_00_in12 = reg_0929;
    91: op1_00_in12 = reg_0555;
    92: op1_00_in12 = reg_0576;
    93: op1_00_in12 = imem04_in[7:4];
    94: op1_00_in12 = reg_0059;
    95: op1_00_in12 = reg_0302;
    96: op1_00_in12 = reg_0561;
    97: op1_00_in12 = reg_1455;
    98: op1_00_in12 = reg_0663;
    99: op1_00_in12 = reg_0449;
    100: op1_00_in12 = reg_0203;
    101: op1_00_in12 = reg_0461;
    102: op1_00_in12 = reg_0829;
    103: op1_00_in12 = reg_0730;
    104: op1_00_in12 = reg_0591;
    105: op1_00_in12 = reg_0776;
    106: op1_00_in12 = reg_0608;
    107: op1_00_in12 = reg_1280;
    108: op1_00_in12 = reg_0872;
    109: op1_00_in12 = reg_1425;
    110: op1_00_in12 = reg_0821;
    111: op1_00_in12 = reg_0094;
    112: op1_00_in12 = reg_0201;
    113: op1_00_in12 = reg_0097;
    114: op1_00_in12 = reg_0390;
    115: op1_00_in12 = reg_1170;
    116: op1_00_in12 = reg_0460;
    117: op1_00_in12 = reg_0295;
    120: op1_00_in12 = reg_0712;
    121: op1_00_in12 = reg_0731;
    122: op1_00_in12 = reg_1209;
    124: op1_00_in12 = reg_0254;
    125: op1_00_in12 = reg_0114;
    126: op1_00_in12 = reg_0009;
    128: op1_00_in12 = reg_0189;
    129: op1_00_in12 = reg_0182;
    130: op1_00_in12 = reg_0022;
    131: op1_00_in12 = reg_1181;
    default: op1_00_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv12 = 1;
    15: op1_00_inv12 = 1;
    32: op1_00_inv12 = 1;
    26: op1_00_inv12 = 1;
    41: op1_00_inv12 = 1;
    52: op1_00_inv12 = 1;
    54: op1_00_inv12 = 1;
    48: op1_00_inv12 = 1;
    60: op1_00_inv12 = 1;
    53: op1_00_inv12 = 1;
    61: op1_00_inv12 = 1;
    40: op1_00_inv12 = 1;
    55: op1_00_inv12 = 1;
    68: op1_00_inv12 = 1;
    87: op1_00_inv12 = 1;
    78: op1_00_inv12 = 1;
    50: op1_00_inv12 = 1;
    86: op1_00_inv12 = 1;
    69: op1_00_inv12 = 1;
    36: op1_00_inv12 = 1;
    88: op1_00_inv12 = 1;
    56: op1_00_inv12 = 1;
    57: op1_00_inv12 = 1;
    51: op1_00_inv12 = 1;
    80: op1_00_inv12 = 1;
    89: op1_00_inv12 = 1;
    63: op1_00_inv12 = 1;
    82: op1_00_inv12 = 1;
    83: op1_00_inv12 = 1;
    90: op1_00_inv12 = 1;
    66: op1_00_inv12 = 1;
    92: op1_00_inv12 = 1;
    93: op1_00_inv12 = 1;
    97: op1_00_inv12 = 1;
    99: op1_00_inv12 = 1;
    100: op1_00_inv12 = 1;
    103: op1_00_inv12 = 1;
    104: op1_00_inv12 = 1;
    107: op1_00_inv12 = 1;
    108: op1_00_inv12 = 1;
    111: op1_00_inv12 = 1;
    112: op1_00_inv12 = 1;
    113: op1_00_inv12 = 1;
    124: op1_00_inv12 = 1;
    125: op1_00_inv12 = 1;
    128: op1_00_inv12 = 1;
    default: op1_00_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の13番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in13 = reg_0172;
    15: op1_00_in13 = reg_0042;
    19: op1_00_in13 = reg_0179;
    11: op1_00_in13 = reg_0151;
    33: op1_00_in13 = reg_0026;
    35: op1_00_in13 = reg_0474;
    32: op1_00_in13 = reg_0420;
    26: op1_00_in13 = reg_0184;
    41: op1_00_in13 = reg_0431;
    38: op1_00_in13 = reg_0377;
    39: op1_00_in13 = reg_0250;
    45: op1_00_in13 = reg_0568;
    52: op1_00_in13 = reg_1068;
    49: op1_00_in13 = reg_0117;
    46: op1_00_in13 = reg_0704;
    58: op1_00_in13 = reg_0189;
    54: op1_00_in13 = reg_0848;
    48: op1_00_in13 = reg_0791;
    60: op1_00_in13 = reg_0350;
    53: op1_00_in13 = reg_0128;
    97: op1_00_in13 = reg_0128;
    61: op1_00_in13 = reg_1200;
    67: op1_00_in13 = reg_1326;
    76: op1_00_in13 = reg_0928;
    71: op1_00_in13 = reg_0035;
    72: op1_00_in13 = reg_0115;
    40: op1_00_in13 = reg_0002;
    55: op1_00_in13 = reg_0008;
    74: op1_00_in13 = reg_0008;
    68: op1_00_in13 = reg_0034;
    87: op1_00_in13 = reg_0061;
    78: op1_00_in13 = reg_0960;
    73: op1_00_in13 = reg_0703;
    59: op1_00_in13 = imem01_in[3:0];
    50: op1_00_in13 = reg_0989;
    86: op1_00_in13 = reg_1518;
    69: op1_00_in13 = reg_0839;
    36: op1_00_in13 = reg_0532;
    120: op1_00_in13 = reg_0532;
    44: op1_00_in13 = reg_0014;
    88: op1_00_in13 = reg_1032;
    47: op1_00_in13 = reg_0157;
    56: op1_00_in13 = reg_0836;
    75: op1_00_in13 = reg_0126;
    42: op1_00_in13 = reg_0133;
    70: op1_00_in13 = reg_0429;
    57: op1_00_in13 = reg_0917;
    77: op1_00_in13 = reg_0578;
    51: op1_00_in13 = reg_0308;
    79: op1_00_in13 = reg_0060;
    43: op1_00_in13 = imem05_in[11:8];
    62: op1_00_in13 = reg_0134;
    80: op1_00_in13 = reg_1448;
    81: op1_00_in13 = reg_0203;
    89: op1_00_in13 = imem04_in[3:0];
    63: op1_00_in13 = reg_0171;
    82: op1_00_in13 = reg_0849;
    83: op1_00_in13 = reg_0476;
    64: op1_00_in13 = reg_0898;
    84: op1_00_in13 = reg_0528;
    65: op1_00_in13 = reg_0550;
    90: op1_00_in13 = reg_0488;
    85: op1_00_in13 = reg_0382;
    66: op1_00_in13 = reg_0925;
    91: op1_00_in13 = reg_0523;
    92: op1_00_in13 = reg_0602;
    93: op1_00_in13 = reg_0032;
    94: op1_00_in13 = imem01_in[15:12];
    95: op1_00_in13 = reg_0300;
    96: op1_00_in13 = reg_0254;
    98: op1_00_in13 = reg_0285;
    99: op1_00_in13 = reg_0861;
    100: op1_00_in13 = reg_0057;
    101: op1_00_in13 = reg_0994;
    102: op1_00_in13 = reg_0745;
    105: op1_00_in13 = reg_0745;
    103: op1_00_in13 = reg_1420;
    104: op1_00_in13 = reg_0592;
    106: op1_00_in13 = reg_1493;
    107: op1_00_in13 = reg_0425;
    108: op1_00_in13 = reg_0888;
    109: op1_00_in13 = reg_0145;
    110: op1_00_in13 = reg_0351;
    111: op1_00_in13 = reg_0698;
    113: op1_00_in13 = reg_0698;
    112: op1_00_in13 = reg_0072;
    114: op1_00_in13 = reg_0971;
    115: op1_00_in13 = imem07_in[7:4];
    116: op1_00_in13 = reg_1418;
    117: op1_00_in13 = reg_0419;
    121: op1_00_in13 = reg_0297;
    122: op1_00_in13 = reg_0730;
    123: op1_00_in13 = reg_0262;
    124: op1_00_in13 = reg_0533;
    125: op1_00_in13 = reg_0361;
    126: op1_00_in13 = imem03_in[7:4];
    128: op1_00_in13 = reg_0428;
    129: op1_00_in13 = reg_0131;
    130: op1_00_in13 = imem07_in[15:12];
    131: op1_00_in13 = reg_0939;
    default: op1_00_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv13 = 1;
    35: op1_00_inv13 = 1;
    32: op1_00_inv13 = 1;
    26: op1_00_inv13 = 1;
    41: op1_00_inv13 = 1;
    38: op1_00_inv13 = 1;
    52: op1_00_inv13 = 1;
    49: op1_00_inv13 = 1;
    58: op1_00_inv13 = 1;
    54: op1_00_inv13 = 1;
    48: op1_00_inv13 = 1;
    60: op1_00_inv13 = 1;
    53: op1_00_inv13 = 1;
    61: op1_00_inv13 = 1;
    76: op1_00_inv13 = 1;
    71: op1_00_inv13 = 1;
    72: op1_00_inv13 = 1;
    74: op1_00_inv13 = 1;
    78: op1_00_inv13 = 1;
    73: op1_00_inv13 = 1;
    59: op1_00_inv13 = 1;
    50: op1_00_inv13 = 1;
    57: op1_00_inv13 = 1;
    77: op1_00_inv13 = 1;
    81: op1_00_inv13 = 1;
    82: op1_00_inv13 = 1;
    83: op1_00_inv13 = 1;
    64: op1_00_inv13 = 1;
    84: op1_00_inv13 = 1;
    65: op1_00_inv13 = 1;
    90: op1_00_inv13 = 1;
    92: op1_00_inv13 = 1;
    93: op1_00_inv13 = 1;
    94: op1_00_inv13 = 1;
    98: op1_00_inv13 = 1;
    99: op1_00_inv13 = 1;
    102: op1_00_inv13 = 1;
    103: op1_00_inv13 = 1;
    104: op1_00_inv13 = 1;
    105: op1_00_inv13 = 1;
    106: op1_00_inv13 = 1;
    107: op1_00_inv13 = 1;
    108: op1_00_inv13 = 1;
    109: op1_00_inv13 = 1;
    111: op1_00_inv13 = 1;
    112: op1_00_inv13 = 1;
    113: op1_00_inv13 = 1;
    114: op1_00_inv13 = 1;
    116: op1_00_inv13 = 1;
    124: op1_00_inv13 = 1;
    129: op1_00_inv13 = 1;
    131: op1_00_inv13 = 1;
    default: op1_00_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の14番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in14 = reg_0155;
    15: op1_00_in14 = reg_0011;
    19: op1_00_in14 = reg_0154;
    11: op1_00_in14 = reg_0130;
    33: op1_00_in14 = reg_0027;
    35: op1_00_in14 = reg_0455;
    32: op1_00_in14 = reg_0421;
    26: op1_00_in14 = reg_0273;
    41: op1_00_in14 = reg_0405;
    38: op1_00_in14 = reg_0025;
    39: op1_00_in14 = reg_0648;
    45: op1_00_in14 = reg_0526;
    52: op1_00_in14 = reg_1069;
    49: op1_00_in14 = imem05_in[3:0];
    46: op1_00_in14 = reg_0673;
    58: op1_00_in14 = reg_0072;
    54: op1_00_in14 = reg_0069;
    102: op1_00_in14 = reg_0069;
    48: op1_00_in14 = reg_0774;
    60: op1_00_in14 = reg_0351;
    76: op1_00_in14 = reg_0351;
    53: op1_00_in14 = reg_0380;
    85: op1_00_in14 = reg_0380;
    61: op1_00_in14 = reg_0370;
    67: op1_00_in14 = reg_0160;
    71: op1_00_in14 = imem05_in[7:4];
    72: op1_00_in14 = reg_0194;
    40: op1_00_in14 = reg_0053;
    55: op1_00_in14 = reg_0024;
    68: op1_00_in14 = reg_0794;
    74: op1_00_in14 = reg_0695;
    87: op1_00_in14 = reg_1151;
    78: op1_00_in14 = reg_1508;
    73: op1_00_in14 = reg_1094;
    59: op1_00_in14 = reg_0547;
    50: op1_00_in14 = reg_0970;
    86: op1_00_in14 = reg_0190;
    69: op1_00_in14 = reg_1392;
    36: op1_00_in14 = reg_0497;
    44: op1_00_in14 = reg_0754;
    88: op1_00_in14 = reg_0745;
    47: op1_00_in14 = reg_0779;
    56: op1_00_in14 = reg_0338;
    75: op1_00_in14 = reg_0106;
    42: op1_00_in14 = reg_0126;
    70: op1_00_in14 = reg_0382;
    57: op1_00_in14 = reg_0611;
    77: op1_00_in14 = reg_1431;
    51: op1_00_in14 = reg_0244;
    79: op1_00_in14 = reg_1322;
    43: op1_00_in14 = reg_0301;
    62: op1_00_in14 = reg_0026;
    80: op1_00_in14 = reg_1149;
    81: op1_00_in14 = reg_0057;
    112: op1_00_in14 = reg_0057;
    89: op1_00_in14 = reg_0034;
    63: op1_00_in14 = reg_0308;
    82: op1_00_in14 = reg_0426;
    83: op1_00_in14 = reg_0431;
    128: op1_00_in14 = reg_0431;
    64: op1_00_in14 = reg_0712;
    84: op1_00_in14 = reg_0568;
    65: op1_00_in14 = reg_0468;
    90: op1_00_in14 = reg_0681;
    66: op1_00_in14 = reg_0859;
    91: op1_00_in14 = reg_0250;
    92: op1_00_in14 = reg_0344;
    93: op1_00_in14 = reg_1372;
    94: op1_00_in14 = reg_1032;
    95: op1_00_in14 = reg_0601;
    96: op1_00_in14 = reg_1343;
    97: op1_00_in14 = reg_0112;
    98: op1_00_in14 = reg_0408;
    99: op1_00_in14 = reg_0014;
    100: op1_00_in14 = reg_0122;
    101: op1_00_in14 = reg_1060;
    103: op1_00_in14 = reg_0780;
    104: op1_00_in14 = reg_0050;
    105: op1_00_in14 = reg_0897;
    106: op1_00_in14 = reg_1074;
    107: op1_00_in14 = imem04_in[7:4];
    108: op1_00_in14 = reg_0492;
    109: op1_00_in14 = reg_0000;
    110: op1_00_in14 = reg_0428;
    111: op1_00_in14 = reg_1143;
    113: op1_00_in14 = reg_0835;
    114: op1_00_in14 = reg_1455;
    115: op1_00_in14 = imem07_in[11:8];
    116: op1_00_in14 = reg_0821;
    117: op1_00_in14 = reg_0119;
    120: op1_00_in14 = reg_0822;
    121: op1_00_in14 = reg_1083;
    122: op1_00_in14 = reg_0696;
    123: op1_00_in14 = reg_1146;
    124: op1_00_in14 = reg_0429;
    125: op1_00_in14 = reg_0228;
    126: op1_00_in14 = reg_0758;
    129: op1_00_in14 = reg_0697;
    130: op1_00_in14 = reg_0103;
    131: op1_00_in14 = reg_1163;
    default: op1_00_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv14 = 1;
    11: op1_00_inv14 = 1;
    33: op1_00_inv14 = 1;
    35: op1_00_inv14 = 1;
    32: op1_00_inv14 = 1;
    26: op1_00_inv14 = 1;
    41: op1_00_inv14 = 1;
    39: op1_00_inv14 = 1;
    52: op1_00_inv14 = 1;
    46: op1_00_inv14 = 1;
    61: op1_00_inv14 = 1;
    76: op1_00_inv14 = 1;
    72: op1_00_inv14 = 1;
    40: op1_00_inv14 = 1;
    74: op1_00_inv14 = 1;
    87: op1_00_inv14 = 1;
    78: op1_00_inv14 = 1;
    73: op1_00_inv14 = 1;
    50: op1_00_inv14 = 1;
    69: op1_00_inv14 = 1;
    88: op1_00_inv14 = 1;
    70: op1_00_inv14 = 1;
    57: op1_00_inv14 = 1;
    62: op1_00_inv14 = 1;
    80: op1_00_inv14 = 1;
    81: op1_00_inv14 = 1;
    89: op1_00_inv14 = 1;
    63: op1_00_inv14 = 1;
    83: op1_00_inv14 = 1;
    64: op1_00_inv14 = 1;
    84: op1_00_inv14 = 1;
    90: op1_00_inv14 = 1;
    85: op1_00_inv14 = 1;
    66: op1_00_inv14 = 1;
    91: op1_00_inv14 = 1;
    93: op1_00_inv14 = 1;
    95: op1_00_inv14 = 1;
    96: op1_00_inv14 = 1;
    97: op1_00_inv14 = 1;
    100: op1_00_inv14 = 1;
    101: op1_00_inv14 = 1;
    103: op1_00_inv14 = 1;
    106: op1_00_inv14 = 1;
    107: op1_00_inv14 = 1;
    111: op1_00_inv14 = 1;
    112: op1_00_inv14 = 1;
    115: op1_00_inv14 = 1;
    117: op1_00_inv14 = 1;
    120: op1_00_inv14 = 1;
    121: op1_00_inv14 = 1;
    122: op1_00_inv14 = 1;
    126: op1_00_inv14 = 1;
    default: op1_00_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の15番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in15 = reg_0134;
    41: op1_00_in15 = reg_0134;
    15: op1_00_in15 = imem02_in[7:4];
    19: op1_00_in15 = reg_0143;
    11: op1_00_in15 = reg_0131;
    33: op1_00_in15 = imem01_in[3:0];
    35: op1_00_in15 = reg_0429;
    32: op1_00_in15 = reg_0412;
    26: op1_00_in15 = reg_0251;
    38: op1_00_in15 = reg_0293;
    39: op1_00_in15 = reg_0649;
    45: op1_00_in15 = reg_0527;
    52: op1_00_in15 = reg_1032;
    49: op1_00_in15 = reg_0173;
    46: op1_00_in15 = reg_0672;
    58: op1_00_in15 = reg_0122;
    81: op1_00_in15 = reg_0122;
    54: op1_00_in15 = reg_0276;
    48: op1_00_in15 = reg_0029;
    60: op1_00_in15 = reg_0059;
    53: op1_00_in15 = reg_0381;
    85: op1_00_in15 = reg_0381;
    61: op1_00_in15 = reg_0341;
    67: op1_00_in15 = reg_0827;
    76: op1_00_in15 = reg_0073;
    71: op1_00_in15 = imem05_in[15:12];
    72: op1_00_in15 = reg_0141;
    55: op1_00_in15 = reg_0068;
    68: op1_00_in15 = reg_0391;
    74: op1_00_in15 = imem03_in[15:12];
    87: op1_00_in15 = reg_0904;
    78: op1_00_in15 = reg_1504;
    73: op1_00_in15 = reg_0030;
    59: op1_00_in15 = reg_0550;
    50: op1_00_in15 = reg_0935;
    86: op1_00_in15 = reg_1301;
    69: op1_00_in15 = reg_0280;
    36: op1_00_in15 = reg_0475;
    44: op1_00_in15 = reg_0193;
    88: op1_00_in15 = reg_1078;
    47: op1_00_in15 = reg_0661;
    56: op1_00_in15 = reg_0339;
    75: op1_00_in15 = reg_0105;
    42: op1_00_in15 = reg_0380;
    70: op1_00_in15 = reg_0496;
    57: op1_00_in15 = reg_0612;
    77: op1_00_in15 = reg_0877;
    51: op1_00_in15 = reg_0271;
    79: op1_00_in15 = reg_0027;
    43: op1_00_in15 = reg_0872;
    62: op1_00_in15 = reg_0917;
    80: op1_00_in15 = imem03_in[11:8];
    89: op1_00_in15 = reg_1338;
    63: op1_00_in15 = reg_0152;
    82: op1_00_in15 = reg_0975;
    83: op1_00_in15 = reg_0203;
    64: op1_00_in15 = reg_0307;
    84: op1_00_in15 = reg_0371;
    65: op1_00_in15 = reg_0469;
    90: op1_00_in15 = reg_1233;
    66: op1_00_in15 = reg_0752;
    91: op1_00_in15 = reg_1027;
    92: op1_00_in15 = reg_0037;
    93: op1_00_in15 = reg_1367;
    107: op1_00_in15 = reg_1367;
    94: op1_00_in15 = reg_0355;
    95: op1_00_in15 = reg_0603;
    96: op1_00_in15 = reg_0712;
    97: op1_00_in15 = reg_1140;
    98: op1_00_in15 = reg_0137;
    99: op1_00_in15 = imem06_in[15:12];
    100: op1_00_in15 = imem01_in[7:4];
    112: op1_00_in15 = imem01_in[7:4];
    101: op1_00_in15 = reg_0135;
    102: op1_00_in15 = reg_0632;
    103: op1_00_in15 = reg_0116;
    105: op1_00_in15 = reg_0802;
    106: op1_00_in15 = reg_0497;
    108: op1_00_in15 = reg_1348;
    109: op1_00_in15 = reg_0180;
    110: op1_00_in15 = reg_0431;
    111: op1_00_in15 = reg_0368;
    113: op1_00_in15 = reg_1312;
    114: op1_00_in15 = reg_0128;
    115: op1_00_in15 = imem07_in[15:12];
    116: op1_00_in15 = reg_1405;
    117: op1_00_in15 = reg_1202;
    120: op1_00_in15 = reg_0495;
    121: op1_00_in15 = reg_1214;
    122: op1_00_in15 = reg_0863;
    123: op1_00_in15 = reg_1151;
    124: op1_00_in15 = reg_1455;
    125: op1_00_in15 = reg_1351;
    126: op1_00_in15 = reg_0759;
    128: op1_00_in15 = reg_0389;
    129: op1_00_in15 = reg_0940;
    130: op1_00_in15 = reg_0087;
    131: op1_00_in15 = reg_0090;
    default: op1_00_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv15 = 1;
    19: op1_00_inv15 = 1;
    33: op1_00_inv15 = 1;
    32: op1_00_inv15 = 1;
    26: op1_00_inv15 = 1;
    41: op1_00_inv15 = 1;
    39: op1_00_inv15 = 1;
    49: op1_00_inv15 = 1;
    61: op1_00_inv15 = 1;
    67: op1_00_inv15 = 1;
    71: op1_00_inv15 = 1;
    68: op1_00_inv15 = 1;
    87: op1_00_inv15 = 1;
    59: op1_00_inv15 = 1;
    50: op1_00_inv15 = 1;
    44: op1_00_inv15 = 1;
    56: op1_00_inv15 = 1;
    42: op1_00_inv15 = 1;
    51: op1_00_inv15 = 1;
    79: op1_00_inv15 = 1;
    43: op1_00_inv15 = 1;
    62: op1_00_inv15 = 1;
    80: op1_00_inv15 = 1;
    83: op1_00_inv15 = 1;
    85: op1_00_inv15 = 1;
    66: op1_00_inv15 = 1;
    91: op1_00_inv15 = 1;
    93: op1_00_inv15 = 1;
    94: op1_00_inv15 = 1;
    95: op1_00_inv15 = 1;
    98: op1_00_inv15 = 1;
    101: op1_00_inv15 = 1;
    102: op1_00_inv15 = 1;
    105: op1_00_inv15 = 1;
    106: op1_00_inv15 = 1;
    108: op1_00_inv15 = 1;
    111: op1_00_inv15 = 1;
    121: op1_00_inv15 = 1;
    123: op1_00_inv15 = 1;
    128: op1_00_inv15 = 1;
    129: op1_00_inv15 = 1;
    130: op1_00_inv15 = 1;
    default: op1_00_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の16番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in16 = reg_0135;
    15: op1_00_in16 = reg_0227;
    19: op1_00_in16 = reg_0121;
    11: op1_00_in16 = reg_0118;
    33: op1_00_in16 = reg_0572;
    35: op1_00_in16 = reg_0390;
    32: op1_00_in16 = reg_0370;
    26: op1_00_in16 = imem06_in[11:8];
    41: op1_00_in16 = reg_0350;
    38: op1_00_in16 = reg_0000;
    39: op1_00_in16 = reg_0601;
    45: op1_00_in16 = reg_0296;
    52: op1_00_in16 = reg_1034;
    49: op1_00_in16 = reg_0992;
    46: op1_00_in16 = reg_0777;
    58: op1_00_in16 = imem01_in[11:8];
    54: op1_00_in16 = imem03_in[3:0];
    48: op1_00_in16 = reg_0366;
    60: op1_00_in16 = reg_0027;
    53: op1_00_in16 = reg_0898;
    61: op1_00_in16 = reg_0095;
    56: op1_00_in16 = reg_0095;
    67: op1_00_in16 = reg_0264;
    93: op1_00_in16 = reg_0264;
    76: op1_00_in16 = reg_0075;
    71: op1_00_in16 = reg_0579;
    72: op1_00_in16 = reg_0528;
    55: op1_00_in16 = reg_0279;
    68: op1_00_in16 = reg_0315;
    74: op1_00_in16 = reg_1000;
    87: op1_00_in16 = reg_1107;
    78: op1_00_in16 = reg_0161;
    73: op1_00_in16 = reg_0413;
    59: op1_00_in16 = reg_0238;
    50: op1_00_in16 = reg_0111;
    86: op1_00_in16 = reg_1208;
    69: op1_00_in16 = reg_0235;
    36: op1_00_in16 = reg_0429;
    44: op1_00_in16 = imem06_in[7:4];
    88: op1_00_in16 = reg_1006;
    47: op1_00_in16 = reg_0285;
    75: op1_00_in16 = reg_0496;
    42: op1_00_in16 = reg_0056;
    70: op1_00_in16 = reg_1433;
    57: op1_00_in16 = reg_0335;
    77: op1_00_in16 = reg_0996;
    51: op1_00_in16 = reg_0023;
    79: op1_00_in16 = imem01_in[3:0];
    81: op1_00_in16 = imem01_in[3:0];
    43: op1_00_in16 = reg_0130;
    62: op1_00_in16 = reg_0822;
    80: op1_00_in16 = reg_1001;
    89: op1_00_in16 = reg_0297;
    63: op1_00_in16 = reg_0214;
    82: op1_00_in16 = reg_1368;
    83: op1_00_in16 = reg_0026;
    64: op1_00_in16 = reg_0153;
    84: op1_00_in16 = reg_0215;
    65: op1_00_in16 = reg_0430;
    90: op1_00_in16 = reg_0421;
    85: op1_00_in16 = imem02_in[7:4];
    66: op1_00_in16 = reg_0110;
    103: op1_00_in16 = reg_0110;
    91: op1_00_in16 = reg_0221;
    92: op1_00_in16 = imem06_in[3:0];
    94: op1_00_in16 = reg_0163;
    95: op1_00_in16 = reg_0449;
    108: op1_00_in16 = reg_0449;
    96: op1_00_in16 = reg_0532;
    97: op1_00_in16 = reg_0829;
    98: op1_00_in16 = reg_0084;
    99: op1_00_in16 = reg_0905;
    100: op1_00_in16 = reg_0547;
    101: op1_00_in16 = reg_0457;
    102: op1_00_in16 = reg_1515;
    105: op1_00_in16 = reg_1078;
    106: op1_00_in16 = reg_1260;
    107: op1_00_in16 = reg_0088;
    109: op1_00_in16 = reg_1495;
    110: op1_00_in16 = reg_0071;
    111: op1_00_in16 = reg_1146;
    112: op1_00_in16 = reg_0010;
    113: op1_00_in16 = reg_1189;
    114: op1_00_in16 = reg_0126;
    115: op1_00_in16 = reg_0993;
    116: op1_00_in16 = reg_0886;
    117: op1_00_in16 = reg_0015;
    120: op1_00_in16 = reg_0778;
    121: op1_00_in16 = reg_0599;
    122: op1_00_in16 = reg_0827;
    123: op1_00_in16 = reg_0236;
    124: op1_00_in16 = reg_0382;
    125: op1_00_in16 = reg_0001;
    126: op1_00_in16 = reg_0233;
    128: op1_00_in16 = reg_0072;
    129: op1_00_in16 = reg_0792;
    130: op1_00_in16 = reg_0994;
    131: op1_00_in16 = reg_0736;
    default: op1_00_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv16 = 1;
    15: op1_00_inv16 = 1;
    11: op1_00_inv16 = 1;
    38: op1_00_inv16 = 1;
    45: op1_00_inv16 = 1;
    52: op1_00_inv16 = 1;
    46: op1_00_inv16 = 1;
    58: op1_00_inv16 = 1;
    54: op1_00_inv16 = 1;
    60: op1_00_inv16 = 1;
    61: op1_00_inv16 = 1;
    76: op1_00_inv16 = 1;
    71: op1_00_inv16 = 1;
    68: op1_00_inv16 = 1;
    74: op1_00_inv16 = 1;
    87: op1_00_inv16 = 1;
    78: op1_00_inv16 = 1;
    73: op1_00_inv16 = 1;
    36: op1_00_inv16 = 1;
    44: op1_00_inv16 = 1;
    88: op1_00_inv16 = 1;
    47: op1_00_inv16 = 1;
    56: op1_00_inv16 = 1;
    75: op1_00_inv16 = 1;
    70: op1_00_inv16 = 1;
    51: op1_00_inv16 = 1;
    79: op1_00_inv16 = 1;
    43: op1_00_inv16 = 1;
    81: op1_00_inv16 = 1;
    89: op1_00_inv16 = 1;
    63: op1_00_inv16 = 1;
    82: op1_00_inv16 = 1;
    83: op1_00_inv16 = 1;
    90: op1_00_inv16 = 1;
    85: op1_00_inv16 = 1;
    66: op1_00_inv16 = 1;
    93: op1_00_inv16 = 1;
    96: op1_00_inv16 = 1;
    99: op1_00_inv16 = 1;
    102: op1_00_inv16 = 1;
    105: op1_00_inv16 = 1;
    106: op1_00_inv16 = 1;
    107: op1_00_inv16 = 1;
    109: op1_00_inv16 = 1;
    110: op1_00_inv16 = 1;
    113: op1_00_inv16 = 1;
    120: op1_00_inv16 = 1;
    122: op1_00_inv16 = 1;
    124: op1_00_inv16 = 1;
    128: op1_00_inv16 = 1;
    default: op1_00_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の17番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in17 = reg_0136;
    15: op1_00_in17 = reg_0216;
    19: op1_00_in17 = reg_0104;
    11: op1_00_in17 = reg_0090;
    33: op1_00_in17 = reg_0553;
    35: op1_00_in17 = reg_0382;
    32: op1_00_in17 = reg_0341;
    26: op1_00_in17 = reg_0396;
    41: op1_00_in17 = reg_0072;
    38: op1_00_in17 = reg_0048;
    39: op1_00_in17 = reg_0602;
    45: op1_00_in17 = reg_0308;
    52: op1_00_in17 = reg_0575;
    49: op1_00_in17 = reg_0334;
    46: op1_00_in17 = reg_0663;
    58: op1_00_in17 = reg_1254;
    54: op1_00_in17 = reg_1149;
    48: op1_00_in17 = reg_0739;
    60: op1_00_in17 = imem01_in[3:0];
    53: op1_00_in17 = reg_0294;
    64: op1_00_in17 = reg_0294;
    61: op1_00_in17 = reg_0209;
    87: op1_00_in17 = reg_0209;
    67: op1_00_in17 = reg_0637;
    76: op1_00_in17 = reg_0060;
    71: op1_00_in17 = reg_0833;
    72: op1_00_in17 = reg_0570;
    55: op1_00_in17 = reg_0280;
    68: op1_00_in17 = reg_0750;
    74: op1_00_in17 = reg_0699;
    78: op1_00_in17 = reg_0718;
    73: op1_00_in17 = reg_0114;
    59: op1_00_in17 = reg_0982;
    50: op1_00_in17 = reg_0112;
    86: op1_00_in17 = reg_0107;
    69: op1_00_in17 = imem03_in[7:4];
    36: op1_00_in17 = reg_0436;
    44: op1_00_in17 = reg_0906;
    88: op1_00_in17 = reg_0255;
    105: op1_00_in17 = reg_0255;
    47: op1_00_in17 = reg_0103;
    56: op1_00_in17 = reg_0210;
    75: op1_00_in17 = reg_0379;
    42: op1_00_in17 = reg_0307;
    70: op1_00_in17 = reg_0897;
    57: op1_00_in17 = imem01_in[15:12];
    79: op1_00_in17 = imem01_in[15:12];
    81: op1_00_in17 = imem01_in[15:12];
    77: op1_00_in17 = reg_0346;
    51: op1_00_in17 = reg_0152;
    43: op1_00_in17 = reg_0274;
    62: op1_00_in17 = reg_0788;
    80: op1_00_in17 = reg_0823;
    89: op1_00_in17 = reg_0488;
    63: op1_00_in17 = reg_0213;
    82: op1_00_in17 = reg_1367;
    83: op1_00_in17 = reg_0161;
    99: op1_00_in17 = reg_0161;
    84: op1_00_in17 = imem07_in[11:8];
    65: op1_00_in17 = reg_0930;
    90: op1_00_in17 = reg_0599;
    85: op1_00_in17 = reg_1098;
    66: op1_00_in17 = reg_0374;
    103: op1_00_in17 = reg_0374;
    91: op1_00_in17 = reg_0485;
    92: op1_00_in17 = reg_0931;
    93: op1_00_in17 = reg_0034;
    94: op1_00_in17 = reg_0550;
    95: op1_00_in17 = reg_0151;
    108: op1_00_in17 = reg_0151;
    96: op1_00_in17 = reg_0822;
    97: op1_00_in17 = reg_0560;
    98: op1_00_in17 = reg_0123;
    100: op1_00_in17 = reg_0743;
    101: op1_00_in17 = reg_0157;
    102: op1_00_in17 = imem03_in[15:12];
    106: op1_00_in17 = reg_1455;
    107: op1_00_in17 = reg_0264;
    109: op1_00_in17 = reg_0142;
    110: op1_00_in17 = reg_0075;
    111: op1_00_in17 = reg_1189;
    112: op1_00_in17 = reg_0746;
    113: op1_00_in17 = reg_0095;
    114: op1_00_in17 = reg_0111;
    115: op1_00_in17 = reg_0667;
    116: op1_00_in17 = reg_0722;
    117: op1_00_in17 = imem07_in[3:0];
    120: op1_00_in17 = reg_0972;
    121: op1_00_in17 = reg_0199;
    122: op1_00_in17 = reg_0115;
    123: op1_00_in17 = reg_0117;
    124: op1_00_in17 = reg_0496;
    125: op1_00_in17 = reg_0004;
    126: op1_00_in17 = reg_0185;
    128: op1_00_in17 = reg_1321;
    129: op1_00_in17 = reg_0318;
    130: op1_00_in17 = reg_0140;
    131: op1_00_in17 = reg_0066;
    default: op1_00_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_00_inv17 = 1;
    35: op1_00_inv17 = 1;
    39: op1_00_inv17 = 1;
    45: op1_00_inv17 = 1;
    49: op1_00_inv17 = 1;
    54: op1_00_inv17 = 1;
    53: op1_00_inv17 = 1;
    67: op1_00_inv17 = 1;
    71: op1_00_inv17 = 1;
    55: op1_00_inv17 = 1;
    68: op1_00_inv17 = 1;
    74: op1_00_inv17 = 1;
    78: op1_00_inv17 = 1;
    59: op1_00_inv17 = 1;
    50: op1_00_inv17 = 1;
    86: op1_00_inv17 = 1;
    69: op1_00_inv17 = 1;
    44: op1_00_inv17 = 1;
    88: op1_00_inv17 = 1;
    42: op1_00_inv17 = 1;
    77: op1_00_inv17 = 1;
    79: op1_00_inv17 = 1;
    81: op1_00_inv17 = 1;
    89: op1_00_inv17 = 1;
    82: op1_00_inv17 = 1;
    83: op1_00_inv17 = 1;
    85: op1_00_inv17 = 1;
    91: op1_00_inv17 = 1;
    93: op1_00_inv17 = 1;
    94: op1_00_inv17 = 1;
    95: op1_00_inv17 = 1;
    96: op1_00_inv17 = 1;
    97: op1_00_inv17 = 1;
    98: op1_00_inv17 = 1;
    99: op1_00_inv17 = 1;
    101: op1_00_inv17 = 1;
    102: op1_00_inv17 = 1;
    107: op1_00_inv17 = 1;
    108: op1_00_inv17 = 1;
    109: op1_00_inv17 = 1;
    110: op1_00_inv17 = 1;
    112: op1_00_inv17 = 1;
    114: op1_00_inv17 = 1;
    115: op1_00_inv17 = 1;
    116: op1_00_inv17 = 1;
    117: op1_00_inv17 = 1;
    123: op1_00_inv17 = 1;
    124: op1_00_inv17 = 1;
    126: op1_00_inv17 = 1;
    128: op1_00_inv17 = 1;
    129: op1_00_inv17 = 1;
    default: op1_00_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の18番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in18 = reg_0122;
    15: op1_00_in18 = reg_0217;
    19: op1_00_in18 = reg_0070;
    109: op1_00_in18 = reg_0070;
    11: op1_00_in18 = reg_0066;
    33: op1_00_in18 = reg_0549;
    35: op1_00_in18 = reg_0322;
    32: op1_00_in18 = reg_0305;
    26: op1_00_in18 = reg_0374;
    67: op1_00_in18 = reg_0374;
    41: op1_00_in18 = reg_0058;
    110: op1_00_in18 = reg_0058;
    38: op1_00_in18 = reg_0505;
    39: op1_00_in18 = reg_0565;
    45: op1_00_in18 = reg_0461;
    52: op1_00_in18 = reg_0984;
    49: op1_00_in18 = reg_0332;
    46: op1_00_in18 = reg_0740;
    58: op1_00_in18 = reg_0788;
    81: op1_00_in18 = reg_0788;
    54: op1_00_in18 = reg_0232;
    48: op1_00_in18 = reg_0408;
    60: op1_00_in18 = reg_0257;
    53: op1_00_in18 = reg_0876;
    61: op1_00_in18 = reg_0061;
    76: op1_00_in18 = reg_0072;
    71: op1_00_in18 = reg_0877;
    72: op1_00_in18 = reg_0345;
    55: op1_00_in18 = reg_1132;
    68: op1_00_in18 = reg_1298;
    74: op1_00_in18 = reg_0444;
    87: op1_00_in18 = reg_0065;
    78: op1_00_in18 = reg_1303;
    73: op1_00_in18 = reg_0228;
    59: op1_00_in18 = reg_0968;
    50: op1_00_in18 = reg_0105;
    86: op1_00_in18 = reg_0882;
    69: op1_00_in18 = reg_0375;
    36: op1_00_in18 = reg_0128;
    106: op1_00_in18 = reg_0128;
    44: op1_00_in18 = reg_0869;
    88: op1_00_in18 = reg_0006;
    47: op1_00_in18 = reg_0114;
    56: op1_00_in18 = reg_0208;
    75: op1_00_in18 = reg_0068;
    42: op1_00_in18 = imem02_in[3:0];
    70: op1_00_in18 = reg_0820;
    100: op1_00_in18 = reg_0820;
    57: op1_00_in18 = reg_1071;
    77: op1_00_in18 = imem05_in[3:0];
    51: op1_00_in18 = reg_0213;
    79: op1_00_in18 = reg_1290;
    43: op1_00_in18 = reg_0037;
    62: op1_00_in18 = reg_1253;
    80: op1_00_in18 = reg_0707;
    89: op1_00_in18 = reg_1233;
    63: op1_00_in18 = reg_0490;
    82: op1_00_in18 = reg_1339;
    83: op1_00_in18 = reg_0277;
    64: op1_00_in18 = reg_0846;
    84: op1_00_in18 = reg_0786;
    65: op1_00_in18 = reg_0149;
    90: op1_00_in18 = reg_0320;
    85: op1_00_in18 = reg_0695;
    66: op1_00_in18 = reg_0528;
    91: op1_00_in18 = reg_1454;
    92: op1_00_in18 = reg_0906;
    93: op1_00_in18 = reg_0797;
    94: op1_00_in18 = reg_0798;
    95: op1_00_in18 = imem06_in[3:0];
    96: op1_00_in18 = reg_0497;
    97: op1_00_in18 = reg_1492;
    98: op1_00_in18 = reg_1182;
    99: op1_00_in18 = reg_0730;
    101: op1_00_in18 = reg_0030;
    102: op1_00_in18 = reg_0783;
    103: op1_00_in18 = reg_0586;
    105: op1_00_in18 = imem03_in[11:8];
    107: op1_00_in18 = reg_0531;
    108: op1_00_in18 = imem06_in[7:4];
    111: op1_00_in18 = reg_0236;
    112: op1_00_in18 = reg_0787;
    113: op1_00_in18 = reg_0420;
    114: op1_00_in18 = reg_0307;
    115: op1_00_in18 = reg_0924;
    116: op1_00_in18 = reg_0405;
    117: op1_00_in18 = reg_0050;
    120: op1_00_in18 = reg_1450;
    121: op1_00_in18 = reg_0451;
    122: op1_00_in18 = reg_0110;
    123: op1_00_in18 = reg_1107;
    124: op1_00_in18 = reg_0745;
    125: op1_00_in18 = reg_0521;
    126: op1_00_in18 = reg_0154;
    128: op1_00_in18 = reg_1322;
    129: op1_00_in18 = reg_0243;
    130: op1_00_in18 = reg_0157;
    131: op1_00_in18 = reg_0347;
    default: op1_00_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv18 = 1;
    15: op1_00_inv18 = 1;
    19: op1_00_inv18 = 1;
    11: op1_00_inv18 = 1;
    33: op1_00_inv18 = 1;
    35: op1_00_inv18 = 1;
    41: op1_00_inv18 = 1;
    38: op1_00_inv18 = 1;
    39: op1_00_inv18 = 1;
    49: op1_00_inv18 = 1;
    46: op1_00_inv18 = 1;
    58: op1_00_inv18 = 1;
    54: op1_00_inv18 = 1;
    48: op1_00_inv18 = 1;
    60: op1_00_inv18 = 1;
    61: op1_00_inv18 = 1;
    76: op1_00_inv18 = 1;
    71: op1_00_inv18 = 1;
    55: op1_00_inv18 = 1;
    68: op1_00_inv18 = 1;
    74: op1_00_inv18 = 1;
    78: op1_00_inv18 = 1;
    59: op1_00_inv18 = 1;
    69: op1_00_inv18 = 1;
    36: op1_00_inv18 = 1;
    44: op1_00_inv18 = 1;
    47: op1_00_inv18 = 1;
    56: op1_00_inv18 = 1;
    75: op1_00_inv18 = 1;
    79: op1_00_inv18 = 1;
    62: op1_00_inv18 = 1;
    80: op1_00_inv18 = 1;
    81: op1_00_inv18 = 1;
    63: op1_00_inv18 = 1;
    82: op1_00_inv18 = 1;
    84: op1_00_inv18 = 1;
    65: op1_00_inv18 = 1;
    90: op1_00_inv18 = 1;
    66: op1_00_inv18 = 1;
    93: op1_00_inv18 = 1;
    94: op1_00_inv18 = 1;
    95: op1_00_inv18 = 1;
    96: op1_00_inv18 = 1;
    97: op1_00_inv18 = 1;
    102: op1_00_inv18 = 1;
    105: op1_00_inv18 = 1;
    109: op1_00_inv18 = 1;
    110: op1_00_inv18 = 1;
    112: op1_00_inv18 = 1;
    114: op1_00_inv18 = 1;
    115: op1_00_inv18 = 1;
    116: op1_00_inv18 = 1;
    117: op1_00_inv18 = 1;
    122: op1_00_inv18 = 1;
    126: op1_00_inv18 = 1;
    129: op1_00_inv18 = 1;
    default: op1_00_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の19番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in19 = reg_0089;
    15: op1_00_in19 = reg_0197;
    19: op1_00_in19 = reg_0048;
    11: op1_00_in19 = reg_0045;
    33: op1_00_in19 = reg_0486;
    35: op1_00_in19 = reg_0306;
    32: op1_00_in19 = reg_0319;
    26: op1_00_in19 = reg_0265;
    41: op1_00_in19 = reg_0005;
    38: op1_00_in19 = reg_0506;
    39: op1_00_in19 = reg_0540;
    45: op1_00_in19 = reg_0270;
    52: op1_00_in19 = reg_0985;
    49: op1_00_in19 = reg_0938;
    46: op1_00_in19 = reg_0618;
    58: op1_00_in19 = reg_0746;
    54: op1_00_in19 = reg_0789;
    48: op1_00_in19 = reg_0621;
    60: op1_00_in19 = reg_0239;
    53: op1_00_in19 = reg_0878;
    61: op1_00_in19 = reg_0035;
    67: op1_00_in19 = reg_0586;
    76: op1_00_in19 = reg_0057;
    71: op1_00_in19 = reg_1168;
    72: op1_00_in19 = reg_0323;
    55: op1_00_in19 = reg_0288;
    68: op1_00_in19 = reg_0735;
    74: op1_00_in19 = reg_1449;
    87: op1_00_in19 = reg_0095;
    78: op1_00_in19 = reg_0141;
    73: op1_00_in19 = reg_0052;
    59: op1_00_in19 = reg_0439;
    50: op1_00_in19 = reg_0380;
    86: op1_00_in19 = reg_0505;
    69: op1_00_in19 = reg_0559;
    36: op1_00_in19 = reg_0105;
    44: op1_00_in19 = reg_0397;
    88: op1_00_in19 = reg_1515;
    47: op1_00_in19 = reg_0028;
    56: op1_00_in19 = reg_0061;
    75: op1_00_in19 = reg_0069;
    42: op1_00_in19 = reg_0848;
    70: op1_00_in19 = reg_0121;
    57: op1_00_in19 = reg_0372;
    77: op1_00_in19 = reg_0986;
    51: op1_00_in19 = reg_0017;
    79: op1_00_in19 = reg_0166;
    43: op1_00_in19 = reg_0194;
    62: op1_00_in19 = reg_1033;
    80: op1_00_in19 = reg_0541;
    81: op1_00_in19 = reg_0754;
    89: op1_00_in19 = reg_0796;
    63: op1_00_in19 = reg_0600;
    82: op1_00_in19 = reg_1340;
    83: op1_00_in19 = reg_0331;
    64: op1_00_in19 = reg_0008;
    84: op1_00_in19 = reg_1440;
    65: op1_00_in19 = reg_0148;
    90: op1_00_in19 = reg_0342;
    85: op1_00_in19 = reg_0563;
    66: op1_00_in19 = reg_0568;
    91: op1_00_in19 = reg_0961;
    92: op1_00_in19 = reg_0316;
    93: op1_00_in19 = reg_1257;
    94: op1_00_in19 = reg_0612;
    95: op1_00_in19 = imem06_in[15:12];
    96: op1_00_in19 = reg_0432;
    97: op1_00_in19 = reg_1098;
    99: op1_00_in19 = reg_0696;
    100: op1_00_in19 = reg_0966;
    101: op1_00_in19 = reg_0287;
    102: op1_00_in19 = reg_0000;
    103: op1_00_in19 = reg_0619;
    105: op1_00_in19 = reg_1145;
    106: op1_00_in19 = reg_0125;
    107: op1_00_in19 = reg_0500;
    108: op1_00_in19 = reg_0730;
    109: op1_00_in19 = reg_1300;
    110: op1_00_in19 = reg_1324;
    111: op1_00_in19 = reg_0209;
    112: op1_00_in19 = reg_0572;
    113: op1_00_in19 = imem05_in[15:12];
    114: op1_00_in19 = reg_0903;
    115: op1_00_in19 = reg_0779;
    116: op1_00_in19 = reg_0134;
    117: op1_00_in19 = reg_0478;
    120: op1_00_in19 = reg_0106;
    121: op1_00_in19 = reg_0033;
    122: op1_00_in19 = reg_0718;
    123: op1_00_in19 = reg_0536;
    124: op1_00_in19 = reg_0897;
    126: op1_00_in19 = reg_0783;
    128: op1_00_in19 = reg_0027;
    129: op1_00_in19 = reg_0603;
    130: op1_00_in19 = reg_0489;
    131: op1_00_in19 = reg_0575;
    default: op1_00_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    35: op1_00_inv19 = 1;
    41: op1_00_inv19 = 1;
    38: op1_00_inv19 = 1;
    52: op1_00_inv19 = 1;
    58: op1_00_inv19 = 1;
    61: op1_00_inv19 = 1;
    67: op1_00_inv19 = 1;
    76: op1_00_inv19 = 1;
    68: op1_00_inv19 = 1;
    74: op1_00_inv19 = 1;
    73: op1_00_inv19 = 1;
    50: op1_00_inv19 = 1;
    86: op1_00_inv19 = 1;
    36: op1_00_inv19 = 1;
    47: op1_00_inv19 = 1;
    56: op1_00_inv19 = 1;
    75: op1_00_inv19 = 1;
    57: op1_00_inv19 = 1;
    79: op1_00_inv19 = 1;
    62: op1_00_inv19 = 1;
    83: op1_00_inv19 = 1;
    64: op1_00_inv19 = 1;
    84: op1_00_inv19 = 1;
    90: op1_00_inv19 = 1;
    85: op1_00_inv19 = 1;
    66: op1_00_inv19 = 1;
    93: op1_00_inv19 = 1;
    95: op1_00_inv19 = 1;
    96: op1_00_inv19 = 1;
    97: op1_00_inv19 = 1;
    99: op1_00_inv19 = 1;
    101: op1_00_inv19 = 1;
    102: op1_00_inv19 = 1;
    105: op1_00_inv19 = 1;
    107: op1_00_inv19 = 1;
    108: op1_00_inv19 = 1;
    109: op1_00_inv19 = 1;
    110: op1_00_inv19 = 1;
    113: op1_00_inv19 = 1;
    115: op1_00_inv19 = 1;
    116: op1_00_inv19 = 1;
    117: op1_00_inv19 = 1;
    120: op1_00_inv19 = 1;
    122: op1_00_inv19 = 1;
    126: op1_00_inv19 = 1;
    128: op1_00_inv19 = 1;
    129: op1_00_inv19 = 1;
    130: op1_00_inv19 = 1;
    default: op1_00_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の20番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in20 = reg_0071;
    15: op1_00_in20 = reg_0184;
    19: op1_00_in20 = reg_0049;
    11: op1_00_in20 = reg_0038;
    33: op1_00_in20 = reg_0468;
    35: op1_00_in20 = reg_0154;
    64: op1_00_in20 = reg_0154;
    105: op1_00_in20 = reg_0154;
    32: op1_00_in20 = reg_0199;
    26: op1_00_in20 = reg_0155;
    41: op1_00_in20 = imem01_in[3:0];
    38: op1_00_in20 = reg_0479;
    86: op1_00_in20 = reg_0479;
    39: op1_00_in20 = reg_0489;
    45: op1_00_in20 = reg_0269;
    52: op1_00_in20 = reg_0966;
    49: op1_00_in20 = reg_0450;
    46: op1_00_in20 = reg_0593;
    58: op1_00_in20 = reg_0747;
    54: op1_00_in20 = reg_0999;
    69: op1_00_in20 = reg_0999;
    48: op1_00_in20 = reg_0051;
    60: op1_00_in20 = reg_0984;
    53: op1_00_in20 = reg_0839;
    42: op1_00_in20 = reg_0839;
    61: op1_00_in20 = imem05_in[11:8];
    67: op1_00_in20 = reg_0526;
    76: op1_00_in20 = reg_1100;
    71: op1_00_in20 = reg_1164;
    72: op1_00_in20 = reg_0289;
    55: op1_00_in20 = reg_0706;
    68: op1_00_in20 = reg_0395;
    74: op1_00_in20 = reg_0185;
    87: op1_00_in20 = reg_0633;
    78: op1_00_in20 = reg_0373;
    73: op1_00_in20 = reg_0084;
    59: op1_00_in20 = reg_0728;
    50: op1_00_in20 = reg_0381;
    36: op1_00_in20 = reg_0381;
    44: op1_00_in20 = reg_0396;
    88: op1_00_in20 = imem03_in[3:0];
    47: op1_00_in20 = reg_0003;
    56: op1_00_in20 = reg_0032;
    75: op1_00_in20 = reg_0801;
    70: op1_00_in20 = reg_0377;
    57: op1_00_in20 = reg_0548;
    77: op1_00_in20 = reg_0303;
    51: op1_00_in20 = reg_0394;
    79: op1_00_in20 = reg_1512;
    43: op1_00_in20 = reg_0195;
    62: op1_00_in20 = reg_0634;
    80: op1_00_in20 = reg_0143;
    126: op1_00_in20 = reg_0143;
    81: op1_00_in20 = reg_0166;
    89: op1_00_in20 = reg_1147;
    63: op1_00_in20 = reg_0186;
    82: op1_00_in20 = reg_0978;
    83: op1_00_in20 = reg_0547;
    84: op1_00_in20 = reg_1183;
    65: op1_00_in20 = reg_0360;
    90: op1_00_in20 = reg_1107;
    85: op1_00_in20 = reg_0699;
    66: op1_00_in20 = reg_0119;
    91: op1_00_in20 = reg_1417;
    92: op1_00_in20 = reg_1420;
    93: op1_00_in20 = reg_1258;
    94: op1_00_in20 = reg_0967;
    112: op1_00_in20 = reg_0967;
    95: op1_00_in20 = reg_0172;
    96: op1_00_in20 = reg_1451;
    97: op1_00_in20 = reg_0008;
    99: op1_00_in20 = reg_1505;
    100: op1_00_in20 = reg_0968;
    101: op1_00_in20 = reg_0441;
    102: op1_00_in20 = reg_0789;
    103: op1_00_in20 = reg_0527;
    106: op1_00_in20 = reg_0382;
    107: op1_00_in20 = reg_1040;
    108: op1_00_in20 = reg_1323;
    109: op1_00_in20 = reg_0178;
    110: op1_00_in20 = reg_0122;
    111: op1_00_in20 = reg_0420;
    123: op1_00_in20 = reg_0420;
    113: op1_00_in20 = reg_0204;
    114: op1_00_in20 = reg_0217;
    115: op1_00_in20 = reg_0030;
    116: op1_00_in20 = reg_0060;
    117: op1_00_in20 = reg_0667;
    120: op1_00_in20 = reg_0496;
    121: op1_00_in20 = reg_0268;
    122: op1_00_in20 = reg_0717;
    124: op1_00_in20 = reg_1098;
    128: op1_00_in20 = imem01_in[15:12];
    129: op1_00_in20 = reg_0565;
    130: op1_00_in20 = reg_0777;
    131: op1_00_in20 = reg_0344;
    default: op1_00_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv20 = 1;
    15: op1_00_inv20 = 1;
    11: op1_00_inv20 = 1;
    32: op1_00_inv20 = 1;
    41: op1_00_inv20 = 1;
    38: op1_00_inv20 = 1;
    39: op1_00_inv20 = 1;
    49: op1_00_inv20 = 1;
    54: op1_00_inv20 = 1;
    48: op1_00_inv20 = 1;
    60: op1_00_inv20 = 1;
    76: op1_00_inv20 = 1;
    72: op1_00_inv20 = 1;
    55: op1_00_inv20 = 1;
    68: op1_00_inv20 = 1;
    78: op1_00_inv20 = 1;
    73: op1_00_inv20 = 1;
    86: op1_00_inv20 = 1;
    69: op1_00_inv20 = 1;
    75: op1_00_inv20 = 1;
    42: op1_00_inv20 = 1;
    51: op1_00_inv20 = 1;
    79: op1_00_inv20 = 1;
    43: op1_00_inv20 = 1;
    80: op1_00_inv20 = 1;
    81: op1_00_inv20 = 1;
    89: op1_00_inv20 = 1;
    84: op1_00_inv20 = 1;
    65: op1_00_inv20 = 1;
    85: op1_00_inv20 = 1;
    91: op1_00_inv20 = 1;
    94: op1_00_inv20 = 1;
    97: op1_00_inv20 = 1;
    101: op1_00_inv20 = 1;
    103: op1_00_inv20 = 1;
    105: op1_00_inv20 = 1;
    106: op1_00_inv20 = 1;
    107: op1_00_inv20 = 1;
    111: op1_00_inv20 = 1;
    114: op1_00_inv20 = 1;
    115: op1_00_inv20 = 1;
    116: op1_00_inv20 = 1;
    117: op1_00_inv20 = 1;
    122: op1_00_inv20 = 1;
    123: op1_00_inv20 = 1;
    124: op1_00_inv20 = 1;
    126: op1_00_inv20 = 1;
    128: op1_00_inv20 = 1;
    129: op1_00_inv20 = 1;
    130: op1_00_inv20 = 1;
    default: op1_00_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の21番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in21 = reg_0075;
    15: op1_00_in21 = reg_0168;
    68: op1_00_in21 = reg_0168;
    19: op1_00_in21 = reg_0025;
    84: op1_00_in21 = reg_0025;
    11: op1_00_in21 = reg_0014;
    33: op1_00_in21 = reg_0469;
    35: op1_00_in21 = reg_0325;
    32: op1_00_in21 = reg_0337;
    26: op1_00_in21 = reg_0171;
    41: op1_00_in21 = reg_0448;
    38: op1_00_in21 = reg_0448;
    39: op1_00_in21 = reg_0477;
    45: op1_00_in21 = reg_0046;
    52: op1_00_in21 = reg_0930;
    79: op1_00_in21 = reg_0930;
    49: op1_00_in21 = reg_0895;
    46: op1_00_in21 = reg_0050;
    58: op1_00_in21 = reg_0161;
    60: op1_00_in21 = reg_0161;
    54: op1_00_in21 = reg_0962;
    48: op1_00_in21 = reg_0001;
    53: op1_00_in21 = reg_0217;
    64: op1_00_in21 = reg_0217;
    61: op1_00_in21 = reg_0204;
    67: op1_00_in21 = reg_0979;
    76: op1_00_in21 = imem01_in[11:8];
    110: op1_00_in21 = imem01_in[11:8];
    71: op1_00_in21 = reg_0333;
    72: op1_00_in21 = reg_0269;
    55: op1_00_in21 = reg_0348;
    74: op1_00_in21 = reg_0144;
    87: op1_00_in21 = reg_0210;
    78: op1_00_in21 = reg_0570;
    59: op1_00_in21 = reg_0726;
    100: op1_00_in21 = reg_0726;
    50: op1_00_in21 = reg_0138;
    86: op1_00_in21 = imem03_in[11:8];
    69: op1_00_in21 = reg_1314;
    36: op1_00_in21 = reg_0342;
    44: op1_00_in21 = reg_0860;
    88: op1_00_in21 = imem03_in[15:12];
    47: op1_00_in21 = reg_0053;
    56: op1_00_in21 = reg_0793;
    75: op1_00_in21 = reg_0281;
    42: op1_00_in21 = reg_0830;
    70: op1_00_in21 = reg_0177;
    57: op1_00_in21 = reg_0239;
    77: op1_00_in21 = reg_0301;
    51: op1_00_in21 = imem07_in[7:4];
    43: op1_00_in21 = reg_0729;
    62: op1_00_in21 = reg_0548;
    80: op1_00_in21 = reg_0180;
    126: op1_00_in21 = reg_0180;
    81: op1_00_in21 = reg_1513;
    89: op1_00_in21 = reg_1065;
    107: op1_00_in21 = reg_1065;
    63: op1_00_in21 = reg_1315;
    82: op1_00_in21 = reg_0462;
    83: op1_00_in21 = reg_0609;
    65: op1_00_in21 = reg_0875;
    90: op1_00_in21 = reg_0021;
    85: op1_00_in21 = reg_0759;
    66: op1_00_in21 = reg_1204;
    91: op1_00_in21 = reg_0459;
    92: op1_00_in21 = reg_0133;
    93: op1_00_in21 = reg_0531;
    94: op1_00_in21 = reg_0383;
    112: op1_00_in21 = reg_0383;
    95: op1_00_in21 = reg_0780;
    96: op1_00_in21 = reg_0128;
    97: op1_00_in21 = reg_0069;
    99: op1_00_in21 = reg_1303;
    101: op1_00_in21 = reg_0366;
    102: op1_00_in21 = reg_0375;
    103: op1_00_in21 = reg_0568;
    105: op1_00_in21 = reg_1448;
    106: op1_00_in21 = reg_0496;
    108: op1_00_in21 = reg_1505;
    109: op1_00_in21 = reg_1009;
    111: op1_00_in21 = reg_0019;
    113: op1_00_in21 = reg_0338;
    114: op1_00_in21 = reg_0255;
    115: op1_00_in21 = reg_0741;
    116: op1_00_in21 = reg_0059;
    117: op1_00_in21 = reg_0922;
    120: op1_00_in21 = reg_1433;
    121: op1_00_in21 = reg_0862;
    122: op1_00_in21 = reg_0398;
    123: op1_00_in21 = reg_1488;
    124: op1_00_in21 = reg_0711;
    128: op1_00_in21 = reg_0576;
    129: op1_00_in21 = imem06_in[3:0];
    130: op1_00_in21 = reg_0030;
    131: op1_00_in21 = reg_0449;
    default: op1_00_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    19: op1_00_inv21 = 1;
    11: op1_00_inv21 = 1;
    32: op1_00_inv21 = 1;
    26: op1_00_inv21 = 1;
    41: op1_00_inv21 = 1;
    39: op1_00_inv21 = 1;
    45: op1_00_inv21 = 1;
    52: op1_00_inv21 = 1;
    49: op1_00_inv21 = 1;
    58: op1_00_inv21 = 1;
    48: op1_00_inv21 = 1;
    60: op1_00_inv21 = 1;
    68: op1_00_inv21 = 1;
    74: op1_00_inv21 = 1;
    78: op1_00_inv21 = 1;
    50: op1_00_inv21 = 1;
    88: op1_00_inv21 = 1;
    47: op1_00_inv21 = 1;
    56: op1_00_inv21 = 1;
    42: op1_00_inv21 = 1;
    70: op1_00_inv21 = 1;
    57: op1_00_inv21 = 1;
    77: op1_00_inv21 = 1;
    81: op1_00_inv21 = 1;
    63: op1_00_inv21 = 1;
    83: op1_00_inv21 = 1;
    84: op1_00_inv21 = 1;
    65: op1_00_inv21 = 1;
    90: op1_00_inv21 = 1;
    66: op1_00_inv21 = 1;
    92: op1_00_inv21 = 1;
    94: op1_00_inv21 = 1;
    95: op1_00_inv21 = 1;
    99: op1_00_inv21 = 1;
    100: op1_00_inv21 = 1;
    102: op1_00_inv21 = 1;
    106: op1_00_inv21 = 1;
    107: op1_00_inv21 = 1;
    115: op1_00_inv21 = 1;
    116: op1_00_inv21 = 1;
    124: op1_00_inv21 = 1;
    128: op1_00_inv21 = 1;
    130: op1_00_inv21 = 1;
    default: op1_00_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の22番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in22 = reg_0057;
    15: op1_00_in22 = reg_0169;
    19: op1_00_in22 = reg_0000;
    11: op1_00_in22 = imem06_in[3:0];
    33: op1_00_in22 = reg_0446;
    35: op1_00_in22 = reg_0069;
    32: op1_00_in22 = reg_0164;
    26: op1_00_in22 = reg_0172;
    108: op1_00_in22 = reg_0172;
    41: op1_00_in22 = reg_0819;
    38: op1_00_in22 = reg_0328;
    39: op1_00_in22 = reg_0449;
    45: op1_00_in22 = imem07_in[3:0];
    52: op1_00_in22 = reg_0092;
    49: op1_00_in22 = reg_0872;
    46: op1_00_in22 = reg_0052;
    58: op1_00_in22 = reg_0553;
    54: op1_00_in22 = reg_0952;
    48: op1_00_in22 = reg_0002;
    60: op1_00_in22 = reg_0967;
    53: op1_00_in22 = reg_0311;
    61: op1_00_in22 = reg_0702;
    67: op1_00_in22 = reg_1225;
    76: op1_00_in22 = reg_1512;
    71: op1_00_in22 = reg_0566;
    72: op1_00_in22 = reg_0215;
    55: op1_00_in22 = reg_0232;
    68: op1_00_in22 = reg_1164;
    74: op1_00_in22 = reg_0789;
    87: op1_00_in22 = reg_0370;
    78: op1_00_in22 = reg_0522;
    59: op1_00_in22 = reg_0403;
    50: op1_00_in22 = reg_0154;
    86: op1_00_in22 = reg_1280;
    69: op1_00_in22 = reg_0954;
    36: op1_00_in22 = reg_0054;
    44: op1_00_in22 = reg_0371;
    88: op1_00_in22 = reg_1000;
    47: op1_00_in22 = reg_0085;
    56: op1_00_in22 = reg_0631;
    75: op1_00_in22 = imem02_in[3:0];
    42: op1_00_in22 = reg_0068;
    70: op1_00_in22 = reg_0199;
    57: op1_00_in22 = reg_0161;
    77: op1_00_in22 = reg_0090;
    51: op1_00_in22 = reg_0299;
    79: op1_00_in22 = reg_0258;
    128: op1_00_in22 = reg_0258;
    43: op1_00_in22 = reg_0860;
    92: op1_00_in22 = reg_0860;
    62: op1_00_in22 = reg_0746;
    80: op1_00_in22 = reg_0989;
    81: op1_00_in22 = reg_0331;
    89: op1_00_in22 = reg_0342;
    63: op1_00_in22 = reg_0894;
    82: op1_00_in22 = reg_0577;
    83: op1_00_in22 = reg_0238;
    64: op1_00_in22 = reg_0227;
    84: op1_00_in22 = reg_0245;
    65: op1_00_in22 = reg_0292;
    90: op1_00_in22 = reg_0210;
    111: op1_00_in22 = reg_0210;
    85: op1_00_in22 = reg_0179;
    66: op1_00_in22 = reg_0185;
    91: op1_00_in22 = reg_1405;
    93: op1_00_in22 = reg_0574;
    94: op1_00_in22 = reg_0360;
    95: op1_00_in22 = reg_0116;
    96: op1_00_in22 = reg_0112;
    97: op1_00_in22 = imem03_in[11:8];
    99: op1_00_in22 = reg_0398;
    100: op1_00_in22 = reg_0146;
    101: op1_00_in22 = reg_0623;
    102: op1_00_in22 = reg_1494;
    103: op1_00_in22 = reg_0571;
    105: op1_00_in22 = reg_0216;
    106: op1_00_in22 = reg_1433;
    107: op1_00_in22 = reg_0320;
    109: op1_00_in22 = reg_0313;
    110: op1_00_in22 = reg_0166;
    112: op1_00_in22 = reg_0362;
    113: op1_00_in22 = reg_0346;
    114: op1_00_in22 = imem03_in[7:4];
    115: op1_00_in22 = reg_0591;
    116: op1_00_in22 = reg_0723;
    117: op1_00_in22 = reg_0310;
    120: op1_00_in22 = reg_0876;
    121: op1_00_in22 = reg_0719;
    122: op1_00_in22 = reg_0586;
    123: op1_00_in22 = imem05_in[7:4];
    124: op1_00_in22 = reg_0848;
    126: op1_00_in22 = reg_0142;
    129: op1_00_in22 = imem06_in[11:8];
    130: op1_00_in22 = reg_0287;
    131: op1_00_in22 = reg_0828;
    default: op1_00_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    19: op1_00_inv22 = 1;
    11: op1_00_inv22 = 1;
    38: op1_00_inv22 = 1;
    45: op1_00_inv22 = 1;
    52: op1_00_inv22 = 1;
    58: op1_00_inv22 = 1;
    54: op1_00_inv22 = 1;
    61: op1_00_inv22 = 1;
    76: op1_00_inv22 = 1;
    71: op1_00_inv22 = 1;
    72: op1_00_inv22 = 1;
    55: op1_00_inv22 = 1;
    87: op1_00_inv22 = 1;
    59: op1_00_inv22 = 1;
    50: op1_00_inv22 = 1;
    86: op1_00_inv22 = 1;
    36: op1_00_inv22 = 1;
    44: op1_00_inv22 = 1;
    88: op1_00_inv22 = 1;
    56: op1_00_inv22 = 1;
    75: op1_00_inv22 = 1;
    57: op1_00_inv22 = 1;
    79: op1_00_inv22 = 1;
    62: op1_00_inv22 = 1;
    89: op1_00_inv22 = 1;
    83: op1_00_inv22 = 1;
    90: op1_00_inv22 = 1;
    66: op1_00_inv22 = 1;
    91: op1_00_inv22 = 1;
    93: op1_00_inv22 = 1;
    97: op1_00_inv22 = 1;
    107: op1_00_inv22 = 1;
    108: op1_00_inv22 = 1;
    109: op1_00_inv22 = 1;
    112: op1_00_inv22 = 1;
    115: op1_00_inv22 = 1;
    120: op1_00_inv22 = 1;
    121: op1_00_inv22 = 1;
    122: op1_00_inv22 = 1;
    123: op1_00_inv22 = 1;
    124: op1_00_inv22 = 1;
    126: op1_00_inv22 = 1;
    129: op1_00_inv22 = 1;
    default: op1_00_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の23番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in23 = reg_0026;
    15: op1_00_in23 = reg_0153;
    19: op1_00_in23 = imem04_in[7:4];
    11: op1_00_in23 = reg_0165;
    33: op1_00_in23 = reg_0430;
    60: op1_00_in23 = reg_0430;
    35: op1_00_in23 = reg_0276;
    32: op1_00_in23 = reg_0117;
    26: op1_00_in23 = reg_0263;
    41: op1_00_in23 = reg_0787;
    38: op1_00_in23 = reg_0329;
    39: op1_00_in23 = reg_0130;
    45: op1_00_in23 = reg_0135;
    52: op1_00_in23 = reg_0724;
    49: op1_00_in23 = reg_0449;
    46: op1_00_in23 = reg_0519;
    48: op1_00_in23 = reg_0519;
    58: op1_00_in23 = reg_0967;
    54: op1_00_in23 = reg_0558;
    53: op1_00_in23 = reg_0312;
    61: op1_00_in23 = reg_0395;
    67: op1_00_in23 = reg_1202;
    76: op1_00_in23 = reg_0331;
    71: op1_00_in23 = reg_0045;
    72: op1_00_in23 = reg_1170;
    55: op1_00_in23 = reg_0790;
    68: op1_00_in23 = reg_0996;
    74: op1_00_in23 = reg_0142;
    87: op1_00_in23 = imem05_in[11:8];
    123: op1_00_in23 = imem05_in[11:8];
    78: op1_00_in23 = reg_0296;
    59: op1_00_in23 = reg_0386;
    50: op1_00_in23 = reg_0830;
    83: op1_00_in23 = reg_0830;
    86: op1_00_in23 = reg_0427;
    69: op1_00_in23 = reg_0246;
    36: op1_00_in23 = imem02_in[11:8];
    44: op1_00_in23 = reg_0109;
    88: op1_00_in23 = reg_0185;
    47: op1_00_in23 = reg_0520;
    56: op1_00_in23 = reg_0175;
    94: op1_00_in23 = reg_0175;
    75: op1_00_in23 = reg_1000;
    42: op1_00_in23 = reg_0069;
    70: op1_00_in23 = reg_0375;
    57: op1_00_in23 = reg_0609;
    77: op1_00_in23 = reg_1484;
    51: op1_00_in23 = reg_0309;
    79: op1_00_in23 = reg_0547;
    43: op1_00_in23 = reg_0859;
    62: op1_00_in23 = reg_0747;
    80: op1_00_in23 = reg_0377;
    81: op1_00_in23 = reg_0222;
    89: op1_00_in23 = reg_0582;
    63: op1_00_in23 = reg_0703;
    84: op1_00_in23 = reg_0703;
    82: op1_00_in23 = reg_1215;
    64: op1_00_in23 = reg_1063;
    65: op1_00_in23 = reg_0044;
    90: op1_00_in23 = imem05_in[7:4];
    85: op1_00_in23 = reg_1449;
    66: op1_00_in23 = imem07_in[3:0];
    91: op1_00_in23 = reg_0476;
    92: op1_00_in23 = reg_1323;
    93: op1_00_in23 = reg_1233;
    95: op1_00_in23 = reg_0527;
    96: op1_00_in23 = reg_0897;
    97: op1_00_in23 = reg_0504;
    99: op1_00_in23 = reg_0586;
    100: op1_00_in23 = reg_0290;
    101: op1_00_in23 = reg_0137;
    102: op1_00_in23 = reg_0070;
    103: op1_00_in23 = reg_1225;
    105: op1_00_in23 = reg_0198;
    106: op1_00_in23 = reg_0473;
    107: op1_00_in23 = reg_0061;
    108: op1_00_in23 = reg_1179;
    109: op1_00_in23 = reg_0288;
    110: op1_00_in23 = reg_0010;
    111: op1_00_in23 = reg_0470;
    112: op1_00_in23 = reg_0092;
    113: op1_00_in23 = reg_0831;
    114: op1_00_in23 = imem03_in[15:12];
    115: op1_00_in23 = reg_0103;
    116: op1_00_in23 = imem01_in[3:0];
    117: op1_00_in23 = reg_0786;
    120: op1_00_in23 = reg_0381;
    121: op1_00_in23 = reg_0211;
    122: op1_00_in23 = reg_0570;
    124: op1_00_in23 = reg_1006;
    126: op1_00_in23 = reg_0349;
    128: op1_00_in23 = reg_0549;
    129: op1_00_in23 = imem06_in[15:12];
    130: op1_00_in23 = reg_0441;
    131: op1_00_in23 = reg_1431;
    default: op1_00_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_00_inv23 = 1;
    19: op1_00_inv23 = 1;
    11: op1_00_inv23 = 1;
    33: op1_00_inv23 = 1;
    32: op1_00_inv23 = 1;
    41: op1_00_inv23 = 1;
    38: op1_00_inv23 = 1;
    39: op1_00_inv23 = 1;
    58: op1_00_inv23 = 1;
    54: op1_00_inv23 = 1;
    48: op1_00_inv23 = 1;
    60: op1_00_inv23 = 1;
    53: op1_00_inv23 = 1;
    67: op1_00_inv23 = 1;
    76: op1_00_inv23 = 1;
    74: op1_00_inv23 = 1;
    87: op1_00_inv23 = 1;
    50: op1_00_inv23 = 1;
    86: op1_00_inv23 = 1;
    69: op1_00_inv23 = 1;
    88: op1_00_inv23 = 1;
    47: op1_00_inv23 = 1;
    42: op1_00_inv23 = 1;
    57: op1_00_inv23 = 1;
    51: op1_00_inv23 = 1;
    43: op1_00_inv23 = 1;
    81: op1_00_inv23 = 1;
    89: op1_00_inv23 = 1;
    82: op1_00_inv23 = 1;
    83: op1_00_inv23 = 1;
    64: op1_00_inv23 = 1;
    84: op1_00_inv23 = 1;
    65: op1_00_inv23 = 1;
    93: op1_00_inv23 = 1;
    95: op1_00_inv23 = 1;
    97: op1_00_inv23 = 1;
    99: op1_00_inv23 = 1;
    100: op1_00_inv23 = 1;
    105: op1_00_inv23 = 1;
    106: op1_00_inv23 = 1;
    107: op1_00_inv23 = 1;
    108: op1_00_inv23 = 1;
    110: op1_00_inv23 = 1;
    112: op1_00_inv23 = 1;
    113: op1_00_inv23 = 1;
    116: op1_00_inv23 = 1;
    120: op1_00_inv23 = 1;
    124: op1_00_inv23 = 1;
    126: op1_00_inv23 = 1;
    129: op1_00_inv23 = 1;
    131: op1_00_inv23 = 1;
    default: op1_00_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の24番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in24 = reg_0027;
    15: op1_00_in24 = reg_0133;
    19: op1_00_in24 = imem04_in[11:8];
    11: op1_00_in24 = reg_0152;
    33: op1_00_in24 = reg_0401;
    35: op1_00_in24 = imem03_in[11:8];
    32: op1_00_in24 = reg_0065;
    26: op1_00_in24 = reg_0323;
    41: op1_00_in24 = reg_0742;
    38: op1_00_in24 = imem04_in[7:4];
    39: op1_00_in24 = reg_0240;
    45: op1_00_in24 = reg_0892;
    52: op1_00_in24 = reg_0899;
    49: op1_00_in24 = imem06_in[3:0];
    46: op1_00_in24 = reg_0521;
    58: op1_00_in24 = reg_0819;
    54: op1_00_in24 = reg_0113;
    48: op1_00_in24 = reg_0520;
    60: op1_00_in24 = reg_0728;
    53: op1_00_in24 = reg_0709;
    61: op1_00_in24 = reg_0347;
    67: op1_00_in24 = reg_0269;
    76: op1_00_in24 = reg_0258;
    71: op1_00_in24 = reg_1181;
    72: op1_00_in24 = imem07_in[3:0];
    55: op1_00_in24 = reg_0789;
    68: op1_00_in24 = reg_0392;
    113: op1_00_in24 = reg_0392;
    74: op1_00_in24 = reg_0965;
    87: op1_00_in24 = reg_0278;
    78: op1_00_in24 = reg_0289;
    59: op1_00_in24 = reg_0385;
    50: op1_00_in24 = reg_0829;
    120: op1_00_in24 = reg_0829;
    86: op1_00_in24 = reg_1384;
    69: op1_00_in24 = reg_0558;
    36: op1_00_in24 = reg_0009;
    44: op1_00_in24 = reg_0636;
    43: op1_00_in24 = reg_0636;
    88: op1_00_in24 = reg_1449;
    47: op1_00_in24 = reg_0123;
    56: op1_00_in24 = reg_0831;
    75: op1_00_in24 = reg_0559;
    114: op1_00_in24 = reg_0559;
    42: op1_00_in24 = reg_0325;
    70: op1_00_in24 = reg_0376;
    57: op1_00_in24 = reg_1152;
    77: op1_00_in24 = reg_0602;
    51: op1_00_in24 = reg_0673;
    79: op1_00_in24 = reg_0746;
    62: op1_00_in24 = imem01_in[7:4];
    80: op1_00_in24 = reg_0070;
    81: op1_00_in24 = reg_0260;
    89: op1_00_in24 = reg_0262;
    63: op1_00_in24 = reg_0140;
    84: op1_00_in24 = reg_0140;
    82: op1_00_in24 = reg_1216;
    83: op1_00_in24 = reg_0612;
    64: op1_00_in24 = reg_0350;
    65: op1_00_in24 = reg_0013;
    90: op1_00_in24 = imem05_in[15:12];
    85: op1_00_in24 = reg_0177;
    66: op1_00_in24 = reg_0310;
    91: op1_00_in24 = reg_0351;
    92: op1_00_in24 = reg_0827;
    93: op1_00_in24 = reg_0500;
    94: op1_00_in24 = reg_0464;
    95: op1_00_in24 = reg_0569;
    96: op1_00_in24 = reg_0007;
    97: op1_00_in24 = reg_0507;
    99: op1_00_in24 = reg_0617;
    100: op1_00_in24 = reg_1511;
    101: op1_00_in24 = reg_0100;
    102: op1_00_in24 = reg_1516;
    103: op1_00_in24 = reg_0419;
    105: op1_00_in24 = reg_0847;
    106: op1_00_in24 = reg_0306;
    107: op1_00_in24 = reg_0368;
    108: op1_00_in24 = reg_0265;
    109: op1_00_in24 = reg_0426;
    110: op1_00_in24 = reg_0985;
    111: op1_00_in24 = imem05_in[11:8];
    112: op1_00_in24 = reg_0901;
    115: op1_00_in24 = reg_0085;
    116: op1_00_in24 = reg_0980;
    117: op1_00_in24 = reg_0457;
    121: op1_00_in24 = reg_1107;
    122: op1_00_in24 = reg_0296;
    123: op1_00_in24 = reg_1259;
    124: op1_00_in24 = reg_0227;
    126: op1_00_in24 = reg_0954;
    128: op1_00_in24 = reg_0241;
    129: op1_00_in24 = reg_0670;
    130: op1_00_in24 = reg_0437;
    131: op1_00_in24 = reg_0039;
    default: op1_00_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_00_inv24 = 1;
    32: op1_00_inv24 = 1;
    26: op1_00_inv24 = 1;
    41: op1_00_inv24 = 1;
    46: op1_00_inv24 = 1;
    58: op1_00_inv24 = 1;
    48: op1_00_inv24 = 1;
    60: op1_00_inv24 = 1;
    67: op1_00_inv24 = 1;
    76: op1_00_inv24 = 1;
    72: op1_00_inv24 = 1;
    87: op1_00_inv24 = 1;
    50: op1_00_inv24 = 1;
    86: op1_00_inv24 = 1;
    69: op1_00_inv24 = 1;
    36: op1_00_inv24 = 1;
    88: op1_00_inv24 = 1;
    42: op1_00_inv24 = 1;
    70: op1_00_inv24 = 1;
    57: op1_00_inv24 = 1;
    77: op1_00_inv24 = 1;
    79: op1_00_inv24 = 1;
    43: op1_00_inv24 = 1;
    62: op1_00_inv24 = 1;
    81: op1_00_inv24 = 1;
    89: op1_00_inv24 = 1;
    63: op1_00_inv24 = 1;
    83: op1_00_inv24 = 1;
    64: op1_00_inv24 = 1;
    91: op1_00_inv24 = 1;
    92: op1_00_inv24 = 1;
    93: op1_00_inv24 = 1;
    95: op1_00_inv24 = 1;
    96: op1_00_inv24 = 1;
    97: op1_00_inv24 = 1;
    99: op1_00_inv24 = 1;
    100: op1_00_inv24 = 1;
    102: op1_00_inv24 = 1;
    103: op1_00_inv24 = 1;
    107: op1_00_inv24 = 1;
    109: op1_00_inv24 = 1;
    112: op1_00_inv24 = 1;
    113: op1_00_inv24 = 1;
    115: op1_00_inv24 = 1;
    116: op1_00_inv24 = 1;
    117: op1_00_inv24 = 1;
    121: op1_00_inv24 = 1;
    122: op1_00_inv24 = 1;
    123: op1_00_inv24 = 1;
    124: op1_00_inv24 = 1;
    128: op1_00_inv24 = 1;
    129: op1_00_inv24 = 1;
    default: op1_00_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の25番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in25 = reg_0005;
    15: op1_00_in25 = reg_0126;
    19: op1_00_in25 = reg_0292;
    11: op1_00_in25 = reg_0132;
    33: op1_00_in25 = reg_0386;
    35: op1_00_in25 = reg_0632;
    32: op1_00_in25 = reg_0211;
    26: op1_00_in25 = reg_0308;
    41: op1_00_in25 = reg_0724;
    38: op1_00_in25 = reg_0721;
    39: op1_00_in25 = reg_0274;
    45: op1_00_in25 = reg_0187;
    52: op1_00_in25 = reg_0875;
    49: op1_00_in25 = imem06_in[7:4];
    46: op1_00_in25 = reg_0124;
    58: op1_00_in25 = reg_0439;
    54: op1_00_in25 = reg_0885;
    60: op1_00_in25 = reg_0400;
    53: op1_00_in25 = reg_1063;
    114: op1_00_in25 = reg_1063;
    61: op1_00_in25 = reg_0700;
    67: op1_00_in25 = reg_1170;
    76: op1_00_in25 = reg_0222;
    65: op1_00_in25 = reg_0222;
    71: op1_00_in25 = reg_1401;
    72: op1_00_in25 = reg_0065;
    55: op1_00_in25 = reg_1003;
    68: op1_00_in25 = reg_0565;
    74: op1_00_in25 = reg_0964;
    87: op1_00_in25 = reg_0733;
    78: op1_00_in25 = reg_0119;
    59: op1_00_in25 = reg_0362;
    50: op1_00_in25 = reg_0800;
    86: op1_00_in25 = reg_1383;
    69: op1_00_in25 = reg_1199;
    36: op1_00_in25 = reg_0326;
    44: op1_00_in25 = reg_0637;
    88: op1_00_in25 = reg_1001;
    56: op1_00_in25 = reg_0701;
    75: op1_00_in25 = reg_0227;
    42: op1_00_in25 = reg_0276;
    70: op1_00_in25 = reg_0180;
    57: op1_00_in25 = reg_0469;
    77: op1_00_in25 = reg_1346;
    51: op1_00_in25 = reg_0159;
    79: op1_00_in25 = reg_0743;
    62: op1_00_in25 = reg_0743;
    43: op1_00_in25 = reg_0263;
    80: op1_00_in25 = reg_0349;
    81: op1_00_in25 = reg_0798;
    89: op1_00_in25 = reg_0337;
    107: op1_00_in25 = reg_0337;
    63: op1_00_in25 = reg_0157;
    82: op1_00_in25 = imem04_in[15:12];
    109: op1_00_in25 = imem04_in[15:12];
    83: op1_00_in25 = reg_0438;
    64: op1_00_in25 = reg_0638;
    84: op1_00_in25 = reg_0170;
    90: op1_00_in25 = reg_0736;
    85: op1_00_in25 = reg_0216;
    66: op1_00_in25 = reg_0851;
    91: op1_00_in25 = reg_0075;
    92: op1_00_in25 = reg_0780;
    93: op1_00_in25 = reg_1147;
    94: op1_00_in25 = reg_0011;
    95: op1_00_in25 = reg_0570;
    96: op1_00_in25 = reg_0279;
    97: op1_00_in25 = reg_0999;
    99: op1_00_in25 = reg_0528;
    100: op1_00_in25 = reg_0385;
    101: op1_00_in25 = reg_0086;
    102: op1_00_in25 = reg_0314;
    103: op1_00_in25 = reg_0244;
    105: op1_00_in25 = reg_0789;
    106: op1_00_in25 = reg_0711;
    108: op1_00_in25 = reg_1508;
    110: op1_00_in25 = reg_0874;
    111: op1_00_in25 = reg_0466;
    112: op1_00_in25 = reg_0335;
    113: op1_00_in25 = reg_0566;
    116: op1_00_in25 = reg_0785;
    117: op1_00_in25 = reg_0139;
    120: op1_00_in25 = reg_0009;
    121: op1_00_in25 = reg_0021;
    122: op1_00_in25 = reg_0371;
    123: op1_00_in25 = reg_0832;
    124: op1_00_in25 = reg_0563;
    126: op1_00_in25 = reg_1092;
    128: op1_00_in25 = reg_0149;
    129: op1_00_in25 = reg_0397;
    130: op1_00_in25 = reg_0052;
    131: op1_00_in25 = imem06_in[3:0];
    default: op1_00_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv25 = 1;
    19: op1_00_inv25 = 1;
    11: op1_00_inv25 = 1;
    35: op1_00_inv25 = 1;
    26: op1_00_inv25 = 1;
    39: op1_00_inv25 = 1;
    45: op1_00_inv25 = 1;
    49: op1_00_inv25 = 1;
    54: op1_00_inv25 = 1;
    60: op1_00_inv25 = 1;
    67: op1_00_inv25 = 1;
    76: op1_00_inv25 = 1;
    71: op1_00_inv25 = 1;
    55: op1_00_inv25 = 1;
    68: op1_00_inv25 = 1;
    74: op1_00_inv25 = 1;
    87: op1_00_inv25 = 1;
    50: op1_00_inv25 = 1;
    56: op1_00_inv25 = 1;
    75: op1_00_inv25 = 1;
    42: op1_00_inv25 = 1;
    70: op1_00_inv25 = 1;
    57: op1_00_inv25 = 1;
    77: op1_00_inv25 = 1;
    51: op1_00_inv25 = 1;
    79: op1_00_inv25 = 1;
    43: op1_00_inv25 = 1;
    62: op1_00_inv25 = 1;
    81: op1_00_inv25 = 1;
    89: op1_00_inv25 = 1;
    63: op1_00_inv25 = 1;
    82: op1_00_inv25 = 1;
    83: op1_00_inv25 = 1;
    84: op1_00_inv25 = 1;
    65: op1_00_inv25 = 1;
    91: op1_00_inv25 = 1;
    93: op1_00_inv25 = 1;
    94: op1_00_inv25 = 1;
    95: op1_00_inv25 = 1;
    99: op1_00_inv25 = 1;
    100: op1_00_inv25 = 1;
    101: op1_00_inv25 = 1;
    103: op1_00_inv25 = 1;
    105: op1_00_inv25 = 1;
    108: op1_00_inv25 = 1;
    111: op1_00_inv25 = 1;
    112: op1_00_inv25 = 1;
    114: op1_00_inv25 = 1;
    121: op1_00_inv25 = 1;
    122: op1_00_inv25 = 1;
    123: op1_00_inv25 = 1;
    126: op1_00_inv25 = 1;
    128: op1_00_inv25 = 1;
    129: op1_00_inv25 = 1;
    130: op1_00_inv25 = 1;
    default: op1_00_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の26番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in26 = imem01_in[15:12];
    15: op1_00_in26 = reg_0106;
    19: op1_00_in26 = reg_0088;
    11: op1_00_in26 = reg_0119;
    33: op1_00_in26 = reg_0362;
    35: op1_00_in26 = reg_0600;
    32: op1_00_in26 = reg_0064;
    26: op1_00_in26 = reg_0295;
    41: op1_00_in26 = reg_0726;
    38: op1_00_in26 = reg_0719;
    39: op1_00_in26 = reg_0151;
    45: op1_00_in26 = reg_0851;
    84: op1_00_in26 = reg_0851;
    52: op1_00_in26 = reg_0078;
    49: op1_00_in26 = imem06_in[15:12];
    58: op1_00_in26 = reg_0147;
    54: op1_00_in26 = reg_0849;
    60: op1_00_in26 = reg_0384;
    53: op1_00_in26 = reg_0349;
    61: op1_00_in26 = reg_0066;
    67: op1_00_in26 = imem07_in[15:12];
    76: op1_00_in26 = reg_0798;
    71: op1_00_in26 = reg_0541;
    72: op1_00_in26 = reg_1439;
    55: op1_00_in26 = reg_0143;
    68: op1_00_in26 = reg_0745;
    74: op1_00_in26 = reg_0952;
    87: op1_00_in26 = reg_0174;
    78: op1_00_in26 = reg_0023;
    59: op1_00_in26 = reg_0360;
    50: op1_00_in26 = reg_0325;
    86: op1_00_in26 = reg_0032;
    69: op1_00_in26 = reg_1092;
    36: op1_00_in26 = reg_0276;
    44: op1_00_in26 = reg_0619;
    88: op1_00_in26 = reg_0707;
    56: op1_00_in26 = reg_0395;
    75: op1_00_in26 = reg_0706;
    42: op1_00_in26 = reg_0312;
    70: op1_00_in26 = reg_0965;
    57: op1_00_in26 = reg_0403;
    112: op1_00_in26 = reg_0403;
    77: op1_00_in26 = reg_0589;
    51: op1_00_in26 = reg_0156;
    79: op1_00_in26 = reg_0609;
    43: op1_00_in26 = reg_0132;
    62: op1_00_in26 = reg_0715;
    80: op1_00_in26 = reg_1231;
    81: op1_00_in26 = reg_0612;
    89: op1_00_in26 = reg_0339;
    63: op1_00_in26 = reg_0923;
    82: op1_00_in26 = reg_0407;
    83: op1_00_in26 = reg_0092;
    64: op1_00_in26 = reg_0999;
    65: op1_00_in26 = reg_0699;
    90: op1_00_in26 = reg_0579;
    85: op1_00_in26 = reg_0847;
    66: op1_00_in26 = reg_1349;
    91: op1_00_in26 = reg_0027;
    92: op1_00_in26 = reg_0110;
    93: op1_00_in26 = reg_0421;
    94: op1_00_in26 = imem02_in[15:12];
    95: op1_00_in26 = reg_1225;
    96: op1_00_in26 = imem03_in[11:8];
    97: op1_00_in26 = reg_0233;
    99: op1_00_in26 = reg_0571;
    100: op1_00_in26 = reg_0899;
    101: op1_00_in26 = reg_0518;
    102: op1_00_in26 = reg_0190;
    103: op1_00_in26 = reg_0754;
    105: op1_00_in26 = reg_1494;
    106: op1_00_in26 = reg_0008;
    107: op1_00_in26 = reg_0096;
    108: op1_00_in26 = reg_0637;
    109: op1_00_in26 = reg_0263;
    110: op1_00_in26 = reg_0576;
    111: op1_00_in26 = reg_0347;
    113: op1_00_in26 = reg_0131;
    114: op1_00_in26 = reg_0198;
    116: op1_00_in26 = reg_0282;
    117: op1_00_in26 = reg_0224;
    120: op1_00_in26 = reg_0227;
    121: op1_00_in26 = reg_1488;
    122: op1_00_in26 = reg_0015;
    123: op1_00_in26 = reg_0445;
    124: op1_00_in26 = imem03_in[3:0];
    126: op1_00_in26 = reg_0108;
    128: op1_00_in26 = reg_1034;
    129: op1_00_in26 = reg_0870;
    130: op1_00_in26 = reg_0086;
    131: op1_00_in26 = reg_0714;
    default: op1_00_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_00_inv26 = 1;
    35: op1_00_inv26 = 1;
    26: op1_00_inv26 = 1;
    38: op1_00_inv26 = 1;
    52: op1_00_inv26 = 1;
    54: op1_00_inv26 = 1;
    60: op1_00_inv26 = 1;
    61: op1_00_inv26 = 1;
    76: op1_00_inv26 = 1;
    71: op1_00_inv26 = 1;
    72: op1_00_inv26 = 1;
    55: op1_00_inv26 = 1;
    68: op1_00_inv26 = 1;
    86: op1_00_inv26 = 1;
    44: op1_00_inv26 = 1;
    88: op1_00_inv26 = 1;
    56: op1_00_inv26 = 1;
    75: op1_00_inv26 = 1;
    42: op1_00_inv26 = 1;
    70: op1_00_inv26 = 1;
    77: op1_00_inv26 = 1;
    62: op1_00_inv26 = 1;
    81: op1_00_inv26 = 1;
    63: op1_00_inv26 = 1;
    64: op1_00_inv26 = 1;
    90: op1_00_inv26 = 1;
    85: op1_00_inv26 = 1;
    66: op1_00_inv26 = 1;
    91: op1_00_inv26 = 1;
    92: op1_00_inv26 = 1;
    94: op1_00_inv26 = 1;
    97: op1_00_inv26 = 1;
    100: op1_00_inv26 = 1;
    102: op1_00_inv26 = 1;
    105: op1_00_inv26 = 1;
    106: op1_00_inv26 = 1;
    108: op1_00_inv26 = 1;
    109: op1_00_inv26 = 1;
    110: op1_00_inv26 = 1;
    111: op1_00_inv26 = 1;
    112: op1_00_inv26 = 1;
    113: op1_00_inv26 = 1;
    114: op1_00_inv26 = 1;
    117: op1_00_inv26 = 1;
    120: op1_00_inv26 = 1;
    126: op1_00_inv26 = 1;
    128: op1_00_inv26 = 1;
    129: op1_00_inv26 = 1;
    130: op1_00_inv26 = 1;
    default: op1_00_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の27番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in27 = reg_0307;
    15: op1_00_in27 = reg_0068;
    19: op1_00_in27 = reg_0262;
    11: op1_00_in27 = reg_0109;
    92: op1_00_in27 = reg_0109;
    33: op1_00_in27 = reg_0365;
    35: op1_00_in27 = reg_0573;
    32: op1_00_in27 = reg_0061;
    26: op1_00_in27 = reg_0119;
    41: op1_00_in27 = reg_0715;
    38: op1_00_in27 = reg_0695;
    39: op1_00_in27 = imem06_in[11:8];
    45: op1_00_in27 = reg_0158;
    66: op1_00_in27 = reg_0158;
    52: op1_00_in27 = reg_0282;
    49: op1_00_in27 = reg_0161;
    58: op1_00_in27 = reg_0402;
    54: op1_00_in27 = imem04_in[3:0];
    60: op1_00_in27 = reg_0871;
    53: op1_00_in27 = reg_0348;
    61: op1_00_in27 = reg_1212;
    67: op1_00_in27 = reg_0230;
    76: op1_00_in27 = reg_0820;
    71: op1_00_in27 = reg_0939;
    72: op1_00_in27 = reg_0162;
    55: op1_00_in27 = reg_0246;
    68: op1_00_in27 = reg_0045;
    74: op1_00_in27 = reg_0558;
    87: op1_00_in27 = reg_0562;
    78: op1_00_in27 = reg_0214;
    59: op1_00_in27 = reg_0047;
    110: op1_00_in27 = reg_0047;
    50: op1_00_in27 = reg_0757;
    86: op1_00_in27 = reg_0263;
    69: op1_00_in27 = reg_0885;
    36: op1_00_in27 = reg_0678;
    44: op1_00_in27 = reg_0586;
    88: op1_00_in27 = reg_1314;
    105: op1_00_in27 = reg_1314;
    56: op1_00_in27 = reg_0347;
    75: op1_00_in27 = reg_0232;
    42: op1_00_in27 = reg_0756;
    70: op1_00_in27 = reg_0963;
    57: op1_00_in27 = reg_0386;
    77: op1_00_in27 = reg_0151;
    51: op1_00_in27 = reg_0921;
    79: op1_00_in27 = reg_1474;
    43: op1_00_in27 = reg_0295;
    62: op1_00_in27 = reg_0572;
    80: op1_00_in27 = reg_1226;
    81: op1_00_in27 = reg_0430;
    89: op1_00_in27 = reg_1189;
    107: op1_00_in27 = reg_1189;
    63: op1_00_in27 = reg_1094;
    82: op1_00_in27 = reg_0598;
    83: op1_00_in27 = reg_0901;
    128: op1_00_in27 = reg_0901;
    64: op1_00_in27 = reg_1300;
    102: op1_00_in27 = reg_1300;
    84: op1_00_in27 = reg_0775;
    65: op1_00_in27 = reg_0612;
    90: op1_00_in27 = reg_0702;
    85: op1_00_in27 = reg_0989;
    91: op1_00_in27 = imem01_in[3:0];
    93: op1_00_in27 = reg_0412;
    94: op1_00_in27 = reg_0474;
    95: op1_00_in27 = reg_0023;
    96: op1_00_in27 = imem03_in[15:12];
    97: op1_00_in27 = reg_0759;
    99: op1_00_in27 = reg_0522;
    100: op1_00_in27 = reg_0875;
    101: op1_00_in27 = reg_0484;
    103: op1_00_in27 = reg_0195;
    106: op1_00_in27 = reg_0217;
    108: op1_00_in27 = reg_0585;
    109: op1_00_in27 = reg_1369;
    111: op1_00_in27 = reg_0996;
    112: op1_00_in27 = reg_0043;
    113: op1_00_in27 = reg_1403;
    114: op1_00_in27 = reg_0847;
    116: op1_00_in27 = reg_0550;
    117: op1_00_in27 = reg_0286;
    120: op1_00_in27 = reg_0632;
    121: op1_00_in27 = imem05_in[7:4];
    122: op1_00_in27 = imem07_in[11:8];
    123: op1_00_in27 = reg_0395;
    124: op1_00_in27 = reg_0190;
    126: op1_00_in27 = reg_0113;
    129: op1_00_in27 = reg_0730;
    130: op1_00_in27 = reg_0404;
    131: op1_00_in27 = reg_0475;
    default: op1_00_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv27 = 1;
    15: op1_00_inv27 = 1;
    19: op1_00_inv27 = 1;
    11: op1_00_inv27 = 1;
    33: op1_00_inv27 = 1;
    35: op1_00_inv27 = 1;
    26: op1_00_inv27 = 1;
    38: op1_00_inv27 = 1;
    39: op1_00_inv27 = 1;
    45: op1_00_inv27 = 1;
    52: op1_00_inv27 = 1;
    58: op1_00_inv27 = 1;
    54: op1_00_inv27 = 1;
    60: op1_00_inv27 = 1;
    53: op1_00_inv27 = 1;
    61: op1_00_inv27 = 1;
    72: op1_00_inv27 = 1;
    55: op1_00_inv27 = 1;
    68: op1_00_inv27 = 1;
    74: op1_00_inv27 = 1;
    50: op1_00_inv27 = 1;
    36: op1_00_inv27 = 1;
    44: op1_00_inv27 = 1;
    75: op1_00_inv27 = 1;
    42: op1_00_inv27 = 1;
    57: op1_00_inv27 = 1;
    43: op1_00_inv27 = 1;
    64: op1_00_inv27 = 1;
    84: op1_00_inv27 = 1;
    65: op1_00_inv27 = 1;
    85: op1_00_inv27 = 1;
    66: op1_00_inv27 = 1;
    91: op1_00_inv27 = 1;
    93: op1_00_inv27 = 1;
    94: op1_00_inv27 = 1;
    96: op1_00_inv27 = 1;
    100: op1_00_inv27 = 1;
    103: op1_00_inv27 = 1;
    105: op1_00_inv27 = 1;
    106: op1_00_inv27 = 1;
    107: op1_00_inv27 = 1;
    108: op1_00_inv27 = 1;
    111: op1_00_inv27 = 1;
    112: op1_00_inv27 = 1;
    113: op1_00_inv27 = 1;
    114: op1_00_inv27 = 1;
    121: op1_00_inv27 = 1;
    123: op1_00_inv27 = 1;
    124: op1_00_inv27 = 1;
    126: op1_00_inv27 = 1;
    128: op1_00_inv27 = 1;
    130: op1_00_inv27 = 1;
    131: op1_00_inv27 = 1;
    default: op1_00_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の28番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in28 = reg_0183;
    15: op1_00_in28 = reg_0069;
    19: op1_00_in28 = reg_0263;
    11: op1_00_in28 = reg_0067;
    33: op1_00_in28 = reg_0320;
    35: op1_00_in28 = reg_0558;
    32: op1_00_in28 = reg_0019;
    26: op1_00_in28 = reg_0269;
    41: op1_00_in28 = reg_0451;
    38: op1_00_in28 = reg_0676;
    39: op1_00_in28 = reg_0754;
    45: op1_00_in28 = reg_0140;
    52: op1_00_in28 = reg_0679;
    49: op1_00_in28 = reg_0780;
    58: op1_00_in28 = reg_0400;
    54: op1_00_in28 = reg_1143;
    60: op1_00_in28 = reg_0868;
    53: op1_00_in28 = reg_1000;
    61: op1_00_in28 = reg_0182;
    67: op1_00_in28 = reg_0892;
    76: op1_00_in28 = reg_1475;
    71: op1_00_in28 = reg_0197;
    72: op1_00_in28 = reg_1415;
    55: op1_00_in28 = imem03_in[11:8];
    68: op1_00_in28 = reg_0477;
    74: op1_00_in28 = reg_1226;
    87: op1_00_in28 = reg_0173;
    78: op1_00_in28 = imem07_in[11:8];
    59: op1_00_in28 = reg_0093;
    50: op1_00_in28 = reg_0732;
    86: op1_00_in28 = reg_1372;
    69: op1_00_in28 = reg_0411;
    36: op1_00_in28 = reg_0288;
    44: op1_00_in28 = reg_0570;
    88: op1_00_in28 = reg_0220;
    124: op1_00_in28 = reg_0220;
    56: op1_00_in28 = imem05_in[15:12];
    75: op1_00_in28 = reg_0378;
    42: op1_00_in28 = reg_0675;
    70: op1_00_in28 = reg_0246;
    57: op1_00_in28 = reg_0875;
    77: op1_00_in28 = reg_0014;
    51: op1_00_in28 = reg_0924;
    79: op1_00_in28 = reg_0967;
    43: op1_00_in28 = reg_0165;
    62: op1_00_in28 = reg_0968;
    80: op1_00_in28 = reg_1208;
    81: op1_00_in28 = reg_0402;
    89: op1_00_in28 = reg_0117;
    107: op1_00_in28 = reg_0117;
    63: op1_00_in28 = reg_0741;
    82: op1_00_in28 = reg_0471;
    83: op1_00_in28 = reg_0724;
    64: op1_00_in28 = reg_1301;
    105: op1_00_in28 = reg_1301;
    84: op1_00_in28 = reg_0774;
    65: op1_00_in28 = reg_0606;
    90: op1_00_in28 = reg_0278;
    85: op1_00_in28 = reg_1003;
    66: op1_00_in28 = reg_0139;
    91: op1_00_in28 = reg_0871;
    92: op1_00_in28 = reg_0636;
    93: op1_00_in28 = reg_1041;
    94: op1_00_in28 = reg_0846;
    95: op1_00_in28 = reg_0152;
    96: op1_00_in28 = reg_0507;
    97: op1_00_in28 = reg_1063;
    99: op1_00_in28 = reg_0132;
    100: op1_00_in28 = reg_0727;
    101: op1_00_in28 = reg_1182;
    102: op1_00_in28 = reg_1149;
    103: op1_00_in28 = reg_0046;
    106: op1_00_in28 = reg_0009;
    108: op1_00_in28 = reg_0527;
    109: op1_00_in28 = reg_0978;
    110: op1_00_in28 = reg_0550;
    111: op1_00_in28 = reg_0701;
    112: op1_00_in28 = reg_0012;
    113: op1_00_in28 = reg_0418;
    114: op1_00_in28 = reg_0556;
    116: op1_00_in28 = reg_0548;
    117: op1_00_in28 = reg_0437;
    120: op1_00_in28 = imem03_in[7:4];
    121: op1_00_in28 = reg_0832;
    122: op1_00_in28 = reg_0478;
    123: op1_00_in28 = reg_1268;
    126: op1_00_in28 = reg_0350;
    128: op1_00_in28 = reg_0175;
    129: op1_00_in28 = reg_0782;
    130: op1_00_in28 = reg_0123;
    131: op1_00_in28 = reg_1420;
    default: op1_00_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_00_inv28 = 1;
    11: op1_00_inv28 = 1;
    32: op1_00_inv28 = 1;
    52: op1_00_inv28 = 1;
    49: op1_00_inv28 = 1;
    58: op1_00_inv28 = 1;
    61: op1_00_inv28 = 1;
    55: op1_00_inv28 = 1;
    74: op1_00_inv28 = 1;
    87: op1_00_inv28 = 1;
    59: op1_00_inv28 = 1;
    50: op1_00_inv28 = 1;
    86: op1_00_inv28 = 1;
    88: op1_00_inv28 = 1;
    75: op1_00_inv28 = 1;
    70: op1_00_inv28 = 1;
    57: op1_00_inv28 = 1;
    80: op1_00_inv28 = 1;
    81: op1_00_inv28 = 1;
    63: op1_00_inv28 = 1;
    82: op1_00_inv28 = 1;
    83: op1_00_inv28 = 1;
    65: op1_00_inv28 = 1;
    90: op1_00_inv28 = 1;
    85: op1_00_inv28 = 1;
    66: op1_00_inv28 = 1;
    91: op1_00_inv28 = 1;
    93: op1_00_inv28 = 1;
    94: op1_00_inv28 = 1;
    100: op1_00_inv28 = 1;
    101: op1_00_inv28 = 1;
    102: op1_00_inv28 = 1;
    106: op1_00_inv28 = 1;
    107: op1_00_inv28 = 1;
    109: op1_00_inv28 = 1;
    113: op1_00_inv28 = 1;
    116: op1_00_inv28 = 1;
    117: op1_00_inv28 = 1;
    122: op1_00_inv28 = 1;
    123: op1_00_inv28 = 1;
    124: op1_00_inv28 = 1;
    128: op1_00_inv28 = 1;
    130: op1_00_inv28 = 1;
    default: op1_00_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の29番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in29 = reg_0294;
    15: op1_00_in29 = reg_0055;
    19: op1_00_in29 = reg_0264;
    11: op1_00_in29 = reg_0046;
    33: op1_00_in29 = reg_0291;
    35: op1_00_in29 = reg_0525;
    32: op1_00_in29 = reg_0020;
    26: op1_00_in29 = reg_0214;
    41: op1_00_in29 = reg_0430;
    38: op1_00_in29 = reg_0552;
    39: op1_00_in29 = reg_0752;
    45: op1_00_in29 = reg_0775;
    66: op1_00_in29 = reg_0775;
    52: op1_00_in29 = reg_0446;
    49: op1_00_in29 = reg_0160;
    58: op1_00_in29 = reg_0401;
    54: op1_00_in29 = reg_0595;
    60: op1_00_in29 = reg_0874;
    57: op1_00_in29 = reg_0874;
    53: op1_00_in29 = reg_0964;
    61: op1_00_in29 = reg_0045;
    67: op1_00_in29 = reg_0245;
    76: op1_00_in29 = reg_1474;
    71: op1_00_in29 = reg_0492;
    72: op1_00_in29 = reg_0025;
    55: op1_00_in29 = reg_0113;
    68: op1_00_in29 = reg_1373;
    74: op1_00_in29 = reg_1092;
    87: op1_00_in29 = reg_0566;
    78: op1_00_in29 = reg_0198;
    42: op1_00_in29 = reg_0198;
    59: op1_00_in29 = reg_0899;
    81: op1_00_in29 = reg_0899;
    50: op1_00_in29 = reg_0573;
    86: op1_00_in29 = reg_1368;
    69: op1_00_in29 = reg_0488;
    36: op1_00_in29 = imem03_in[7:4];
    44: op1_00_in29 = reg_0526;
    88: op1_00_in29 = reg_1300;
    56: op1_00_in29 = reg_0565;
    75: op1_00_in29 = reg_0640;
    70: op1_00_in29 = reg_0885;
    80: op1_00_in29 = reg_0885;
    64: op1_00_in29 = reg_0885;
    77: op1_00_in29 = reg_0458;
    126: op1_00_in29 = reg_0458;
    51: op1_00_in29 = reg_0139;
    79: op1_00_in29 = reg_0438;
    43: op1_00_in29 = reg_0461;
    62: op1_00_in29 = reg_0434;
    89: op1_00_in29 = reg_0370;
    63: op1_00_in29 = reg_0593;
    82: op1_00_in29 = reg_1041;
    83: op1_00_in29 = reg_0078;
    84: op1_00_in29 = reg_0030;
    65: op1_00_in29 = reg_0255;
    90: op1_00_in29 = reg_1168;
    85: op1_00_in29 = reg_1517;
    91: op1_00_in29 = reg_1255;
    92: op1_00_in29 = reg_0584;
    93: op1_00_in29 = reg_1004;
    94: op1_00_in29 = reg_0561;
    95: op1_00_in29 = imem07_in[3:0];
    96: op1_00_in29 = reg_0840;
    97: op1_00_in29 = reg_1425;
    99: op1_00_in29 = reg_0119;
    100: op1_00_in29 = reg_0464;
    102: op1_00_in29 = reg_0378;
    103: op1_00_in29 = reg_0022;
    105: op1_00_in29 = reg_0558;
    106: op1_00_in29 = reg_0279;
    107: op1_00_in29 = reg_0536;
    108: op1_00_in29 = reg_0132;
    109: op1_00_in29 = reg_1203;
    110: op1_00_in29 = reg_0548;
    111: op1_00_in29 = reg_1401;
    112: op1_00_in29 = reg_0662;
    113: op1_00_in29 = reg_0601;
    114: op1_00_in29 = reg_0965;
    116: op1_00_in29 = reg_0746;
    117: op1_00_in29 = reg_0415;
    120: op1_00_in29 = imem03_in[11:8];
    121: op1_00_in29 = reg_0136;
    122: op1_00_in29 = reg_1060;
    123: op1_00_in29 = reg_1059;
    124: op1_00_in29 = reg_0507;
    128: op1_00_in29 = reg_0727;
    129: op1_00_in29 = reg_0696;
    131: op1_00_in29 = reg_0782;
    default: op1_00_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    11: op1_00_inv29 = 1;
    33: op1_00_inv29 = 1;
    35: op1_00_inv29 = 1;
    26: op1_00_inv29 = 1;
    41: op1_00_inv29 = 1;
    39: op1_00_inv29 = 1;
    49: op1_00_inv29 = 1;
    58: op1_00_inv29 = 1;
    60: op1_00_inv29 = 1;
    53: op1_00_inv29 = 1;
    61: op1_00_inv29 = 1;
    67: op1_00_inv29 = 1;
    68: op1_00_inv29 = 1;
    87: op1_00_inv29 = 1;
    59: op1_00_inv29 = 1;
    50: op1_00_inv29 = 1;
    69: op1_00_inv29 = 1;
    56: op1_00_inv29 = 1;
    42: op1_00_inv29 = 1;
    70: op1_00_inv29 = 1;
    57: op1_00_inv29 = 1;
    43: op1_00_inv29 = 1;
    62: op1_00_inv29 = 1;
    80: op1_00_inv29 = 1;
    81: op1_00_inv29 = 1;
    82: op1_00_inv29 = 1;
    83: op1_00_inv29 = 1;
    64: op1_00_inv29 = 1;
    84: op1_00_inv29 = 1;
    91: op1_00_inv29 = 1;
    97: op1_00_inv29 = 1;
    102: op1_00_inv29 = 1;
    105: op1_00_inv29 = 1;
    109: op1_00_inv29 = 1;
    110: op1_00_inv29 = 1;
    113: op1_00_inv29 = 1;
    114: op1_00_inv29 = 1;
    116: op1_00_inv29 = 1;
    121: op1_00_inv29 = 1;
    122: op1_00_inv29 = 1;
    123: op1_00_inv29 = 1;
    124: op1_00_inv29 = 1;
    126: op1_00_inv29 = 1;
    129: op1_00_inv29 = 1;
    131: op1_00_inv29 = 1;
    default: op1_00_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の30番目の入力
  always @ ( * ) begin
    case ( state )
    20: op1_00_in30 = reg_0047;
    15: op1_00_in30 = reg_0024;
    19: op1_00_in30 = reg_0247;
    69: op1_00_in30 = reg_0247;
    11: op1_00_in30 = reg_0023;
    33: op1_00_in30 = reg_0277;
    35: op1_00_in30 = reg_0504;
    70: op1_00_in30 = reg_0504;
    32: op1_00_in30 = imem05_in[7:4];
    26: op1_00_in30 = reg_0022;
    41: op1_00_in30 = reg_0148;
    38: op1_00_in30 = reg_0420;
    107: op1_00_in30 = reg_0420;
    39: op1_00_in30 = reg_0720;
    129: op1_00_in30 = reg_0720;
    45: op1_00_in30 = reg_0740;
    52: op1_00_in30 = imem02_in[7:4];
    112: op1_00_in30 = imem02_in[7:4];
    49: op1_00_in30 = reg_0979;
    58: op1_00_in30 = reg_0899;
    79: op1_00_in30 = reg_0899;
    54: op1_00_in30 = reg_0577;
    60: op1_00_in30 = reg_0079;
    53: op1_00_in30 = reg_0962;
    61: op1_00_in30 = reg_1181;
    67: op1_00_in30 = reg_1349;
    76: op1_00_in30 = reg_1452;
    71: op1_00_in30 = reg_1348;
    72: op1_00_in30 = reg_0667;
    55: op1_00_in30 = reg_0506;
    68: op1_00_in30 = reg_0274;
    74: op1_00_in30 = reg_0113;
    87: op1_00_in30 = reg_0564;
    78: op1_00_in30 = reg_1056;
    59: op1_00_in30 = reg_0901;
    81: op1_00_in30 = reg_0901;
    50: op1_00_in30 = reg_0677;
    86: op1_00_in30 = imem04_in[3:0];
    36: op1_00_in30 = imem03_in[15:12];
    44: op1_00_in30 = reg_0529;
    88: op1_00_in30 = reg_1231;
    56: op1_00_in30 = reg_0539;
    75: op1_00_in30 = reg_0234;
    42: op1_00_in30 = reg_0707;
    57: op1_00_in30 = reg_0080;
    77: op1_00_in30 = reg_0192;
    51: op1_00_in30 = reg_0791;
    43: op1_00_in30 = reg_0460;
    62: op1_00_in30 = reg_0727;
    80: op1_00_in30 = reg_0882;
    64: op1_00_in30 = reg_0882;
    89: op1_00_in30 = imem05_in[11:8];
    63: op1_00_in30 = reg_0591;
    82: op1_00_in30 = reg_0454;
    83: op1_00_in30 = reg_0042;
    84: op1_00_in30 = reg_0284;
    65: op1_00_in30 = reg_0497;
    90: op1_00_in30 = reg_1169;
    85: op1_00_in30 = reg_0349;
    66: op1_00_in30 = reg_0003;
    91: op1_00_in30 = reg_1253;
    92: op1_00_in30 = reg_0619;
    93: op1_00_in30 = reg_0451;
    94: op1_00_in30 = reg_0436;
    95: op1_00_in30 = reg_0299;
    96: op1_00_in30 = reg_0889;
    97: op1_00_in30 = reg_1033;
    99: op1_00_in30 = reg_0244;
    100: op1_00_in30 = reg_0400;
    128: op1_00_in30 = reg_0400;
    102: op1_00_in30 = reg_1009;
    103: op1_00_in30 = imem07_in[15:12];
    105: op1_00_in30 = reg_0178;
    106: op1_00_in30 = reg_0632;
    108: op1_00_in30 = reg_0396;
    109: op1_00_in30 = reg_0681;
    110: op1_00_in30 = reg_0241;
    111: op1_00_in30 = reg_1373;
    113: op1_00_in30 = reg_0393;
    114: op1_00_in30 = reg_0314;
    116: op1_00_in30 = reg_0260;
    117: op1_00_in30 = reg_0100;
    120: op1_00_in30 = reg_0179;
    121: op1_00_in30 = reg_0702;
    122: op1_00_in30 = reg_1345;
    123: op1_00_in30 = reg_0793;
    124: op1_00_in30 = reg_0198;
    126: op1_00_in30 = reg_0790;
    131: op1_00_in30 = reg_1437;
    default: op1_00_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    20: op1_00_inv30 = 1;
    19: op1_00_inv30 = 1;
    11: op1_00_inv30 = 1;
    35: op1_00_inv30 = 1;
    32: op1_00_inv30 = 1;
    41: op1_00_inv30 = 1;
    38: op1_00_inv30 = 1;
    52: op1_00_inv30 = 1;
    49: op1_00_inv30 = 1;
    58: op1_00_inv30 = 1;
    60: op1_00_inv30 = 1;
    61: op1_00_inv30 = 1;
    67: op1_00_inv30 = 1;
    71: op1_00_inv30 = 1;
    55: op1_00_inv30 = 1;
    50: op1_00_inv30 = 1;
    69: op1_00_inv30 = 1;
    75: op1_00_inv30 = 1;
    42: op1_00_inv30 = 1;
    77: op1_00_inv30 = 1;
    43: op1_00_inv30 = 1;
    62: op1_00_inv30 = 1;
    81: op1_00_inv30 = 1;
    63: op1_00_inv30 = 1;
    65: op1_00_inv30 = 1;
    66: op1_00_inv30 = 1;
    91: op1_00_inv30 = 1;
    94: op1_00_inv30 = 1;
    100: op1_00_inv30 = 1;
    107: op1_00_inv30 = 1;
    110: op1_00_inv30 = 1;
    124: op1_00_inv30 = 1;
    126: op1_00_inv30 = 1;
    129: op1_00_inv30 = 1;
    default: op1_00_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_00_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_00_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の0番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in00 = imem06_in[11:8];
    52: op1_01_in00 = imem02_in[15:12];
    90: op1_01_in00 = imem02_in[15:12];
    91: op1_01_in00 = imem02_in[15:12];
    112: op1_01_in00 = imem02_in[15:12];
    49: op1_01_in00 = imem07_in[11:8];
    5: op1_01_in00 = imem07_in[11:8];
    53: op1_01_in00 = reg_0362;
    67: op1_01_in00 = imem03_in[3:0];
    61: op1_01_in00 = reg_0616;
    54: op1_01_in00 = imem07_in[3:0];
    22: op1_01_in00 = imem07_in[3:0];
    72: op1_01_in00 = reg_0555;
    58: op1_01_in00 = imem07_in[15:12];
    68: op1_01_in00 = reg_0233;
    96: op1_01_in00 = reg_0233;
    55: op1_01_in00 = reg_0594;
    73: op1_01_in00 = reg_0697;
    71: op1_01_in00 = reg_0615;
    48: op1_01_in00 = reg_0742;
    110: op1_01_in00 = reg_0742;
    86: op1_01_in00 = reg_1184;
    69: op1_01_in00 = reg_0709;
    59: op1_01_in00 = reg_1099;
    50: op1_01_in00 = reg_0282;
    60: op1_01_in00 = reg_0042;
    33: op1_01_in00 = imem07_in[7:4];
    25: op1_01_in00 = imem07_in[7:4];
    24: op1_01_in00 = imem07_in[7:4];
    46: op1_01_in00 = reg_0234;
    74: op1_01_in00 = reg_0582;
    47: op1_01_in00 = reg_0527;
    75: op1_01_in00 = reg_0147;
    44: op1_01_in00 = reg_0338;
    56: op1_01_in00 = reg_0104;
    87: op1_01_in00 = reg_0975;
    40: op1_01_in00 = reg_0310;
    37: op1_01_in00 = reg_0465;
    76: op1_01_in00 = imem00_in[3:0];
    84: op1_01_in00 = imem00_in[3:0];
    115: op1_01_in00 = imem00_in[3:0];
    127: op1_01_in00 = imem00_in[3:0];
    57: op1_01_in00 = reg_0270;
    70: op1_01_in00 = reg_0889;
    77: op1_01_in00 = reg_0369;
    4: op1_01_in00 = reg_0003;
    28: op1_01_in00 = reg_0002;
    88: op1_01_in00 = reg_1325;
    34: op1_01_in00 = reg_0029;
    51: op1_01_in00 = reg_0923;
    78: op1_01_in00 = imem00_in[15:12];
    82: op1_01_in00 = imem00_in[15:12];
    85: op1_01_in00 = imem00_in[15:12];
    92: op1_01_in00 = imem00_in[15:12];
    117: op1_01_in00 = imem00_in[15:12];
    118: op1_01_in00 = imem00_in[15:12];
    119: op1_01_in00 = imem00_in[15:12];
    42: op1_01_in00 = reg_0819;
    79: op1_01_in00 = reg_1502;
    35: op1_01_in00 = reg_0438;
    62: op1_01_in00 = reg_0445;
    121: op1_01_in00 = reg_0445;
    80: op1_01_in00 = imem00_in[7:4];
    104: op1_01_in00 = imem00_in[7:4];
    122: op1_01_in00 = imem00_in[7:4];
    125: op1_01_in00 = imem00_in[7:4];
    130: op1_01_in00 = imem00_in[7:4];
    81: op1_01_in00 = reg_0983;
    89: op1_01_in00 = reg_0481;
    63: op1_01_in00 = reg_0743;
    83: op1_01_in00 = reg_0044;
    39: op1_01_in00 = reg_0330;
    64: op1_01_in00 = reg_0363;
    65: op1_01_in00 = reg_0474;
    66: op1_01_in00 = reg_0866;
    93: op1_01_in00 = reg_0097;
    94: op1_01_in00 = reg_0054;
    95: op1_01_in00 = imem00_in[11:8];
    98: op1_01_in00 = imem00_in[11:8];
    101: op1_01_in00 = imem00_in[11:8];
    97: op1_01_in00 = reg_0198;
    99: op1_01_in00 = reg_1204;
    100: op1_01_in00 = reg_0078;
    102: op1_01_in00 = imem05_in[7:4];
    103: op1_01_in00 = reg_0489;
    105: op1_01_in00 = reg_1208;
    106: op1_01_in00 = imem03_in[11:8];
    107: op1_01_in00 = reg_0020;
    27: op1_01_in00 = reg_0247;
    108: op1_01_in00 = reg_0977;
    109: op1_01_in00 = reg_0969;
    38: op1_01_in00 = reg_0442;
    111: op1_01_in00 = reg_0344;
    113: op1_01_in00 = reg_0130;
    114: op1_01_in00 = reg_0349;
    29: op1_01_in00 = reg_0186;
    116: op1_01_in00 = reg_0383;
    43: op1_01_in00 = imem04_in[15:12];
    120: op1_01_in00 = reg_0706;
    123: op1_01_in00 = reg_0604;
    124: op1_01_in00 = reg_1001;
    126: op1_01_in00 = reg_0443;
    128: op1_01_in00 = reg_0077;
    129: op1_01_in00 = reg_0752;
    131: op1_01_in00 = reg_0271;
    default: op1_01_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv00 = 1;
    53: op1_01_inv00 = 1;
    67: op1_01_inv00 = 1;
    72: op1_01_inv00 = 1;
    58: op1_01_inv00 = 1;
    59: op1_01_inv00 = 1;
    50: op1_01_inv00 = 1;
    60: op1_01_inv00 = 1;
    74: op1_01_inv00 = 1;
    56: op1_01_inv00 = 1;
    87: op1_01_inv00 = 1;
    76: op1_01_inv00 = 1;
    57: op1_01_inv00 = 1;
    88: op1_01_inv00 = 1;
    34: op1_01_inv00 = 1;
    51: op1_01_inv00 = 1;
    78: op1_01_inv00 = 1;
    42: op1_01_inv00 = 1;
    63: op1_01_inv00 = 1;
    83: op1_01_inv00 = 1;
    39: op1_01_inv00 = 1;
    85: op1_01_inv00 = 1;
    92: op1_01_inv00 = 1;
    25: op1_01_inv00 = 1;
    93: op1_01_inv00 = 1;
    94: op1_01_inv00 = 1;
    95: op1_01_inv00 = 1;
    97: op1_01_inv00 = 1;
    98: op1_01_inv00 = 1;
    99: op1_01_inv00 = 1;
    100: op1_01_inv00 = 1;
    101: op1_01_inv00 = 1;
    104: op1_01_inv00 = 1;
    109: op1_01_inv00 = 1;
    110: op1_01_inv00 = 1;
    38: op1_01_inv00 = 1;
    111: op1_01_inv00 = 1;
    112: op1_01_inv00 = 1;
    113: op1_01_inv00 = 1;
    5: op1_01_inv00 = 1;
    114: op1_01_inv00 = 1;
    115: op1_01_inv00 = 1;
    119: op1_01_inv00 = 1;
    124: op1_01_inv00 = 1;
    125: op1_01_inv00 = 1;
    127: op1_01_inv00 = 1;
    129: op1_01_inv00 = 1;
    131: op1_01_inv00 = 1;
    default: op1_01_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の1番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in01 = reg_0119;
    47: op1_01_in01 = reg_0119;
    52: op1_01_in01 = reg_1098;
    49: op1_01_in01 = reg_0465;
    53: op1_01_in01 = reg_0047;
    67: op1_01_in01 = reg_0830;
    61: op1_01_in01 = reg_0615;
    72: op1_01_in01 = reg_0701;
    123: op1_01_in01 = reg_0701;
    58: op1_01_in01 = reg_0998;
    68: op1_01_in01 = reg_0972;
    55: op1_01_in01 = reg_0463;
    73: op1_01_in01 = reg_0090;
    71: op1_01_in01 = reg_0791;
    85: op1_01_in01 = reg_0791;
    48: op1_01_in01 = reg_0430;
    86: op1_01_in01 = reg_0954;
    69: op1_01_in01 = reg_1063;
    59: op1_01_in01 = imem00_in[15:12];
    95: op1_01_in01 = imem00_in[15:12];
    50: op1_01_in01 = reg_0679;
    60: op1_01_in01 = reg_0041;
    33: op1_01_in01 = reg_0593;
    46: op1_01_in01 = imem03_in[7:4];
    74: op1_01_in01 = reg_0340;
    75: op1_01_in01 = reg_0148;
    44: op1_01_in01 = reg_0097;
    109: op1_01_in01 = reg_0097;
    56: op1_01_in01 = reg_0506;
    87: op1_01_in01 = reg_1369;
    40: op1_01_in01 = reg_0298;
    37: op1_01_in01 = reg_0665;
    76: op1_01_in01 = reg_0983;
    57: op1_01_in01 = reg_0271;
    70: op1_01_in01 = reg_0474;
    22: op1_01_in01 = reg_0001;
    77: op1_01_in01 = reg_0582;
    4: op1_01_in01 = imem07_in[3:0];
    28: op1_01_in01 = reg_0003;
    88: op1_01_in01 = reg_0443;
    34: op1_01_in01 = imem07_in[7:4];
    51: op1_01_in01 = reg_0140;
    78: op1_01_in01 = reg_0806;
    101: op1_01_in01 = reg_0806;
    42: op1_01_in01 = reg_0120;
    79: op1_01_in01 = reg_0210;
    35: op1_01_in01 = reg_0162;
    62: op1_01_in01 = reg_1242;
    80: op1_01_in01 = reg_1278;
    81: op1_01_in01 = reg_0907;
    89: op1_01_in01 = reg_0263;
    63: op1_01_in01 = reg_0161;
    82: op1_01_in01 = reg_1490;
    83: op1_01_in01 = reg_0012;
    39: op1_01_in01 = reg_0744;
    64: op1_01_in01 = reg_0093;
    84: op1_01_in01 = reg_0868;
    65: op1_01_in01 = reg_0494;
    90: op1_01_in01 = reg_1002;
    66: op1_01_in01 = reg_0803;
    91: op1_01_in01 = reg_0878;
    92: op1_01_in01 = reg_0725;
    98: op1_01_in01 = reg_0725;
    25: op1_01_in01 = reg_0031;
    93: op1_01_in01 = reg_1189;
    94: op1_01_in01 = reg_0326;
    96: op1_01_in01 = reg_0154;
    97: op1_01_in01 = reg_0312;
    99: op1_01_in01 = reg_0018;
    100: op1_01_in01 = reg_0257;
    128: op1_01_in01 = reg_0257;
    102: op1_01_in01 = reg_0197;
    103: op1_01_in01 = reg_1094;
    104: op1_01_in01 = imem00_in[11:8];
    105: op1_01_in01 = reg_0104;
    106: op1_01_in01 = imem03_in[15:12];
    107: op1_01_in01 = imem05_in[3:0];
    27: op1_01_in01 = reg_0296;
    108: op1_01_in01 = reg_0213;
    110: op1_01_in01 = reg_0468;
    38: op1_01_in01 = reg_0739;
    111: op1_01_in01 = reg_0206;
    113: op1_01_in01 = reg_0206;
    112: op1_01_in01 = reg_0606;
    5: op1_01_in01 = imem07_in[15:12];
    114: op1_01_in01 = reg_0952;
    29: op1_01_in01 = reg_0085;
    115: op1_01_in01 = reg_1277;
    116: op1_01_in01 = reg_0899;
    117: op1_01_in01 = reg_1081;
    118: op1_01_in01 = reg_1244;
    43: op1_01_in01 = reg_0199;
    119: op1_01_in01 = reg_1470;
    120: op1_01_in01 = reg_1000;
    121: op1_01_in01 = reg_0205;
    122: op1_01_in01 = reg_0959;
    124: op1_01_in01 = reg_0783;
    125: op1_01_in01 = reg_0748;
    126: op1_01_in01 = reg_0411;
    127: op1_01_in01 = reg_0581;
    129: op1_01_in01 = reg_0827;
    130: op1_01_in01 = reg_0640;
    131: op1_01_in01 = reg_1467;
    24: op1_01_in01 = reg_0100;
    default: op1_01_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_01_inv01 = 1;
    49: op1_01_inv01 = 1;
    53: op1_01_inv01 = 1;
    67: op1_01_inv01 = 1;
    61: op1_01_inv01 = 1;
    72: op1_01_inv01 = 1;
    58: op1_01_inv01 = 1;
    68: op1_01_inv01 = 1;
    73: op1_01_inv01 = 1;
    71: op1_01_inv01 = 1;
    86: op1_01_inv01 = 1;
    69: op1_01_inv01 = 1;
    60: op1_01_inv01 = 1;
    47: op1_01_inv01 = 1;
    75: op1_01_inv01 = 1;
    56: op1_01_inv01 = 1;
    76: op1_01_inv01 = 1;
    22: op1_01_inv01 = 1;
    4: op1_01_inv01 = 1;
    28: op1_01_inv01 = 1;
    88: op1_01_inv01 = 1;
    34: op1_01_inv01 = 1;
    78: op1_01_inv01 = 1;
    42: op1_01_inv01 = 1;
    35: op1_01_inv01 = 1;
    80: op1_01_inv01 = 1;
    81: op1_01_inv01 = 1;
    83: op1_01_inv01 = 1;
    39: op1_01_inv01 = 1;
    64: op1_01_inv01 = 1;
    65: op1_01_inv01 = 1;
    25: op1_01_inv01 = 1;
    93: op1_01_inv01 = 1;
    95: op1_01_inv01 = 1;
    96: op1_01_inv01 = 1;
    97: op1_01_inv01 = 1;
    99: op1_01_inv01 = 1;
    102: op1_01_inv01 = 1;
    106: op1_01_inv01 = 1;
    108: op1_01_inv01 = 1;
    110: op1_01_inv01 = 1;
    38: op1_01_inv01 = 1;
    112: op1_01_inv01 = 1;
    5: op1_01_inv01 = 1;
    117: op1_01_inv01 = 1;
    118: op1_01_inv01 = 1;
    43: op1_01_inv01 = 1;
    122: op1_01_inv01 = 1;
    129: op1_01_inv01 = 1;
    24: op1_01_inv01 = 1;
    default: op1_01_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の2番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in02 = reg_0067;
    52: op1_01_in02 = reg_0606;
    49: op1_01_in02 = reg_0741;
    53: op1_01_in02 = reg_0724;
    67: op1_01_in02 = reg_0557;
    61: op1_01_in02 = reg_0669;
    72: op1_01_in02 = reg_0672;
    58: op1_01_in02 = reg_0496;
    68: op1_01_in02 = reg_0128;
    55: op1_01_in02 = reg_0978;
    73: op1_01_in02 = reg_0197;
    71: op1_01_in02 = reg_1278;
    48: op1_01_in02 = reg_0402;
    35: op1_01_in02 = reg_0402;
    128: op1_01_in02 = reg_0402;
    86: op1_01_in02 = reg_1093;
    69: op1_01_in02 = reg_1149;
    59: op1_01_in02 = reg_1242;
    50: op1_01_in02 = reg_0254;
    60: op1_01_in02 = reg_0446;
    33: op1_01_in02 = reg_0361;
    46: op1_01_in02 = imem03_in[15:12];
    74: op1_01_in02 = imem04_in[7:4];
    47: op1_01_in02 = reg_0244;
    75: op1_01_in02 = reg_0146;
    44: op1_01_in02 = reg_0094;
    56: op1_01_in02 = reg_0000;
    87: op1_01_in02 = reg_0535;
    40: op1_01_in02 = imem07_in[7:4];
    37: op1_01_in02 = reg_0287;
    76: op1_01_in02 = reg_0841;
    127: op1_01_in02 = reg_0841;
    57: op1_01_in02 = reg_0152;
    70: op1_01_in02 = reg_0326;
    22: op1_01_in02 = reg_0004;
    77: op1_01_in02 = reg_0340;
    28: op1_01_in02 = reg_0050;
    88: op1_01_in02 = imem04_in[15:12];
    34: op1_01_in02 = reg_0103;
    51: op1_01_in02 = reg_0031;
    78: op1_01_in02 = reg_0218;
    42: op1_01_in02 = reg_0258;
    79: op1_01_in02 = reg_1430;
    62: op1_01_in02 = reg_0523;
    80: op1_01_in02 = reg_1277;
    81: op1_01_in02 = reg_1281;
    89: op1_01_in02 = reg_0088;
    63: op1_01_in02 = reg_0553;
    82: op1_01_in02 = reg_0615;
    83: op1_01_in02 = imem01_in[15:12];
    39: op1_01_in02 = reg_0487;
    64: op1_01_in02 = reg_0292;
    84: op1_01_in02 = reg_1079;
    65: op1_01_in02 = reg_0433;
    85: op1_01_in02 = reg_0907;
    90: op1_01_in02 = reg_0495;
    66: op1_01_in02 = reg_1052;
    91: op1_01_in02 = reg_0829;
    92: op1_01_in02 = reg_0445;
    25: op1_01_in02 = reg_0030;
    93: op1_01_in02 = reg_0633;
    94: op1_01_in02 = reg_0778;
    95: op1_01_in02 = reg_0501;
    98: op1_01_in02 = reg_0501;
    96: op1_01_in02 = reg_0444;
    97: op1_01_in02 = reg_0789;
    99: op1_01_in02 = imem07_in[3:0];
    100: op1_01_in02 = reg_0044;
    101: op1_01_in02 = reg_0580;
    102: op1_01_in02 = reg_0492;
    103: op1_01_in02 = reg_0779;
    104: op1_01_in02 = reg_0748;
    115: op1_01_in02 = reg_0748;
    105: op1_01_in02 = reg_0541;
    106: op1_01_in02 = reg_0677;
    107: op1_01_in02 = imem05_in[11:8];
    27: op1_01_in02 = reg_0132;
    108: op1_01_in02 = reg_0015;
    109: op1_01_in02 = reg_1312;
    110: op1_01_in02 = reg_0715;
    38: op1_01_in02 = reg_0593;
    111: op1_01_in02 = reg_0014;
    112: op1_01_in02 = reg_0456;
    113: op1_01_in02 = imem06_in[15:12];
    114: op1_01_in02 = reg_0558;
    29: op1_01_in02 = reg_0123;
    116: op1_01_in02 = reg_0078;
    117: op1_01_in02 = reg_0843;
    118: op1_01_in02 = reg_0638;
    43: op1_01_in02 = reg_0305;
    119: op1_01_in02 = reg_1081;
    120: op1_01_in02 = reg_1425;
    121: op1_01_in02 = reg_0831;
    122: op1_01_in02 = reg_0958;
    123: op1_01_in02 = reg_0630;
    124: op1_01_in02 = reg_0234;
    125: op1_01_in02 = reg_1141;
    126: op1_01_in02 = imem04_in[3:0];
    129: op1_01_in02 = reg_0194;
    130: op1_01_in02 = reg_1028;
    131: op1_01_in02 = reg_0720;
    24: op1_01_in02 = reg_0229;
    default: op1_01_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_01_inv02 = 1;
    53: op1_01_inv02 = 1;
    67: op1_01_inv02 = 1;
    61: op1_01_inv02 = 1;
    73: op1_01_inv02 = 1;
    71: op1_01_inv02 = 1;
    48: op1_01_inv02 = 1;
    50: op1_01_inv02 = 1;
    60: op1_01_inv02 = 1;
    74: op1_01_inv02 = 1;
    47: op1_01_inv02 = 1;
    75: op1_01_inv02 = 1;
    44: op1_01_inv02 = 1;
    40: op1_01_inv02 = 1;
    57: op1_01_inv02 = 1;
    70: op1_01_inv02 = 1;
    88: op1_01_inv02 = 1;
    34: op1_01_inv02 = 1;
    42: op1_01_inv02 = 1;
    79: op1_01_inv02 = 1;
    35: op1_01_inv02 = 1;
    62: op1_01_inv02 = 1;
    80: op1_01_inv02 = 1;
    81: op1_01_inv02 = 1;
    63: op1_01_inv02 = 1;
    39: op1_01_inv02 = 1;
    64: op1_01_inv02 = 1;
    65: op1_01_inv02 = 1;
    90: op1_01_inv02 = 1;
    66: op1_01_inv02 = 1;
    92: op1_01_inv02 = 1;
    94: op1_01_inv02 = 1;
    95: op1_01_inv02 = 1;
    96: op1_01_inv02 = 1;
    98: op1_01_inv02 = 1;
    100: op1_01_inv02 = 1;
    101: op1_01_inv02 = 1;
    102: op1_01_inv02 = 1;
    27: op1_01_inv02 = 1;
    108: op1_01_inv02 = 1;
    109: op1_01_inv02 = 1;
    110: op1_01_inv02 = 1;
    111: op1_01_inv02 = 1;
    114: op1_01_inv02 = 1;
    29: op1_01_inv02 = 1;
    117: op1_01_inv02 = 1;
    118: op1_01_inv02 = 1;
    121: op1_01_inv02 = 1;
    126: op1_01_inv02 = 1;
    127: op1_01_inv02 = 1;
    129: op1_01_inv02 = 1;
    default: op1_01_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の3番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in03 = reg_0213;
    52: op1_01_in03 = reg_0922;
    49: op1_01_in03 = reg_0413;
    53: op1_01_in03 = reg_0868;
    67: op1_01_in03 = reg_0177;
    61: op1_01_in03 = reg_1081;
    72: op1_01_in03 = reg_1278;
    58: op1_01_in03 = reg_0394;
    68: op1_01_in03 = reg_0127;
    55: op1_01_in03 = imem04_in[3:0];
    73: op1_01_in03 = reg_0601;
    71: op1_01_in03 = reg_1279;
    48: op1_01_in03 = reg_0092;
    86: op1_01_in03 = reg_0479;
    69: op1_01_in03 = imem03_in[7:4];
    59: op1_01_in03 = reg_0804;
    50: op1_01_in03 = reg_0255;
    60: op1_01_in03 = reg_0399;
    33: op1_01_in03 = reg_0228;
    34: op1_01_in03 = reg_0228;
    46: op1_01_in03 = reg_0556;
    74: op1_01_in03 = reg_0626;
    47: op1_01_in03 = reg_0268;
    75: op1_01_in03 = reg_0901;
    44: op1_01_in03 = reg_0237;
    56: op1_01_in03 = reg_0425;
    87: op1_01_in03 = reg_1257;
    40: op1_01_in03 = imem07_in[11:8];
    99: op1_01_in03 = imem07_in[11:8];
    37: op1_01_in03 = reg_0442;
    76: op1_01_in03 = reg_1078;
    57: op1_01_in03 = reg_0230;
    70: op1_01_in03 = reg_0973;
    77: op1_01_in03 = reg_0487;
    28: op1_01_in03 = imem07_in[15:12];
    88: op1_01_in03 = reg_1312;
    51: op1_01_in03 = reg_0029;
    78: op1_01_in03 = reg_0523;
    66: op1_01_in03 = reg_0523;
    42: op1_01_in03 = reg_0238;
    79: op1_01_in03 = reg_1268;
    35: op1_01_in03 = reg_0400;
    62: op1_01_in03 = reg_0476;
    80: op1_01_in03 = reg_1079;
    81: op1_01_in03 = reg_1242;
    89: op1_01_in03 = reg_1040;
    63: op1_01_in03 = reg_0982;
    82: op1_01_in03 = reg_0580;
    83: op1_01_in03 = reg_0332;
    39: op1_01_in03 = reg_0463;
    64: op1_01_in03 = reg_0012;
    84: op1_01_in03 = reg_1489;
    104: op1_01_in03 = reg_1489;
    65: op1_01_in03 = reg_0971;
    94: op1_01_in03 = reg_0971;
    85: op1_01_in03 = reg_1277;
    90: op1_01_in03 = reg_1207;
    91: op1_01_in03 = reg_0897;
    92: op1_01_in03 = reg_0841;
    95: op1_01_in03 = reg_0841;
    25: op1_01_in03 = reg_0102;
    93: op1_01_in03 = reg_0016;
    96: op1_01_in03 = reg_0216;
    120: op1_01_in03 = reg_0216;
    97: op1_01_in03 = reg_1494;
    98: op1_01_in03 = reg_0907;
    118: op1_01_in03 = reg_0907;
    100: op1_01_in03 = reg_0447;
    101: op1_01_in03 = reg_0153;
    102: op1_01_in03 = reg_0240;
    103: op1_01_in03 = reg_0465;
    105: op1_01_in03 = reg_0025;
    106: op1_01_in03 = reg_0559;
    107: op1_01_in03 = reg_0466;
    27: op1_01_in03 = imem06_in[11:8];
    108: op1_01_in03 = imem07_in[3:0];
    109: op1_01_in03 = reg_1151;
    110: op1_01_in03 = reg_0430;
    38: op1_01_in03 = reg_0100;
    111: op1_01_in03 = imem06_in[7:4];
    112: op1_01_in03 = reg_1260;
    113: op1_01_in03 = reg_0729;
    114: op1_01_in03 = reg_1092;
    115: op1_01_in03 = reg_0806;
    125: op1_01_in03 = reg_0806;
    116: op1_01_in03 = reg_1071;
    117: op1_01_in03 = reg_0486;
    43: op1_01_in03 = reg_0719;
    119: op1_01_in03 = reg_0748;
    122: op1_01_in03 = reg_0748;
    121: op1_01_in03 = reg_0182;
    123: op1_01_in03 = reg_1401;
    124: op1_01_in03 = reg_0142;
    126: op1_01_in03 = reg_0032;
    127: op1_01_in03 = reg_0387;
    128: op1_01_in03 = reg_0044;
    129: op1_01_in03 = reg_0374;
    130: op1_01_in03 = reg_0485;
    131: op1_01_in03 = reg_0752;
    24: op1_01_in03 = reg_0135;
    default: op1_01_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv03 = 1;
    49: op1_01_inv03 = 1;
    53: op1_01_inv03 = 1;
    61: op1_01_inv03 = 1;
    55: op1_01_inv03 = 1;
    71: op1_01_inv03 = 1;
    69: op1_01_inv03 = 1;
    59: op1_01_inv03 = 1;
    50: op1_01_inv03 = 1;
    60: op1_01_inv03 = 1;
    46: op1_01_inv03 = 1;
    47: op1_01_inv03 = 1;
    44: op1_01_inv03 = 1;
    56: op1_01_inv03 = 1;
    40: op1_01_inv03 = 1;
    57: op1_01_inv03 = 1;
    77: op1_01_inv03 = 1;
    28: op1_01_inv03 = 1;
    88: op1_01_inv03 = 1;
    51: op1_01_inv03 = 1;
    78: op1_01_inv03 = 1;
    42: op1_01_inv03 = 1;
    79: op1_01_inv03 = 1;
    62: op1_01_inv03 = 1;
    80: op1_01_inv03 = 1;
    83: op1_01_inv03 = 1;
    39: op1_01_inv03 = 1;
    64: op1_01_inv03 = 1;
    84: op1_01_inv03 = 1;
    90: op1_01_inv03 = 1;
    91: op1_01_inv03 = 1;
    92: op1_01_inv03 = 1;
    93: op1_01_inv03 = 1;
    94: op1_01_inv03 = 1;
    96: op1_01_inv03 = 1;
    100: op1_01_inv03 = 1;
    101: op1_01_inv03 = 1;
    104: op1_01_inv03 = 1;
    107: op1_01_inv03 = 1;
    109: op1_01_inv03 = 1;
    38: op1_01_inv03 = 1;
    111: op1_01_inv03 = 1;
    113: op1_01_inv03 = 1;
    114: op1_01_inv03 = 1;
    115: op1_01_inv03 = 1;
    116: op1_01_inv03 = 1;
    118: op1_01_inv03 = 1;
    43: op1_01_inv03 = 1;
    120: op1_01_inv03 = 1;
    122: op1_01_inv03 = 1;
    124: op1_01_inv03 = 1;
    125: op1_01_inv03 = 1;
    126: op1_01_inv03 = 1;
    127: op1_01_inv03 = 1;
    129: op1_01_inv03 = 1;
    24: op1_01_inv03 = 1;
    default: op1_01_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の4番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in04 = reg_0018;
    52: op1_01_in04 = reg_0456;
    49: op1_01_in04 = reg_0623;
    53: op1_01_in04 = reg_0290;
    67: op1_01_in04 = reg_0375;
    61: op1_01_in04 = reg_0842;
    72: op1_01_in04 = reg_1079;
    71: op1_01_in04 = reg_1079;
    58: op1_01_in04 = reg_0245;
    68: op1_01_in04 = reg_0106;
    55: op1_01_in04 = imem04_in[7:4];
    73: op1_01_in04 = reg_0274;
    48: op1_01_in04 = reg_0283;
    86: op1_01_in04 = imem03_in[15:12];
    69: op1_01_in04 = reg_0350;
    59: op1_01_in04 = reg_0805;
    98: op1_01_in04 = reg_0805;
    50: op1_01_in04 = imem02_in[3:0];
    60: op1_01_in04 = reg_0256;
    33: op1_01_in04 = reg_0003;
    46: op1_01_in04 = reg_0104;
    74: op1_01_in04 = reg_0587;
    47: op1_01_in04 = reg_0213;
    75: op1_01_in04 = reg_0896;
    44: op1_01_in04 = reg_0117;
    56: op1_01_in04 = reg_0411;
    87: op1_01_in04 = reg_1233;
    40: op1_01_in04 = reg_0140;
    37: op1_01_in04 = imem07_in[11:8];
    108: op1_01_in04 = imem07_in[11:8];
    76: op1_01_in04 = reg_1490;
    57: op1_01_in04 = reg_0191;
    70: op1_01_in04 = reg_0127;
    77: op1_01_in04 = reg_0719;
    88: op1_01_in04 = reg_0535;
    34: op1_01_in04 = reg_0051;
    51: op1_01_in04 = reg_0408;
    78: op1_01_in04 = reg_0249;
    42: op1_01_in04 = reg_0241;
    79: op1_01_in04 = reg_1269;
    35: op1_01_in04 = reg_0384;
    62: op1_01_in04 = reg_0172;
    80: op1_01_in04 = reg_1081;
    81: op1_01_in04 = reg_0613;
    115: op1_01_in04 = reg_0613;
    89: op1_01_in04 = reg_1004;
    63: op1_01_in04 = reg_0715;
    82: op1_01_in04 = reg_1470;
    83: op1_01_in04 = reg_1493;
    39: op1_01_in04 = reg_0695;
    64: op1_01_in04 = reg_0605;
    84: op1_01_in04 = reg_1241;
    65: op1_01_in04 = reg_0126;
    85: op1_01_in04 = reg_0445;
    90: op1_01_in04 = reg_0433;
    66: op1_01_in04 = reg_1028;
    91: op1_01_in04 = reg_0294;
    92: op1_01_in04 = reg_0153;
    25: op1_01_in04 = reg_0103;
    93: op1_01_in04 = reg_1488;
    94: op1_01_in04 = reg_0111;
    95: op1_01_in04 = reg_0554;
    96: op1_01_in04 = reg_0198;
    120: op1_01_in04 = reg_0198;
    97: op1_01_in04 = reg_0965;
    99: op1_01_in04 = reg_0498;
    100: op1_01_in04 = reg_1071;
    101: op1_01_in04 = reg_1053;
    117: op1_01_in04 = reg_1053;
    102: op1_01_in04 = reg_1346;
    103: op1_01_in04 = reg_0663;
    104: op1_01_in04 = reg_1491;
    105: op1_01_in04 = reg_0291;
    106: op1_01_in04 = reg_0233;
    107: op1_01_in04 = reg_0347;
    27: op1_01_in04 = reg_0270;
    109: op1_01_in04 = reg_0236;
    110: op1_01_in04 = reg_1456;
    38: op1_01_in04 = reg_0050;
    111: op1_01_in04 = imem06_in[11:8];
    112: op1_01_in04 = reg_0659;
    113: op1_01_in04 = reg_0906;
    114: op1_01_in04 = reg_0107;
    116: op1_01_in04 = imem02_in[11:8];
    128: op1_01_in04 = imem02_in[11:8];
    118: op1_01_in04 = reg_0615;
    43: op1_01_in04 = reg_0337;
    119: op1_01_in04 = reg_1141;
    121: op1_01_in04 = reg_0131;
    122: op1_01_in04 = reg_1487;
    123: op1_01_in04 = reg_0266;
    124: op1_01_in04 = reg_1517;
    125: op1_01_in04 = reg_0804;
    126: op1_01_in04 = reg_0534;
    127: op1_01_in04 = reg_0748;
    129: op1_01_in04 = reg_0585;
    130: op1_01_in04 = reg_1453;
    131: op1_01_in04 = reg_0115;
    24: op1_01_in04 = reg_0001;
    default: op1_01_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv04 = 1;
    53: op1_01_inv04 = 1;
    58: op1_01_inv04 = 1;
    55: op1_01_inv04 = 1;
    59: op1_01_inv04 = 1;
    50: op1_01_inv04 = 1;
    33: op1_01_inv04 = 1;
    46: op1_01_inv04 = 1;
    47: op1_01_inv04 = 1;
    75: op1_01_inv04 = 1;
    44: op1_01_inv04 = 1;
    56: op1_01_inv04 = 1;
    76: op1_01_inv04 = 1;
    70: op1_01_inv04 = 1;
    77: op1_01_inv04 = 1;
    88: op1_01_inv04 = 1;
    34: op1_01_inv04 = 1;
    78: op1_01_inv04 = 1;
    42: op1_01_inv04 = 1;
    35: op1_01_inv04 = 1;
    89: op1_01_inv04 = 1;
    82: op1_01_inv04 = 1;
    83: op1_01_inv04 = 1;
    39: op1_01_inv04 = 1;
    64: op1_01_inv04 = 1;
    84: op1_01_inv04 = 1;
    90: op1_01_inv04 = 1;
    66: op1_01_inv04 = 1;
    92: op1_01_inv04 = 1;
    25: op1_01_inv04 = 1;
    94: op1_01_inv04 = 1;
    95: op1_01_inv04 = 1;
    98: op1_01_inv04 = 1;
    99: op1_01_inv04 = 1;
    102: op1_01_inv04 = 1;
    107: op1_01_inv04 = 1;
    108: op1_01_inv04 = 1;
    110: op1_01_inv04 = 1;
    116: op1_01_inv04 = 1;
    43: op1_01_inv04 = 1;
    121: op1_01_inv04 = 1;
    122: op1_01_inv04 = 1;
    124: op1_01_inv04 = 1;
    127: op1_01_inv04 = 1;
    129: op1_01_inv04 = 1;
    131: op1_01_inv04 = 1;
    24: op1_01_inv04 = 1;
    default: op1_01_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の5番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in05 = imem07_in[7:4];
    52: op1_01_in05 = reg_0989;
    49: op1_01_in05 = reg_0114;
    53: op1_01_in05 = reg_0291;
    67: op1_01_in05 = reg_0350;
    61: op1_01_in05 = reg_1242;
    85: op1_01_in05 = reg_1242;
    72: op1_01_in05 = reg_0842;
    71: op1_01_in05 = reg_0842;
    58: op1_01_in05 = reg_0673;
    86: op1_01_in05 = reg_0673;
    68: op1_01_in05 = reg_0390;
    55: op1_01_in05 = reg_1077;
    73: op1_01_in05 = reg_0393;
    48: op1_01_in05 = reg_0010;
    69: op1_01_in05 = reg_1325;
    59: op1_01_in05 = reg_1053;
    50: op1_01_in05 = reg_0922;
    60: op1_01_in05 = reg_0475;
    33: op1_01_in05 = reg_0053;
    46: op1_01_in05 = reg_0504;
    74: op1_01_in05 = reg_1299;
    47: op1_01_in05 = reg_0923;
    75: op1_01_in05 = reg_0874;
    44: op1_01_in05 = reg_0211;
    56: op1_01_in05 = reg_0463;
    87: op1_01_in05 = reg_0281;
    40: op1_01_in05 = reg_0779;
    37: op1_01_in05 = reg_0592;
    103: op1_01_in05 = reg_0592;
    76: op1_01_in05 = reg_0552;
    126: op1_01_in05 = reg_0552;
    57: op1_01_in05 = reg_1097;
    70: op1_01_in05 = reg_0382;
    77: op1_01_in05 = reg_0117;
    88: op1_01_in05 = reg_1339;
    34: op1_01_in05 = reg_0052;
    51: op1_01_in05 = reg_0415;
    78: op1_01_in05 = reg_0987;
    42: op1_01_in05 = reg_0746;
    79: op1_01_in05 = reg_0395;
    107: op1_01_in05 = reg_0395;
    35: op1_01_in05 = reg_0047;
    62: op1_01_in05 = reg_0136;
    66: op1_01_in05 = reg_0136;
    80: op1_01_in05 = reg_0580;
    81: op1_01_in05 = reg_0803;
    89: op1_01_in05 = reg_0342;
    63: op1_01_in05 = reg_0968;
    82: op1_01_in05 = reg_0523;
    83: op1_01_in05 = reg_0169;
    39: op1_01_in05 = reg_0595;
    64: op1_01_in05 = reg_0530;
    84: op1_01_in05 = reg_0841;
    115: op1_01_in05 = reg_0841;
    65: op1_01_in05 = reg_0106;
    90: op1_01_in05 = reg_1451;
    91: op1_01_in05 = reg_0217;
    92: op1_01_in05 = reg_1405;
    25: op1_01_in05 = reg_0321;
    93: op1_01_in05 = reg_0035;
    94: op1_01_in05 = reg_0878;
    95: op1_01_in05 = reg_0640;
    96: op1_01_in05 = reg_0783;
    97: op1_01_in05 = reg_1184;
    98: op1_01_in05 = reg_0554;
    99: op1_01_in05 = reg_1414;
    100: op1_01_in05 = imem02_in[3:0];
    101: op1_01_in05 = reg_1227;
    130: op1_01_in05 = reg_1227;
    102: op1_01_in05 = reg_0799;
    104: op1_01_in05 = reg_0805;
    105: op1_01_in05 = reg_1139;
    106: op1_01_in05 = reg_0699;
    27: op1_01_in05 = reg_0023;
    108: op1_01_in05 = reg_0478;
    109: op1_01_in05 = reg_1503;
    110: op1_01_in05 = reg_0147;
    38: op1_01_in05 = reg_0051;
    111: op1_01_in05 = reg_1058;
    112: op1_01_in05 = reg_0666;
    113: op1_01_in05 = reg_0397;
    114: op1_01_in05 = reg_0880;
    116: op1_01_in05 = reg_0889;
    117: op1_01_in05 = reg_0440;
    118: op1_01_in05 = reg_1028;
    43: op1_01_in05 = reg_0065;
    119: op1_01_in05 = reg_0804;
    120: op1_01_in05 = reg_1001;
    121: op1_01_in05 = reg_0939;
    122: op1_01_in05 = reg_1491;
    123: op1_01_in05 = reg_1514;
    124: op1_01_in05 = reg_1313;
    125: op1_01_in05 = reg_1205;
    127: op1_01_in05 = reg_1490;
    128: op1_01_in05 = reg_0327;
    129: op1_01_in05 = reg_0373;
    131: op1_01_in05 = reg_0116;
    24: op1_01_in05 = reg_0084;
    default: op1_01_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_01_inv05 = 1;
    67: op1_01_inv05 = 1;
    61: op1_01_inv05 = 1;
    68: op1_01_inv05 = 1;
    73: op1_01_inv05 = 1;
    71: op1_01_inv05 = 1;
    60: op1_01_inv05 = 1;
    46: op1_01_inv05 = 1;
    74: op1_01_inv05 = 1;
    47: op1_01_inv05 = 1;
    44: op1_01_inv05 = 1;
    56: op1_01_inv05 = 1;
    37: op1_01_inv05 = 1;
    76: op1_01_inv05 = 1;
    57: op1_01_inv05 = 1;
    51: op1_01_inv05 = 1;
    78: op1_01_inv05 = 1;
    42: op1_01_inv05 = 1;
    35: op1_01_inv05 = 1;
    81: op1_01_inv05 = 1;
    89: op1_01_inv05 = 1;
    63: op1_01_inv05 = 1;
    83: op1_01_inv05 = 1;
    90: op1_01_inv05 = 1;
    91: op1_01_inv05 = 1;
    25: op1_01_inv05 = 1;
    93: op1_01_inv05 = 1;
    94: op1_01_inv05 = 1;
    95: op1_01_inv05 = 1;
    98: op1_01_inv05 = 1;
    101: op1_01_inv05 = 1;
    103: op1_01_inv05 = 1;
    104: op1_01_inv05 = 1;
    27: op1_01_inv05 = 1;
    108: op1_01_inv05 = 1;
    109: op1_01_inv05 = 1;
    113: op1_01_inv05 = 1;
    115: op1_01_inv05 = 1;
    116: op1_01_inv05 = 1;
    118: op1_01_inv05 = 1;
    119: op1_01_inv05 = 1;
    122: op1_01_inv05 = 1;
    125: op1_01_inv05 = 1;
    127: op1_01_inv05 = 1;
    129: op1_01_inv05 = 1;
    130: op1_01_inv05 = 1;
    24: op1_01_inv05 = 1;
    default: op1_01_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の6番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in06 = reg_0228;
    25: op1_01_in06 = reg_0228;
    52: op1_01_in06 = reg_0970;
    49: op1_01_in06 = reg_0520;
    53: op1_01_in06 = reg_0044;
    67: op1_01_in06 = reg_0638;
    61: op1_01_in06 = reg_1053;
    72: op1_01_in06 = imem00_in[3:0];
    71: op1_01_in06 = imem00_in[3:0];
    58: op1_01_in06 = reg_0158;
    68: op1_01_in06 = reg_0055;
    112: op1_01_in06 = reg_0055;
    55: op1_01_in06 = reg_0420;
    73: op1_01_in06 = reg_0828;
    48: op1_01_in06 = reg_0553;
    86: op1_01_in06 = reg_0288;
    69: op1_01_in06 = reg_0180;
    59: op1_01_in06 = reg_0155;
    50: op1_01_in06 = reg_0589;
    60: op1_01_in06 = reg_0474;
    33: op1_01_in06 = reg_0518;
    46: op1_01_in06 = reg_0574;
    74: op1_01_in06 = reg_0204;
    47: op1_01_in06 = imem07_in[11:8];
    57: op1_01_in06 = imem07_in[11:8];
    75: op1_01_in06 = reg_0079;
    44: op1_01_in06 = reg_0016;
    56: op1_01_in06 = reg_0464;
    87: op1_01_in06 = reg_0454;
    40: op1_01_in06 = reg_0286;
    37: op1_01_in06 = reg_0100;
    76: op1_01_in06 = reg_1469;
    70: op1_01_in06 = reg_0056;
    77: op1_01_in06 = reg_0021;
    43: op1_01_in06 = reg_0021;
    88: op1_01_in06 = reg_1340;
    34: op1_01_in06 = reg_0084;
    51: op1_01_in06 = reg_0623;
    78: op1_01_in06 = reg_0460;
    42: op1_01_in06 = reg_0726;
    79: op1_01_in06 = reg_0646;
    35: op1_01_in06 = reg_0291;
    62: op1_01_in06 = reg_1227;
    95: op1_01_in06 = reg_1227;
    80: op1_01_in06 = reg_0806;
    81: op1_01_in06 = reg_1027;
    89: op1_01_in06 = reg_0304;
    63: op1_01_in06 = reg_0438;
    82: op1_01_in06 = reg_0250;
    83: op1_01_in06 = reg_0276;
    39: op1_01_in06 = reg_0596;
    64: op1_01_in06 = reg_0455;
    84: op1_01_in06 = reg_0459;
    65: op1_01_in06 = reg_0897;
    85: op1_01_in06 = reg_0580;
    90: op1_01_in06 = reg_0128;
    66: op1_01_in06 = reg_0249;
    101: op1_01_in06 = reg_0249;
    91: op1_01_in06 = imem03_in[3:0];
    92: op1_01_in06 = reg_0202;
    93: op1_01_in06 = imem05_in[7:4];
    94: op1_01_in06 = reg_0380;
    96: op1_01_in06 = reg_0556;
    97: op1_01_in06 = reg_0142;
    98: op1_01_in06 = reg_1052;
    99: op1_01_in06 = reg_0461;
    100: op1_01_in06 = reg_0668;
    102: op1_01_in06 = reg_0151;
    103: op1_01_in06 = reg_0103;
    104: op1_01_in06 = reg_0555;
    105: op1_01_in06 = reg_0348;
    106: op1_01_in06 = reg_0732;
    107: op1_01_in06 = reg_0272;
    27: op1_01_in06 = reg_0015;
    108: op1_01_in06 = reg_1315;
    109: op1_01_in06 = imem05_in[15:12];
    110: op1_01_in06 = reg_1511;
    38: op1_01_in06 = reg_0003;
    111: op1_01_in06 = reg_0270;
    113: op1_01_in06 = reg_1326;
    114: op1_01_in06 = reg_0707;
    115: op1_01_in06 = reg_0615;
    116: op1_01_in06 = reg_0322;
    117: op1_01_in06 = reg_0416;
    118: op1_01_in06 = reg_1230;
    119: op1_01_in06 = reg_0805;
    120: op1_01_in06 = reg_0783;
    121: op1_01_in06 = reg_0266;
    122: op1_01_in06 = reg_0613;
    123: op1_01_in06 = reg_0303;
    124: op1_01_in06 = reg_0756;
    125: op1_01_in06 = reg_1405;
    126: op1_01_in06 = reg_1203;
    127: op1_01_in06 = reg_1489;
    128: op1_01_in06 = reg_0879;
    129: op1_01_in06 = reg_0527;
    130: op1_01_in06 = reg_1205;
    131: op1_01_in06 = reg_0109;
    24: op1_01_in06 = reg_0053;
    default: op1_01_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv06 = 1;
    53: op1_01_inv06 = 1;
    61: op1_01_inv06 = 1;
    72: op1_01_inv06 = 1;
    58: op1_01_inv06 = 1;
    68: op1_01_inv06 = 1;
    55: op1_01_inv06 = 1;
    73: op1_01_inv06 = 1;
    71: op1_01_inv06 = 1;
    48: op1_01_inv06 = 1;
    86: op1_01_inv06 = 1;
    69: op1_01_inv06 = 1;
    59: op1_01_inv06 = 1;
    60: op1_01_inv06 = 1;
    33: op1_01_inv06 = 1;
    46: op1_01_inv06 = 1;
    74: op1_01_inv06 = 1;
    47: op1_01_inv06 = 1;
    75: op1_01_inv06 = 1;
    57: op1_01_inv06 = 1;
    34: op1_01_inv06 = 1;
    51: op1_01_inv06 = 1;
    78: op1_01_inv06 = 1;
    42: op1_01_inv06 = 1;
    89: op1_01_inv06 = 1;
    63: op1_01_inv06 = 1;
    82: op1_01_inv06 = 1;
    39: op1_01_inv06 = 1;
    64: op1_01_inv06 = 1;
    84: op1_01_inv06 = 1;
    85: op1_01_inv06 = 1;
    25: op1_01_inv06 = 1;
    96: op1_01_inv06 = 1;
    98: op1_01_inv06 = 1;
    99: op1_01_inv06 = 1;
    100: op1_01_inv06 = 1;
    103: op1_01_inv06 = 1;
    104: op1_01_inv06 = 1;
    105: op1_01_inv06 = 1;
    106: op1_01_inv06 = 1;
    27: op1_01_inv06 = 1;
    108: op1_01_inv06 = 1;
    109: op1_01_inv06 = 1;
    112: op1_01_inv06 = 1;
    113: op1_01_inv06 = 1;
    116: op1_01_inv06 = 1;
    117: op1_01_inv06 = 1;
    120: op1_01_inv06 = 1;
    121: op1_01_inv06 = 1;
    122: op1_01_inv06 = 1;
    123: op1_01_inv06 = 1;
    125: op1_01_inv06 = 1;
    127: op1_01_inv06 = 1;
    129: op1_01_inv06 = 1;
    default: op1_01_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の7番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in07 = reg_0223;
    52: op1_01_in07 = reg_0971;
    49: op1_01_in07 = reg_0123;
    53: op1_01_in07 = reg_0041;
    67: op1_01_in07 = reg_0234;
    61: op1_01_in07 = reg_1027;
    104: op1_01_in07 = reg_1027;
    72: op1_01_in07 = reg_0805;
    58: op1_01_in07 = reg_0791;
    68: op1_01_in07 = reg_0711;
    55: op1_01_in07 = reg_0421;
    73: op1_01_in07 = reg_0206;
    71: op1_01_in07 = reg_0293;
    85: op1_01_in07 = reg_0293;
    48: op1_01_in07 = imem02_in[3:0];
    86: op1_01_in07 = reg_1282;
    114: op1_01_in07 = reg_1282;
    69: op1_01_in07 = reg_0964;
    59: op1_01_in07 = reg_0249;
    95: op1_01_in07 = reg_0249;
    50: op1_01_in07 = reg_0563;
    60: op1_01_in07 = reg_0933;
    33: op1_01_in07 = reg_0520;
    46: op1_01_in07 = reg_0537;
    74: op1_01_in07 = reg_1298;
    47: op1_01_in07 = reg_0225;
    75: op1_01_in07 = reg_0043;
    44: op1_01_in07 = reg_0578;
    56: op1_01_in07 = reg_1198;
    87: op1_01_in07 = reg_0932;
    40: op1_01_in07 = reg_0366;
    37: op1_01_in07 = reg_0114;
    76: op1_01_in07 = reg_0523;
    98: op1_01_in07 = reg_0523;
    57: op1_01_in07 = reg_0668;
    70: op1_01_in07 = reg_0708;
    77: op1_01_in07 = reg_0470;
    88: op1_01_in07 = reg_1338;
    34: op1_01_in07 = reg_0087;
    51: op1_01_in07 = reg_0591;
    78: op1_01_in07 = reg_1417;
    81: op1_01_in07 = reg_1417;
    42: op1_01_in07 = reg_0727;
    79: op1_01_in07 = reg_0565;
    35: op1_01_in07 = reg_0282;
    62: op1_01_in07 = reg_0725;
    80: op1_01_in07 = reg_1471;
    89: op1_01_in07 = reg_0338;
    63: op1_01_in07 = reg_0726;
    82: op1_01_in07 = reg_1028;
    83: op1_01_in07 = reg_0055;
    39: op1_01_in07 = reg_0368;
    64: op1_01_in07 = reg_0560;
    84: op1_01_in07 = reg_0928;
    65: op1_01_in07 = reg_0294;
    90: op1_01_in07 = reg_1433;
    66: op1_01_in07 = reg_0459;
    91: op1_01_in07 = reg_0506;
    92: op1_01_in07 = reg_0352;
    25: op1_01_in07 = reg_0186;
    93: op1_01_in07 = reg_0315;
    94: op1_01_in07 = reg_0473;
    96: op1_01_in07 = reg_0965;
    97: op1_01_in07 = reg_1313;
    99: op1_01_in07 = reg_0478;
    100: op1_01_in07 = reg_0455;
    101: op1_01_in07 = reg_1229;
    102: op1_01_in07 = reg_0861;
    103: op1_01_in07 = reg_0051;
    105: op1_01_in07 = reg_0427;
    106: op1_01_in07 = reg_1145;
    107: op1_01_in07 = reg_0205;
    27: op1_01_in07 = reg_0252;
    108: op1_01_in07 = reg_1056;
    109: op1_01_in07 = reg_1430;
    110: op1_01_in07 = reg_0385;
    38: op1_01_in07 = reg_0085;
    111: op1_01_in07 = reg_0870;
    112: op1_01_in07 = reg_0532;
    113: op1_01_in07 = reg_0863;
    115: op1_01_in07 = reg_1053;
    116: op1_01_in07 = reg_1235;
    117: op1_01_in07 = reg_0405;
    118: op1_01_in07 = reg_0987;
    43: op1_01_in07 = reg_0032;
    119: op1_01_in07 = reg_1052;
    120: op1_01_in07 = reg_0312;
    121: op1_01_in07 = reg_1169;
    122: op1_01_in07 = reg_0615;
    123: op1_01_in07 = reg_0736;
    124: op1_01_in07 = reg_0558;
    125: op1_01_in07 = reg_0881;
    126: op1_01_in07 = reg_1215;
    127: op1_01_in07 = reg_0803;
    128: op1_01_in07 = reg_0608;
    129: op1_01_in07 = reg_0570;
    130: op1_01_in07 = reg_1206;
    131: op1_01_in07 = reg_0718;
    default: op1_01_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv07 = 1;
    52: op1_01_inv07 = 1;
    49: op1_01_inv07 = 1;
    61: op1_01_inv07 = 1;
    58: op1_01_inv07 = 1;
    86: op1_01_inv07 = 1;
    59: op1_01_inv07 = 1;
    60: op1_01_inv07 = 1;
    46: op1_01_inv07 = 1;
    74: op1_01_inv07 = 1;
    47: op1_01_inv07 = 1;
    75: op1_01_inv07 = 1;
    56: op1_01_inv07 = 1;
    87: op1_01_inv07 = 1;
    40: op1_01_inv07 = 1;
    76: op1_01_inv07 = 1;
    57: op1_01_inv07 = 1;
    34: op1_01_inv07 = 1;
    51: op1_01_inv07 = 1;
    78: op1_01_inv07 = 1;
    35: op1_01_inv07 = 1;
    62: op1_01_inv07 = 1;
    80: op1_01_inv07 = 1;
    81: op1_01_inv07 = 1;
    89: op1_01_inv07 = 1;
    83: op1_01_inv07 = 1;
    64: op1_01_inv07 = 1;
    65: op1_01_inv07 = 1;
    66: op1_01_inv07 = 1;
    91: op1_01_inv07 = 1;
    92: op1_01_inv07 = 1;
    95: op1_01_inv07 = 1;
    96: op1_01_inv07 = 1;
    97: op1_01_inv07 = 1;
    98: op1_01_inv07 = 1;
    102: op1_01_inv07 = 1;
    105: op1_01_inv07 = 1;
    106: op1_01_inv07 = 1;
    107: op1_01_inv07 = 1;
    108: op1_01_inv07 = 1;
    109: op1_01_inv07 = 1;
    110: op1_01_inv07 = 1;
    38: op1_01_inv07 = 1;
    111: op1_01_inv07 = 1;
    117: op1_01_inv07 = 1;
    118: op1_01_inv07 = 1;
    43: op1_01_inv07 = 1;
    121: op1_01_inv07 = 1;
    122: op1_01_inv07 = 1;
    126: op1_01_inv07 = 1;
    127: op1_01_inv07 = 1;
    128: op1_01_inv07 = 1;
    131: op1_01_inv07 = 1;
    default: op1_01_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の8番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in08 = reg_0225;
    108: op1_01_in08 = reg_0225;
    52: op1_01_in08 = reg_0626;
    53: op1_01_in08 = reg_0446;
    67: op1_01_in08 = reg_0180;
    61: op1_01_in08 = reg_0460;
    72: op1_01_in08 = reg_0961;
    66: op1_01_in08 = reg_0961;
    58: op1_01_in08 = reg_0140;
    68: op1_01_in08 = reg_0306;
    55: op1_01_in08 = reg_0414;
    73: op1_01_in08 = reg_0458;
    71: op1_01_in08 = reg_1229;
    48: op1_01_in08 = imem02_in[11:8];
    86: op1_01_in08 = reg_0426;
    69: op1_01_in08 = reg_0190;
    59: op1_01_in08 = reg_1205;
    85: op1_01_in08 = reg_1205;
    50: op1_01_in08 = reg_0561;
    60: op1_01_in08 = reg_0380;
    33: op1_01_in08 = reg_0124;
    46: op1_01_in08 = reg_0534;
    74: op1_01_in08 = reg_0877;
    47: op1_01_in08 = reg_0893;
    75: op1_01_in08 = reg_0744;
    44: op1_01_in08 = reg_0393;
    56: op1_01_in08 = reg_0466;
    87: op1_01_in08 = reg_0064;
    40: op1_01_in08 = reg_0623;
    37: op1_01_in08 = reg_0321;
    76: op1_01_in08 = reg_1028;
    98: op1_01_in08 = reg_1028;
    57: op1_01_in08 = reg_0224;
    70: op1_01_in08 = reg_0279;
    77: op1_01_in08 = reg_0587;
    88: op1_01_in08 = reg_0297;
    34: op1_01_in08 = reg_0519;
    51: op1_01_in08 = reg_0001;
    78: op1_01_in08 = reg_0722;
    42: op1_01_in08 = reg_0439;
    79: op1_01_in08 = reg_0938;
    35: op1_01_in08 = reg_0044;
    62: op1_01_in08 = reg_0435;
    80: op1_01_in08 = reg_1469;
    81: op1_01_in08 = reg_0881;
    89: op1_01_in08 = reg_1488;
    63: op1_01_in08 = reg_0147;
    82: op1_01_in08 = reg_1027;
    83: op1_01_in08 = reg_0390;
    39: op1_01_in08 = reg_0304;
    64: op1_01_in08 = reg_1343;
    84: op1_01_in08 = reg_0883;
    65: op1_01_in08 = reg_0009;
    90: op1_01_in08 = reg_1032;
    91: op1_01_in08 = reg_0840;
    92: op1_01_in08 = reg_0387;
    25: op1_01_in08 = reg_0002;
    93: op1_01_in08 = reg_0204;
    94: op1_01_in08 = reg_0007;
    95: op1_01_in08 = reg_1230;
    96: op1_01_in08 = reg_1184;
    97: op1_01_in08 = reg_0048;
    99: op1_01_in08 = reg_0219;
    100: op1_01_in08 = reg_0588;
    101: op1_01_in08 = reg_1432;
    102: op1_01_in08 = reg_0207;
    103: op1_01_in08 = reg_0004;
    104: op1_01_in08 = reg_1454;
    105: op1_01_in08 = imem04_in[7:4];
    106: op1_01_in08 = reg_0330;
    107: op1_01_in08 = reg_1164;
    27: op1_01_in08 = reg_0230;
    109: op1_01_in08 = reg_0996;
    110: op1_01_in08 = reg_0362;
    38: op1_01_in08 = reg_0084;
    111: op1_01_in08 = reg_1420;
    112: op1_01_in08 = reg_0898;
    113: op1_01_in08 = reg_0717;
    114: op1_01_in08 = imem04_in[15:12];
    115: op1_01_in08 = reg_0293;
    116: op1_01_in08 = reg_0056;
    117: op1_01_in08 = reg_0122;
    118: op1_01_in08 = reg_1206;
    43: op1_01_in08 = reg_0391;
    119: op1_01_in08 = reg_0250;
    120: op1_01_in08 = reg_1494;
    121: op1_01_in08 = reg_0090;
    122: op1_01_in08 = reg_0486;
    123: op1_01_in08 = reg_0275;
    124: op1_01_in08 = reg_1093;
    125: op1_01_in08 = reg_0887;
    126: op1_01_in08 = reg_1233;
    127: op1_01_in08 = reg_1102;
    128: op1_01_in08 = reg_0975;
    129: op1_01_in08 = reg_1228;
    130: op1_01_in08 = reg_0524;
    131: op1_01_in08 = reg_0636;
    default: op1_01_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv08 = 1;
    53: op1_01_inv08 = 1;
    67: op1_01_inv08 = 1;
    61: op1_01_inv08 = 1;
    58: op1_01_inv08 = 1;
    68: op1_01_inv08 = 1;
    71: op1_01_inv08 = 1;
    59: op1_01_inv08 = 1;
    60: op1_01_inv08 = 1;
    74: op1_01_inv08 = 1;
    56: op1_01_inv08 = 1;
    40: op1_01_inv08 = 1;
    76: op1_01_inv08 = 1;
    57: op1_01_inv08 = 1;
    70: op1_01_inv08 = 1;
    34: op1_01_inv08 = 1;
    51: op1_01_inv08 = 1;
    78: op1_01_inv08 = 1;
    35: op1_01_inv08 = 1;
    89: op1_01_inv08 = 1;
    63: op1_01_inv08 = 1;
    82: op1_01_inv08 = 1;
    65: op1_01_inv08 = 1;
    85: op1_01_inv08 = 1;
    90: op1_01_inv08 = 1;
    93: op1_01_inv08 = 1;
    95: op1_01_inv08 = 1;
    98: op1_01_inv08 = 1;
    99: op1_01_inv08 = 1;
    101: op1_01_inv08 = 1;
    104: op1_01_inv08 = 1;
    105: op1_01_inv08 = 1;
    107: op1_01_inv08 = 1;
    108: op1_01_inv08 = 1;
    110: op1_01_inv08 = 1;
    111: op1_01_inv08 = 1;
    112: op1_01_inv08 = 1;
    113: op1_01_inv08 = 1;
    114: op1_01_inv08 = 1;
    118: op1_01_inv08 = 1;
    119: op1_01_inv08 = 1;
    121: op1_01_inv08 = 1;
    122: op1_01_inv08 = 1;
    123: op1_01_inv08 = 1;
    125: op1_01_inv08 = 1;
    127: op1_01_inv08 = 1;
    130: op1_01_inv08 = 1;
    default: op1_01_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の9番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in09 = reg_0198;
    52: op1_01_in09 = reg_0055;
    53: op1_01_in09 = reg_0662;
    67: op1_01_in09 = reg_0789;
    61: op1_01_in09 = reg_0409;
    72: op1_01_in09 = reg_1432;
    58: op1_01_in09 = reg_0775;
    68: op1_01_in09 = reg_0630;
    55: op1_01_in09 = reg_0412;
    73: op1_01_in09 = reg_0751;
    71: op1_01_in09 = reg_0987;
    48: op1_01_in09 = reg_0563;
    86: op1_01_in09 = reg_0411;
    69: op1_01_in09 = reg_0597;
    59: op1_01_in09 = reg_0459;
    101: op1_01_in09 = reg_0459;
    50: op1_01_in09 = reg_0532;
    60: op1_01_in09 = reg_0381;
    46: op1_01_in09 = reg_0463;
    74: op1_01_in09 = reg_0733;
    47: op1_01_in09 = reg_0170;
    75: op1_01_in09 = reg_0456;
    44: op1_01_in09 = reg_0745;
    56: op1_01_in09 = reg_0467;
    87: op1_01_in09 = reg_0095;
    40: op1_01_in09 = reg_0618;
    37: op1_01_in09 = reg_0050;
    76: op1_01_in09 = reg_0221;
    82: op1_01_in09 = reg_0221;
    57: op1_01_in09 = reg_0704;
    70: op1_01_in09 = reg_0311;
    77: op1_01_in09 = reg_1430;
    88: op1_01_in09 = reg_1203;
    34: op1_01_in09 = reg_0124;
    78: op1_01_in09 = reg_0388;
    42: op1_01_in09 = reg_0434;
    79: op1_01_in09 = reg_0318;
    35: op1_01_in09 = reg_0012;
    62: op1_01_in09 = reg_0387;
    80: op1_01_in09 = reg_1470;
    81: op1_01_in09 = reg_0887;
    89: op1_01_in09 = reg_0736;
    121: op1_01_in09 = reg_0736;
    63: op1_01_in09 = reg_0148;
    83: op1_01_in09 = reg_0473;
    39: op1_01_in09 = reg_0262;
    64: op1_01_in09 = reg_0256;
    84: op1_01_in09 = reg_0722;
    65: op1_01_in09 = reg_0024;
    85: op1_01_in09 = reg_0229;
    90: op1_01_in09 = reg_0380;
    66: op1_01_in09 = reg_0352;
    91: op1_01_in09 = reg_0759;
    92: op1_01_in09 = reg_0389;
    25: op1_01_in09 = reg_0004;
    93: op1_01_in09 = reg_0205;
    94: op1_01_in09 = reg_1392;
    95: op1_01_in09 = reg_1406;
    130: op1_01_in09 = reg_1406;
    96: op1_01_in09 = reg_0957;
    97: op1_01_in09 = reg_1093;
    98: op1_01_in09 = reg_1027;
    122: op1_01_in09 = reg_1027;
    99: op1_01_in09 = reg_0703;
    100: op1_01_in09 = reg_0839;
    128: op1_01_in09 = reg_0839;
    102: op1_01_in09 = imem06_in[3:0];
    104: op1_01_in09 = reg_1227;
    105: op1_01_in09 = reg_0032;
    114: op1_01_in09 = reg_0032;
    106: op1_01_in09 = reg_1448;
    107: op1_01_in09 = reg_0648;
    27: op1_01_in09 = reg_0231;
    108: op1_01_in09 = reg_0457;
    109: op1_01_in09 = reg_0649;
    110: op1_01_in09 = reg_0464;
    38: op1_01_in09 = reg_0520;
    111: op1_01_in09 = reg_0696;
    112: op1_01_in09 = reg_0495;
    113: op1_01_in09 = reg_0636;
    115: op1_01_in09 = reg_0485;
    116: op1_01_in09 = reg_0900;
    117: op1_01_in09 = reg_0917;
    118: op1_01_in09 = reg_0460;
    43: op1_01_in09 = reg_0748;
    119: op1_01_in09 = reg_0293;
    120: op1_01_in09 = reg_1184;
    123: op1_01_in09 = reg_0393;
    124: op1_01_in09 = reg_1208;
    125: op1_01_in09 = reg_0883;
    126: op1_01_in09 = reg_0407;
    127: op1_01_in09 = reg_0616;
    129: op1_01_in09 = reg_0419;
    131: op1_01_in09 = reg_0141;
    default: op1_01_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_01_inv09 = 1;
    61: op1_01_inv09 = 1;
    55: op1_01_inv09 = 1;
    73: op1_01_inv09 = 1;
    71: op1_01_inv09 = 1;
    48: op1_01_inv09 = 1;
    86: op1_01_inv09 = 1;
    69: op1_01_inv09 = 1;
    50: op1_01_inv09 = 1;
    46: op1_01_inv09 = 1;
    47: op1_01_inv09 = 1;
    75: op1_01_inv09 = 1;
    87: op1_01_inv09 = 1;
    37: op1_01_inv09 = 1;
    57: op1_01_inv09 = 1;
    77: op1_01_inv09 = 1;
    88: op1_01_inv09 = 1;
    34: op1_01_inv09 = 1;
    42: op1_01_inv09 = 1;
    79: op1_01_inv09 = 1;
    35: op1_01_inv09 = 1;
    62: op1_01_inv09 = 1;
    81: op1_01_inv09 = 1;
    89: op1_01_inv09 = 1;
    39: op1_01_inv09 = 1;
    64: op1_01_inv09 = 1;
    84: op1_01_inv09 = 1;
    65: op1_01_inv09 = 1;
    66: op1_01_inv09 = 1;
    91: op1_01_inv09 = 1;
    93: op1_01_inv09 = 1;
    94: op1_01_inv09 = 1;
    97: op1_01_inv09 = 1;
    105: op1_01_inv09 = 1;
    27: op1_01_inv09 = 1;
    109: op1_01_inv09 = 1;
    110: op1_01_inv09 = 1;
    111: op1_01_inv09 = 1;
    113: op1_01_inv09 = 1;
    114: op1_01_inv09 = 1;
    115: op1_01_inv09 = 1;
    116: op1_01_inv09 = 1;
    43: op1_01_inv09 = 1;
    121: op1_01_inv09 = 1;
    122: op1_01_inv09 = 1;
    126: op1_01_inv09 = 1;
    127: op1_01_inv09 = 1;
    129: op1_01_inv09 = 1;
    default: op1_01_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の10番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in10 = reg_0187;
    52: op1_01_in10 = reg_0897;
    53: op1_01_in10 = reg_0629;
    67: op1_01_in10 = reg_0261;
    61: op1_01_in10 = reg_0388;
    72: op1_01_in10 = reg_0459;
    58: op1_01_in10 = reg_0665;
    68: op1_01_in10 = reg_0191;
    55: op1_01_in10 = reg_0598;
    73: op1_01_in10 = reg_1105;
    71: op1_01_in10 = reg_0155;
    48: op1_01_in10 = reg_0532;
    86: op1_01_in10 = reg_0898;
    69: op1_01_in10 = reg_1301;
    59: op1_01_in10 = reg_0928;
    85: op1_01_in10 = reg_0928;
    50: op1_01_in10 = reg_0495;
    60: op1_01_in10 = reg_0153;
    46: op1_01_in10 = reg_0406;
    74: op1_01_in10 = reg_0347;
    47: op1_01_in10 = reg_0186;
    75: op1_01_in10 = reg_1344;
    44: op1_01_in10 = reg_0344;
    56: op1_01_in10 = reg_0798;
    87: op1_01_in10 = reg_0420;
    40: op1_01_in10 = reg_0137;
    37: op1_01_in10 = reg_0051;
    76: op1_01_in10 = reg_0249;
    57: op1_01_in10 = reg_0310;
    70: op1_01_in10 = reg_0313;
    77: op1_01_in10 = reg_0833;
    88: op1_01_in10 = reg_1200;
    78: op1_01_in10 = reg_0026;
    42: op1_01_in10 = reg_0162;
    79: op1_01_in10 = reg_0631;
    35: op1_01_in10 = reg_0662;
    62: op1_01_in10 = reg_0122;
    80: op1_01_in10 = reg_0250;
    81: op1_01_in10 = reg_0351;
    89: op1_01_in10 = reg_0205;
    63: op1_01_in10 = reg_0403;
    82: op1_01_in10 = reg_1454;
    119: op1_01_in10 = reg_1454;
    83: op1_01_in10 = reg_0474;
    39: op1_01_in10 = reg_0094;
    64: op1_01_in10 = reg_0972;
    84: op1_01_in10 = reg_0416;
    65: op1_01_in10 = reg_0068;
    90: op1_01_in10 = reg_0379;
    66: op1_01_in10 = reg_0201;
    91: op1_01_in10 = reg_0185;
    92: op1_01_in10 = reg_0059;
    93: op1_01_in10 = reg_1268;
    94: op1_01_in10 = imem03_in[7:4];
    95: op1_01_in10 = reg_0821;
    96: op1_01_in10 = reg_0108;
    97: op1_01_in10 = reg_0378;
    98: op1_01_in10 = reg_1459;
    99: op1_01_in10 = reg_0225;
    100: op1_01_in10 = reg_0497;
    101: op1_01_in10 = reg_0524;
    104: op1_01_in10 = reg_0524;
    102: op1_01_in10 = reg_0161;
    105: op1_01_in10 = reg_1369;
    106: op1_01_in10 = reg_0311;
    107: op1_01_in10 = reg_0562;
    109: op1_01_in10 = reg_0562;
    27: op1_01_in10 = reg_0246;
    108: op1_01_in10 = reg_0923;
    110: op1_01_in10 = reg_0079;
    111: op1_01_in10 = reg_0984;
    112: op1_01_in10 = reg_0973;
    113: op1_01_in10 = reg_0570;
    114: op1_01_in10 = reg_0129;
    115: op1_01_in10 = reg_1201;
    116: op1_01_in10 = reg_1207;
    117: op1_01_in10 = reg_0723;
    118: op1_01_in10 = reg_1417;
    43: op1_01_in10 = reg_0702;
    120: op1_01_in10 = reg_1518;
    121: op1_01_in10 = reg_0888;
    122: op1_01_in10 = reg_0485;
    123: op1_01_in10 = reg_0602;
    124: op1_01_in10 = reg_0104;
    125: op1_01_in10 = reg_0352;
    126: op1_01_in10 = reg_0969;
    127: op1_01_in10 = reg_0805;
    128: op1_01_in10 = reg_0900;
    129: op1_01_in10 = reg_0165;
    130: op1_01_in10 = reg_1393;
    131: op1_01_in10 = reg_0586;
    default: op1_01_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv10 = 1;
    67: op1_01_inv10 = 1;
    55: op1_01_inv10 = 1;
    73: op1_01_inv10 = 1;
    71: op1_01_inv10 = 1;
    86: op1_01_inv10 = 1;
    60: op1_01_inv10 = 1;
    47: op1_01_inv10 = 1;
    44: op1_01_inv10 = 1;
    56: op1_01_inv10 = 1;
    87: op1_01_inv10 = 1;
    40: op1_01_inv10 = 1;
    76: op1_01_inv10 = 1;
    78: op1_01_inv10 = 1;
    79: op1_01_inv10 = 1;
    62: op1_01_inv10 = 1;
    80: op1_01_inv10 = 1;
    81: op1_01_inv10 = 1;
    63: op1_01_inv10 = 1;
    84: op1_01_inv10 = 1;
    85: op1_01_inv10 = 1;
    90: op1_01_inv10 = 1;
    91: op1_01_inv10 = 1;
    93: op1_01_inv10 = 1;
    95: op1_01_inv10 = 1;
    96: op1_01_inv10 = 1;
    98: op1_01_inv10 = 1;
    100: op1_01_inv10 = 1;
    101: op1_01_inv10 = 1;
    104: op1_01_inv10 = 1;
    107: op1_01_inv10 = 1;
    110: op1_01_inv10 = 1;
    111: op1_01_inv10 = 1;
    116: op1_01_inv10 = 1;
    117: op1_01_inv10 = 1;
    118: op1_01_inv10 = 1;
    122: op1_01_inv10 = 1;
    123: op1_01_inv10 = 1;
    124: op1_01_inv10 = 1;
    126: op1_01_inv10 = 1;
    127: op1_01_inv10 = 1;
    128: op1_01_inv10 = 1;
    129: op1_01_inv10 = 1;
    130: op1_01_inv10 = 1;
    default: op1_01_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の11番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in11 = reg_0170;
    27: op1_01_in11 = reg_0170;
    52: op1_01_in11 = reg_0900;
    53: op1_01_in11 = reg_0922;
    67: op1_01_in11 = reg_1314;
    61: op1_01_in11 = reg_0350;
    124: op1_01_in11 = reg_0350;
    72: op1_01_in11 = reg_0821;
    101: op1_01_in11 = reg_0821;
    58: op1_01_in11 = reg_0285;
    68: op1_01_in11 = reg_0198;
    55: op1_01_in11 = reg_0454;
    73: op1_01_in11 = reg_0780;
    71: op1_01_in11 = reg_1405;
    48: op1_01_in11 = reg_0533;
    86: op1_01_in11 = reg_0696;
    69: op1_01_in11 = reg_0178;
    59: op1_01_in11 = reg_0188;
    50: op1_01_in11 = reg_0473;
    60: op1_01_in11 = reg_0306;
    46: op1_01_in11 = imem04_in[11:8];
    74: op1_01_in11 = reg_0174;
    47: op1_01_in11 = reg_0157;
    75: op1_01_in11 = reg_0254;
    44: op1_01_in11 = reg_0345;
    56: op1_01_in11 = reg_0721;
    87: op1_01_in11 = reg_1503;
    40: op1_01_in11 = reg_0102;
    37: op1_01_in11 = reg_0001;
    76: op1_01_in11 = reg_0189;
    57: op1_01_in11 = reg_0867;
    70: op1_01_in11 = reg_0758;
    77: op1_01_in11 = reg_0992;
    88: op1_01_in11 = reg_0488;
    78: op1_01_in11 = imem01_in[15:12];
    42: op1_01_in11 = reg_0146;
    79: op1_01_in11 = reg_0799;
    35: op1_01_in11 = imem02_in[3:0];
    62: op1_01_in11 = reg_0335;
    80: op1_01_in11 = reg_0987;
    81: op1_01_in11 = reg_0722;
    89: op1_01_in11 = reg_1299;
    63: op1_01_in11 = reg_0401;
    82: op1_01_in11 = reg_1227;
    98: op1_01_in11 = reg_1227;
    122: op1_01_in11 = reg_1227;
    83: op1_01_in11 = reg_0433;
    128: op1_01_in11 = reg_0433;
    39: op1_01_in11 = reg_0065;
    64: op1_01_in11 = reg_0934;
    84: op1_01_in11 = reg_1321;
    65: op1_01_in11 = reg_0801;
    85: op1_01_in11 = reg_0351;
    95: op1_01_in11 = reg_0351;
    90: op1_01_in11 = reg_1492;
    66: op1_01_in11 = reg_0435;
    91: op1_01_in11 = reg_0444;
    92: op1_01_in11 = reg_0058;
    93: op1_01_in11 = reg_0648;
    94: op1_01_in11 = reg_0330;
    96: op1_01_in11 = reg_0104;
    97: op1_01_in11 = reg_0291;
    99: op1_01_in11 = reg_0299;
    100: op1_01_in11 = reg_0429;
    102: op1_01_in11 = reg_1437;
    104: op1_01_in11 = reg_0881;
    118: op1_01_in11 = reg_0881;
    105: op1_01_in11 = reg_1368;
    106: op1_01_in11 = reg_0142;
    107: op1_01_in11 = reg_0391;
    108: op1_01_in11 = reg_0465;
    109: op1_01_in11 = reg_1180;
    110: op1_01_in11 = reg_0402;
    111: op1_01_in11 = reg_1467;
    112: op1_01_in11 = reg_1451;
    113: op1_01_in11 = reg_0308;
    114: op1_01_in11 = reg_0297;
    115: op1_01_in11 = reg_1432;
    116: op1_01_in11 = reg_0436;
    117: op1_01_in11 = imem01_in[11:8];
    43: op1_01_in11 = reg_0175;
    119: op1_01_in11 = reg_0459;
    120: op1_01_in11 = reg_0957;
    121: op1_01_in11 = reg_0196;
    123: op1_01_in11 = reg_0565;
    125: op1_01_in11 = reg_0201;
    126: op1_01_in11 = reg_0599;
    127: op1_01_in11 = reg_1230;
    129: op1_01_in11 = reg_1202;
    130: op1_01_in11 = reg_0202;
    131: op1_01_in11 = reg_0622;
    default: op1_01_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv11 = 1;
    52: op1_01_inv11 = 1;
    53: op1_01_inv11 = 1;
    61: op1_01_inv11 = 1;
    55: op1_01_inv11 = 1;
    71: op1_01_inv11 = 1;
    86: op1_01_inv11 = 1;
    69: op1_01_inv11 = 1;
    59: op1_01_inv11 = 1;
    50: op1_01_inv11 = 1;
    75: op1_01_inv11 = 1;
    56: op1_01_inv11 = 1;
    40: op1_01_inv11 = 1;
    37: op1_01_inv11 = 1;
    76: op1_01_inv11 = 1;
    57: op1_01_inv11 = 1;
    77: op1_01_inv11 = 1;
    78: op1_01_inv11 = 1;
    42: op1_01_inv11 = 1;
    79: op1_01_inv11 = 1;
    35: op1_01_inv11 = 1;
    62: op1_01_inv11 = 1;
    81: op1_01_inv11 = 1;
    89: op1_01_inv11 = 1;
    63: op1_01_inv11 = 1;
    82: op1_01_inv11 = 1;
    39: op1_01_inv11 = 1;
    64: op1_01_inv11 = 1;
    65: op1_01_inv11 = 1;
    66: op1_01_inv11 = 1;
    91: op1_01_inv11 = 1;
    92: op1_01_inv11 = 1;
    94: op1_01_inv11 = 1;
    96: op1_01_inv11 = 1;
    97: op1_01_inv11 = 1;
    101: op1_01_inv11 = 1;
    102: op1_01_inv11 = 1;
    106: op1_01_inv11 = 1;
    107: op1_01_inv11 = 1;
    109: op1_01_inv11 = 1;
    111: op1_01_inv11 = 1;
    112: op1_01_inv11 = 1;
    115: op1_01_inv11 = 1;
    116: op1_01_inv11 = 1;
    118: op1_01_inv11 = 1;
    43: op1_01_inv11 = 1;
    121: op1_01_inv11 = 1;
    122: op1_01_inv11 = 1;
    123: op1_01_inv11 = 1;
    124: op1_01_inv11 = 1;
    127: op1_01_inv11 = 1;
    128: op1_01_inv11 = 1;
    129: op1_01_inv11 = 1;
    130: op1_01_inv11 = 1;
    default: op1_01_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の12番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in12 = reg_0156;
    52: op1_01_in12 = reg_0876;
    53: op1_01_in12 = reg_0587;
    67: op1_01_in12 = reg_1313;
    61: op1_01_in12 = reg_0352;
    130: op1_01_in12 = reg_0352;
    72: op1_01_in12 = reg_0928;
    58: op1_01_in12 = reg_0114;
    68: op1_01_in12 = reg_0376;
    55: op1_01_in12 = reg_0862;
    73: op1_01_in12 = reg_0120;
    71: op1_01_in12 = reg_0886;
    104: op1_01_in12 = reg_0886;
    48: op1_01_in12 = reg_0326;
    86: op1_01_in12 = reg_0975;
    69: op1_01_in12 = reg_0506;
    59: op1_01_in12 = reg_0722;
    82: op1_01_in12 = reg_0722;
    50: op1_01_in12 = reg_0991;
    60: op1_01_in12 = reg_0878;
    46: op1_01_in12 = reg_0904;
    74: op1_01_in12 = reg_0272;
    47: op1_01_in12 = reg_0140;
    75: op1_01_in12 = reg_0776;
    44: op1_01_in12 = reg_0702;
    56: op1_01_in12 = reg_0369;
    87: op1_01_in12 = imem05_in[11:8];
    40: op1_01_in12 = reg_0361;
    37: op1_01_in12 = reg_0002;
    76: op1_01_in12 = reg_0405;
    57: op1_01_in12 = reg_0298;
    70: op1_01_in12 = reg_0227;
    77: op1_01_in12 = reg_0346;
    88: op1_01_in12 = reg_1215;
    78: op1_01_in12 = reg_0553;
    42: op1_01_in12 = reg_0402;
    79: op1_01_in12 = reg_0449;
    35: op1_01_in12 = reg_0254;
    62: op1_01_in12 = reg_0175;
    80: op1_01_in12 = reg_0961;
    81: op1_01_in12 = reg_0189;
    95: op1_01_in12 = reg_0189;
    125: op1_01_in12 = reg_0189;
    89: op1_01_in12 = reg_1431;
    63: op1_01_in12 = reg_0385;
    83: op1_01_in12 = reg_1455;
    39: op1_01_in12 = reg_0064;
    64: op1_01_in12 = reg_0935;
    84: op1_01_in12 = reg_1100;
    65: op1_01_in12 = reg_0802;
    85: op1_01_in12 = reg_0431;
    90: op1_01_in12 = reg_0069;
    66: op1_01_in12 = reg_0388;
    91: op1_01_in12 = reg_1448;
    92: op1_01_in12 = reg_0005;
    93: op1_01_in12 = reg_0174;
    94: op1_01_in12 = reg_1447;
    96: op1_01_in12 = reg_0882;
    97: op1_01_in12 = reg_0288;
    98: op1_01_in12 = reg_0155;
    99: op1_01_in12 = reg_0457;
    100: op1_01_in12 = reg_0971;
    116: op1_01_in12 = reg_0971;
    101: op1_01_in12 = reg_0927;
    102: op1_01_in12 = reg_0751;
    105: op1_01_in12 = reg_0088;
    106: op1_01_in12 = reg_0627;
    107: op1_01_in12 = reg_0182;
    27: op1_01_in12 = reg_0245;
    108: op1_01_in12 = reg_0285;
    109: op1_01_in12 = reg_0940;
    110: op1_01_in12 = reg_0634;
    111: op1_01_in12 = reg_0584;
    112: op1_01_in12 = reg_0105;
    113: op1_01_in12 = reg_0289;
    114: op1_01_in12 = reg_1203;
    115: op1_01_in12 = reg_0229;
    117: op1_01_in12 = reg_0980;
    118: op1_01_in12 = reg_0887;
    43: op1_01_in12 = reg_0221;
    119: op1_01_in12 = reg_0476;
    120: op1_01_in12 = reg_0104;
    121: op1_01_in12 = reg_0240;
    122: op1_01_in12 = reg_1206;
    123: op1_01_in12 = imem06_in[3:0];
    124: op1_01_in12 = reg_0458;
    126: op1_01_in12 = reg_1041;
    127: op1_01_in12 = reg_1418;
    128: op1_01_in12 = reg_1451;
    129: op1_01_in12 = reg_0754;
    131: op1_01_in12 = reg_0419;
    default: op1_01_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv12 = 1;
    72: op1_01_inv12 = 1;
    58: op1_01_inv12 = 1;
    68: op1_01_inv12 = 1;
    55: op1_01_inv12 = 1;
    73: op1_01_inv12 = 1;
    71: op1_01_inv12 = 1;
    48: op1_01_inv12 = 1;
    59: op1_01_inv12 = 1;
    50: op1_01_inv12 = 1;
    60: op1_01_inv12 = 1;
    46: op1_01_inv12 = 1;
    75: op1_01_inv12 = 1;
    44: op1_01_inv12 = 1;
    87: op1_01_inv12 = 1;
    37: op1_01_inv12 = 1;
    88: op1_01_inv12 = 1;
    42: op1_01_inv12 = 1;
    79: op1_01_inv12 = 1;
    62: op1_01_inv12 = 1;
    89: op1_01_inv12 = 1;
    63: op1_01_inv12 = 1;
    83: op1_01_inv12 = 1;
    39: op1_01_inv12 = 1;
    84: op1_01_inv12 = 1;
    85: op1_01_inv12 = 1;
    66: op1_01_inv12 = 1;
    91: op1_01_inv12 = 1;
    93: op1_01_inv12 = 1;
    98: op1_01_inv12 = 1;
    99: op1_01_inv12 = 1;
    100: op1_01_inv12 = 1;
    101: op1_01_inv12 = 1;
    104: op1_01_inv12 = 1;
    105: op1_01_inv12 = 1;
    106: op1_01_inv12 = 1;
    107: op1_01_inv12 = 1;
    108: op1_01_inv12 = 1;
    109: op1_01_inv12 = 1;
    113: op1_01_inv12 = 1;
    114: op1_01_inv12 = 1;
    116: op1_01_inv12 = 1;
    43: op1_01_inv12 = 1;
    119: op1_01_inv12 = 1;
    121: op1_01_inv12 = 1;
    124: op1_01_inv12 = 1;
    127: op1_01_inv12 = 1;
    128: op1_01_inv12 = 1;
    default: op1_01_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の13番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in13 = reg_0139;
    52: op1_01_in13 = reg_0845;
    53: op1_01_in13 = imem02_in[7:4];
    67: op1_01_in13 = reg_1226;
    61: op1_01_in13 = reg_0005;
    72: op1_01_in13 = reg_0352;
    58: op1_01_in13 = reg_0521;
    40: op1_01_in13 = reg_0521;
    68: op1_01_in13 = reg_0180;
    55: op1_01_in13 = reg_0837;
    73: op1_01_in13 = reg_0192;
    71: op1_01_in13 = reg_0722;
    48: op1_01_in13 = reg_0778;
    75: op1_01_in13 = reg_0778;
    86: op1_01_in13 = reg_0263;
    69: op1_01_in13 = reg_0507;
    59: op1_01_in13 = reg_0201;
    50: op1_01_in13 = reg_0432;
    60: op1_01_in13 = reg_0830;
    46: op1_01_in13 = reg_0368;
    74: op1_01_in13 = reg_1404;
    47: op1_01_in13 = reg_0030;
    44: op1_01_in13 = reg_0174;
    56: op1_01_in13 = reg_0341;
    87: op1_01_in13 = imem05_in[15:12];
    37: op1_01_in13 = reg_0483;
    76: op1_01_in13 = reg_0389;
    57: op1_01_in13 = reg_0299;
    70: op1_01_in13 = imem03_in[7:4];
    77: op1_01_in13 = reg_0131;
    88: op1_01_in13 = reg_0681;
    78: op1_01_in13 = reg_0550;
    42: op1_01_in13 = reg_0401;
    79: op1_01_in13 = reg_0038;
    35: op1_01_in13 = reg_0256;
    62: op1_01_in13 = reg_0695;
    80: op1_01_in13 = reg_0821;
    122: op1_01_in13 = reg_0821;
    81: op1_01_in13 = reg_0409;
    89: op1_01_in13 = reg_1163;
    63: op1_01_in13 = reg_0091;
    82: op1_01_in13 = reg_0387;
    83: op1_01_in13 = reg_0105;
    39: op1_01_in13 = reg_0061;
    64: op1_01_in13 = reg_0126;
    84: op1_01_in13 = reg_0611;
    65: op1_01_in13 = reg_0279;
    85: op1_01_in13 = reg_0075;
    90: op1_01_in13 = reg_0154;
    66: op1_01_in13 = reg_0058;
    91: op1_01_in13 = reg_0557;
    92: op1_01_in13 = reg_0917;
    93: op1_01_in13 = reg_0066;
    94: op1_01_in13 = reg_0177;
    95: op1_01_in13 = reg_0410;
    96: op1_01_in13 = reg_0541;
    97: op1_01_in13 = reg_1282;
    98: op1_01_in13 = reg_0459;
    127: op1_01_in13 = reg_0459;
    99: op1_01_in13 = reg_1350;
    100: op1_01_in13 = reg_1458;
    101: op1_01_in13 = reg_1393;
    102: op1_01_in13 = reg_0860;
    104: op1_01_in13 = reg_0188;
    130: op1_01_in13 = reg_0188;
    105: op1_01_in13 = reg_0034;
    106: op1_01_in13 = reg_1300;
    107: op1_01_in13 = reg_0630;
    27: op1_01_in13 = reg_0156;
    108: op1_01_in13 = reg_0442;
    109: op1_01_in13 = reg_0303;
    110: op1_01_in13 = reg_0895;
    111: op1_01_in13 = reg_0617;
    112: op1_01_in13 = reg_0684;
    116: op1_01_in13 = reg_0684;
    113: op1_01_in13 = reg_0214;
    114: op1_01_in13 = reg_0281;
    115: op1_01_in13 = reg_0155;
    117: op1_01_in13 = reg_0635;
    118: op1_01_in13 = reg_0886;
    43: op1_01_in13 = reg_0445;
    119: op1_01_in13 = reg_0881;
    120: op1_01_in13 = reg_0885;
    121: op1_01_in13 = reg_1348;
    123: op1_01_in13 = reg_0929;
    124: op1_01_in13 = reg_0025;
    125: op1_01_in13 = reg_0203;
    126: op1_01_in13 = reg_0320;
    128: op1_01_in13 = reg_0106;
    129: op1_01_in13 = reg_0215;
    131: op1_01_in13 = reg_0754;
    default: op1_01_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv13 = 1;
    52: op1_01_inv13 = 1;
    67: op1_01_inv13 = 1;
    72: op1_01_inv13 = 1;
    58: op1_01_inv13 = 1;
    68: op1_01_inv13 = 1;
    55: op1_01_inv13 = 1;
    71: op1_01_inv13 = 1;
    86: op1_01_inv13 = 1;
    69: op1_01_inv13 = 1;
    59: op1_01_inv13 = 1;
    60: op1_01_inv13 = 1;
    47: op1_01_inv13 = 1;
    56: op1_01_inv13 = 1;
    87: op1_01_inv13 = 1;
    57: op1_01_inv13 = 1;
    70: op1_01_inv13 = 1;
    77: op1_01_inv13 = 1;
    88: op1_01_inv13 = 1;
    79: op1_01_inv13 = 1;
    62: op1_01_inv13 = 1;
    81: op1_01_inv13 = 1;
    63: op1_01_inv13 = 1;
    83: op1_01_inv13 = 1;
    39: op1_01_inv13 = 1;
    64: op1_01_inv13 = 1;
    90: op1_01_inv13 = 1;
    66: op1_01_inv13 = 1;
    94: op1_01_inv13 = 1;
    97: op1_01_inv13 = 1;
    98: op1_01_inv13 = 1;
    101: op1_01_inv13 = 1;
    102: op1_01_inv13 = 1;
    104: op1_01_inv13 = 1;
    105: op1_01_inv13 = 1;
    106: op1_01_inv13 = 1;
    107: op1_01_inv13 = 1;
    108: op1_01_inv13 = 1;
    109: op1_01_inv13 = 1;
    113: op1_01_inv13 = 1;
    114: op1_01_inv13 = 1;
    115: op1_01_inv13 = 1;
    116: op1_01_inv13 = 1;
    118: op1_01_inv13 = 1;
    119: op1_01_inv13 = 1;
    120: op1_01_inv13 = 1;
    121: op1_01_inv13 = 1;
    122: op1_01_inv13 = 1;
    125: op1_01_inv13 = 1;
    127: op1_01_inv13 = 1;
    129: op1_01_inv13 = 1;
    131: op1_01_inv13 = 1;
    default: op1_01_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の14番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in14 = reg_0123;
    52: op1_01_in14 = reg_0154;
    53: op1_01_in14 = imem02_in[15:12];
    67: op1_01_in14 = reg_1092;
    61: op1_01_in14 = imem01_in[3:0];
    72: op1_01_in14 = reg_0188;
    68: op1_01_in14 = reg_0963;
    55: op1_01_in14 = reg_0117;
    73: op1_01_in14 = reg_0925;
    71: op1_01_in14 = reg_0189;
    48: op1_01_in14 = reg_0127;
    86: op1_01_in14 = imem04_in[15:12];
    69: op1_01_in14 = reg_0525;
    60: op1_01_in14 = reg_0525;
    59: op1_01_in14 = reg_0387;
    81: op1_01_in14 = reg_0387;
    50: op1_01_in14 = reg_0778;
    46: op1_01_in14 = reg_0164;
    105: op1_01_in14 = reg_0164;
    74: op1_01_in14 = imem05_in[7:4];
    47: op1_01_in14 = reg_0665;
    75: op1_01_in14 = reg_1458;
    44: op1_01_in14 = reg_0523;
    56: op1_01_in14 = reg_0596;
    87: op1_01_in14 = reg_0333;
    40: op1_01_in14 = reg_0483;
    76: op1_01_in14 = reg_0060;
    85: op1_01_in14 = reg_0060;
    57: op1_01_in14 = reg_0851;
    70: op1_01_in14 = reg_0704;
    77: op1_01_in14 = reg_1180;
    88: op1_01_in14 = reg_0500;
    78: op1_01_in14 = reg_0746;
    42: op1_01_in14 = reg_0383;
    79: op1_01_in14 = imem06_in[7:4];
    35: op1_01_in14 = reg_0631;
    62: op1_01_in14 = reg_1253;
    80: op1_01_in14 = reg_0886;
    89: op1_01_in14 = reg_0392;
    63: op1_01_in14 = reg_0047;
    82: op1_01_in14 = reg_0071;
    83: op1_01_in14 = reg_0629;
    39: op1_01_in14 = imem05_in[11:8];
    64: op1_01_in14 = reg_0900;
    84: op1_01_in14 = reg_0335;
    65: op1_01_in14 = reg_0756;
    90: op1_01_in14 = reg_0789;
    66: op1_01_in14 = reg_0723;
    92: op1_01_in14 = reg_0723;
    91: op1_01_in14 = reg_0600;
    93: op1_01_in14 = reg_0701;
    94: op1_01_in14 = reg_0180;
    95: op1_01_in14 = reg_0405;
    96: op1_01_in14 = reg_0348;
    97: op1_01_in14 = reg_1280;
    98: op1_01_in14 = reg_1405;
    122: op1_01_in14 = reg_1405;
    99: op1_01_in14 = reg_0923;
    100: op1_01_in14 = reg_0128;
    101: op1_01_in14 = reg_0881;
    102: op1_01_in14 = reg_1504;
    104: op1_01_in14 = reg_0409;
    130: op1_01_in14 = reg_0409;
    106: op1_01_in14 = reg_0329;
    107: op1_01_in14 = reg_0564;
    27: op1_01_in14 = reg_0287;
    108: op1_01_in14 = reg_0621;
    109: op1_01_in14 = reg_0090;
    110: op1_01_in14 = reg_0447;
    111: op1_01_in14 = reg_0528;
    112: op1_01_in14 = reg_0829;
    113: op1_01_in14 = reg_0015;
    114: op1_01_in14 = reg_1214;
    115: op1_01_in14 = reg_1406;
    116: op1_01_in14 = reg_0560;
    117: op1_01_in14 = reg_1290;
    118: op1_01_in14 = reg_0431;
    43: op1_01_in14 = reg_0567;
    119: op1_01_in14 = reg_0352;
    120: op1_01_in14 = reg_0448;
    121: op1_01_in14 = reg_0589;
    123: op1_01_in14 = reg_1437;
    124: op1_01_in14 = reg_0673;
    125: op1_01_in14 = reg_0072;
    126: op1_01_in14 = reg_0698;
    127: op1_01_in14 = reg_0476;
    128: op1_01_in14 = reg_0105;
    129: op1_01_in14 = reg_0018;
    131: op1_01_in14 = reg_0396;
    default: op1_01_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv14 = 1;
    53: op1_01_inv14 = 1;
    67: op1_01_inv14 = 1;
    55: op1_01_inv14 = 1;
    59: op1_01_inv14 = 1;
    60: op1_01_inv14 = 1;
    46: op1_01_inv14 = 1;
    74: op1_01_inv14 = 1;
    47: op1_01_inv14 = 1;
    44: op1_01_inv14 = 1;
    56: op1_01_inv14 = 1;
    87: op1_01_inv14 = 1;
    77: op1_01_inv14 = 1;
    88: op1_01_inv14 = 1;
    42: op1_01_inv14 = 1;
    35: op1_01_inv14 = 1;
    81: op1_01_inv14 = 1;
    82: op1_01_inv14 = 1;
    83: op1_01_inv14 = 1;
    64: op1_01_inv14 = 1;
    84: op1_01_inv14 = 1;
    65: op1_01_inv14 = 1;
    90: op1_01_inv14 = 1;
    66: op1_01_inv14 = 1;
    91: op1_01_inv14 = 1;
    94: op1_01_inv14 = 1;
    104: op1_01_inv14 = 1;
    105: op1_01_inv14 = 1;
    107: op1_01_inv14 = 1;
    109: op1_01_inv14 = 1;
    114: op1_01_inv14 = 1;
    117: op1_01_inv14 = 1;
    119: op1_01_inv14 = 1;
    120: op1_01_inv14 = 1;
    121: op1_01_inv14 = 1;
    123: op1_01_inv14 = 1;
    124: op1_01_inv14 = 1;
    127: op1_01_inv14 = 1;
    130: op1_01_inv14 = 1;
    131: op1_01_inv14 = 1;
    default: op1_01_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の15番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in15 = reg_0100;
    52: op1_01_in15 = reg_0325;
    53: op1_01_in15 = reg_0475;
    67: op1_01_in15 = reg_0104;
    61: op1_01_in15 = reg_1255;
    72: op1_01_in15 = reg_0440;
    68: op1_01_in15 = reg_0314;
    55: op1_01_in15 = reg_0208;
    73: op1_01_in15 = reg_1334;
    71: op1_01_in15 = reg_0405;
    48: op1_01_in15 = reg_0055;
    86: op1_01_in15 = reg_1258;
    69: op1_01_in15 = reg_0573;
    59: op1_01_in15 = reg_0353;
    98: op1_01_in15 = reg_0353;
    50: op1_01_in15 = reg_0970;
    60: op1_01_in15 = reg_0734;
    46: op1_01_in15 = reg_0065;
    74: op1_01_in15 = imem05_in[15:12];
    47: op1_01_in15 = reg_0661;
    75: op1_01_in15 = reg_0125;
    44: op1_01_in15 = reg_0650;
    56: op1_01_in15 = reg_0199;
    87: op1_01_in15 = reg_0347;
    40: op1_01_in15 = reg_0484;
    76: op1_01_in15 = reg_0059;
    57: op1_01_in15 = reg_0775;
    70: op1_01_in15 = reg_0177;
    77: op1_01_in15 = reg_0794;
    88: op1_01_in15 = reg_1147;
    78: op1_01_in15 = reg_0609;
    42: op1_01_in15 = reg_0365;
    79: op1_01_in15 = imem06_in[11:8];
    35: op1_01_in15 = reg_0561;
    62: op1_01_in15 = reg_0550;
    80: op1_01_in15 = reg_0722;
    81: op1_01_in15 = reg_0072;
    82: op1_01_in15 = reg_0072;
    89: op1_01_in15 = reg_0491;
    63: op1_01_in15 = reg_0078;
    83: op1_01_in15 = reg_0876;
    39: op1_01_in15 = reg_0749;
    64: op1_01_in15 = reg_0705;
    84: op1_01_in15 = reg_0161;
    65: op1_01_in15 = reg_0525;
    85: op1_01_in15 = reg_0917;
    125: op1_01_in15 = reg_0917;
    90: op1_01_in15 = reg_0375;
    66: op1_01_in15 = reg_0785;
    91: op1_01_in15 = reg_0144;
    92: op1_01_in15 = imem01_in[7:4];
    93: op1_01_in15 = reg_1181;
    94: op1_01_in15 = reg_0556;
    95: op1_01_in15 = reg_0387;
    96: op1_01_in15 = imem04_in[11:8];
    97: op1_01_in15 = reg_0411;
    99: op1_01_in15 = reg_0489;
    100: op1_01_in15 = reg_0106;
    101: op1_01_in15 = reg_0431;
    102: op1_01_in15 = reg_0374;
    104: op1_01_in15 = reg_0410;
    105: op1_01_in15 = reg_0731;
    106: op1_01_in15 = reg_0350;
    107: op1_01_in15 = reg_1070;
    27: op1_01_in15 = reg_0441;
    108: op1_01_in15 = reg_0593;
    109: op1_01_in15 = reg_0888;
    110: op1_01_in15 = imem02_in[3:0];
    111: op1_01_in15 = reg_0529;
    112: op1_01_in15 = reg_0800;
    113: op1_01_in15 = reg_0022;
    129: op1_01_in15 = reg_0022;
    114: op1_01_in15 = reg_1082;
    115: op1_01_in15 = reg_0928;
    116: op1_01_in15 = reg_0294;
    117: op1_01_in15 = reg_0553;
    118: op1_01_in15 = reg_0203;
    43: op1_01_in15 = reg_0566;
    119: op1_01_in15 = reg_0389;
    120: op1_01_in15 = reg_0378;
    121: op1_01_in15 = reg_0799;
    122: op1_01_in15 = reg_0476;
    123: op1_01_in15 = reg_0751;
    124: op1_01_in15 = reg_1280;
    126: op1_01_in15 = reg_0262;
    127: op1_01_in15 = reg_0927;
    128: op1_01_in15 = reg_0253;
    130: op1_01_in15 = reg_0073;
    131: op1_01_in15 = reg_0023;
    default: op1_01_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    67: op1_01_inv15 = 1;
    73: op1_01_inv15 = 1;
    69: op1_01_inv15 = 1;
    50: op1_01_inv15 = 1;
    60: op1_01_inv15 = 1;
    75: op1_01_inv15 = 1;
    44: op1_01_inv15 = 1;
    56: op1_01_inv15 = 1;
    87: op1_01_inv15 = 1;
    40: op1_01_inv15 = 1;
    76: op1_01_inv15 = 1;
    42: op1_01_inv15 = 1;
    79: op1_01_inv15 = 1;
    35: op1_01_inv15 = 1;
    80: op1_01_inv15 = 1;
    81: op1_01_inv15 = 1;
    89: op1_01_inv15 = 1;
    63: op1_01_inv15 = 1;
    39: op1_01_inv15 = 1;
    84: op1_01_inv15 = 1;
    65: op1_01_inv15 = 1;
    85: op1_01_inv15 = 1;
    90: op1_01_inv15 = 1;
    91: op1_01_inv15 = 1;
    92: op1_01_inv15 = 1;
    93: op1_01_inv15 = 1;
    95: op1_01_inv15 = 1;
    97: op1_01_inv15 = 1;
    98: op1_01_inv15 = 1;
    99: op1_01_inv15 = 1;
    100: op1_01_inv15 = 1;
    104: op1_01_inv15 = 1;
    106: op1_01_inv15 = 1;
    109: op1_01_inv15 = 1;
    110: op1_01_inv15 = 1;
    113: op1_01_inv15 = 1;
    116: op1_01_inv15 = 1;
    117: op1_01_inv15 = 1;
    118: op1_01_inv15 = 1;
    43: op1_01_inv15 = 1;
    122: op1_01_inv15 = 1;
    123: op1_01_inv15 = 1;
    124: op1_01_inv15 = 1;
    125: op1_01_inv15 = 1;
    130: op1_01_inv15 = 1;
    default: op1_01_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の16番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in16 = reg_0085;
    52: op1_01_in16 = imem03_in[3:0];
    53: op1_01_in16 = reg_0990;
    67: op1_01_in16 = reg_0885;
    61: op1_01_in16 = reg_0575;
    72: op1_01_in16 = reg_0134;
    101: op1_01_in16 = reg_0134;
    68: op1_01_in16 = reg_0190;
    55: op1_01_in16 = reg_0064;
    73: op1_01_in16 = imem06_in[11:8];
    71: op1_01_in16 = reg_0611;
    66: op1_01_in16 = reg_0611;
    48: op1_01_in16 = reg_0897;
    86: op1_01_in16 = reg_0796;
    114: op1_01_in16 = reg_0796;
    69: op1_01_in16 = reg_0443;
    59: op1_01_in16 = reg_0351;
    50: op1_01_in16 = reg_0128;
    60: op1_01_in16 = reg_0630;
    46: op1_01_in16 = reg_0150;
    74: op1_01_in16 = reg_0318;
    47: op1_01_in16 = reg_0287;
    75: op1_01_in16 = reg_0878;
    44: op1_01_in16 = reg_0602;
    56: op1_01_in16 = reg_0319;
    87: op1_01_in16 = reg_0184;
    40: op1_01_in16 = reg_0124;
    76: op1_01_in16 = reg_0058;
    81: op1_01_in16 = reg_0058;
    57: op1_01_in16 = reg_0774;
    70: op1_01_in16 = reg_1425;
    77: op1_01_in16 = reg_1514;
    88: op1_01_in16 = reg_0320;
    78: op1_01_in16 = reg_0819;
    42: op1_01_in16 = reg_0363;
    79: op1_01_in16 = reg_0261;
    35: op1_01_in16 = reg_0531;
    105: op1_01_in16 = reg_0531;
    62: op1_01_in16 = reg_0238;
    80: op1_01_in16 = reg_0435;
    89: op1_01_in16 = reg_1181;
    63: op1_01_in16 = reg_0079;
    82: op1_01_in16 = reg_1321;
    83: op1_01_in16 = reg_0153;
    39: op1_01_in16 = reg_0750;
    64: op1_01_in16 = reg_0876;
    84: op1_01_in16 = reg_1290;
    65: op1_01_in16 = reg_0677;
    85: op1_01_in16 = reg_1256;
    90: op1_01_in16 = reg_0964;
    91: op1_01_in16 = reg_0377;
    92: op1_01_in16 = reg_1254;
    93: op1_01_in16 = reg_1404;
    94: op1_01_in16 = reg_1184;
    95: op1_01_in16 = reg_0389;
    96: op1_01_in16 = reg_0467;
    97: op1_01_in16 = imem04_in[15:12];
    98: op1_01_in16 = reg_0722;
    99: op1_01_in16 = reg_0223;
    100: op1_01_in16 = reg_0382;
    102: op1_01_in16 = reg_0622;
    104: op1_01_in16 = reg_0071;
    106: op1_01_in16 = reg_1149;
    107: op1_01_in16 = reg_0938;
    27: op1_01_in16 = reg_0442;
    108: op1_01_in16 = reg_0592;
    109: op1_01_in16 = reg_0130;
    110: op1_01_in16 = reg_0530;
    111: op1_01_in16 = reg_0979;
    112: op1_01_in16 = reg_0069;
    113: op1_01_in16 = imem07_in[15:12];
    115: op1_01_in16 = reg_0428;
    116: op1_01_in16 = reg_0007;
    117: op1_01_in16 = reg_0746;
    118: op1_01_in16 = reg_0060;
    43: op1_01_in16 = reg_0182;
    119: op1_01_in16 = reg_1324;
    120: op1_01_in16 = reg_1280;
    121: op1_01_in16 = reg_0864;
    122: op1_01_in16 = reg_0927;
    123: op1_01_in16 = reg_0863;
    124: op1_01_in16 = imem04_in[7:4];
    125: op1_01_in16 = imem01_in[7:4];
    126: op1_01_in16 = reg_0836;
    127: op1_01_in16 = reg_0887;
    128: op1_01_in16 = reg_0068;
    129: op1_01_in16 = imem07_in[11:8];
    130: op1_01_in16 = imem01_in[11:8];
    131: op1_01_in16 = reg_0215;
    default: op1_01_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    15: op1_01_inv16 = 1;
    67: op1_01_inv16 = 1;
    55: op1_01_inv16 = 1;
    73: op1_01_inv16 = 1;
    71: op1_01_inv16 = 1;
    48: op1_01_inv16 = 1;
    69: op1_01_inv16 = 1;
    46: op1_01_inv16 = 1;
    75: op1_01_inv16 = 1;
    44: op1_01_inv16 = 1;
    56: op1_01_inv16 = 1;
    57: op1_01_inv16 = 1;
    42: op1_01_inv16 = 1;
    35: op1_01_inv16 = 1;
    62: op1_01_inv16 = 1;
    80: op1_01_inv16 = 1;
    83: op1_01_inv16 = 1;
    64: op1_01_inv16 = 1;
    65: op1_01_inv16 = 1;
    66: op1_01_inv16 = 1;
    92: op1_01_inv16 = 1;
    94: op1_01_inv16 = 1;
    98: op1_01_inv16 = 1;
    107: op1_01_inv16 = 1;
    27: op1_01_inv16 = 1;
    108: op1_01_inv16 = 1;
    111: op1_01_inv16 = 1;
    114: op1_01_inv16 = 1;
    116: op1_01_inv16 = 1;
    117: op1_01_inv16 = 1;
    119: op1_01_inv16 = 1;
    121: op1_01_inv16 = 1;
    122: op1_01_inv16 = 1;
    123: op1_01_inv16 = 1;
    124: op1_01_inv16 = 1;
    125: op1_01_inv16 = 1;
    127: op1_01_inv16 = 1;
    128: op1_01_inv16 = 1;
    130: op1_01_inv16 = 1;
    131: op1_01_inv16 = 1;
    default: op1_01_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の17番目の入力
  always @ ( * ) begin
    case ( state )
    15: op1_01_in17 = reg_0050;
    52: op1_01_in17 = reg_1092;
    53: op1_01_in17 = reg_0991;
    67: op1_01_in17 = reg_0504;
    61: op1_01_in17 = reg_0550;
    72: op1_01_in17 = reg_0073;
    68: op1_01_in17 = reg_0597;
    55: op1_01_in17 = reg_0032;
    73: op1_01_in17 = reg_0115;
    71: op1_01_in17 = reg_1290;
    48: op1_01_in17 = reg_0898;
    86: op1_01_in17 = reg_0094;
    69: op1_01_in17 = reg_1258;
    59: op1_01_in17 = reg_0071;
    50: op1_01_in17 = reg_0125;
    60: op1_01_in17 = reg_1145;
    46: op1_01_in17 = reg_0211;
    74: op1_01_in17 = reg_0601;
    47: op1_01_in17 = reg_0408;
    75: op1_01_in17 = reg_0380;
    44: op1_01_in17 = reg_0603;
    56: op1_01_in17 = reg_0368;
    87: op1_01_in17 = reg_0346;
    76: op1_01_in17 = reg_0372;
    57: op1_01_in17 = reg_0029;
    70: op1_01_in17 = reg_1325;
    77: op1_01_in17 = reg_0872;
    88: op1_01_in17 = reg_0342;
    78: op1_01_in17 = reg_0430;
    42: op1_01_in17 = reg_0047;
    79: op1_01_in17 = reg_0192;
    35: op1_01_in17 = reg_0475;
    62: op1_01_in17 = reg_0241;
    80: op1_01_in17 = reg_0405;
    127: op1_01_in17 = reg_0405;
    81: op1_01_in17 = reg_1321;
    89: op1_01_in17 = reg_1180;
    63: op1_01_in17 = reg_0282;
    82: op1_01_in17 = reg_0005;
    83: op1_01_in17 = reg_0306;
    39: op1_01_in17 = reg_0700;
    64: op1_01_in17 = reg_0878;
    84: op1_01_in17 = reg_0448;
    65: op1_01_in17 = reg_0675;
    85: op1_01_in17 = reg_0547;
    90: op1_01_in17 = reg_0142;
    91: op1_01_in17 = reg_0142;
    66: op1_01_in17 = reg_1256;
    92: op1_01_in17 = reg_0166;
    93: op1_01_in17 = reg_0986;
    94: op1_01_in17 = reg_0964;
    95: op1_01_in17 = reg_0203;
    96: op1_01_in17 = reg_0493;
    97: op1_01_in17 = reg_0467;
    98: op1_01_in17 = reg_0435;
    115: op1_01_in17 = reg_0435;
    99: op1_01_in17 = reg_0139;
    100: op1_01_in17 = reg_0628;
    101: op1_01_in17 = reg_0388;
    102: op1_01_in17 = reg_0526;
    104: op1_01_in17 = reg_0075;
    105: op1_01_in17 = reg_1215;
    106: op1_01_in17 = reg_0458;
    107: op1_01_in17 = reg_0792;
    27: op1_01_in17 = reg_0413;
    108: op1_01_in17 = reg_0084;
    109: op1_01_in17 = imem06_in[7:4];
    121: op1_01_in17 = imem06_in[7:4];
    110: op1_01_in17 = reg_0607;
    111: op1_01_in17 = reg_0323;
    112: op1_01_in17 = reg_0279;
    113: op1_01_in17 = reg_0478;
    114: op1_01_in17 = reg_1041;
    116: op1_01_in17 = reg_1078;
    117: op1_01_in17 = reg_0610;
    118: op1_01_in17 = reg_0057;
    43: op1_01_in17 = reg_0541;
    119: op1_01_in17 = imem01_in[11:8];
    120: op1_01_in17 = imem04_in[11:8];
    122: op1_01_in17 = reg_0886;
    123: op1_01_in17 = reg_0717;
    124: op1_01_in17 = reg_0534;
    125: op1_01_in17 = reg_0966;
    126: op1_01_in17 = reg_1312;
    128: op1_01_in17 = reg_0227;
    129: op1_01_in17 = imem07_in[15:12];
    130: op1_01_in17 = reg_0163;
    131: op1_01_in17 = reg_0213;
    default: op1_01_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_01_inv17 = 1;
    68: op1_01_inv17 = 1;
    71: op1_01_inv17 = 1;
    48: op1_01_inv17 = 1;
    86: op1_01_inv17 = 1;
    59: op1_01_inv17 = 1;
    60: op1_01_inv17 = 1;
    46: op1_01_inv17 = 1;
    75: op1_01_inv17 = 1;
    76: op1_01_inv17 = 1;
    70: op1_01_inv17 = 1;
    77: op1_01_inv17 = 1;
    88: op1_01_inv17 = 1;
    78: op1_01_inv17 = 1;
    42: op1_01_inv17 = 1;
    79: op1_01_inv17 = 1;
    89: op1_01_inv17 = 1;
    63: op1_01_inv17 = 1;
    83: op1_01_inv17 = 1;
    90: op1_01_inv17 = 1;
    66: op1_01_inv17 = 1;
    92: op1_01_inv17 = 1;
    94: op1_01_inv17 = 1;
    98: op1_01_inv17 = 1;
    101: op1_01_inv17 = 1;
    104: op1_01_inv17 = 1;
    106: op1_01_inv17 = 1;
    107: op1_01_inv17 = 1;
    27: op1_01_inv17 = 1;
    110: op1_01_inv17 = 1;
    112: op1_01_inv17 = 1;
    114: op1_01_inv17 = 1;
    116: op1_01_inv17 = 1;
    43: op1_01_inv17 = 1;
    119: op1_01_inv17 = 1;
    120: op1_01_inv17 = 1;
    124: op1_01_inv17 = 1;
    126: op1_01_inv17 = 1;
    128: op1_01_inv17 = 1;
    129: op1_01_inv17 = 1;
    130: op1_01_inv17 = 1;
    131: op1_01_inv17 = 1;
    default: op1_01_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の18番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in18 = reg_1063;
    53: op1_01_in18 = reg_0436;
    67: op1_01_in18 = reg_0480;
    61: op1_01_in18 = reg_0548;
    72: op1_01_in18 = reg_0059;
    68: op1_01_in18 = reg_0246;
    55: op1_01_in18 = reg_0033;
    73: op1_01_in18 = reg_0619;
    71: op1_01_in18 = reg_0448;
    48: op1_01_in18 = reg_0705;
    86: op1_01_in18 = reg_1147;
    69: op1_01_in18 = reg_1198;
    59: op1_01_in18 = reg_0073;
    95: op1_01_in18 = reg_0073;
    50: op1_01_in18 = reg_0111;
    60: op1_01_in18 = reg_0025;
    46: op1_01_in18 = reg_0745;
    74: op1_01_in18 = reg_0861;
    47: op1_01_in18 = reg_0413;
    75: op1_01_in18 = reg_0381;
    44: op1_01_in18 = reg_0564;
    56: op1_01_in18 = reg_0019;
    87: op1_01_in18 = reg_0066;
    76: op1_01_in18 = reg_1291;
    57: op1_01_in18 = reg_0030;
    70: op1_01_in18 = reg_0145;
    77: op1_01_in18 = reg_1373;
    88: op1_01_in18 = reg_0319;
    78: op1_01_in18 = reg_1457;
    42: op1_01_in18 = imem01_in[3:0];
    79: op1_01_in18 = reg_1509;
    35: op1_01_in18 = reg_0474;
    62: op1_01_in18 = reg_0439;
    80: op1_01_in18 = reg_0203;
    81: op1_01_in18 = reg_0089;
    89: op1_01_in18 = reg_1404;
    63: op1_01_in18 = reg_0042;
    82: op1_01_in18 = reg_0917;
    118: op1_01_in18 = reg_0917;
    127: op1_01_in18 = reg_0917;
    83: op1_01_in18 = reg_0379;
    39: op1_01_in18 = reg_0173;
    64: op1_01_in18 = reg_0327;
    84: op1_01_in18 = reg_0277;
    65: op1_01_in18 = reg_0707;
    85: op1_01_in18 = reg_0609;
    90: op1_01_in18 = reg_0070;
    66: op1_01_in18 = reg_0547;
    91: op1_01_in18 = reg_1517;
    92: op1_01_in18 = reg_0787;
    93: op1_01_in18 = reg_0303;
    94: op1_01_in18 = reg_0142;
    96: op1_01_in18 = reg_1214;
    97: op1_01_in18 = reg_1372;
    98: op1_01_in18 = reg_0388;
    99: op1_01_in18 = reg_0777;
    100: op1_01_in18 = reg_0631;
    101: op1_01_in18 = reg_0057;
    102: op1_01_in18 = reg_0522;
    104: op1_01_in18 = reg_1322;
    105: op1_01_in18 = reg_0796;
    106: op1_01_in18 = reg_1282;
    107: op1_01_in18 = reg_1163;
    27: op1_01_in18 = reg_0228;
    108: op1_01_in18 = reg_0521;
    109: op1_01_in18 = reg_1105;
    110: op1_01_in18 = reg_0276;
    111: op1_01_in18 = reg_1204;
    112: op1_01_in18 = reg_0563;
    113: op1_01_in18 = reg_1060;
    114: op1_01_in18 = reg_1419;
    115: op1_01_in18 = reg_0410;
    116: op1_01_in18 = reg_1091;
    117: op1_01_in18 = reg_0241;
    43: op1_01_in18 = reg_0490;
    119: op1_01_in18 = reg_0577;
    120: op1_01_in18 = reg_0534;
    121: op1_01_in18 = reg_0270;
    122: op1_01_in18 = reg_0202;
    123: op1_01_in18 = reg_0637;
    124: op1_01_in18 = reg_1369;
    125: op1_01_in18 = reg_0047;
    126: op1_01_in18 = reg_0256;
    128: op1_01_in18 = reg_0006;
    129: op1_01_in18 = reg_0394;
    130: op1_01_in18 = reg_0549;
    131: op1_01_in18 = imem07_in[7:4];
    default: op1_01_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    68: op1_01_inv18 = 1;
    55: op1_01_inv18 = 1;
    71: op1_01_inv18 = 1;
    86: op1_01_inv18 = 1;
    69: op1_01_inv18 = 1;
    59: op1_01_inv18 = 1;
    50: op1_01_inv18 = 1;
    47: op1_01_inv18 = 1;
    75: op1_01_inv18 = 1;
    56: op1_01_inv18 = 1;
    87: op1_01_inv18 = 1;
    77: op1_01_inv18 = 1;
    78: op1_01_inv18 = 1;
    79: op1_01_inv18 = 1;
    62: op1_01_inv18 = 1;
    80: op1_01_inv18 = 1;
    89: op1_01_inv18 = 1;
    63: op1_01_inv18 = 1;
    82: op1_01_inv18 = 1;
    64: op1_01_inv18 = 1;
    84: op1_01_inv18 = 1;
    90: op1_01_inv18 = 1;
    91: op1_01_inv18 = 1;
    92: op1_01_inv18 = 1;
    94: op1_01_inv18 = 1;
    99: op1_01_inv18 = 1;
    100: op1_01_inv18 = 1;
    104: op1_01_inv18 = 1;
    105: op1_01_inv18 = 1;
    106: op1_01_inv18 = 1;
    107: op1_01_inv18 = 1;
    110: op1_01_inv18 = 1;
    112: op1_01_inv18 = 1;
    115: op1_01_inv18 = 1;
    116: op1_01_inv18 = 1;
    43: op1_01_inv18 = 1;
    119: op1_01_inv18 = 1;
    121: op1_01_inv18 = 1;
    122: op1_01_inv18 = 1;
    124: op1_01_inv18 = 1;
    127: op1_01_inv18 = 1;
    default: op1_01_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の19番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in19 = reg_0697;
    53: op1_01_in19 = reg_0054;
    67: op1_01_in19 = imem04_in[7:4];
    61: op1_01_in19 = reg_0259;
    72: op1_01_in19 = reg_0122;
    68: op1_01_in19 = reg_1301;
    55: op1_01_in19 = reg_0793;
    73: op1_01_in19 = reg_0570;
    71: op1_01_in19 = reg_1255;
    48: op1_01_in19 = reg_0846;
    86: op1_01_in19 = reg_0406;
    69: op1_01_in19 = reg_1083;
    59: op1_01_in19 = reg_0723;
    82: op1_01_in19 = reg_0723;
    50: op1_01_in19 = reg_0379;
    60: op1_01_in19 = reg_0952;
    46: op1_01_in19 = reg_0733;
    74: op1_01_in19 = reg_0040;
    47: op1_01_in19 = reg_0618;
    75: op1_01_in19 = reg_0695;
    44: op1_01_in19 = reg_0182;
    56: op1_01_in19 = reg_0032;
    87: op1_01_in19 = reg_0491;
    43: op1_01_in19 = reg_0491;
    76: op1_01_in19 = imem01_in[7:4];
    42: op1_01_in19 = imem01_in[7:4];
    80: op1_01_in19 = imem01_in[7:4];
    57: op1_01_in19 = reg_0665;
    70: op1_01_in19 = reg_0142;
    77: op1_01_in19 = reg_0243;
    88: op1_01_in19 = reg_0835;
    78: op1_01_in19 = reg_0726;
    79: op1_01_in19 = reg_1323;
    35: op1_01_in19 = reg_0456;
    62: op1_01_in19 = reg_0438;
    81: op1_01_in19 = reg_0446;
    89: op1_01_in19 = reg_0940;
    63: op1_01_in19 = reg_0044;
    83: op1_01_in19 = reg_0531;
    39: op1_01_in19 = reg_0176;
    64: op1_01_in19 = reg_0069;
    84: op1_01_in19 = reg_0258;
    125: op1_01_in19 = reg_0258;
    65: op1_01_in19 = reg_0709;
    85: op1_01_in19 = reg_1474;
    90: op1_01_in19 = reg_0627;
    66: op1_01_in19 = reg_0609;
    91: op1_01_in19 = reg_0048;
    92: op1_01_in19 = reg_0242;
    93: op1_01_in19 = reg_0090;
    94: op1_01_in19 = reg_0070;
    95: op1_01_in19 = reg_1322;
    96: op1_01_in19 = reg_1082;
    97: op1_01_in19 = reg_1198;
    98: op1_01_in19 = reg_0058;
    99: op1_01_in19 = reg_0779;
    100: op1_01_in19 = reg_1091;
    101: op1_01_in19 = reg_1324;
    102: op1_01_in19 = reg_0296;
    104: op1_01_in19 = reg_0089;
    105: op1_01_in19 = reg_0421;
    106: op1_01_in19 = reg_0348;
    107: op1_01_in19 = reg_0197;
    27: op1_01_in19 = reg_0229;
    109: op1_01_in19 = reg_1064;
    110: op1_01_in19 = reg_1074;
    111: op1_01_in19 = reg_1202;
    112: op1_01_in19 = imem03_in[3:0];
    116: op1_01_in19 = imem03_in[3:0];
    113: op1_01_in19 = reg_0703;
    114: op1_01_in19 = reg_0369;
    115: op1_01_in19 = reg_0134;
    117: op1_01_in19 = reg_0434;
    118: op1_01_in19 = imem01_in[3:0];
    127: op1_01_in19 = imem01_in[3:0];
    119: op1_01_in19 = reg_0982;
    120: op1_01_in19 = reg_1368;
    121: op1_01_in19 = reg_0333;
    122: op1_01_in19 = reg_0351;
    123: op1_01_in19 = reg_0979;
    124: op1_01_in19 = reg_0328;
    126: op1_01_in19 = reg_1151;
    128: op1_01_in19 = imem03_in[15:12];
    129: op1_01_in19 = reg_0922;
    130: op1_01_in19 = reg_0222;
    131: op1_01_in19 = reg_1010;
    default: op1_01_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    68: op1_01_inv19 = 1;
    73: op1_01_inv19 = 1;
    48: op1_01_inv19 = 1;
    69: op1_01_inv19 = 1;
    59: op1_01_inv19 = 1;
    50: op1_01_inv19 = 1;
    74: op1_01_inv19 = 1;
    56: op1_01_inv19 = 1;
    87: op1_01_inv19 = 1;
    57: op1_01_inv19 = 1;
    70: op1_01_inv19 = 1;
    42: op1_01_inv19 = 1;
    62: op1_01_inv19 = 1;
    81: op1_01_inv19 = 1;
    89: op1_01_inv19 = 1;
    63: op1_01_inv19 = 1;
    39: op1_01_inv19 = 1;
    84: op1_01_inv19 = 1;
    65: op1_01_inv19 = 1;
    90: op1_01_inv19 = 1;
    93: op1_01_inv19 = 1;
    95: op1_01_inv19 = 1;
    96: op1_01_inv19 = 1;
    97: op1_01_inv19 = 1;
    100: op1_01_inv19 = 1;
    107: op1_01_inv19 = 1;
    109: op1_01_inv19 = 1;
    112: op1_01_inv19 = 1;
    113: op1_01_inv19 = 1;
    114: op1_01_inv19 = 1;
    116: op1_01_inv19 = 1;
    118: op1_01_inv19 = 1;
    120: op1_01_inv19 = 1;
    123: op1_01_inv19 = 1;
    124: op1_01_inv19 = 1;
    125: op1_01_inv19 = 1;
    default: op1_01_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の20番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in20 = reg_0232;
    53: op1_01_in20 = reg_0776;
    67: op1_01_in20 = imem04_in[11:8];
    61: op1_01_in20 = reg_0161;
    72: op1_01_in20 = reg_1100;
    68: op1_01_in20 = reg_0107;
    55: op1_01_in20 = reg_0391;
    73: op1_01_in20 = reg_1228;
    71: op1_01_in20 = reg_0549;
    48: op1_01_in20 = reg_0830;
    86: op1_01_in20 = reg_0407;
    69: op1_01_in20 = reg_0412;
    105: op1_01_in20 = reg_0412;
    59: op1_01_in20 = reg_1031;
    50: op1_01_in20 = reg_0056;
    60: op1_01_in20 = imem03_in[7:4];
    46: op1_01_in20 = reg_0833;
    74: op1_01_in20 = reg_0014;
    47: op1_01_in20 = reg_0361;
    75: op1_01_in20 = reg_0069;
    44: op1_01_in20 = reg_0332;
    56: op1_01_in20 = reg_0631;
    87: op1_01_in20 = reg_0167;
    76: op1_01_in20 = reg_0553;
    57: op1_01_in20 = reg_0623;
    70: op1_01_in20 = reg_0964;
    77: op1_01_in20 = reg_1346;
    88: op1_01_in20 = reg_0063;
    78: op1_01_in20 = reg_0147;
    42: op1_01_in20 = reg_0080;
    79: op1_01_in20 = reg_1504;
    35: op1_01_in20 = reg_0452;
    62: op1_01_in20 = reg_0726;
    80: op1_01_in20 = imem01_in[15:12];
    81: op1_01_in20 = reg_0788;
    89: op1_01_in20 = reg_0939;
    63: op1_01_in20 = reg_0011;
    82: op1_01_in20 = imem01_in[7:4];
    83: op1_01_in20 = reg_0563;
    39: op1_01_in20 = reg_0523;
    64: op1_01_in20 = reg_0279;
    84: op1_01_in20 = reg_0550;
    65: op1_01_in20 = reg_1139;
    85: op1_01_in20 = reg_0966;
    90: op1_01_in20 = reg_0220;
    66: op1_01_in20 = reg_0715;
    91: op1_01_in20 = reg_1226;
    92: op1_01_in20 = reg_0820;
    93: op1_01_in20 = reg_0872;
    94: op1_01_in20 = reg_1518;
    95: op1_01_in20 = reg_0089;
    96: op1_01_in20 = reg_1147;
    97: op1_01_in20 = reg_0681;
    98: op1_01_in20 = imem01_in[3:0];
    99: op1_01_in20 = reg_0465;
    100: op1_01_in20 = reg_0009;
    101: op1_01_in20 = reg_0267;
    102: op1_01_in20 = reg_0244;
    104: op1_01_in20 = reg_0917;
    106: op1_01_in20 = reg_0427;
    107: op1_01_in20 = reg_0130;
    27: op1_01_in20 = reg_0219;
    109: op1_01_in20 = reg_0795;
    110: op1_01_in20 = reg_0494;
    111: op1_01_in20 = reg_0215;
    112: op1_01_in20 = imem03_in[11:8];
    113: op1_01_in20 = reg_0851;
    114: op1_01_in20 = reg_1151;
    115: op1_01_in20 = reg_0388;
    116: op1_01_in20 = reg_0377;
    117: op1_01_in20 = reg_0149;
    118: op1_01_in20 = reg_0985;
    43: op1_01_in20 = reg_0418;
    119: op1_01_in20 = reg_1152;
    120: op1_01_in20 = reg_0088;
    121: op1_01_in20 = reg_1334;
    122: op1_01_in20 = reg_0189;
    123: op1_01_in20 = reg_0195;
    124: op1_01_in20 = reg_0462;
    125: op1_01_in20 = reg_0899;
    126: op1_01_in20 = reg_0096;
    127: op1_01_in20 = reg_0746;
    128: op1_01_in20 = reg_0732;
    129: op1_01_in20 = reg_0231;
    130: op1_01_in20 = reg_0260;
    131: op1_01_in20 = reg_0922;
    default: op1_01_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_01_inv20 = 1;
    67: op1_01_inv20 = 1;
    73: op1_01_inv20 = 1;
    71: op1_01_inv20 = 1;
    69: op1_01_inv20 = 1;
    50: op1_01_inv20 = 1;
    60: op1_01_inv20 = 1;
    74: op1_01_inv20 = 1;
    47: op1_01_inv20 = 1;
    76: op1_01_inv20 = 1;
    70: op1_01_inv20 = 1;
    78: op1_01_inv20 = 1;
    42: op1_01_inv20 = 1;
    79: op1_01_inv20 = 1;
    35: op1_01_inv20 = 1;
    62: op1_01_inv20 = 1;
    80: op1_01_inv20 = 1;
    81: op1_01_inv20 = 1;
    89: op1_01_inv20 = 1;
    63: op1_01_inv20 = 1;
    64: op1_01_inv20 = 1;
    65: op1_01_inv20 = 1;
    92: op1_01_inv20 = 1;
    97: op1_01_inv20 = 1;
    98: op1_01_inv20 = 1;
    100: op1_01_inv20 = 1;
    101: op1_01_inv20 = 1;
    105: op1_01_inv20 = 1;
    106: op1_01_inv20 = 1;
    27: op1_01_inv20 = 1;
    114: op1_01_inv20 = 1;
    116: op1_01_inv20 = 1;
    118: op1_01_inv20 = 1;
    43: op1_01_inv20 = 1;
    119: op1_01_inv20 = 1;
    121: op1_01_inv20 = 1;
    122: op1_01_inv20 = 1;
    125: op1_01_inv20 = 1;
    126: op1_01_inv20 = 1;
    127: op1_01_inv20 = 1;
    129: op1_01_inv20 = 1;
    130: op1_01_inv20 = 1;
    default: op1_01_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の21番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in21 = reg_1003;
    53: op1_01_in21 = reg_0972;
    67: op1_01_in21 = imem04_in[15:12];
    61: op1_01_in21 = reg_0966;
    72: op1_01_in21 = reg_0553;
    68: op1_01_in21 = imem03_in[7:4];
    55: op1_01_in21 = reg_0579;
    73: op1_01_in21 = reg_0171;
    71: op1_01_in21 = reg_0550;
    48: op1_01_in21 = reg_0802;
    86: op1_01_in21 = reg_0451;
    69: op1_01_in21 = reg_0599;
    59: op1_01_in21 = reg_1034;
    50: op1_01_in21 = reg_0708;
    60: op1_01_in21 = reg_1208;
    46: op1_01_in21 = reg_0832;
    74: op1_01_in21 = reg_1105;
    47: op1_01_in21 = reg_0228;
    75: op1_01_in21 = reg_0325;
    44: op1_01_in21 = reg_0540;
    56: op1_01_in21 = reg_0391;
    87: op1_01_in21 = reg_0697;
    76: op1_01_in21 = reg_0547;
    57: op1_01_in21 = reg_0103;
    70: op1_01_in21 = reg_0597;
    77: op1_01_in21 = reg_0799;
    88: op1_01_in21 = reg_0633;
    78: op1_01_in21 = reg_0402;
    42: op1_01_in21 = reg_0078;
    79: op1_01_in21 = reg_0717;
    35: op1_01_in21 = reg_0138;
    62: op1_01_in21 = reg_0383;
    80: op1_01_in21 = reg_1254;
    81: op1_01_in21 = reg_0277;
    89: op1_01_in21 = reg_0794;
    63: op1_01_in21 = reg_0010;
    82: op1_01_in21 = reg_0448;
    83: op1_01_in21 = reg_1132;
    39: op1_01_in21 = reg_0648;
    64: op1_01_in21 = reg_0312;
    84: op1_01_in21 = reg_0222;
    65: op1_01_in21 = reg_0143;
    85: op1_01_in21 = reg_0968;
    90: op1_01_in21 = reg_1231;
    66: op1_01_in21 = reg_0147;
    91: op1_01_in21 = reg_0880;
    92: op1_01_in21 = reg_1473;
    93: op1_01_in21 = reg_0318;
    94: op1_01_in21 = reg_0954;
    95: op1_01_in21 = reg_0027;
    96: op1_01_in21 = reg_0407;
    97: op1_01_in21 = reg_0500;
    98: op1_01_in21 = reg_0985;
    99: op1_01_in21 = reg_0404;
    100: op1_01_in21 = reg_0227;
    101: op1_01_in21 = imem01_in[15:12];
    102: op1_01_in21 = reg_0165;
    104: op1_01_in21 = imem01_in[7:4];
    105: op1_01_in21 = reg_0406;
    106: op1_01_in21 = imem04_in[7:4];
    107: op1_01_in21 = reg_0039;
    27: op1_01_in21 = reg_0052;
    109: op1_01_in21 = reg_0192;
    110: op1_01_in21 = reg_0970;
    111: op1_01_in21 = reg_0015;
    112: op1_01_in21 = reg_1063;
    113: op1_01_in21 = reg_0775;
    114: op1_01_in21 = reg_0096;
    115: op1_01_in21 = reg_0075;
    116: op1_01_in21 = reg_1145;
    117: op1_01_in21 = reg_0148;
    118: op1_01_in21 = reg_0874;
    43: op1_01_in21 = reg_0302;
    119: op1_01_in21 = reg_0241;
    120: op1_01_in21 = reg_0531;
    121: op1_01_in21 = reg_0782;
    122: op1_01_in21 = reg_0389;
    123: op1_01_in21 = reg_0152;
    124: op1_01_in21 = reg_0421;
    125: op1_01_in21 = reg_0901;
    126: op1_01_in21 = reg_0536;
    127: op1_01_in21 = reg_0747;
    128: op1_01_in21 = reg_0154;
    129: op1_01_in21 = reg_1056;
    130: op1_01_in21 = reg_0609;
    131: op1_01_in21 = reg_0050;
    default: op1_01_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    67: op1_01_inv21 = 1;
    72: op1_01_inv21 = 1;
    68: op1_01_inv21 = 1;
    71: op1_01_inv21 = 1;
    48: op1_01_inv21 = 1;
    59: op1_01_inv21 = 1;
    50: op1_01_inv21 = 1;
    74: op1_01_inv21 = 1;
    47: op1_01_inv21 = 1;
    75: op1_01_inv21 = 1;
    77: op1_01_inv21 = 1;
    88: op1_01_inv21 = 1;
    42: op1_01_inv21 = 1;
    79: op1_01_inv21 = 1;
    62: op1_01_inv21 = 1;
    80: op1_01_inv21 = 1;
    81: op1_01_inv21 = 1;
    89: op1_01_inv21 = 1;
    63: op1_01_inv21 = 1;
    83: op1_01_inv21 = 1;
    39: op1_01_inv21 = 1;
    64: op1_01_inv21 = 1;
    84: op1_01_inv21 = 1;
    65: op1_01_inv21 = 1;
    85: op1_01_inv21 = 1;
    90: op1_01_inv21 = 1;
    66: op1_01_inv21 = 1;
    91: op1_01_inv21 = 1;
    93: op1_01_inv21 = 1;
    96: op1_01_inv21 = 1;
    97: op1_01_inv21 = 1;
    98: op1_01_inv21 = 1;
    105: op1_01_inv21 = 1;
    106: op1_01_inv21 = 1;
    107: op1_01_inv21 = 1;
    116: op1_01_inv21 = 1;
    117: op1_01_inv21 = 1;
    118: op1_01_inv21 = 1;
    119: op1_01_inv21 = 1;
    120: op1_01_inv21 = 1;
    125: op1_01_inv21 = 1;
    126: op1_01_inv21 = 1;
    127: op1_01_inv21 = 1;
    default: op1_01_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の22番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in22 = reg_0964;
    53: op1_01_in22 = reg_0105;
    67: op1_01_in22 = reg_1383;
    61: op1_01_in22 = reg_0147;
    72: op1_01_in22 = reg_0093;
    81: op1_01_in22 = reg_0093;
    68: op1_01_in22 = reg_0330;
    55: op1_01_in22 = reg_0750;
    73: op1_01_in22 = reg_0152;
    71: op1_01_in22 = reg_0239;
    48: op1_01_in22 = reg_0800;
    86: op1_01_in22 = reg_0342;
    69: op1_01_in22 = reg_0796;
    97: op1_01_in22 = reg_0796;
    59: op1_01_in22 = reg_0576;
    50: op1_01_in22 = reg_0006;
    60: op1_01_in22 = reg_0113;
    46: op1_01_in22 = reg_0701;
    74: op1_01_in22 = reg_0399;
    47: op1_01_in22 = reg_0002;
    99: op1_01_in22 = reg_0002;
    75: op1_01_in22 = reg_0279;
    44: op1_01_in22 = reg_0490;
    56: op1_01_in22 = reg_0748;
    87: op1_01_in22 = reg_1402;
    76: op1_01_in22 = reg_0747;
    57: op1_01_in22 = reg_0051;
    70: op1_01_in22 = reg_1208;
    77: op1_01_in22 = reg_0864;
    88: op1_01_in22 = imem05_in[11:8];
    78: op1_01_in22 = reg_0384;
    42: op1_01_in22 = reg_0282;
    101: op1_01_in22 = reg_0282;
    79: op1_01_in22 = reg_0617;
    35: op1_01_in22 = reg_0112;
    62: op1_01_in22 = reg_0091;
    80: op1_01_in22 = reg_0166;
    89: op1_01_in22 = reg_0450;
    63: op1_01_in22 = reg_0744;
    82: op1_01_in22 = reg_0754;
    83: op1_01_in22 = reg_1494;
    39: op1_01_in22 = reg_0649;
    64: op1_01_in22 = reg_0227;
    84: op1_01_in22 = reg_0743;
    65: op1_01_in22 = reg_0891;
    85: op1_01_in22 = reg_0819;
    90: op1_01_in22 = reg_0107;
    66: op1_01_in22 = reg_0149;
    91: op1_01_in22 = reg_0218;
    92: op1_01_in22 = reg_0438;
    93: op1_01_in22 = reg_1485;
    94: op1_01_in22 = reg_1093;
    95: op1_01_in22 = reg_0267;
    96: op1_01_in22 = reg_0454;
    98: op1_01_in22 = reg_1254;
    104: op1_01_in22 = reg_1254;
    100: op1_01_in22 = imem03_in[7:4];
    102: op1_01_in22 = reg_1204;
    105: op1_01_in22 = reg_1041;
    106: op1_01_in22 = reg_1340;
    107: op1_01_in22 = imem06_in[15:12];
    109: op1_01_in22 = reg_0870;
    110: op1_01_in22 = reg_1458;
    111: op1_01_in22 = reg_1170;
    112: op1_01_in22 = reg_0198;
    113: op1_01_in22 = reg_0031;
    114: op1_01_in22 = reg_0035;
    115: op1_01_in22 = reg_0058;
    116: op1_01_in22 = reg_0185;
    117: op1_01_in22 = reg_0868;
    118: op1_01_in22 = reg_0930;
    43: op1_01_in22 = reg_0300;
    119: op1_01_in22 = reg_0820;
    120: op1_01_in22 = reg_0297;
    121: op1_01_in22 = reg_0860;
    122: op1_01_in22 = reg_0060;
    123: op1_01_in22 = reg_0212;
    124: op1_01_in22 = reg_0451;
    125: op1_01_in22 = reg_0595;
    126: op1_01_in22 = reg_0065;
    127: op1_01_in22 = reg_0241;
    128: op1_01_in22 = reg_0573;
    129: op1_01_in22 = reg_0224;
    130: op1_01_in22 = reg_1475;
    131: op1_01_in22 = reg_0231;
    default: op1_01_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_01_inv22 = 1;
    67: op1_01_inv22 = 1;
    61: op1_01_inv22 = 1;
    68: op1_01_inv22 = 1;
    55: op1_01_inv22 = 1;
    71: op1_01_inv22 = 1;
    48: op1_01_inv22 = 1;
    46: op1_01_inv22 = 1;
    74: op1_01_inv22 = 1;
    75: op1_01_inv22 = 1;
    44: op1_01_inv22 = 1;
    70: op1_01_inv22 = 1;
    77: op1_01_inv22 = 1;
    88: op1_01_inv22 = 1;
    42: op1_01_inv22 = 1;
    35: op1_01_inv22 = 1;
    62: op1_01_inv22 = 1;
    80: op1_01_inv22 = 1;
    81: op1_01_inv22 = 1;
    63: op1_01_inv22 = 1;
    82: op1_01_inv22 = 1;
    39: op1_01_inv22 = 1;
    84: op1_01_inv22 = 1;
    90: op1_01_inv22 = 1;
    91: op1_01_inv22 = 1;
    97: op1_01_inv22 = 1;
    98: op1_01_inv22 = 1;
    99: op1_01_inv22 = 1;
    102: op1_01_inv22 = 1;
    104: op1_01_inv22 = 1;
    105: op1_01_inv22 = 1;
    107: op1_01_inv22 = 1;
    112: op1_01_inv22 = 1;
    117: op1_01_inv22 = 1;
    43: op1_01_inv22 = 1;
    119: op1_01_inv22 = 1;
    121: op1_01_inv22 = 1;
    122: op1_01_inv22 = 1;
    123: op1_01_inv22 = 1;
    124: op1_01_inv22 = 1;
    125: op1_01_inv22 = 1;
    128: op1_01_inv22 = 1;
    129: op1_01_inv22 = 1;
    131: op1_01_inv22 = 1;
    default: op1_01_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の23番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in23 = reg_0957;
    53: op1_01_in23 = reg_0876;
    67: op1_01_in23 = reg_0263;
    61: op1_01_in23 = reg_0899;
    72: op1_01_in23 = imem01_in[11:8];
    68: op1_01_in23 = reg_0790;
    55: op1_01_in23 = reg_0733;
    73: op1_01_in23 = reg_0213;
    71: op1_01_in23 = reg_0743;
    48: op1_01_in23 = reg_0758;
    86: op1_01_in23 = reg_0340;
    69: op1_01_in23 = reg_0797;
    59: op1_01_in23 = reg_0610;
    50: op1_01_in23 = reg_0068;
    60: op1_01_in23 = reg_0505;
    46: op1_01_in23 = reg_0697;
    74: op1_01_in23 = reg_0795;
    47: op1_01_in23 = reg_0084;
    75: op1_01_in23 = imem02_in[3:0];
    44: op1_01_in23 = reg_0888;
    56: op1_01_in23 = reg_0831;
    87: op1_01_in23 = reg_0477;
    76: op1_01_in23 = reg_0242;
    57: op1_01_in23 = reg_0002;
    70: op1_01_in23 = reg_0884;
    77: op1_01_in23 = reg_0449;
    88: op1_01_in23 = reg_0578;
    78: op1_01_in23 = reg_0386;
    42: op1_01_in23 = reg_0043;
    79: op1_01_in23 = reg_0571;
    35: op1_01_in23 = reg_0106;
    62: op1_01_in23 = reg_0724;
    80: op1_01_in23 = reg_0550;
    81: op1_01_in23 = reg_0463;
    89: op1_01_in23 = reg_0937;
    63: op1_01_in23 = reg_1029;
    82: op1_01_in23 = reg_0963;
    83: op1_01_in23 = reg_1000;
    39: op1_01_in23 = reg_0603;
    64: op1_01_in23 = reg_0235;
    84: op1_01_in23 = reg_0260;
    65: op1_01_in23 = reg_0559;
    85: op1_01_in23 = reg_0403;
    90: op1_01_in23 = reg_0882;
    66: op1_01_in23 = reg_0148;
    92: op1_01_in23 = reg_0148;
    91: op1_01_in23 = reg_0291;
    93: op1_01_in23 = reg_0576;
    94: op1_01_in23 = reg_0178;
    95: op1_01_in23 = imem01_in[3:0];
    115: op1_01_in23 = imem01_in[3:0];
    96: op1_01_in23 = reg_1004;
    97: op1_01_in23 = reg_1147;
    98: op1_01_in23 = reg_0785;
    99: op1_01_in23 = reg_0085;
    100: op1_01_in23 = reg_0840;
    101: op1_01_in23 = reg_1253;
    127: op1_01_in23 = reg_1253;
    102: op1_01_in23 = reg_0583;
    104: op1_01_in23 = reg_1290;
    105: op1_01_in23 = reg_1040;
    106: op1_01_in23 = reg_1372;
    107: op1_01_in23 = reg_0826;
    109: op1_01_in23 = reg_0859;
    110: op1_01_in23 = reg_1450;
    111: op1_01_in23 = imem07_in[3:0];
    112: op1_01_in23 = reg_0191;
    113: op1_01_in23 = reg_0663;
    114: op1_01_in23 = reg_0470;
    116: op1_01_in23 = reg_0177;
    117: op1_01_in23 = reg_0727;
    125: op1_01_in23 = reg_0727;
    118: op1_01_in23 = reg_0553;
    43: op1_01_in23 = reg_0090;
    119: op1_01_in23 = reg_0715;
    120: op1_01_in23 = reg_0488;
    121: op1_01_in23 = reg_0863;
    122: op1_01_in23 = reg_0058;
    123: op1_01_in23 = reg_0214;
    124: op1_01_in23 = reg_0368;
    126: op1_01_in23 = reg_0019;
    128: op1_01_in23 = reg_0706;
    129: op1_01_in23 = reg_0623;
    130: op1_01_in23 = reg_0469;
    131: op1_01_in23 = reg_0100;
    default: op1_01_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_01_inv23 = 1;
    53: op1_01_inv23 = 1;
    67: op1_01_inv23 = 1;
    72: op1_01_inv23 = 1;
    71: op1_01_inv23 = 1;
    86: op1_01_inv23 = 1;
    69: op1_01_inv23 = 1;
    59: op1_01_inv23 = 1;
    50: op1_01_inv23 = 1;
    60: op1_01_inv23 = 1;
    74: op1_01_inv23 = 1;
    44: op1_01_inv23 = 1;
    87: op1_01_inv23 = 1;
    76: op1_01_inv23 = 1;
    70: op1_01_inv23 = 1;
    78: op1_01_inv23 = 1;
    35: op1_01_inv23 = 1;
    80: op1_01_inv23 = 1;
    81: op1_01_inv23 = 1;
    63: op1_01_inv23 = 1;
    82: op1_01_inv23 = 1;
    83: op1_01_inv23 = 1;
    64: op1_01_inv23 = 1;
    90: op1_01_inv23 = 1;
    91: op1_01_inv23 = 1;
    92: op1_01_inv23 = 1;
    93: op1_01_inv23 = 1;
    95: op1_01_inv23 = 1;
    96: op1_01_inv23 = 1;
    97: op1_01_inv23 = 1;
    102: op1_01_inv23 = 1;
    105: op1_01_inv23 = 1;
    106: op1_01_inv23 = 1;
    107: op1_01_inv23 = 1;
    112: op1_01_inv23 = 1;
    113: op1_01_inv23 = 1;
    115: op1_01_inv23 = 1;
    116: op1_01_inv23 = 1;
    117: op1_01_inv23 = 1;
    119: op1_01_inv23 = 1;
    120: op1_01_inv23 = 1;
    121: op1_01_inv23 = 1;
    123: op1_01_inv23 = 1;
    124: op1_01_inv23 = 1;
    125: op1_01_inv23 = 1;
    128: op1_01_inv23 = 1;
    130: op1_01_inv23 = 1;
    default: op1_01_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の24番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in24 = reg_0246;
    53: op1_01_in24 = reg_0009;
    67: op1_01_in24 = reg_1367;
    61: op1_01_in24 = reg_0871;
    72: op1_01_in24 = reg_1475;
    68: op1_01_in24 = reg_0488;
    55: op1_01_in24 = reg_0828;
    73: op1_01_in24 = reg_0017;
    71: op1_01_in24 = reg_0572;
    48: op1_01_in24 = reg_0757;
    86: op1_01_in24 = reg_0338;
    69: op1_01_in24 = reg_1419;
    59: op1_01_in24 = reg_0609;
    50: op1_01_in24 = reg_0069;
    60: op1_01_in24 = reg_0481;
    70: op1_01_in24 = reg_0481;
    46: op1_01_in24 = reg_0445;
    74: op1_01_in24 = imem06_in[15:12];
    75: op1_01_in24 = reg_0312;
    44: op1_01_in24 = reg_0302;
    56: op1_01_in24 = reg_0832;
    87: op1_01_in24 = reg_0275;
    76: op1_01_in24 = reg_0238;
    57: op1_01_in24 = reg_0053;
    77: op1_01_in24 = reg_0861;
    88: op1_01_in24 = reg_1430;
    78: op1_01_in24 = reg_0365;
    42: op1_01_in24 = reg_0042;
    79: op1_01_in24 = reg_0296;
    35: op1_01_in24 = reg_0380;
    62: op1_01_in24 = reg_0078;
    80: op1_01_in24 = reg_0830;
    84: op1_01_in24 = reg_0830;
    81: op1_01_in24 = reg_0163;
    89: op1_01_in24 = reg_0090;
    63: op1_01_in24 = reg_0605;
    82: op1_01_in24 = reg_1512;
    83: op1_01_in24 = reg_0328;
    39: op1_01_in24 = reg_0316;
    64: op1_01_in24 = reg_1064;
    65: op1_01_in24 = reg_0954;
    85: op1_01_in24 = reg_0092;
    90: op1_01_in24 = reg_0426;
    66: op1_01_in24 = reg_0403;
    91: op1_01_in24 = reg_0790;
    92: op1_01_in24 = reg_0401;
    93: op1_01_in24 = reg_0274;
    94: op1_01_in24 = reg_0108;
    95: op1_01_in24 = reg_0553;
    98: op1_01_in24 = reg_0553;
    96: op1_01_in24 = reg_0369;
    97: op1_01_in24 = reg_0421;
    99: op1_01_in24 = reg_0520;
    100: op1_01_in24 = reg_0185;
    101: op1_01_in24 = reg_0874;
    102: op1_01_in24 = reg_1202;
    104: op1_01_in24 = reg_0930;
    105: op1_01_in24 = reg_0199;
    106: op1_01_in24 = reg_0694;
    107: op1_01_in24 = reg_1058;
    109: op1_01_in24 = reg_0265;
    110: op1_01_in24 = reg_0496;
    111: op1_01_in24 = reg_1415;
    112: op1_01_in24 = reg_0789;
    113: op1_01_in24 = reg_0442;
    114: op1_01_in24 = imem05_in[7:4];
    115: op1_01_in24 = imem01_in[11:8];
    116: op1_01_in24 = reg_0557;
    117: op1_01_in24 = reg_0335;
    118: op1_01_in24 = reg_0550;
    43: op1_01_in24 = reg_0873;
    119: op1_01_in24 = reg_0434;
    120: op1_01_in24 = reg_1233;
    121: op1_01_in24 = reg_1508;
    122: op1_01_in24 = reg_1321;
    123: op1_01_in24 = reg_0022;
    124: op1_01_in24 = reg_0932;
    125: op1_01_in24 = reg_0634;
    126: op1_01_in24 = reg_0210;
    127: op1_01_in24 = reg_0091;
    128: op1_01_in24 = reg_0597;
    129: op1_01_in24 = reg_0621;
    130: op1_01_in24 = reg_1452;
    131: op1_01_in24 = reg_0703;
    default: op1_01_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_01_inv24 = 1;
    53: op1_01_inv24 = 1;
    61: op1_01_inv24 = 1;
    68: op1_01_inv24 = 1;
    71: op1_01_inv24 = 1;
    86: op1_01_inv24 = 1;
    50: op1_01_inv24 = 1;
    60: op1_01_inv24 = 1;
    46: op1_01_inv24 = 1;
    74: op1_01_inv24 = 1;
    75: op1_01_inv24 = 1;
    44: op1_01_inv24 = 1;
    87: op1_01_inv24 = 1;
    76: op1_01_inv24 = 1;
    70: op1_01_inv24 = 1;
    78: op1_01_inv24 = 1;
    79: op1_01_inv24 = 1;
    81: op1_01_inv24 = 1;
    82: op1_01_inv24 = 1;
    39: op1_01_inv24 = 1;
    64: op1_01_inv24 = 1;
    85: op1_01_inv24 = 1;
    90: op1_01_inv24 = 1;
    91: op1_01_inv24 = 1;
    92: op1_01_inv24 = 1;
    93: op1_01_inv24 = 1;
    94: op1_01_inv24 = 1;
    99: op1_01_inv24 = 1;
    100: op1_01_inv24 = 1;
    101: op1_01_inv24 = 1;
    105: op1_01_inv24 = 1;
    107: op1_01_inv24 = 1;
    110: op1_01_inv24 = 1;
    111: op1_01_inv24 = 1;
    113: op1_01_inv24 = 1;
    115: op1_01_inv24 = 1;
    116: op1_01_inv24 = 1;
    117: op1_01_inv24 = 1;
    118: op1_01_inv24 = 1;
    121: op1_01_inv24 = 1;
    122: op1_01_inv24 = 1;
    125: op1_01_inv24 = 1;
    126: op1_01_inv24 = 1;
    127: op1_01_inv24 = 1;
    128: op1_01_inv24 = 1;
    129: op1_01_inv24 = 1;
    130: op1_01_inv24 = 1;
    131: op1_01_inv24 = 1;
    default: op1_01_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の25番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in25 = reg_0448;
    53: op1_01_in25 = reg_0830;
    67: op1_01_in25 = reg_0252;
    61: op1_01_in25 = imem02_in[7:4];
    72: op1_01_in25 = reg_1474;
    68: op1_01_in25 = reg_1368;
    55: op1_01_in25 = reg_0831;
    73: op1_01_in25 = reg_1439;
    71: op1_01_in25 = reg_0434;
    48: op1_01_in25 = reg_0677;
    86: op1_01_in25 = reg_1151;
    69: op1_01_in25 = reg_0698;
    59: op1_01_in25 = reg_0715;
    50: op1_01_in25 = reg_0802;
    60: op1_01_in25 = reg_0479;
    46: op1_01_in25 = reg_0066;
    74: op1_01_in25 = reg_1065;
    75: op1_01_in25 = reg_0191;
    44: op1_01_in25 = reg_0301;
    56: op1_01_in25 = reg_1169;
    87: op1_01_in25 = reg_0575;
    76: op1_01_in25 = reg_0798;
    57: op1_01_in25 = reg_0086;
    70: op1_01_in25 = reg_0348;
    77: op1_01_in25 = reg_0317;
    88: op1_01_in25 = reg_0347;
    78: op1_01_in25 = reg_0363;
    42: op1_01_in25 = reg_0044;
    79: op1_01_in25 = reg_0289;
    35: op1_01_in25 = reg_0343;
    62: op1_01_in25 = reg_0290;
    80: op1_01_in25 = reg_0147;
    81: op1_01_in25 = reg_0550;
    89: op1_01_in25 = reg_1485;
    63: op1_01_in25 = reg_0455;
    82: op1_01_in25 = reg_1513;
    83: op1_01_in25 = reg_0709;
    39: op1_01_in25 = reg_0450;
    64: op1_01_in25 = reg_0963;
    84: op1_01_in25 = reg_0430;
    65: op1_01_in25 = reg_0329;
    85: op1_01_in25 = reg_0727;
    90: op1_01_in25 = reg_0032;
    66: op1_01_in25 = reg_0401;
    91: op1_01_in25 = reg_0427;
    92: op1_01_in25 = reg_0386;
    93: op1_01_in25 = reg_0861;
    94: op1_01_in25 = reg_0884;
    95: op1_01_in25 = reg_0463;
    98: op1_01_in25 = reg_0463;
    96: op1_01_in25 = reg_0862;
    97: op1_01_in25 = reg_0414;
    100: op1_01_in25 = reg_0444;
    101: op1_01_in25 = reg_0576;
    102: op1_01_in25 = reg_0396;
    104: op1_01_in25 = reg_0047;
    105: op1_01_in25 = reg_0454;
    106: op1_01_in25 = reg_0281;
    107: op1_01_in25 = reg_0269;
    109: op1_01_in25 = reg_0116;
    110: op1_01_in25 = reg_1140;
    111: op1_01_in25 = reg_0894;
    112: op1_01_in25 = reg_0375;
    113: op1_01_in25 = reg_0739;
    114: op1_01_in25 = reg_0251;
    115: op1_01_in25 = reg_1032;
    116: op1_01_in25 = reg_0312;
    117: op1_01_in25 = reg_0080;
    118: op1_01_in25 = reg_0260;
    43: op1_01_in25 = reg_0196;
    119: op1_01_in25 = reg_0726;
    120: op1_01_in25 = reg_0421;
    121: op1_01_in25 = reg_0115;
    122: op1_01_in25 = reg_1322;
    123: op1_01_in25 = imem07_in[7:4];
    124: op1_01_in25 = reg_1502;
    125: op1_01_in25 = reg_0041;
    126: op1_01_in25 = reg_0470;
    127: op1_01_in25 = reg_0162;
    128: op1_01_in25 = reg_1063;
    129: op1_01_in25 = reg_0321;
    130: op1_01_in25 = reg_1034;
    131: op1_01_in25 = reg_0223;
    default: op1_01_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_01_inv25 = 1;
    72: op1_01_inv25 = 1;
    55: op1_01_inv25 = 1;
    71: op1_01_inv25 = 1;
    48: op1_01_inv25 = 1;
    86: op1_01_inv25 = 1;
    50: op1_01_inv25 = 1;
    60: op1_01_inv25 = 1;
    74: op1_01_inv25 = 1;
    75: op1_01_inv25 = 1;
    56: op1_01_inv25 = 1;
    76: op1_01_inv25 = 1;
    57: op1_01_inv25 = 1;
    70: op1_01_inv25 = 1;
    88: op1_01_inv25 = 1;
    78: op1_01_inv25 = 1;
    42: op1_01_inv25 = 1;
    79: op1_01_inv25 = 1;
    89: op1_01_inv25 = 1;
    39: op1_01_inv25 = 1;
    64: op1_01_inv25 = 1;
    85: op1_01_inv25 = 1;
    92: op1_01_inv25 = 1;
    93: op1_01_inv25 = 1;
    95: op1_01_inv25 = 1;
    97: op1_01_inv25 = 1;
    98: op1_01_inv25 = 1;
    101: op1_01_inv25 = 1;
    104: op1_01_inv25 = 1;
    116: op1_01_inv25 = 1;
    118: op1_01_inv25 = 1;
    43: op1_01_inv25 = 1;
    120: op1_01_inv25 = 1;
    127: op1_01_inv25 = 1;
    129: op1_01_inv25 = 1;
    130: op1_01_inv25 = 1;
    default: op1_01_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の26番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in26 = reg_0882;
    53: op1_01_in26 = reg_0829;
    67: op1_01_in26 = reg_0396;
    61: op1_01_in26 = reg_0533;
    72: op1_01_in26 = reg_1452;
    68: op1_01_in26 = reg_1367;
    55: op1_01_in26 = reg_0346;
    73: op1_01_in26 = reg_0391;
    71: op1_01_in26 = reg_0148;
    48: op1_01_in26 = reg_0675;
    86: op1_01_in26 = reg_0536;
    69: op1_01_in26 = reg_0340;
    59: op1_01_in26 = reg_0572;
    50: op1_01_in26 = reg_0311;
    60: op1_01_in26 = reg_0427;
    46: op1_01_in26 = reg_0317;
    74: op1_01_in26 = reg_0718;
    75: op1_01_in26 = reg_0999;
    44: op1_01_in26 = reg_0197;
    39: op1_01_in26 = reg_0197;
    56: op1_01_in26 = reg_0445;
    87: op1_01_in26 = reg_1348;
    76: op1_01_in26 = reg_1475;
    57: op1_01_in26 = reg_0519;
    70: op1_01_in26 = reg_0898;
    77: op1_01_in26 = reg_1064;
    88: op1_01_in26 = reg_0272;
    78: op1_01_in26 = reg_0257;
    42: op1_01_in26 = reg_0041;
    79: op1_01_in26 = reg_0119;
    35: op1_01_in26 = reg_0322;
    62: op1_01_in26 = reg_0169;
    80: op1_01_in26 = reg_0149;
    84: op1_01_in26 = reg_0149;
    81: op1_01_in26 = reg_0966;
    89: op1_01_in26 = reg_1484;
    63: op1_01_in26 = reg_0589;
    82: op1_01_in26 = reg_0047;
    66: op1_01_in26 = reg_0047;
    83: op1_01_in26 = reg_0261;
    64: op1_01_in26 = reg_0962;
    65: op1_01_in26 = reg_1301;
    85: op1_01_in26 = reg_0874;
    90: op1_01_in26 = reg_0088;
    91: op1_01_in26 = imem04_in[11:8];
    92: op1_01_in26 = reg_0362;
    93: op1_01_in26 = reg_0014;
    94: op1_01_in26 = reg_0288;
    95: op1_01_in26 = reg_0549;
    96: op1_01_in26 = reg_0836;
    97: op1_01_in26 = reg_0320;
    98: op1_01_in26 = reg_0550;
    100: op1_01_in26 = reg_1449;
    101: op1_01_in26 = reg_0547;
    102: op1_01_in26 = reg_0067;
    104: op1_01_in26 = reg_0093;
    105: op1_01_in26 = reg_0451;
    106: op1_01_in26 = reg_0407;
    107: op1_01_in26 = reg_1420;
    109: op1_01_in26 = reg_0714;
    121: op1_01_in26 = reg_0714;
    110: op1_01_in26 = reg_0684;
    111: op1_01_in26 = reg_0299;
    112: op1_01_in26 = reg_0965;
    113: op1_01_in26 = reg_0620;
    114: op1_01_in26 = reg_0697;
    115: op1_01_in26 = reg_0985;
    116: op1_01_in26 = reg_0191;
    117: op1_01_in26 = reg_0078;
    118: op1_01_in26 = reg_1473;
    43: op1_01_in26 = reg_0273;
    119: op1_01_in26 = reg_0290;
    120: op1_01_in26 = reg_1041;
    122: op1_01_in26 = reg_0122;
    123: op1_01_in26 = reg_0394;
    124: op1_01_in26 = reg_0021;
    125: op1_01_in26 = reg_0895;
    126: op1_01_in26 = imem05_in[7:4];
    127: op1_01_in26 = reg_0044;
    128: op1_01_in26 = reg_1184;
    129: op1_01_in26 = reg_0052;
    130: op1_01_in26 = reg_0363;
    131: op1_01_in26 = reg_0465;
    default: op1_01_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    61: op1_01_inv26 = 1;
    48: op1_01_inv26 = 1;
    86: op1_01_inv26 = 1;
    69: op1_01_inv26 = 1;
    59: op1_01_inv26 = 1;
    50: op1_01_inv26 = 1;
    60: op1_01_inv26 = 1;
    74: op1_01_inv26 = 1;
    75: op1_01_inv26 = 1;
    44: op1_01_inv26 = 1;
    87: op1_01_inv26 = 1;
    76: op1_01_inv26 = 1;
    70: op1_01_inv26 = 1;
    77: op1_01_inv26 = 1;
    78: op1_01_inv26 = 1;
    62: op1_01_inv26 = 1;
    89: op1_01_inv26 = 1;
    39: op1_01_inv26 = 1;
    84: op1_01_inv26 = 1;
    85: op1_01_inv26 = 1;
    66: op1_01_inv26 = 1;
    92: op1_01_inv26 = 1;
    95: op1_01_inv26 = 1;
    97: op1_01_inv26 = 1;
    98: op1_01_inv26 = 1;
    104: op1_01_inv26 = 1;
    106: op1_01_inv26 = 1;
    107: op1_01_inv26 = 1;
    109: op1_01_inv26 = 1;
    115: op1_01_inv26 = 1;
    117: op1_01_inv26 = 1;
    119: op1_01_inv26 = 1;
    122: op1_01_inv26 = 1;
    123: op1_01_inv26 = 1;
    124: op1_01_inv26 = 1;
    125: op1_01_inv26 = 1;
    131: op1_01_inv26 = 1;
    default: op1_01_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の27番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in27 = reg_0880;
    53: op1_01_in27 = reg_0802;
    67: op1_01_in27 = reg_0464;
    119: op1_01_in27 = reg_0464;
    61: op1_01_in27 = reg_1139;
    72: op1_01_in27 = reg_0726;
    68: op1_01_in27 = reg_0493;
    55: op1_01_in27 = reg_0392;
    73: op1_01_in27 = reg_0491;
    71: op1_01_in27 = reg_0401;
    115: op1_01_in27 = reg_0401;
    48: op1_01_in27 = reg_0235;
    86: op1_01_in27 = reg_1502;
    69: op1_01_in27 = reg_0487;
    59: op1_01_in27 = reg_0967;
    50: op1_01_in27 = reg_0312;
    60: op1_01_in27 = reg_0411;
    46: op1_01_in27 = reg_0940;
    74: op1_01_in27 = reg_1303;
    121: op1_01_in27 = reg_1303;
    75: op1_01_in27 = reg_0328;
    44: op1_01_in27 = reg_0130;
    39: op1_01_in27 = reg_0130;
    56: op1_01_in27 = reg_0173;
    87: op1_01_in27 = reg_0589;
    76: op1_01_in27 = reg_0715;
    57: op1_01_in27 = reg_0123;
    70: op1_01_in27 = reg_1312;
    77: op1_01_in27 = reg_0192;
    88: op1_01_in27 = reg_1104;
    78: op1_01_in27 = reg_0278;
    42: op1_01_in27 = reg_0012;
    79: op1_01_in27 = reg_0165;
    35: op1_01_in27 = reg_0307;
    62: op1_01_in27 = reg_0253;
    80: op1_01_in27 = reg_0148;
    81: op1_01_in27 = reg_1457;
    89: op1_01_in27 = reg_0799;
    63: op1_01_in27 = reg_0587;
    82: op1_01_in27 = reg_0743;
    83: op1_01_in27 = reg_0216;
    64: op1_01_in27 = reg_0952;
    84: op1_01_in27 = reg_0365;
    65: op1_01_in27 = reg_1093;
    85: op1_01_in27 = reg_0011;
    90: op1_01_in27 = reg_1258;
    66: op1_01_in27 = reg_0899;
    91: op1_01_in27 = reg_0577;
    92: op1_01_in27 = reg_0875;
    93: op1_01_in27 = imem06_in[7:4];
    94: op1_01_in27 = reg_0348;
    95: op1_01_in27 = reg_0548;
    96: op1_01_in27 = reg_0016;
    97: op1_01_in27 = reg_0097;
    98: op1_01_in27 = reg_0747;
    100: op1_01_in27 = reg_0261;
    101: op1_01_in27 = reg_0549;
    102: op1_01_in27 = reg_0213;
    104: op1_01_in27 = reg_0239;
    105: op1_01_in27 = reg_0340;
    106: op1_01_in27 = reg_1040;
    107: op1_01_in27 = reg_1326;
    109: op1_01_in27 = reg_0636;
    110: op1_01_in27 = reg_0824;
    111: op1_01_in27 = reg_0457;
    112: op1_01_in27 = reg_1447;
    113: op1_01_in27 = reg_0591;
    114: op1_01_in27 = reg_1403;
    116: op1_01_in27 = reg_0143;
    117: op1_01_in27 = reg_0077;
    118: op1_01_in27 = reg_0434;
    43: op1_01_in27 = reg_0449;
    120: op1_01_in27 = reg_1077;
    122: op1_01_in27 = reg_0026;
    123: op1_01_in27 = reg_0993;
    124: op1_01_in27 = reg_0210;
    125: op1_01_in27 = imem02_in[3:0];
    126: op1_01_in27 = reg_0332;
    127: op1_01_in27 = imem02_in[15:12];
    128: op1_01_in27 = reg_0964;
    129: op1_01_in27 = reg_0086;
    130: op1_01_in27 = reg_0079;
    131: op1_01_in27 = reg_0665;
    default: op1_01_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_01_inv27 = 1;
    53: op1_01_inv27 = 1;
    72: op1_01_inv27 = 1;
    73: op1_01_inv27 = 1;
    71: op1_01_inv27 = 1;
    48: op1_01_inv27 = 1;
    59: op1_01_inv27 = 1;
    60: op1_01_inv27 = 1;
    44: op1_01_inv27 = 1;
    56: op1_01_inv27 = 1;
    57: op1_01_inv27 = 1;
    88: op1_01_inv27 = 1;
    78: op1_01_inv27 = 1;
    42: op1_01_inv27 = 1;
    35: op1_01_inv27 = 1;
    80: op1_01_inv27 = 1;
    89: op1_01_inv27 = 1;
    82: op1_01_inv27 = 1;
    83: op1_01_inv27 = 1;
    39: op1_01_inv27 = 1;
    64: op1_01_inv27 = 1;
    84: op1_01_inv27 = 1;
    65: op1_01_inv27 = 1;
    85: op1_01_inv27 = 1;
    66: op1_01_inv27 = 1;
    91: op1_01_inv27 = 1;
    93: op1_01_inv27 = 1;
    94: op1_01_inv27 = 1;
    96: op1_01_inv27 = 1;
    97: op1_01_inv27 = 1;
    98: op1_01_inv27 = 1;
    100: op1_01_inv27 = 1;
    101: op1_01_inv27 = 1;
    104: op1_01_inv27 = 1;
    105: op1_01_inv27 = 1;
    106: op1_01_inv27 = 1;
    107: op1_01_inv27 = 1;
    109: op1_01_inv27 = 1;
    110: op1_01_inv27 = 1;
    112: op1_01_inv27 = 1;
    113: op1_01_inv27 = 1;
    114: op1_01_inv27 = 1;
    115: op1_01_inv27 = 1;
    117: op1_01_inv27 = 1;
    126: op1_01_inv27 = 1;
    127: op1_01_inv27 = 1;
    129: op1_01_inv27 = 1;
    130: op1_01_inv27 = 1;
    131: op1_01_inv27 = 1;
    default: op1_01_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の28番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in28 = reg_0328;
    53: op1_01_in28 = reg_1132;
    67: op1_01_in28 = reg_0421;
    61: op1_01_in28 = reg_1260;
    72: op1_01_in28 = reg_0899;
    68: op1_01_in28 = reg_0252;
    55: op1_01_in28 = reg_0996;
    73: op1_01_in28 = reg_1416;
    71: op1_01_in28 = reg_0895;
    48: op1_01_in28 = reg_0349;
    86: op1_01_in28 = reg_0175;
    69: op1_01_in28 = reg_0368;
    59: op1_01_in28 = reg_0968;
    50: op1_01_in28 = reg_0734;
    60: op1_01_in28 = reg_0247;
    91: op1_01_in28 = reg_0247;
    46: op1_01_in28 = reg_0090;
    74: op1_01_in28 = reg_0636;
    121: op1_01_in28 = reg_0636;
    75: op1_01_in28 = reg_0444;
    44: op1_01_in28 = reg_0272;
    56: op1_01_in28 = reg_0392;
    87: op1_01_in28 = reg_0151;
    43: op1_01_in28 = reg_0151;
    76: op1_01_in28 = reg_0434;
    57: op1_01_in28 = reg_0124;
    70: op1_01_in28 = reg_0534;
    77: op1_01_in28 = reg_1420;
    88: op1_01_in28 = reg_0182;
    78: op1_01_in28 = reg_0043;
    42: op1_01_in28 = reg_0446;
    79: op1_01_in28 = reg_1202;
    35: op1_01_in28 = reg_0154;
    62: op1_01_in28 = reg_0456;
    80: op1_01_in28 = reg_0727;
    81: op1_01_in28 = reg_0149;
    89: op1_01_in28 = imem06_in[3:0];
    63: op1_01_in28 = reg_0560;
    82: op1_01_in28 = reg_0468;
    83: op1_01_in28 = reg_0145;
    39: op1_01_in28 = reg_0240;
    64: op1_01_in28 = reg_0597;
    84: op1_01_in28 = reg_0874;
    65: op1_01_in28 = reg_1092;
    85: op1_01_in28 = reg_0169;
    90: op1_01_in28 = reg_1083;
    66: op1_01_in28 = reg_0902;
    92: op1_01_in28 = reg_0292;
    93: op1_01_in28 = imem06_in[15:12];
    94: op1_01_in28 = imem04_in[3:0];
    95: op1_01_in28 = reg_0610;
    96: op1_01_in28 = reg_0021;
    97: op1_01_in28 = reg_0862;
    98: op1_01_in28 = reg_0239;
    100: op1_01_in28 = reg_0177;
    101: op1_01_in28 = reg_0743;
    102: op1_01_in28 = reg_0015;
    104: op1_01_in28 = reg_0572;
    105: op1_01_in28 = reg_0262;
    106: op1_01_in28 = reg_0033;
    107: op1_01_in28 = reg_1467;
    109: op1_01_in28 = reg_0398;
    110: op1_01_in28 = reg_0227;
    111: op1_01_in28 = reg_0139;
    112: op1_01_in28 = reg_0178;
    113: op1_01_in28 = reg_0050;
    114: op1_01_in28 = reg_0938;
    115: op1_01_in28 = reg_0553;
    116: op1_01_in28 = reg_0891;
    117: op1_01_in28 = reg_0162;
    118: op1_01_in28 = reg_1513;
    119: op1_01_in28 = reg_0335;
    120: op1_01_in28 = reg_1419;
    122: op1_01_in28 = imem01_in[7:4];
    123: op1_01_in28 = reg_1055;
    124: op1_01_in28 = imem05_in[7:4];
    125: op1_01_in28 = imem02_in[15:12];
    126: op1_01_in28 = reg_0890;
    127: op1_01_in28 = reg_0846;
    128: op1_01_in28 = reg_1516;
    129: op1_01_in28 = reg_0483;
    130: op1_01_in28 = reg_0257;
    131: op1_01_in28 = reg_0442;
    default: op1_01_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_01_inv28 = 1;
    67: op1_01_inv28 = 1;
    61: op1_01_inv28 = 1;
    55: op1_01_inv28 = 1;
    71: op1_01_inv28 = 1;
    48: op1_01_inv28 = 1;
    69: op1_01_inv28 = 1;
    59: op1_01_inv28 = 1;
    60: op1_01_inv28 = 1;
    46: op1_01_inv28 = 1;
    74: op1_01_inv28 = 1;
    75: op1_01_inv28 = 1;
    44: op1_01_inv28 = 1;
    87: op1_01_inv28 = 1;
    76: op1_01_inv28 = 1;
    57: op1_01_inv28 = 1;
    42: op1_01_inv28 = 1;
    80: op1_01_inv28 = 1;
    81: op1_01_inv28 = 1;
    89: op1_01_inv28 = 1;
    83: op1_01_inv28 = 1;
    64: op1_01_inv28 = 1;
    65: op1_01_inv28 = 1;
    85: op1_01_inv28 = 1;
    91: op1_01_inv28 = 1;
    94: op1_01_inv28 = 1;
    95: op1_01_inv28 = 1;
    97: op1_01_inv28 = 1;
    101: op1_01_inv28 = 1;
    105: op1_01_inv28 = 1;
    107: op1_01_inv28 = 1;
    109: op1_01_inv28 = 1;
    110: op1_01_inv28 = 1;
    114: op1_01_inv28 = 1;
    118: op1_01_inv28 = 1;
    119: op1_01_inv28 = 1;
    121: op1_01_inv28 = 1;
    122: op1_01_inv28 = 1;
    123: op1_01_inv28 = 1;
    124: op1_01_inv28 = 1;
    125: op1_01_inv28 = 1;
    126: op1_01_inv28 = 1;
    127: op1_01_inv28 = 1;
    129: op1_01_inv28 = 1;
    130: op1_01_inv28 = 1;
    default: op1_01_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の29番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in29 = reg_0849;
    53: op1_01_in29 = reg_0311;
    67: op1_01_in29 = reg_0414;
    61: op1_01_in29 = reg_0997;
    72: op1_01_in29 = reg_0724;
    68: op1_01_in29 = reg_1147;
    55: op1_01_in29 = reg_0565;
    73: op1_01_in29 = reg_0245;
    71: op1_01_in29 = reg_0874;
    48: op1_01_in29 = reg_0177;
    86: op1_01_in29 = reg_0578;
    69: op1_01_in29 = reg_0835;
    59: op1_01_in29 = reg_0093;
    115: op1_01_in29 = reg_0093;
    50: op1_01_in29 = reg_0678;
    60: op1_01_in29 = imem04_in[15:12];
    46: op1_01_in29 = reg_0168;
    110: op1_01_in29 = reg_0168;
    74: op1_01_in29 = reg_0398;
    75: op1_01_in29 = reg_0557;
    44: op1_01_in29 = reg_0195;
    56: op1_01_in29 = reg_0566;
    87: op1_01_in29 = reg_0861;
    76: op1_01_in29 = reg_1452;
    70: op1_01_in29 = reg_1372;
    77: op1_01_in29 = reg_1509;
    88: op1_01_in29 = reg_0630;
    78: op1_01_in29 = reg_0679;
    42: op1_01_in29 = reg_0589;
    79: op1_01_in29 = reg_0015;
    35: op1_01_in29 = reg_0133;
    62: op1_01_in29 = reg_0455;
    80: op1_01_in29 = reg_0896;
    119: op1_01_in29 = reg_0896;
    81: op1_01_in29 = reg_0400;
    89: op1_01_in29 = reg_1437;
    63: op1_01_in29 = imem02_in[15:12];
    82: op1_01_in29 = reg_0430;
    83: op1_01_in29 = reg_0964;
    39: op1_01_in29 = reg_0251;
    64: op1_01_in29 = reg_1300;
    84: op1_01_in29 = reg_0088;
    65: op1_01_in29 = reg_0882;
    85: op1_01_in29 = reg_0456;
    90: op1_01_in29 = reg_0796;
    66: op1_01_in29 = imem01_in[7:4];
    91: op1_01_in29 = reg_0263;
    92: op1_01_in29 = reg_0335;
    93: op1_01_in29 = reg_1467;
    94: op1_01_in29 = reg_0181;
    95: op1_01_in29 = reg_0238;
    96: op1_01_in29 = imem05_in[3:0];
    97: op1_01_in29 = reg_0836;
    98: op1_01_in29 = reg_0241;
    100: op1_01_in29 = reg_0823;
    101: op1_01_in29 = reg_0612;
    102: op1_01_in29 = imem07_in[7:4];
    104: op1_01_in29 = reg_0434;
    105: op1_01_in29 = reg_0719;
    106: op1_01_in29 = reg_0064;
    107: op1_01_in29 = reg_0110;
    109: op1_01_in29 = reg_0374;
    111: op1_01_in29 = reg_0774;
    112: op1_01_in29 = reg_1208;
    113: op1_01_in29 = reg_0002;
    114: op1_01_in29 = reg_0601;
    116: op1_01_in29 = reg_0789;
    117: op1_01_in29 = reg_0012;
    118: op1_01_in29 = reg_0363;
    43: op1_01_in29 = reg_0037;
    120: op1_01_in29 = reg_0117;
    121: op1_01_in29 = reg_0568;
    122: op1_01_in29 = imem01_in[11:8];
    123: op1_01_in29 = reg_1315;
    124: op1_01_in29 = reg_0538;
    125: op1_01_in29 = reg_0322;
    126: op1_01_in29 = reg_0395;
    127: op1_01_in29 = reg_0588;
    128: op1_01_in29 = reg_1518;
    130: op1_01_in29 = reg_0403;
    131: op1_01_in29 = reg_0741;
    default: op1_01_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    67: op1_01_inv29 = 1;
    61: op1_01_inv29 = 1;
    71: op1_01_inv29 = 1;
    86: op1_01_inv29 = 1;
    69: op1_01_inv29 = 1;
    60: op1_01_inv29 = 1;
    46: op1_01_inv29 = 1;
    74: op1_01_inv29 = 1;
    44: op1_01_inv29 = 1;
    56: op1_01_inv29 = 1;
    87: op1_01_inv29 = 1;
    76: op1_01_inv29 = 1;
    88: op1_01_inv29 = 1;
    78: op1_01_inv29 = 1;
    79: op1_01_inv29 = 1;
    35: op1_01_inv29 = 1;
    80: op1_01_inv29 = 1;
    81: op1_01_inv29 = 1;
    89: op1_01_inv29 = 1;
    63: op1_01_inv29 = 1;
    83: op1_01_inv29 = 1;
    39: op1_01_inv29 = 1;
    65: op1_01_inv29 = 1;
    90: op1_01_inv29 = 1;
    66: op1_01_inv29 = 1;
    91: op1_01_inv29 = 1;
    93: op1_01_inv29 = 1;
    95: op1_01_inv29 = 1;
    98: op1_01_inv29 = 1;
    101: op1_01_inv29 = 1;
    102: op1_01_inv29 = 1;
    104: op1_01_inv29 = 1;
    109: op1_01_inv29 = 1;
    110: op1_01_inv29 = 1;
    114: op1_01_inv29 = 1;
    115: op1_01_inv29 = 1;
    116: op1_01_inv29 = 1;
    121: op1_01_inv29 = 1;
    123: op1_01_inv29 = 1;
    125: op1_01_inv29 = 1;
    126: op1_01_inv29 = 1;
    128: op1_01_inv29 = 1;
    default: op1_01_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の30番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_01_in30 = reg_0000;
    53: op1_01_in30 = reg_0756;
    67: op1_01_in30 = reg_0406;
    61: op1_01_in30 = reg_0473;
    72: op1_01_in30 = reg_0595;
    68: op1_01_in30 = reg_0932;
    55: op1_01_in30 = reg_1181;
    73: op1_01_in30 = reg_0703;
    71: op1_01_in30 = reg_0078;
    48: op1_01_in30 = reg_1000;
    86: op1_01_in30 = reg_0832;
    69: op1_01_in30 = reg_0336;
    59: op1_01_in30 = reg_0277;
    50: op1_01_in30 = reg_0121;
    60: op1_01_in30 = reg_0536;
    46: op1_01_in30 = reg_0864;
    74: op1_01_in30 = reg_0568;
    75: op1_01_in30 = reg_1449;
    44: op1_01_in30 = imem06_in[15:12];
    56: op1_01_in30 = reg_0315;
    87: op1_01_in30 = reg_0828;
    76: op1_01_in30 = reg_1457;
    70: op1_01_in30 = reg_1369;
    77: op1_01_in30 = reg_0863;
    88: op1_01_in30 = reg_0939;
    78: op1_01_in30 = reg_0662;
    42: op1_01_in30 = reg_0587;
    62: op1_01_in30 = reg_0587;
    79: op1_01_in30 = reg_0022;
    35: op1_01_in30 = reg_0007;
    80: op1_01_in30 = reg_0077;
    81: op1_01_in30 = reg_0257;
    89: op1_01_in30 = reg_1334;
    63: op1_01_in30 = reg_0497;
    82: op1_01_in30 = reg_0438;
    104: op1_01_in30 = reg_0438;
    83: op1_01_in30 = reg_0349;
    39: op1_01_in30 = reg_0206;
    64: op1_01_in30 = reg_1199;
    84: op1_01_in30 = reg_1071;
    65: op1_01_in30 = reg_0880;
    85: op1_01_in30 = reg_1344;
    90: op1_01_in30 = reg_1040;
    66: op1_01_in30 = imem01_in[11:8];
    91: op1_01_in30 = reg_1258;
    92: op1_01_in30 = reg_0079;
    93: op1_01_in30 = reg_0860;
    94: op1_01_in30 = reg_0731;
    95: op1_01_in30 = reg_0798;
    96: op1_01_in30 = imem05_in[7:4];
    97: op1_01_in30 = reg_0209;
    98: op1_01_in30 = reg_0742;
    100: op1_01_in30 = reg_0600;
    101: op1_01_in30 = reg_0469;
    102: op1_01_in30 = reg_1414;
    105: op1_01_in30 = reg_1151;
    106: op1_01_in30 = reg_0210;
    107: op1_01_in30 = reg_0141;
    109: op1_01_in30 = reg_0617;
    110: op1_01_in30 = imem03_in[11:8];
    111: op1_01_in30 = reg_0739;
    112: op1_01_in30 = reg_0104;
    113: op1_01_in30 = reg_0052;
    114: op1_01_in30 = reg_0602;
    115: op1_01_in30 = reg_0468;
    116: op1_01_in30 = reg_0070;
    117: op1_01_in30 = imem02_in[3:0];
    118: op1_01_in30 = reg_0901;
    43: op1_01_in30 = reg_0038;
    119: op1_01_in30 = imem02_in[7:4];
    120: op1_01_in30 = reg_0095;
    121: op1_01_in30 = reg_0371;
    122: op1_01_in30 = reg_0269;
    123: op1_01_in30 = reg_0894;
    124: op1_01_in30 = reg_1168;
    125: op1_01_in30 = reg_0659;
    126: op1_01_in30 = reg_0346;
    127: op1_01_in30 = reg_0472;
    128: op1_01_in30 = reg_1313;
    130: op1_01_in30 = reg_0042;
    131: op1_01_in30 = reg_0415;
    default: op1_01_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_01_inv30 = 1;
    72: op1_01_inv30 = 1;
    55: op1_01_inv30 = 1;
    71: op1_01_inv30 = 1;
    69: op1_01_inv30 = 1;
    59: op1_01_inv30 = 1;
    50: op1_01_inv30 = 1;
    46: op1_01_inv30 = 1;
    75: op1_01_inv30 = 1;
    44: op1_01_inv30 = 1;
    56: op1_01_inv30 = 1;
    87: op1_01_inv30 = 1;
    70: op1_01_inv30 = 1;
    77: op1_01_inv30 = 1;
    88: op1_01_inv30 = 1;
    79: op1_01_inv30 = 1;
    63: op1_01_inv30 = 1;
    83: op1_01_inv30 = 1;
    39: op1_01_inv30 = 1;
    84: op1_01_inv30 = 1;
    65: op1_01_inv30 = 1;
    66: op1_01_inv30 = 1;
    91: op1_01_inv30 = 1;
    92: op1_01_inv30 = 1;
    95: op1_01_inv30 = 1;
    96: op1_01_inv30 = 1;
    100: op1_01_inv30 = 1;
    106: op1_01_inv30 = 1;
    107: op1_01_inv30 = 1;
    111: op1_01_inv30 = 1;
    112: op1_01_inv30 = 1;
    114: op1_01_inv30 = 1;
    115: op1_01_inv30 = 1;
    116: op1_01_inv30 = 1;
    117: op1_01_inv30 = 1;
    43: op1_01_inv30 = 1;
    119: op1_01_inv30 = 1;
    120: op1_01_inv30 = 1;
    125: op1_01_inv30 = 1;
    130: op1_01_inv30 = 1;
    131: op1_01_inv30 = 1;
    default: op1_01_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_01_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の0番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in00 = reg_1065;
    53: op1_02_in00 = reg_0184;
    72: op1_02_in00 = reg_1279;
    49: op1_02_in00 = reg_0297;
    55: op1_02_in00 = reg_0582;
    73: op1_02_in00 = reg_0096;
    69: op1_02_in00 = reg_0563;
    86: op1_02_in00 = imem04_in[11:8];
    54: op1_02_in00 = reg_0158;
    59: op1_02_in00 = reg_0824;
    71: op1_02_in00 = reg_0219;
    61: op1_02_in00 = reg_0353;
    50: op1_02_in00 = reg_0614;
    68: op1_02_in00 = reg_1199;
    48: op1_02_in00 = reg_0209;
    74: op1_02_in00 = reg_1404;
    46: op1_02_in00 = reg_0094;
    47: op1_02_in00 = reg_0459;
    75: op1_02_in00 = reg_0724;
    56: op1_02_in00 = reg_1170;
    87: op1_02_in00 = reg_1018;
    37: op1_02_in00 = reg_0286;
    33: op1_02_in00 = imem00_in[11:8];
    103: op1_02_in00 = imem00_in[11:8];
    60: op1_02_in00 = reg_0458;
    76: op1_02_in00 = reg_0836;
    57: op1_02_in00 = reg_0968;
    98: op1_02_in00 = reg_0968;
    101: op1_02_in00 = reg_0968;
    115: op1_02_in00 = reg_0968;
    70: op1_02_in00 = reg_0472;
    77: op1_02_in00 = reg_0827;
    44: op1_02_in00 = reg_0391;
    58: op1_02_in00 = reg_0153;
    88: op1_02_in00 = reg_0847;
    78: op1_02_in00 = reg_0907;
    28: op1_02_in00 = reg_0053;
    51: op1_02_in00 = reg_0489;
    34: op1_02_in00 = imem07_in[3:0];
    79: op1_02_in00 = reg_0332;
    84: op1_02_in00 = reg_0332;
    22: op1_02_in00 = reg_0030;
    42: op1_02_in00 = reg_0581;
    4: op1_02_in00 = imem07_in[15:12];
    80: op1_02_in00 = imem06_in[3:0];
    62: op1_02_in00 = reg_0613;
    81: op1_02_in00 = reg_0077;
    40: op1_02_in00 = reg_0299;
    89: op1_02_in00 = reg_0377;
    63: op1_02_in00 = reg_0555;
    82: op1_02_in00 = reg_1092;
    83: op1_02_in00 = reg_1299;
    64: op1_02_in00 = reg_0885;
    112: op1_02_in00 = reg_0885;
    65: op1_02_in00 = reg_0213;
    85: op1_02_in00 = imem06_in[15:12];
    90: op1_02_in00 = reg_1449;
    66: op1_02_in00 = reg_0561;
    91: op1_02_in00 = imem05_in[3:0];
    67: op1_02_in00 = reg_0161;
    92: op1_02_in00 = reg_0162;
    93: op1_02_in00 = reg_0863;
    94: op1_02_in00 = reg_0694;
    95: op1_02_in00 = reg_0742;
    96: op1_02_in00 = reg_0833;
    97: op1_02_in00 = reg_0536;
    99: op1_02_in00 = imem00_in[7:4];
    100: op1_02_in00 = reg_0191;
    102: op1_02_in00 = reg_0994;
    104: op1_02_in00 = reg_0901;
    105: op1_02_in00 = reg_0117;
    106: op1_02_in00 = reg_0370;
    107: op1_02_in00 = imem00_in[3:0];
    108: op1_02_in00 = imem00_in[3:0];
    109: op1_02_in00 = reg_0323;
    110: op1_02_in00 = reg_0759;
    38: op1_02_in00 = reg_0740;
    111: op1_02_in00 = imem00_in[15:12];
    113: op1_02_in00 = imem00_in[15:12];
    129: op1_02_in00 = imem00_in[15:12];
    131: op1_02_in00 = imem00_in[15:12];
    114: op1_02_in00 = reg_1346;
    29: op1_02_in00 = reg_0156;
    116: op1_02_in00 = reg_1518;
    117: op1_02_in00 = imem02_in[11:8];
    118: op1_02_in00 = reg_0727;
    25: op1_02_in00 = reg_0123;
    119: op1_02_in00 = reg_0889;
    120: op1_02_in00 = imem05_in[15:12];
    5: op1_02_in00 = imem07_in[7:4];
    121: op1_02_in00 = reg_0023;
    122: op1_02_in00 = reg_0871;
    123: op1_02_in00 = reg_0921;
    124: op1_02_in00 = reg_0251;
    125: op1_02_in00 = reg_0712;
    126: op1_02_in00 = reg_0733;
    127: op1_02_in00 = reg_1207;
    43: op1_02_in00 = reg_0414;
    128: op1_02_in00 = reg_0505;
    130: op1_02_in00 = reg_0895;
    default: op1_02_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv00 = 1;
    72: op1_02_inv00 = 1;
    73: op1_02_inv00 = 1;
    69: op1_02_inv00 = 1;
    68: op1_02_inv00 = 1;
    56: op1_02_inv00 = 1;
    87: op1_02_inv00 = 1;
    33: op1_02_inv00 = 1;
    60: op1_02_inv00 = 1;
    76: op1_02_inv00 = 1;
    70: op1_02_inv00 = 1;
    51: op1_02_inv00 = 1;
    22: op1_02_inv00 = 1;
    42: op1_02_inv00 = 1;
    81: op1_02_inv00 = 1;
    89: op1_02_inv00 = 1;
    63: op1_02_inv00 = 1;
    83: op1_02_inv00 = 1;
    65: op1_02_inv00 = 1;
    85: op1_02_inv00 = 1;
    67: op1_02_inv00 = 1;
    92: op1_02_inv00 = 1;
    95: op1_02_inv00 = 1;
    96: op1_02_inv00 = 1;
    97: op1_02_inv00 = 1;
    98: op1_02_inv00 = 1;
    101: op1_02_inv00 = 1;
    105: op1_02_inv00 = 1;
    106: op1_02_inv00 = 1;
    108: op1_02_inv00 = 1;
    110: op1_02_inv00 = 1;
    38: op1_02_inv00 = 1;
    111: op1_02_inv00 = 1;
    113: op1_02_inv00 = 1;
    115: op1_02_inv00 = 1;
    29: op1_02_inv00 = 1;
    116: op1_02_inv00 = 1;
    117: op1_02_inv00 = 1;
    118: op1_02_inv00 = 1;
    25: op1_02_inv00 = 1;
    120: op1_02_inv00 = 1;
    5: op1_02_inv00 = 1;
    121: op1_02_inv00 = 1;
    122: op1_02_inv00 = 1;
    123: op1_02_inv00 = 1;
    124: op1_02_inv00 = 1;
    127: op1_02_inv00 = 1;
    128: op1_02_inv00 = 1;
    129: op1_02_inv00 = 1;
    default: op1_02_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の1番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in01 = reg_0407;
    43: op1_02_in01 = reg_0407;
    53: op1_02_in01 = reg_0039;
    72: op1_02_in01 = reg_1080;
    113: op1_02_in01 = reg_1080;
    131: op1_02_in01 = reg_1080;
    49: op1_02_in01 = reg_0673;
    55: op1_02_in01 = reg_1144;
    73: op1_02_in01 = reg_0675;
    69: op1_02_in01 = reg_0562;
    86: op1_02_in01 = reg_0252;
    54: op1_02_in01 = reg_0031;
    59: op1_02_in01 = reg_1100;
    71: op1_02_in01 = reg_0824;
    62: op1_02_in01 = reg_0824;
    61: op1_02_in01 = reg_0351;
    50: op1_02_in01 = reg_0580;
    68: op1_02_in01 = reg_0178;
    48: op1_02_in01 = reg_0034;
    74: op1_02_in01 = reg_0940;
    46: op1_02_in01 = reg_0021;
    47: op1_02_in01 = reg_0215;
    75: op1_02_in01 = reg_0896;
    56: op1_02_in01 = reg_0191;
    87: op1_02_in01 = reg_0256;
    37: op1_02_in01 = imem07_in[7:4];
    34: op1_02_in01 = imem07_in[7:4];
    33: op1_02_in01 = reg_0524;
    60: op1_02_in01 = imem04_in[15:12];
    76: op1_02_in01 = reg_0096;
    57: op1_02_in01 = reg_0146;
    70: op1_02_in01 = reg_0971;
    127: op1_02_in01 = reg_0971;
    77: op1_02_in01 = reg_0669;
    44: op1_02_in01 = reg_0748;
    58: op1_02_in01 = reg_0877;
    119: op1_02_in01 = reg_0877;
    88: op1_02_in01 = reg_0783;
    78: op1_02_in01 = reg_1277;
    28: op1_02_in01 = imem07_in[3:0];
    22: op1_02_in01 = imem07_in[3:0];
    40: op1_02_in01 = imem07_in[3:0];
    25: op1_02_in01 = imem07_in[3:0];
    51: op1_02_in01 = reg_0465;
    79: op1_02_in01 = reg_1235;
    42: op1_02_in01 = reg_0843;
    80: op1_02_in01 = reg_0115;
    81: op1_02_in01 = reg_0282;
    89: op1_02_in01 = reg_0965;
    63: op1_02_in01 = reg_0615;
    82: op1_02_in01 = reg_0882;
    83: op1_02_in01 = reg_1298;
    64: op1_02_in01 = reg_0505;
    84: op1_02_in01 = reg_0184;
    65: op1_02_in01 = reg_1150;
    85: op1_02_in01 = reg_0860;
    90: op1_02_in01 = reg_0261;
    66: op1_02_in01 = reg_0233;
    91: op1_02_in01 = reg_0206;
    67: op1_02_in01 = reg_0609;
    92: op1_02_in01 = reg_0013;
    93: op1_02_in01 = reg_0827;
    94: op1_02_in01 = reg_0094;
    95: op1_02_in01 = reg_1473;
    96: op1_02_in01 = reg_0272;
    97: op1_02_in01 = reg_0064;
    98: op1_02_in01 = reg_0438;
    99: op1_02_in01 = imem00_in[11:8];
    100: op1_02_in01 = reg_0180;
    101: op1_02_in01 = reg_0148;
    102: op1_02_in01 = reg_0135;
    103: op1_02_in01 = reg_0725;
    104: op1_02_in01 = reg_0875;
    105: op1_02_in01 = reg_1502;
    106: op1_02_in01 = imem05_in[3:0];
    107: op1_02_in01 = reg_0672;
    111: op1_02_in01 = reg_0672;
    108: op1_02_in01 = imem00_in[15:12];
    109: op1_02_in01 = reg_0296;
    110: op1_02_in01 = reg_0823;
    38: op1_02_in01 = reg_0408;
    112: op1_02_in01 = reg_0350;
    114: op1_02_in01 = reg_0344;
    115: op1_02_in01 = reg_0078;
    29: op1_02_in01 = reg_0158;
    116: op1_02_in01 = reg_1313;
    117: op1_02_in01 = reg_0423;
    118: op1_02_in01 = reg_0257;
    120: op1_02_in01 = reg_0708;
    5: op1_02_in01 = imem07_in[15:12];
    121: op1_02_in01 = reg_0046;
    122: op1_02_in01 = reg_0576;
    123: op1_02_in01 = reg_0775;
    124: op1_02_in01 = reg_1059;
    125: op1_02_in01 = reg_0822;
    126: op1_02_in01 = reg_0173;
    128: op1_02_in01 = reg_0756;
    129: op1_02_in01 = reg_1079;
    130: op1_02_in01 = imem02_in[7:4];
    default: op1_02_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_02_inv01 = 1;
    69: op1_02_inv01 = 1;
    54: op1_02_inv01 = 1;
    61: op1_02_inv01 = 1;
    48: op1_02_inv01 = 1;
    75: op1_02_inv01 = 1;
    56: op1_02_inv01 = 1;
    60: op1_02_inv01 = 1;
    76: op1_02_inv01 = 1;
    70: op1_02_inv01 = 1;
    58: op1_02_inv01 = 1;
    78: op1_02_inv01 = 1;
    28: op1_02_inv01 = 1;
    34: op1_02_inv01 = 1;
    22: op1_02_inv01 = 1;
    80: op1_02_inv01 = 1;
    62: op1_02_inv01 = 1;
    89: op1_02_inv01 = 1;
    82: op1_02_inv01 = 1;
    83: op1_02_inv01 = 1;
    91: op1_02_inv01 = 1;
    67: op1_02_inv01 = 1;
    92: op1_02_inv01 = 1;
    97: op1_02_inv01 = 1;
    98: op1_02_inv01 = 1;
    101: op1_02_inv01 = 1;
    104: op1_02_inv01 = 1;
    108: op1_02_inv01 = 1;
    109: op1_02_inv01 = 1;
    110: op1_02_inv01 = 1;
    111: op1_02_inv01 = 1;
    112: op1_02_inv01 = 1;
    113: op1_02_inv01 = 1;
    115: op1_02_inv01 = 1;
    117: op1_02_inv01 = 1;
    118: op1_02_inv01 = 1;
    120: op1_02_inv01 = 1;
    123: op1_02_inv01 = 1;
    125: op1_02_inv01 = 1;
    43: op1_02_inv01 = 1;
    128: op1_02_inv01 = 1;
    130: op1_02_inv01 = 1;
    default: op1_02_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の2番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in02 = reg_0451;
    53: op1_02_in02 = reg_0752;
    72: op1_02_in02 = reg_1078;
    62: op1_02_in02 = reg_1078;
    49: op1_02_in02 = reg_0158;
    55: op1_02_in02 = reg_0534;
    73: op1_02_in02 = reg_0750;
    44: op1_02_in02 = reg_0750;
    69: op1_02_in02 = reg_0433;
    86: op1_02_in02 = reg_1338;
    54: op1_02_in02 = reg_0030;
    25: op1_02_in02 = reg_0030;
    59: op1_02_in02 = imem00_in[7:4];
    71: op1_02_in02 = reg_0791;
    61: op1_02_in02 = reg_0058;
    50: op1_02_in02 = reg_0555;
    68: op1_02_in02 = reg_0506;
    48: op1_02_in02 = reg_0799;
    74: op1_02_in02 = imem05_in[15:12];
    46: op1_02_in02 = reg_0392;
    47: op1_02_in02 = reg_0214;
    75: op1_02_in02 = reg_0290;
    56: op1_02_in02 = reg_1094;
    87: op1_02_in02 = reg_0436;
    37: op1_02_in02 = reg_0408;
    40: op1_02_in02 = reg_0408;
    33: op1_02_in02 = reg_0267;
    60: op1_02_in02 = reg_0535;
    76: op1_02_in02 = reg_0237;
    57: op1_02_in02 = reg_0724;
    70: op1_02_in02 = imem02_in[3:0];
    77: op1_02_in02 = reg_0116;
    80: op1_02_in02 = reg_0116;
    58: op1_02_in02 = reg_0829;
    88: op1_02_in02 = reg_0375;
    100: op1_02_in02 = reg_0375;
    78: op1_02_in02 = reg_1243;
    51: op1_02_in02 = reg_0366;
    123: op1_02_in02 = reg_0366;
    34: op1_02_in02 = reg_0442;
    79: op1_02_in02 = reg_0561;
    22: op1_02_in02 = imem07_in[11:8];
    42: op1_02_in02 = reg_0248;
    81: op1_02_in02 = reg_0044;
    115: op1_02_in02 = reg_0044;
    89: op1_02_in02 = reg_1184;
    63: op1_02_in02 = reg_0445;
    82: op1_02_in02 = reg_0505;
    83: op1_02_in02 = reg_0273;
    64: op1_02_in02 = reg_0348;
    84: op1_02_in02 = reg_0626;
    65: op1_02_in02 = reg_0993;
    85: op1_02_in02 = reg_1035;
    90: op1_02_in02 = reg_1001;
    66: op1_02_in02 = reg_0494;
    91: op1_02_in02 = imem06_in[11:8];
    67: op1_02_in02 = reg_0819;
    92: op1_02_in02 = reg_1071;
    93: op1_02_in02 = reg_1505;
    94: op1_02_in02 = reg_0407;
    95: op1_02_in02 = reg_1475;
    96: op1_02_in02 = reg_1164;
    97: op1_02_in02 = reg_0063;
    98: op1_02_in02 = reg_0727;
    99: op1_02_in02 = reg_1278;
    101: op1_02_in02 = reg_1513;
    102: op1_02_in02 = reg_0219;
    103: op1_02_in02 = reg_1101;
    104: op1_02_in02 = reg_0464;
    105: op1_02_in02 = reg_0370;
    106: op1_02_in02 = imem05_in[7:4];
    107: op1_02_in02 = reg_0638;
    108: op1_02_in02 = reg_0319;
    109: op1_02_in02 = reg_0583;
    110: op1_02_in02 = reg_0311;
    38: op1_02_in02 = reg_0620;
    111: op1_02_in02 = reg_0725;
    112: op1_02_in02 = reg_1009;
    113: op1_02_in02 = reg_0983;
    114: op1_02_in02 = imem06_in[15:12];
    29: op1_02_in02 = reg_0139;
    116: op1_02_in02 = reg_0957;
    117: op1_02_in02 = reg_0056;
    118: op1_02_in02 = reg_0402;
    119: op1_02_in02 = reg_1235;
    120: op1_02_in02 = reg_0833;
    121: op1_02_in02 = reg_0215;
    122: op1_02_in02 = reg_0902;
    124: op1_02_in02 = reg_0340;
    125: op1_02_in02 = reg_0390;
    126: op1_02_in02 = reg_0491;
    127: op1_02_in02 = reg_0973;
    43: op1_02_in02 = reg_0599;
    128: op1_02_in02 = reg_1231;
    129: op1_02_in02 = reg_1279;
    130: op1_02_in02 = reg_0497;
    131: op1_02_in02 = reg_0926;
    default: op1_02_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_02_inv02 = 1;
    86: op1_02_inv02 = 1;
    59: op1_02_inv02 = 1;
    71: op1_02_inv02 = 1;
    50: op1_02_inv02 = 1;
    74: op1_02_inv02 = 1;
    75: op1_02_inv02 = 1;
    87: op1_02_inv02 = 1;
    37: op1_02_inv02 = 1;
    33: op1_02_inv02 = 1;
    60: op1_02_inv02 = 1;
    76: op1_02_inv02 = 1;
    70: op1_02_inv02 = 1;
    77: op1_02_inv02 = 1;
    44: op1_02_inv02 = 1;
    51: op1_02_inv02 = 1;
    34: op1_02_inv02 = 1;
    79: op1_02_inv02 = 1;
    42: op1_02_inv02 = 1;
    80: op1_02_inv02 = 1;
    81: op1_02_inv02 = 1;
    89: op1_02_inv02 = 1;
    83: op1_02_inv02 = 1;
    64: op1_02_inv02 = 1;
    84: op1_02_inv02 = 1;
    85: op1_02_inv02 = 1;
    90: op1_02_inv02 = 1;
    91: op1_02_inv02 = 1;
    67: op1_02_inv02 = 1;
    92: op1_02_inv02 = 1;
    94: op1_02_inv02 = 1;
    95: op1_02_inv02 = 1;
    96: op1_02_inv02 = 1;
    97: op1_02_inv02 = 1;
    98: op1_02_inv02 = 1;
    99: op1_02_inv02 = 1;
    100: op1_02_inv02 = 1;
    102: op1_02_inv02 = 1;
    103: op1_02_inv02 = 1;
    106: op1_02_inv02 = 1;
    108: op1_02_inv02 = 1;
    109: op1_02_inv02 = 1;
    110: op1_02_inv02 = 1;
    38: op1_02_inv02 = 1;
    111: op1_02_inv02 = 1;
    112: op1_02_inv02 = 1;
    115: op1_02_inv02 = 1;
    116: op1_02_inv02 = 1;
    117: op1_02_inv02 = 1;
    25: op1_02_inv02 = 1;
    119: op1_02_inv02 = 1;
    120: op1_02_inv02 = 1;
    121: op1_02_inv02 = 1;
    122: op1_02_inv02 = 1;
    123: op1_02_inv02 = 1;
    127: op1_02_inv02 = 1;
    128: op1_02_inv02 = 1;
    129: op1_02_inv02 = 1;
    130: op1_02_inv02 = 1;
    131: op1_02_inv02 = 1;
    default: op1_02_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の3番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in03 = reg_0319;
    53: op1_02_in03 = reg_0780;
    72: op1_02_in03 = reg_0841;
    49: op1_02_in03 = reg_0157;
    55: op1_02_in03 = reg_0268;
    73: op1_02_in03 = reg_1299;
    69: op1_02_in03 = reg_0126;
    127: op1_02_in03 = reg_0126;
    86: op1_02_in03 = reg_1257;
    54: op1_02_in03 = reg_0592;
    59: op1_02_in03 = imem00_in[11:8];
    71: op1_02_in03 = reg_0672;
    99: op1_02_in03 = reg_0672;
    61: op1_02_in03 = reg_0089;
    50: op1_02_in03 = reg_0844;
    68: op1_02_in03 = imem03_in[15:12];
    48: op1_02_in03 = reg_0749;
    74: op1_02_in03 = reg_0090;
    46: op1_02_in03 = reg_0745;
    47: op1_02_in03 = imem07_in[7:4];
    121: op1_02_in03 = imem07_in[7:4];
    75: op1_02_in03 = reg_0277;
    56: op1_02_in03 = reg_1057;
    87: op1_02_in03 = reg_1458;
    37: op1_02_in03 = reg_0415;
    33: op1_02_in03 = reg_0249;
    60: op1_02_in03 = reg_0263;
    76: op1_02_in03 = reg_0064;
    57: op1_02_in03 = reg_0871;
    70: op1_02_in03 = imem02_in[11:8];
    77: op1_02_in03 = reg_0636;
    44: op1_02_in03 = reg_0346;
    83: op1_02_in03 = reg_0346;
    58: op1_02_in03 = reg_0325;
    88: op1_02_in03 = reg_0964;
    78: op1_02_in03 = reg_1241;
    51: op1_02_in03 = reg_0740;
    34: op1_02_in03 = reg_0404;
    79: op1_02_in03 = reg_0055;
    22: op1_02_in03 = reg_0051;
    42: op1_02_in03 = reg_0725;
    80: op1_02_in03 = reg_0586;
    62: op1_02_in03 = reg_1027;
    81: op1_02_in03 = reg_0662;
    40: op1_02_in03 = reg_0413;
    89: op1_02_in03 = reg_0070;
    63: op1_02_in03 = reg_1278;
    107: op1_02_in03 = reg_1278;
    82: op1_02_in03 = reg_0480;
    64: op1_02_in03 = reg_0425;
    84: op1_02_in03 = reg_0845;
    65: op1_02_in03 = imem07_in[11:8];
    85: op1_02_in03 = reg_0718;
    93: op1_02_in03 = reg_0718;
    90: op1_02_in03 = reg_0143;
    66: op1_02_in03 = reg_0429;
    91: op1_02_in03 = reg_0825;
    67: op1_02_in03 = reg_0438;
    95: op1_02_in03 = reg_0438;
    92: op1_02_in03 = imem02_in[7:4];
    94: op1_02_in03 = reg_0471;
    96: op1_02_in03 = reg_0992;
    97: op1_02_in03 = reg_0065;
    98: op1_02_in03 = reg_0400;
    104: op1_02_in03 = reg_0400;
    100: op1_02_in03 = reg_1494;
    101: op1_02_in03 = reg_0362;
    102: op1_02_in03 = reg_1056;
    103: op1_02_in03 = reg_1487;
    105: op1_02_in03 = imem05_in[15:12];
    106: op1_02_in03 = reg_0833;
    108: op1_02_in03 = reg_1281;
    109: op1_02_in03 = reg_0023;
    110: op1_02_in03 = reg_0312;
    38: op1_02_in03 = reg_0123;
    111: op1_02_in03 = reg_1490;
    131: op1_02_in03 = reg_1490;
    112: op1_02_in03 = imem04_in[3:0];
    113: op1_02_in03 = reg_0805;
    114: op1_02_in03 = reg_1437;
    115: op1_02_in03 = reg_0012;
    29: op1_02_in03 = reg_0465;
    116: op1_02_in03 = reg_0952;
    117: op1_02_in03 = reg_1493;
    118: op1_02_in03 = reg_1071;
    25: op1_02_in03 = reg_0102;
    119: op1_02_in03 = reg_0588;
    120: op1_02_in03 = reg_0205;
    122: op1_02_in03 = reg_0163;
    123: op1_02_in03 = reg_0739;
    124: op1_02_in03 = reg_0649;
    125: op1_02_in03 = reg_0472;
    126: op1_02_in03 = reg_0131;
    43: op1_02_in03 = imem04_in[7:4];
    128: op1_02_in03 = reg_0885;
    129: op1_02_in03 = reg_0501;
    130: op1_02_in03 = reg_0533;
    default: op1_02_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv03 = 1;
    72: op1_02_inv03 = 1;
    73: op1_02_inv03 = 1;
    69: op1_02_inv03 = 1;
    59: op1_02_inv03 = 1;
    61: op1_02_inv03 = 1;
    50: op1_02_inv03 = 1;
    68: op1_02_inv03 = 1;
    48: op1_02_inv03 = 1;
    46: op1_02_inv03 = 1;
    47: op1_02_inv03 = 1;
    56: op1_02_inv03 = 1;
    87: op1_02_inv03 = 1;
    60: op1_02_inv03 = 1;
    76: op1_02_inv03 = 1;
    57: op1_02_inv03 = 1;
    44: op1_02_inv03 = 1;
    58: op1_02_inv03 = 1;
    51: op1_02_inv03 = 1;
    34: op1_02_inv03 = 1;
    79: op1_02_inv03 = 1;
    80: op1_02_inv03 = 1;
    62: op1_02_inv03 = 1;
    81: op1_02_inv03 = 1;
    89: op1_02_inv03 = 1;
    84: op1_02_inv03 = 1;
    85: op1_02_inv03 = 1;
    94: op1_02_inv03 = 1;
    95: op1_02_inv03 = 1;
    96: op1_02_inv03 = 1;
    99: op1_02_inv03 = 1;
    101: op1_02_inv03 = 1;
    102: op1_02_inv03 = 1;
    104: op1_02_inv03 = 1;
    105: op1_02_inv03 = 1;
    108: op1_02_inv03 = 1;
    113: op1_02_inv03 = 1;
    115: op1_02_inv03 = 1;
    118: op1_02_inv03 = 1;
    25: op1_02_inv03 = 1;
    119: op1_02_inv03 = 1;
    121: op1_02_inv03 = 1;
    123: op1_02_inv03 = 1;
    124: op1_02_inv03 = 1;
    125: op1_02_inv03 = 1;
    126: op1_02_inv03 = 1;
    43: op1_02_inv03 = 1;
    130: op1_02_inv03 = 1;
    131: op1_02_inv03 = 1;
    default: op1_02_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の4番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in04 = reg_0208;
    53: op1_02_in04 = reg_0784;
    72: op1_02_in04 = imem00_in[7:4];
    49: op1_02_in04 = imem07_in[3:0];
    54: op1_02_in04 = imem07_in[3:0];
    55: op1_02_in04 = reg_0462;
    73: op1_02_in04 = reg_1430;
    69: op1_02_in04 = imem02_in[11:8];
    86: op1_02_in04 = reg_0488;
    59: op1_02_in04 = reg_1242;
    71: op1_02_in04 = reg_0866;
    61: op1_02_in04 = imem01_in[11:8];
    50: op1_02_in04 = reg_0821;
    68: op1_02_in04 = reg_0790;
    48: op1_02_in04 = reg_0701;
    74: op1_02_in04 = reg_1485;
    46: op1_02_in04 = reg_0733;
    47: op1_02_in04 = reg_0703;
    75: op1_02_in04 = reg_0043;
    56: op1_02_in04 = reg_0668;
    87: op1_02_in04 = reg_1455;
    37: op1_02_in04 = reg_0618;
    33: op1_02_in04 = reg_0250;
    60: op1_02_in04 = reg_0493;
    76: op1_02_in04 = reg_0063;
    57: op1_02_in04 = reg_0080;
    70: op1_02_in04 = reg_0105;
    77: op1_02_in04 = reg_0374;
    44: op1_02_in04 = reg_0173;
    58: op1_02_in04 = reg_0280;
    88: op1_02_in04 = reg_0142;
    78: op1_02_in04 = reg_1471;
    51: op1_02_in04 = reg_0415;
    34: op1_02_in04 = reg_0415;
    79: op1_02_in04 = reg_0255;
    42: op1_02_in04 = reg_0172;
    80: op1_02_in04 = reg_0619;
    62: op1_02_in04 = reg_0405;
    81: op1_02_in04 = reg_1493;
    40: op1_02_in04 = reg_0593;
    89: op1_02_in04 = reg_0627;
    63: op1_02_in04 = reg_1279;
    82: op1_02_in04 = reg_0831;
    83: op1_02_in04 = imem05_in[3:0];
    97: op1_02_in04 = imem05_in[3:0];
    64: op1_02_in04 = reg_1340;
    84: op1_02_in04 = reg_0456;
    65: op1_02_in04 = reg_0674;
    85: op1_02_in04 = reg_1303;
    90: op1_02_in04 = reg_0789;
    66: op1_02_in04 = reg_0776;
    91: op1_02_in04 = reg_0795;
    67: op1_02_in04 = reg_0147;
    92: op1_02_in04 = reg_0169;
    93: op1_02_in04 = reg_0636;
    94: op1_02_in04 = reg_0537;
    95: op1_02_in04 = reg_1457;
    96: op1_02_in04 = reg_0649;
    98: op1_02_in04 = reg_0662;
    99: op1_02_in04 = reg_0616;
    100: op1_02_in04 = reg_0965;
    101: op1_02_in04 = reg_0727;
    102: op1_02_in04 = reg_0170;
    103: op1_02_in04 = reg_0615;
    104: op1_02_in04 = reg_0728;
    105: op1_02_in04 = reg_0986;
    106: op1_02_in04 = reg_1431;
    107: op1_02_in04 = reg_0804;
    108: op1_02_in04 = reg_1278;
    109: op1_02_in04 = imem07_in[11:8];
    121: op1_02_in04 = imem07_in[11:8];
    110: op1_02_in04 = reg_0191;
    38: op1_02_in04 = reg_0124;
    111: op1_02_in04 = reg_0907;
    131: op1_02_in04 = reg_0907;
    112: op1_02_in04 = reg_1368;
    113: op1_02_in04 = reg_0640;
    114: op1_02_in04 = reg_0751;
    115: op1_02_in04 = imem02_in[15:12];
    118: op1_02_in04 = imem02_in[15:12];
    29: op1_02_in04 = reg_0103;
    116: op1_02_in04 = reg_0329;
    117: op1_02_in04 = reg_0532;
    25: op1_02_in04 = reg_0028;
    119: op1_02_in04 = reg_0778;
    120: op1_02_in04 = reg_0700;
    122: op1_02_in04 = reg_0548;
    123: op1_02_in04 = reg_0408;
    124: op1_02_in04 = reg_0066;
    125: op1_02_in04 = reg_0494;
    126: op1_02_in04 = reg_1403;
    127: op1_02_in04 = reg_0628;
    43: op1_02_in04 = reg_0199;
    128: op1_02_in04 = reg_0638;
    129: op1_02_in04 = reg_1052;
    130: op1_02_in04 = reg_0436;
    default: op1_02_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv04 = 1;
    53: op1_02_inv04 = 1;
    72: op1_02_inv04 = 1;
    73: op1_02_inv04 = 1;
    54: op1_02_inv04 = 1;
    59: op1_02_inv04 = 1;
    74: op1_02_inv04 = 1;
    46: op1_02_inv04 = 1;
    47: op1_02_inv04 = 1;
    75: op1_02_inv04 = 1;
    33: op1_02_inv04 = 1;
    60: op1_02_inv04 = 1;
    77: op1_02_inv04 = 1;
    58: op1_02_inv04 = 1;
    88: op1_02_inv04 = 1;
    34: op1_02_inv04 = 1;
    80: op1_02_inv04 = 1;
    62: op1_02_inv04 = 1;
    81: op1_02_inv04 = 1;
    89: op1_02_inv04 = 1;
    64: op1_02_inv04 = 1;
    65: op1_02_inv04 = 1;
    85: op1_02_inv04 = 1;
    90: op1_02_inv04 = 1;
    66: op1_02_inv04 = 1;
    91: op1_02_inv04 = 1;
    94: op1_02_inv04 = 1;
    96: op1_02_inv04 = 1;
    97: op1_02_inv04 = 1;
    98: op1_02_inv04 = 1;
    100: op1_02_inv04 = 1;
    101: op1_02_inv04 = 1;
    104: op1_02_inv04 = 1;
    106: op1_02_inv04 = 1;
    107: op1_02_inv04 = 1;
    109: op1_02_inv04 = 1;
    110: op1_02_inv04 = 1;
    113: op1_02_inv04 = 1;
    114: op1_02_inv04 = 1;
    115: op1_02_inv04 = 1;
    29: op1_02_inv04 = 1;
    25: op1_02_inv04 = 1;
    120: op1_02_inv04 = 1;
    121: op1_02_inv04 = 1;
    122: op1_02_inv04 = 1;
    123: op1_02_inv04 = 1;
    124: op1_02_inv04 = 1;
    127: op1_02_inv04 = 1;
    128: op1_02_inv04 = 1;
    129: op1_02_inv04 = 1;
    default: op1_02_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の5番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in05 = reg_0062;
    53: op1_02_in05 = reg_0906;
    72: op1_02_in05 = reg_1052;
    113: op1_02_in05 = reg_1052;
    49: op1_02_in05 = reg_0779;
    55: op1_02_in05 = imem04_in[7:4];
    73: op1_02_in05 = reg_1431;
    69: op1_02_in05 = reg_0712;
    86: op1_02_in05 = reg_1147;
    59: op1_02_in05 = reg_1230;
    71: op1_02_in05 = reg_1243;
    61: op1_02_in05 = reg_0175;
    44: op1_02_in05 = reg_0175;
    50: op1_02_in05 = reg_0485;
    68: op1_02_in05 = reg_1383;
    48: op1_02_in05 = imem05_in[3:0];
    74: op1_02_in05 = reg_0601;
    46: op1_02_in05 = reg_0833;
    47: op1_02_in05 = reg_0170;
    65: op1_02_in05 = reg_0170;
    75: op1_02_in05 = reg_0013;
    56: op1_02_in05 = reg_0224;
    87: op1_02_in05 = reg_0382;
    37: op1_02_in05 = reg_0137;
    33: op1_02_in05 = reg_0220;
    42: op1_02_in05 = reg_0220;
    60: op1_02_in05 = reg_1257;
    76: op1_02_in05 = reg_0065;
    57: op1_02_in05 = reg_0042;
    104: op1_02_in05 = reg_0042;
    70: op1_02_in05 = reg_1433;
    77: op1_02_in05 = reg_0979;
    80: op1_02_in05 = reg_0979;
    58: op1_02_in05 = reg_0732;
    88: op1_02_in05 = reg_1516;
    78: op1_02_in05 = reg_0250;
    51: op1_02_in05 = reg_0028;
    34: op1_02_in05 = reg_0413;
    79: op1_02_in05 = reg_1207;
    62: op1_02_in05 = reg_0353;
    81: op1_02_in05 = reg_0590;
    40: op1_02_in05 = reg_0361;
    25: op1_02_in05 = reg_0361;
    89: op1_02_in05 = reg_0048;
    63: op1_02_in05 = reg_1080;
    82: op1_02_in05 = reg_0734;
    83: op1_02_in05 = reg_1104;
    64: op1_02_in05 = reg_1200;
    84: op1_02_in05 = reg_0608;
    85: op1_02_in05 = reg_0141;
    90: op1_02_in05 = reg_0375;
    66: op1_02_in05 = reg_0778;
    130: op1_02_in05 = reg_0778;
    91: op1_02_in05 = reg_0908;
    67: op1_02_in05 = reg_0148;
    92: op1_02_in05 = reg_0138;
    93: op1_02_in05 = reg_0398;
    94: op1_02_in05 = reg_0304;
    95: op1_02_in05 = reg_0146;
    96: op1_02_in05 = reg_0392;
    97: op1_02_in05 = reg_0466;
    98: op1_02_in05 = imem02_in[11:8];
    99: op1_02_in05 = reg_0293;
    100: op1_02_in05 = reg_1184;
    101: op1_02_in05 = reg_0257;
    102: op1_02_in05 = reg_0139;
    103: op1_02_in05 = reg_0555;
    105: op1_02_in05 = reg_0367;
    106: op1_02_in05 = reg_0205;
    107: op1_02_in05 = reg_0907;
    108: op1_02_in05 = reg_1490;
    109: op1_02_in05 = reg_0867;
    110: op1_02_in05 = reg_0144;
    111: op1_02_in05 = reg_0554;
    112: op1_02_in05 = reg_0493;
    114: op1_02_in05 = reg_0863;
    115: op1_02_in05 = reg_0659;
    29: op1_02_in05 = reg_0186;
    116: op1_02_in05 = reg_0291;
    117: op1_02_in05 = reg_0822;
    118: op1_02_in05 = reg_0254;
    119: op1_02_in05 = reg_0127;
    120: op1_02_in05 = reg_0562;
    121: op1_02_in05 = reg_0498;
    122: op1_02_in05 = reg_0610;
    123: op1_02_in05 = reg_0621;
    124: op1_02_in05 = reg_0630;
    125: op1_02_in05 = reg_0326;
    126: op1_02_in05 = reg_0301;
    127: op1_02_in05 = reg_0380;
    43: op1_02_in05 = reg_0016;
    128: op1_02_in05 = reg_1280;
    129: op1_02_in05 = reg_0221;
    131: op1_02_in05 = reg_0248;
    default: op1_02_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv05 = 1;
    72: op1_02_inv05 = 1;
    55: op1_02_inv05 = 1;
    69: op1_02_inv05 = 1;
    86: op1_02_inv05 = 1;
    59: op1_02_inv05 = 1;
    61: op1_02_inv05 = 1;
    68: op1_02_inv05 = 1;
    75: op1_02_inv05 = 1;
    56: op1_02_inv05 = 1;
    87: op1_02_inv05 = 1;
    33: op1_02_inv05 = 1;
    60: op1_02_inv05 = 1;
    76: op1_02_inv05 = 1;
    57: op1_02_inv05 = 1;
    70: op1_02_inv05 = 1;
    77: op1_02_inv05 = 1;
    78: op1_02_inv05 = 1;
    34: op1_02_inv05 = 1;
    79: op1_02_inv05 = 1;
    42: op1_02_inv05 = 1;
    62: op1_02_inv05 = 1;
    81: op1_02_inv05 = 1;
    63: op1_02_inv05 = 1;
    64: op1_02_inv05 = 1;
    85: op1_02_inv05 = 1;
    66: op1_02_inv05 = 1;
    67: op1_02_inv05 = 1;
    93: op1_02_inv05 = 1;
    94: op1_02_inv05 = 1;
    99: op1_02_inv05 = 1;
    100: op1_02_inv05 = 1;
    101: op1_02_inv05 = 1;
    102: op1_02_inv05 = 1;
    103: op1_02_inv05 = 1;
    106: op1_02_inv05 = 1;
    109: op1_02_inv05 = 1;
    110: op1_02_inv05 = 1;
    112: op1_02_inv05 = 1;
    113: op1_02_inv05 = 1;
    114: op1_02_inv05 = 1;
    29: op1_02_inv05 = 1;
    124: op1_02_inv05 = 1;
    128: op1_02_inv05 = 1;
    130: op1_02_inv05 = 1;
    default: op1_02_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の6番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in06 = reg_0020;
    43: op1_02_in06 = reg_0020;
    53: op1_02_in06 = reg_0398;
    72: op1_02_in06 = reg_1417;
    49: op1_02_in06 = reg_0775;
    55: op1_02_in06 = imem04_in[15:12];
    73: op1_02_in06 = reg_0136;
    69: op1_02_in06 = reg_0711;
    86: op1_02_in06 = reg_0412;
    59: op1_02_in06 = reg_0203;
    71: op1_02_in06 = reg_1244;
    61: op1_02_in06 = reg_1290;
    50: op1_02_in06 = reg_0202;
    68: op1_02_in06 = reg_1216;
    48: op1_02_in06 = imem05_in[11:8];
    74: op1_02_in06 = reg_0274;
    46: op1_02_in06 = reg_0174;
    47: op1_02_in06 = reg_0309;
    75: op1_02_in06 = reg_0679;
    56: op1_02_in06 = reg_0894;
    87: op1_02_in06 = reg_1032;
    37: op1_02_in06 = reg_0592;
    33: op1_02_in06 = reg_0221;
    113: op1_02_in06 = reg_0221;
    60: op1_02_in06 = reg_1214;
    76: op1_02_in06 = reg_0370;
    57: op1_02_in06 = reg_0662;
    70: op1_02_in06 = reg_0390;
    84: op1_02_in06 = reg_0390;
    77: op1_02_in06 = reg_1204;
    44: op1_02_in06 = reg_0648;
    58: op1_02_in06 = reg_0573;
    88: op1_02_in06 = reg_0597;
    78: op1_02_in06 = reg_1230;
    129: op1_02_in06 = reg_1230;
    51: op1_02_in06 = reg_0001;
    34: op1_02_in06 = reg_0623;
    79: op1_02_in06 = reg_1450;
    42: op1_02_in06 = reg_0188;
    80: op1_02_in06 = reg_0244;
    62: op1_02_in06 = reg_0351;
    81: op1_02_in06 = reg_1103;
    40: op1_02_in06 = reg_0003;
    89: op1_02_in06 = reg_0329;
    63: op1_02_in06 = reg_1081;
    82: op1_02_in06 = reg_1312;
    83: op1_02_in06 = reg_0986;
    64: op1_02_in06 = reg_0676;
    65: op1_02_in06 = reg_1345;
    85: op1_02_in06 = reg_0373;
    90: op1_02_in06 = reg_1517;
    66: op1_02_in06 = reg_0934;
    115: op1_02_in06 = reg_0934;
    91: op1_02_in06 = reg_0905;
    67: op1_02_in06 = reg_0146;
    92: op1_02_in06 = reg_0561;
    93: op1_02_in06 = reg_0374;
    94: op1_02_in06 = reg_0305;
    95: op1_02_in06 = reg_0365;
    96: op1_02_in06 = reg_0564;
    97: op1_02_in06 = reg_0332;
    98: op1_02_in06 = reg_0456;
    99: op1_02_in06 = reg_0961;
    100: op1_02_in06 = reg_0349;
    101: op1_02_in06 = reg_0042;
    102: op1_02_in06 = reg_0366;
    103: op1_02_in06 = reg_1229;
    104: op1_02_in06 = reg_0044;
    105: op1_02_in06 = reg_0205;
    106: op1_02_in06 = reg_1164;
    107: op1_02_in06 = reg_0841;
    108: op1_02_in06 = reg_0803;
    109: op1_02_in06 = reg_0963;
    110: op1_02_in06 = reg_0180;
    111: op1_02_in06 = reg_1052;
    112: op1_02_in06 = reg_0088;
    114: op1_02_in06 = reg_0859;
    29: op1_02_in06 = reg_0086;
    116: op1_02_in06 = imem04_in[3:0];
    117: op1_02_in06 = reg_0900;
    118: op1_02_in06 = reg_0133;
    25: op1_02_in06 = reg_0228;
    119: op1_02_in06 = reg_1433;
    120: op1_02_in06 = reg_1070;
    124: op1_02_in06 = reg_1070;
    121: op1_02_in06 = reg_0394;
    122: op1_02_in06 = reg_0787;
    123: op1_02_in06 = reg_0618;
    125: op1_02_in06 = reg_0382;
    126: op1_02_in06 = reg_0318;
    127: op1_02_in06 = reg_0829;
    128: op1_02_in06 = imem04_in[11:8];
    130: op1_02_in06 = reg_0970;
    131: op1_02_in06 = reg_0059;
    default: op1_02_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_02_inv06 = 1;
    49: op1_02_inv06 = 1;
    69: op1_02_inv06 = 1;
    86: op1_02_inv06 = 1;
    59: op1_02_inv06 = 1;
    61: op1_02_inv06 = 1;
    50: op1_02_inv06 = 1;
    48: op1_02_inv06 = 1;
    46: op1_02_inv06 = 1;
    47: op1_02_inv06 = 1;
    56: op1_02_inv06 = 1;
    37: op1_02_inv06 = 1;
    33: op1_02_inv06 = 1;
    60: op1_02_inv06 = 1;
    76: op1_02_inv06 = 1;
    57: op1_02_inv06 = 1;
    70: op1_02_inv06 = 1;
    77: op1_02_inv06 = 1;
    58: op1_02_inv06 = 1;
    88: op1_02_inv06 = 1;
    34: op1_02_inv06 = 1;
    42: op1_02_inv06 = 1;
    81: op1_02_inv06 = 1;
    40: op1_02_inv06 = 1;
    89: op1_02_inv06 = 1;
    64: op1_02_inv06 = 1;
    84: op1_02_inv06 = 1;
    65: op1_02_inv06 = 1;
    85: op1_02_inv06 = 1;
    91: op1_02_inv06 = 1;
    67: op1_02_inv06 = 1;
    92: op1_02_inv06 = 1;
    95: op1_02_inv06 = 1;
    96: op1_02_inv06 = 1;
    99: op1_02_inv06 = 1;
    100: op1_02_inv06 = 1;
    104: op1_02_inv06 = 1;
    105: op1_02_inv06 = 1;
    106: op1_02_inv06 = 1;
    107: op1_02_inv06 = 1;
    110: op1_02_inv06 = 1;
    112: op1_02_inv06 = 1;
    115: op1_02_inv06 = 1;
    116: op1_02_inv06 = 1;
    117: op1_02_inv06 = 1;
    25: op1_02_inv06 = 1;
    125: op1_02_inv06 = 1;
    127: op1_02_inv06 = 1;
    128: op1_02_inv06 = 1;
    default: op1_02_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の7番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in07 = imem05_in[3:0];
    53: op1_02_in07 = reg_0863;
    72: op1_02_in07 = reg_0459;
    49: op1_02_in07 = reg_0031;
    55: op1_02_in07 = reg_0414;
    73: op1_02_in07 = reg_1168;
    69: op1_02_in07 = reg_0153;
    108: op1_02_in07 = reg_0153;
    86: op1_02_in07 = reg_1077;
    59: op1_02_in07 = reg_0460;
    99: op1_02_in07 = reg_0460;
    71: op1_02_in07 = reg_0806;
    61: op1_02_in07 = reg_0448;
    50: op1_02_in07 = reg_0203;
    68: op1_02_in07 = reg_1200;
    48: op1_02_in07 = reg_0650;
    44: op1_02_in07 = reg_0650;
    74: op1_02_in07 = reg_0393;
    46: op1_02_in07 = reg_0221;
    47: op1_02_in07 = reg_0674;
    75: op1_02_in07 = reg_1103;
    56: op1_02_in07 = reg_0299;
    87: op1_02_in07 = reg_0307;
    37: op1_02_in07 = reg_0102;
    123: op1_02_in07 = reg_0102;
    33: op1_02_in07 = reg_0202;
    60: op1_02_in07 = reg_1082;
    76: op1_02_in07 = reg_0737;
    57: op1_02_in07 = reg_0254;
    92: op1_02_in07 = reg_0254;
    70: op1_02_in07 = reg_0712;
    77: op1_02_in07 = reg_0583;
    58: op1_02_in07 = reg_0677;
    88: op1_02_in07 = reg_1093;
    78: op1_02_in07 = reg_1418;
    103: op1_02_in07 = reg_1418;
    51: op1_02_in07 = reg_0002;
    34: op1_02_in07 = reg_0618;
    79: op1_02_in07 = reg_0112;
    42: op1_02_in07 = reg_0189;
    80: op1_02_in07 = reg_0270;
    62: op1_02_in07 = reg_0917;
    81: op1_02_in07 = reg_0256;
    89: op1_02_in07 = reg_1301;
    63: op1_02_in07 = reg_1244;
    82: op1_02_in07 = reg_0534;
    83: op1_02_in07 = reg_1514;
    64: op1_02_in07 = reg_0969;
    84: op1_02_in07 = reg_0473;
    65: op1_02_in07 = reg_0158;
    85: op1_02_in07 = reg_0345;
    93: op1_02_in07 = reg_0345;
    90: op1_02_in07 = reg_0314;
    66: op1_02_in07 = reg_0127;
    91: op1_02_in07 = reg_0870;
    67: op1_02_in07 = reg_0402;
    94: op1_02_in07 = reg_0836;
    95: op1_02_in07 = reg_0092;
    96: op1_02_in07 = reg_0302;
    97: op1_02_in07 = reg_0278;
    98: op1_02_in07 = reg_0934;
    100: op1_02_in07 = reg_0597;
    101: op1_02_in07 = imem02_in[3:0];
    102: op1_02_in07 = reg_0591;
    104: op1_02_in07 = reg_0013;
    105: op1_02_in07 = reg_1164;
    106: op1_02_in07 = reg_0831;
    107: op1_02_in07 = reg_0486;
    109: op1_02_in07 = reg_0324;
    110: op1_02_in07 = reg_0556;
    111: op1_02_in07 = reg_1454;
    112: op1_02_in07 = reg_1215;
    113: op1_02_in07 = reg_1405;
    114: op1_02_in07 = reg_1323;
    115: op1_02_in07 = reg_0055;
    29: op1_02_in07 = imem07_in[3:0];
    116: op1_02_in07 = imem04_in[11:8];
    117: op1_02_in07 = reg_0495;
    118: op1_02_in07 = reg_1074;
    25: op1_02_in07 = reg_0135;
    119: op1_02_in07 = reg_0684;
    120: op1_02_in07 = reg_0939;
    121: op1_02_in07 = reg_1095;
    122: op1_02_in07 = reg_0743;
    124: op1_02_in07 = reg_0792;
    125: op1_02_in07 = reg_0496;
    130: op1_02_in07 = reg_0496;
    126: op1_02_in07 = reg_0275;
    127: op1_02_in07 = reg_0745;
    43: op1_02_in07 = reg_0035;
    128: op1_02_in07 = reg_1384;
    129: op1_02_in07 = reg_1205;
    131: op1_02_in07 = reg_0616;
    default: op1_02_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_02_inv07 = 1;
    72: op1_02_inv07 = 1;
    49: op1_02_inv07 = 1;
    55: op1_02_inv07 = 1;
    73: op1_02_inv07 = 1;
    86: op1_02_inv07 = 1;
    71: op1_02_inv07 = 1;
    50: op1_02_inv07 = 1;
    46: op1_02_inv07 = 1;
    47: op1_02_inv07 = 1;
    56: op1_02_inv07 = 1;
    60: op1_02_inv07 = 1;
    76: op1_02_inv07 = 1;
    77: op1_02_inv07 = 1;
    44: op1_02_inv07 = 1;
    88: op1_02_inv07 = 1;
    51: op1_02_inv07 = 1;
    79: op1_02_inv07 = 1;
    42: op1_02_inv07 = 1;
    62: op1_02_inv07 = 1;
    81: op1_02_inv07 = 1;
    63: op1_02_inv07 = 1;
    83: op1_02_inv07 = 1;
    65: op1_02_inv07 = 1;
    85: op1_02_inv07 = 1;
    90: op1_02_inv07 = 1;
    66: op1_02_inv07 = 1;
    67: op1_02_inv07 = 1;
    93: op1_02_inv07 = 1;
    94: op1_02_inv07 = 1;
    95: op1_02_inv07 = 1;
    97: op1_02_inv07 = 1;
    100: op1_02_inv07 = 1;
    104: op1_02_inv07 = 1;
    106: op1_02_inv07 = 1;
    108: op1_02_inv07 = 1;
    110: op1_02_inv07 = 1;
    113: op1_02_inv07 = 1;
    29: op1_02_inv07 = 1;
    116: op1_02_inv07 = 1;
    117: op1_02_inv07 = 1;
    25: op1_02_inv07 = 1;
    120: op1_02_inv07 = 1;
    124: op1_02_inv07 = 1;
    126: op1_02_inv07 = 1;
    128: op1_02_inv07 = 1;
    130: op1_02_inv07 = 1;
    131: op1_02_inv07 = 1;
    default: op1_02_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の8番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in08 = reg_0331;
    53: op1_02_in08 = reg_0374;
    72: op1_02_in08 = reg_1405;
    49: op1_02_in08 = reg_0441;
    55: op1_02_in08 = reg_0407;
    73: op1_02_in08 = reg_0700;
    69: op1_02_in08 = reg_0009;
    86: op1_02_in08 = reg_0305;
    59: op1_02_in08 = reg_0926;
    71: op1_02_in08 = reg_0805;
    61: op1_02_in08 = reg_1291;
    50: op1_02_in08 = reg_0987;
    68: op1_02_in08 = reg_1077;
    48: op1_02_in08 = reg_0992;
    74: op1_02_in08 = reg_0130;
    46: op1_02_in08 = reg_0601;
    47: op1_02_in08 = reg_0157;
    65: op1_02_in08 = reg_0157;
    75: op1_02_in08 = reg_0607;
    56: op1_02_in08 = reg_0170;
    87: op1_02_in08 = reg_0829;
    119: op1_02_in08 = reg_0829;
    37: op1_02_in08 = reg_0103;
    33: op1_02_in08 = reg_0201;
    60: op1_02_in08 = reg_0414;
    76: op1_02_in08 = reg_0395;
    57: op1_02_in08 = reg_0255;
    70: op1_02_in08 = reg_0708;
    77: op1_02_in08 = reg_0269;
    44: op1_02_in08 = reg_0603;
    58: op1_02_in08 = reg_0198;
    88: op1_02_in08 = reg_0880;
    78: op1_02_in08 = reg_0459;
    99: op1_02_in08 = reg_0459;
    129: op1_02_in08 = reg_0459;
    51: op1_02_in08 = reg_0052;
    34: op1_02_in08 = reg_0593;
    79: op1_02_in08 = reg_0106;
    42: op1_02_in08 = reg_0135;
    80: op1_02_in08 = reg_0271;
    62: op1_02_in08 = reg_0785;
    81: op1_02_in08 = reg_0473;
    89: op1_02_in08 = reg_0481;
    63: op1_02_in08 = reg_0803;
    82: op1_02_in08 = reg_0263;
    83: op1_02_in08 = reg_0090;
    96: op1_02_in08 = reg_0090;
    64: op1_02_in08 = reg_0599;
    112: op1_02_in08 = reg_0599;
    84: op1_02_in08 = reg_0326;
    85: op1_02_in08 = reg_0289;
    90: op1_02_in08 = reg_1314;
    66: op1_02_in08 = reg_0126;
    91: op1_02_in08 = reg_1209;
    67: op1_02_in08 = reg_0401;
    92: op1_02_in08 = reg_0712;
    93: op1_02_in08 = reg_0171;
    94: op1_02_in08 = reg_0339;
    95: op1_02_in08 = reg_0595;
    97: op1_02_in08 = reg_0346;
    98: op1_02_in08 = reg_0561;
    100: op1_02_in08 = reg_1301;
    101: op1_02_in08 = imem02_in[7:4];
    102: op1_02_in08 = reg_0100;
    103: op1_02_in08 = reg_1406;
    104: op1_02_in08 = imem02_in[11:8];
    105: op1_02_in08 = reg_0996;
    106: op1_02_in08 = reg_0562;
    107: op1_02_in08 = reg_1053;
    108: op1_02_in08 = reg_1459;
    109: op1_02_in08 = reg_1010;
    110: op1_02_in08 = reg_1184;
    111: op1_02_in08 = reg_0821;
    113: op1_02_in08 = reg_0887;
    114: op1_02_in08 = reg_1504;
    115: op1_02_in08 = reg_0254;
    29: op1_02_in08 = imem07_in[11:8];
    116: op1_02_in08 = reg_0493;
    117: op1_02_in08 = reg_1207;
    118: op1_02_in08 = reg_0497;
    120: op1_02_in08 = reg_1163;
    124: op1_02_in08 = reg_1163;
    121: op1_02_in08 = reg_0993;
    122: op1_02_in08 = reg_0609;
    123: op1_02_in08 = reg_0235;
    125: op1_02_in08 = reg_1433;
    130: op1_02_in08 = reg_1433;
    126: op1_02_in08 = reg_0393;
    127: op1_02_in08 = reg_0801;
    43: op1_02_in08 = reg_0794;
    128: op1_02_in08 = reg_0721;
    131: op1_02_in08 = reg_0486;
    default: op1_02_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_02_inv08 = 1;
    73: op1_02_inv08 = 1;
    69: op1_02_inv08 = 1;
    59: op1_02_inv08 = 1;
    50: op1_02_inv08 = 1;
    47: op1_02_inv08 = 1;
    75: op1_02_inv08 = 1;
    87: op1_02_inv08 = 1;
    76: op1_02_inv08 = 1;
    70: op1_02_inv08 = 1;
    77: op1_02_inv08 = 1;
    44: op1_02_inv08 = 1;
    58: op1_02_inv08 = 1;
    88: op1_02_inv08 = 1;
    34: op1_02_inv08 = 1;
    80: op1_02_inv08 = 1;
    89: op1_02_inv08 = 1;
    82: op1_02_inv08 = 1;
    65: op1_02_inv08 = 1;
    90: op1_02_inv08 = 1;
    91: op1_02_inv08 = 1;
    67: op1_02_inv08 = 1;
    92: op1_02_inv08 = 1;
    100: op1_02_inv08 = 1;
    103: op1_02_inv08 = 1;
    104: op1_02_inv08 = 1;
    106: op1_02_inv08 = 1;
    108: op1_02_inv08 = 1;
    109: op1_02_inv08 = 1;
    111: op1_02_inv08 = 1;
    112: op1_02_inv08 = 1;
    114: op1_02_inv08 = 1;
    118: op1_02_inv08 = 1;
    121: op1_02_inv08 = 1;
    123: op1_02_inv08 = 1;
    125: op1_02_inv08 = 1;
    43: op1_02_inv08 = 1;
    default: op1_02_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の9番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in09 = reg_0175;
    53: op1_02_in09 = reg_0371;
    72: op1_02_in09 = reg_0188;
    49: op1_02_in09 = reg_0741;
    55: op1_02_in09 = reg_0599;
    73: op1_02_in09 = reg_0176;
    105: op1_02_in09 = reg_0176;
    69: op1_02_in09 = reg_0632;
    86: op1_02_in09 = reg_0487;
    59: op1_02_in09 = reg_0886;
    71: op1_02_in09 = reg_0803;
    61: op1_02_in09 = reg_1033;
    50: op1_02_in09 = reg_0926;
    68: op1_02_in09 = reg_0796;
    48: op1_02_in09 = reg_0538;
    74: op1_02_in09 = reg_0118;
    46: op1_02_in09 = reg_0604;
    47: op1_02_in09 = reg_0031;
    75: op1_02_in09 = reg_0455;
    56: op1_02_in09 = reg_0674;
    87: op1_02_in09 = reg_0311;
    37: op1_02_in09 = reg_0321;
    33: op1_02_in09 = reg_0445;
    60: op1_02_in09 = reg_0969;
    76: op1_02_in09 = reg_1259;
    57: op1_02_in09 = reg_0133;
    70: op1_02_in09 = reg_0306;
    77: op1_02_in09 = reg_0067;
    44: op1_02_in09 = reg_0567;
    58: op1_02_in09 = reg_0709;
    88: op1_02_in09 = reg_0350;
    78: op1_02_in09 = reg_0428;
    51: op1_02_in09 = reg_0053;
    123: op1_02_in09 = reg_0053;
    34: op1_02_in09 = reg_0004;
    79: op1_02_in09 = reg_0878;
    42: op1_02_in09 = imem00_in[3:0];
    80: op1_02_in09 = reg_0022;
    62: op1_02_in09 = reg_0166;
    81: op1_02_in09 = reg_0474;
    89: op1_02_in09 = reg_0291;
    63: op1_02_in09 = reg_1028;
    82: op1_02_in09 = reg_0462;
    83: op1_02_in09 = reg_0601;
    64: op1_02_in09 = reg_0451;
    84: op1_02_in09 = reg_0973;
    65: op1_02_in09 = reg_0224;
    85: op1_02_in09 = reg_0270;
    90: op1_02_in09 = reg_1300;
    66: op1_02_in09 = reg_0900;
    91: op1_02_in09 = reg_1509;
    67: op1_02_in09 = reg_0360;
    92: op1_02_in09 = reg_0532;
    93: op1_02_in09 = reg_0289;
    94: op1_02_in09 = reg_1107;
    95: op1_02_in09 = reg_0042;
    96: op1_02_in09 = reg_0275;
    97: op1_02_in09 = reg_1268;
    98: op1_02_in09 = reg_1343;
    99: op1_02_in09 = reg_0435;
    100: op1_02_in09 = reg_1093;
    101: op1_02_in09 = reg_0276;
    102: op1_02_in09 = reg_0114;
    103: op1_02_in09 = reg_1405;
    104: op1_02_in09 = reg_0138;
    106: op1_02_in09 = reg_0173;
    107: op1_02_in09 = reg_0250;
    108: op1_02_in09 = reg_0249;
    109: op1_02_in09 = reg_1315;
    110: op1_02_in09 = reg_0142;
    111: op1_02_in09 = reg_0202;
    113: op1_02_in09 = reg_0202;
    112: op1_02_in09 = reg_0199;
    114: op1_02_in09 = reg_1508;
    115: op1_02_in09 = reg_1493;
    29: op1_02_in09 = reg_0123;
    116: op1_02_in09 = reg_0264;
    117: op1_02_in09 = reg_0429;
    118: op1_02_in09 = reg_0436;
    119: op1_02_in09 = reg_0379;
    120: op1_02_in09 = reg_0888;
    121: op1_02_in09 = reg_0478;
    122: op1_02_in09 = reg_0241;
    124: op1_02_in09 = reg_0418;
    125: op1_02_in09 = reg_0628;
    126: op1_02_in09 = reg_0207;
    127: op1_02_in09 = reg_0848;
    43: op1_02_in09 = reg_0344;
    128: op1_02_in09 = reg_0936;
    129: op1_02_in09 = reg_0928;
    130: op1_02_in09 = reg_0684;
    131: op1_02_in09 = reg_0523;
    default: op1_02_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    49: op1_02_inv09 = 1;
    55: op1_02_inv09 = 1;
    73: op1_02_inv09 = 1;
    50: op1_02_inv09 = 1;
    74: op1_02_inv09 = 1;
    47: op1_02_inv09 = 1;
    75: op1_02_inv09 = 1;
    56: op1_02_inv09 = 1;
    87: op1_02_inv09 = 1;
    37: op1_02_inv09 = 1;
    70: op1_02_inv09 = 1;
    77: op1_02_inv09 = 1;
    44: op1_02_inv09 = 1;
    88: op1_02_inv09 = 1;
    34: op1_02_inv09 = 1;
    42: op1_02_inv09 = 1;
    80: op1_02_inv09 = 1;
    62: op1_02_inv09 = 1;
    63: op1_02_inv09 = 1;
    82: op1_02_inv09 = 1;
    64: op1_02_inv09 = 1;
    84: op1_02_inv09 = 1;
    65: op1_02_inv09 = 1;
    85: op1_02_inv09 = 1;
    90: op1_02_inv09 = 1;
    67: op1_02_inv09 = 1;
    96: op1_02_inv09 = 1;
    98: op1_02_inv09 = 1;
    99: op1_02_inv09 = 1;
    102: op1_02_inv09 = 1;
    103: op1_02_inv09 = 1;
    104: op1_02_inv09 = 1;
    105: op1_02_inv09 = 1;
    107: op1_02_inv09 = 1;
    109: op1_02_inv09 = 1;
    112: op1_02_inv09 = 1;
    113: op1_02_inv09 = 1;
    114: op1_02_inv09 = 1;
    29: op1_02_inv09 = 1;
    117: op1_02_inv09 = 1;
    119: op1_02_inv09 = 1;
    121: op1_02_inv09 = 1;
    123: op1_02_inv09 = 1;
    124: op1_02_inv09 = 1;
    125: op1_02_inv09 = 1;
    128: op1_02_inv09 = 1;
    129: op1_02_inv09 = 1;
    default: op1_02_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の10番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in10 = reg_0832;
    53: op1_02_in10 = reg_0116;
    72: op1_02_in10 = reg_0405;
    49: op1_02_in10 = reg_0415;
    55: op1_02_in10 = reg_0936;
    73: op1_02_in10 = reg_0646;
    69: op1_02_in10 = reg_0755;
    86: op1_02_in10 = reg_0719;
    59: op1_02_in10 = reg_0431;
    71: op1_02_in10 = imem00_in[3:0];
    61: op1_02_in10 = reg_1034;
    50: op1_02_in10 = reg_0886;
    68: op1_02_in10 = reg_0798;
    60: op1_02_in10 = reg_0798;
    122: op1_02_in10 = reg_0798;
    48: op1_02_in10 = reg_0090;
    74: op1_02_in10 = reg_0575;
    46: op1_02_in10 = reg_0066;
    47: op1_02_in10 = reg_0287;
    75: op1_02_in10 = reg_0588;
    56: op1_02_in10 = reg_0169;
    87: op1_02_in10 = reg_0191;
    37: op1_02_in10 = reg_0087;
    51: op1_02_in10 = reg_0087;
    33: op1_02_in10 = reg_0121;
    76: op1_02_in10 = reg_0346;
    57: op1_02_in10 = reg_0606;
    70: op1_02_in10 = reg_1392;
    77: op1_02_in10 = reg_0046;
    44: op1_02_in10 = reg_0566;
    106: op1_02_in10 = reg_0566;
    58: op1_02_in10 = reg_0235;
    88: op1_02_in10 = reg_0480;
    78: op1_02_in10 = reg_0435;
    34: op1_02_in10 = reg_0002;
    79: op1_02_in10 = reg_0848;
    42: op1_02_in10 = imem00_in[15:12];
    80: op1_02_in10 = imem07_in[7:4];
    62: op1_02_in10 = reg_1254;
    81: op1_02_in10 = reg_0432;
    89: op1_02_in10 = reg_1282;
    63: op1_02_in10 = reg_1206;
    82: op1_02_in10 = reg_1198;
    83: op1_02_in10 = reg_0206;
    64: op1_02_in10 = reg_0904;
    84: op1_02_in10 = reg_0972;
    65: op1_02_in10 = reg_0774;
    85: op1_02_in10 = reg_0152;
    90: op1_02_in10 = reg_1301;
    66: op1_02_in10 = reg_0877;
    91: op1_02_in10 = reg_0860;
    67: op1_02_in10 = reg_0363;
    92: op1_02_in10 = reg_1458;
    93: op1_02_in10 = reg_0269;
    94: op1_02_in10 = reg_1488;
    95: op1_02_in10 = reg_0041;
    96: op1_02_in10 = reg_1348;
    97: op1_02_in10 = reg_0392;
    98: op1_02_in10 = reg_0256;
    99: op1_02_in10 = reg_0058;
    100: op1_02_in10 = reg_0350;
    101: op1_02_in10 = reg_0934;
    102: op1_02_in10 = reg_0028;
    103: op1_02_in10 = reg_0351;
    107: op1_02_in10 = reg_0351;
    104: op1_02_in10 = reg_0254;
    105: op1_02_in10 = reg_0649;
    108: op1_02_in10 = reg_0155;
    109: op1_02_in10 = reg_1056;
    110: op1_02_in10 = reg_0349;
    111: op1_02_in10 = reg_0353;
    112: op1_02_in10 = reg_0342;
    113: op1_02_in10 = reg_0188;
    114: op1_02_in10 = reg_0716;
    115: op1_02_in10 = reg_1074;
    116: op1_02_in10 = reg_0731;
    117: op1_02_in10 = reg_0776;
    118: op1_02_in10 = reg_0776;
    119: op1_02_in10 = reg_0897;
    120: op1_02_in10 = reg_0799;
    121: op1_02_in10 = reg_0922;
    123: op1_02_in10 = reg_0521;
    124: op1_02_in10 = reg_0736;
    125: op1_02_in10 = reg_1098;
    126: op1_02_in10 = imem06_in[7:4];
    127: op1_02_in10 = reg_0279;
    43: op1_02_in10 = reg_0250;
    128: op1_02_in10 = reg_0236;
    129: op1_02_in10 = reg_0883;
    130: op1_02_in10 = reg_0876;
    131: op1_02_in10 = reg_1459;
    default: op1_02_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_02_inv10 = 1;
    69: op1_02_inv10 = 1;
    86: op1_02_inv10 = 1;
    71: op1_02_inv10 = 1;
    68: op1_02_inv10 = 1;
    74: op1_02_inv10 = 1;
    46: op1_02_inv10 = 1;
    47: op1_02_inv10 = 1;
    75: op1_02_inv10 = 1;
    60: op1_02_inv10 = 1;
    76: op1_02_inv10 = 1;
    70: op1_02_inv10 = 1;
    77: op1_02_inv10 = 1;
    58: op1_02_inv10 = 1;
    88: op1_02_inv10 = 1;
    78: op1_02_inv10 = 1;
    51: op1_02_inv10 = 1;
    79: op1_02_inv10 = 1;
    81: op1_02_inv10 = 1;
    89: op1_02_inv10 = 1;
    63: op1_02_inv10 = 1;
    83: op1_02_inv10 = 1;
    64: op1_02_inv10 = 1;
    84: op1_02_inv10 = 1;
    85: op1_02_inv10 = 1;
    90: op1_02_inv10 = 1;
    94: op1_02_inv10 = 1;
    95: op1_02_inv10 = 1;
    96: op1_02_inv10 = 1;
    97: op1_02_inv10 = 1;
    99: op1_02_inv10 = 1;
    101: op1_02_inv10 = 1;
    102: op1_02_inv10 = 1;
    103: op1_02_inv10 = 1;
    104: op1_02_inv10 = 1;
    106: op1_02_inv10 = 1;
    107: op1_02_inv10 = 1;
    108: op1_02_inv10 = 1;
    114: op1_02_inv10 = 1;
    115: op1_02_inv10 = 1;
    116: op1_02_inv10 = 1;
    117: op1_02_inv10 = 1;
    118: op1_02_inv10 = 1;
    124: op1_02_inv10 = 1;
    125: op1_02_inv10 = 1;
    129: op1_02_inv10 = 1;
    131: op1_02_inv10 = 1;
    default: op1_02_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の11番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in11 = reg_0649;
    73: op1_02_in11 = reg_0649;
    53: op1_02_in11 = reg_0622;
    72: op1_02_in11 = reg_0122;
    49: op1_02_in11 = reg_0103;
    55: op1_02_in11 = reg_0320;
    69: op1_02_in11 = reg_0191;
    86: op1_02_in11 = reg_0338;
    59: op1_02_in11 = reg_0389;
    71: op1_02_in11 = imem00_in[11:8];
    61: op1_02_in11 = reg_0634;
    50: op1_02_in11 = reg_0641;
    42: op1_02_in11 = reg_0641;
    68: op1_02_in11 = reg_0451;
    48: op1_02_in11 = reg_0197;
    74: op1_02_in11 = reg_0864;
    46: op1_02_in11 = reg_0182;
    47: op1_02_in11 = reg_0366;
    75: op1_02_in11 = reg_0495;
    56: op1_02_in11 = reg_0413;
    87: op1_02_in11 = reg_0840;
    33: op1_02_in11 = reg_0440;
    60: op1_02_in11 = reg_0341;
    64: op1_02_in11 = reg_0341;
    76: op1_02_in11 = reg_0045;
    57: op1_02_in11 = reg_0587;
    70: op1_02_in11 = reg_0069;
    77: op1_02_in11 = reg_0215;
    85: op1_02_in11 = reg_0215;
    44: op1_02_in11 = reg_0333;
    58: op1_02_in11 = reg_1145;
    88: op1_02_in11 = reg_0481;
    78: op1_02_in11 = reg_0203;
    51: op1_02_in11 = reg_0520;
    123: op1_02_in11 = reg_0520;
    34: op1_02_in11 = reg_0087;
    79: op1_02_in11 = reg_1515;
    80: op1_02_in11 = imem07_in[11:8];
    62: op1_02_in11 = reg_1033;
    81: op1_02_in11 = reg_0970;
    89: op1_02_in11 = reg_0790;
    63: op1_02_in11 = reg_0959;
    82: op1_02_in11 = reg_0681;
    83: op1_02_in11 = reg_0038;
    84: op1_02_in11 = reg_0126;
    65: op1_02_in11 = reg_0030;
    90: op1_02_in11 = reg_0178;
    66: op1_02_in11 = reg_0839;
    91: op1_02_in11 = reg_0172;
    67: op1_02_in11 = reg_0047;
    92: op1_02_in11 = reg_0111;
    93: op1_02_in11 = reg_0271;
    94: op1_02_in11 = reg_0470;
    95: op1_02_in11 = reg_0011;
    96: op1_02_in11 = reg_0799;
    97: op1_02_in11 = reg_0630;
    98: op1_02_in11 = reg_0472;
    99: op1_02_in11 = reg_0057;
    100: op1_02_in11 = reg_0427;
    101: op1_02_in11 = reg_0055;
    102: op1_02_in11 = reg_0228;
    103: op1_02_in11 = reg_0352;
    107: op1_02_in11 = reg_0352;
    104: op1_02_in11 = reg_0455;
    105: op1_02_in11 = reg_0174;
    106: op1_02_in11 = reg_0940;
    108: op1_02_in11 = reg_1418;
    109: op1_02_in11 = reg_0703;
    110: op1_02_in11 = reg_0597;
    111: op1_02_in11 = reg_0351;
    112: op1_02_in11 = reg_0061;
    113: op1_02_in11 = reg_0189;
    114: op1_02_in11 = reg_0718;
    115: op1_02_in11 = reg_0900;
    116: op1_02_in11 = reg_0797;
    117: op1_02_in11 = reg_1451;
    118: op1_02_in11 = reg_0778;
    119: op1_02_in11 = reg_0800;
    125: op1_02_in11 = reg_0800;
    120: op1_02_in11 = reg_0151;
    121: op1_02_in11 = reg_1440;
    122: op1_02_in11 = reg_1474;
    124: op1_02_in11 = reg_0888;
    126: op1_02_in11 = reg_0397;
    127: op1_02_in11 = imem03_in[11:8];
    43: op1_02_in11 = reg_0523;
    128: op1_02_in11 = reg_0731;
    129: op1_02_in11 = reg_0722;
    130: op1_02_in11 = reg_0745;
    131: op1_02_in11 = reg_1230;
    default: op1_02_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv11 = 1;
    53: op1_02_inv11 = 1;
    49: op1_02_inv11 = 1;
    73: op1_02_inv11 = 1;
    69: op1_02_inv11 = 1;
    61: op1_02_inv11 = 1;
    50: op1_02_inv11 = 1;
    74: op1_02_inv11 = 1;
    60: op1_02_inv11 = 1;
    57: op1_02_inv11 = 1;
    70: op1_02_inv11 = 1;
    77: op1_02_inv11 = 1;
    44: op1_02_inv11 = 1;
    88: op1_02_inv11 = 1;
    34: op1_02_inv11 = 1;
    79: op1_02_inv11 = 1;
    81: op1_02_inv11 = 1;
    89: op1_02_inv11 = 1;
    64: op1_02_inv11 = 1;
    90: op1_02_inv11 = 1;
    66: op1_02_inv11 = 1;
    91: op1_02_inv11 = 1;
    67: op1_02_inv11 = 1;
    95: op1_02_inv11 = 1;
    96: op1_02_inv11 = 1;
    97: op1_02_inv11 = 1;
    98: op1_02_inv11 = 1;
    99: op1_02_inv11 = 1;
    102: op1_02_inv11 = 1;
    104: op1_02_inv11 = 1;
    105: op1_02_inv11 = 1;
    106: op1_02_inv11 = 1;
    113: op1_02_inv11 = 1;
    116: op1_02_inv11 = 1;
    117: op1_02_inv11 = 1;
    120: op1_02_inv11 = 1;
    122: op1_02_inv11 = 1;
    124: op1_02_inv11 = 1;
    125: op1_02_inv11 = 1;
    126: op1_02_inv11 = 1;
    127: op1_02_inv11 = 1;
    43: op1_02_inv11 = 1;
    128: op1_02_inv11 = 1;
    130: op1_02_inv11 = 1;
    default: op1_02_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の12番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in12 = reg_0066;
    53: op1_02_in12 = reg_0067;
    72: op1_02_in12 = reg_0175;
    49: op1_02_in12 = reg_0100;
    55: op1_02_in12 = reg_0340;
    73: op1_02_in12 = reg_1403;
    69: op1_02_in12 = reg_0154;
    86: op1_02_in12 = reg_0339;
    59: op1_02_in12 = reg_0089;
    99: op1_02_in12 = reg_0089;
    71: op1_02_in12 = imem00_in[15:12];
    61: op1_02_in12 = reg_0601;
    50: op1_02_in12 = reg_0638;
    68: op1_02_in12 = reg_0262;
    48: op1_02_in12 = reg_0272;
    74: op1_02_in12 = reg_0037;
    46: op1_02_in12 = imem05_in[11:8];
    47: op1_02_in12 = reg_0738;
    75: op1_02_in12 = reg_1207;
    56: op1_02_in12 = reg_0623;
    87: op1_02_in12 = reg_0710;
    33: op1_02_in12 = imem01_in[3:0];
    60: op1_02_in12 = reg_0096;
    76: op1_02_in12 = reg_0418;
    57: op1_02_in12 = reg_0563;
    70: op1_02_in12 = reg_0802;
    77: op1_02_in12 = reg_0213;
    44: op1_02_in12 = reg_0541;
    58: op1_02_in12 = reg_0177;
    88: op1_02_in12 = reg_0479;
    78: op1_02_in12 = reg_0073;
    51: op1_02_in12 = reg_0123;
    79: op1_02_in12 = reg_0313;
    42: op1_02_in12 = reg_0640;
    80: op1_02_in12 = reg_1441;
    62: op1_02_in12 = reg_0547;
    81: op1_02_in12 = reg_0379;
    89: op1_02_in12 = reg_0425;
    63: op1_02_in12 = reg_0881;
    82: op1_02_in12 = reg_0414;
    116: op1_02_in12 = reg_0414;
    83: op1_02_in12 = imem06_in[7:4];
    64: op1_02_in12 = reg_0596;
    84: op1_02_in12 = reg_0876;
    65: op1_02_in12 = reg_0366;
    85: op1_02_in12 = reg_0018;
    90: op1_02_in12 = reg_0104;
    66: op1_02_in12 = reg_0695;
    91: op1_02_in12 = reg_0109;
    67: op1_02_in12 = reg_0093;
    92: op1_02_in12 = reg_0631;
    93: op1_02_in12 = reg_0023;
    94: op1_02_in12 = imem05_in[3:0];
    95: op1_02_in12 = imem02_in[7:4];
    96: op1_02_in12 = reg_0038;
    97: op1_02_in12 = reg_0794;
    98: op1_02_in12 = reg_0382;
    100: op1_02_in12 = imem04_in[7:4];
    101: op1_02_in12 = reg_0532;
    102: op1_02_in12 = reg_0085;
    103: op1_02_in12 = reg_0059;
    104: op1_02_in12 = reg_0497;
    105: op1_02_in12 = reg_0562;
    106: op1_02_in12 = reg_1169;
    107: op1_02_in12 = reg_0431;
    108: op1_02_in12 = reg_1406;
    109: op1_02_in12 = reg_0170;
    110: op1_02_in12 = reg_1093;
    111: op1_02_in12 = reg_0352;
    112: op1_02_in12 = reg_1419;
    113: op1_02_in12 = reg_0134;
    114: op1_02_in12 = reg_1303;
    115: op1_02_in12 = reg_0429;
    117: op1_02_in12 = reg_0628;
    118: op1_02_in12 = reg_0972;
    119: op1_02_in12 = reg_0903;
    120: op1_02_in12 = reg_0206;
    121: op1_02_in12 = reg_1349;
    122: op1_02_in12 = reg_0967;
    124: op1_02_in12 = reg_0492;
    125: op1_02_in12 = reg_1006;
    126: op1_02_in12 = reg_0925;
    127: op1_02_in12 = reg_0185;
    43: op1_02_in12 = reg_0445;
    128: op1_02_in12 = reg_0797;
    129: op1_02_in12 = reg_0201;
    130: op1_02_in12 = reg_1492;
    131: op1_02_in12 = reg_0821;
    default: op1_02_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_02_inv12 = 1;
    72: op1_02_inv12 = 1;
    49: op1_02_inv12 = 1;
    55: op1_02_inv12 = 1;
    86: op1_02_inv12 = 1;
    71: op1_02_inv12 = 1;
    50: op1_02_inv12 = 1;
    68: op1_02_inv12 = 1;
    48: op1_02_inv12 = 1;
    74: op1_02_inv12 = 1;
    47: op1_02_inv12 = 1;
    75: op1_02_inv12 = 1;
    33: op1_02_inv12 = 1;
    57: op1_02_inv12 = 1;
    77: op1_02_inv12 = 1;
    88: op1_02_inv12 = 1;
    78: op1_02_inv12 = 1;
    51: op1_02_inv12 = 1;
    80: op1_02_inv12 = 1;
    89: op1_02_inv12 = 1;
    63: op1_02_inv12 = 1;
    82: op1_02_inv12 = 1;
    83: op1_02_inv12 = 1;
    90: op1_02_inv12 = 1;
    66: op1_02_inv12 = 1;
    93: op1_02_inv12 = 1;
    95: op1_02_inv12 = 1;
    98: op1_02_inv12 = 1;
    99: op1_02_inv12 = 1;
    101: op1_02_inv12 = 1;
    104: op1_02_inv12 = 1;
    105: op1_02_inv12 = 1;
    106: op1_02_inv12 = 1;
    110: op1_02_inv12 = 1;
    111: op1_02_inv12 = 1;
    119: op1_02_inv12 = 1;
    120: op1_02_inv12 = 1;
    124: op1_02_inv12 = 1;
    126: op1_02_inv12 = 1;
    127: op1_02_inv12 = 1;
    43: op1_02_inv12 = 1;
    128: op1_02_inv12 = 1;
    129: op1_02_inv12 = 1;
    130: op1_02_inv12 = 1;
    131: op1_02_inv12 = 1;
    default: op1_02_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の13番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in13 = reg_0316;
    53: op1_02_in13 = reg_0214;
    72: op1_02_in13 = reg_0372;
    49: op1_02_in13 = reg_0050;
    55: op1_02_in13 = reg_0096;
    73: op1_02_in13 = reg_0938;
    69: op1_02_in13 = reg_0709;
    86: op1_02_in13 = reg_1488;
    59: op1_02_in13 = reg_0005;
    71: op1_02_in13 = reg_0293;
    61: op1_02_in13 = reg_0549;
    50: op1_02_in13 = reg_0201;
    68: op1_02_in13 = reg_0097;
    48: op1_02_in13 = reg_0205;
    74: op1_02_in13 = reg_1035;
    46: op1_02_in13 = reg_0539;
    44: op1_02_in13 = reg_0539;
    47: op1_02_in13 = reg_0519;
    75: op1_02_in13 = reg_0494;
    56: op1_02_in13 = reg_0620;
    87: op1_02_in13 = reg_1449;
    33: op1_02_in13 = imem01_in[7:4];
    60: op1_02_in13 = reg_0164;
    76: op1_02_in13 = reg_0300;
    57: op1_02_in13 = reg_0561;
    70: op1_02_in13 = reg_0281;
    77: op1_02_in13 = imem07_in[7:4];
    58: op1_02_in13 = reg_1003;
    88: op1_02_in13 = reg_0478;
    78: op1_02_in13 = reg_1068;
    79: op1_02_in13 = reg_0999;
    42: op1_02_in13 = reg_0431;
    129: op1_02_in13 = reg_0431;
    80: op1_02_in13 = reg_1440;
    62: op1_02_in13 = reg_0242;
    81: op1_02_in13 = reg_0897;
    89: op1_02_in13 = imem04_in[15:12];
    63: op1_02_in13 = reg_0188;
    111: op1_02_in13 = reg_0188;
    82: op1_02_in13 = reg_0232;
    83: op1_02_in13 = reg_1426;
    64: op1_02_in13 = reg_0199;
    84: op1_02_in13 = reg_0381;
    65: op1_02_in13 = reg_0740;
    85: op1_02_in13 = imem07_in[11:8];
    90: op1_02_in13 = reg_0885;
    66: op1_02_in13 = reg_0632;
    91: op1_02_in13 = reg_0398;
    67: op1_02_in13 = imem01_in[3:0];
    92: op1_02_in13 = reg_0380;
    93: op1_02_in13 = reg_0152;
    94: op1_02_in13 = reg_0204;
    95: op1_02_in13 = reg_0475;
    96: op1_02_in13 = imem06_in[3:0];
    97: op1_02_in13 = reg_0196;
    98: op1_02_in13 = reg_0496;
    99: op1_02_in13 = reg_0027;
    100: op1_02_in13 = reg_0129;
    101: op1_02_in13 = reg_1074;
    102: op1_02_in13 = reg_0084;
    103: op1_02_in13 = reg_1324;
    104: op1_02_in13 = reg_0973;
    105: op1_02_in13 = reg_0391;
    106: op1_02_in13 = reg_0477;
    107: op1_02_in13 = reg_0388;
    108: op1_02_in13 = reg_0821;
    109: op1_02_in13 = reg_0309;
    110: op1_02_in13 = reg_1199;
    112: op1_02_in13 = reg_0698;
    113: op1_02_in13 = reg_0059;
    114: op1_02_in13 = reg_0636;
    115: op1_02_in13 = reg_0776;
    116: op1_02_in13 = reg_0412;
    117: op1_02_in13 = reg_0876;
    118: op1_02_in13 = reg_1451;
    119: op1_02_in13 = reg_0006;
    120: op1_02_in13 = imem06_in[11:8];
    121: op1_02_in13 = reg_0157;
    122: op1_02_in13 = reg_0968;
    124: op1_02_in13 = reg_0240;
    125: op1_02_in13 = reg_0227;
    126: op1_02_in13 = reg_0870;
    127: op1_02_in13 = reg_0154;
    43: op1_02_in13 = reg_0649;
    128: op1_02_in13 = reg_0531;
    130: op1_02_in13 = reg_1098;
    131: op1_02_in13 = reg_0476;
    default: op1_02_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv13 = 1;
    53: op1_02_inv13 = 1;
    72: op1_02_inv13 = 1;
    55: op1_02_inv13 = 1;
    69: op1_02_inv13 = 1;
    71: op1_02_inv13 = 1;
    50: op1_02_inv13 = 1;
    74: op1_02_inv13 = 1;
    47: op1_02_inv13 = 1;
    56: op1_02_inv13 = 1;
    60: op1_02_inv13 = 1;
    57: op1_02_inv13 = 1;
    70: op1_02_inv13 = 1;
    77: op1_02_inv13 = 1;
    44: op1_02_inv13 = 1;
    58: op1_02_inv13 = 1;
    88: op1_02_inv13 = 1;
    42: op1_02_inv13 = 1;
    80: op1_02_inv13 = 1;
    64: op1_02_inv13 = 1;
    85: op1_02_inv13 = 1;
    91: op1_02_inv13 = 1;
    92: op1_02_inv13 = 1;
    94: op1_02_inv13 = 1;
    95: op1_02_inv13 = 1;
    96: op1_02_inv13 = 1;
    97: op1_02_inv13 = 1;
    98: op1_02_inv13 = 1;
    102: op1_02_inv13 = 1;
    103: op1_02_inv13 = 1;
    104: op1_02_inv13 = 1;
    105: op1_02_inv13 = 1;
    107: op1_02_inv13 = 1;
    110: op1_02_inv13 = 1;
    112: op1_02_inv13 = 1;
    118: op1_02_inv13 = 1;
    121: op1_02_inv13 = 1;
    122: op1_02_inv13 = 1;
    126: op1_02_inv13 = 1;
    127: op1_02_inv13 = 1;
    43: op1_02_inv13 = 1;
    128: op1_02_inv13 = 1;
    default: op1_02_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の14番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in14 = reg_0317;
    53: op1_02_in14 = imem07_in[11:8];
    72: op1_02_in14 = reg_0728;
    49: op1_02_in14 = reg_0003;
    55: op1_02_in14 = reg_0095;
    73: op1_02_in14 = reg_0196;
    69: op1_02_in14 = reg_0704;
    79: op1_02_in14 = reg_0704;
    86: op1_02_in14 = reg_0035;
    59: op1_02_in14 = reg_0786;
    71: op1_02_in14 = reg_1027;
    61: op1_02_in14 = reg_0610;
    50: op1_02_in14 = reg_0410;
    68: op1_02_in14 = reg_0065;
    48: op1_02_in14 = reg_0207;
    74: op1_02_in14 = reg_1468;
    46: op1_02_in14 = reg_0183;
    47: op1_02_in14 = reg_0484;
    75: op1_02_in14 = reg_1450;
    56: op1_02_in14 = reg_0591;
    87: op1_02_in14 = reg_1063;
    127: op1_02_in14 = reg_1063;
    33: op1_02_in14 = reg_0335;
    60: op1_02_in14 = reg_0209;
    76: op1_02_in14 = reg_0873;
    57: op1_02_in14 = reg_1140;
    70: op1_02_in14 = reg_0311;
    77: op1_02_in14 = reg_0490;
    85: op1_02_in14 = reg_0490;
    44: op1_02_in14 = reg_0491;
    58: op1_02_in14 = reg_0448;
    88: op1_02_in14 = reg_0218;
    78: op1_02_in14 = imem01_in[3:0];
    113: op1_02_in14 = imem01_in[3:0];
    42: op1_02_in14 = reg_0409;
    80: op1_02_in14 = reg_0225;
    62: op1_02_in14 = reg_0239;
    81: op1_02_in14 = reg_0531;
    89: op1_02_in14 = reg_0263;
    63: op1_02_in14 = reg_0387;
    82: op1_02_in14 = reg_0487;
    83: op1_02_in14 = reg_0870;
    64: op1_02_in14 = reg_0304;
    84: op1_02_in14 = reg_0712;
    65: op1_02_in14 = reg_0623;
    90: op1_02_in14 = reg_0880;
    66: op1_02_in14 = reg_0068;
    91: op1_02_in14 = reg_0141;
    67: op1_02_in14 = reg_0078;
    92: op1_02_in14 = reg_0560;
    117: op1_02_in14 = reg_0560;
    93: op1_02_in14 = reg_0212;
    94: op1_02_in14 = reg_0832;
    95: op1_02_in14 = reg_0455;
    96: op1_02_in14 = reg_0195;
    97: op1_02_in14 = reg_0603;
    98: op1_02_in14 = reg_0380;
    99: op1_02_in14 = reg_0267;
    100: op1_02_in14 = reg_0467;
    101: op1_02_in14 = reg_0436;
    102: op1_02_in14 = reg_0520;
    103: op1_02_in14 = imem01_in[11:8];
    104: op1_02_in14 = reg_0128;
    105: op1_02_in14 = reg_1104;
    106: op1_02_in14 = reg_0301;
    107: op1_02_in14 = reg_0060;
    108: op1_02_in14 = reg_0352;
    109: op1_02_in14 = reg_0924;
    110: op1_02_in14 = reg_0885;
    111: op1_02_in14 = reg_0722;
    112: op1_02_in14 = reg_0582;
    114: op1_02_in14 = reg_0619;
    115: op1_02_in14 = reg_0326;
    116: op1_02_in14 = reg_1041;
    118: op1_02_in14 = reg_0105;
    119: op1_02_in14 = imem03_in[11:8];
    120: op1_02_in14 = reg_1334;
    121: op1_02_in14 = reg_0777;
    122: op1_02_in14 = reg_0439;
    124: op1_02_in14 = reg_1348;
    125: op1_02_in14 = reg_0006;
    126: op1_02_in14 = reg_0696;
    43: op1_02_in14 = reg_0650;
    128: op1_02_in14 = reg_1200;
    129: op1_02_in14 = reg_0435;
    130: op1_02_in14 = reg_0848;
    131: op1_02_in14 = reg_0927;
    default: op1_02_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_02_inv14 = 1;
    49: op1_02_inv14 = 1;
    86: op1_02_inv14 = 1;
    59: op1_02_inv14 = 1;
    71: op1_02_inv14 = 1;
    50: op1_02_inv14 = 1;
    48: op1_02_inv14 = 1;
    74: op1_02_inv14 = 1;
    46: op1_02_inv14 = 1;
    75: op1_02_inv14 = 1;
    70: op1_02_inv14 = 1;
    77: op1_02_inv14 = 1;
    44: op1_02_inv14 = 1;
    42: op1_02_inv14 = 1;
    62: op1_02_inv14 = 1;
    83: op1_02_inv14 = 1;
    67: op1_02_inv14 = 1;
    92: op1_02_inv14 = 1;
    93: op1_02_inv14 = 1;
    94: op1_02_inv14 = 1;
    96: op1_02_inv14 = 1;
    100: op1_02_inv14 = 1;
    101: op1_02_inv14 = 1;
    102: op1_02_inv14 = 1;
    105: op1_02_inv14 = 1;
    107: op1_02_inv14 = 1;
    108: op1_02_inv14 = 1;
    109: op1_02_inv14 = 1;
    114: op1_02_inv14 = 1;
    115: op1_02_inv14 = 1;
    116: op1_02_inv14 = 1;
    117: op1_02_inv14 = 1;
    119: op1_02_inv14 = 1;
    120: op1_02_inv14 = 1;
    124: op1_02_inv14 = 1;
    125: op1_02_inv14 = 1;
    127: op1_02_inv14 = 1;
    128: op1_02_inv14 = 1;
    129: op1_02_inv14 = 1;
    default: op1_02_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の15番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in15 = reg_0167;
    53: op1_02_in15 = reg_0490;
    72: op1_02_in15 = reg_0093;
    49: op1_02_in15 = reg_0086;
    55: op1_02_in15 = reg_0211;
    73: op1_02_in15 = reg_0797;
    69: op1_02_in15 = reg_1149;
    86: op1_02_in15 = reg_0736;
    59: op1_02_in15 = reg_1253;
    71: op1_02_in15 = reg_0221;
    61: op1_02_in15 = reg_0787;
    50: op1_02_in15 = reg_0405;
    68: op1_02_in15 = reg_0150;
    48: op1_02_in15 = reg_0037;
    74: op1_02_in15 = reg_0720;
    46: op1_02_in15 = reg_0090;
    75: op1_02_in15 = reg_0629;
    56: op1_02_in15 = reg_0321;
    87: op1_02_in15 = reg_0962;
    33: op1_02_in15 = reg_0549;
    60: op1_02_in15 = reg_0016;
    76: op1_02_in15 = reg_1484;
    57: op1_02_in15 = imem02_in[7:4];
    70: op1_02_in15 = reg_0312;
    77: op1_02_in15 = reg_0461;
    44: op1_02_in15 = reg_0303;
    58: op1_02_in15 = reg_0107;
    88: op1_02_in15 = reg_0348;
    78: op1_02_in15 = reg_0331;
    79: op1_02_in15 = reg_0177;
    42: op1_02_in15 = reg_0072;
    80: op1_02_in15 = reg_0921;
    62: op1_02_in15 = reg_0609;
    81: op1_02_in15 = imem02_in[11:8];
    89: op1_02_in15 = reg_1372;
    100: op1_02_in15 = reg_1372;
    63: op1_02_in15 = reg_0027;
    82: op1_02_in15 = reg_0835;
    83: op1_02_in15 = reg_0860;
    64: op1_02_in15 = reg_0837;
    84: op1_02_in15 = reg_0307;
    65: op1_02_in15 = reg_0593;
    85: op1_02_in15 = reg_1439;
    90: op1_02_in15 = imem03_in[15:12];
    66: op1_02_in15 = reg_0313;
    91: op1_02_in15 = reg_0619;
    67: op1_02_in15 = reg_0290;
    92: op1_02_in15 = reg_1492;
    93: op1_02_in15 = reg_0214;
    94: op1_02_in15 = reg_0333;
    95: op1_02_in15 = reg_0934;
    96: op1_02_in15 = reg_1468;
    97: op1_02_in15 = reg_0449;
    98: op1_02_in15 = reg_0473;
    99: op1_02_in15 = imem01_in[7:4];
    101: op1_02_in15 = reg_0776;
    102: op1_02_in15 = reg_0483;
    103: op1_02_in15 = reg_0576;
    104: op1_02_in15 = reg_0127;
    105: op1_02_in15 = reg_0182;
    106: op1_02_in15 = reg_0794;
    107: op1_02_in15 = imem01_in[15:12];
    108: op1_02_in15 = reg_0416;
    109: op1_02_in15 = reg_0465;
    110: op1_02_in15 = reg_0882;
    111: op1_02_in15 = reg_0428;
    112: op1_02_in15 = reg_0268;
    113: op1_02_in15 = reg_1034;
    114: op1_02_in15 = reg_0568;
    115: op1_02_in15 = reg_0628;
    116: op1_02_in15 = reg_0199;
    117: op1_02_in15 = reg_0695;
    118: op1_02_in15 = reg_0684;
    119: op1_02_in15 = reg_1145;
    120: op1_02_in15 = reg_0870;
    121: op1_02_in15 = reg_0775;
    122: op1_02_in15 = reg_0438;
    124: op1_02_in15 = reg_1346;
    125: op1_02_in15 = imem03_in[11:8];
    126: op1_02_in15 = reg_0984;
    127: op1_02_in15 = reg_1425;
    43: op1_02_in15 = reg_0567;
    128: op1_02_in15 = reg_0796;
    129: op1_02_in15 = reg_0058;
    130: op1_02_in15 = reg_1006;
    131: op1_02_in15 = reg_0886;
    default: op1_02_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_02_inv15 = 1;
    49: op1_02_inv15 = 1;
    55: op1_02_inv15 = 1;
    73: op1_02_inv15 = 1;
    69: op1_02_inv15 = 1;
    71: op1_02_inv15 = 1;
    68: op1_02_inv15 = 1;
    56: op1_02_inv15 = 1;
    76: op1_02_inv15 = 1;
    70: op1_02_inv15 = 1;
    44: op1_02_inv15 = 1;
    88: op1_02_inv15 = 1;
    62: op1_02_inv15 = 1;
    81: op1_02_inv15 = 1;
    89: op1_02_inv15 = 1;
    64: op1_02_inv15 = 1;
    84: op1_02_inv15 = 1;
    65: op1_02_inv15 = 1;
    90: op1_02_inv15 = 1;
    91: op1_02_inv15 = 1;
    67: op1_02_inv15 = 1;
    92: op1_02_inv15 = 1;
    93: op1_02_inv15 = 1;
    94: op1_02_inv15 = 1;
    96: op1_02_inv15 = 1;
    97: op1_02_inv15 = 1;
    99: op1_02_inv15 = 1;
    100: op1_02_inv15 = 1;
    101: op1_02_inv15 = 1;
    102: op1_02_inv15 = 1;
    103: op1_02_inv15 = 1;
    105: op1_02_inv15 = 1;
    106: op1_02_inv15 = 1;
    107: op1_02_inv15 = 1;
    109: op1_02_inv15 = 1;
    110: op1_02_inv15 = 1;
    111: op1_02_inv15 = 1;
    112: op1_02_inv15 = 1;
    113: op1_02_inv15 = 1;
    115: op1_02_inv15 = 1;
    116: op1_02_inv15 = 1;
    120: op1_02_inv15 = 1;
    121: op1_02_inv15 = 1;
    122: op1_02_inv15 = 1;
    124: op1_02_inv15 = 1;
    129: op1_02_inv15 = 1;
    130: op1_02_inv15 = 1;
    131: op1_02_inv15 = 1;
    default: op1_02_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の16番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in16 = reg_0070;
    53: op1_02_in16 = reg_1094;
    72: op1_02_in16 = reg_0258;
    49: op1_02_in16 = reg_0521;
    55: op1_02_in16 = reg_0209;
    73: op1_02_in16 = reg_0151;
    124: op1_02_in16 = reg_0151;
    69: op1_02_in16 = imem03_in[3:0];
    86: op1_02_in16 = reg_0251;
    59: op1_02_in16 = imem01_in[15:12];
    71: op1_02_in16 = reg_1229;
    61: op1_02_in16 = reg_0259;
    50: op1_02_in16 = reg_0353;
    68: op1_02_in16 = reg_0063;
    48: op1_02_in16 = reg_0014;
    74: op1_02_in16 = imem06_in[7:4];
    46: op1_02_in16 = reg_0196;
    75: op1_02_in16 = reg_0390;
    56: op1_02_in16 = reg_0085;
    87: op1_02_in16 = reg_1184;
    33: op1_02_in16 = reg_0548;
    60: op1_02_in16 = reg_0033;
    76: op1_02_in16 = reg_0275;
    57: op1_02_in16 = reg_0494;
    70: op1_02_in16 = reg_0758;
    77: op1_02_in16 = reg_1415;
    44: op1_02_in16 = reg_0090;
    58: op1_02_in16 = reg_0113;
    88: op1_02_in16 = reg_0425;
    78: op1_02_in16 = reg_0743;
    79: op1_02_in16 = reg_1425;
    42: op1_02_in16 = reg_0060;
    80: op1_02_in16 = reg_0924;
    62: op1_02_in16 = reg_1151;
    81: op1_02_in16 = reg_0217;
    89: op1_02_in16 = reg_1368;
    63: op1_02_in16 = reg_0822;
    82: op1_02_in16 = reg_0337;
    83: op1_02_in16 = reg_0869;
    64: op1_02_in16 = reg_0836;
    84: op1_02_in16 = reg_0008;
    92: op1_02_in16 = reg_0008;
    65: op1_02_in16 = reg_0103;
    85: op1_02_in16 = reg_0892;
    90: op1_02_in16 = reg_0348;
    110: op1_02_in16 = reg_0348;
    66: op1_02_in16 = reg_0525;
    91: op1_02_in16 = reg_0617;
    67: op1_02_in16 = reg_0291;
    93: op1_02_in16 = reg_0213;
    94: op1_02_in16 = reg_0184;
    95: op1_02_in16 = reg_0532;
    96: op1_02_in16 = reg_0795;
    97: op1_02_in16 = imem06_in[3:0];
    98: op1_02_in16 = reg_1492;
    99: op1_02_in16 = reg_1152;
    100: op1_02_in16 = reg_1369;
    101: op1_02_in16 = reg_0778;
    103: op1_02_in16 = reg_0401;
    104: op1_02_in16 = reg_1140;
    105: op1_02_in16 = reg_0564;
    106: op1_02_in16 = reg_1373;
    107: op1_02_in16 = reg_0183;
    108: op1_02_in16 = reg_0387;
    109: op1_02_in16 = reg_0284;
    111: op1_02_in16 = reg_0431;
    112: op1_02_in16 = reg_0256;
    113: op1_02_in16 = reg_0930;
    114: op1_02_in16 = reg_0570;
    115: op1_02_in16 = reg_0878;
    116: op1_02_in16 = reg_1077;
    117: op1_02_in16 = reg_0800;
    118: op1_02_in16 = reg_0628;
    119: op1_02_in16 = reg_0444;
    120: op1_02_in16 = reg_0730;
    121: op1_02_in16 = reg_0286;
    122: op1_02_in16 = reg_1032;
    125: op1_02_in16 = reg_1000;
    126: op1_02_in16 = reg_0863;
    127: op1_02_in16 = reg_0823;
    43: op1_02_in16 = reg_0566;
    128: op1_02_in16 = reg_0969;
    129: op1_02_in16 = reg_1321;
    130: op1_02_in16 = reg_0024;
    131: op1_02_in16 = reg_0201;
    default: op1_02_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_02_inv16 = 1;
    73: op1_02_inv16 = 1;
    59: op1_02_inv16 = 1;
    71: op1_02_inv16 = 1;
    48: op1_02_inv16 = 1;
    46: op1_02_inv16 = 1;
    33: op1_02_inv16 = 1;
    70: op1_02_inv16 = 1;
    44: op1_02_inv16 = 1;
    88: op1_02_inv16 = 1;
    42: op1_02_inv16 = 1;
    62: op1_02_inv16 = 1;
    63: op1_02_inv16 = 1;
    83: op1_02_inv16 = 1;
    85: op1_02_inv16 = 1;
    90: op1_02_inv16 = 1;
    66: op1_02_inv16 = 1;
    92: op1_02_inv16 = 1;
    94: op1_02_inv16 = 1;
    95: op1_02_inv16 = 1;
    96: op1_02_inv16 = 1;
    101: op1_02_inv16 = 1;
    104: op1_02_inv16 = 1;
    105: op1_02_inv16 = 1;
    106: op1_02_inv16 = 1;
    107: op1_02_inv16 = 1;
    109: op1_02_inv16 = 1;
    110: op1_02_inv16 = 1;
    112: op1_02_inv16 = 1;
    114: op1_02_inv16 = 1;
    115: op1_02_inv16 = 1;
    121: op1_02_inv16 = 1;
    124: op1_02_inv16 = 1;
    126: op1_02_inv16 = 1;
    127: op1_02_inv16 = 1;
    43: op1_02_inv16 = 1;
    129: op1_02_inv16 = 1;
    130: op1_02_inv16 = 1;
    131: op1_02_inv16 = 1;
    default: op1_02_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の17番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in17 = reg_0890;
    53: op1_02_in17 = reg_1057;
    72: op1_02_in17 = reg_0331;
    60: op1_02_in17 = reg_0331;
    55: op1_02_in17 = reg_0064;
    73: op1_02_in17 = reg_0207;
    69: op1_02_in17 = imem03_in[15:12];
    86: op1_02_in17 = reg_1430;
    59: op1_02_in17 = reg_0258;
    113: op1_02_in17 = reg_0258;
    71: op1_02_in17 = reg_0961;
    61: op1_02_in17 = reg_0260;
    33: op1_02_in17 = reg_0260;
    50: op1_02_in17 = reg_0351;
    68: op1_02_in17 = reg_0061;
    48: op1_02_in17 = reg_0782;
    74: op1_02_in17 = reg_0984;
    46: op1_02_in17 = reg_0184;
    75: op1_02_in17 = reg_1392;
    56: op1_02_in17 = reg_0084;
    87: op1_02_in17 = reg_0964;
    127: op1_02_in17 = reg_0964;
    76: op1_02_in17 = reg_0864;
    57: op1_02_in17 = reg_0970;
    70: op1_02_in17 = reg_0191;
    77: op1_02_in17 = reg_0922;
    44: op1_02_in17 = reg_0873;
    58: op1_02_in17 = reg_0480;
    88: op1_02_in17 = reg_0443;
    78: op1_02_in17 = reg_1457;
    79: op1_02_in17 = reg_0199;
    42: op1_02_in17 = reg_0026;
    80: op1_02_in17 = reg_0139;
    62: op1_02_in17 = reg_0553;
    81: op1_02_in17 = reg_0279;
    89: op1_02_in17 = reg_0034;
    63: op1_02_in17 = reg_0695;
    104: op1_02_in17 = reg_0695;
    115: op1_02_in17 = reg_0695;
    82: op1_02_in17 = reg_0236;
    83: op1_02_in17 = reg_0752;
    64: op1_02_in17 = reg_0835;
    84: op1_02_in17 = reg_1078;
    65: op1_02_in17 = reg_0052;
    85: op1_02_in17 = reg_0245;
    90: op1_02_in17 = reg_0467;
    66: op1_02_in17 = reg_0573;
    91: op1_02_in17 = reg_0570;
    67: op1_02_in17 = reg_0282;
    92: op1_02_in17 = reg_0168;
    93: op1_02_in17 = imem07_in[7:4];
    94: op1_02_in17 = reg_0251;
    95: op1_02_in17 = reg_1207;
    96: op1_02_in17 = reg_0905;
    97: op1_02_in17 = imem06_in[11:8];
    98: op1_02_in17 = imem03_in[11:8];
    99: op1_02_in17 = reg_0576;
    100: op1_02_in17 = reg_0164;
    101: op1_02_in17 = reg_0127;
    103: op1_02_in17 = reg_0242;
    105: op1_02_in17 = reg_1180;
    106: op1_02_in17 = reg_0130;
    107: op1_02_in17 = reg_0548;
    108: op1_02_in17 = reg_0073;
    109: op1_02_in17 = reg_0285;
    110: op1_02_in17 = reg_0426;
    111: op1_02_in17 = reg_0410;
    112: op1_02_in17 = reg_0211;
    114: op1_02_in17 = reg_0345;
    116: op1_02_in17 = reg_1065;
    117: op1_02_in17 = reg_0903;
    118: op1_02_in17 = reg_0876;
    119: op1_02_in17 = reg_0177;
    120: op1_02_in17 = reg_1437;
    121: op1_02_in17 = reg_0591;
    122: op1_02_in17 = reg_0385;
    124: op1_02_in17 = imem06_in[7:4];
    125: op1_02_in17 = reg_0220;
    126: op1_02_in17 = reg_1504;
    43: op1_02_in17 = reg_0333;
    128: op1_02_in17 = reg_0599;
    129: op1_02_in17 = reg_1322;
    130: op1_02_in17 = reg_0068;
    131: op1_02_in17 = reg_0416;
    default: op1_02_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv17 = 1;
    53: op1_02_inv17 = 1;
    55: op1_02_inv17 = 1;
    73: op1_02_inv17 = 1;
    86: op1_02_inv17 = 1;
    61: op1_02_inv17 = 1;
    46: op1_02_inv17 = 1;
    75: op1_02_inv17 = 1;
    87: op1_02_inv17 = 1;
    33: op1_02_inv17 = 1;
    76: op1_02_inv17 = 1;
    77: op1_02_inv17 = 1;
    44: op1_02_inv17 = 1;
    88: op1_02_inv17 = 1;
    78: op1_02_inv17 = 1;
    62: op1_02_inv17 = 1;
    89: op1_02_inv17 = 1;
    82: op1_02_inv17 = 1;
    64: op1_02_inv17 = 1;
    84: op1_02_inv17 = 1;
    65: op1_02_inv17 = 1;
    90: op1_02_inv17 = 1;
    67: op1_02_inv17 = 1;
    92: op1_02_inv17 = 1;
    93: op1_02_inv17 = 1;
    95: op1_02_inv17 = 1;
    97: op1_02_inv17 = 1;
    99: op1_02_inv17 = 1;
    100: op1_02_inv17 = 1;
    101: op1_02_inv17 = 1;
    105: op1_02_inv17 = 1;
    107: op1_02_inv17 = 1;
    112: op1_02_inv17 = 1;
    113: op1_02_inv17 = 1;
    115: op1_02_inv17 = 1;
    116: op1_02_inv17 = 1;
    117: op1_02_inv17 = 1;
    118: op1_02_inv17 = 1;
    124: op1_02_inv17 = 1;
    125: op1_02_inv17 = 1;
    126: op1_02_inv17 = 1;
    127: op1_02_inv17 = 1;
    43: op1_02_inv17 = 1;
    130: op1_02_inv17 = 1;
    131: op1_02_inv17 = 1;
    default: op1_02_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の18番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in18 = reg_0888;
    53: op1_02_in18 = reg_0994;
    72: op1_02_in18 = imem01_in[15:12];
    55: op1_02_in18 = reg_0021;
    68: op1_02_in18 = reg_0021;
    73: op1_02_in18 = reg_0037;
    69: op1_02_in18 = reg_1325;
    86: op1_02_in18 = reg_1431;
    59: op1_02_in18 = reg_1151;
    71: op1_02_in18 = reg_1432;
    61: op1_02_in18 = reg_0238;
    50: op1_02_in18 = reg_0071;
    48: op1_02_in18 = reg_0783;
    74: op1_02_in18 = reg_0161;
    96: op1_02_in18 = reg_0161;
    46: op1_02_in18 = reg_0130;
    75: op1_02_in18 = reg_0024;
    56: op1_02_in18 = reg_0483;
    87: op1_02_in18 = reg_1516;
    33: op1_02_in18 = reg_0242;
    60: op1_02_in18 = reg_0332;
    43: op1_02_in18 = reg_0332;
    76: op1_02_in18 = reg_0828;
    57: op1_02_in18 = reg_0972;
    70: op1_02_in18 = reg_1425;
    77: op1_02_in18 = reg_0225;
    44: op1_02_in18 = reg_0197;
    58: op1_02_in18 = reg_0329;
    88: op1_02_in18 = imem04_in[7:4];
    110: op1_02_in18 = imem04_in[7:4];
    78: op1_02_in18 = reg_0726;
    79: op1_02_in18 = imem03_in[7:4];
    130: op1_02_in18 = imem03_in[7:4];
    42: op1_02_in18 = reg_0595;
    80: op1_02_in18 = reg_0664;
    62: op1_02_in18 = reg_0728;
    81: op1_02_in18 = reg_0154;
    89: op1_02_in18 = reg_1338;
    63: op1_02_in18 = imem01_in[7:4];
    82: op1_02_in18 = reg_0065;
    64: op1_02_in18 = reg_0065;
    83: op1_02_in18 = reg_0827;
    84: op1_02_in18 = reg_0255;
    65: op1_02_in18 = reg_1182;
    85: op1_02_in18 = reg_0441;
    90: op1_02_in18 = reg_0062;
    66: op1_02_in18 = reg_0121;
    91: op1_02_in18 = reg_1228;
    67: op1_02_in18 = reg_0043;
    92: op1_02_in18 = reg_1515;
    93: op1_02_in18 = reg_1439;
    121: op1_02_in18 = reg_1439;
    94: op1_02_in18 = reg_0649;
    95: op1_02_in18 = reg_0054;
    97: op1_02_in18 = reg_0908;
    98: op1_02_in18 = imem03_in[15:12];
    99: op1_02_in18 = reg_0553;
    100: op1_02_in18 = reg_1258;
    101: op1_02_in18 = reg_0684;
    103: op1_02_in18 = reg_0239;
    104: op1_02_in18 = reg_1006;
    105: op1_02_in18 = reg_1163;
    106: op1_02_in18 = reg_0207;
    107: op1_02_in18 = reg_0260;
    108: op1_02_in18 = reg_0072;
    111: op1_02_in18 = reg_0072;
    109: op1_02_in18 = reg_0442;
    112: op1_02_in18 = reg_0420;
    113: op1_02_in18 = reg_0787;
    114: op1_02_in18 = reg_0323;
    115: op1_02_in18 = reg_0800;
    116: op1_02_in18 = reg_0340;
    117: op1_02_in18 = reg_0632;
    118: op1_02_in18 = reg_0306;
    119: op1_02_in18 = reg_0965;
    120: op1_02_in18 = reg_0271;
    122: op1_02_in18 = reg_0078;
    124: op1_02_in18 = reg_0270;
    125: op1_02_in18 = reg_0507;
    126: op1_02_in18 = reg_0115;
    127: op1_02_in18 = reg_0142;
    128: op1_02_in18 = reg_1040;
    129: op1_02_in18 = reg_1100;
    131: op1_02_in18 = reg_0410;
    default: op1_02_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv18 = 1;
    53: op1_02_inv18 = 1;
    73: op1_02_inv18 = 1;
    69: op1_02_inv18 = 1;
    71: op1_02_inv18 = 1;
    50: op1_02_inv18 = 1;
    68: op1_02_inv18 = 1;
    46: op1_02_inv18 = 1;
    75: op1_02_inv18 = 1;
    56: op1_02_inv18 = 1;
    70: op1_02_inv18 = 1;
    77: op1_02_inv18 = 1;
    44: op1_02_inv18 = 1;
    88: op1_02_inv18 = 1;
    78: op1_02_inv18 = 1;
    79: op1_02_inv18 = 1;
    80: op1_02_inv18 = 1;
    81: op1_02_inv18 = 1;
    89: op1_02_inv18 = 1;
    63: op1_02_inv18 = 1;
    83: op1_02_inv18 = 1;
    64: op1_02_inv18 = 1;
    65: op1_02_inv18 = 1;
    85: op1_02_inv18 = 1;
    90: op1_02_inv18 = 1;
    66: op1_02_inv18 = 1;
    67: op1_02_inv18 = 1;
    92: op1_02_inv18 = 1;
    94: op1_02_inv18 = 1;
    97: op1_02_inv18 = 1;
    98: op1_02_inv18 = 1;
    99: op1_02_inv18 = 1;
    100: op1_02_inv18 = 1;
    101: op1_02_inv18 = 1;
    103: op1_02_inv18 = 1;
    105: op1_02_inv18 = 1;
    108: op1_02_inv18 = 1;
    110: op1_02_inv18 = 1;
    113: op1_02_inv18 = 1;
    114: op1_02_inv18 = 1;
    115: op1_02_inv18 = 1;
    118: op1_02_inv18 = 1;
    120: op1_02_inv18 = 1;
    121: op1_02_inv18 = 1;
    127: op1_02_inv18 = 1;
    43: op1_02_inv18 = 1;
    128: op1_02_inv18 = 1;
    129: op1_02_inv18 = 1;
    default: op1_02_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の19番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in19 = reg_0873;
    53: op1_02_in19 = reg_0993;
    72: op1_02_in19 = reg_0715;
    59: op1_02_in19 = reg_0715;
    55: op1_02_in19 = reg_0034;
    73: op1_02_in19 = reg_0195;
    69: op1_02_in19 = reg_0143;
    86: op1_02_in19 = reg_1268;
    71: op1_02_in19 = reg_0524;
    61: op1_02_in19 = reg_0241;
    33: op1_02_in19 = reg_0241;
    113: op1_02_in19 = reg_0241;
    50: op1_02_in19 = reg_0122;
    111: op1_02_in19 = reg_0122;
    68: op1_02_in19 = reg_0578;
    48: op1_02_in19 = reg_0193;
    74: op1_02_in19 = reg_0373;
    46: op1_02_in19 = reg_0206;
    106: op1_02_in19 = reg_0206;
    75: op1_02_in19 = reg_0069;
    87: op1_02_in19 = reg_1518;
    60: op1_02_in19 = reg_0736;
    76: op1_02_in19 = reg_0037;
    57: op1_02_in19 = reg_0626;
    70: op1_02_in19 = reg_1033;
    77: op1_02_in19 = reg_0140;
    44: op1_02_in19 = reg_0118;
    58: op1_02_in19 = reg_1143;
    88: op1_02_in19 = imem04_in[15:12];
    78: op1_02_in19 = reg_0895;
    79: op1_02_in19 = reg_0541;
    130: op1_02_in19 = reg_0541;
    42: op1_02_in19 = reg_0450;
    80: op1_02_in19 = reg_0284;
    62: op1_02_in19 = reg_0402;
    81: op1_02_in19 = reg_0710;
    89: op1_02_in19 = reg_0531;
    63: op1_02_in19 = reg_0331;
    82: op1_02_in19 = reg_0470;
    83: op1_02_in19 = reg_1035;
    64: op1_02_in19 = reg_0211;
    84: op1_02_in19 = reg_1495;
    85: op1_02_in19 = reg_0366;
    90: op1_02_in19 = reg_1368;
    66: op1_02_in19 = reg_1064;
    91: op1_02_in19 = reg_0419;
    67: op1_02_in19 = reg_0011;
    92: op1_02_in19 = imem03_in[7:4];
    117: op1_02_in19 = imem03_in[7:4];
    93: op1_02_in19 = reg_0498;
    94: op1_02_in19 = reg_0182;
    95: op1_02_in19 = reg_0971;
    96: op1_02_in19 = reg_0730;
    97: op1_02_in19 = reg_0870;
    98: op1_02_in19 = reg_0505;
    99: op1_02_in19 = reg_0743;
    100: op1_02_in19 = reg_0978;
    101: op1_02_in19 = reg_0628;
    103: op1_02_in19 = reg_0238;
    104: op1_02_in19 = reg_0068;
    105: op1_02_in19 = reg_1514;
    107: op1_02_in19 = reg_0798;
    108: op1_02_in19 = reg_1321;
    109: op1_02_in19 = reg_0051;
    110: op1_02_in19 = reg_1144;
    112: op1_02_in19 = reg_0633;
    114: op1_02_in19 = reg_0296;
    115: op1_02_in19 = reg_1091;
    116: op1_02_in19 = reg_0268;
    118: op1_02_in19 = reg_0829;
    119: op1_02_in19 = reg_1184;
    120: op1_02_in19 = reg_0984;
    121: op1_02_in19 = reg_0002;
    122: op1_02_in19 = reg_0403;
    124: op1_02_in19 = reg_0929;
    125: op1_02_in19 = reg_0191;
    126: op1_02_in19 = reg_0718;
    127: op1_02_in19 = reg_0314;
    43: op1_02_in19 = reg_0317;
    128: op1_02_in19 = reg_1419;
    129: op1_02_in19 = imem01_in[3:0];
    131: op1_02_in19 = reg_0134;
    default: op1_02_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_02_inv19 = 1;
    73: op1_02_inv19 = 1;
    69: op1_02_inv19 = 1;
    86: op1_02_inv19 = 1;
    50: op1_02_inv19 = 1;
    46: op1_02_inv19 = 1;
    76: op1_02_inv19 = 1;
    70: op1_02_inv19 = 1;
    58: op1_02_inv19 = 1;
    78: op1_02_inv19 = 1;
    81: op1_02_inv19 = 1;
    63: op1_02_inv19 = 1;
    82: op1_02_inv19 = 1;
    64: op1_02_inv19 = 1;
    84: op1_02_inv19 = 1;
    85: op1_02_inv19 = 1;
    93: op1_02_inv19 = 1;
    95: op1_02_inv19 = 1;
    96: op1_02_inv19 = 1;
    101: op1_02_inv19 = 1;
    103: op1_02_inv19 = 1;
    106: op1_02_inv19 = 1;
    108: op1_02_inv19 = 1;
    110: op1_02_inv19 = 1;
    112: op1_02_inv19 = 1;
    114: op1_02_inv19 = 1;
    121: op1_02_inv19 = 1;
    43: op1_02_inv19 = 1;
    128: op1_02_inv19 = 1;
    129: op1_02_inv19 = 1;
    130: op1_02_inv19 = 1;
    default: op1_02_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の20番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in20 = reg_0130;
    53: op1_02_in20 = reg_0995;
    72: op1_02_in20 = reg_1452;
    55: op1_02_in20 = reg_0792;
    73: op1_02_in20 = reg_0377;
    69: op1_02_in20 = reg_0144;
    86: op1_02_in20 = reg_1169;
    59: op1_02_in20 = reg_0819;
    42: op1_02_in20 = reg_0819;
    71: op1_02_in20 = reg_1405;
    61: op1_02_in20 = reg_0609;
    50: op1_02_in20 = reg_0612;
    68: op1_02_in20 = reg_1299;
    48: op1_02_in20 = reg_0192;
    74: op1_02_in20 = reg_0295;
    46: op1_02_in20 = reg_0039;
    76: op1_02_in20 = reg_0039;
    75: op1_02_in20 = imem02_in[3:0];
    87: op1_02_in20 = reg_1314;
    33: op1_02_in20 = reg_0222;
    67: op1_02_in20 = reg_0222;
    60: op1_02_in20 = reg_0828;
    57: op1_02_in20 = reg_0125;
    70: op1_02_in20 = reg_0962;
    79: op1_02_in20 = reg_0962;
    77: op1_02_in20 = reg_0779;
    44: op1_02_in20 = reg_0861;
    58: op1_02_in20 = reg_0534;
    88: op1_02_in20 = reg_1312;
    116: op1_02_in20 = reg_1312;
    78: op1_02_in20 = reg_0010;
    80: op1_02_in20 = reg_0285;
    62: op1_02_in20 = reg_0403;
    81: op1_02_in20 = reg_0216;
    89: op1_02_in20 = reg_0552;
    63: op1_02_in20 = reg_0238;
    82: op1_02_in20 = reg_0370;
    83: op1_02_in20 = reg_0717;
    64: op1_02_in20 = reg_0020;
    84: op1_02_in20 = imem03_in[7:4];
    85: op1_02_in20 = reg_0741;
    90: op1_02_in20 = reg_0535;
    66: op1_02_in20 = reg_1325;
    91: op1_02_in20 = reg_0165;
    92: op1_02_in20 = reg_0121;
    93: op1_02_in20 = reg_1414;
    94: op1_02_in20 = reg_0564;
    95: op1_02_in20 = reg_1458;
    96: op1_02_in20 = reg_0751;
    97: op1_02_in20 = reg_0960;
    98: op1_02_in20 = reg_0889;
    99: op1_02_in20 = reg_0966;
    100: op1_02_in20 = reg_0297;
    101: op1_02_in20 = reg_0007;
    103: op1_02_in20 = reg_0241;
    104: op1_02_in20 = reg_0227;
    115: op1_02_in20 = reg_0227;
    105: op1_02_in20 = reg_0090;
    106: op1_02_in20 = imem06_in[11:8];
    107: op1_02_in20 = reg_0742;
    108: op1_02_in20 = reg_0027;
    109: op1_02_in20 = reg_0004;
    110: op1_02_in20 = reg_1369;
    111: op1_02_in20 = imem01_in[3:0];
    112: op1_02_in20 = imem05_in[15:12];
    113: op1_02_in20 = reg_0798;
    114: op1_02_in20 = reg_0371;
    117: op1_02_in20 = reg_0559;
    118: op1_02_in20 = reg_0745;
    119: op1_02_in20 = reg_0070;
    120: op1_02_in20 = reg_1467;
    122: op1_02_in20 = reg_0044;
    124: op1_02_in20 = reg_0870;
    125: op1_02_in20 = reg_0375;
    126: op1_02_in20 = reg_0714;
    127: op1_02_in20 = reg_0349;
    43: op1_02_in20 = reg_0315;
    128: op1_02_in20 = reg_0582;
    129: op1_02_in20 = reg_0610;
    130: op1_02_in20 = reg_0246;
    131: op1_02_in20 = reg_0389;
    default: op1_02_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv20 = 1;
    53: op1_02_inv20 = 1;
    72: op1_02_inv20 = 1;
    69: op1_02_inv20 = 1;
    50: op1_02_inv20 = 1;
    68: op1_02_inv20 = 1;
    75: op1_02_inv20 = 1;
    87: op1_02_inv20 = 1;
    33: op1_02_inv20 = 1;
    60: op1_02_inv20 = 1;
    57: op1_02_inv20 = 1;
    70: op1_02_inv20 = 1;
    88: op1_02_inv20 = 1;
    78: op1_02_inv20 = 1;
    79: op1_02_inv20 = 1;
    62: op1_02_inv20 = 1;
    81: op1_02_inv20 = 1;
    89: op1_02_inv20 = 1;
    63: op1_02_inv20 = 1;
    64: op1_02_inv20 = 1;
    84: op1_02_inv20 = 1;
    85: op1_02_inv20 = 1;
    67: op1_02_inv20 = 1;
    92: op1_02_inv20 = 1;
    93: op1_02_inv20 = 1;
    95: op1_02_inv20 = 1;
    96: op1_02_inv20 = 1;
    97: op1_02_inv20 = 1;
    99: op1_02_inv20 = 1;
    101: op1_02_inv20 = 1;
    103: op1_02_inv20 = 1;
    105: op1_02_inv20 = 1;
    107: op1_02_inv20 = 1;
    108: op1_02_inv20 = 1;
    109: op1_02_inv20 = 1;
    110: op1_02_inv20 = 1;
    111: op1_02_inv20 = 1;
    112: op1_02_inv20 = 1;
    114: op1_02_inv20 = 1;
    117: op1_02_inv20 = 1;
    118: op1_02_inv20 = 1;
    119: op1_02_inv20 = 1;
    125: op1_02_inv20 = 1;
    126: op1_02_inv20 = 1;
    127: op1_02_inv20 = 1;
    128: op1_02_inv20 = 1;
    131: op1_02_inv20 = 1;
    default: op1_02_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の21番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in21 = reg_0206;
    53: op1_02_in21 = reg_0867;
    72: op1_02_in21 = reg_0147;
    55: op1_02_in21 = reg_0793;
    73: op1_02_in21 = reg_0120;
    69: op1_02_in21 = reg_0891;
    81: op1_02_in21 = reg_0891;
    86: op1_02_in21 = reg_0992;
    59: op1_02_in21 = reg_0930;
    71: op1_02_in21 = reg_0476;
    61: op1_02_in21 = reg_0982;
    50: op1_02_in21 = reg_0609;
    68: op1_02_in21 = reg_0251;
    48: op1_02_in21 = imem06_in[7:4];
    74: op1_02_in21 = reg_0165;
    46: op1_02_in21 = reg_0195;
    75: op1_02_in21 = reg_0840;
    87: op1_02_in21 = reg_1313;
    33: op1_02_in21 = reg_0451;
    60: op1_02_in21 = reg_0832;
    76: op1_02_in21 = reg_1426;
    57: op1_02_in21 = reg_0056;
    70: op1_02_in21 = reg_0478;
    77: op1_02_in21 = reg_0665;
    44: op1_02_in21 = reg_0754;
    114: op1_02_in21 = reg_0754;
    58: op1_02_in21 = reg_0595;
    88: op1_02_in21 = reg_1383;
    78: op1_02_in21 = reg_0679;
    79: op1_02_in21 = reg_0143;
    42: op1_02_in21 = reg_0167;
    80: op1_02_in21 = reg_0740;
    62: op1_02_in21 = reg_0383;
    89: op1_02_in21 = reg_1200;
    63: op1_02_in21 = reg_1151;
    82: op1_02_in21 = reg_0708;
    83: op1_02_in21 = reg_0585;
    126: op1_02_in21 = reg_0585;
    64: op1_02_in21 = reg_0033;
    84: op1_02_in21 = imem03_in[11:8];
    85: op1_02_in21 = reg_0415;
    90: op1_02_in21 = reg_1339;
    66: op1_02_in21 = reg_0349;
    91: op1_02_in21 = reg_1202;
    67: op1_02_in21 = reg_0662;
    92: op1_02_in21 = reg_0154;
    98: op1_02_in21 = reg_0154;
    93: op1_02_in21 = reg_0298;
    94: op1_02_in21 = reg_0697;
    95: op1_02_in21 = reg_0105;
    96: op1_02_in21 = reg_0720;
    97: op1_02_in21 = reg_1326;
    99: op1_02_in21 = reg_0968;
    100: op1_02_in21 = reg_1214;
    101: op1_02_in21 = reg_0024;
    103: op1_02_in21 = reg_0830;
    104: op1_02_in21 = imem03_in[15:12];
    105: op1_02_in21 = reg_0736;
    106: op1_02_in21 = reg_0795;
    107: op1_02_in21 = reg_1474;
    108: op1_02_in21 = imem01_in[15:12];
    109: op1_02_in21 = reg_0003;
    110: op1_02_in21 = reg_1367;
    111: op1_02_in21 = imem01_in[7:4];
    112: op1_02_in21 = reg_0367;
    113: op1_02_in21 = reg_0820;
    115: op1_02_in21 = reg_0168;
    116: op1_02_in21 = reg_0256;
    117: op1_02_in21 = reg_0709;
    118: op1_02_in21 = reg_0897;
    119: op1_02_in21 = reg_0314;
    120: op1_02_in21 = reg_0869;
    122: op1_02_in21 = reg_0041;
    124: op1_02_in21 = reg_0974;
    125: op1_02_in21 = reg_1494;
    127: op1_02_in21 = reg_0954;
    43: op1_02_in21 = reg_0318;
    128: op1_02_in21 = reg_0268;
    129: op1_02_in21 = reg_0787;
    130: op1_02_in21 = reg_0732;
    131: op1_02_in21 = reg_0060;
    default: op1_02_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_02_inv21 = 1;
    59: op1_02_inv21 = 1;
    71: op1_02_inv21 = 1;
    61: op1_02_inv21 = 1;
    68: op1_02_inv21 = 1;
    74: op1_02_inv21 = 1;
    46: op1_02_inv21 = 1;
    75: op1_02_inv21 = 1;
    57: op1_02_inv21 = 1;
    70: op1_02_inv21 = 1;
    44: op1_02_inv21 = 1;
    58: op1_02_inv21 = 1;
    79: op1_02_inv21 = 1;
    63: op1_02_inv21 = 1;
    82: op1_02_inv21 = 1;
    85: op1_02_inv21 = 1;
    66: op1_02_inv21 = 1;
    91: op1_02_inv21 = 1;
    93: op1_02_inv21 = 1;
    97: op1_02_inv21 = 1;
    98: op1_02_inv21 = 1;
    100: op1_02_inv21 = 1;
    103: op1_02_inv21 = 1;
    104: op1_02_inv21 = 1;
    105: op1_02_inv21 = 1;
    107: op1_02_inv21 = 1;
    108: op1_02_inv21 = 1;
    109: op1_02_inv21 = 1;
    111: op1_02_inv21 = 1;
    114: op1_02_inv21 = 1;
    115: op1_02_inv21 = 1;
    116: op1_02_inv21 = 1;
    119: op1_02_inv21 = 1;
    122: op1_02_inv21 = 1;
    128: op1_02_inv21 = 1;
    default: op1_02_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の22番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in22 = imem06_in[15:12];
    48: op1_02_in22 = imem06_in[15:12];
    53: op1_02_in22 = reg_0156;
    72: op1_02_in22 = reg_0899;
    55: op1_02_in22 = reg_0733;
    73: op1_02_in22 = reg_0192;
    69: op1_02_in22 = reg_0142;
    86: op1_02_in22 = reg_0648;
    59: op1_02_in22 = reg_0402;
    71: op1_02_in22 = reg_0928;
    61: op1_02_in22 = reg_0439;
    50: op1_02_in22 = reg_0335;
    68: op1_02_in22 = reg_0273;
    74: op1_02_in22 = reg_0583;
    46: op1_02_in22 = reg_0161;
    33: op1_02_in22 = reg_0161;
    75: op1_02_in22 = reg_0699;
    87: op1_02_in22 = reg_1226;
    127: op1_02_in22 = reg_1226;
    60: op1_02_in22 = reg_0646;
    76: op1_02_in22 = reg_0133;
    57: op1_02_in22 = reg_0845;
    70: op1_02_in22 = reg_0840;
    77: op1_02_in22 = reg_0441;
    44: op1_02_in22 = imem06_in[7:4];
    58: op1_02_in22 = reg_0268;
    88: op1_02_in22 = reg_1372;
    78: op1_02_in22 = reg_1139;
    79: op1_02_in22 = reg_0180;
    42: op1_02_in22 = reg_0120;
    108: op1_02_in22 = reg_0120;
    80: op1_02_in22 = reg_0404;
    62: op1_02_in22 = reg_0362;
    81: op1_02_in22 = reg_0789;
    89: op1_02_in22 = reg_0094;
    63: op1_02_in22 = reg_1152;
    82: op1_02_in22 = reg_0205;
    83: op1_02_in22 = reg_0586;
    64: op1_02_in22 = reg_0793;
    84: op1_02_in22 = reg_0179;
    85: op1_02_in22 = reg_0592;
    90: op1_02_in22 = reg_0978;
    66: op1_02_in22 = reg_1301;
    91: op1_02_in22 = reg_0270;
    67: op1_02_in22 = reg_0606;
    92: op1_02_in22 = reg_0311;
    93: op1_02_in22 = reg_0135;
    94: op1_02_in22 = reg_0938;
    95: op1_02_in22 = reg_0876;
    96: op1_02_in22 = reg_0859;
    97: op1_02_in22 = reg_0720;
    98: op1_02_in22 = reg_0573;
    99: op1_02_in22 = reg_0360;
    100: op1_02_in22 = reg_1040;
    101: op1_02_in22 = reg_0563;
    103: op1_02_in22 = reg_0798;
    104: op1_02_in22 = reg_0216;
    105: op1_02_in22 = reg_0450;
    106: op1_02_in22 = reg_0908;
    107: op1_02_in22 = reg_1457;
    109: op1_02_in22 = reg_0002;
    110: op1_02_in22 = reg_0493;
    111: op1_02_in22 = reg_0985;
    112: op1_02_in22 = reg_0333;
    113: op1_02_in22 = reg_1473;
    114: op1_02_in22 = reg_0046;
    115: op1_02_in22 = imem03_in[3:0];
    116: op1_02_in22 = reg_0117;
    117: op1_02_in22 = reg_0597;
    118: op1_02_in22 = reg_0560;
    119: op1_02_in22 = reg_0957;
    120: op1_02_in22 = reg_1505;
    122: op1_02_in22 = reg_0012;
    124: op1_02_in22 = reg_0696;
    125: op1_02_in22 = reg_0965;
    126: op1_02_in22 = reg_0571;
    43: op1_02_in22 = reg_0540;
    128: op1_02_in22 = reg_0932;
    129: op1_02_in22 = reg_0609;
    130: op1_02_in22 = reg_1003;
    131: op1_02_in22 = reg_0072;
    default: op1_02_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_02_inv22 = 1;
    72: op1_02_inv22 = 1;
    69: op1_02_inv22 = 1;
    86: op1_02_inv22 = 1;
    74: op1_02_inv22 = 1;
    46: op1_02_inv22 = 1;
    75: op1_02_inv22 = 1;
    33: op1_02_inv22 = 1;
    60: op1_02_inv22 = 1;
    44: op1_02_inv22 = 1;
    88: op1_02_inv22 = 1;
    78: op1_02_inv22 = 1;
    42: op1_02_inv22 = 1;
    80: op1_02_inv22 = 1;
    62: op1_02_inv22 = 1;
    81: op1_02_inv22 = 1;
    82: op1_02_inv22 = 1;
    85: op1_02_inv22 = 1;
    92: op1_02_inv22 = 1;
    97: op1_02_inv22 = 1;
    98: op1_02_inv22 = 1;
    99: op1_02_inv22 = 1;
    101: op1_02_inv22 = 1;
    103: op1_02_inv22 = 1;
    104: op1_02_inv22 = 1;
    108: op1_02_inv22 = 1;
    109: op1_02_inv22 = 1;
    110: op1_02_inv22 = 1;
    113: op1_02_inv22 = 1;
    116: op1_02_inv22 = 1;
    117: op1_02_inv22 = 1;
    118: op1_02_inv22 = 1;
    119: op1_02_inv22 = 1;
    124: op1_02_inv22 = 1;
    125: op1_02_inv22 = 1;
    126: op1_02_inv22 = 1;
    128: op1_02_inv22 = 1;
    131: op1_02_inv22 = 1;
    default: op1_02_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の23番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in23 = reg_1105;
    53: op1_02_in23 = reg_0921;
    72: op1_02_in23 = reg_0257;
    55: op1_02_in23 = reg_1059;
    73: op1_02_in23 = reg_0870;
    69: op1_02_in23 = reg_1003;
    79: op1_02_in23 = reg_1003;
    86: op1_02_in23 = reg_0604;
    59: op1_02_in23 = reg_0385;
    71: op1_02_in23 = reg_0883;
    61: op1_02_in23 = reg_0430;
    50: op1_02_in23 = reg_0595;
    68: op1_02_in23 = reg_0702;
    48: op1_02_in23 = reg_0133;
    74: op1_02_in23 = reg_0215;
    46: op1_02_in23 = imem06_in[11:8];
    75: op1_02_in23 = reg_0198;
    87: op1_02_in23 = reg_0884;
    33: op1_02_in23 = reg_0147;
    60: op1_02_in23 = reg_0745;
    76: op1_02_in23 = reg_0161;
    57: op1_02_in23 = reg_0311;
    70: op1_02_in23 = reg_0488;
    77: op1_02_in23 = reg_0413;
    44: op1_02_in23 = reg_0141;
    58: op1_02_in23 = reg_1198;
    88: op1_02_in23 = reg_1368;
    78: op1_02_in23 = reg_0276;
    42: op1_02_in23 = reg_0258;
    80: op1_02_in23 = reg_0415;
    62: op1_02_in23 = reg_0360;
    81: op1_02_in23 = reg_0375;
    89: op1_02_in23 = reg_0412;
    63: op1_02_in23 = reg_0080;
    82: op1_02_in23 = reg_0750;
    127: op1_02_in23 = reg_0750;
    83: op1_02_in23 = reg_0528;
    64: op1_02_in23 = reg_0205;
    84: op1_02_in23 = reg_1448;
    85: op1_02_in23 = reg_0051;
    90: op1_02_in23 = reg_0552;
    66: op1_02_in23 = reg_0558;
    91: op1_02_in23 = reg_0023;
    67: op1_02_in23 = reg_0533;
    92: op1_02_in23 = reg_0789;
    93: op1_02_in23 = reg_1440;
    94: op1_02_in23 = reg_0418;
    95: op1_02_in23 = reg_0307;
    96: op1_02_in23 = reg_0752;
    97: op1_02_in23 = reg_0116;
    98: op1_02_in23 = reg_1063;
    99: op1_02_in23 = reg_0899;
    100: op1_02_in23 = reg_0232;
    101: op1_02_in23 = reg_0168;
    103: op1_02_in23 = reg_0742;
    129: op1_02_in23 = reg_0742;
    104: op1_02_in23 = reg_0847;
    105: op1_02_in23 = reg_0197;
    106: op1_02_in23 = reg_0192;
    107: op1_02_in23 = reg_1456;
    108: op1_02_in23 = reg_1256;
    109: op1_02_in23 = reg_0519;
    110: op1_02_in23 = reg_0034;
    111: op1_02_in23 = reg_0547;
    112: op1_02_in23 = reg_0272;
    113: op1_02_in23 = reg_1474;
    114: op1_02_in23 = reg_0214;
    115: op1_02_in23 = reg_0699;
    116: op1_02_in23 = reg_0063;
    117: op1_02_in23 = reg_0177;
    118: op1_02_in23 = reg_0903;
    119: op1_02_in23 = reg_0952;
    120: op1_02_in23 = reg_1504;
    122: op1_02_in23 = reg_0011;
    124: op1_02_in23 = reg_1323;
    125: op1_02_in23 = reg_0314;
    126: op1_02_in23 = reg_0569;
    43: op1_02_in23 = imem05_in[7:4];
    128: op1_02_in23 = reg_0633;
    130: op1_02_in23 = reg_0573;
    131: op1_02_in23 = reg_1324;
    default: op1_02_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_02_inv23 = 1;
    55: op1_02_inv23 = 1;
    86: op1_02_inv23 = 1;
    59: op1_02_inv23 = 1;
    71: op1_02_inv23 = 1;
    68: op1_02_inv23 = 1;
    48: op1_02_inv23 = 1;
    74: op1_02_inv23 = 1;
    46: op1_02_inv23 = 1;
    75: op1_02_inv23 = 1;
    33: op1_02_inv23 = 1;
    76: op1_02_inv23 = 1;
    57: op1_02_inv23 = 1;
    77: op1_02_inv23 = 1;
    78: op1_02_inv23 = 1;
    79: op1_02_inv23 = 1;
    62: op1_02_inv23 = 1;
    81: op1_02_inv23 = 1;
    89: op1_02_inv23 = 1;
    63: op1_02_inv23 = 1;
    64: op1_02_inv23 = 1;
    93: op1_02_inv23 = 1;
    97: op1_02_inv23 = 1;
    98: op1_02_inv23 = 1;
    103: op1_02_inv23 = 1;
    104: op1_02_inv23 = 1;
    105: op1_02_inv23 = 1;
    106: op1_02_inv23 = 1;
    107: op1_02_inv23 = 1;
    108: op1_02_inv23 = 1;
    109: op1_02_inv23 = 1;
    114: op1_02_inv23 = 1;
    119: op1_02_inv23 = 1;
    120: op1_02_inv23 = 1;
    122: op1_02_inv23 = 1;
    126: op1_02_inv23 = 1;
    43: op1_02_inv23 = 1;
    128: op1_02_inv23 = 1;
    129: op1_02_inv23 = 1;
    131: op1_02_inv23 = 1;
    default: op1_02_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の24番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in24 = reg_0192;
    53: op1_02_in24 = reg_0437;
    72: op1_02_in24 = reg_0077;
    55: op1_02_in24 = reg_0831;
    73: op1_02_in24 = imem06_in[15:12];
    69: op1_02_in24 = reg_0349;
    86: op1_02_in24 = reg_0173;
    59: op1_02_in24 = reg_0362;
    71: op1_02_in24 = reg_0353;
    61: op1_02_in24 = reg_0726;
    50: op1_02_in24 = reg_0695;
    68: op1_02_in24 = imem05_in[7:4];
    48: op1_02_in24 = reg_0907;
    74: op1_02_in24 = imem07_in[15:12];
    46: op1_02_in24 = reg_0859;
    75: op1_02_in24 = reg_0232;
    87: op1_02_in24 = reg_0288;
    33: op1_02_in24 = reg_0403;
    60: op1_02_in24 = reg_1181;
    76: op1_02_in24 = reg_1303;
    57: op1_02_in24 = reg_0734;
    70: op1_02_in24 = reg_1312;
    77: op1_02_in24 = reg_0321;
    44: op1_02_in24 = reg_0397;
    58: op1_02_in24 = reg_1077;
    90: op1_02_in24 = reg_1077;
    88: op1_02_in24 = reg_0088;
    78: op1_02_in24 = reg_0934;
    79: op1_02_in24 = reg_0965;
    42: op1_02_in24 = reg_0746;
    80: op1_02_in24 = reg_0623;
    62: op1_02_in24 = reg_0093;
    81: op1_02_in24 = reg_1003;
    92: op1_02_in24 = reg_1003;
    89: op1_02_in24 = reg_0407;
    63: op1_02_in24 = reg_0283;
    82: op1_02_in24 = reg_1298;
    83: op1_02_in24 = reg_0529;
    64: op1_02_in24 = reg_0750;
    84: op1_02_in24 = reg_0557;
    85: op1_02_in24 = reg_0001;
    66: op1_02_in24 = reg_0328;
    91: op1_02_in24 = reg_0215;
    67: op1_02_in24 = reg_0253;
    93: op1_02_in24 = reg_0703;
    94: op1_02_in24 = reg_0872;
    95: op1_02_in24 = reg_0306;
    96: op1_02_in24 = reg_1501;
    97: op1_02_in24 = reg_0398;
    98: op1_02_in24 = reg_0177;
    99: op1_02_in24 = reg_0335;
    100: op1_02_in24 = reg_0582;
    101: op1_02_in24 = reg_1515;
    103: op1_02_in24 = reg_0468;
    104: op1_02_in24 = reg_0311;
    105: op1_02_in24 = reg_0344;
    106: op1_02_in24 = reg_0316;
    107: op1_02_in24 = reg_0147;
    108: op1_02_in24 = reg_0874;
    110: op1_02_in24 = reg_0531;
    111: op1_02_in24 = reg_0260;
    112: op1_02_in24 = reg_0066;
    113: op1_02_in24 = reg_0819;
    114: op1_02_in24 = reg_1170;
    115: op1_02_in24 = reg_0732;
    116: op1_02_in24 = reg_1502;
    117: op1_02_in24 = reg_0847;
    118: op1_02_in24 = reg_1078;
    119: op1_02_in24 = reg_0756;
    120: op1_02_in24 = reg_0780;
    122: op1_02_in24 = reg_0662;
    124: op1_02_in24 = reg_0752;
    125: op1_02_in24 = reg_0627;
    126: op1_02_in24 = reg_0296;
    127: op1_02_in24 = reg_0673;
    43: op1_02_in24 = reg_0251;
    128: op1_02_in24 = reg_0021;
    129: op1_02_in24 = reg_0715;
    130: op1_02_in24 = reg_0597;
    131: op1_02_in24 = imem01_in[11:8];
    default: op1_02_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_02_inv24 = 1;
    55: op1_02_inv24 = 1;
    73: op1_02_inv24 = 1;
    86: op1_02_inv24 = 1;
    61: op1_02_inv24 = 1;
    50: op1_02_inv24 = 1;
    68: op1_02_inv24 = 1;
    48: op1_02_inv24 = 1;
    74: op1_02_inv24 = 1;
    75: op1_02_inv24 = 1;
    87: op1_02_inv24 = 1;
    60: op1_02_inv24 = 1;
    57: op1_02_inv24 = 1;
    70: op1_02_inv24 = 1;
    44: op1_02_inv24 = 1;
    58: op1_02_inv24 = 1;
    88: op1_02_inv24 = 1;
    78: op1_02_inv24 = 1;
    79: op1_02_inv24 = 1;
    89: op1_02_inv24 = 1;
    83: op1_02_inv24 = 1;
    84: op1_02_inv24 = 1;
    66: op1_02_inv24 = 1;
    91: op1_02_inv24 = 1;
    92: op1_02_inv24 = 1;
    94: op1_02_inv24 = 1;
    98: op1_02_inv24 = 1;
    103: op1_02_inv24 = 1;
    104: op1_02_inv24 = 1;
    105: op1_02_inv24 = 1;
    114: op1_02_inv24 = 1;
    115: op1_02_inv24 = 1;
    117: op1_02_inv24 = 1;
    119: op1_02_inv24 = 1;
    120: op1_02_inv24 = 1;
    122: op1_02_inv24 = 1;
    124: op1_02_inv24 = 1;
    125: op1_02_inv24 = 1;
    126: op1_02_inv24 = 1;
    129: op1_02_inv24 = 1;
    130: op1_02_inv24 = 1;
    131: op1_02_inv24 = 1;
    default: op1_02_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の25番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in25 = reg_0870;
    53: op1_02_in25 = reg_0137;
    72: op1_02_in25 = reg_0079;
    55: op1_02_in25 = reg_0700;
    73: op1_02_in25 = reg_0109;
    69: op1_02_in25 = reg_0597;
    86: op1_02_in25 = reg_0045;
    59: op1_02_in25 = reg_0360;
    71: op1_02_in25 = reg_0188;
    61: op1_02_in25 = reg_0148;
    50: op1_02_in25 = imem01_in[3:0];
    68: op1_02_in25 = imem05_in[15:12];
    48: op1_02_in25 = reg_0696;
    74: op1_02_in25 = reg_0461;
    46: op1_02_in25 = reg_0714;
    75: op1_02_in25 = reg_0375;
    87: op1_02_in25 = imem04_in[15:12];
    33: op1_02_in25 = reg_0401;
    60: op1_02_in25 = reg_1180;
    76: op1_02_in25 = reg_0637;
    57: op1_02_in25 = reg_0556;
    70: op1_02_in25 = reg_1384;
    77: op1_02_in25 = reg_0361;
    44: op1_02_in25 = reg_0396;
    58: op1_02_in25 = reg_1082;
    88: op1_02_in25 = reg_0034;
    78: op1_02_in25 = reg_0981;
    79: op1_02_in25 = reg_0048;
    42: op1_02_in25 = reg_0742;
    80: op1_02_in25 = reg_0620;
    62: op1_02_in25 = reg_0875;
    81: op1_02_in25 = reg_0329;
    119: op1_02_in25 = reg_0329;
    89: op1_02_in25 = reg_0598;
    63: op1_02_in25 = reg_0184;
    82: op1_02_in25 = reg_1431;
    83: op1_02_in25 = reg_1228;
    64: op1_02_in25 = reg_0736;
    84: op1_02_in25 = reg_0962;
    85: op1_02_in25 = reg_0085;
    90: op1_02_in25 = reg_1065;
    66: op1_02_in25 = reg_1282;
    91: op1_02_in25 = imem07_in[11:8];
    114: op1_02_in25 = imem07_in[11:8];
    67: op1_02_in25 = reg_1343;
    92: op1_02_in25 = reg_0954;
    93: op1_02_in25 = reg_0851;
    94: op1_02_in25 = reg_0118;
    95: op1_02_in25 = reg_0745;
    96: op1_02_in25 = reg_0635;
    97: op1_02_in25 = reg_0374;
    98: op1_02_in25 = reg_0198;
    99: op1_02_in25 = reg_0077;
    100: op1_02_in25 = reg_0340;
    101: op1_02_in25 = imem03_in[3:0];
    103: op1_02_in25 = reg_0469;
    111: op1_02_in25 = reg_0469;
    104: op1_02_in25 = reg_0191;
    105: op1_02_in25 = reg_0589;
    106: op1_02_in25 = reg_0974;
    107: op1_02_in25 = reg_0146;
    108: op1_02_in25 = reg_1290;
    110: op1_02_in25 = reg_0297;
    112: op1_02_in25 = reg_0604;
    113: op1_02_in25 = reg_0149;
    115: op1_02_in25 = reg_0847;
    116: op1_02_in25 = imem05_in[3:0];
    117: op1_02_in25 = reg_0312;
    118: op1_02_in25 = reg_0563;
    120: op1_02_in25 = reg_0716;
    122: op1_02_in25 = imem02_in[7:4];
    124: op1_02_in25 = reg_0115;
    125: op1_02_in25 = reg_1447;
    126: op1_02_in25 = reg_0119;
    127: op1_02_in25 = reg_1325;
    43: op1_02_in25 = reg_0197;
    128: op1_02_in25 = reg_0035;
    129: op1_02_in25 = reg_0434;
    130: op1_02_in25 = reg_0220;
    131: op1_02_in25 = reg_0577;
    default: op1_02_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv25 = 1;
    53: op1_02_inv25 = 1;
    55: op1_02_inv25 = 1;
    86: op1_02_inv25 = 1;
    59: op1_02_inv25 = 1;
    71: op1_02_inv25 = 1;
    61: op1_02_inv25 = 1;
    50: op1_02_inv25 = 1;
    68: op1_02_inv25 = 1;
    48: op1_02_inv25 = 1;
    75: op1_02_inv25 = 1;
    33: op1_02_inv25 = 1;
    57: op1_02_inv25 = 1;
    70: op1_02_inv25 = 1;
    44: op1_02_inv25 = 1;
    88: op1_02_inv25 = 1;
    78: op1_02_inv25 = 1;
    79: op1_02_inv25 = 1;
    62: op1_02_inv25 = 1;
    63: op1_02_inv25 = 1;
    64: op1_02_inv25 = 1;
    85: op1_02_inv25 = 1;
    90: op1_02_inv25 = 1;
    66: op1_02_inv25 = 1;
    91: op1_02_inv25 = 1;
    67: op1_02_inv25 = 1;
    92: op1_02_inv25 = 1;
    94: op1_02_inv25 = 1;
    97: op1_02_inv25 = 1;
    98: op1_02_inv25 = 1;
    99: op1_02_inv25 = 1;
    101: op1_02_inv25 = 1;
    103: op1_02_inv25 = 1;
    105: op1_02_inv25 = 1;
    107: op1_02_inv25 = 1;
    108: op1_02_inv25 = 1;
    110: op1_02_inv25 = 1;
    112: op1_02_inv25 = 1;
    114: op1_02_inv25 = 1;
    120: op1_02_inv25 = 1;
    125: op1_02_inv25 = 1;
    126: op1_02_inv25 = 1;
    43: op1_02_inv25 = 1;
    128: op1_02_inv25 = 1;
    129: op1_02_inv25 = 1;
    131: op1_02_inv25 = 1;
    default: op1_02_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の26番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in26 = reg_0720;
    53: op1_02_in26 = reg_0103;
    72: op1_02_in26 = reg_0010;
    55: op1_02_in26 = reg_0346;
    73: op1_02_in26 = reg_0141;
    69: op1_02_in26 = reg_0329;
    86: op1_02_in26 = reg_0167;
    59: op1_02_in26 = reg_0363;
    71: op1_02_in26 = reg_0440;
    61: op1_02_in26 = reg_0402;
    50: op1_02_in26 = reg_0602;
    68: op1_02_in26 = reg_0347;
    48: op1_02_in26 = reg_0870;
    74: op1_02_in26 = reg_0922;
    46: op1_02_in26 = reg_0670;
    75: op1_02_in26 = reg_0376;
    87: op1_02_in26 = reg_1372;
    33: op1_02_in26 = reg_0384;
    60: op1_02_in26 = reg_0318;
    76: op1_02_in26 = reg_0622;
    57: op1_02_in26 = reg_0707;
    70: op1_02_in26 = reg_0032;
    77: op1_02_in26 = reg_0050;
    44: op1_02_in26 = reg_0371;
    58: op1_02_in26 = reg_0798;
    88: op1_02_in26 = reg_1258;
    78: op1_02_in26 = reg_1207;
    79: op1_02_in26 = reg_1384;
    42: op1_02_in26 = reg_0728;
    80: op1_02_in26 = reg_0100;
    62: op1_02_in26 = reg_0290;
    103: op1_02_in26 = reg_0290;
    81: op1_02_in26 = reg_0558;
    89: op1_02_in26 = reg_1040;
    63: op1_02_in26 = reg_0606;
    82: op1_02_in26 = reg_0832;
    83: op1_02_in26 = reg_1202;
    64: op1_02_in26 = reg_0649;
    84: op1_02_in26 = reg_0375;
    85: op1_02_in26 = reg_0520;
    90: op1_02_in26 = reg_0369;
    66: op1_02_in26 = reg_0348;
    91: op1_02_in26 = reg_0490;
    67: op1_02_in26 = reg_0474;
    92: op1_02_in26 = reg_0597;
    93: op1_02_in26 = reg_0457;
    94: op1_02_in26 = reg_0014;
    95: op1_02_in26 = reg_1492;
    96: op1_02_in26 = reg_0110;
    97: op1_02_in26 = reg_0526;
    98: op1_02_in26 = reg_1001;
    99: op1_02_in26 = reg_0043;
    100: op1_02_in26 = reg_0837;
    101: op1_02_in26 = imem03_in[7:4];
    104: op1_02_in26 = reg_0234;
    105: op1_02_in26 = reg_0151;
    106: op1_02_in26 = reg_0751;
    107: op1_02_in26 = reg_0901;
    108: op1_02_in26 = reg_0401;
    110: op1_02_in26 = reg_0598;
    111: op1_02_in26 = reg_0146;
    112: op1_02_in26 = reg_0045;
    113: op1_02_in26 = reg_0386;
    114: op1_02_in26 = reg_0963;
    115: op1_02_in26 = reg_0145;
    116: op1_02_in26 = imem05_in[11:8];
    128: op1_02_in26 = imem05_in[11:8];
    117: op1_02_in26 = reg_0144;
    118: op1_02_in26 = reg_0632;
    119: op1_02_in26 = reg_0178;
    120: op1_02_in26 = reg_0717;
    122: op1_02_in26 = reg_0456;
    124: op1_02_in26 = reg_0637;
    125: op1_02_in26 = reg_0756;
    126: op1_02_in26 = reg_0165;
    127: op1_02_in26 = reg_1282;
    43: op1_02_in26 = reg_0196;
    129: op1_02_in26 = reg_1034;
    130: op1_02_in26 = reg_0177;
    131: op1_02_in26 = reg_0239;
    default: op1_02_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv26 = 1;
    53: op1_02_inv26 = 1;
    72: op1_02_inv26 = 1;
    73: op1_02_inv26 = 1;
    59: op1_02_inv26 = 1;
    50: op1_02_inv26 = 1;
    48: op1_02_inv26 = 1;
    74: op1_02_inv26 = 1;
    87: op1_02_inv26 = 1;
    33: op1_02_inv26 = 1;
    76: op1_02_inv26 = 1;
    70: op1_02_inv26 = 1;
    77: op1_02_inv26 = 1;
    58: op1_02_inv26 = 1;
    42: op1_02_inv26 = 1;
    62: op1_02_inv26 = 1;
    89: op1_02_inv26 = 1;
    83: op1_02_inv26 = 1;
    90: op1_02_inv26 = 1;
    94: op1_02_inv26 = 1;
    96: op1_02_inv26 = 1;
    98: op1_02_inv26 = 1;
    99: op1_02_inv26 = 1;
    103: op1_02_inv26 = 1;
    104: op1_02_inv26 = 1;
    105: op1_02_inv26 = 1;
    106: op1_02_inv26 = 1;
    107: op1_02_inv26 = 1;
    111: op1_02_inv26 = 1;
    113: op1_02_inv26 = 1;
    115: op1_02_inv26 = 1;
    117: op1_02_inv26 = 1;
    118: op1_02_inv26 = 1;
    122: op1_02_inv26 = 1;
    126: op1_02_inv26 = 1;
    128: op1_02_inv26 = 1;
    129: op1_02_inv26 = 1;
    default: op1_02_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の27番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in27 = reg_0714;
    53: op1_02_in27 = reg_0114;
    72: op1_02_in27 = reg_0997;
    55: op1_02_in27 = reg_0646;
    73: op1_02_in27 = reg_0584;
    69: op1_02_in27 = reg_0882;
    86: op1_02_in27 = reg_0334;
    59: op1_02_in27 = reg_0047;
    71: op1_02_in27 = reg_0409;
    61: op1_02_in27 = reg_0400;
    50: op1_02_in27 = reg_0576;
    131: op1_02_in27 = reg_0576;
    68: op1_02_in27 = reg_1168;
    48: op1_02_in27 = reg_0622;
    74: op1_02_in27 = reg_0892;
    46: op1_02_in27 = reg_0669;
    75: op1_02_in27 = reg_1003;
    87: op1_02_in27 = reg_1369;
    33: op1_02_in27 = reg_0383;
    60: op1_02_in27 = reg_0940;
    76: op1_02_in27 = reg_0528;
    97: op1_02_in27 = reg_0528;
    57: op1_02_in27 = reg_1064;
    70: op1_02_in27 = reg_0263;
    77: op1_02_in27 = reg_0085;
    44: op1_02_in27 = reg_0822;
    58: op1_02_in27 = reg_0452;
    88: op1_02_in27 = reg_0462;
    78: op1_02_in27 = reg_0127;
    79: op1_02_in27 = reg_0181;
    42: op1_02_in27 = reg_0727;
    80: op1_02_in27 = reg_0228;
    62: op1_02_in27 = reg_0457;
    81: op1_02_in27 = reg_1093;
    89: op1_02_in27 = reg_0342;
    63: op1_02_in27 = reg_0532;
    82: op1_02_in27 = reg_0879;
    83: op1_02_in27 = reg_0371;
    64: op1_02_in27 = reg_0066;
    84: op1_02_in27 = reg_0377;
    85: op1_02_in27 = reg_0484;
    90: op1_02_in27 = reg_0862;
    66: op1_02_in27 = reg_0425;
    91: op1_02_in27 = reg_1097;
    67: op1_02_in27 = reg_0472;
    92: op1_02_in27 = reg_0448;
    93: op1_02_in27 = reg_0158;
    94: op1_02_in27 = imem06_in[7:4];
    95: op1_02_in27 = reg_0802;
    96: op1_02_in27 = reg_0718;
    98: op1_02_in27 = reg_0375;
    99: op1_02_in27 = reg_0042;
    100: op1_02_in27 = reg_0719;
    101: op1_02_in27 = imem03_in[15:12];
    103: op1_02_in27 = reg_1513;
    104: op1_02_in27 = reg_0180;
    105: op1_02_in27 = reg_0828;
    106: op1_02_in27 = reg_1504;
    107: op1_02_in27 = reg_0595;
    108: op1_02_in27 = reg_0463;
    110: op1_02_in27 = reg_0969;
    111: op1_02_in27 = reg_1511;
    112: op1_02_in27 = reg_0792;
    113: op1_02_in27 = reg_0175;
    114: op1_02_in27 = reg_1095;
    115: op1_02_in27 = reg_0143;
    116: op1_02_in27 = reg_0204;
    117: op1_02_in27 = reg_0000;
    118: op1_02_in27 = imem03_in[7:4];
    119: op1_02_in27 = reg_1009;
    120: op1_02_in27 = reg_0374;
    122: op1_02_in27 = reg_0475;
    124: op1_02_in27 = reg_0373;
    125: op1_02_in27 = reg_0962;
    126: op1_02_in27 = reg_1204;
    127: op1_02_in27 = reg_0427;
    43: op1_02_in27 = reg_0240;
    128: op1_02_in27 = reg_0832;
    129: op1_02_in27 = reg_0362;
    130: op1_02_in27 = reg_1033;
    default: op1_02_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_02_inv27 = 1;
    73: op1_02_inv27 = 1;
    71: op1_02_inv27 = 1;
    61: op1_02_inv27 = 1;
    74: op1_02_inv27 = 1;
    75: op1_02_inv27 = 1;
    87: op1_02_inv27 = 1;
    57: op1_02_inv27 = 1;
    77: op1_02_inv27 = 1;
    44: op1_02_inv27 = 1;
    58: op1_02_inv27 = 1;
    78: op1_02_inv27 = 1;
    79: op1_02_inv27 = 1;
    42: op1_02_inv27 = 1;
    80: op1_02_inv27 = 1;
    89: op1_02_inv27 = 1;
    63: op1_02_inv27 = 1;
    84: op1_02_inv27 = 1;
    85: op1_02_inv27 = 1;
    90: op1_02_inv27 = 1;
    67: op1_02_inv27 = 1;
    93: op1_02_inv27 = 1;
    94: op1_02_inv27 = 1;
    95: op1_02_inv27 = 1;
    96: op1_02_inv27 = 1;
    97: op1_02_inv27 = 1;
    98: op1_02_inv27 = 1;
    99: op1_02_inv27 = 1;
    105: op1_02_inv27 = 1;
    106: op1_02_inv27 = 1;
    107: op1_02_inv27 = 1;
    108: op1_02_inv27 = 1;
    111: op1_02_inv27 = 1;
    114: op1_02_inv27 = 1;
    115: op1_02_inv27 = 1;
    117: op1_02_inv27 = 1;
    118: op1_02_inv27 = 1;
    120: op1_02_inv27 = 1;
    122: op1_02_inv27 = 1;
    125: op1_02_inv27 = 1;
    126: op1_02_inv27 = 1;
    127: op1_02_inv27 = 1;
    128: op1_02_inv27 = 1;
    129: op1_02_inv27 = 1;
    131: op1_02_inv27 = 1;
    default: op1_02_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の28番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in28 = reg_0670;
    53: op1_02_in28 = reg_0028;
    72: op1_02_in28 = reg_0561;
    55: op1_02_in28 = reg_0996;
    73: op1_02_in28 = reg_0570;
    76: op1_02_in28 = reg_0570;
    69: op1_02_in28 = reg_0880;
    86: op1_02_in28 = reg_1403;
    59: op1_02_in28 = reg_0093;
    71: op1_02_in28 = reg_0410;
    61: op1_02_in28 = reg_0365;
    50: op1_02_in28 = reg_0966;
    68: op1_02_in28 = reg_0565;
    48: op1_02_in28 = reg_0046;
    74: op1_02_in28 = reg_0851;
    46: op1_02_in28 = reg_0635;
    75: op1_02_in28 = imem03_in[3:0];
    87: op1_02_in28 = reg_0088;
    33: op1_02_in28 = reg_0363;
    103: op1_02_in28 = reg_0363;
    60: op1_02_in28 = reg_0207;
    57: op1_02_in28 = reg_0049;
    70: op1_02_in28 = reg_1367;
    77: op1_02_in28 = reg_0483;
    44: op1_02_in28 = reg_0718;
    58: op1_02_in28 = reg_0304;
    88: op1_02_in28 = reg_1083;
    78: op1_02_in28 = reg_0126;
    79: op1_02_in28 = reg_0978;
    42: op1_02_in28 = reg_0451;
    80: op1_02_in28 = reg_0001;
    62: op1_02_in28 = reg_0742;
    81: op1_02_in28 = reg_1199;
    125: op1_02_in28 = reg_1199;
    89: op1_02_in28 = reg_0368;
    63: op1_02_in28 = reg_0588;
    82: op1_02_in28 = reg_1169;
    83: op1_02_in28 = reg_1179;
    64: op1_02_in28 = reg_1180;
    84: op1_02_in28 = reg_1517;
    90: op1_02_in28 = reg_0339;
    66: op1_02_in28 = reg_0426;
    91: op1_02_in28 = reg_1439;
    67: op1_02_in28 = reg_0326;
    92: op1_02_in28 = reg_0350;
    93: op1_02_in28 = reg_0139;
    94: op1_02_in28 = reg_1105;
    95: op1_02_in28 = reg_0294;
    96: op1_02_in28 = reg_1303;
    97: op1_02_in28 = reg_0345;
    98: op1_02_in28 = reg_1184;
    99: op1_02_in28 = imem02_in[7:4];
    100: op1_02_in28 = reg_0932;
    101: op1_02_in28 = reg_0377;
    104: op1_02_in28 = reg_1494;
    117: op1_02_in28 = reg_1494;
    105: op1_02_in28 = reg_0317;
    106: op1_02_in28 = reg_0717;
    107: op1_02_in28 = reg_0875;
    108: op1_02_in28 = reg_0549;
    110: op1_02_in28 = reg_0033;
    111: op1_02_in28 = reg_1513;
    112: op1_02_in28 = reg_0418;
    113: op1_02_in28 = reg_0400;
    114: op1_02_in28 = reg_1057;
    115: op1_02_in28 = reg_0000;
    130: op1_02_in28 = reg_0000;
    116: op1_02_in28 = reg_0338;
    118: op1_02_in28 = reg_0444;
    119: op1_02_in28 = imem04_in[11:8];
    127: op1_02_in28 = imem04_in[11:8];
    120: op1_02_in28 = reg_0586;
    122: op1_02_in28 = reg_0184;
    124: op1_02_in28 = reg_0624;
    126: op1_02_in28 = reg_0977;
    43: op1_02_in28 = reg_0273;
    128: op1_02_in28 = reg_0833;
    129: op1_02_in28 = reg_0595;
    131: op1_02_in28 = reg_0463;
    default: op1_02_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_02_inv28 = 1;
    55: op1_02_inv28 = 1;
    73: op1_02_inv28 = 1;
    69: op1_02_inv28 = 1;
    59: op1_02_inv28 = 1;
    48: op1_02_inv28 = 1;
    33: op1_02_inv28 = 1;
    76: op1_02_inv28 = 1;
    57: op1_02_inv28 = 1;
    70: op1_02_inv28 = 1;
    77: op1_02_inv28 = 1;
    78: op1_02_inv28 = 1;
    79: op1_02_inv28 = 1;
    89: op1_02_inv28 = 1;
    83: op1_02_inv28 = 1;
    91: op1_02_inv28 = 1;
    92: op1_02_inv28 = 1;
    94: op1_02_inv28 = 1;
    97: op1_02_inv28 = 1;
    98: op1_02_inv28 = 1;
    100: op1_02_inv28 = 1;
    101: op1_02_inv28 = 1;
    103: op1_02_inv28 = 1;
    105: op1_02_inv28 = 1;
    108: op1_02_inv28 = 1;
    111: op1_02_inv28 = 1;
    112: op1_02_inv28 = 1;
    114: op1_02_inv28 = 1;
    115: op1_02_inv28 = 1;
    118: op1_02_inv28 = 1;
    119: op1_02_inv28 = 1;
    120: op1_02_inv28 = 1;
    122: op1_02_inv28 = 1;
    127: op1_02_inv28 = 1;
    130: op1_02_inv28 = 1;
    default: op1_02_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の29番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in29 = reg_0634;
    53: op1_02_in29 = reg_0003;
    72: op1_02_in29 = reg_1344;
    55: op1_02_in29 = reg_0997;
    73: op1_02_in29 = reg_0419;
    69: op1_02_in29 = reg_0247;
    86: op1_02_in29 = reg_1402;
    59: op1_02_in29 = reg_0291;
    71: op1_02_in29 = reg_0405;
    61: op1_02_in29 = reg_0363;
    50: op1_02_in29 = reg_0434;
    68: op1_02_in29 = reg_0697;
    48: op1_02_in29 = reg_0017;
    74: op1_02_in29 = reg_0159;
    46: op1_02_in29 = reg_0637;
    75: op1_02_in29 = reg_0597;
    87: op1_02_in29 = reg_0252;
    33: op1_02_in29 = reg_0093;
    60: op1_02_in29 = reg_0039;
    76: op1_02_in29 = reg_0345;
    57: op1_02_in29 = reg_0348;
    70: op1_02_in29 = reg_1257;
    44: op1_02_in29 = reg_0529;
    58: op1_02_in29 = reg_0338;
    88: op1_02_in29 = reg_0681;
    78: op1_02_in29 = reg_0111;
    79: op1_02_in29 = reg_1215;
    42: op1_02_in29 = reg_0438;
    80: op1_02_in29 = reg_0521;
    62: op1_02_in29 = reg_0532;
    81: op1_02_in29 = reg_1208;
    125: op1_02_in29 = reg_1208;
    89: op1_02_in29 = reg_0719;
    63: op1_02_in29 = reg_0590;
    82: op1_02_in29 = reg_0996;
    83: op1_02_in29 = reg_0023;
    64: op1_02_in29 = reg_0183;
    84: op1_02_in29 = reg_0246;
    90: op1_02_in29 = reg_1237;
    66: op1_02_in29 = reg_0698;
    91: op1_02_in29 = reg_0868;
    67: op1_02_in29 = reg_0973;
    92: op1_02_in29 = reg_1149;
    93: op1_02_in29 = reg_0366;
    94: op1_02_in29 = reg_1030;
    95: op1_02_in29 = reg_0069;
    96: op1_02_in29 = reg_0526;
    97: op1_02_in29 = reg_1179;
    98: op1_02_in29 = reg_1517;
    99: op1_02_in29 = reg_0399;
    100: op1_02_in29 = reg_0209;
    101: op1_02_in29 = reg_0709;
    118: op1_02_in29 = reg_0709;
    103: op1_02_in29 = reg_0899;
    104: op1_02_in29 = reg_1495;
    105: op1_02_in29 = reg_0206;
    106: op1_02_in29 = reg_0714;
    107: op1_02_in29 = reg_0043;
    108: op1_02_in29 = reg_0550;
    110: op1_02_in29 = reg_0232;
    111: op1_02_in29 = reg_0383;
    112: op1_02_in29 = reg_0601;
    113: op1_02_in29 = reg_0162;
    114: op1_02_in29 = reg_0994;
    115: op1_02_in29 = reg_0375;
    116: op1_02_in29 = reg_0466;
    117: op1_02_in29 = reg_0965;
    119: op1_02_in29 = reg_0656;
    120: op1_02_in29 = reg_0584;
    122: op1_02_in29 = reg_1235;
    124: op1_02_in29 = reg_0569;
    126: op1_02_in29 = reg_0152;
    127: op1_02_in29 = reg_1258;
    43: op1_02_in29 = reg_0151;
    128: op1_02_in29 = reg_0890;
    129: op1_02_in29 = reg_0080;
    130: op1_02_in29 = reg_0180;
    131: op1_02_in29 = reg_0163;
    default: op1_02_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    52: op1_02_inv29 = 1;
    53: op1_02_inv29 = 1;
    72: op1_02_inv29 = 1;
    59: op1_02_inv29 = 1;
    71: op1_02_inv29 = 1;
    48: op1_02_inv29 = 1;
    74: op1_02_inv29 = 1;
    33: op1_02_inv29 = 1;
    57: op1_02_inv29 = 1;
    44: op1_02_inv29 = 1;
    79: op1_02_inv29 = 1;
    80: op1_02_inv29 = 1;
    62: op1_02_inv29 = 1;
    81: op1_02_inv29 = 1;
    63: op1_02_inv29 = 1;
    64: op1_02_inv29 = 1;
    84: op1_02_inv29 = 1;
    67: op1_02_inv29 = 1;
    92: op1_02_inv29 = 1;
    93: op1_02_inv29 = 1;
    95: op1_02_inv29 = 1;
    98: op1_02_inv29 = 1;
    99: op1_02_inv29 = 1;
    100: op1_02_inv29 = 1;
    101: op1_02_inv29 = 1;
    103: op1_02_inv29 = 1;
    104: op1_02_inv29 = 1;
    106: op1_02_inv29 = 1;
    107: op1_02_inv29 = 1;
    110: op1_02_inv29 = 1;
    111: op1_02_inv29 = 1;
    114: op1_02_inv29 = 1;
    115: op1_02_inv29 = 1;
    116: op1_02_inv29 = 1;
    122: op1_02_inv29 = 1;
    124: op1_02_inv29 = 1;
    125: op1_02_inv29 = 1;
    126: op1_02_inv29 = 1;
    43: op1_02_inv29 = 1;
    130: op1_02_inv29 = 1;
    default: op1_02_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の30番目の入力
  always @ ( * ) begin
    case ( state )
    52: op1_02_in30 = reg_0584;
    53: op1_02_in30 = reg_0483;
    72: op1_02_in30 = reg_0332;
    55: op1_02_in30 = reg_0992;
    73: op1_02_in30 = reg_0023;
    69: op1_02_in30 = reg_1369;
    86: op1_02_in30 = reg_0939;
    59: op1_02_in30 = reg_0278;
    71: op1_02_in30 = reg_0387;
    61: op1_02_in30 = reg_0047;
    50: op1_02_in30 = reg_0727;
    68: op1_02_in30 = reg_0540;
    48: op1_02_in30 = reg_0162;
    42: op1_02_in30 = reg_0162;
    74: op1_02_in30 = reg_0921;
    46: op1_02_in30 = reg_0261;
    75: op1_02_in30 = reg_1301;
    84: op1_02_in30 = reg_1301;
    87: op1_02_in30 = reg_1215;
    33: op1_02_in30 = reg_0080;
    60: op1_02_in30 = reg_1035;
    76: op1_02_in30 = imem07_in[7:4];
    57: op1_02_in30 = reg_0790;
    70: op1_02_in30 = reg_0978;
    44: op1_02_in30 = reg_0527;
    58: op1_02_in30 = reg_0019;
    88: op1_02_in30 = reg_1082;
    78: op1_02_in30 = reg_0824;
    79: op1_02_in30 = reg_1200;
    80: op1_02_in30 = reg_0520;
    62: op1_02_in30 = reg_0253;
    81: op1_02_in30 = reg_0104;
    89: op1_02_in30 = reg_0336;
    63: op1_02_in30 = reg_0589;
    82: op1_02_in30 = reg_0174;
    83: op1_02_in30 = reg_0022;
    64: op1_02_in30 = reg_0418;
    90: op1_02_in30 = reg_0211;
    66: op1_02_in30 = reg_0582;
    91: op1_02_in30 = reg_0786;
    67: op1_02_in30 = reg_0126;
    92: op1_02_in30 = reg_0707;
    93: op1_02_in30 = reg_0213;
    94: op1_02_in30 = reg_1467;
    95: op1_02_in30 = reg_0279;
    96: op1_02_in30 = reg_0528;
    97: op1_02_in30 = reg_0270;
    98: op1_02_in30 = reg_0329;
    99: op1_02_in30 = reg_1018;
    100: op1_02_in30 = imem05_in[7:4];
    101: op1_02_in30 = reg_0823;
    103: op1_02_in30 = reg_0899;
    104: op1_02_in30 = reg_0954;
    105: op1_02_in30 = imem06_in[15:12];
    106: op1_02_in30 = reg_0398;
    107: op1_02_in30 = reg_0895;
    108: op1_02_in30 = reg_1474;
    110: op1_02_in30 = reg_0698;
    111: op1_02_in30 = reg_0363;
    112: op1_02_in30 = reg_0274;
    113: op1_02_in30 = reg_0402;
    114: op1_02_in30 = reg_0140;
    115: op1_02_in30 = reg_1495;
    130: op1_02_in30 = reg_1495;
    116: op1_02_in30 = reg_0333;
    117: op1_02_in30 = reg_0142;
    118: op1_02_in30 = reg_1000;
    119: op1_02_in30 = reg_0340;
    120: op1_02_in30 = reg_0619;
    122: op1_02_in30 = reg_0879;
    124: op1_02_in30 = reg_0132;
    125: op1_02_in30 = reg_0107;
    126: op1_02_in30 = reg_0214;
    127: op1_02_in30 = reg_0574;
    43: op1_02_in30 = reg_0204;
    128: op1_02_in30 = reg_0040;
    129: op1_02_in30 = reg_0896;
    131: op1_02_in30 = reg_0331;
    default: op1_02_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_02_inv30 = 1;
    55: op1_02_inv30 = 1;
    69: op1_02_inv30 = 1;
    86: op1_02_inv30 = 1;
    59: op1_02_inv30 = 1;
    71: op1_02_inv30 = 1;
    68: op1_02_inv30 = 1;
    74: op1_02_inv30 = 1;
    75: op1_02_inv30 = 1;
    87: op1_02_inv30 = 1;
    33: op1_02_inv30 = 1;
    60: op1_02_inv30 = 1;
    76: op1_02_inv30 = 1;
    44: op1_02_inv30 = 1;
    88: op1_02_inv30 = 1;
    78: op1_02_inv30 = 1;
    79: op1_02_inv30 = 1;
    81: op1_02_inv30 = 1;
    63: op1_02_inv30 = 1;
    82: op1_02_inv30 = 1;
    83: op1_02_inv30 = 1;
    64: op1_02_inv30 = 1;
    84: op1_02_inv30 = 1;
    91: op1_02_inv30 = 1;
    67: op1_02_inv30 = 1;
    92: op1_02_inv30 = 1;
    99: op1_02_inv30 = 1;
    101: op1_02_inv30 = 1;
    103: op1_02_inv30 = 1;
    104: op1_02_inv30 = 1;
    105: op1_02_inv30 = 1;
    106: op1_02_inv30 = 1;
    110: op1_02_inv30 = 1;
    112: op1_02_inv30 = 1;
    114: op1_02_inv30 = 1;
    115: op1_02_inv30 = 1;
    116: op1_02_inv30 = 1;
    118: op1_02_inv30 = 1;
    119: op1_02_inv30 = 1;
    120: op1_02_inv30 = 1;
    122: op1_02_inv30 = 1;
    43: op1_02_inv30 = 1;
    128: op1_02_inv30 = 1;
    default: op1_02_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_02_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#2の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_02_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の0番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in00 = reg_0451;
    42: op1_03_in00 = reg_0451;
    72: op1_03_in00 = reg_0565;
    55: op1_03_in00 = reg_0295;
    73: op1_03_in00 = reg_0937;
    86: op1_03_in00 = reg_0185;
    49: op1_03_in00 = reg_0716;
    69: op1_03_in00 = reg_0055;
    61: op1_03_in00 = reg_0554;
    54: op1_03_in00 = reg_0285;
    71: op1_03_in00 = reg_0748;
    50: op1_03_in00 = reg_0253;
    68: op1_03_in00 = reg_0113;
    48: op1_03_in00 = reg_0902;
    52: op1_03_in00 = imem00_in[7:4];
    92: op1_03_in00 = imem00_in[7:4];
    109: op1_03_in00 = imem00_in[7:4];
    123: op1_03_in00 = imem00_in[7:4];
    74: op1_03_in00 = reg_0066;
    75: op1_03_in00 = reg_0540;
    87: op1_03_in00 = reg_0497;
    56: op1_03_in00 = reg_0022;
    46: op1_03_in00 = reg_0012;
    60: op1_03_in00 = reg_0313;
    76: op1_03_in00 = reg_1509;
    59: op1_03_in00 = reg_0219;
    33: op1_03_in00 = reg_0366;
    57: op1_03_in00 = reg_0332;
    77: op1_03_in00 = imem00_in[3:0];
    81: op1_03_in00 = imem00_in[3:0];
    93: op1_03_in00 = imem00_in[3:0];
    114: op1_03_in00 = imem00_in[3:0];
    121: op1_03_in00 = imem00_in[3:0];
    70: op1_03_in00 = imem01_in[11:8];
    58: op1_03_in00 = reg_0718;
    44: op1_03_in00 = reg_0799;
    78: op1_03_in00 = reg_0701;
    88: op1_03_in00 = reg_0104;
    51: op1_03_in00 = reg_0043;
    28: op1_03_in00 = reg_0001;
    79: op1_03_in00 = reg_1277;
    22: op1_03_in00 = imem07_in[11:8];
    4: op1_03_in00 = imem07_in[11:8];
    37: op1_03_in00 = reg_0139;
    80: op1_03_in00 = reg_0395;
    62: op1_03_in00 = reg_0042;
    34: op1_03_in00 = imem07_in[7:4];
    47: op1_03_in00 = reg_0371;
    89: op1_03_in00 = imem02_in[7:4];
    63: op1_03_in00 = reg_0152;
    97: op1_03_in00 = reg_0152;
    82: op1_03_in00 = reg_0182;
    83: op1_03_in00 = reg_0698;
    64: op1_03_in00 = reg_0899;
    40: op1_03_in00 = reg_0603;
    84: op1_03_in00 = reg_0604;
    65: op1_03_in00 = reg_0559;
    85: op1_03_in00 = reg_0791;
    90: op1_03_in00 = reg_0312;
    66: op1_03_in00 = reg_1346;
    91: op1_03_in00 = reg_0725;
    67: op1_03_in00 = reg_0569;
    94: op1_03_in00 = reg_0720;
    95: op1_03_in00 = imem03_in[11:8];
    96: op1_03_in00 = reg_0570;
    98: op1_03_in00 = reg_1301;
    99: op1_03_in00 = reg_0138;
    100: op1_03_in00 = imem05_in[11:8];
    101: op1_03_in00 = reg_0143;
    102: op1_03_in00 = imem00_in[11:8];
    103: op1_03_in00 = reg_0092;
    104: op1_03_in00 = reg_0048;
    105: op1_03_in00 = reg_0931;
    106: op1_03_in00 = reg_0141;
    107: op1_03_in00 = reg_0447;
    108: op1_03_in00 = reg_0572;
    110: op1_03_in00 = reg_0582;
    111: op1_03_in00 = reg_0595;
    38: op1_03_in00 = reg_0299;
    112: op1_03_in00 = reg_0575;
    113: op1_03_in00 = imem02_in[15:12];
    115: op1_03_in00 = reg_0965;
    116: op1_03_in00 = reg_0184;
    117: op1_03_in00 = reg_0954;
    118: op1_03_in00 = reg_1425;
    119: op1_03_in00 = reg_0129;
    120: op1_03_in00 = reg_0527;
    29: op1_03_in00 = reg_0137;
    122: op1_03_in00 = reg_0276;
    124: op1_03_in00 = reg_1204;
    125: op1_03_in00 = reg_0880;
    126: op1_03_in00 = reg_0213;
    127: op1_03_in00 = imem05_in[3:0];
    128: op1_03_in00 = reg_0996;
    129: op1_03_in00 = reg_0403;
    130: op1_03_in00 = reg_0556;
    43: op1_03_in00 = reg_0330;
    131: op1_03_in00 = reg_0550;
    default: op1_03_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv00 = 1;
    86: op1_03_inv00 = 1;
    50: op1_03_inv00 = 1;
    74: op1_03_inv00 = 1;
    46: op1_03_inv00 = 1;
    60: op1_03_inv00 = 1;
    76: op1_03_inv00 = 1;
    59: op1_03_inv00 = 1;
    77: op1_03_inv00 = 1;
    70: op1_03_inv00 = 1;
    58: op1_03_inv00 = 1;
    88: op1_03_inv00 = 1;
    51: op1_03_inv00 = 1;
    22: op1_03_inv00 = 1;
    37: op1_03_inv00 = 1;
    80: op1_03_inv00 = 1;
    42: op1_03_inv00 = 1;
    82: op1_03_inv00 = 1;
    83: op1_03_inv00 = 1;
    40: op1_03_inv00 = 1;
    84: op1_03_inv00 = 1;
    65: op1_03_inv00 = 1;
    85: op1_03_inv00 = 1;
    92: op1_03_inv00 = 1;
    97: op1_03_inv00 = 1;
    98: op1_03_inv00 = 1;
    100: op1_03_inv00 = 1;
    102: op1_03_inv00 = 1;
    104: op1_03_inv00 = 1;
    105: op1_03_inv00 = 1;
    106: op1_03_inv00 = 1;
    108: op1_03_inv00 = 1;
    38: op1_03_inv00 = 1;
    112: op1_03_inv00 = 1;
    113: op1_03_inv00 = 1;
    115: op1_03_inv00 = 1;
    118: op1_03_inv00 = 1;
    121: op1_03_inv00 = 1;
    125: op1_03_inv00 = 1;
    127: op1_03_inv00 = 1;
    129: op1_03_inv00 = 1;
    130: op1_03_inv00 = 1;
    43: op1_03_inv00 = 1;
    default: op1_03_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の1番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in01 = reg_0904;
    72: op1_03_in01 = reg_0566;
    55: op1_03_in01 = reg_0171;
    73: op1_03_in01 = reg_0070;
    86: op1_03_in01 = reg_0154;
    49: op1_03_in01 = reg_0670;
    69: op1_03_in01 = reg_0876;
    61: op1_03_in01 = reg_0616;
    81: op1_03_in01 = reg_0616;
    54: op1_03_in01 = reg_0741;
    71: op1_03_in01 = reg_0824;
    50: op1_03_in01 = reg_0530;
    68: op1_03_in01 = reg_0880;
    48: op1_03_in01 = reg_0013;
    46: op1_03_in01 = reg_0013;
    62: op1_03_in01 = reg_0013;
    52: op1_03_in01 = imem00_in[11:8];
    74: op1_03_in01 = reg_0541;
    75: op1_03_in01 = reg_0541;
    87: op1_03_in01 = reg_0390;
    99: op1_03_in01 = reg_0390;
    56: op1_03_in01 = reg_1183;
    60: op1_03_in01 = reg_0525;
    76: op1_03_in01 = reg_0264;
    59: op1_03_in01 = reg_1101;
    33: op1_03_in01 = imem07_in[7:4];
    57: op1_03_in01 = reg_0736;
    77: op1_03_in01 = reg_1079;
    70: op1_03_in01 = reg_0147;
    58: op1_03_in01 = reg_0636;
    44: op1_03_in01 = reg_0578;
    78: op1_03_in01 = reg_0640;
    88: op1_03_in01 = reg_0448;
    51: op1_03_in01 = imem02_in[3:0];
    129: op1_03_in01 = imem02_in[3:0];
    28: op1_03_in01 = imem07_in[3:0];
    79: op1_03_in01 = reg_1490;
    37: op1_03_in01 = reg_0663;
    80: op1_03_in01 = reg_0347;
    34: op1_03_in01 = reg_0284;
    42: op1_03_in01 = reg_0439;
    47: op1_03_in01 = reg_0110;
    89: op1_03_in01 = reg_0472;
    63: op1_03_in01 = reg_0214;
    82: op1_03_in01 = reg_0564;
    83: op1_03_in01 = reg_0236;
    64: op1_03_in01 = reg_0292;
    111: op1_03_in01 = reg_0292;
    40: op1_03_in01 = reg_0567;
    84: op1_03_in01 = reg_0391;
    65: op1_03_in01 = reg_0964;
    85: op1_03_in01 = reg_0866;
    90: op1_03_in01 = reg_1184;
    115: op1_03_in01 = reg_1184;
    66: op1_03_in01 = reg_0151;
    91: op1_03_in01 = reg_0638;
    67: op1_03_in01 = reg_1225;
    92: op1_03_in01 = imem00_in[15:12];
    93: op1_03_in01 = imem00_in[7:4];
    114: op1_03_in01 = imem00_in[7:4];
    94: op1_03_in01 = reg_1505;
    95: op1_03_in01 = reg_0506;
    96: op1_03_in01 = reg_0979;
    97: op1_03_in01 = reg_0022;
    98: op1_03_in01 = reg_0558;
    100: op1_03_in01 = reg_1059;
    101: op1_03_in01 = reg_0234;
    102: op1_03_in01 = reg_1278;
    103: op1_03_in01 = reg_0595;
    104: op1_03_in01 = reg_1325;
    105: op1_03_in01 = reg_1467;
    106: op1_03_in01 = reg_0373;
    107: op1_03_in01 = reg_0889;
    113: op1_03_in01 = reg_0889;
    108: op1_03_in01 = reg_1456;
    109: op1_03_in01 = reg_1243;
    110: op1_03_in01 = reg_0268;
    38: op1_03_in01 = reg_0672;
    112: op1_03_in01 = reg_1346;
    116: op1_03_in01 = reg_0996;
    117: op1_03_in01 = reg_0505;
    118: op1_03_in01 = reg_1001;
    119: op1_03_in01 = reg_1367;
    120: op1_03_in01 = reg_0568;
    121: op1_03_in01 = reg_0983;
    29: op1_03_in01 = reg_0413;
    122: op1_03_in01 = reg_0254;
    123: op1_03_in01 = reg_1099;
    124: op1_03_in01 = reg_0195;
    125: op1_03_in01 = reg_0291;
    126: op1_03_in01 = reg_0018;
    127: op1_03_in01 = reg_0575;
    128: op1_03_in01 = reg_0992;
    130: op1_03_in01 = reg_1517;
    43: op1_03_in01 = reg_0582;
    131: op1_03_in01 = reg_0610;
    default: op1_03_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv01 = 1;
    86: op1_03_inv01 = 1;
    69: op1_03_inv01 = 1;
    61: op1_03_inv01 = 1;
    54: op1_03_inv01 = 1;
    71: op1_03_inv01 = 1;
    68: op1_03_inv01 = 1;
    48: op1_03_inv01 = 1;
    52: op1_03_inv01 = 1;
    56: op1_03_inv01 = 1;
    46: op1_03_inv01 = 1;
    70: op1_03_inv01 = 1;
    44: op1_03_inv01 = 1;
    78: op1_03_inv01 = 1;
    51: op1_03_inv01 = 1;
    79: op1_03_inv01 = 1;
    80: op1_03_inv01 = 1;
    62: op1_03_inv01 = 1;
    63: op1_03_inv01 = 1;
    64: op1_03_inv01 = 1;
    40: op1_03_inv01 = 1;
    85: op1_03_inv01 = 1;
    66: op1_03_inv01 = 1;
    92: op1_03_inv01 = 1;
    93: op1_03_inv01 = 1;
    95: op1_03_inv01 = 1;
    96: op1_03_inv01 = 1;
    97: op1_03_inv01 = 1;
    99: op1_03_inv01 = 1;
    101: op1_03_inv01 = 1;
    103: op1_03_inv01 = 1;
    105: op1_03_inv01 = 1;
    107: op1_03_inv01 = 1;
    108: op1_03_inv01 = 1;
    109: op1_03_inv01 = 1;
    110: op1_03_inv01 = 1;
    38: op1_03_inv01 = 1;
    112: op1_03_inv01 = 1;
    115: op1_03_inv01 = 1;
    116: op1_03_inv01 = 1;
    117: op1_03_inv01 = 1;
    121: op1_03_inv01 = 1;
    122: op1_03_inv01 = 1;
    125: op1_03_inv01 = 1;
    126: op1_03_inv01 = 1;
    129: op1_03_inv01 = 1;
    130: op1_03_inv01 = 1;
    43: op1_03_inv01 = 1;
    131: op1_03_inv01 = 1;
    default: op1_03_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の2番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in02 = reg_0304;
    72: op1_03_in02 = reg_1403;
    55: op1_03_in02 = reg_0419;
    73: op1_03_in02 = reg_0197;
    86: op1_03_in02 = reg_0706;
    49: op1_03_in02 = reg_0583;
    69: op1_03_in02 = reg_0878;
    61: op1_03_in02 = reg_0615;
    102: op1_03_in02 = reg_0615;
    54: op1_03_in02 = reg_0593;
    71: op1_03_in02 = reg_0791;
    50: op1_03_in02 = reg_0981;
    68: op1_03_in02 = reg_0884;
    48: op1_03_in02 = reg_0662;
    52: op1_03_in02 = reg_0581;
    74: op1_03_in02 = imem05_in[11:8];
    75: op1_03_in02 = reg_0939;
    87: op1_03_in02 = reg_0475;
    56: op1_03_in02 = reg_0893;
    46: op1_03_in02 = reg_0628;
    60: op1_03_in02 = reg_0556;
    76: op1_03_in02 = reg_1326;
    59: op1_03_in02 = reg_1102;
    33: op1_03_in02 = imem07_in[15:12];
    97: op1_03_in02 = imem07_in[15:12];
    57: op1_03_in02 = reg_0737;
    77: op1_03_in02 = reg_1490;
    91: op1_03_in02 = reg_1490;
    70: op1_03_in02 = reg_0386;
    58: op1_03_in02 = reg_0637;
    44: op1_03_in02 = reg_0393;
    78: op1_03_in02 = reg_1278;
    88: op1_03_in02 = reg_0481;
    51: op1_03_in02 = imem02_in[15:12];
    79: op1_03_in02 = reg_0841;
    37: op1_03_in02 = imem07_in[11:8];
    80: op1_03_in02 = reg_0346;
    62: op1_03_in02 = reg_0699;
    34: op1_03_in02 = reg_0285;
    42: op1_03_in02 = reg_0161;
    47: op1_03_in02 = reg_0524;
    81: op1_03_in02 = reg_1281;
    89: op1_03_in02 = reg_0432;
    63: op1_03_in02 = reg_0491;
    82: op1_03_in02 = reg_1402;
    83: op1_03_in02 = reg_0904;
    64: op1_03_in02 = reg_0277;
    40: op1_03_in02 = reg_0066;
    84: op1_03_in02 = reg_0334;
    65: op1_03_in02 = reg_1314;
    90: op1_03_in02 = reg_1314;
    85: op1_03_in02 = reg_0616;
    66: op1_03_in02 = reg_0828;
    67: op1_03_in02 = reg_0171;
    92: op1_03_in02 = reg_1243;
    93: op1_03_in02 = reg_0638;
    94: op1_03_in02 = reg_0172;
    95: op1_03_in02 = reg_0559;
    96: op1_03_in02 = reg_0296;
    98: op1_03_in02 = reg_1199;
    99: op1_03_in02 = reg_0433;
    100: op1_03_in02 = reg_1431;
    101: op1_03_in02 = reg_0142;
    103: op1_03_in02 = reg_0335;
    104: op1_03_in02 = reg_0426;
    105: op1_03_in02 = reg_0720;
    106: op1_03_in02 = reg_0624;
    107: op1_03_in02 = reg_0607;
    108: op1_03_in02 = reg_0147;
    109: op1_03_in02 = reg_1277;
    110: op1_03_in02 = reg_0487;
    111: op1_03_in02 = reg_0080;
    38: op1_03_in02 = reg_0661;
    112: op1_03_in02 = reg_0799;
    113: op1_03_in02 = reg_0721;
    114: op1_03_in02 = reg_1242;
    115: op1_03_in02 = reg_1516;
    116: op1_03_in02 = reg_0831;
    117: op1_03_in02 = reg_1301;
    118: op1_03_in02 = reg_0311;
    119: op1_03_in02 = reg_0264;
    120: op1_03_in02 = reg_0345;
    121: op1_03_in02 = reg_1081;
    29: op1_03_in02 = reg_0123;
    122: op1_03_in02 = reg_0839;
    123: op1_03_in02 = reg_1141;
    124: op1_03_in02 = reg_0152;
    125: op1_03_in02 = reg_0313;
    126: op1_03_in02 = imem07_in[3:0];
    127: op1_03_in02 = reg_0206;
    128: op1_03_in02 = reg_0793;
    129: op1_03_in02 = imem02_in[11:8];
    130: op1_03_in02 = reg_0627;
    43: op1_03_in02 = reg_0471;
    131: op1_03_in02 = reg_0222;
    default: op1_03_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv02 = 1;
    55: op1_03_inv02 = 1;
    73: op1_03_inv02 = 1;
    54: op1_03_inv02 = 1;
    71: op1_03_inv02 = 1;
    50: op1_03_inv02 = 1;
    48: op1_03_inv02 = 1;
    52: op1_03_inv02 = 1;
    75: op1_03_inv02 = 1;
    60: op1_03_inv02 = 1;
    76: op1_03_inv02 = 1;
    77: op1_03_inv02 = 1;
    44: op1_03_inv02 = 1;
    78: op1_03_inv02 = 1;
    88: op1_03_inv02 = 1;
    51: op1_03_inv02 = 1;
    79: op1_03_inv02 = 1;
    37: op1_03_inv02 = 1;
    80: op1_03_inv02 = 1;
    62: op1_03_inv02 = 1;
    42: op1_03_inv02 = 1;
    47: op1_03_inv02 = 1;
    89: op1_03_inv02 = 1;
    63: op1_03_inv02 = 1;
    83: op1_03_inv02 = 1;
    64: op1_03_inv02 = 1;
    40: op1_03_inv02 = 1;
    84: op1_03_inv02 = 1;
    65: op1_03_inv02 = 1;
    66: op1_03_inv02 = 1;
    67: op1_03_inv02 = 1;
    94: op1_03_inv02 = 1;
    96: op1_03_inv02 = 1;
    100: op1_03_inv02 = 1;
    101: op1_03_inv02 = 1;
    102: op1_03_inv02 = 1;
    104: op1_03_inv02 = 1;
    106: op1_03_inv02 = 1;
    107: op1_03_inv02 = 1;
    109: op1_03_inv02 = 1;
    111: op1_03_inv02 = 1;
    38: op1_03_inv02 = 1;
    112: op1_03_inv02 = 1;
    114: op1_03_inv02 = 1;
    116: op1_03_inv02 = 1;
    118: op1_03_inv02 = 1;
    119: op1_03_inv02 = 1;
    121: op1_03_inv02 = 1;
    29: op1_03_inv02 = 1;
    125: op1_03_inv02 = 1;
    127: op1_03_inv02 = 1;
    131: op1_03_inv02 = 1;
    default: op1_03_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の3番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in03 = reg_0837;
    72: op1_03_in03 = reg_0538;
    55: op1_03_in03 = reg_0308;
    73: op1_03_in03 = reg_0274;
    86: op1_03_in03 = reg_0847;
    49: op1_03_in03 = reg_0244;
    67: op1_03_in03 = reg_0244;
    69: op1_03_in03 = reg_0381;
    61: op1_03_in03 = reg_0614;
    54: op1_03_in03 = reg_0591;
    71: op1_03_in03 = reg_1079;
    50: op1_03_in03 = reg_0991;
    68: op1_03_in03 = reg_0504;
    48: op1_03_in03 = reg_0553;
    52: op1_03_in03 = reg_1100;
    74: op1_03_in03 = reg_0576;
    75: op1_03_in03 = reg_0301;
    87: op1_03_in03 = reg_0971;
    56: op1_03_in03 = reg_0310;
    46: op1_03_in03 = reg_0631;
    60: op1_03_in03 = reg_0707;
    76: op1_03_in03 = reg_1334;
    59: op1_03_in03 = imem00_in[7:4];
    33: op1_03_in03 = reg_0361;
    57: op1_03_in03 = reg_0702;
    77: op1_03_in03 = reg_0350;
    70: op1_03_in03 = reg_0290;
    58: op1_03_in03 = imem06_in[3:0];
    44: op1_03_in03 = reg_0344;
    78: op1_03_in03 = reg_1279;
    109: op1_03_in03 = reg_1279;
    88: op1_03_in03 = reg_0025;
    51: op1_03_in03 = reg_0588;
    79: op1_03_in03 = reg_0615;
    37: op1_03_in03 = imem07_in[15:12];
    126: op1_03_in03 = imem07_in[15:12];
    80: op1_03_in03 = reg_0646;
    62: op1_03_in03 = reg_0632;
    34: op1_03_in03 = reg_0442;
    42: op1_03_in03 = reg_0146;
    47: op1_03_in03 = reg_0636;
    81: op1_03_in03 = reg_1081;
    89: op1_03_in03 = reg_0436;
    63: op1_03_in03 = reg_1057;
    82: op1_03_in03 = reg_1404;
    83: op1_03_in03 = reg_0065;
    64: op1_03_in03 = reg_0699;
    40: op1_03_in03 = reg_0045;
    84: op1_03_in03 = reg_1180;
    65: op1_03_in03 = reg_0627;
    85: op1_03_in03 = reg_0907;
    90: op1_03_in03 = reg_0957;
    130: op1_03_in03 = reg_0957;
    66: op1_03_in03 = reg_0317;
    91: op1_03_in03 = reg_0580;
    92: op1_03_in03 = reg_0613;
    123: op1_03_in03 = reg_0613;
    93: op1_03_in03 = reg_1281;
    94: op1_03_in03 = reg_0110;
    95: op1_03_in03 = reg_0179;
    96: op1_03_in03 = reg_0295;
    97: op1_03_in03 = reg_1055;
    98: op1_03_in03 = reg_0107;
    99: op1_03_in03 = reg_0326;
    100: op1_03_in03 = reg_0184;
    101: op1_03_in03 = reg_1517;
    102: op1_03_in03 = reg_0805;
    103: op1_03_in03 = reg_0162;
    104: op1_03_in03 = reg_0411;
    105: op1_03_in03 = reg_0827;
    106: op1_03_in03 = reg_0570;
    107: op1_03_in03 = reg_0169;
    108: op1_03_in03 = reg_0148;
    110: op1_03_in03 = reg_0236;
    111: op1_03_in03 = reg_0634;
    38: op1_03_in03 = reg_0287;
    112: op1_03_in03 = reg_0864;
    113: op1_03_in03 = reg_1002;
    114: op1_03_in03 = reg_0581;
    115: op1_03_in03 = reg_0329;
    116: op1_03_in03 = reg_0648;
    117: op1_03_in03 = reg_0880;
    118: op1_03_in03 = reg_0191;
    119: op1_03_in03 = reg_0034;
    120: op1_03_in03 = reg_0419;
    121: op1_03_in03 = reg_0638;
    122: op1_03_in03 = reg_0744;
    124: op1_03_in03 = reg_0212;
    125: op1_03_in03 = reg_0790;
    127: op1_03_in03 = reg_0039;
    128: op1_03_in03 = reg_0604;
    129: op1_03_in03 = imem02_in[15:12];
    43: op1_03_in03 = reg_0454;
    131: op1_03_in03 = reg_0743;
    default: op1_03_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv03 = 1;
    73: op1_03_inv03 = 1;
    86: op1_03_inv03 = 1;
    49: op1_03_inv03 = 1;
    69: op1_03_inv03 = 1;
    61: op1_03_inv03 = 1;
    74: op1_03_inv03 = 1;
    75: op1_03_inv03 = 1;
    46: op1_03_inv03 = 1;
    76: op1_03_inv03 = 1;
    33: op1_03_inv03 = 1;
    57: op1_03_inv03 = 1;
    58: op1_03_inv03 = 1;
    88: op1_03_inv03 = 1;
    51: op1_03_inv03 = 1;
    80: op1_03_inv03 = 1;
    34: op1_03_inv03 = 1;
    47: op1_03_inv03 = 1;
    63: op1_03_inv03 = 1;
    82: op1_03_inv03 = 1;
    83: op1_03_inv03 = 1;
    64: op1_03_inv03 = 1;
    40: op1_03_inv03 = 1;
    84: op1_03_inv03 = 1;
    65: op1_03_inv03 = 1;
    66: op1_03_inv03 = 1;
    93: op1_03_inv03 = 1;
    95: op1_03_inv03 = 1;
    98: op1_03_inv03 = 1;
    99: op1_03_inv03 = 1;
    100: op1_03_inv03 = 1;
    101: op1_03_inv03 = 1;
    106: op1_03_inv03 = 1;
    109: op1_03_inv03 = 1;
    110: op1_03_inv03 = 1;
    38: op1_03_inv03 = 1;
    113: op1_03_inv03 = 1;
    114: op1_03_inv03 = 1;
    115: op1_03_inv03 = 1;
    116: op1_03_inv03 = 1;
    117: op1_03_inv03 = 1;
    121: op1_03_inv03 = 1;
    124: op1_03_inv03 = 1;
    128: op1_03_inv03 = 1;
    130: op1_03_inv03 = 1;
    43: op1_03_inv03 = 1;
    131: op1_03_inv03 = 1;
    default: op1_03_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の4番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in04 = reg_0338;
    72: op1_03_in04 = reg_0450;
    55: op1_03_in04 = imem06_in[7:4];
    73: op1_03_in04 = reg_0118;
    86: op1_03_in04 = reg_0823;
    49: op1_03_in04 = reg_0490;
    69: op1_03_in04 = reg_0705;
    61: op1_03_in04 = reg_0748;
    54: op1_03_in04 = reg_0103;
    71: op1_03_in04 = reg_0842;
    50: op1_03_in04 = reg_0326;
    89: op1_03_in04 = reg_0326;
    68: op1_03_in04 = reg_0479;
    48: op1_03_in04 = reg_0256;
    52: op1_03_in04 = reg_0843;
    74: op1_03_in04 = reg_0492;
    75: op1_03_in04 = reg_0274;
    87: op1_03_in04 = reg_0127;
    56: op1_03_in04 = reg_0186;
    46: op1_03_in04 = reg_0531;
    60: op1_03_in04 = reg_0706;
    76: op1_03_in04 = reg_0869;
    59: op1_03_in04 = reg_1079;
    78: op1_03_in04 = reg_1079;
    93: op1_03_in04 = reg_1079;
    33: op1_03_in04 = reg_0053;
    57: op1_03_in04 = reg_1168;
    77: op1_03_in04 = reg_0121;
    70: op1_03_in04 = reg_0606;
    58: op1_03_in04 = reg_0619;
    44: op1_03_in04 = reg_0702;
    88: op1_03_in04 = reg_0291;
    51: op1_03_in04 = reg_0590;
    79: op1_03_in04 = reg_0580;
    37: op1_03_in04 = reg_0404;
    80: op1_03_in04 = reg_0649;
    62: op1_03_in04 = reg_0608;
    34: op1_03_in04 = reg_0618;
    42: op1_03_in04 = reg_0400;
    47: op1_03_in04 = reg_0624;
    81: op1_03_in04 = reg_1487;
    63: op1_03_in04 = reg_1055;
    82: op1_03_in04 = reg_0940;
    83: op1_03_in04 = reg_0420;
    64: op1_03_in04 = imem02_in[7:4];
    40: op1_03_in04 = reg_0131;
    84: op1_03_in04 = reg_1403;
    65: op1_03_in04 = reg_0957;
    85: op1_03_in04 = reg_0672;
    90: op1_03_in04 = reg_0952;
    66: op1_03_in04 = reg_0040;
    112: op1_03_in04 = reg_0040;
    91: op1_03_in04 = reg_0555;
    67: op1_03_in04 = reg_1202;
    96: op1_03_in04 = reg_1202;
    92: op1_03_in04 = reg_0616;
    94: op1_03_in04 = reg_0109;
    95: op1_03_in04 = reg_0330;
    97: op1_03_in04 = reg_0219;
    98: op1_03_in04 = reg_0350;
    99: op1_03_in04 = reg_0970;
    100: op1_03_in04 = reg_0272;
    101: op1_03_in04 = reg_0627;
    102: op1_03_in04 = reg_0523;
    103: op1_03_in04 = reg_0402;
    104: op1_03_in04 = imem04_in[7:4];
    105: op1_03_in04 = reg_1501;
    106: op1_03_in04 = reg_1225;
    107: op1_03_in04 = reg_0399;
    108: op1_03_in04 = reg_1511;
    109: op1_03_in04 = reg_0153;
    110: op1_03_in04 = reg_0904;
    111: op1_03_in04 = reg_0012;
    38: op1_03_in04 = reg_0366;
    113: op1_03_in04 = reg_1235;
    114: op1_03_in04 = reg_0958;
    115: op1_03_in04 = reg_1199;
    116: op1_03_in04 = reg_0604;
    117: op1_03_in04 = reg_0313;
    118: op1_03_in04 = reg_1184;
    119: op1_03_in04 = reg_0694;
    120: op1_03_in04 = reg_0152;
    121: op1_03_in04 = reg_1278;
    122: op1_03_in04 = reg_0822;
    123: op1_03_in04 = reg_0841;
    124: op1_03_in04 = imem07_in[7:4];
    125: op1_03_in04 = reg_0425;
    126: op1_03_in04 = reg_0169;
    127: op1_03_in04 = reg_1299;
    128: op1_03_in04 = reg_0045;
    129: op1_03_in04 = reg_0495;
    130: op1_03_in04 = reg_0505;
    43: op1_03_in04 = reg_0699;
    131: op1_03_in04 = reg_0609;
    default: op1_03_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv04 = 1;
    55: op1_03_inv04 = 1;
    50: op1_03_inv04 = 1;
    48: op1_03_inv04 = 1;
    74: op1_03_inv04 = 1;
    75: op1_03_inv04 = 1;
    56: op1_03_inv04 = 1;
    60: op1_03_inv04 = 1;
    76: op1_03_inv04 = 1;
    33: op1_03_inv04 = 1;
    70: op1_03_inv04 = 1;
    58: op1_03_inv04 = 1;
    78: op1_03_inv04 = 1;
    37: op1_03_inv04 = 1;
    80: op1_03_inv04 = 1;
    34: op1_03_inv04 = 1;
    42: op1_03_inv04 = 1;
    81: op1_03_inv04 = 1;
    63: op1_03_inv04 = 1;
    64: op1_03_inv04 = 1;
    84: op1_03_inv04 = 1;
    65: op1_03_inv04 = 1;
    85: op1_03_inv04 = 1;
    90: op1_03_inv04 = 1;
    67: op1_03_inv04 = 1;
    92: op1_03_inv04 = 1;
    93: op1_03_inv04 = 1;
    94: op1_03_inv04 = 1;
    96: op1_03_inv04 = 1;
    97: op1_03_inv04 = 1;
    98: op1_03_inv04 = 1;
    100: op1_03_inv04 = 1;
    101: op1_03_inv04 = 1;
    105: op1_03_inv04 = 1;
    109: op1_03_inv04 = 1;
    114: op1_03_inv04 = 1;
    119: op1_03_inv04 = 1;
    120: op1_03_inv04 = 1;
    121: op1_03_inv04 = 1;
    123: op1_03_inv04 = 1;
    126: op1_03_inv04 = 1;
    127: op1_03_inv04 = 1;
    130: op1_03_inv04 = 1;
    131: op1_03_inv04 = 1;
    default: op1_03_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の5番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in05 = reg_0095;
    72: op1_03_in05 = reg_0183;
    55: op1_03_in05 = imem06_in[11:8];
    73: op1_03_in05 = reg_0240;
    86: op1_03_in05 = reg_0378;
    49: op1_03_in05 = reg_0704;
    69: op1_03_in05 = reg_0845;
    61: op1_03_in05 = reg_0701;
    54: op1_03_in05 = reg_0053;
    71: op1_03_in05 = imem00_in[3:0];
    50: op1_03_in05 = reg_0106;
    68: op1_03_in05 = imem03_in[11:8];
    48: op1_03_in05 = reg_0631;
    52: op1_03_in05 = reg_0250;
    74: op1_03_in05 = reg_0575;
    75: op1_03_in05 = reg_0393;
    87: op1_03_in05 = reg_0897;
    56: op1_03_in05 = reg_0921;
    46: op1_03_in05 = reg_0473;
    60: op1_03_in05 = reg_0000;
    76: op1_03_in05 = reg_1501;
    59: op1_03_in05 = reg_0842;
    33: op1_03_in05 = reg_0518;
    57: op1_03_in05 = reg_0174;
    77: op1_03_in05 = reg_0552;
    70: op1_03_in05 = reg_0605;
    58: op1_03_in05 = reg_0526;
    44: op1_03_in05 = reg_0221;
    78: op1_03_in05 = reg_1080;
    88: op1_03_in05 = reg_1282;
    51: op1_03_in05 = reg_0981;
    79: op1_03_in05 = reg_0806;
    37: op1_03_in05 = reg_0413;
    80: op1_03_in05 = imem05_in[3:0];
    62: op1_03_in05 = reg_0456;
    34: op1_03_in05 = reg_0592;
    42: op1_03_in05 = reg_0320;
    47: op1_03_in05 = reg_0585;
    81: op1_03_in05 = reg_1244;
    85: op1_03_in05 = reg_1244;
    89: op1_03_in05 = reg_0970;
    63: op1_03_in05 = reg_0185;
    82: op1_03_in05 = reg_0794;
    83: op1_03_in05 = reg_0272;
    64: op1_03_in05 = imem02_in[15:12];
    111: op1_03_in05 = imem02_in[15:12];
    40: op1_03_in05 = reg_0333;
    84: op1_03_in05 = reg_1401;
    65: op1_03_in05 = reg_0246;
    90: op1_03_in05 = reg_0048;
    66: op1_03_in05 = reg_0974;
    91: op1_03_in05 = reg_1053;
    67: op1_03_in05 = reg_1179;
    96: op1_03_in05 = reg_1179;
    92: op1_03_in05 = reg_1028;
    93: op1_03_in05 = reg_1490;
    94: op1_03_in05 = reg_0619;
    95: op1_03_in05 = reg_0823;
    97: op1_03_in05 = reg_0225;
    98: op1_03_in05 = reg_0541;
    99: op1_03_in05 = reg_0111;
    100: op1_03_in05 = reg_0700;
    101: op1_03_in05 = reg_1301;
    102: op1_03_in05 = reg_0293;
    103: op1_03_in05 = reg_0042;
    104: op1_03_in05 = reg_1383;
    105: op1_03_in05 = reg_0780;
    106: op1_03_in05 = reg_0754;
    107: op1_03_in05 = reg_0879;
    108: op1_03_in05 = reg_0386;
    109: op1_03_in05 = reg_1453;
    110: op1_03_in05 = reg_0019;
    38: op1_03_in05 = reg_0738;
    112: op1_03_in05 = imem06_in[15:12];
    113: op1_03_in05 = reg_0423;
    114: op1_03_in05 = reg_1277;
    121: op1_03_in05 = reg_1277;
    115: op1_03_in05 = reg_1208;
    116: op1_03_in05 = reg_0392;
    117: op1_03_in05 = reg_0288;
    118: op1_03_in05 = reg_0957;
    119: op1_03_in05 = reg_1147;
    120: op1_03_in05 = reg_0215;
    122: op1_03_in05 = reg_0900;
    123: op1_03_in05 = reg_0554;
    124: op1_03_in05 = reg_1057;
    125: op1_03_in05 = reg_0411;
    126: op1_03_in05 = reg_0791;
    127: op1_03_in05 = imem06_in[3:0];
    128: op1_03_in05 = reg_0630;
    129: op1_03_in05 = reg_0008;
    130: op1_03_in05 = reg_0290;
    43: op1_03_in05 = reg_0633;
    131: op1_03_in05 = reg_0612;
    default: op1_03_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    49: op1_03_inv05 = 1;
    54: op1_03_inv05 = 1;
    68: op1_03_inv05 = 1;
    74: op1_03_inv05 = 1;
    75: op1_03_inv05 = 1;
    87: op1_03_inv05 = 1;
    56: op1_03_inv05 = 1;
    76: op1_03_inv05 = 1;
    57: op1_03_inv05 = 1;
    70: op1_03_inv05 = 1;
    44: op1_03_inv05 = 1;
    78: op1_03_inv05 = 1;
    37: op1_03_inv05 = 1;
    80: op1_03_inv05 = 1;
    62: op1_03_inv05 = 1;
    42: op1_03_inv05 = 1;
    47: op1_03_inv05 = 1;
    81: op1_03_inv05 = 1;
    63: op1_03_inv05 = 1;
    82: op1_03_inv05 = 1;
    85: op1_03_inv05 = 1;
    67: op1_03_inv05 = 1;
    95: op1_03_inv05 = 1;
    99: op1_03_inv05 = 1;
    100: op1_03_inv05 = 1;
    104: op1_03_inv05 = 1;
    105: op1_03_inv05 = 1;
    107: op1_03_inv05 = 1;
    108: op1_03_inv05 = 1;
    109: op1_03_inv05 = 1;
    110: op1_03_inv05 = 1;
    38: op1_03_inv05 = 1;
    113: op1_03_inv05 = 1;
    115: op1_03_inv05 = 1;
    116: op1_03_inv05 = 1;
    117: op1_03_inv05 = 1;
    118: op1_03_inv05 = 1;
    119: op1_03_inv05 = 1;
    120: op1_03_inv05 = 1;
    121: op1_03_inv05 = 1;
    122: op1_03_inv05 = 1;
    124: op1_03_inv05 = 1;
    126: op1_03_inv05 = 1;
    128: op1_03_inv05 = 1;
    43: op1_03_inv05 = 1;
    131: op1_03_inv05 = 1;
    default: op1_03_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の6番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in06 = reg_0181;
    72: op1_03_in06 = reg_0090;
    55: op1_03_in06 = reg_1179;
    73: op1_03_in06 = reg_0449;
    86: op1_03_in06 = reg_0891;
    49: op1_03_in06 = reg_0187;
    69: op1_03_in06 = reg_0327;
    61: op1_03_in06 = reg_0672;
    54: op1_03_in06 = reg_0086;
    71: op1_03_in06 = reg_0523;
    79: op1_03_in06 = reg_0523;
    50: op1_03_in06 = reg_0897;
    68: op1_03_in06 = reg_1280;
    48: op1_03_in06 = reg_0605;
    52: op1_03_in06 = reg_1028;
    91: op1_03_in06 = reg_1028;
    74: op1_03_in06 = reg_0631;
    75: op1_03_in06 = reg_0240;
    87: op1_03_in06 = reg_0560;
    56: op1_03_in06 = reg_0169;
    46: op1_03_in06 = imem02_in[15:12];
    60: op1_03_in06 = reg_0190;
    76: op1_03_in06 = reg_0984;
    59: op1_03_in06 = reg_1243;
    57: op1_03_in06 = reg_0066;
    77: op1_03_in06 = reg_1471;
    85: op1_03_in06 = reg_1471;
    70: op1_03_in06 = reg_0532;
    58: op1_03_in06 = reg_1225;
    44: op1_03_in06 = reg_0648;
    78: op1_03_in06 = reg_1081;
    88: op1_03_in06 = reg_0427;
    51: op1_03_in06 = reg_0990;
    37: op1_03_in06 = reg_0623;
    80: op1_03_in06 = imem05_in[15:12];
    62: op1_03_in06 = reg_0590;
    34: op1_03_in06 = reg_0103;
    42: op1_03_in06 = imem01_in[7:4];
    47: op1_03_in06 = reg_0568;
    81: op1_03_in06 = reg_1242;
    89: op1_03_in06 = reg_0972;
    63: op1_03_in06 = reg_0994;
    82: op1_03_in06 = reg_0450;
    83: op1_03_in06 = reg_0578;
    64: op1_03_in06 = reg_1029;
    40: op1_03_in06 = reg_0316;
    84: op1_03_in06 = reg_1404;
    65: op1_03_in06 = reg_1300;
    90: op1_03_in06 = reg_1226;
    66: op1_03_in06 = reg_0929;
    67: op1_03_in06 = reg_0023;
    92: op1_03_in06 = reg_0221;
    93: op1_03_in06 = reg_1487;
    94: op1_03_in06 = reg_0528;
    95: op1_03_in06 = reg_0145;
    96: op1_03_in06 = imem07_in[11:8];
    106: op1_03_in06 = imem07_in[11:8];
    97: op1_03_in06 = reg_0170;
    98: op1_03_in06 = reg_1139;
    99: op1_03_in06 = reg_0382;
    100: op1_03_in06 = reg_0701;
    101: op1_03_in06 = reg_1092;
    102: op1_03_in06 = reg_1027;
    103: op1_03_in06 = reg_0041;
    104: op1_03_in06 = reg_0088;
    105: op1_03_in06 = reg_0718;
    107: op1_03_in06 = reg_0276;
    108: op1_03_in06 = reg_0383;
    109: op1_03_in06 = reg_1227;
    110: op1_03_in06 = imem05_in[3:0];
    111: op1_03_in06 = reg_0846;
    38: op1_03_in06 = reg_0321;
    112: op1_03_in06 = reg_0795;
    43: op1_03_in06 = reg_0795;
    113: op1_03_in06 = reg_1018;
    114: op1_03_in06 = reg_1279;
    115: op1_03_in06 = reg_0882;
    116: op1_03_in06 = reg_0045;
    117: op1_03_in06 = imem04_in[15:12];
    118: op1_03_in06 = reg_1447;
    119: op1_03_in06 = reg_0421;
    120: op1_03_in06 = imem07_in[3:0];
    121: op1_03_in06 = reg_1099;
    122: op1_03_in06 = reg_1207;
    123: op1_03_in06 = reg_1052;
    124: op1_03_in06 = reg_1315;
    125: op1_03_in06 = imem04_in[7:4];
    126: op1_03_in06 = reg_1095;
    127: op1_03_in06 = reg_0263;
    128: op1_03_in06 = reg_1514;
    129: op1_03_in06 = reg_0606;
    130: op1_03_in06 = reg_0376;
    131: op1_03_in06 = reg_0149;
    default: op1_03_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_03_inv06 = 1;
    86: op1_03_inv06 = 1;
    49: op1_03_inv06 = 1;
    61: op1_03_inv06 = 1;
    48: op1_03_inv06 = 1;
    52: op1_03_inv06 = 1;
    74: op1_03_inv06 = 1;
    56: op1_03_inv06 = 1;
    59: op1_03_inv06 = 1;
    77: op1_03_inv06 = 1;
    70: op1_03_inv06 = 1;
    78: op1_03_inv06 = 1;
    88: op1_03_inv06 = 1;
    51: op1_03_inv06 = 1;
    37: op1_03_inv06 = 1;
    80: op1_03_inv06 = 1;
    62: op1_03_inv06 = 1;
    34: op1_03_inv06 = 1;
    42: op1_03_inv06 = 1;
    81: op1_03_inv06 = 1;
    82: op1_03_inv06 = 1;
    83: op1_03_inv06 = 1;
    64: op1_03_inv06 = 1;
    84: op1_03_inv06 = 1;
    65: op1_03_inv06 = 1;
    85: op1_03_inv06 = 1;
    91: op1_03_inv06 = 1;
    95: op1_03_inv06 = 1;
    99: op1_03_inv06 = 1;
    101: op1_03_inv06 = 1;
    102: op1_03_inv06 = 1;
    106: op1_03_inv06 = 1;
    107: op1_03_inv06 = 1;
    109: op1_03_inv06 = 1;
    38: op1_03_inv06 = 1;
    114: op1_03_inv06 = 1;
    116: op1_03_inv06 = 1;
    117: op1_03_inv06 = 1;
    118: op1_03_inv06 = 1;
    122: op1_03_inv06 = 1;
    123: op1_03_inv06 = 1;
    124: op1_03_inv06 = 1;
    127: op1_03_inv06 = 1;
    128: op1_03_inv06 = 1;
    129: op1_03_inv06 = 1;
    130: op1_03_inv06 = 1;
    default: op1_03_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の7番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in07 = reg_0208;
    72: op1_03_in07 = reg_0872;
    100: op1_03_in07 = reg_0872;
    55: op1_03_in07 = reg_0214;
    73: op1_03_in07 = reg_0317;
    86: op1_03_in07 = reg_0377;
    49: op1_03_in07 = reg_0672;
    69: op1_03_in07 = reg_0800;
    61: op1_03_in07 = reg_0202;
    54: op1_03_in07 = reg_0084;
    71: op1_03_in07 = reg_0221;
    50: op1_03_in07 = reg_0711;
    68: op1_03_in07 = reg_0443;
    48: op1_03_in07 = reg_0607;
    52: op1_03_in07 = reg_0136;
    74: op1_03_in07 = reg_0206;
    75: op1_03_in07 = reg_1346;
    87: op1_03_in07 = reg_1392;
    56: op1_03_in07 = reg_0777;
    46: op1_03_in07 = reg_0626;
    60: op1_03_in07 = reg_1226;
    76: op1_03_in07 = reg_0714;
    59: op1_03_in07 = reg_1053;
    57: op1_03_in07 = reg_0566;
    77: op1_03_in07 = reg_1470;
    70: op1_03_in07 = reg_0456;
    58: op1_03_in07 = reg_0295;
    44: op1_03_in07 = reg_0649;
    78: op1_03_in07 = reg_1491;
    88: op1_03_in07 = imem04_in[7:4];
    51: op1_03_in07 = reg_0054;
    79: op1_03_in07 = reg_0293;
    37: op1_03_in07 = reg_0003;
    80: op1_03_in07 = reg_0334;
    62: op1_03_in07 = reg_0561;
    34: op1_03_in07 = reg_0050;
    42: op1_03_in07 = reg_0283;
    47: op1_03_in07 = reg_0570;
    81: op1_03_in07 = reg_0580;
    89: op1_03_in07 = reg_0007;
    63: op1_03_in07 = reg_0629;
    82: op1_03_in07 = reg_1486;
    83: op1_03_in07 = reg_0750;
    64: op1_03_in07 = reg_0605;
    40: op1_03_in07 = reg_0300;
    84: op1_03_in07 = reg_0986;
    65: op1_03_in07 = reg_1093;
    85: op1_03_in07 = reg_0523;
    90: op1_03_in07 = reg_1208;
    66: op1_03_in07 = reg_0783;
    91: op1_03_in07 = reg_1230;
    67: op1_03_in07 = reg_0046;
    92: op1_03_in07 = reg_0249;
    93: op1_03_in07 = reg_0806;
    94: op1_03_in07 = reg_0529;
    95: op1_03_in07 = reg_0143;
    96: op1_03_in07 = reg_1097;
    97: op1_03_in07 = reg_0309;
    98: op1_03_in07 = reg_1282;
    99: op1_03_in07 = reg_0496;
    101: op1_03_in07 = reg_0178;
    102: op1_03_in07 = reg_1227;
    103: op1_03_in07 = reg_0011;
    104: op1_03_in07 = reg_0297;
    105: op1_03_in07 = reg_0398;
    106: op1_03_in07 = imem07_in[15:12];
    107: op1_03_in07 = reg_0934;
    108: op1_03_in07 = reg_0091;
    109: op1_03_in07 = reg_0961;
    110: op1_03_in07 = imem05_in[15:12];
    111: op1_03_in07 = reg_0608;
    38: op1_03_in07 = reg_0004;
    112: op1_03_in07 = reg_1467;
    113: op1_03_in07 = reg_0975;
    114: op1_03_in07 = reg_1141;
    115: op1_03_in07 = reg_0025;
    116: op1_03_in07 = reg_0564;
    117: op1_03_in07 = reg_0181;
    118: op1_03_in07 = reg_0113;
    119: op1_03_in07 = reg_1040;
    120: op1_03_in07 = imem07_in[7:4];
    121: op1_03_in07 = reg_1490;
    122: op1_03_in07 = reg_0432;
    123: op1_03_in07 = reg_1201;
    124: op1_03_in07 = reg_0298;
    125: op1_03_in07 = reg_1258;
    126: op1_03_in07 = reg_1057;
    127: op1_03_in07 = reg_0720;
    128: op1_03_in07 = reg_0303;
    129: op1_03_in07 = reg_0138;
    130: op1_03_in07 = reg_1092;
    43: op1_03_in07 = imem04_in[11:8];
    131: op1_03_in07 = reg_0148;
    default: op1_03_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_03_inv07 = 1;
    73: op1_03_inv07 = 1;
    49: op1_03_inv07 = 1;
    69: op1_03_inv07 = 1;
    48: op1_03_inv07 = 1;
    75: op1_03_inv07 = 1;
    87: op1_03_inv07 = 1;
    56: op1_03_inv07 = 1;
    57: op1_03_inv07 = 1;
    77: op1_03_inv07 = 1;
    58: op1_03_inv07 = 1;
    88: op1_03_inv07 = 1;
    62: op1_03_inv07 = 1;
    42: op1_03_inv07 = 1;
    82: op1_03_inv07 = 1;
    83: op1_03_inv07 = 1;
    64: op1_03_inv07 = 1;
    84: op1_03_inv07 = 1;
    65: op1_03_inv07 = 1;
    85: op1_03_inv07 = 1;
    90: op1_03_inv07 = 1;
    91: op1_03_inv07 = 1;
    92: op1_03_inv07 = 1;
    95: op1_03_inv07 = 1;
    96: op1_03_inv07 = 1;
    97: op1_03_inv07 = 1;
    98: op1_03_inv07 = 1;
    100: op1_03_inv07 = 1;
    102: op1_03_inv07 = 1;
    103: op1_03_inv07 = 1;
    104: op1_03_inv07 = 1;
    107: op1_03_inv07 = 1;
    109: op1_03_inv07 = 1;
    111: op1_03_inv07 = 1;
    38: op1_03_inv07 = 1;
    112: op1_03_inv07 = 1;
    114: op1_03_inv07 = 1;
    116: op1_03_inv07 = 1;
    117: op1_03_inv07 = 1;
    118: op1_03_inv07 = 1;
    121: op1_03_inv07 = 1;
    123: op1_03_inv07 = 1;
    124: op1_03_inv07 = 1;
    125: op1_03_inv07 = 1;
    126: op1_03_inv07 = 1;
    129: op1_03_inv07 = 1;
    130: op1_03_inv07 = 1;
    43: op1_03_inv07 = 1;
    131: op1_03_inv07 = 1;
    default: op1_03_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の8番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in08 = reg_0063;
    72: op1_03_in08 = reg_0301;
    55: op1_03_in08 = reg_0162;
    73: op1_03_in08 = reg_0751;
    112: op1_03_in08 = reg_0751;
    86: op1_03_in08 = reg_1003;
    49: op1_03_in08 = reg_0674;
    69: op1_03_in08 = reg_0279;
    61: op1_03_in08 = reg_0958;
    54: op1_03_in08 = reg_0520;
    71: op1_03_in08 = reg_1230;
    50: op1_03_in08 = reg_0307;
    68: op1_03_in08 = reg_0488;
    48: op1_03_in08 = imem02_in[3:0];
    103: op1_03_in08 = imem02_in[3:0];
    52: op1_03_in08 = reg_0485;
    74: op1_03_in08 = reg_0037;
    75: op1_03_in08 = reg_0631;
    87: op1_03_in08 = reg_0255;
    56: op1_03_in08 = reg_0465;
    46: op1_03_in08 = reg_0128;
    60: op1_03_in08 = reg_0107;
    76: op1_03_in08 = reg_1302;
    59: op1_03_in08 = reg_0523;
    57: op1_03_in08 = reg_0745;
    77: op1_03_in08 = reg_0250;
    70: op1_03_in08 = reg_0326;
    58: op1_03_in08 = reg_0419;
    44: op1_03_in08 = reg_0567;
    78: op1_03_in08 = reg_1244;
    88: op1_03_in08 = imem04_in[15:12];
    51: op1_03_in08 = reg_0778;
    79: op1_03_in08 = reg_1027;
    85: op1_03_in08 = reg_1027;
    37: op1_03_in08 = reg_0086;
    38: op1_03_in08 = reg_0086;
    80: op1_03_in08 = reg_1402;
    62: op1_03_in08 = reg_0612;
    34: op1_03_in08 = reg_0002;
    42: op1_03_in08 = reg_0486;
    47: op1_03_in08 = reg_0528;
    81: op1_03_in08 = reg_0218;
    89: op1_03_in08 = reg_1006;
    63: op1_03_in08 = reg_0667;
    82: op1_03_in08 = reg_1485;
    83: op1_03_in08 = reg_0702;
    64: op1_03_in08 = reg_0607;
    40: op1_03_in08 = reg_0275;
    84: op1_03_in08 = reg_0302;
    128: op1_03_in08 = reg_0302;
    65: op1_03_in08 = reg_1199;
    90: op1_03_in08 = reg_0104;
    118: op1_03_in08 = reg_0104;
    66: op1_03_in08 = reg_0906;
    91: op1_03_in08 = reg_1205;
    67: op1_03_in08 = reg_0214;
    92: op1_03_in08 = reg_0460;
    93: op1_03_in08 = reg_0804;
    94: op1_03_in08 = reg_0571;
    95: op1_03_in08 = reg_0180;
    96: op1_03_in08 = reg_0394;
    97: op1_03_in08 = reg_1345;
    98: op1_03_in08 = imem04_in[11:8];
    99: op1_03_in08 = reg_0684;
    100: op1_03_in08 = reg_1486;
    101: op1_03_in08 = reg_0113;
    130: op1_03_in08 = reg_0113;
    102: op1_03_in08 = reg_0249;
    104: op1_03_in08 = reg_1203;
    105: op1_03_in08 = reg_0373;
    106: op1_03_in08 = reg_0324;
    107: op1_03_in08 = reg_0254;
    108: op1_03_in08 = reg_0875;
    109: op1_03_in08 = reg_0821;
    110: op1_03_in08 = reg_1059;
    111: op1_03_in08 = reg_0712;
    113: op1_03_in08 = reg_0390;
    114: op1_03_in08 = reg_1490;
    115: op1_03_in08 = reg_0411;
    116: op1_03_in08 = reg_0697;
    117: op1_03_in08 = reg_0493;
    119: op1_03_in08 = reg_0097;
    120: op1_03_in08 = reg_0994;
    126: op1_03_in08 = reg_0994;
    121: op1_03_in08 = reg_1489;
    122: op1_03_in08 = reg_1451;
    123: op1_03_in08 = reg_0155;
    124: op1_03_in08 = reg_1056;
    125: op1_03_in08 = reg_0297;
    127: op1_03_in08 = reg_0827;
    129: op1_03_in08 = reg_0056;
    43: op1_03_in08 = reg_0319;
    131: op1_03_in08 = reg_1032;
    default: op1_03_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv08 = 1;
    69: op1_03_inv08 = 1;
    61: op1_03_inv08 = 1;
    54: op1_03_inv08 = 1;
    68: op1_03_inv08 = 1;
    48: op1_03_inv08 = 1;
    74: op1_03_inv08 = 1;
    75: op1_03_inv08 = 1;
    60: op1_03_inv08 = 1;
    76: op1_03_inv08 = 1;
    70: op1_03_inv08 = 1;
    51: op1_03_inv08 = 1;
    80: op1_03_inv08 = 1;
    34: op1_03_inv08 = 1;
    42: op1_03_inv08 = 1;
    47: op1_03_inv08 = 1;
    89: op1_03_inv08 = 1;
    82: op1_03_inv08 = 1;
    83: op1_03_inv08 = 1;
    40: op1_03_inv08 = 1;
    84: op1_03_inv08 = 1;
    85: op1_03_inv08 = 1;
    91: op1_03_inv08 = 1;
    93: op1_03_inv08 = 1;
    95: op1_03_inv08 = 1;
    96: op1_03_inv08 = 1;
    97: op1_03_inv08 = 1;
    98: op1_03_inv08 = 1;
    101: op1_03_inv08 = 1;
    105: op1_03_inv08 = 1;
    107: op1_03_inv08 = 1;
    109: op1_03_inv08 = 1;
    110: op1_03_inv08 = 1;
    111: op1_03_inv08 = 1;
    38: op1_03_inv08 = 1;
    114: op1_03_inv08 = 1;
    116: op1_03_inv08 = 1;
    117: op1_03_inv08 = 1;
    118: op1_03_inv08 = 1;
    120: op1_03_inv08 = 1;
    126: op1_03_inv08 = 1;
    127: op1_03_inv08 = 1;
    130: op1_03_inv08 = 1;
    131: op1_03_inv08 = 1;
    default: op1_03_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の9番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in09 = reg_0032;
    88: op1_03_in09 = reg_0032;
    72: op1_03_in09 = reg_0130;
    55: op1_03_in09 = reg_1060;
    73: op1_03_in09 = reg_0780;
    86: op1_03_in09 = reg_1314;
    49: op1_03_in09 = reg_0156;
    69: op1_03_in09 = reg_0313;
    61: op1_03_in09 = reg_1148;
    54: op1_03_in09 = reg_0123;
    71: op1_03_in09 = reg_0460;
    50: op1_03_in09 = reg_0006;
    68: op1_03_in09 = reg_0247;
    48: op1_03_in09 = reg_0590;
    52: op1_03_in09 = reg_0202;
    74: op1_03_in09 = reg_0458;
    75: op1_03_in09 = reg_0797;
    87: op1_03_in09 = reg_0312;
    56: op1_03_in09 = reg_0738;
    46: op1_03_in09 = reg_0381;
    60: op1_03_in09 = reg_0504;
    76: op1_03_in09 = reg_0373;
    59: op1_03_in09 = reg_0293;
    57: op1_03_in09 = reg_1181;
    77: op1_03_in09 = reg_0221;
    79: op1_03_in09 = reg_0221;
    85: op1_03_in09 = reg_0221;
    70: op1_03_in09 = reg_0972;
    58: op1_03_in09 = reg_0289;
    44: op1_03_in09 = reg_0564;
    78: op1_03_in09 = imem00_in[15:12];
    51: op1_03_in09 = reg_0056;
    37: op1_03_in09 = reg_0520;
    80: op1_03_in09 = reg_1401;
    62: op1_03_in09 = reg_1260;
    34: op1_03_in09 = reg_0053;
    42: op1_03_in09 = reg_0253;
    47: op1_03_in09 = reg_0529;
    81: op1_03_in09 = reg_0250;
    89: op1_03_in09 = reg_0068;
    63: op1_03_in09 = reg_0704;
    82: op1_03_in09 = reg_0275;
    83: op1_03_in09 = reg_0733;
    64: op1_03_in09 = reg_0169;
    40: op1_03_in09 = reg_0251;
    84: op1_03_in09 = reg_0197;
    65: op1_03_in09 = reg_0108;
    90: op1_03_in09 = reg_0882;
    130: op1_03_in09 = reg_0882;
    66: op1_03_in09 = reg_0730;
    91: op1_03_in09 = reg_1417;
    67: op1_03_in09 = reg_0213;
    92: op1_03_in09 = reg_0351;
    93: op1_03_in09 = reg_0615;
    94: op1_03_in09 = reg_0570;
    95: op1_03_in09 = reg_0965;
    96: op1_03_in09 = reg_0498;
    97: op1_03_in09 = reg_0157;
    98: op1_03_in09 = reg_0577;
    99: op1_03_in09 = reg_0878;
    100: op1_03_in09 = reg_0196;
    101: op1_03_in09 = reg_0884;
    102: op1_03_in09 = reg_0987;
    103: op1_03_in09 = reg_0607;
    104: op1_03_in09 = reg_0488;
    105: op1_03_in09 = reg_0584;
    106: op1_03_in09 = reg_1414;
    107: op1_03_in09 = reg_1207;
    108: op1_03_in09 = reg_0400;
    109: op1_03_in09 = reg_0881;
    110: op1_03_in09 = reg_0278;
    111: op1_03_in09 = reg_0973;
    38: op1_03_in09 = reg_0084;
    112: op1_03_in09 = reg_0863;
    113: op1_03_in09 = reg_0898;
    114: op1_03_in09 = reg_0804;
    115: op1_03_in09 = imem04_in[3:0];
    116: op1_03_in09 = reg_1404;
    117: op1_03_in09 = reg_0034;
    118: op1_03_in09 = reg_0350;
    119: op1_03_in09 = reg_0268;
    120: op1_03_in09 = reg_0478;
    121: op1_03_in09 = reg_0907;
    122: op1_03_in09 = reg_0126;
    123: op1_03_in09 = reg_0821;
    124: op1_03_in09 = reg_0457;
    125: op1_03_in09 = reg_1215;
    126: op1_03_in09 = reg_1055;
    127: op1_03_in09 = reg_0109;
    128: op1_03_in09 = reg_0300;
    129: op1_03_in09 = reg_0588;
    43: op1_03_in09 = reg_0487;
    131: op1_03_in09 = reg_1253;
    default: op1_03_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_03_inv09 = 1;
    73: op1_03_inv09 = 1;
    49: op1_03_inv09 = 1;
    61: op1_03_inv09 = 1;
    71: op1_03_inv09 = 1;
    48: op1_03_inv09 = 1;
    52: op1_03_inv09 = 1;
    74: op1_03_inv09 = 1;
    56: op1_03_inv09 = 1;
    60: op1_03_inv09 = 1;
    76: op1_03_inv09 = 1;
    57: op1_03_inv09 = 1;
    70: op1_03_inv09 = 1;
    58: op1_03_inv09 = 1;
    44: op1_03_inv09 = 1;
    51: op1_03_inv09 = 1;
    37: op1_03_inv09 = 1;
    62: op1_03_inv09 = 1;
    81: op1_03_inv09 = 1;
    89: op1_03_inv09 = 1;
    63: op1_03_inv09 = 1;
    82: op1_03_inv09 = 1;
    64: op1_03_inv09 = 1;
    84: op1_03_inv09 = 1;
    85: op1_03_inv09 = 1;
    90: op1_03_inv09 = 1;
    66: op1_03_inv09 = 1;
    67: op1_03_inv09 = 1;
    94: op1_03_inv09 = 1;
    97: op1_03_inv09 = 1;
    99: op1_03_inv09 = 1;
    104: op1_03_inv09 = 1;
    105: op1_03_inv09 = 1;
    106: op1_03_inv09 = 1;
    109: op1_03_inv09 = 1;
    111: op1_03_inv09 = 1;
    38: op1_03_inv09 = 1;
    113: op1_03_inv09 = 1;
    114: op1_03_inv09 = 1;
    115: op1_03_inv09 = 1;
    116: op1_03_inv09 = 1;
    119: op1_03_inv09 = 1;
    125: op1_03_inv09 = 1;
    127: op1_03_inv09 = 1;
    129: op1_03_inv09 = 1;
    130: op1_03_inv09 = 1;
    43: op1_03_inv09 = 1;
    default: op1_03_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の10番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in10 = reg_0736;
    72: op1_03_in10 = reg_0118;
    55: op1_03_in10 = reg_0994;
    73: op1_03_in10 = reg_0755;
    86: op1_03_in10 = reg_0954;
    49: op1_03_in10 = imem07_in[7:4];
    69: op1_03_in10 = reg_0757;
    61: op1_03_in10 = reg_0725;
    54: op1_03_in10 = reg_0124;
    71: op1_03_in10 = reg_0928;
    50: op1_03_in10 = reg_0829;
    68: op1_03_in10 = reg_0263;
    48: op1_03_in10 = reg_0494;
    52: op1_03_in10 = reg_0926;
    74: op1_03_in10 = reg_1035;
    75: op1_03_in10 = reg_0864;
    87: op1_03_in10 = reg_1000;
    56: op1_03_in10 = reg_0408;
    46: op1_03_in10 = reg_0138;
    60: op1_03_in10 = reg_0506;
    76: op1_03_in10 = reg_0571;
    59: op1_03_in10 = reg_0221;
    57: op1_03_in10 = reg_0540;
    77: op1_03_in10 = reg_1432;
    70: op1_03_in10 = reg_0125;
    58: op1_03_in10 = reg_0119;
    44: op1_03_in10 = reg_0066;
    78: op1_03_in10 = reg_1471;
    88: op1_03_in10 = reg_0264;
    51: op1_03_in10 = reg_0845;
    79: op1_03_in10 = reg_0460;
    37: op1_03_in10 = reg_0484;
    80: op1_03_in10 = reg_0939;
    116: op1_03_in10 = reg_0939;
    62: op1_03_in10 = imem02_in[15:12];
    34: op1_03_in10 = reg_0086;
    42: op1_03_in10 = reg_0626;
    47: op1_03_in10 = reg_0295;
    94: op1_03_in10 = reg_0295;
    81: op1_03_in10 = reg_1028;
    89: op1_03_in10 = reg_0233;
    63: op1_03_in10 = reg_0299;
    82: op1_03_in10 = reg_0130;
    83: op1_03_in10 = reg_1168;
    64: op1_03_in10 = reg_0562;
    40: op1_03_in10 = reg_0205;
    84: op1_03_in10 = reg_0601;
    65: op1_03_in10 = reg_0113;
    85: op1_03_in10 = reg_0485;
    90: op1_03_in10 = reg_1325;
    66: op1_03_in10 = reg_0960;
    91: op1_03_in10 = reg_0155;
    67: op1_03_in10 = reg_0015;
    92: op1_03_in10 = reg_0431;
    93: op1_03_in10 = reg_0805;
    95: op1_03_in10 = reg_1516;
    96: op1_03_in10 = reg_0461;
    106: op1_03_in10 = reg_0461;
    97: op1_03_in10 = reg_0139;
    98: op1_03_in10 = reg_1372;
    99: op1_03_in10 = reg_0560;
    100: op1_03_in10 = reg_0243;
    101: op1_03_in10 = reg_0378;
    102: op1_03_in10 = reg_1201;
    103: op1_03_in10 = reg_0056;
    104: op1_03_in10 = reg_1215;
    105: op1_03_in10 = reg_0622;
    107: op1_03_in10 = reg_1458;
    108: op1_03_in10 = reg_0079;
    109: op1_03_in10 = reg_0883;
    110: op1_03_in10 = reg_0996;
    111: op1_03_in10 = reg_1450;
    112: op1_03_in10 = reg_0752;
    113: op1_03_in10 = reg_0472;
    114: op1_03_in10 = reg_0803;
    115: op1_03_in10 = imem04_in[7:4];
    117: op1_03_in10 = reg_0552;
    118: op1_03_in10 = reg_0707;
    119: op1_03_in10 = reg_0368;
    120: op1_03_in10 = reg_0298;
    121: op1_03_in10 = reg_1053;
    122: op1_03_in10 = reg_0111;
    123: op1_03_in10 = reg_1405;
    124: op1_03_in10 = reg_1350;
    125: op1_03_in10 = reg_0500;
    126: op1_03_in10 = reg_0457;
    127: op1_03_in10 = reg_0398;
    128: op1_03_in10 = reg_0393;
    129: op1_03_in10 = reg_1493;
    130: op1_03_in10 = reg_1149;
    43: op1_03_in10 = reg_0096;
    131: op1_03_in10 = reg_0385;
    default: op1_03_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv10 = 1;
    55: op1_03_inv10 = 1;
    49: op1_03_inv10 = 1;
    69: op1_03_inv10 = 1;
    54: op1_03_inv10 = 1;
    68: op1_03_inv10 = 1;
    74: op1_03_inv10 = 1;
    87: op1_03_inv10 = 1;
    56: op1_03_inv10 = 1;
    60: op1_03_inv10 = 1;
    70: op1_03_inv10 = 1;
    44: op1_03_inv10 = 1;
    78: op1_03_inv10 = 1;
    88: op1_03_inv10 = 1;
    51: op1_03_inv10 = 1;
    79: op1_03_inv10 = 1;
    37: op1_03_inv10 = 1;
    63: op1_03_inv10 = 1;
    82: op1_03_inv10 = 1;
    64: op1_03_inv10 = 1;
    65: op1_03_inv10 = 1;
    85: op1_03_inv10 = 1;
    90: op1_03_inv10 = 1;
    66: op1_03_inv10 = 1;
    67: op1_03_inv10 = 1;
    99: op1_03_inv10 = 1;
    104: op1_03_inv10 = 1;
    108: op1_03_inv10 = 1;
    109: op1_03_inv10 = 1;
    111: op1_03_inv10 = 1;
    114: op1_03_inv10 = 1;
    121: op1_03_inv10 = 1;
    122: op1_03_inv10 = 1;
    123: op1_03_inv10 = 1;
    126: op1_03_inv10 = 1;
    127: op1_03_inv10 = 1;
    128: op1_03_inv10 = 1;
    130: op1_03_inv10 = 1;
    131: op1_03_inv10 = 1;
    default: op1_03_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の11番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in11 = reg_0735;
    72: op1_03_in11 = reg_1348;
    55: op1_03_in11 = reg_0998;
    73: op1_03_in11 = reg_0720;
    66: op1_03_in11 = reg_0720;
    86: op1_03_in11 = reg_1300;
    49: op1_03_in11 = reg_0777;
    69: op1_03_in11 = reg_0218;
    61: op1_03_in11 = reg_0060;
    54: op1_03_in11 = imem07_in[3:0];
    71: op1_03_in11 = reg_0886;
    50: op1_03_in11 = reg_0279;
    68: op1_03_in11 = reg_1372;
    48: op1_03_in11 = reg_0473;
    52: op1_03_in11 = reg_0188;
    74: op1_03_in11 = reg_0192;
    75: op1_03_in11 = reg_0014;
    87: op1_03_in11 = reg_0999;
    56: op1_03_in11 = reg_0621;
    46: op1_03_in11 = reg_0903;
    60: op1_03_in11 = reg_0849;
    76: op1_03_in11 = reg_0323;
    59: op1_03_in11 = reg_1205;
    121: op1_03_in11 = reg_1205;
    57: op1_03_in11 = reg_0539;
    77: op1_03_in11 = reg_0460;
    70: op1_03_in11 = reg_0105;
    58: op1_03_in11 = reg_1202;
    44: op1_03_in11 = reg_0333;
    78: op1_03_in11 = reg_1469;
    88: op1_03_in11 = reg_1340;
    51: op1_03_in11 = reg_0846;
    79: op1_03_in11 = reg_0887;
    80: op1_03_in11 = reg_0492;
    62: op1_03_in11 = reg_1207;
    42: op1_03_in11 = reg_0629;
    47: op1_03_in11 = reg_0165;
    81: op1_03_in11 = reg_1206;
    89: op1_03_in11 = reg_0710;
    63: op1_03_in11 = reg_0140;
    82: op1_03_in11 = reg_0118;
    83: op1_03_in11 = reg_1163;
    64: op1_03_in11 = reg_0560;
    40: op1_03_in11 = reg_0751;
    84: op1_03_in11 = reg_0602;
    65: op1_03_in11 = reg_1282;
    85: op1_03_in11 = reg_1454;
    90: op1_03_in11 = reg_0790;
    91: op1_03_in11 = reg_1418;
    67: op1_03_in11 = reg_0490;
    92: op1_03_in11 = reg_0440;
    93: op1_03_in11 = reg_0640;
    94: op1_03_in11 = reg_0308;
    95: op1_03_in11 = reg_0627;
    96: op1_03_in11 = reg_0994;
    97: op1_03_in11 = reg_1094;
    98: op1_03_in11 = reg_0493;
    99: op1_03_in11 = reg_1006;
    100: op1_03_in11 = reg_0151;
    101: op1_03_in11 = reg_0541;
    102: op1_03_in11 = reg_0883;
    103: op1_03_in11 = reg_0390;
    104: op1_03_in11 = reg_1233;
    105: op1_03_in11 = reg_0619;
    106: op1_03_in11 = reg_1055;
    107: op1_03_in11 = reg_0382;
    108: op1_03_in11 = reg_0402;
    109: op1_03_in11 = reg_0431;
    110: op1_03_in11 = reg_0174;
    111: op1_03_in11 = reg_1433;
    112: op1_03_in11 = reg_0780;
    113: op1_03_in11 = reg_1451;
    114: op1_03_in11 = reg_0250;
    115: op1_03_in11 = imem04_in[11:8];
    116: op1_03_in11 = reg_1169;
    117: op1_03_in11 = reg_0094;
    118: op1_03_in11 = reg_0291;
    119: op1_03_in11 = reg_0719;
    120: op1_03_in11 = reg_0892;
    122: op1_03_in11 = reg_0684;
    123: op1_03_in11 = reg_0202;
    124: op1_03_in11 = reg_1349;
    125: op1_03_in11 = reg_0421;
    126: op1_03_in11 = reg_0159;
    127: op1_03_in11 = reg_0622;
    128: op1_03_in11 = reg_0243;
    129: op1_03_in11 = reg_0497;
    130: op1_03_in11 = reg_0559;
    43: op1_03_in11 = reg_0129;
    131: op1_03_in11 = reg_0365;
    default: op1_03_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv11 = 1;
    72: op1_03_inv11 = 1;
    55: op1_03_inv11 = 1;
    73: op1_03_inv11 = 1;
    86: op1_03_inv11 = 1;
    69: op1_03_inv11 = 1;
    54: op1_03_inv11 = 1;
    71: op1_03_inv11 = 1;
    48: op1_03_inv11 = 1;
    52: op1_03_inv11 = 1;
    87: op1_03_inv11 = 1;
    56: op1_03_inv11 = 1;
    60: op1_03_inv11 = 1;
    76: op1_03_inv11 = 1;
    57: op1_03_inv11 = 1;
    77: op1_03_inv11 = 1;
    58: op1_03_inv11 = 1;
    44: op1_03_inv11 = 1;
    78: op1_03_inv11 = 1;
    88: op1_03_inv11 = 1;
    79: op1_03_inv11 = 1;
    42: op1_03_inv11 = 1;
    81: op1_03_inv11 = 1;
    89: op1_03_inv11 = 1;
    63: op1_03_inv11 = 1;
    84: op1_03_inv11 = 1;
    90: op1_03_inv11 = 1;
    66: op1_03_inv11 = 1;
    96: op1_03_inv11 = 1;
    97: op1_03_inv11 = 1;
    98: op1_03_inv11 = 1;
    100: op1_03_inv11 = 1;
    101: op1_03_inv11 = 1;
    102: op1_03_inv11 = 1;
    109: op1_03_inv11 = 1;
    110: op1_03_inv11 = 1;
    112: op1_03_inv11 = 1;
    113: op1_03_inv11 = 1;
    114: op1_03_inv11 = 1;
    115: op1_03_inv11 = 1;
    117: op1_03_inv11 = 1;
    118: op1_03_inv11 = 1;
    119: op1_03_inv11 = 1;
    121: op1_03_inv11 = 1;
    122: op1_03_inv11 = 1;
    123: op1_03_inv11 = 1;
    126: op1_03_inv11 = 1;
    130: op1_03_inv11 = 1;
    43: op1_03_inv11 = 1;
    default: op1_03_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の12番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in12 = reg_0175;
    72: op1_03_in12 = imem05_in[3:0];
    55: op1_03_in12 = imem07_in[11:8];
    73: op1_03_in12 = reg_0859;
    86: op1_03_in12 = reg_1092;
    49: op1_03_in12 = reg_0775;
    97: op1_03_in12 = reg_0775;
    69: op1_03_in12 = reg_0191;
    61: op1_03_in12 = imem01_in[3:0];
    71: op1_03_in12 = reg_0202;
    50: op1_03_in12 = reg_0276;
    68: op1_03_in12 = reg_1369;
    48: op1_03_in12 = reg_0970;
    52: op1_03_in12 = reg_0722;
    74: op1_03_in12 = reg_0730;
    75: op1_03_in12 = reg_1105;
    87: op1_03_in12 = reg_0444;
    56: op1_03_in12 = reg_0028;
    46: op1_03_in12 = reg_0006;
    60: op1_03_in12 = reg_0582;
    76: op1_03_in12 = reg_0132;
    59: op1_03_in12 = reg_0459;
    57: op1_03_in12 = reg_0937;
    77: op1_03_in12 = reg_1405;
    70: op1_03_in12 = reg_0382;
    58: op1_03_in12 = reg_1179;
    44: op1_03_in12 = reg_0332;
    64: op1_03_in12 = reg_0332;
    78: op1_03_in12 = reg_1470;
    88: op1_03_in12 = reg_0252;
    51: op1_03_in12 = reg_0007;
    79: op1_03_in12 = reg_0883;
    80: op1_03_in12 = reg_1373;
    62: op1_03_in12 = reg_0432;
    42: op1_03_in12 = reg_0628;
    47: op1_03_in12 = reg_0461;
    81: op1_03_in12 = reg_0961;
    89: op1_03_in12 = reg_0179;
    63: op1_03_in12 = reg_0158;
    82: op1_03_in12 = reg_0602;
    83: op1_03_in12 = reg_0992;
    40: op1_03_in12 = reg_0141;
    84: op1_03_in12 = reg_1346;
    65: op1_03_in12 = reg_0790;
    85: op1_03_in12 = reg_0249;
    90: op1_03_in12 = reg_0348;
    66: op1_03_in12 = reg_0869;
    91: op1_03_in12 = reg_1406;
    67: op1_03_in12 = reg_0230;
    92: op1_03_in12 = reg_0410;
    93: op1_03_in12 = reg_1053;
    94: op1_03_in12 = reg_0152;
    95: op1_03_in12 = reg_0329;
    96: op1_03_in12 = reg_0298;
    98: op1_03_in12 = reg_1258;
    99: op1_03_in12 = reg_0068;
    100: op1_03_in12 = reg_0206;
    101: op1_03_in12 = reg_0218;
    102: op1_03_in12 = reg_0886;
    103: op1_03_in12 = reg_0256;
    104: op1_03_in12 = reg_0500;
    105: op1_03_in12 = reg_0617;
    106: op1_03_in12 = reg_0667;
    107: op1_03_in12 = reg_0629;
    108: op1_03_in12 = reg_0041;
    109: op1_03_in12 = reg_0416;
    110: op1_03_in12 = reg_0604;
    111: op1_03_in12 = reg_1140;
    112: op1_03_in12 = reg_0716;
    113: op1_03_in12 = reg_0128;
    114: op1_03_in12 = reg_0987;
    115: op1_03_in12 = reg_0656;
    116: op1_03_in12 = reg_0302;
    117: op1_03_in12 = reg_0414;
    118: op1_03_in12 = reg_0288;
    119: op1_03_in12 = reg_0096;
    120: op1_03_in12 = reg_0703;
    121: op1_03_in12 = reg_0229;
    122: op1_03_in12 = reg_0381;
    123: op1_03_in12 = reg_0189;
    124: op1_03_in12 = reg_0159;
    125: op1_03_in12 = reg_0471;
    126: op1_03_in12 = reg_0224;
    127: op1_03_in12 = reg_0522;
    128: op1_03_in12 = reg_0799;
    129: op1_03_in12 = reg_0433;
    130: op1_03_in12 = reg_0291;
    43: op1_03_in12 = reg_0209;
    131: op1_03_in12 = reg_0092;
    default: op1_03_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv12 = 1;
    72: op1_03_inv12 = 1;
    55: op1_03_inv12 = 1;
    73: op1_03_inv12 = 1;
    86: op1_03_inv12 = 1;
    49: op1_03_inv12 = 1;
    69: op1_03_inv12 = 1;
    71: op1_03_inv12 = 1;
    68: op1_03_inv12 = 1;
    74: op1_03_inv12 = 1;
    75: op1_03_inv12 = 1;
    56: op1_03_inv12 = 1;
    46: op1_03_inv12 = 1;
    59: op1_03_inv12 = 1;
    77: op1_03_inv12 = 1;
    70: op1_03_inv12 = 1;
    58: op1_03_inv12 = 1;
    88: op1_03_inv12 = 1;
    51: op1_03_inv12 = 1;
    80: op1_03_inv12 = 1;
    42: op1_03_inv12 = 1;
    89: op1_03_inv12 = 1;
    63: op1_03_inv12 = 1;
    64: op1_03_inv12 = 1;
    66: op1_03_inv12 = 1;
    91: op1_03_inv12 = 1;
    67: op1_03_inv12 = 1;
    95: op1_03_inv12 = 1;
    98: op1_03_inv12 = 1;
    100: op1_03_inv12 = 1;
    101: op1_03_inv12 = 1;
    105: op1_03_inv12 = 1;
    106: op1_03_inv12 = 1;
    108: op1_03_inv12 = 1;
    110: op1_03_inv12 = 1;
    112: op1_03_inv12 = 1;
    113: op1_03_inv12 = 1;
    117: op1_03_inv12 = 1;
    118: op1_03_inv12 = 1;
    120: op1_03_inv12 = 1;
    121: op1_03_inv12 = 1;
    122: op1_03_inv12 = 1;
    124: op1_03_inv12 = 1;
    125: op1_03_inv12 = 1;
    127: op1_03_inv12 = 1;
    131: op1_03_inv12 = 1;
    default: op1_03_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の13番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in13 = reg_0831;
    72: op1_03_in13 = imem05_in[7:4];
    83: op1_03_in13 = imem05_in[7:4];
    55: op1_03_in13 = imem07_in[15:12];
    73: op1_03_in13 = reg_0133;
    86: op1_03_in13 = reg_0504;
    49: op1_03_in13 = reg_0284;
    69: op1_03_in13 = reg_0677;
    61: op1_03_in13 = imem01_in[15:12];
    71: op1_03_in13 = reg_0351;
    79: op1_03_in13 = reg_0351;
    50: op1_03_in13 = reg_0313;
    68: op1_03_in13 = reg_1368;
    48: op1_03_in13 = reg_0973;
    52: op1_03_in13 = reg_0428;
    74: op1_03_in13 = reg_0160;
    75: op1_03_in13 = reg_1064;
    87: op1_03_in13 = reg_1449;
    56: op1_03_in13 = reg_0361;
    46: op1_03_in13 = reg_0314;
    60: op1_03_in13 = reg_1144;
    76: op1_03_in13 = reg_0171;
    59: op1_03_in13 = reg_1141;
    57: op1_03_in13 = reg_0939;
    77: op1_03_in13 = reg_0202;
    91: op1_03_in13 = reg_0202;
    70: op1_03_in13 = reg_0876;
    58: op1_03_in13 = reg_0067;
    44: op1_03_in13 = imem05_in[3:0];
    78: op1_03_in13 = reg_0523;
    88: op1_03_in13 = reg_1198;
    51: op1_03_in13 = reg_0800;
    80: op1_03_in13 = reg_1348;
    62: op1_03_in13 = reg_0326;
    42: op1_03_in13 = reg_0561;
    47: op1_03_in13 = reg_0270;
    81: op1_03_in13 = reg_1417;
    89: op1_03_in13 = reg_1447;
    63: op1_03_in13 = reg_0923;
    82: op1_03_in13 = reg_0799;
    64: op1_03_in13 = reg_0631;
    84: op1_03_in13 = reg_0631;
    111: op1_03_in13 = reg_0631;
    40: op1_03_in13 = imem06_in[11:8];
    65: op1_03_in13 = reg_1280;
    85: op1_03_in13 = reg_1229;
    90: op1_03_in13 = reg_0467;
    66: op1_03_in13 = reg_0586;
    67: op1_03_in13 = reg_0378;
    92: op1_03_in13 = reg_0405;
    93: op1_03_in13 = reg_1028;
    94: op1_03_in13 = reg_0212;
    95: op1_03_in13 = reg_1093;
    96: op1_03_in13 = reg_0219;
    97: op1_03_in13 = reg_0465;
    98: op1_03_in13 = reg_1233;
    99: op1_03_in13 = reg_0009;
    100: op1_03_in13 = reg_0037;
    101: op1_03_in13 = imem04_in[7:4];
    102: op1_03_in13 = reg_0353;
    103: op1_03_in13 = reg_0432;
    104: op1_03_in13 = reg_0796;
    105: op1_03_in13 = reg_1202;
    106: op1_03_in13 = reg_0703;
    107: op1_03_in13 = reg_1433;
    108: op1_03_in13 = reg_1068;
    109: op1_03_in13 = reg_0410;
    110: op1_03_in13 = reg_0872;
    116: op1_03_in13 = reg_0872;
    112: op1_03_in13 = reg_0194;
    113: op1_03_in13 = reg_0629;
    114: op1_03_in13 = reg_1432;
    115: op1_03_in13 = reg_1258;
    117: op1_03_in13 = reg_0598;
    118: op1_03_in13 = reg_1325;
    119: op1_03_in13 = reg_0211;
    120: op1_03_in13 = reg_1350;
    121: op1_03_in13 = reg_0459;
    122: op1_03_in13 = reg_0306;
    123: op1_03_in13 = reg_0071;
    124: op1_03_in13 = reg_0156;
    125: op1_03_in13 = reg_0232;
    126: op1_03_in13 = reg_0775;
    127: op1_03_in13 = reg_0323;
    128: op1_03_in13 = reg_0828;
    129: op1_03_in13 = reg_1455;
    130: op1_03_in13 = imem04_in[11:8];
    43: op1_03_in13 = reg_0061;
    131: op1_03_in13 = reg_0595;
    default: op1_03_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv13 = 1;
    72: op1_03_inv13 = 1;
    55: op1_03_inv13 = 1;
    73: op1_03_inv13 = 1;
    69: op1_03_inv13 = 1;
    71: op1_03_inv13 = 1;
    50: op1_03_inv13 = 1;
    68: op1_03_inv13 = 1;
    48: op1_03_inv13 = 1;
    74: op1_03_inv13 = 1;
    87: op1_03_inv13 = 1;
    57: op1_03_inv13 = 1;
    77: op1_03_inv13 = 1;
    44: op1_03_inv13 = 1;
    78: op1_03_inv13 = 1;
    88: op1_03_inv13 = 1;
    79: op1_03_inv13 = 1;
    80: op1_03_inv13 = 1;
    89: op1_03_inv13 = 1;
    63: op1_03_inv13 = 1;
    64: op1_03_inv13 = 1;
    40: op1_03_inv13 = 1;
    65: op1_03_inv13 = 1;
    67: op1_03_inv13 = 1;
    92: op1_03_inv13 = 1;
    93: op1_03_inv13 = 1;
    96: op1_03_inv13 = 1;
    97: op1_03_inv13 = 1;
    98: op1_03_inv13 = 1;
    100: op1_03_inv13 = 1;
    101: op1_03_inv13 = 1;
    103: op1_03_inv13 = 1;
    108: op1_03_inv13 = 1;
    112: op1_03_inv13 = 1;
    116: op1_03_inv13 = 1;
    118: op1_03_inv13 = 1;
    119: op1_03_inv13 = 1;
    120: op1_03_inv13 = 1;
    121: op1_03_inv13 = 1;
    126: op1_03_inv13 = 1;
    128: op1_03_inv13 = 1;
    129: op1_03_inv13 = 1;
    131: op1_03_inv13 = 1;
    default: op1_03_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の14番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in14 = reg_0832;
    72: op1_03_in14 = reg_0449;
    55: op1_03_in14 = reg_0226;
    73: op1_03_in14 = imem06_in[15:12];
    86: op1_03_in14 = reg_0426;
    49: op1_03_in14 = reg_0286;
    69: op1_03_in14 = reg_0227;
    61: op1_03_in14 = reg_0695;
    122: op1_03_in14 = reg_0695;
    71: op1_03_in14 = reg_0428;
    50: op1_03_in14 = reg_0758;
    68: op1_03_in14 = reg_1367;
    48: op1_03_in14 = reg_0626;
    52: op1_03_in14 = reg_0440;
    74: op1_03_in14 = imem06_in[11:8];
    100: op1_03_in14 = imem06_in[11:8];
    75: op1_03_in14 = reg_0720;
    87: op1_03_in14 = reg_1425;
    56: op1_03_in14 = reg_0051;
    46: op1_03_in14 = reg_0313;
    60: op1_03_in14 = imem04_in[11:8];
    76: op1_03_in14 = reg_0419;
    59: op1_03_in14 = reg_1148;
    57: op1_03_in14 = reg_0477;
    77: op1_03_in14 = reg_0431;
    70: op1_03_in14 = reg_0705;
    58: op1_03_in14 = reg_0213;
    44: op1_03_in14 = reg_0367;
    78: op1_03_in14 = reg_0250;
    88: op1_03_in14 = reg_0500;
    51: op1_03_in14 = reg_0281;
    79: op1_03_in14 = reg_1321;
    80: op1_03_in14 = reg_0631;
    62: op1_03_in14 = reg_0971;
    42: op1_03_in14 = reg_0472;
    64: op1_03_in14 = reg_0472;
    47: op1_03_in14 = reg_0046;
    81: op1_03_in14 = reg_1418;
    89: op1_03_in14 = imem03_in[3:0];
    63: op1_03_in14 = reg_0489;
    82: op1_03_in14 = reg_0207;
    83: op1_03_in14 = reg_0491;
    40: op1_03_in14 = reg_0115;
    84: op1_03_in14 = reg_0039;
    65: op1_03_in14 = reg_0425;
    85: op1_03_in14 = reg_1417;
    90: op1_03_in14 = reg_0263;
    66: op1_03_in14 = reg_0622;
    91: op1_03_in14 = reg_0409;
    67: op1_03_in14 = reg_0600;
    92: op1_03_in14 = reg_0059;
    93: op1_03_in14 = reg_1230;
    94: op1_03_in14 = reg_0018;
    95: op1_03_in14 = reg_1226;
    96: op1_03_in14 = reg_0029;
    97: op1_03_in14 = reg_0740;
    98: op1_03_in14 = reg_0796;
    99: op1_03_in14 = reg_0168;
    101: op1_03_in14 = reg_0032;
    102: op1_03_in14 = reg_0188;
    103: op1_03_in14 = reg_0429;
    104: op1_03_in14 = reg_1041;
    105: op1_03_in14 = reg_0371;
    106: op1_03_in14 = reg_0140;
    107: op1_03_in14 = reg_1140;
    108: op1_03_in14 = reg_1071;
    109: op1_03_in14 = reg_0075;
    110: op1_03_in14 = reg_0318;
    111: op1_03_in14 = reg_0306;
    112: op1_03_in14 = reg_0624;
    113: op1_03_in14 = reg_0628;
    114: op1_03_in14 = reg_0524;
    115: op1_03_in14 = reg_0681;
    116: op1_03_in14 = reg_0393;
    117: op1_03_in14 = reg_1040;
    118: op1_03_in14 = reg_0790;
    119: op1_03_in14 = reg_1502;
    120: op1_03_in14 = reg_0157;
    121: op1_03_in14 = reg_0821;
    123: op1_03_in14 = reg_0058;
    124: op1_03_in14 = reg_0139;
    125: op1_03_in14 = reg_1143;
    126: op1_03_in14 = reg_0774;
    127: op1_03_in14 = reg_0132;
    128: op1_03_in14 = imem06_in[7:4];
    129: op1_03_in14 = reg_0126;
    130: op1_03_in14 = reg_0694;
    43: op1_03_in14 = reg_0019;
    131: op1_03_in14 = reg_0175;
    default: op1_03_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv14 = 1;
    86: op1_03_inv14 = 1;
    48: op1_03_inv14 = 1;
    52: op1_03_inv14 = 1;
    75: op1_03_inv14 = 1;
    46: op1_03_inv14 = 1;
    60: op1_03_inv14 = 1;
    76: op1_03_inv14 = 1;
    59: op1_03_inv14 = 1;
    57: op1_03_inv14 = 1;
    70: op1_03_inv14 = 1;
    58: op1_03_inv14 = 1;
    78: op1_03_inv14 = 1;
    88: op1_03_inv14 = 1;
    80: op1_03_inv14 = 1;
    63: op1_03_inv14 = 1;
    82: op1_03_inv14 = 1;
    64: op1_03_inv14 = 1;
    40: op1_03_inv14 = 1;
    65: op1_03_inv14 = 1;
    90: op1_03_inv14 = 1;
    66: op1_03_inv14 = 1;
    91: op1_03_inv14 = 1;
    67: op1_03_inv14 = 1;
    93: op1_03_inv14 = 1;
    95: op1_03_inv14 = 1;
    96: op1_03_inv14 = 1;
    98: op1_03_inv14 = 1;
    99: op1_03_inv14 = 1;
    101: op1_03_inv14 = 1;
    103: op1_03_inv14 = 1;
    108: op1_03_inv14 = 1;
    109: op1_03_inv14 = 1;
    110: op1_03_inv14 = 1;
    115: op1_03_inv14 = 1;
    118: op1_03_inv14 = 1;
    119: op1_03_inv14 = 1;
    121: op1_03_inv14 = 1;
    122: op1_03_inv14 = 1;
    124: op1_03_inv14 = 1;
    125: op1_03_inv14 = 1;
    127: op1_03_inv14 = 1;
    129: op1_03_inv14 = 1;
    default: op1_03_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の15番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in15 = reg_0700;
    72: op1_03_in15 = reg_0317;
    55: op1_03_in15 = reg_0851;
    73: op1_03_in15 = reg_1302;
    86: op1_03_in15 = reg_0534;
    49: op1_03_in15 = reg_0366;
    126: op1_03_in15 = reg_0366;
    69: op1_03_in15 = reg_0830;
    61: op1_03_in15 = reg_0166;
    71: op1_03_in15 = reg_0409;
    50: op1_03_in15 = reg_0573;
    68: op1_03_in15 = reg_0462;
    48: op1_03_in15 = reg_0934;
    52: op1_03_in15 = reg_0352;
    74: op1_03_in15 = reg_0373;
    75: op1_03_in15 = reg_0859;
    87: op1_03_in15 = reg_0000;
    46: op1_03_in15 = reg_0732;
    60: op1_03_in15 = reg_0396;
    76: op1_03_in15 = reg_0308;
    59: op1_03_in15 = reg_0926;
    57: op1_03_in15 = reg_0196;
    77: op1_03_in15 = reg_0416;
    70: op1_03_in15 = reg_0306;
    58: op1_03_in15 = reg_1170;
    94: op1_03_in15 = reg_1170;
    44: op1_03_in15 = reg_0873;
    78: op1_03_in15 = reg_0293;
    88: op1_03_in15 = reg_0421;
    51: op1_03_in15 = reg_0757;
    79: op1_03_in15 = reg_0122;
    80: op1_03_in15 = reg_0151;
    62: op1_03_in15 = reg_0105;
    42: op1_03_in15 = reg_0436;
    47: op1_03_in15 = reg_0215;
    81: op1_03_in15 = reg_0928;
    89: op1_03_in15 = imem03_in[7:4];
    63: op1_03_in15 = reg_0139;
    82: op1_03_in15 = imem06_in[3:0];
    83: op1_03_in15 = reg_0182;
    64: op1_03_in15 = reg_0495;
    40: op1_03_in15 = reg_0109;
    84: op1_03_in15 = reg_0014;
    65: op1_03_in15 = reg_0531;
    85: op1_03_in15 = reg_1405;
    121: op1_03_in15 = reg_1405;
    90: op1_03_in15 = reg_1372;
    66: op1_03_in15 = reg_0979;
    91: op1_03_in15 = reg_0677;
    67: op1_03_in15 = reg_0673;
    92: op1_03_in15 = reg_0058;
    93: op1_03_in15 = reg_1201;
    95: op1_03_in15 = reg_0104;
    96: op1_03_in15 = reg_0284;
    97: op1_03_in15 = reg_0415;
    98: op1_03_in15 = reg_0598;
    99: op1_03_in15 = imem03_in[11:8];
    100: op1_03_in15 = imem06_in[15:12];
    101: op1_03_in15 = reg_1369;
    102: op1_03_in15 = reg_0201;
    103: op1_03_in15 = reg_0778;
    104: op1_03_in15 = reg_1040;
    105: op1_03_in15 = reg_0754;
    106: op1_03_in15 = reg_0170;
    107: op1_03_in15 = imem02_in[3:0];
    108: op1_03_in15 = imem02_in[7:4];
    109: op1_03_in15 = reg_1321;
    110: op1_03_in15 = reg_0393;
    111: op1_03_in15 = reg_1492;
    112: op1_03_in15 = reg_0289;
    113: op1_03_in15 = reg_0381;
    114: op1_03_in15 = reg_0887;
    115: op1_03_in15 = reg_0414;
    116: op1_03_in15 = reg_0206;
    117: op1_03_in15 = reg_1004;
    118: op1_03_in15 = reg_1280;
    119: op1_03_in15 = reg_0021;
    43: op1_03_in15 = reg_0021;
    120: op1_03_in15 = reg_0738;
    122: op1_03_in15 = reg_0294;
    123: op1_03_in15 = reg_0005;
    124: op1_03_in15 = reg_0030;
    125: op1_03_in15 = reg_0268;
    127: op1_03_in15 = reg_1204;
    128: op1_03_in15 = reg_0670;
    129: op1_03_in15 = reg_0496;
    130: op1_03_in15 = reg_1257;
    131: op1_03_in15 = reg_0044;
    default: op1_03_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv15 = 1;
    73: op1_03_inv15 = 1;
    49: op1_03_inv15 = 1;
    61: op1_03_inv15 = 1;
    68: op1_03_inv15 = 1;
    48: op1_03_inv15 = 1;
    75: op1_03_inv15 = 1;
    87: op1_03_inv15 = 1;
    76: op1_03_inv15 = 1;
    59: op1_03_inv15 = 1;
    57: op1_03_inv15 = 1;
    58: op1_03_inv15 = 1;
    44: op1_03_inv15 = 1;
    78: op1_03_inv15 = 1;
    62: op1_03_inv15 = 1;
    42: op1_03_inv15 = 1;
    81: op1_03_inv15 = 1;
    89: op1_03_inv15 = 1;
    63: op1_03_inv15 = 1;
    82: op1_03_inv15 = 1;
    83: op1_03_inv15 = 1;
    64: op1_03_inv15 = 1;
    40: op1_03_inv15 = 1;
    84: op1_03_inv15 = 1;
    65: op1_03_inv15 = 1;
    66: op1_03_inv15 = 1;
    92: op1_03_inv15 = 1;
    94: op1_03_inv15 = 1;
    96: op1_03_inv15 = 1;
    97: op1_03_inv15 = 1;
    101: op1_03_inv15 = 1;
    102: op1_03_inv15 = 1;
    106: op1_03_inv15 = 1;
    109: op1_03_inv15 = 1;
    110: op1_03_inv15 = 1;
    111: op1_03_inv15 = 1;
    112: op1_03_inv15 = 1;
    115: op1_03_inv15 = 1;
    122: op1_03_inv15 = 1;
    123: op1_03_inv15 = 1;
    125: op1_03_inv15 = 1;
    126: op1_03_inv15 = 1;
    128: op1_03_inv15 = 1;
    129: op1_03_inv15 = 1;
    130: op1_03_inv15 = 1;
    131: op1_03_inv15 = 1;
    default: op1_03_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の16番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in16 = imem05_in[7:4];
    72: op1_03_in16 = reg_0038;
    55: op1_03_in16 = reg_0030;
    73: op1_03_in16 = reg_0141;
    86: op1_03_in16 = reg_0694;
    49: op1_03_in16 = reg_0740;
    69: op1_03_in16 = reg_0154;
    61: op1_03_in16 = reg_1290;
    71: op1_03_in16 = reg_0410;
    50: op1_03_in16 = reg_0678;
    68: op1_03_in16 = reg_0466;
    48: op1_03_in16 = reg_0106;
    52: op1_03_in16 = reg_0072;
    74: op1_03_in16 = reg_0584;
    75: op1_03_in16 = reg_0752;
    87: op1_03_in16 = reg_1003;
    46: op1_03_in16 = reg_0573;
    60: op1_03_in16 = reg_0463;
    76: op1_03_in16 = reg_0289;
    59: op1_03_in16 = reg_0201;
    57: op1_03_in16 = reg_0240;
    77: op1_03_in16 = reg_0405;
    70: op1_03_in16 = reg_0839;
    58: op1_03_in16 = reg_0490;
    44: op1_03_in16 = reg_0197;
    78: op1_03_in16 = reg_1453;
    88: op1_03_in16 = reg_0414;
    51: op1_03_in16 = imem03_in[3:0];
    79: op1_03_in16 = reg_1291;
    91: op1_03_in16 = reg_1291;
    80: op1_03_in16 = reg_0207;
    62: op1_03_in16 = reg_0712;
    42: op1_03_in16 = reg_0776;
    47: op1_03_in16 = reg_0923;
    81: op1_03_in16 = reg_0189;
    89: op1_03_in16 = imem03_in[11:8];
    63: op1_03_in16 = reg_0224;
    82: op1_03_in16 = imem06_in[7:4];
    83: op1_03_in16 = reg_0566;
    64: op1_03_in16 = reg_0626;
    40: op1_03_in16 = reg_0717;
    84: op1_03_in16 = imem06_in[3:0];
    65: op1_03_in16 = imem04_in[3:0];
    118: op1_03_in16 = imem04_in[3:0];
    85: op1_03_in16 = reg_0887;
    90: op1_03_in16 = reg_1368;
    66: op1_03_in16 = reg_1225;
    67: op1_03_in16 = reg_0025;
    92: op1_03_in16 = reg_0026;
    93: op1_03_in16 = reg_0229;
    94: op1_03_in16 = imem07_in[7:4];
    95: op1_03_in16 = reg_0350;
    96: op1_03_in16 = reg_0286;
    97: op1_03_in16 = reg_0413;
    98: op1_03_in16 = reg_0471;
    99: op1_03_in16 = reg_0889;
    100: op1_03_in16 = reg_0906;
    101: op1_03_in16 = reg_0164;
    102: op1_03_in16 = reg_0389;
    103: op1_03_in16 = reg_1450;
    104: op1_03_in16 = reg_1077;
    105: op1_03_in16 = reg_0195;
    106: op1_03_in16 = reg_0921;
    107: op1_03_in16 = reg_1091;
    108: op1_03_in16 = reg_0721;
    109: op1_03_in16 = imem01_in[3:0];
    123: op1_03_in16 = imem01_in[3:0];
    110: op1_03_in16 = reg_0037;
    111: op1_03_in16 = reg_0253;
    112: op1_03_in16 = reg_0396;
    113: op1_03_in16 = reg_0379;
    114: op1_03_in16 = reg_0353;
    115: op1_03_in16 = reg_1143;
    116: op1_03_in16 = reg_0565;
    117: op1_03_in16 = reg_0320;
    119: op1_03_in16 = reg_0470;
    120: op1_03_in16 = reg_0102;
    121: op1_03_in16 = reg_0476;
    122: op1_03_in16 = reg_1078;
    124: op1_03_in16 = reg_0442;
    125: op1_03_in16 = reg_0096;
    126: op1_03_in16 = reg_0741;
    127: op1_03_in16 = reg_0583;
    128: op1_03_in16 = reg_1334;
    129: op1_03_in16 = reg_1433;
    130: op1_03_in16 = reg_1258;
    43: op1_03_in16 = reg_0792;
    131: op1_03_in16 = reg_1068;
    default: op1_03_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv16 = 1;
    55: op1_03_inv16 = 1;
    73: op1_03_inv16 = 1;
    49: op1_03_inv16 = 1;
    52: op1_03_inv16 = 1;
    74: op1_03_inv16 = 1;
    75: op1_03_inv16 = 1;
    60: op1_03_inv16 = 1;
    77: op1_03_inv16 = 1;
    70: op1_03_inv16 = 1;
    78: op1_03_inv16 = 1;
    51: op1_03_inv16 = 1;
    62: op1_03_inv16 = 1;
    81: op1_03_inv16 = 1;
    63: op1_03_inv16 = 1;
    64: op1_03_inv16 = 1;
    40: op1_03_inv16 = 1;
    84: op1_03_inv16 = 1;
    65: op1_03_inv16 = 1;
    90: op1_03_inv16 = 1;
    66: op1_03_inv16 = 1;
    91: op1_03_inv16 = 1;
    93: op1_03_inv16 = 1;
    95: op1_03_inv16 = 1;
    96: op1_03_inv16 = 1;
    98: op1_03_inv16 = 1;
    99: op1_03_inv16 = 1;
    106: op1_03_inv16 = 1;
    112: op1_03_inv16 = 1;
    114: op1_03_inv16 = 1;
    115: op1_03_inv16 = 1;
    117: op1_03_inv16 = 1;
    119: op1_03_inv16 = 1;
    120: op1_03_inv16 = 1;
    121: op1_03_inv16 = 1;
    122: op1_03_inv16 = 1;
    124: op1_03_inv16 = 1;
    125: op1_03_inv16 = 1;
    126: op1_03_inv16 = 1;
    128: op1_03_inv16 = 1;
    129: op1_03_inv16 = 1;
    default: op1_03_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の17番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in17 = imem05_in[15:12];
    72: op1_03_in17 = reg_1105;
    55: op1_03_in17 = reg_0437;
    73: op1_03_in17 = reg_0585;
    86: op1_03_in17 = imem04_in[15:12];
    49: op1_03_in17 = reg_0415;
    69: op1_03_in17 = reg_0444;
    61: op1_03_in17 = reg_1254;
    71: op1_03_in17 = reg_0071;
    50: op1_03_in17 = reg_0632;
    107: op1_03_in17 = reg_0632;
    68: op1_03_in17 = reg_0681;
    48: op1_03_in17 = reg_0381;
    52: op1_03_in17 = reg_0089;
    74: op1_03_in17 = reg_0619;
    75: op1_03_in17 = reg_0172;
    87: op1_03_in17 = reg_0070;
    46: op1_03_in17 = reg_0227;
    60: op1_03_in17 = reg_0493;
    76: op1_03_in17 = reg_0023;
    105: op1_03_in17 = reg_0023;
    59: op1_03_in17 = reg_0189;
    57: op1_03_in17 = reg_0273;
    77: op1_03_in17 = reg_0134;
    70: op1_03_in17 = reg_0846;
    58: op1_03_in17 = reg_0629;
    44: op1_03_in17 = reg_0243;
    78: op1_03_in17 = reg_0987;
    88: op1_03_in17 = reg_0598;
    51: op1_03_in17 = imem03_in[7:4];
    79: op1_03_in17 = reg_0785;
    80: op1_03_in17 = reg_0206;
    62: op1_03_in17 = reg_0878;
    42: op1_03_in17 = reg_0343;
    47: op1_03_in17 = reg_0922;
    81: op1_03_in17 = reg_0428;
    89: op1_03_in17 = imem03_in[15:12];
    63: op1_03_in17 = reg_0664;
    82: op1_03_in17 = reg_1435;
    83: op1_03_in17 = reg_0131;
    64: op1_03_in17 = reg_0105;
    40: op1_03_in17 = reg_0461;
    84: op1_03_in17 = reg_0974;
    65: op1_03_in17 = imem04_in[11:8];
    85: op1_03_in17 = reg_0722;
    90: op1_03_in17 = reg_0264;
    66: op1_03_in17 = reg_0132;
    91: op1_03_in17 = reg_1255;
    67: op1_03_in17 = reg_0186;
    92: op1_03_in17 = reg_0728;
    93: op1_03_in17 = reg_0155;
    94: op1_03_in17 = imem07_in[15:12];
    95: op1_03_in17 = reg_0032;
    118: op1_03_in17 = reg_0032;
    96: op1_03_in17 = reg_0002;
    97: op1_03_in17 = reg_0050;
    98: op1_03_in17 = reg_0537;
    99: op1_03_in17 = reg_1447;
    100: op1_03_in17 = reg_1334;
    101: op1_03_in17 = reg_1257;
    102: op1_03_in17 = reg_0026;
    103: op1_03_in17 = reg_0106;
    104: op1_03_in17 = reg_0451;
    106: op1_03_in17 = reg_0223;
    108: op1_03_in17 = reg_0530;
    109: op1_03_in17 = reg_0576;
    110: op1_03_in17 = imem06_in[7:4];
    111: op1_03_in17 = reg_0848;
    112: op1_03_in17 = reg_0152;
    113: op1_03_in17 = reg_0897;
    114: op1_03_in17 = reg_0188;
    115: op1_03_in17 = reg_1312;
    116: op1_03_in17 = imem06_in[3:0];
    117: op1_03_in17 = reg_0369;
    119: op1_03_in17 = imem05_in[11:8];
    120: op1_03_in17 = reg_0103;
    121: op1_03_in17 = reg_0928;
    122: op1_03_in17 = reg_0255;
    123: op1_03_in17 = imem01_in[11:8];
    124: op1_03_in17 = reg_0740;
    125: op1_03_in17 = reg_1488;
    126: op1_03_in17 = reg_0621;
    127: op1_03_in17 = reg_0067;
    128: op1_03_in17 = reg_0696;
    129: op1_03_in17 = reg_0684;
    130: op1_03_in17 = reg_0462;
    43: op1_03_in17 = reg_0794;
    131: op1_03_in17 = reg_0662;
    default: op1_03_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv17 = 1;
    72: op1_03_inv17 = 1;
    73: op1_03_inv17 = 1;
    49: op1_03_inv17 = 1;
    71: op1_03_inv17 = 1;
    48: op1_03_inv17 = 1;
    75: op1_03_inv17 = 1;
    76: op1_03_inv17 = 1;
    57: op1_03_inv17 = 1;
    78: op1_03_inv17 = 1;
    88: op1_03_inv17 = 1;
    51: op1_03_inv17 = 1;
    80: op1_03_inv17 = 1;
    42: op1_03_inv17 = 1;
    47: op1_03_inv17 = 1;
    89: op1_03_inv17 = 1;
    82: op1_03_inv17 = 1;
    84: op1_03_inv17 = 1;
    65: op1_03_inv17 = 1;
    66: op1_03_inv17 = 1;
    67: op1_03_inv17 = 1;
    94: op1_03_inv17 = 1;
    95: op1_03_inv17 = 1;
    97: op1_03_inv17 = 1;
    98: op1_03_inv17 = 1;
    103: op1_03_inv17 = 1;
    104: op1_03_inv17 = 1;
    105: op1_03_inv17 = 1;
    106: op1_03_inv17 = 1;
    108: op1_03_inv17 = 1;
    109: op1_03_inv17 = 1;
    110: op1_03_inv17 = 1;
    111: op1_03_inv17 = 1;
    113: op1_03_inv17 = 1;
    115: op1_03_inv17 = 1;
    116: op1_03_inv17 = 1;
    117: op1_03_inv17 = 1;
    121: op1_03_inv17 = 1;
    123: op1_03_inv17 = 1;
    124: op1_03_inv17 = 1;
    125: op1_03_inv17 = 1;
    128: op1_03_inv17 = 1;
    129: op1_03_inv17 = 1;
    130: op1_03_inv17 = 1;
    43: op1_03_inv17 = 1;
    default: op1_03_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の18番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in18 = reg_0347;
    72: op1_03_in18 = reg_0195;
    55: op1_03_in18 = reg_0051;
    73: op1_03_in18 = reg_0586;
    86: op1_03_in18 = reg_0252;
    49: op1_03_in18 = reg_0413;
    69: op1_03_in18 = reg_0704;
    61: op1_03_in18 = reg_1034;
    71: op1_03_in18 = reg_0075;
    50: op1_03_in18 = reg_0707;
    68: op1_03_in18 = reg_0421;
    48: op1_03_in18 = reg_0055;
    52: op1_03_in18 = reg_0917;
    102: op1_03_in18 = reg_0917;
    74: op1_03_in18 = reg_0529;
    75: op1_03_in18 = reg_1065;
    87: op1_03_in18 = reg_1516;
    46: op1_03_in18 = reg_0198;
    99: op1_03_in18 = reg_0198;
    60: op1_03_in18 = reg_0978;
    76: op1_03_in18 = reg_0215;
    112: op1_03_in18 = reg_0215;
    59: op1_03_in18 = reg_0416;
    57: op1_03_in18 = reg_0014;
    77: op1_03_in18 = reg_0387;
    70: op1_03_in18 = reg_0007;
    58: op1_03_in18 = reg_0867;
    44: op1_03_in18 = reg_0118;
    78: op1_03_in18 = reg_1205;
    88: op1_03_in18 = reg_1041;
    51: op1_03_in18 = reg_0444;
    79: op1_03_in18 = reg_1512;
    80: op1_03_in18 = reg_0466;
    62: op1_03_in18 = reg_0069;
    42: op1_03_in18 = reg_0342;
    47: op1_03_in18 = reg_0230;
    81: op1_03_in18 = reg_0431;
    89: op1_03_in18 = reg_0891;
    63: op1_03_in18 = reg_0286;
    82: op1_03_in18 = reg_1467;
    83: op1_03_in18 = reg_1180;
    64: op1_03_in18 = reg_0056;
    40: op1_03_in18 = reg_0459;
    84: op1_03_in18 = reg_0859;
    65: op1_03_in18 = imem04_in[15:12];
    85: op1_03_in18 = reg_0189;
    90: op1_03_in18 = reg_0462;
    66: op1_03_in18 = reg_0023;
    91: op1_03_in18 = reg_1511;
    67: op1_03_in18 = reg_0922;
    92: op1_03_in18 = reg_0871;
    93: op1_03_in18 = reg_1405;
    94: op1_03_in18 = reg_0324;
    95: op1_03_in18 = reg_1368;
    96: op1_03_in18 = reg_0052;
    97: op1_03_in18 = reg_0085;
    98: op1_03_in18 = reg_1077;
    100: op1_03_in18 = reg_1209;
    101: op1_03_in18 = reg_1198;
    103: op1_03_in18 = reg_0629;
    104: op1_03_in18 = reg_0320;
    105: op1_03_in18 = reg_0212;
    106: op1_03_in18 = reg_0224;
    107: op1_03_in18 = imem03_in[7:4];
    108: op1_03_in18 = reg_0846;
    109: op1_03_in18 = reg_0401;
    123: op1_03_in18 = reg_0401;
    110: op1_03_in18 = imem06_in[15:12];
    116: op1_03_in18 = imem06_in[15:12];
    111: op1_03_in18 = reg_1091;
    113: op1_03_in18 = reg_0294;
    114: op1_03_in18 = reg_1322;
    115: op1_03_in18 = reg_0236;
    117: op1_03_in18 = reg_0062;
    118: op1_03_in18 = reg_0535;
    119: op1_03_in18 = reg_0346;
    120: op1_03_in18 = reg_1351;
    121: op1_03_in18 = reg_0089;
    122: op1_03_in18 = reg_0632;
    124: op1_03_in18 = reg_0228;
    125: op1_03_in18 = reg_0210;
    126: op1_03_in18 = reg_0620;
    127: op1_03_in18 = reg_0152;
    128: op1_03_in18 = reg_0984;
    129: op1_03_in18 = reg_0628;
    130: op1_03_in18 = reg_0488;
    43: op1_03_in18 = reg_0749;
    131: op1_03_in18 = imem02_in[11:8];
    default: op1_03_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_03_inv18 = 1;
    49: op1_03_inv18 = 1;
    69: op1_03_inv18 = 1;
    71: op1_03_inv18 = 1;
    68: op1_03_inv18 = 1;
    48: op1_03_inv18 = 1;
    52: op1_03_inv18 = 1;
    76: op1_03_inv18 = 1;
    70: op1_03_inv18 = 1;
    58: op1_03_inv18 = 1;
    44: op1_03_inv18 = 1;
    78: op1_03_inv18 = 1;
    88: op1_03_inv18 = 1;
    51: op1_03_inv18 = 1;
    79: op1_03_inv18 = 1;
    42: op1_03_inv18 = 1;
    89: op1_03_inv18 = 1;
    63: op1_03_inv18 = 1;
    83: op1_03_inv18 = 1;
    64: op1_03_inv18 = 1;
    65: op1_03_inv18 = 1;
    85: op1_03_inv18 = 1;
    90: op1_03_inv18 = 1;
    66: op1_03_inv18 = 1;
    91: op1_03_inv18 = 1;
    92: op1_03_inv18 = 1;
    93: op1_03_inv18 = 1;
    95: op1_03_inv18 = 1;
    96: op1_03_inv18 = 1;
    98: op1_03_inv18 = 1;
    99: op1_03_inv18 = 1;
    102: op1_03_inv18 = 1;
    103: op1_03_inv18 = 1;
    107: op1_03_inv18 = 1;
    113: op1_03_inv18 = 1;
    117: op1_03_inv18 = 1;
    118: op1_03_inv18 = 1;
    120: op1_03_inv18 = 1;
    123: op1_03_inv18 = 1;
    125: op1_03_inv18 = 1;
    128: op1_03_inv18 = 1;
    131: op1_03_inv18 = 1;
    default: op1_03_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の19番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in19 = reg_0066;
    72: op1_03_in19 = imem06_in[3:0];
    55: op1_03_in19 = reg_0003;
    73: op1_03_in19 = reg_0624;
    86: op1_03_in19 = reg_1215;
    49: op1_03_in19 = reg_0623;
    69: op1_03_in19 = reg_1149;
    61: op1_03_in19 = reg_0576;
    71: op1_03_in19 = reg_1324;
    50: op1_03_in19 = imem03_in[7:4];
    68: op1_03_in19 = reg_0407;
    48: op1_03_in19 = reg_0903;
    52: op1_03_in19 = reg_0610;
    74: op1_03_in19 = reg_0568;
    75: op1_03_in19 = reg_0585;
    87: op1_03_in19 = reg_1517;
    46: op1_03_in19 = reg_0375;
    60: op1_03_in19 = reg_1200;
    90: op1_03_in19 = reg_1200;
    76: op1_03_in19 = reg_0022;
    59: op1_03_in19 = reg_0134;
    57: op1_03_in19 = reg_0754;
    77: op1_03_in19 = reg_0075;
    70: op1_03_in19 = reg_0068;
    58: op1_03_in19 = reg_0299;
    44: op1_03_in19 = reg_0240;
    78: op1_03_in19 = reg_0460;
    88: op1_03_in19 = reg_0537;
    51: op1_03_in19 = reg_0377;
    79: op1_03_in19 = reg_1511;
    80: op1_03_in19 = reg_1437;
    62: op1_03_in19 = reg_0801;
    42: op1_03_in19 = reg_0055;
    64: op1_03_in19 = reg_0055;
    47: op1_03_in19 = imem07_in[3:0];
    81: op1_03_in19 = reg_0387;
    89: op1_03_in19 = reg_0314;
    63: op1_03_in19 = reg_0739;
    82: op1_03_in19 = reg_0795;
    83: op1_03_in19 = reg_1404;
    40: op1_03_in19 = reg_0152;
    84: op1_03_in19 = reg_1504;
    65: op1_03_in19 = reg_0252;
    85: op1_03_in19 = reg_0435;
    66: op1_03_in19 = reg_1055;
    91: op1_03_in19 = reg_0930;
    109: op1_03_in19 = reg_0930;
    67: op1_03_in19 = reg_1351;
    92: op1_03_in19 = reg_1512;
    93: op1_03_in19 = reg_0883;
    94: op1_03_in19 = reg_0868;
    95: op1_03_in19 = reg_0535;
    96: op1_03_in19 = reg_0085;
    98: op1_03_in19 = reg_1143;
    99: op1_03_in19 = reg_0312;
    100: op1_03_in19 = reg_0984;
    101: op1_03_in19 = reg_0574;
    102: op1_03_in19 = imem01_in[15:12];
    103: op1_03_in19 = reg_0878;
    104: op1_03_in19 = reg_0339;
    105: op1_03_in19 = reg_0213;
    106: op1_03_in19 = reg_0777;
    107: op1_03_in19 = reg_0505;
    108: op1_03_in19 = reg_0934;
    110: op1_03_in19 = reg_1105;
    111: op1_03_in19 = reg_0069;
    112: op1_03_in19 = imem07_in[11:8];
    113: op1_03_in19 = reg_0007;
    114: op1_03_in19 = reg_1255;
    115: op1_03_in19 = reg_0117;
    116: op1_03_in19 = reg_0825;
    117: op1_03_in19 = reg_1312;
    118: op1_03_in19 = reg_0731;
    119: op1_03_in19 = reg_0205;
    120: op1_03_in19 = reg_0002;
    121: op1_03_in19 = reg_0005;
    122: op1_03_in19 = reg_0006;
    123: op1_03_in19 = reg_0222;
    124: op1_03_in19 = reg_1439;
    125: op1_03_in19 = imem05_in[15:12];
    126: op1_03_in19 = reg_0592;
    127: op1_03_in19 = reg_0018;
    128: op1_03_in19 = reg_0720;
    129: op1_03_in19 = reg_0307;
    130: op1_03_in19 = reg_0281;
    43: op1_03_in19 = reg_0603;
    131: op1_03_in19 = reg_0105;
    default: op1_03_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv19 = 1;
    55: op1_03_inv19 = 1;
    73: op1_03_inv19 = 1;
    86: op1_03_inv19 = 1;
    69: op1_03_inv19 = 1;
    61: op1_03_inv19 = 1;
    71: op1_03_inv19 = 1;
    50: op1_03_inv19 = 1;
    68: op1_03_inv19 = 1;
    48: op1_03_inv19 = 1;
    52: op1_03_inv19 = 1;
    74: op1_03_inv19 = 1;
    75: op1_03_inv19 = 1;
    87: op1_03_inv19 = 1;
    76: op1_03_inv19 = 1;
    59: op1_03_inv19 = 1;
    57: op1_03_inv19 = 1;
    77: op1_03_inv19 = 1;
    58: op1_03_inv19 = 1;
    44: op1_03_inv19 = 1;
    79: op1_03_inv19 = 1;
    62: op1_03_inv19 = 1;
    42: op1_03_inv19 = 1;
    47: op1_03_inv19 = 1;
    81: op1_03_inv19 = 1;
    63: op1_03_inv19 = 1;
    82: op1_03_inv19 = 1;
    64: op1_03_inv19 = 1;
    40: op1_03_inv19 = 1;
    84: op1_03_inv19 = 1;
    65: op1_03_inv19 = 1;
    85: op1_03_inv19 = 1;
    66: op1_03_inv19 = 1;
    67: op1_03_inv19 = 1;
    92: op1_03_inv19 = 1;
    93: op1_03_inv19 = 1;
    94: op1_03_inv19 = 1;
    96: op1_03_inv19 = 1;
    98: op1_03_inv19 = 1;
    99: op1_03_inv19 = 1;
    102: op1_03_inv19 = 1;
    111: op1_03_inv19 = 1;
    113: op1_03_inv19 = 1;
    116: op1_03_inv19 = 1;
    117: op1_03_inv19 = 1;
    118: op1_03_inv19 = 1;
    119: op1_03_inv19 = 1;
    121: op1_03_inv19 = 1;
    122: op1_03_inv19 = 1;
    124: op1_03_inv19 = 1;
    125: op1_03_inv19 = 1;
    126: op1_03_inv19 = 1;
    128: op1_03_inv19 = 1;
    130: op1_03_inv19 = 1;
    131: op1_03_inv19 = 1;
    default: op1_03_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の20番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in20 = reg_0045;
    72: op1_03_in20 = reg_1064;
    55: op1_03_in20 = reg_0002;
    73: op1_03_in20 = reg_0526;
    86: op1_03_in20 = reg_1233;
    49: op1_03_in20 = reg_0137;
    69: op1_03_in20 = reg_0177;
    61: op1_03_in20 = reg_0601;
    71: op1_03_in20 = reg_0026;
    50: op1_03_in20 = reg_0349;
    89: op1_03_in20 = reg_0349;
    68: op1_03_in20 = reg_0796;
    48: op1_03_in20 = reg_0294;
    52: op1_03_in20 = reg_0609;
    74: op1_03_in20 = reg_0570;
    75: op1_03_in20 = reg_0373;
    87: op1_03_in20 = reg_1300;
    46: op1_03_in20 = reg_0235;
    60: op1_03_in20 = reg_0412;
    76: op1_03_in20 = reg_1170;
    59: op1_03_in20 = reg_0071;
    57: op1_03_in20 = reg_0751;
    77: op1_03_in20 = reg_1321;
    85: op1_03_in20 = reg_1321;
    70: op1_03_in20 = reg_0325;
    58: op1_03_in20 = reg_0309;
    44: op1_03_in20 = reg_0274;
    78: op1_03_in20 = reg_1405;
    88: op1_03_in20 = reg_0199;
    51: op1_03_in20 = reg_0049;
    79: op1_03_in20 = reg_0093;
    80: op1_03_in20 = reg_0752;
    62: op1_03_in20 = reg_0802;
    42: op1_03_in20 = reg_0024;
    47: op1_03_in20 = imem07_in[15:12];
    66: op1_03_in20 = imem07_in[15:12];
    112: op1_03_in20 = imem07_in[15:12];
    81: op1_03_in20 = reg_0073;
    63: op1_03_in20 = reg_0361;
    82: op1_03_in20 = reg_0160;
    83: op1_03_in20 = reg_0303;
    64: op1_03_in20 = reg_0711;
    40: op1_03_in20 = reg_0018;
    84: op1_03_in20 = reg_0635;
    65: op1_03_in20 = reg_0978;
    90: op1_03_in20 = reg_1147;
    95: op1_03_in20 = reg_1147;
    91: op1_03_in20 = reg_0047;
    67: op1_03_in20 = reg_0170;
    92: op1_03_in20 = reg_1511;
    93: op1_03_in20 = reg_0886;
    94: op1_03_in20 = reg_0703;
    96: op1_03_in20 = reg_0520;
    98: op1_03_in20 = reg_0337;
    99: op1_03_in20 = reg_1495;
    100: op1_03_in20 = reg_0859;
    101: op1_03_in20 = reg_0500;
    102: op1_03_in20 = reg_0372;
    103: op1_03_in20 = reg_0829;
    104: op1_03_in20 = reg_1151;
    105: op1_03_in20 = imem07_in[7:4];
    106: op1_03_in20 = reg_0029;
    107: op1_03_in20 = reg_0759;
    108: op1_03_in20 = reg_1074;
    109: op1_03_in20 = reg_0163;
    110: op1_03_in20 = reg_0908;
    111: op1_03_in20 = reg_0734;
    113: op1_03_in20 = reg_0168;
    114: op1_03_in20 = reg_0282;
    115: op1_03_in20 = reg_0538;
    125: op1_03_in20 = reg_0538;
    116: op1_03_in20 = reg_0397;
    117: op1_03_in20 = reg_0536;
    118: op1_03_in20 = reg_1258;
    119: op1_03_in20 = reg_0604;
    120: op1_03_in20 = reg_0053;
    124: op1_03_in20 = reg_0053;
    121: op1_03_in20 = reg_0723;
    122: op1_03_in20 = imem03_in[3:0];
    123: op1_03_in20 = reg_0612;
    126: op1_03_in20 = reg_0001;
    127: op1_03_in20 = reg_0135;
    128: op1_03_in20 = reg_0110;
    129: op1_03_in20 = reg_0897;
    130: op1_03_in20 = reg_1214;
    43: op1_03_in20 = reg_0334;
    131: op1_03_in20 = reg_0846;
    default: op1_03_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv20 = 1;
    55: op1_03_inv20 = 1;
    86: op1_03_inv20 = 1;
    49: op1_03_inv20 = 1;
    69: op1_03_inv20 = 1;
    61: op1_03_inv20 = 1;
    48: op1_03_inv20 = 1;
    74: op1_03_inv20 = 1;
    75: op1_03_inv20 = 1;
    87: op1_03_inv20 = 1;
    46: op1_03_inv20 = 1;
    76: op1_03_inv20 = 1;
    88: op1_03_inv20 = 1;
    62: op1_03_inv20 = 1;
    47: op1_03_inv20 = 1;
    81: op1_03_inv20 = 1;
    89: op1_03_inv20 = 1;
    63: op1_03_inv20 = 1;
    83: op1_03_inv20 = 1;
    64: op1_03_inv20 = 1;
    90: op1_03_inv20 = 1;
    66: op1_03_inv20 = 1;
    91: op1_03_inv20 = 1;
    92: op1_03_inv20 = 1;
    96: op1_03_inv20 = 1;
    98: op1_03_inv20 = 1;
    101: op1_03_inv20 = 1;
    102: op1_03_inv20 = 1;
    103: op1_03_inv20 = 1;
    104: op1_03_inv20 = 1;
    105: op1_03_inv20 = 1;
    106: op1_03_inv20 = 1;
    107: op1_03_inv20 = 1;
    110: op1_03_inv20 = 1;
    115: op1_03_inv20 = 1;
    117: op1_03_inv20 = 1;
    120: op1_03_inv20 = 1;
    123: op1_03_inv20 = 1;
    125: op1_03_inv20 = 1;
    126: op1_03_inv20 = 1;
    127: op1_03_inv20 = 1;
    128: op1_03_inv20 = 1;
    129: op1_03_inv20 = 1;
    default: op1_03_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の21番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in21 = reg_0940;
    72: op1_03_in21 = reg_1435;
    55: op1_03_in21 = reg_0085;
    73: op1_03_in21 = reg_0527;
    86: op1_03_in21 = reg_1147;
    49: op1_03_in21 = reg_0028;
    69: op1_03_in21 = imem03_in[11:8];
    122: op1_03_in21 = imem03_in[11:8];
    61: op1_03_in21 = reg_0548;
    79: op1_03_in21 = reg_0548;
    71: op1_03_in21 = reg_0005;
    50: op1_03_in21 = reg_0348;
    51: op1_03_in21 = reg_0348;
    68: op1_03_in21 = reg_0795;
    48: op1_03_in21 = reg_0845;
    52: op1_03_in21 = imem01_in[11:8];
    74: op1_03_in21 = reg_0345;
    75: op1_03_in21 = reg_0624;
    87: op1_03_in21 = reg_1208;
    46: op1_03_in21 = reg_0233;
    60: op1_03_in21 = reg_0406;
    76: op1_03_in21 = reg_0963;
    59: op1_03_in21 = reg_0072;
    57: op1_03_in21 = reg_0194;
    77: op1_03_in21 = reg_0026;
    70: op1_03_in21 = reg_0276;
    62: op1_03_in21 = reg_0276;
    58: op1_03_in21 = reg_0297;
    67: op1_03_in21 = reg_0297;
    44: op1_03_in21 = reg_0783;
    78: op1_03_in21 = reg_0883;
    88: op1_03_in21 = reg_0451;
    80: op1_03_in21 = reg_0827;
    42: op1_03_in21 = reg_0281;
    47: op1_03_in21 = reg_0156;
    81: op1_03_in21 = reg_0060;
    89: op1_03_in21 = reg_1199;
    63: op1_03_in21 = reg_0228;
    82: op1_03_in21 = reg_0720;
    83: op1_03_in21 = reg_0300;
    64: op1_03_in21 = reg_0876;
    40: op1_03_in21 = reg_0252;
    84: op1_03_in21 = reg_0115;
    65: op1_03_in21 = reg_1077;
    101: op1_03_in21 = reg_1077;
    85: op1_03_in21 = reg_0057;
    90: op1_03_in21 = reg_0421;
    66: op1_03_in21 = reg_0600;
    91: op1_03_in21 = reg_0093;
    92: op1_03_in21 = reg_0549;
    93: op1_03_in21 = reg_0188;
    94: op1_03_in21 = reg_1345;
    95: op1_03_in21 = reg_0537;
    96: op1_03_in21 = reg_0483;
    98: op1_03_in21 = reg_1107;
    99: op1_03_in21 = reg_0190;
    100: op1_03_in21 = reg_1035;
    102: op1_03_in21 = reg_0282;
    103: op1_03_in21 = reg_0801;
    104: op1_03_in21 = reg_0096;
    105: op1_03_in21 = reg_1055;
    106: op1_03_in21 = reg_0661;
    107: op1_03_in21 = reg_0677;
    108: op1_03_in21 = reg_1207;
    109: op1_03_in21 = reg_0222;
    110: op1_03_in21 = reg_0974;
    111: op1_03_in21 = reg_0759;
    112: op1_03_in21 = reg_1097;
    113: op1_03_in21 = imem03_in[3:0];
    114: op1_03_in21 = reg_1290;
    115: op1_03_in21 = reg_0278;
    116: op1_03_in21 = reg_0161;
    117: op1_03_in21 = reg_0064;
    118: op1_03_in21 = reg_0462;
    119: op1_03_in21 = reg_0173;
    120: op1_03_in21 = reg_0004;
    121: op1_03_in21 = imem01_in[3:0];
    123: op1_03_in21 = reg_1474;
    124: op1_03_in21 = reg_0123;
    125: op1_03_in21 = reg_0832;
    127: op1_03_in21 = reg_0169;
    128: op1_03_in21 = reg_0718;
    129: op1_03_in21 = reg_0802;
    130: op1_03_in21 = reg_0796;
    43: op1_03_in21 = reg_0316;
    131: op1_03_in21 = reg_1018;
    default: op1_03_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv21 = 1;
    55: op1_03_inv21 = 1;
    73: op1_03_inv21 = 1;
    61: op1_03_inv21 = 1;
    71: op1_03_inv21 = 1;
    52: op1_03_inv21 = 1;
    74: op1_03_inv21 = 1;
    87: op1_03_inv21 = 1;
    46: op1_03_inv21 = 1;
    60: op1_03_inv21 = 1;
    76: op1_03_inv21 = 1;
    59: op1_03_inv21 = 1;
    77: op1_03_inv21 = 1;
    70: op1_03_inv21 = 1;
    58: op1_03_inv21 = 1;
    44: op1_03_inv21 = 1;
    80: op1_03_inv21 = 1;
    62: op1_03_inv21 = 1;
    42: op1_03_inv21 = 1;
    47: op1_03_inv21 = 1;
    81: op1_03_inv21 = 1;
    82: op1_03_inv21 = 1;
    83: op1_03_inv21 = 1;
    40: op1_03_inv21 = 1;
    85: op1_03_inv21 = 1;
    90: op1_03_inv21 = 1;
    66: op1_03_inv21 = 1;
    91: op1_03_inv21 = 1;
    67: op1_03_inv21 = 1;
    95: op1_03_inv21 = 1;
    96: op1_03_inv21 = 1;
    99: op1_03_inv21 = 1;
    100: op1_03_inv21 = 1;
    103: op1_03_inv21 = 1;
    104: op1_03_inv21 = 1;
    105: op1_03_inv21 = 1;
    106: op1_03_inv21 = 1;
    108: op1_03_inv21 = 1;
    110: op1_03_inv21 = 1;
    114: op1_03_inv21 = 1;
    116: op1_03_inv21 = 1;
    117: op1_03_inv21 = 1;
    118: op1_03_inv21 = 1;
    119: op1_03_inv21 = 1;
    124: op1_03_inv21 = 1;
    125: op1_03_inv21 = 1;
    128: op1_03_inv21 = 1;
    129: op1_03_inv21 = 1;
    130: op1_03_inv21 = 1;
    43: op1_03_inv21 = 1;
    default: op1_03_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の22番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in22 = reg_0272;
    72: op1_03_in22 = reg_0133;
    55: op1_03_in22 = reg_0086;
    73: op1_03_in22 = reg_0522;
    86: op1_03_in22 = reg_0412;
    49: op1_03_in22 = reg_0050;
    69: op1_03_in22 = reg_1033;
    61: op1_03_in22 = reg_0259;
    71: op1_03_in22 = reg_0448;
    50: op1_03_in22 = reg_0234;
    68: op1_03_in22 = reg_0862;
    48: op1_03_in22 = reg_0009;
    52: op1_03_in22 = reg_0160;
    74: op1_03_in22 = reg_0979;
    75: op1_03_in22 = reg_0529;
    87: op1_03_in22 = reg_0108;
    46: op1_03_in22 = reg_0349;
    60: op1_03_in22 = reg_0598;
    90: op1_03_in22 = reg_0598;
    76: op1_03_in22 = reg_0034;
    59: op1_03_in22 = reg_0060;
    57: op1_03_in22 = reg_0906;
    77: op1_03_in22 = reg_0267;
    70: op1_03_in22 = reg_0758;
    58: op1_03_in22 = reg_0157;
    47: op1_03_in22 = reg_0157;
    94: op1_03_in22 = reg_0157;
    44: op1_03_in22 = reg_0195;
    78: op1_03_in22 = reg_0409;
    88: op1_03_in22 = reg_0342;
    51: op1_03_in22 = reg_0185;
    79: op1_03_in22 = reg_0743;
    109: op1_03_in22 = reg_0743;
    80: op1_03_in22 = imem06_in[7:4];
    62: op1_03_in22 = reg_0732;
    42: op1_03_in22 = reg_0280;
    81: op1_03_in22 = reg_0072;
    89: op1_03_in22 = reg_1208;
    63: op1_03_in22 = reg_0519;
    82: op1_03_in22 = reg_1323;
    83: op1_03_in22 = reg_0601;
    64: op1_03_in22 = reg_0848;
    40: op1_03_in22 = reg_0230;
    84: op1_03_in22 = reg_0373;
    65: op1_03_in22 = reg_1082;
    85: op1_03_in22 = reg_1322;
    66: op1_03_in22 = reg_0673;
    91: op1_03_in22 = reg_0547;
    67: op1_03_in22 = reg_1349;
    92: op1_03_in22 = reg_0550;
    93: op1_03_in22 = reg_0389;
    95: op1_03_in22 = reg_1077;
    96: op1_03_in22 = reg_0484;
    98: op1_03_in22 = reg_0019;
    99: op1_03_in22 = reg_1300;
    100: op1_03_in22 = reg_0716;
    101: op1_03_in22 = reg_0097;
    102: op1_03_in22 = reg_1031;
    103: op1_03_in22 = reg_1392;
    104: op1_03_in22 = reg_0211;
    105: op1_03_in22 = reg_0922;
    106: op1_03_in22 = reg_0738;
    107: op1_03_in22 = reg_0750;
    108: op1_03_in22 = reg_0436;
    110: op1_03_in22 = reg_1326;
    111: op1_03_in22 = reg_0444;
    112: op1_03_in22 = reg_0867;
    113: op1_03_in22 = reg_0677;
    114: op1_03_in22 = reg_0463;
    115: op1_03_in22 = reg_0395;
    116: op1_03_in22 = reg_1467;
    117: op1_03_in22 = reg_0063;
    118: op1_03_in22 = reg_0552;
    119: op1_03_in22 = reg_1403;
    120: op1_03_in22 = reg_0123;
    121: op1_03_in22 = reg_0982;
    122: op1_03_in22 = imem03_in[15:12];
    123: op1_03_in22 = reg_0819;
    125: op1_03_in22 = reg_0367;
    127: op1_03_in22 = reg_0498;
    128: op1_03_in22 = reg_0637;
    129: op1_03_in22 = reg_0801;
    130: op1_03_in22 = reg_0414;
    43: op1_03_in22 = reg_0317;
    131: op1_03_in22 = reg_0934;
    default: op1_03_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    49: op1_03_inv22 = 1;
    69: op1_03_inv22 = 1;
    61: op1_03_inv22 = 1;
    71: op1_03_inv22 = 1;
    48: op1_03_inv22 = 1;
    52: op1_03_inv22 = 1;
    75: op1_03_inv22 = 1;
    46: op1_03_inv22 = 1;
    60: op1_03_inv22 = 1;
    77: op1_03_inv22 = 1;
    70: op1_03_inv22 = 1;
    44: op1_03_inv22 = 1;
    78: op1_03_inv22 = 1;
    88: op1_03_inv22 = 1;
    62: op1_03_inv22 = 1;
    47: op1_03_inv22 = 1;
    89: op1_03_inv22 = 1;
    82: op1_03_inv22 = 1;
    64: op1_03_inv22 = 1;
    40: op1_03_inv22 = 1;
    65: op1_03_inv22 = 1;
    90: op1_03_inv22 = 1;
    66: op1_03_inv22 = 1;
    67: op1_03_inv22 = 1;
    94: op1_03_inv22 = 1;
    96: op1_03_inv22 = 1;
    102: op1_03_inv22 = 1;
    105: op1_03_inv22 = 1;
    106: op1_03_inv22 = 1;
    107: op1_03_inv22 = 1;
    108: op1_03_inv22 = 1;
    109: op1_03_inv22 = 1;
    110: op1_03_inv22 = 1;
    113: op1_03_inv22 = 1;
    115: op1_03_inv22 = 1;
    116: op1_03_inv22 = 1;
    118: op1_03_inv22 = 1;
    119: op1_03_inv22 = 1;
    122: op1_03_inv22 = 1;
    125: op1_03_inv22 = 1;
    128: op1_03_inv22 = 1;
    43: op1_03_inv22 = 1;
    default: op1_03_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の23番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in23 = reg_0207;
    72: op1_03_in23 = reg_1302;
    55: op1_03_in23 = reg_0087;
    73: op1_03_in23 = reg_0023;
    86: op1_03_in23 = reg_0969;
    90: op1_03_in23 = reg_0969;
    49: op1_03_in23 = reg_0001;
    69: op1_03_in23 = reg_0000;
    61: op1_03_in23 = reg_0258;
    71: op1_03_in23 = reg_1291;
    50: op1_03_in23 = reg_0789;
    68: op1_03_in23 = reg_0164;
    48: op1_03_in23 = reg_0154;
    52: op1_03_in23 = reg_1090;
    74: op1_03_in23 = reg_0171;
    75: op1_03_in23 = reg_0570;
    87: op1_03_in23 = reg_0113;
    46: op1_03_in23 = reg_0049;
    60: op1_03_in23 = reg_0798;
    76: op1_03_in23 = reg_0997;
    59: op1_03_in23 = reg_0175;
    57: op1_03_in23 = reg_0960;
    77: op1_03_in23 = reg_0917;
    70: op1_03_in23 = reg_0191;
    58: op1_03_in23 = reg_0169;
    47: op1_03_in23 = reg_0169;
    44: op1_03_in23 = reg_0730;
    78: op1_03_in23 = reg_1100;
    88: op1_03_in23 = reg_0337;
    51: op1_03_in23 = reg_1003;
    79: op1_03_in23 = reg_0609;
    109: op1_03_in23 = reg_0609;
    80: op1_03_in23 = reg_0398;
    62: op1_03_in23 = reg_0525;
    42: op1_03_in23 = reg_0314;
    81: op1_03_in23 = reg_0058;
    89: op1_03_in23 = reg_0480;
    63: op1_03_in23 = reg_1182;
    82: op1_03_in23 = reg_0780;
    83: op1_03_in23 = reg_0130;
    64: op1_03_in23 = reg_0800;
    40: op1_03_in23 = reg_0324;
    84: op1_03_in23 = reg_0624;
    65: op1_03_in23 = reg_0466;
    125: op1_03_in23 = reg_0466;
    85: op1_03_in23 = reg_0005;
    66: op1_03_in23 = reg_0674;
    91: op1_03_in23 = reg_0610;
    92: op1_03_in23 = reg_0610;
    67: op1_03_in23 = reg_0031;
    93: op1_03_in23 = reg_1322;
    94: op1_03_in23 = reg_0489;
    95: op1_03_in23 = reg_0342;
    96: op1_03_in23 = reg_0123;
    98: op1_03_in23 = reg_0210;
    99: op1_03_in23 = reg_0329;
    100: op1_03_in23 = reg_1303;
    101: op1_03_in23 = reg_0033;
    102: op1_03_in23 = reg_0166;
    103: op1_03_in23 = reg_0848;
    104: op1_03_in23 = reg_0536;
    105: op1_03_in23 = reg_0703;
    106: op1_03_in23 = reg_0415;
    107: op1_03_in23 = reg_0330;
    108: op1_03_in23 = reg_0054;
    110: op1_03_in23 = reg_1508;
    111: op1_03_in23 = reg_0709;
    112: op1_03_in23 = reg_0963;
    113: op1_03_in23 = reg_0233;
    114: op1_03_in23 = reg_0547;
    115: op1_03_in23 = reg_0251;
    116: op1_03_in23 = reg_1179;
    117: op1_03_in23 = reg_0016;
    118: op1_03_in23 = reg_1203;
    119: op1_03_in23 = reg_0937;
    121: op1_03_in23 = reg_0902;
    122: op1_03_in23 = reg_1132;
    123: op1_03_in23 = reg_0726;
    127: op1_03_in23 = reg_0738;
    128: op1_03_in23 = reg_0584;
    129: op1_03_in23 = reg_1006;
    130: op1_03_in23 = reg_1041;
    43: op1_03_in23 = reg_0538;
    131: op1_03_in23 = reg_0254;
    default: op1_03_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv23 = 1;
    55: op1_03_inv23 = 1;
    73: op1_03_inv23 = 1;
    86: op1_03_inv23 = 1;
    61: op1_03_inv23 = 1;
    68: op1_03_inv23 = 1;
    48: op1_03_inv23 = 1;
    75: op1_03_inv23 = 1;
    77: op1_03_inv23 = 1;
    44: op1_03_inv23 = 1;
    79: op1_03_inv23 = 1;
    42: op1_03_inv23 = 1;
    47: op1_03_inv23 = 1;
    81: op1_03_inv23 = 1;
    40: op1_03_inv23 = 1;
    65: op1_03_inv23 = 1;
    90: op1_03_inv23 = 1;
    66: op1_03_inv23 = 1;
    93: op1_03_inv23 = 1;
    95: op1_03_inv23 = 1;
    96: op1_03_inv23 = 1;
    98: op1_03_inv23 = 1;
    99: op1_03_inv23 = 1;
    104: op1_03_inv23 = 1;
    111: op1_03_inv23 = 1;
    114: op1_03_inv23 = 1;
    115: op1_03_inv23 = 1;
    116: op1_03_inv23 = 1;
    130: op1_03_inv23 = 1;
    43: op1_03_inv23 = 1;
    131: op1_03_inv23 = 1;
    default: op1_03_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の24番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in24 = reg_0752;
    72: op1_03_in24 = reg_0194;
    55: op1_03_in24 = reg_0519;
    73: op1_03_in24 = reg_0015;
    86: op1_03_in24 = reg_0061;
    49: op1_03_in24 = reg_0053;
    69: op1_03_in24 = reg_0789;
    61: op1_03_in24 = reg_0743;
    71: op1_03_in24 = reg_1253;
    50: op1_03_in24 = reg_1003;
    68: op1_03_in24 = reg_0129;
    48: op1_03_in24 = reg_0279;
    52: op1_03_in24 = reg_1033;
    111: op1_03_in24 = reg_1033;
    74: op1_03_in24 = reg_0419;
    75: op1_03_in24 = reg_1228;
    87: op1_03_in24 = reg_0885;
    46: op1_03_in24 = reg_0600;
    60: op1_03_in24 = reg_0454;
    76: op1_03_in24 = reg_0391;
    59: op1_03_in24 = reg_0335;
    78: op1_03_in24 = reg_0335;
    57: op1_03_in24 = reg_0398;
    77: op1_03_in24 = reg_1100;
    70: op1_03_in24 = reg_0677;
    58: op1_03_in24 = reg_0779;
    44: op1_03_in24 = reg_0141;
    88: op1_03_in24 = reg_0117;
    51: op1_03_in24 = reg_0891;
    79: op1_03_in24 = reg_0238;
    109: op1_03_in24 = reg_0238;
    80: op1_03_in24 = reg_0529;
    84: op1_03_in24 = reg_0529;
    62: op1_03_in24 = reg_0121;
    42: op1_03_in24 = reg_0313;
    47: op1_03_in24 = reg_0465;
    81: op1_03_in24 = imem01_in[7:4];
    89: op1_03_in24 = reg_0025;
    82: op1_03_in24 = reg_0110;
    83: op1_03_in24 = reg_0797;
    64: op1_03_in24 = reg_0280;
    40: op1_03_in24 = imem07_in[3:0];
    65: op1_03_in24 = reg_0552;
    85: op1_03_in24 = reg_0679;
    90: op1_03_in24 = reg_1077;
    66: op1_03_in24 = reg_0297;
    91: op1_03_in24 = reg_0260;
    67: op1_03_in24 = reg_0664;
    92: op1_03_in24 = reg_0609;
    93: op1_03_in24 = reg_0089;
    94: op1_03_in24 = reg_0139;
    95: op1_03_in24 = reg_0097;
    98: op1_03_in24 = reg_0035;
    99: op1_03_in24 = reg_0104;
    100: op1_03_in24 = reg_0637;
    110: op1_03_in24 = reg_0637;
    101: op1_03_in24 = reg_1419;
    102: op1_03_in24 = reg_0463;
    103: op1_03_in24 = reg_0217;
    104: op1_03_in24 = reg_0095;
    105: op1_03_in24 = reg_0457;
    106: op1_03_in24 = reg_0114;
    107: op1_03_in24 = reg_1001;
    108: op1_03_in24 = reg_0128;
    112: op1_03_in24 = reg_0994;
    113: op1_03_in24 = reg_1000;
    114: op1_03_in24 = reg_0747;
    115: op1_03_in24 = reg_0831;
    116: op1_03_in24 = reg_0780;
    117: op1_03_in24 = reg_0210;
    118: op1_03_in24 = reg_1233;
    119: op1_03_in24 = reg_1514;
    121: op1_03_in24 = reg_0093;
    122: op1_03_in24 = reg_0048;
    123: op1_03_in24 = reg_0147;
    125: op1_03_in24 = reg_0445;
    127: op1_03_in24 = reg_1183;
    128: op1_03_in24 = reg_0624;
    129: op1_03_in24 = reg_0069;
    130: op1_03_in24 = reg_0537;
    43: op1_03_in24 = reg_0489;
    131: op1_03_in24 = reg_1493;
    default: op1_03_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_03_inv24 = 1;
    86: op1_03_inv24 = 1;
    49: op1_03_inv24 = 1;
    71: op1_03_inv24 = 1;
    50: op1_03_inv24 = 1;
    68: op1_03_inv24 = 1;
    48: op1_03_inv24 = 1;
    74: op1_03_inv24 = 1;
    75: op1_03_inv24 = 1;
    87: op1_03_inv24 = 1;
    76: op1_03_inv24 = 1;
    57: op1_03_inv24 = 1;
    77: op1_03_inv24 = 1;
    70: op1_03_inv24 = 1;
    58: op1_03_inv24 = 1;
    44: op1_03_inv24 = 1;
    78: op1_03_inv24 = 1;
    88: op1_03_inv24 = 1;
    79: op1_03_inv24 = 1;
    89: op1_03_inv24 = 1;
    82: op1_03_inv24 = 1;
    40: op1_03_inv24 = 1;
    65: op1_03_inv24 = 1;
    91: op1_03_inv24 = 1;
    93: op1_03_inv24 = 1;
    100: op1_03_inv24 = 1;
    103: op1_03_inv24 = 1;
    104: op1_03_inv24 = 1;
    107: op1_03_inv24 = 1;
    108: op1_03_inv24 = 1;
    110: op1_03_inv24 = 1;
    116: op1_03_inv24 = 1;
    119: op1_03_inv24 = 1;
    121: op1_03_inv24 = 1;
    122: op1_03_inv24 = 1;
    123: op1_03_inv24 = 1;
    130: op1_03_inv24 = 1;
    131: op1_03_inv24 = 1;
    default: op1_03_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の25番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in25 = reg_0195;
    72: op1_03_in25 = reg_0619;
    110: op1_03_in25 = reg_0619;
    73: op1_03_in25 = reg_1170;
    86: op1_03_in25 = reg_0262;
    49: op1_03_in25 = reg_0085;
    69: op1_03_in25 = reg_0261;
    61: op1_03_in25 = reg_0553;
    71: op1_03_in25 = reg_0260;
    50: op1_03_in25 = reg_0965;
    68: op1_03_in25 = reg_0065;
    48: op1_03_in25 = reg_0276;
    52: op1_03_in25 = reg_0602;
    74: op1_03_in25 = reg_1202;
    75: op1_03_in25 = reg_1225;
    87: op1_03_in25 = imem04_in[11:8];
    46: op1_03_in25 = reg_0180;
    60: op1_03_in25 = reg_0452;
    76: op1_03_in25 = reg_1440;
    59: op1_03_in25 = reg_1068;
    57: op1_03_in25 = reg_0374;
    77: op1_03_in25 = imem01_in[15:12];
    70: op1_03_in25 = reg_0678;
    58: op1_03_in25 = reg_0774;
    44: op1_03_in25 = reg_0860;
    78: op1_03_in25 = reg_0788;
    88: op1_03_in25 = reg_1502;
    51: op1_03_in25 = reg_0889;
    79: op1_03_in25 = reg_0241;
    80: op1_03_in25 = reg_0569;
    62: op1_03_in25 = reg_0557;
    42: op1_03_in25 = reg_0732;
    122: op1_03_in25 = reg_0732;
    47: op1_03_in25 = reg_0437;
    81: op1_03_in25 = reg_0463;
    89: op1_03_in25 = reg_0443;
    82: op1_03_in25 = reg_0714;
    83: op1_03_in25 = reg_0449;
    64: op1_03_in25 = reg_0757;
    40: op1_03_in25 = imem07_in[15:12];
    84: op1_03_in25 = reg_0212;
    65: op1_03_in25 = reg_0396;
    85: op1_03_in25 = reg_0982;
    90: op1_03_in25 = reg_1065;
    66: op1_03_in25 = reg_1350;
    105: op1_03_in25 = reg_1350;
    91: op1_03_in25 = reg_0742;
    67: op1_03_in25 = reg_0442;
    92: op1_03_in25 = reg_0242;
    93: op1_03_in25 = reg_0026;
    94: op1_03_in25 = reg_0777;
    95: op1_03_in25 = reg_0582;
    98: op1_03_in25 = reg_0470;
    99: op1_03_in25 = reg_0350;
    100: op1_03_in25 = reg_0617;
    101: op1_03_in25 = reg_1143;
    102: op1_03_in25 = reg_0610;
    103: op1_03_in25 = reg_0009;
    104: op1_03_in25 = reg_0420;
    106: op1_03_in25 = reg_0361;
    107: op1_03_in25 = reg_0312;
    108: op1_03_in25 = reg_0127;
    109: op1_03_in25 = reg_0469;
    111: op1_03_in25 = reg_0311;
    112: op1_03_in25 = reg_0310;
    113: op1_03_in25 = reg_0220;
    114: op1_03_in25 = reg_0222;
    115: op1_03_in25 = reg_0648;
    116: op1_03_in25 = reg_1508;
    117: op1_03_in25 = imem05_in[15:12];
    118: op1_03_in25 = reg_1147;
    119: op1_03_in25 = reg_0418;
    121: op1_03_in25 = reg_0549;
    123: op1_03_in25 = reg_1034;
    125: op1_03_in25 = reg_0395;
    127: op1_03_in25 = reg_1057;
    128: op1_03_in25 = reg_0571;
    129: op1_03_in25 = imem03_in[11:8];
    130: op1_03_in25 = reg_0451;
    43: op1_03_in25 = reg_0490;
    131: op1_03_in25 = reg_1207;
    default: op1_03_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv25 = 1;
    86: op1_03_inv25 = 1;
    50: op1_03_inv25 = 1;
    68: op1_03_inv25 = 1;
    75: op1_03_inv25 = 1;
    46: op1_03_inv25 = 1;
    60: op1_03_inv25 = 1;
    76: op1_03_inv25 = 1;
    57: op1_03_inv25 = 1;
    78: op1_03_inv25 = 1;
    51: op1_03_inv25 = 1;
    79: op1_03_inv25 = 1;
    62: op1_03_inv25 = 1;
    42: op1_03_inv25 = 1;
    89: op1_03_inv25 = 1;
    82: op1_03_inv25 = 1;
    40: op1_03_inv25 = 1;
    65: op1_03_inv25 = 1;
    85: op1_03_inv25 = 1;
    99: op1_03_inv25 = 1;
    100: op1_03_inv25 = 1;
    104: op1_03_inv25 = 1;
    108: op1_03_inv25 = 1;
    109: op1_03_inv25 = 1;
    110: op1_03_inv25 = 1;
    111: op1_03_inv25 = 1;
    115: op1_03_inv25 = 1;
    116: op1_03_inv25 = 1;
    118: op1_03_inv25 = 1;
    119: op1_03_inv25 = 1;
    121: op1_03_inv25 = 1;
    122: op1_03_inv25 = 1;
    125: op1_03_inv25 = 1;
    127: op1_03_inv25 = 1;
    129: op1_03_inv25 = 1;
    43: op1_03_inv25 = 1;
    default: op1_03_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の26番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in26 = reg_0929;
    72: op1_03_in26 = reg_0526;
    73: op1_03_in26 = reg_1439;
    86: op1_03_in26 = reg_0096;
    49: op1_03_in26 = reg_0518;
    69: op1_03_in26 = reg_0965;
    61: op1_03_in26 = reg_0982;
    71: op1_03_in26 = reg_0547;
    52: op1_03_in26 = reg_0547;
    50: op1_03_in26 = reg_0144;
    68: op1_03_in26 = reg_0794;
    48: op1_03_in26 = reg_0314;
    74: op1_03_in26 = reg_1179;
    75: op1_03_in26 = reg_0132;
    87: op1_03_in26 = reg_0034;
    46: op1_03_in26 = reg_0220;
    60: op1_03_in26 = reg_0369;
    130: op1_03_in26 = reg_0369;
    76: op1_03_in26 = reg_1415;
    59: op1_03_in26 = reg_1031;
    57: op1_03_in26 = reg_0115;
    77: op1_03_in26 = reg_0747;
    70: op1_03_in26 = reg_0121;
    58: op1_03_in26 = reg_0593;
    44: op1_03_in26 = reg_0109;
    116: op1_03_in26 = reg_0109;
    78: op1_03_in26 = imem01_in[3:0];
    88: op1_03_in26 = reg_1503;
    51: op1_03_in26 = reg_0107;
    79: op1_03_in26 = reg_1473;
    102: op1_03_in26 = reg_1473;
    80: op1_03_in26 = reg_1228;
    62: op1_03_in26 = reg_0706;
    42: op1_03_in26 = reg_0525;
    47: op1_03_in26 = reg_0741;
    81: op1_03_in26 = reg_0549;
    89: op1_03_in26 = reg_0535;
    82: op1_03_in26 = reg_0637;
    83: op1_03_in26 = reg_0984;
    64: op1_03_in26 = reg_0573;
    40: op1_03_in26 = reg_0791;
    84: op1_03_in26 = reg_0214;
    65: op1_03_in26 = reg_0797;
    85: op1_03_in26 = reg_1512;
    90: op1_03_in26 = reg_0582;
    66: op1_03_in26 = reg_1347;
    91: op1_03_in26 = reg_1475;
    67: op1_03_in26 = reg_0413;
    92: op1_03_in26 = reg_0830;
    93: op1_03_in26 = imem01_in[11:8];
    94: op1_03_in26 = reg_0775;
    95: op1_03_in26 = imem04_in[11:8];
    98: op1_03_in26 = imem05_in[3:0];
    99: op1_03_in26 = reg_0707;
    100: op1_03_in26 = reg_0529;
    101: op1_03_in26 = reg_0062;
    103: op1_03_in26 = reg_0279;
    104: op1_03_in26 = reg_0019;
    105: op1_03_in26 = reg_0156;
    106: op1_03_in26 = reg_0053;
    107: op1_03_in26 = reg_0180;
    108: op1_03_in26 = reg_0106;
    109: op1_03_in26 = reg_1456;
    110: op1_03_in26 = reg_1202;
    111: op1_03_in26 = reg_0143;
    112: op1_03_in26 = reg_1056;
    113: op1_03_in26 = reg_0783;
    114: op1_03_in26 = reg_0743;
    115: op1_03_in26 = reg_0649;
    117: op1_03_in26 = reg_0986;
    118: op1_03_in26 = reg_0421;
    119: op1_03_in26 = reg_0450;
    121: op1_03_in26 = reg_0438;
    122: op1_03_in26 = reg_0154;
    123: op1_03_in26 = reg_0386;
    125: op1_03_in26 = reg_0251;
    127: op1_03_in26 = reg_0084;
    128: op1_03_in26 = reg_0323;
    129: op1_03_in26 = reg_1145;
    43: op1_03_in26 = reg_0477;
    131: op1_03_in26 = reg_0970;
    default: op1_03_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv26 = 1;
    73: op1_03_inv26 = 1;
    86: op1_03_inv26 = 1;
    69: op1_03_inv26 = 1;
    71: op1_03_inv26 = 1;
    87: op1_03_inv26 = 1;
    46: op1_03_inv26 = 1;
    60: op1_03_inv26 = 1;
    57: op1_03_inv26 = 1;
    70: op1_03_inv26 = 1;
    58: op1_03_inv26 = 1;
    78: op1_03_inv26 = 1;
    88: op1_03_inv26 = 1;
    79: op1_03_inv26 = 1;
    80: op1_03_inv26 = 1;
    62: op1_03_inv26 = 1;
    47: op1_03_inv26 = 1;
    89: op1_03_inv26 = 1;
    82: op1_03_inv26 = 1;
    40: op1_03_inv26 = 1;
    84: op1_03_inv26 = 1;
    65: op1_03_inv26 = 1;
    90: op1_03_inv26 = 1;
    66: op1_03_inv26 = 1;
    91: op1_03_inv26 = 1;
    92: op1_03_inv26 = 1;
    93: op1_03_inv26 = 1;
    94: op1_03_inv26 = 1;
    95: op1_03_inv26 = 1;
    100: op1_03_inv26 = 1;
    103: op1_03_inv26 = 1;
    105: op1_03_inv26 = 1;
    106: op1_03_inv26 = 1;
    108: op1_03_inv26 = 1;
    109: op1_03_inv26 = 1;
    111: op1_03_inv26 = 1;
    112: op1_03_inv26 = 1;
    113: op1_03_inv26 = 1;
    114: op1_03_inv26 = 1;
    115: op1_03_inv26 = 1;
    116: op1_03_inv26 = 1;
    118: op1_03_inv26 = 1;
    119: op1_03_inv26 = 1;
    121: op1_03_inv26 = 1;
    130: op1_03_inv26 = 1;
    default: op1_03_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の27番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in27 = reg_0979;
    100: op1_03_in27 = reg_0979;
    72: op1_03_in27 = reg_0529;
    73: op1_03_in27 = reg_1440;
    86: op1_03_in27 = reg_1189;
    49: op1_03_in27 = reg_0520;
    69: op1_03_in27 = reg_0962;
    61: op1_03_in27 = reg_0469;
    71: op1_03_in27 = reg_0548;
    50: op1_03_in27 = reg_0957;
    68: op1_03_in27 = reg_0315;
    48: op1_03_in27 = reg_0312;
    52: op1_03_in27 = reg_0242;
    74: op1_03_in27 = reg_0023;
    75: op1_03_in27 = reg_0171;
    87: op1_03_in27 = reg_1258;
    46: op1_03_in27 = reg_0880;
    60: op1_03_in27 = reg_0341;
    76: op1_03_in27 = reg_0025;
    59: op1_03_in27 = imem01_in[11:8];
    57: op1_03_in27 = reg_0671;
    77: op1_03_in27 = reg_0610;
    70: op1_03_in27 = imem03_in[15:12];
    58: op1_03_in27 = reg_0103;
    67: op1_03_in27 = reg_0103;
    44: op1_03_in27 = reg_0524;
    78: op1_03_in27 = imem01_in[7:4];
    88: op1_03_in27 = reg_0470;
    51: op1_03_in27 = reg_0113;
    79: op1_03_in27 = reg_1475;
    80: op1_03_in27 = reg_0295;
    62: op1_03_in27 = reg_0377;
    42: op1_03_in27 = reg_0734;
    47: op1_03_in27 = reg_0740;
    81: op1_03_in27 = reg_0747;
    89: op1_03_in27 = reg_0978;
    82: op1_03_in27 = reg_0194;
    83: op1_03_in27 = reg_0195;
    110: op1_03_in27 = reg_0195;
    64: op1_03_in27 = reg_0557;
    40: op1_03_in27 = reg_0775;
    84: op1_03_in27 = reg_0017;
    65: op1_03_in27 = reg_0305;
    85: op1_03_in27 = reg_0550;
    90: op1_03_in27 = reg_0836;
    66: op1_03_in27 = reg_0924;
    91: op1_03_in27 = reg_0572;
    92: op1_03_in27 = reg_1474;
    93: op1_03_in27 = reg_1090;
    94: op1_03_in27 = reg_0661;
    95: op1_03_in27 = reg_0262;
    98: op1_03_in27 = reg_0736;
    99: op1_03_in27 = reg_0378;
    101: op1_03_in27 = reg_0837;
    102: op1_03_in27 = reg_0715;
    103: op1_03_in27 = reg_0168;
    104: op1_03_in27 = imem05_in[7:4];
    105: op1_03_in27 = reg_0923;
    106: op1_03_in27 = reg_0483;
    107: op1_03_in27 = reg_1516;
    108: op1_03_in27 = reg_0382;
    109: op1_03_in27 = reg_0147;
    111: op1_03_in27 = reg_0234;
    112: op1_03_in27 = reg_1350;
    113: op1_03_in27 = reg_0823;
    114: op1_03_in27 = reg_0260;
    115: op1_03_in27 = reg_0604;
    116: op1_03_in27 = reg_0585;
    117: op1_03_in27 = reg_0346;
    118: op1_03_in27 = reg_0598;
    119: op1_03_in27 = reg_0601;
    121: op1_03_in27 = reg_1452;
    122: op1_03_in27 = reg_0709;
    123: op1_03_in27 = reg_0362;
    125: op1_03_in27 = reg_0996;
    127: op1_03_in27 = reg_0994;
    128: op1_03_in27 = reg_0244;
    129: op1_03_in27 = reg_0444;
    130: op1_03_in27 = reg_1151;
    43: op1_03_in27 = reg_0872;
    131: op1_03_in27 = reg_1455;
    default: op1_03_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv27 = 1;
    73: op1_03_inv27 = 1;
    49: op1_03_inv27 = 1;
    61: op1_03_inv27 = 1;
    48: op1_03_inv27 = 1;
    52: op1_03_inv27 = 1;
    74: op1_03_inv27 = 1;
    75: op1_03_inv27 = 1;
    87: op1_03_inv27 = 1;
    76: op1_03_inv27 = 1;
    59: op1_03_inv27 = 1;
    57: op1_03_inv27 = 1;
    77: op1_03_inv27 = 1;
    51: op1_03_inv27 = 1;
    80: op1_03_inv27 = 1;
    62: op1_03_inv27 = 1;
    81: op1_03_inv27 = 1;
    89: op1_03_inv27 = 1;
    83: op1_03_inv27 = 1;
    40: op1_03_inv27 = 1;
    84: op1_03_inv27 = 1;
    66: op1_03_inv27 = 1;
    91: op1_03_inv27 = 1;
    93: op1_03_inv27 = 1;
    94: op1_03_inv27 = 1;
    98: op1_03_inv27 = 1;
    100: op1_03_inv27 = 1;
    102: op1_03_inv27 = 1;
    105: op1_03_inv27 = 1;
    106: op1_03_inv27 = 1;
    107: op1_03_inv27 = 1;
    111: op1_03_inv27 = 1;
    113: op1_03_inv27 = 1;
    114: op1_03_inv27 = 1;
    116: op1_03_inv27 = 1;
    119: op1_03_inv27 = 1;
    121: op1_03_inv27 = 1;
    122: op1_03_inv27 = 1;
    125: op1_03_inv27 = 1;
    127: op1_03_inv27 = 1;
    129: op1_03_inv27 = 1;
    default: op1_03_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の28番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in28 = reg_0193;
    72: op1_03_in28 = reg_0568;
    73: op1_03_in28 = reg_0673;
    86: op1_03_in28 = reg_0236;
    69: op1_03_in28 = reg_1313;
    61: op1_03_in28 = reg_0930;
    71: op1_03_in28 = reg_0747;
    50: op1_03_in28 = reg_0220;
    129: op1_03_in28 = reg_0220;
    68: op1_03_in28 = reg_0750;
    48: op1_03_in28 = reg_0313;
    52: op1_03_in28 = reg_0742;
    74: op1_03_in28 = reg_0152;
    75: op1_03_in28 = reg_0289;
    87: op1_03_in28 = reg_0978;
    46: op1_03_in28 = reg_0884;
    60: op1_03_in28 = reg_0199;
    76: op1_03_in28 = reg_0186;
    59: op1_03_in28 = reg_0610;
    57: op1_03_in28 = reg_0635;
    77: op1_03_in28 = reg_0238;
    70: op1_03_in28 = reg_0177;
    58: op1_03_in28 = reg_0361;
    44: op1_03_in28 = reg_0264;
    78: op1_03_in28 = reg_0093;
    88: op1_03_in28 = reg_0702;
    51: op1_03_in28 = reg_0882;
    79: op1_03_in28 = reg_0966;
    91: op1_03_in28 = reg_0966;
    80: op1_03_in28 = reg_0308;
    62: op1_03_in28 = reg_0376;
    42: op1_03_in28 = reg_0573;
    47: op1_03_in28 = reg_0415;
    81: op1_03_in28 = reg_0260;
    89: op1_03_in28 = reg_0462;
    82: op1_03_in28 = reg_0374;
    83: op1_03_in28 = reg_0906;
    64: op1_03_in28 = reg_0707;
    40: op1_03_in28 = reg_0465;
    84: op1_03_in28 = imem07_in[3:0];
    65: op1_03_in28 = reg_0862;
    85: op1_03_in28 = reg_0787;
    90: op1_03_in28 = reg_0904;
    66: op1_03_in28 = reg_1094;
    67: op1_03_in28 = reg_0100;
    92: op1_03_in28 = reg_0726;
    93: op1_03_in28 = reg_0963;
    94: op1_03_in28 = reg_0284;
    95: op1_03_in28 = reg_0836;
    98: op1_03_in28 = reg_0315;
    99: op1_03_in28 = reg_0541;
    100: op1_03_in28 = reg_0396;
    110: op1_03_in28 = reg_0396;
    101: op1_03_in28 = reg_0835;
    102: op1_03_in28 = reg_1452;
    103: op1_03_in28 = reg_1515;
    104: op1_03_in28 = reg_1431;
    105: op1_03_in28 = reg_0139;
    107: op1_03_in28 = reg_1314;
    108: op1_03_in28 = reg_1433;
    109: op1_03_in28 = reg_0727;
    111: op1_03_in28 = reg_0000;
    112: op1_03_in28 = reg_1345;
    113: op1_03_in28 = reg_0312;
    114: op1_03_in28 = reg_0239;
    115: op1_03_in28 = reg_0392;
    116: op1_03_in28 = reg_0624;
    117: op1_03_in28 = reg_0733;
    118: op1_03_in28 = reg_0320;
    119: op1_03_in28 = reg_0196;
    121: op1_03_in28 = reg_1456;
    122: op1_03_in28 = reg_0706;
    123: op1_03_in28 = reg_0363;
    125: op1_03_in28 = reg_0066;
    127: op1_03_in28 = reg_0231;
    128: op1_03_in28 = reg_0067;
    130: op1_03_in28 = reg_0633;
    43: op1_03_in28 = reg_0251;
    131: op1_03_in28 = reg_0127;
    default: op1_03_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv28 = 1;
    86: op1_03_inv28 = 1;
    48: op1_03_inv28 = 1;
    52: op1_03_inv28 = 1;
    46: op1_03_inv28 = 1;
    59: op1_03_inv28 = 1;
    57: op1_03_inv28 = 1;
    77: op1_03_inv28 = 1;
    70: op1_03_inv28 = 1;
    44: op1_03_inv28 = 1;
    62: op1_03_inv28 = 1;
    42: op1_03_inv28 = 1;
    65: op1_03_inv28 = 1;
    85: op1_03_inv28 = 1;
    92: op1_03_inv28 = 1;
    94: op1_03_inv28 = 1;
    95: op1_03_inv28 = 1;
    98: op1_03_inv28 = 1;
    100: op1_03_inv28 = 1;
    101: op1_03_inv28 = 1;
    102: op1_03_inv28 = 1;
    103: op1_03_inv28 = 1;
    104: op1_03_inv28 = 1;
    107: op1_03_inv28 = 1;
    110: op1_03_inv28 = 1;
    112: op1_03_inv28 = 1;
    118: op1_03_inv28 = 1;
    119: op1_03_inv28 = 1;
    122: op1_03_inv28 = 1;
    123: op1_03_inv28 = 1;
    125: op1_03_inv28 = 1;
    130: op1_03_inv28 = 1;
    43: op1_03_inv28 = 1;
    default: op1_03_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の29番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in29 = reg_1058;
    72: op1_03_in29 = reg_0570;
    44: op1_03_in29 = reg_0570;
    73: op1_03_in29 = reg_0299;
    86: op1_03_in29 = reg_0932;
    69: op1_03_in29 = reg_0957;
    61: op1_03_in29 = reg_0385;
    71: op1_03_in29 = reg_0420;
    50: op1_03_in29 = reg_0882;
    68: op1_03_in29 = reg_0737;
    48: op1_03_in29 = reg_0678;
    52: op1_03_in29 = reg_0572;
    74: op1_03_in29 = reg_0213;
    75: op1_03_in29 = reg_1179;
    87: op1_03_in29 = reg_1214;
    46: op1_03_in29 = reg_0506;
    60: op1_03_in29 = reg_0340;
    76: op1_03_in29 = reg_0667;
    59: op1_03_in29 = reg_0241;
    57: op1_03_in29 = reg_0619;
    77: op1_03_in29 = reg_0830;
    70: op1_03_in29 = reg_0185;
    58: op1_03_in29 = reg_0228;
    78: op1_03_in29 = reg_0331;
    88: op1_03_in29 = reg_0466;
    51: op1_03_in29 = reg_0884;
    79: op1_03_in29 = reg_0968;
    80: op1_03_in29 = reg_1204;
    62: op1_03_in29 = reg_0963;
    42: op1_03_in29 = reg_0216;
    47: op1_03_in29 = reg_0591;
    81: op1_03_in29 = reg_1475;
    89: op1_03_in29 = reg_1233;
    82: op1_03_in29 = reg_0141;
    83: op1_03_in29 = reg_0925;
    64: op1_03_in29 = reg_0706;
    40: op1_03_in29 = reg_0287;
    84: op1_03_in29 = imem07_in[15:12];
    65: op1_03_in29 = reg_0835;
    95: op1_03_in29 = reg_0835;
    85: op1_03_in29 = reg_0874;
    90: op1_03_in29 = reg_0117;
    66: op1_03_in29 = reg_0465;
    91: op1_03_in29 = reg_0430;
    67: op1_03_in29 = reg_0002;
    92: op1_03_in29 = reg_1456;
    93: op1_03_in29 = reg_0930;
    94: op1_03_in29 = reg_0285;
    98: op1_03_in29 = reg_0735;
    99: op1_03_in29 = reg_0313;
    100: op1_03_in29 = reg_0977;
    101: op1_03_in29 = imem05_in[7:4];
    102: op1_03_in29 = reg_0290;
    103: op1_03_in29 = imem03_in[11:8];
    104: op1_03_in29 = reg_1268;
    105: op1_03_in29 = reg_0224;
    107: op1_03_in29 = reg_0597;
    108: op1_03_in29 = reg_0379;
    109: op1_03_in29 = reg_0400;
    110: op1_03_in29 = reg_0046;
    111: op1_03_in29 = reg_0556;
    112: op1_03_in29 = reg_0158;
    113: op1_03_in29 = reg_0191;
    114: op1_03_in29 = reg_0612;
    115: op1_03_in29 = reg_0334;
    116: op1_03_in29 = reg_0296;
    117: op1_03_in29 = reg_0272;
    118: op1_03_in29 = reg_0452;
    119: op1_03_in29 = reg_0602;
    121: op1_03_in29 = reg_1511;
    122: op1_03_in29 = reg_0261;
    123: op1_03_in29 = reg_0899;
    125: op1_03_in29 = reg_1403;
    127: op1_03_in29 = reg_0124;
    128: op1_03_in29 = reg_0152;
    129: op1_03_in29 = reg_0557;
    130: op1_03_in29 = reg_1503;
    43: op1_03_in29 = reg_0240;
    131: op1_03_in29 = reg_0126;
    default: op1_03_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_03_inv29 = 1;
    73: op1_03_inv29 = 1;
    86: op1_03_inv29 = 1;
    69: op1_03_inv29 = 1;
    61: op1_03_inv29 = 1;
    71: op1_03_inv29 = 1;
    68: op1_03_inv29 = 1;
    48: op1_03_inv29 = 1;
    52: op1_03_inv29 = 1;
    75: op1_03_inv29 = 1;
    87: op1_03_inv29 = 1;
    46: op1_03_inv29 = 1;
    59: op1_03_inv29 = 1;
    77: op1_03_inv29 = 1;
    70: op1_03_inv29 = 1;
    58: op1_03_inv29 = 1;
    44: op1_03_inv29 = 1;
    88: op1_03_inv29 = 1;
    79: op1_03_inv29 = 1;
    80: op1_03_inv29 = 1;
    62: op1_03_inv29 = 1;
    47: op1_03_inv29 = 1;
    89: op1_03_inv29 = 1;
    82: op1_03_inv29 = 1;
    83: op1_03_inv29 = 1;
    85: op1_03_inv29 = 1;
    94: op1_03_inv29 = 1;
    95: op1_03_inv29 = 1;
    101: op1_03_inv29 = 1;
    110: op1_03_inv29 = 1;
    114: op1_03_inv29 = 1;
    115: op1_03_inv29 = 1;
    117: op1_03_inv29 = 1;
    118: op1_03_inv29 = 1;
    121: op1_03_inv29 = 1;
    122: op1_03_inv29 = 1;
    123: op1_03_inv29 = 1;
    125: op1_03_inv29 = 1;
    127: op1_03_inv29 = 1;
    129: op1_03_inv29 = 1;
    130: op1_03_inv29 = 1;
    131: op1_03_inv29 = 1;
    default: op1_03_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の30番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_03_in30 = reg_0907;
    72: op1_03_in30 = reg_0323;
    73: op1_03_in30 = reg_0170;
    86: op1_03_in30 = reg_0016;
    90: op1_03_in30 = reg_0016;
    69: op1_03_in30 = reg_1300;
    61: op1_03_in30 = reg_0383;
    71: op1_03_in30 = reg_0241;
    50: op1_03_in30 = reg_0480;
    68: op1_03_in30 = reg_0702;
    48: op1_03_in30 = reg_0706;
    52: op1_03_in30 = reg_0967;
    114: op1_03_in30 = reg_0967;
    74: op1_03_in30 = reg_0017;
    75: op1_03_in30 = reg_0017;
    87: op1_03_in30 = reg_0537;
    46: op1_03_in30 = reg_0507;
    51: op1_03_in30 = reg_0507;
    60: op1_03_in30 = reg_0487;
    76: op1_03_in30 = reg_0225;
    59: op1_03_in30 = reg_0161;
    57: op1_03_in30 = reg_0119;
    77: op1_03_in30 = reg_0742;
    70: op1_03_in30 = reg_0199;
    58: op1_03_in30 = reg_0003;
    44: op1_03_in30 = reg_0132;
    78: op1_03_in30 = reg_0550;
    88: op1_03_in30 = reg_0332;
    79: op1_03_in30 = reg_0819;
    80: op1_03_in30 = reg_0583;
    62: op1_03_in30 = reg_0220;
    42: op1_03_in30 = reg_0288;
    47: op1_03_in30 = reg_0050;
    81: op1_03_in30 = reg_0430;
    89: op1_03_in30 = reg_1214;
    82: op1_03_in30 = reg_0373;
    83: op1_03_in30 = reg_0133;
    64: op1_03_in30 = imem03_in[3:0];
    40: op1_03_in30 = reg_0284;
    84: op1_03_in30 = reg_0461;
    65: op1_03_in30 = reg_0097;
    85: op1_03_in30 = imem01_in[3:0];
    66: op1_03_in30 = reg_0029;
    91: op1_03_in30 = reg_0726;
    67: op1_03_in30 = reg_0600;
    92: op1_03_in30 = reg_0402;
    93: op1_03_in30 = reg_0331;
    94: op1_03_in30 = reg_0441;
    95: op1_03_in30 = reg_0339;
    98: op1_03_in30 = reg_0833;
    99: op1_03_in30 = reg_0348;
    100: op1_03_in30 = reg_0152;
    101: op1_03_in30 = reg_0367;
    102: op1_03_in30 = reg_0868;
    103: op1_03_in30 = reg_0328;
    104: op1_03_in30 = reg_0831;
    105: op1_03_in30 = reg_0779;
    107: op1_03_in30 = reg_0558;
    108: op1_03_in30 = reg_1492;
    109: op1_03_in30 = reg_0724;
    110: op1_03_in30 = reg_0015;
    111: op1_03_in30 = reg_1184;
    112: op1_03_in30 = reg_0921;
    113: op1_03_in30 = reg_0234;
    115: op1_03_in30 = reg_0477;
    116: op1_03_in30 = reg_0295;
    117: op1_03_in30 = reg_0176;
    118: op1_03_in30 = reg_0342;
    119: op1_03_in30 = imem06_in[3:0];
    121: op1_03_in30 = reg_1034;
    122: op1_03_in30 = reg_0177;
    123: op1_03_in30 = reg_0092;
    125: op1_03_in30 = reg_1401;
    127: op1_03_in30 = reg_1347;
    128: op1_03_in30 = imem07_in[11:8];
    129: op1_03_in30 = reg_0198;
    130: op1_03_in30 = reg_0210;
    43: op1_03_in30 = reg_0040;
    131: op1_03_in30 = reg_0112;
    default: op1_03_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_03_inv30 = 1;
    86: op1_03_inv30 = 1;
    69: op1_03_inv30 = 1;
    71: op1_03_inv30 = 1;
    68: op1_03_inv30 = 1;
    48: op1_03_inv30 = 1;
    52: op1_03_inv30 = 1;
    87: op1_03_inv30 = 1;
    60: op1_03_inv30 = 1;
    59: op1_03_inv30 = 1;
    77: op1_03_inv30 = 1;
    70: op1_03_inv30 = 1;
    44: op1_03_inv30 = 1;
    78: op1_03_inv30 = 1;
    88: op1_03_inv30 = 1;
    51: op1_03_inv30 = 1;
    62: op1_03_inv30 = 1;
    42: op1_03_inv30 = 1;
    47: op1_03_inv30 = 1;
    89: op1_03_inv30 = 1;
    82: op1_03_inv30 = 1;
    83: op1_03_inv30 = 1;
    40: op1_03_inv30 = 1;
    84: op1_03_inv30 = 1;
    85: op1_03_inv30 = 1;
    66: op1_03_inv30 = 1;
    91: op1_03_inv30 = 1;
    67: op1_03_inv30 = 1;
    98: op1_03_inv30 = 1;
    100: op1_03_inv30 = 1;
    101: op1_03_inv30 = 1;
    102: op1_03_inv30 = 1;
    105: op1_03_inv30 = 1;
    108: op1_03_inv30 = 1;
    111: op1_03_inv30 = 1;
    113: op1_03_inv30 = 1;
    114: op1_03_inv30 = 1;
    115: op1_03_inv30 = 1;
    121: op1_03_inv30 = 1;
    122: op1_03_inv30 = 1;
    125: op1_03_inv30 = 1;
    131: op1_03_inv30 = 1;
    default: op1_03_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_03_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#3の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_03_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in00 = reg_0616;
    55: op1_04_in00 = reg_0191;
    53: op1_04_in00 = reg_0011;
    73: op1_04_in00 = reg_0578;
    64: op1_04_in00 = reg_0578;
    86: op1_04_in00 = reg_1368;
    49: op1_04_in00 = reg_0299;
    61: op1_04_in00 = reg_0866;
    69: op1_04_in00 = reg_0662;
    54: op1_04_in00 = reg_0309;
    50: op1_04_in00 = reg_0238;
    71: op1_04_in00 = reg_0554;
    82: op1_04_in00 = reg_0554;
    68: op1_04_in00 = reg_0704;
    74: op1_04_in00 = reg_0748;
    75: op1_04_in00 = reg_0841;
    87: op1_04_in00 = reg_0999;
    56: op1_04_in00 = reg_1097;
    46: op1_04_in00 = reg_0386;
    60: op1_04_in00 = reg_0411;
    99: op1_04_in00 = reg_0411;
    76: op1_04_in00 = reg_0580;
    48: op1_04_in00 = reg_0969;
    33: op1_04_in00 = reg_0286;
    57: op1_04_in00 = reg_0244;
    77: op1_04_in00 = reg_0421;
    70: op1_04_in00 = reg_0895;
    52: op1_04_in00 = imem00_in[3:0];
    96: op1_04_in00 = imem00_in[3:0];
    97: op1_04_in00 = imem00_in[3:0];
    106: op1_04_in00 = imem00_in[3:0];
    58: op1_04_in00 = reg_0582;
    78: op1_04_in00 = reg_0153;
    88: op1_04_in00 = imem03_in[7:4];
    51: op1_04_in00 = reg_0669;
    79: op1_04_in00 = reg_0938;
    59: op1_04_in00 = reg_0871;
    28: op1_04_in00 = reg_0085;
    80: op1_04_in00 = imem00_in[11:8];
    62: op1_04_in00 = reg_0541;
    37: op1_04_in00 = reg_0030;
    44: op1_04_in00 = reg_0464;
    81: op1_04_in00 = reg_0823;
    22: op1_04_in00 = reg_0114;
    34: op1_04_in00 = reg_0157;
    63: op1_04_in00 = reg_0555;
    89: op1_04_in00 = reg_0824;
    4: op1_04_in00 = imem07_in[15:12];
    40: op1_04_in00 = imem07_in[15:12];
    128: op1_04_in00 = imem07_in[15:12];
    83: op1_04_in00 = reg_0780;
    47: op1_04_in00 = reg_0289;
    84: op1_04_in00 = reg_0589;
    65: op1_04_in00 = reg_0169;
    85: op1_04_in00 = reg_0043;
    90: op1_04_in00 = imem00_in[15:12];
    126: op1_04_in00 = imem00_in[15:12];
    66: op1_04_in00 = reg_0219;
    91: op1_04_in00 = reg_1091;
    42: op1_04_in00 = imem06_in[15:12];
    67: op1_04_in00 = reg_0425;
    92: op1_04_in00 = reg_0384;
    102: op1_04_in00 = reg_0384;
    93: op1_04_in00 = reg_0830;
    94: op1_04_in00 = reg_1079;
    95: op1_04_in00 = reg_0633;
    98: op1_04_in00 = reg_0832;
    100: op1_04_in00 = reg_0214;
    101: op1_04_in00 = reg_0457;
    103: op1_04_in00 = reg_0233;
    104: op1_04_in00 = reg_0173;
    105: op1_04_in00 = imem00_in[7:4];
    120: op1_04_in00 = imem00_in[7:4];
    124: op1_04_in00 = imem00_in[7:4];
    107: op1_04_in00 = reg_1092;
    108: op1_04_in00 = reg_0711;
    109: op1_04_in00 = reg_0403;
    110: op1_04_in00 = imem07_in[3:0];
    111: op1_04_in00 = reg_1516;
    112: op1_04_in00 = reg_0924;
    113: op1_04_in00 = reg_1495;
    38: op1_04_in00 = reg_0738;
    114: op1_04_in00 = reg_0439;
    115: op1_04_in00 = reg_0302;
    116: op1_04_in00 = reg_0165;
    117: op1_04_in00 = reg_0992;
    118: op1_04_in00 = imem05_in[3:0];
    119: op1_04_in00 = reg_1058;
    121: op1_04_in00 = reg_0360;
    122: op1_04_in00 = reg_0216;
    29: op1_04_in00 = reg_0321;
    123: op1_04_in00 = reg_0727;
    125: op1_04_in00 = reg_0301;
    127: op1_04_in00 = reg_0158;
    129: op1_04_in00 = reg_0783;
    130: op1_04_in00 = imem05_in[7:4];
    131: op1_04_in00 = reg_0628;
    default: op1_04_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv00 = 1;
    53: op1_04_inv00 = 1;
    49: op1_04_inv00 = 1;
    69: op1_04_inv00 = 1;
    50: op1_04_inv00 = 1;
    71: op1_04_inv00 = 1;
    74: op1_04_inv00 = 1;
    75: op1_04_inv00 = 1;
    56: op1_04_inv00 = 1;
    46: op1_04_inv00 = 1;
    60: op1_04_inv00 = 1;
    48: op1_04_inv00 = 1;
    77: op1_04_inv00 = 1;
    52: op1_04_inv00 = 1;
    88: op1_04_inv00 = 1;
    51: op1_04_inv00 = 1;
    28: op1_04_inv00 = 1;
    62: op1_04_inv00 = 1;
    89: op1_04_inv00 = 1;
    47: op1_04_inv00 = 1;
    40: op1_04_inv00 = 1;
    90: op1_04_inv00 = 1;
    66: op1_04_inv00 = 1;
    42: op1_04_inv00 = 1;
    92: op1_04_inv00 = 1;
    96: op1_04_inv00 = 1;
    97: op1_04_inv00 = 1;
    98: op1_04_inv00 = 1;
    99: op1_04_inv00 = 1;
    100: op1_04_inv00 = 1;
    102: op1_04_inv00 = 1;
    105: op1_04_inv00 = 1;
    106: op1_04_inv00 = 1;
    107: op1_04_inv00 = 1;
    108: op1_04_inv00 = 1;
    111: op1_04_inv00 = 1;
    116: op1_04_inv00 = 1;
    119: op1_04_inv00 = 1;
    121: op1_04_inv00 = 1;
    29: op1_04_inv00 = 1;
    123: op1_04_inv00 = 1;
    124: op1_04_inv00 = 1;
    125: op1_04_inv00 = 1;
    129: op1_04_inv00 = 1;
    131: op1_04_inv00 = 1;
    default: op1_04_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in01 = reg_0615;
    71: op1_04_in01 = reg_0615;
    80: op1_04_in01 = reg_0615;
    55: op1_04_in01 = reg_1095;
    53: op1_04_in01 = reg_0010;
    73: op1_04_in01 = reg_0204;
    86: op1_04_in01 = reg_1367;
    49: op1_04_in01 = reg_0673;
    54: op1_04_in01 = reg_0673;
    61: op1_04_in01 = reg_0669;
    69: op1_04_in01 = reg_0699;
    50: op1_04_in01 = reg_0980;
    68: op1_04_in01 = reg_0376;
    74: op1_04_in01 = reg_0701;
    75: op1_04_in01 = reg_1489;
    87: op1_04_in01 = reg_0328;
    56: op1_04_in01 = reg_1060;
    46: op1_04_in01 = reg_0078;
    60: op1_04_in01 = imem04_in[3:0];
    99: op1_04_in01 = imem04_in[3:0];
    76: op1_04_in01 = imem00_in[11:8];
    120: op1_04_in01 = imem00_in[11:8];
    124: op1_04_in01 = imem00_in[11:8];
    48: op1_04_in01 = reg_0936;
    33: op1_04_in01 = imem07_in[3:0];
    22: op1_04_in01 = imem07_in[3:0];
    57: op1_04_in01 = reg_0165;
    47: op1_04_in01 = reg_0165;
    77: op1_04_in01 = reg_0414;
    70: op1_04_in01 = reg_0896;
    52: op1_04_in01 = reg_0614;
    58: op1_04_in01 = reg_1144;
    78: op1_04_in01 = reg_0294;
    88: op1_04_in01 = imem03_in[15:12];
    51: op1_04_in01 = reg_0634;
    79: op1_04_in01 = reg_0576;
    59: op1_04_in01 = reg_0868;
    28: op1_04_in01 = imem07_in[7:4];
    37: op1_04_in01 = imem07_in[7:4];
    62: op1_04_in01 = reg_0937;
    44: op1_04_in01 = reg_0696;
    81: op1_04_in01 = reg_1517;
    111: op1_04_in01 = reg_1517;
    34: op1_04_in01 = reg_0465;
    63: op1_04_in01 = reg_0616;
    82: op1_04_in01 = reg_1510;
    89: op1_04_in01 = reg_1029;
    83: op1_04_in01 = reg_0115;
    64: op1_04_in01 = reg_0750;
    84: op1_04_in01 = reg_0797;
    40: op1_04_in01 = reg_0139;
    65: op1_04_in01 = reg_0589;
    85: op1_04_in01 = reg_0044;
    90: op1_04_in01 = reg_0638;
    66: op1_04_in01 = reg_0580;
    91: op1_04_in01 = reg_0068;
    42: op1_04_in01 = reg_0396;
    67: op1_04_in01 = reg_0443;
    92: op1_04_in01 = reg_0385;
    93: op1_04_in01 = reg_0966;
    94: op1_04_in01 = reg_0806;
    95: op1_04_in01 = reg_1488;
    96: op1_04_in01 = reg_1099;
    97: op1_04_in01 = reg_0926;
    98: op1_04_in01 = reg_0347;
    100: op1_04_in01 = imem07_in[11:8];
    101: op1_04_in01 = reg_1347;
    102: op1_04_in01 = reg_0363;
    103: op1_04_in01 = reg_0185;
    104: op1_04_in01 = reg_0182;
    105: op1_04_in01 = reg_0319;
    106: op1_04_in01 = imem00_in[7:4];
    107: op1_04_in01 = reg_0882;
    108: op1_04_in01 = reg_0253;
    109: op1_04_in01 = reg_0012;
    110: op1_04_in01 = reg_0998;
    112: op1_04_in01 = reg_1094;
    113: op1_04_in01 = reg_1184;
    38: op1_04_in01 = reg_0413;
    114: op1_04_in01 = reg_1456;
    115: op1_04_in01 = reg_0873;
    116: op1_04_in01 = reg_1202;
    117: op1_04_in01 = reg_0831;
    118: op1_04_in01 = imem06_in[7:4];
    119: op1_04_in01 = reg_0795;
    121: op1_04_in01 = reg_0091;
    122: op1_04_in01 = reg_1001;
    29: op1_04_in01 = reg_0028;
    123: op1_04_in01 = reg_0335;
    125: op1_04_in01 = reg_0130;
    126: op1_04_in01 = reg_0640;
    127: op1_04_in01 = reg_0924;
    128: op1_04_in01 = reg_0394;
    129: op1_04_in01 = reg_0823;
    130: op1_04_in01 = imem05_in[15:12];
    131: op1_04_in01 = reg_0695;
    default: op1_04_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_04_inv01 = 1;
    73: op1_04_inv01 = 1;
    50: op1_04_inv01 = 1;
    71: op1_04_inv01 = 1;
    68: op1_04_inv01 = 1;
    46: op1_04_inv01 = 1;
    48: op1_04_inv01 = 1;
    33: op1_04_inv01 = 1;
    52: op1_04_inv01 = 1;
    58: op1_04_inv01 = 1;
    88: op1_04_inv01 = 1;
    79: op1_04_inv01 = 1;
    62: op1_04_inv01 = 1;
    44: op1_04_inv01 = 1;
    34: op1_04_inv01 = 1;
    63: op1_04_inv01 = 1;
    89: op1_04_inv01 = 1;
    83: op1_04_inv01 = 1;
    84: op1_04_inv01 = 1;
    65: op1_04_inv01 = 1;
    90: op1_04_inv01 = 1;
    66: op1_04_inv01 = 1;
    67: op1_04_inv01 = 1;
    93: op1_04_inv01 = 1;
    94: op1_04_inv01 = 1;
    95: op1_04_inv01 = 1;
    96: op1_04_inv01 = 1;
    97: op1_04_inv01 = 1;
    98: op1_04_inv01 = 1;
    99: op1_04_inv01 = 1;
    100: op1_04_inv01 = 1;
    103: op1_04_inv01 = 1;
    104: op1_04_inv01 = 1;
    105: op1_04_inv01 = 1;
    106: op1_04_inv01 = 1;
    112: op1_04_inv01 = 1;
    113: op1_04_inv01 = 1;
    114: op1_04_inv01 = 1;
    115: op1_04_inv01 = 1;
    117: op1_04_inv01 = 1;
    121: op1_04_inv01 = 1;
    122: op1_04_inv01 = 1;
    123: op1_04_inv01 = 1;
    124: op1_04_inv01 = 1;
    127: op1_04_inv01 = 1;
    130: op1_04_inv01 = 1;
    default: op1_04_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in02 = reg_0748;
    55: op1_04_in02 = reg_1057;
    53: op1_04_in02 = reg_0486;
    73: op1_04_in02 = reg_0251;
    86: op1_04_in02 = imem04_in[11:8];
    67: op1_04_in02 = imem04_in[11:8];
    49: op1_04_in02 = reg_0157;
    61: op1_04_in02 = reg_1278;
    66: op1_04_in02 = reg_1278;
    69: op1_04_in02 = reg_0744;
    54: op1_04_in02 = reg_0158;
    50: op1_04_in02 = reg_0985;
    71: op1_04_in02 = reg_1277;
    68: op1_04_in02 = reg_1139;
    74: op1_04_in02 = reg_1079;
    75: op1_04_in02 = reg_0350;
    87: op1_04_in02 = reg_0233;
    65: op1_04_in02 = reg_0233;
    56: op1_04_in02 = imem07_in[11:8];
    33: op1_04_in02 = imem07_in[11:8];
    46: op1_04_in02 = reg_0079;
    60: op1_04_in02 = imem04_in[15:12];
    76: op1_04_in02 = reg_0983;
    48: op1_04_in02 = reg_0488;
    57: op1_04_in02 = reg_1202;
    77: op1_04_in02 = reg_0598;
    70: op1_04_in02 = reg_0088;
    52: op1_04_in02 = reg_1099;
    58: op1_04_in02 = reg_0535;
    78: op1_04_in02 = reg_0009;
    88: op1_04_in02 = reg_0699;
    51: op1_04_in02 = reg_0635;
    79: op1_04_in02 = reg_0196;
    59: op1_04_in02 = reg_0874;
    28: op1_04_in02 = imem07_in[15:12];
    80: op1_04_in02 = reg_1469;
    96: op1_04_in02 = reg_1469;
    62: op1_04_in02 = reg_0939;
    37: op1_04_in02 = reg_0408;
    44: op1_04_in02 = reg_0420;
    81: op1_04_in02 = reg_0314;
    22: op1_04_in02 = imem07_in[7:4];
    34: op1_04_in02 = imem07_in[3:0];
    63: op1_04_in02 = reg_1078;
    82: op1_04_in02 = reg_0907;
    89: op1_04_in02 = reg_1343;
    83: op1_04_in02 = reg_0717;
    47: op1_04_in02 = reg_0459;
    64: op1_04_in02 = reg_0204;
    84: op1_04_in02 = reg_0206;
    40: op1_04_in02 = reg_0140;
    85: op1_04_in02 = reg_0010;
    90: op1_04_in02 = reg_0804;
    91: op1_04_in02 = reg_0217;
    42: op1_04_in02 = reg_0859;
    92: op1_04_in02 = reg_0162;
    93: op1_04_in02 = reg_0146;
    94: op1_04_in02 = reg_0580;
    95: op1_04_in02 = reg_0205;
    97: op1_04_in02 = reg_0501;
    98: op1_04_in02 = reg_0992;
    99: op1_04_in02 = reg_0577;
    100: op1_04_in02 = reg_1414;
    101: op1_04_in02 = reg_0923;
    102: op1_04_in02 = reg_0400;
    103: op1_04_in02 = reg_1063;
    104: op1_04_in02 = reg_0045;
    105: op1_04_in02 = reg_1101;
    106: op1_04_in02 = reg_0248;
    107: op1_04_in02 = reg_0884;
    108: op1_04_in02 = reg_0824;
    131: op1_04_in02 = reg_0824;
    109: op1_04_in02 = reg_0662;
    110: op1_04_in02 = reg_0893;
    111: op1_04_in02 = reg_1314;
    112: op1_04_in02 = reg_0029;
    113: op1_04_in02 = reg_1231;
    38: op1_04_in02 = reg_0591;
    114: op1_04_in02 = reg_0149;
    115: op1_04_in02 = reg_0492;
    116: op1_04_in02 = reg_0371;
    117: op1_04_in02 = reg_0649;
    118: op1_04_in02 = imem06_in[11:8];
    119: op1_04_in02 = reg_0730;
    120: op1_04_in02 = reg_1470;
    121: op1_04_in02 = reg_0896;
    122: op1_04_in02 = reg_0783;
    29: op1_04_in02 = reg_0229;
    123: op1_04_in02 = reg_0402;
    124: op1_04_in02 = reg_1279;
    125: op1_04_in02 = reg_0575;
    126: op1_04_in02 = reg_1027;
    127: op1_04_in02 = reg_1094;
    128: op1_04_in02 = reg_0003;
    129: op1_04_in02 = reg_0145;
    130: op1_04_in02 = reg_0986;
    default: op1_04_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_04_inv02 = 1;
    86: op1_04_inv02 = 1;
    49: op1_04_inv02 = 1;
    69: op1_04_inv02 = 1;
    54: op1_04_inv02 = 1;
    74: op1_04_inv02 = 1;
    56: op1_04_inv02 = 1;
    46: op1_04_inv02 = 1;
    48: op1_04_inv02 = 1;
    33: op1_04_inv02 = 1;
    52: op1_04_inv02 = 1;
    58: op1_04_inv02 = 1;
    88: op1_04_inv02 = 1;
    51: op1_04_inv02 = 1;
    79: op1_04_inv02 = 1;
    59: op1_04_inv02 = 1;
    62: op1_04_inv02 = 1;
    37: op1_04_inv02 = 1;
    44: op1_04_inv02 = 1;
    81: op1_04_inv02 = 1;
    22: op1_04_inv02 = 1;
    34: op1_04_inv02 = 1;
    63: op1_04_inv02 = 1;
    82: op1_04_inv02 = 1;
    89: op1_04_inv02 = 1;
    47: op1_04_inv02 = 1;
    64: op1_04_inv02 = 1;
    40: op1_04_inv02 = 1;
    67: op1_04_inv02 = 1;
    94: op1_04_inv02 = 1;
    95: op1_04_inv02 = 1;
    96: op1_04_inv02 = 1;
    97: op1_04_inv02 = 1;
    98: op1_04_inv02 = 1;
    100: op1_04_inv02 = 1;
    101: op1_04_inv02 = 1;
    104: op1_04_inv02 = 1;
    105: op1_04_inv02 = 1;
    107: op1_04_inv02 = 1;
    108: op1_04_inv02 = 1;
    110: op1_04_inv02 = 1;
    111: op1_04_inv02 = 1;
    38: op1_04_inv02 = 1;
    117: op1_04_inv02 = 1;
    118: op1_04_inv02 = 1;
    120: op1_04_inv02 = 1;
    122: op1_04_inv02 = 1;
    123: op1_04_inv02 = 1;
    125: op1_04_inv02 = 1;
    126: op1_04_inv02 = 1;
    130: op1_04_inv02 = 1;
    131: op1_04_inv02 = 1;
    default: op1_04_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in03 = reg_1081;
    63: op1_04_in03 = reg_1081;
    55: op1_04_in03 = reg_1055;
    53: op1_04_in03 = reg_0667;
    73: op1_04_in03 = reg_0173;
    86: op1_04_in03 = imem04_in[15:12];
    49: op1_04_in03 = imem07_in[7:4];
    61: op1_04_in03 = reg_1080;
    69: op1_04_in03 = reg_0997;
    54: op1_04_in03 = reg_0774;
    50: op1_04_in03 = reg_0819;
    71: op1_04_in03 = reg_1279;
    105: op1_04_in03 = reg_1279;
    68: op1_04_in03 = reg_0220;
    74: op1_04_in03 = reg_1487;
    97: op1_04_in03 = reg_1487;
    75: op1_04_in03 = reg_0805;
    87: op1_04_in03 = reg_0699;
    56: op1_04_in03 = reg_0703;
    46: op1_04_in03 = reg_0044;
    60: op1_04_in03 = reg_0396;
    76: op1_04_in03 = reg_1277;
    48: op1_04_in03 = reg_0341;
    33: op1_04_in03 = reg_0592;
    57: op1_04_in03 = reg_1179;
    77: op1_04_in03 = reg_0796;
    70: op1_04_in03 = reg_0277;
    52: op1_04_in03 = reg_1078;
    58: op1_04_in03 = reg_0462;
    78: op1_04_in03 = reg_1392;
    88: op1_04_in03 = reg_0185;
    51: op1_04_in03 = reg_0619;
    79: op1_04_in03 = reg_0449;
    59: op1_04_in03 = reg_0042;
    80: op1_04_in03 = reg_1053;
    62: op1_04_in03 = reg_0167;
    37: op1_04_in03 = reg_0618;
    44: op1_04_in03 = reg_0467;
    81: op1_04_in03 = reg_0957;
    22: op1_04_in03 = reg_0004;
    34: op1_04_in03 = reg_0408;
    82: op1_04_in03 = imem00_in[3:0];
    89: op1_04_in03 = reg_0390;
    83: op1_04_in03 = reg_0636;
    47: op1_04_in03 = reg_0269;
    64: op1_04_in03 = reg_0347;
    84: op1_04_in03 = reg_1437;
    40: op1_04_in03 = reg_0031;
    127: op1_04_in03 = reg_0031;
    65: op1_04_in03 = reg_0473;
    85: op1_04_in03 = reg_0013;
    90: op1_04_in03 = reg_0554;
    66: op1_04_in03 = reg_0843;
    91: op1_04_in03 = reg_0255;
    42: op1_04_in03 = reg_0372;
    67: op1_04_in03 = reg_1368;
    92: op1_04_in03 = reg_0290;
    93: op1_04_in03 = reg_0402;
    102: op1_04_in03 = reg_0402;
    94: op1_04_in03 = reg_1454;
    95: op1_04_in03 = reg_0182;
    98: op1_04_in03 = reg_0182;
    96: op1_04_in03 = reg_0926;
    99: op1_04_in03 = reg_0032;
    100: op1_04_in03 = reg_0159;
    101: op1_04_in03 = reg_0286;
    103: op1_04_in03 = reg_1001;
    104: op1_04_in03 = reg_0564;
    106: op1_04_in03 = reg_0866;
    107: op1_04_in03 = reg_1149;
    108: op1_04_in03 = reg_0069;
    109: op1_04_in03 = reg_0877;
    110: op1_04_in03 = reg_0498;
    111: op1_04_in03 = reg_1199;
    112: op1_04_in03 = reg_0665;
    113: op1_04_in03 = reg_0178;
    38: op1_04_in03 = reg_0051;
    114: op1_04_in03 = reg_0148;
    115: op1_04_in03 = reg_0275;
    116: op1_04_in03 = reg_0977;
    117: op1_04_in03 = reg_0604;
    118: op1_04_in03 = reg_1036;
    119: op1_04_in03 = reg_1420;
    120: op1_04_in03 = reg_0248;
    121: op1_04_in03 = reg_0403;
    122: op1_04_in03 = reg_0191;
    29: op1_04_in03 = reg_0219;
    123: op1_04_in03 = reg_0010;
    124: op1_04_in03 = reg_0748;
    125: op1_04_in03 = reg_1346;
    126: op1_04_in03 = reg_1459;
    128: op1_04_in03 = reg_0993;
    129: op1_04_in03 = reg_0556;
    130: op1_04_in03 = reg_0251;
    131: op1_04_in03 = reg_0848;
    default: op1_04_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv03 = 1;
    55: op1_04_inv03 = 1;
    86: op1_04_inv03 = 1;
    61: op1_04_inv03 = 1;
    50: op1_04_inv03 = 1;
    74: op1_04_inv03 = 1;
    75: op1_04_inv03 = 1;
    56: op1_04_inv03 = 1;
    46: op1_04_inv03 = 1;
    60: op1_04_inv03 = 1;
    76: op1_04_inv03 = 1;
    70: op1_04_inv03 = 1;
    58: op1_04_inv03 = 1;
    78: op1_04_inv03 = 1;
    80: op1_04_inv03 = 1;
    37: op1_04_inv03 = 1;
    44: op1_04_inv03 = 1;
    81: op1_04_inv03 = 1;
    22: op1_04_inv03 = 1;
    34: op1_04_inv03 = 1;
    82: op1_04_inv03 = 1;
    83: op1_04_inv03 = 1;
    47: op1_04_inv03 = 1;
    65: op1_04_inv03 = 1;
    85: op1_04_inv03 = 1;
    42: op1_04_inv03 = 1;
    67: op1_04_inv03 = 1;
    94: op1_04_inv03 = 1;
    97: op1_04_inv03 = 1;
    98: op1_04_inv03 = 1;
    99: op1_04_inv03 = 1;
    100: op1_04_inv03 = 1;
    101: op1_04_inv03 = 1;
    102: op1_04_inv03 = 1;
    104: op1_04_inv03 = 1;
    107: op1_04_inv03 = 1;
    108: op1_04_inv03 = 1;
    110: op1_04_inv03 = 1;
    111: op1_04_inv03 = 1;
    112: op1_04_inv03 = 1;
    113: op1_04_inv03 = 1;
    114: op1_04_inv03 = 1;
    117: op1_04_inv03 = 1;
    119: op1_04_inv03 = 1;
    122: op1_04_inv03 = 1;
    29: op1_04_inv03 = 1;
    126: op1_04_inv03 = 1;
    127: op1_04_inv03 = 1;
    128: op1_04_inv03 = 1;
    129: op1_04_inv03 = 1;
    130: op1_04_inv03 = 1;
    default: op1_04_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in04 = imem00_in[7:4];
    82: op1_04_in04 = imem00_in[7:4];
    55: op1_04_in04 = imem07_in[3:0];
    53: op1_04_in04 = reg_0668;
    73: op1_04_in04 = reg_0646;
    86: op1_04_in04 = reg_1198;
    49: op1_04_in04 = imem07_in[15:12];
    61: op1_04_in04 = reg_0293;
    69: op1_04_in04 = reg_0976;
    54: op1_04_in04 = reg_0030;
    50: op1_04_in04 = reg_0430;
    71: op1_04_in04 = reg_1242;
    68: op1_04_in04 = reg_0505;
    74: op1_04_in04 = reg_0552;
    75: op1_04_in04 = reg_1470;
    87: op1_04_in04 = reg_0710;
    56: op1_04_in04 = reg_0704;
    46: op1_04_in04 = reg_0011;
    60: op1_04_in04 = reg_0263;
    76: op1_04_in04 = reg_1490;
    48: op1_04_in04 = reg_0262;
    33: op1_04_in04 = reg_0102;
    57: op1_04_in04 = reg_0269;
    77: op1_04_in04 = reg_0033;
    70: op1_04_in04 = reg_0044;
    52: op1_04_in04 = reg_0841;
    58: op1_04_in04 = reg_1077;
    78: op1_04_in04 = reg_0695;
    88: op1_04_in04 = reg_0330;
    51: op1_04_in04 = reg_0419;
    79: op1_04_in04 = reg_0828;
    59: op1_04_in04 = reg_0041;
    80: op1_04_in04 = reg_1027;
    62: op1_04_in04 = reg_0872;
    37: op1_04_in04 = reg_0593;
    44: op1_04_in04 = reg_0412;
    81: op1_04_in04 = reg_0048;
    22: op1_04_in04 = reg_0050;
    34: op1_04_in04 = reg_0003;
    63: op1_04_in04 = reg_0806;
    89: op1_04_in04 = imem02_in[7:4];
    83: op1_04_in04 = reg_0374;
    47: op1_04_in04 = reg_0152;
    64: op1_04_in04 = reg_1164;
    84: op1_04_in04 = reg_1435;
    40: op1_04_in04 = reg_0465;
    65: op1_04_in04 = reg_0475;
    85: op1_04_in04 = reg_0895;
    90: op1_04_in04 = reg_0555;
    66: op1_04_in04 = reg_0804;
    97: op1_04_in04 = reg_0804;
    91: op1_04_in04 = reg_0999;
    42: op1_04_in04 = reg_0636;
    67: op1_04_in04 = reg_0252;
    92: op1_04_in04 = reg_0447;
    93: op1_04_in04 = reg_0401;
    94: op1_04_in04 = reg_1459;
    95: op1_04_in04 = reg_1181;
    96: op1_04_in04 = reg_1278;
    98: op1_04_in04 = reg_1403;
    99: op1_04_in04 = reg_1369;
    100: op1_04_in04 = reg_0031;
    101: op1_04_in04 = reg_0437;
    102: op1_04_in04 = reg_1071;
    103: op1_04_in04 = reg_0311;
    104: op1_04_in04 = reg_1070;
    105: op1_04_in04 = reg_0640;
    106: op1_04_in04 = reg_1277;
    107: op1_04_in04 = reg_1009;
    108: op1_04_in04 = reg_1515;
    109: op1_04_in04 = reg_0879;
    110: op1_04_in04 = reg_1010;
    111: op1_04_in04 = reg_0178;
    112: op1_04_in04 = reg_0366;
    113: op1_04_in04 = reg_0107;
    38: op1_04_in04 = reg_0483;
    114: op1_04_in04 = reg_0146;
    115: op1_04_in04 = reg_0243;
    116: op1_04_in04 = reg_0067;
    117: op1_04_in04 = reg_0701;
    118: op1_04_in04 = reg_0905;
    119: op1_04_in04 = reg_1326;
    120: op1_04_in04 = reg_1081;
    121: op1_04_in04 = reg_0634;
    122: op1_04_in04 = reg_0180;
    29: op1_04_in04 = reg_0186;
    123: op1_04_in04 = reg_1068;
    124: op1_04_in04 = reg_1141;
    125: op1_04_in04 = imem06_in[7:4];
    126: op1_04_in04 = reg_0249;
    127: op1_04_in04 = reg_0664;
    128: op1_04_in04 = reg_0994;
    129: op1_04_in04 = reg_0965;
    130: op1_04_in04 = reg_0996;
    131: op1_04_in04 = reg_1078;
    default: op1_04_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv04 = 1;
    55: op1_04_inv04 = 1;
    53: op1_04_inv04 = 1;
    73: op1_04_inv04 = 1;
    86: op1_04_inv04 = 1;
    49: op1_04_inv04 = 1;
    61: op1_04_inv04 = 1;
    50: op1_04_inv04 = 1;
    74: op1_04_inv04 = 1;
    46: op1_04_inv04 = 1;
    60: op1_04_inv04 = 1;
    76: op1_04_inv04 = 1;
    78: op1_04_inv04 = 1;
    80: op1_04_inv04 = 1;
    44: op1_04_inv04 = 1;
    22: op1_04_inv04 = 1;
    34: op1_04_inv04 = 1;
    63: op1_04_inv04 = 1;
    47: op1_04_inv04 = 1;
    64: op1_04_inv04 = 1;
    84: op1_04_inv04 = 1;
    65: op1_04_inv04 = 1;
    91: op1_04_inv04 = 1;
    42: op1_04_inv04 = 1;
    95: op1_04_inv04 = 1;
    96: op1_04_inv04 = 1;
    99: op1_04_inv04 = 1;
    103: op1_04_inv04 = 1;
    105: op1_04_inv04 = 1;
    107: op1_04_inv04 = 1;
    109: op1_04_inv04 = 1;
    110: op1_04_inv04 = 1;
    111: op1_04_inv04 = 1;
    112: op1_04_inv04 = 1;
    38: op1_04_inv04 = 1;
    116: op1_04_inv04 = 1;
    117: op1_04_inv04 = 1;
    118: op1_04_inv04 = 1;
    120: op1_04_inv04 = 1;
    121: op1_04_inv04 = 1;
    122: op1_04_inv04 = 1;
    29: op1_04_inv04 = 1;
    125: op1_04_inv04 = 1;
    127: op1_04_inv04 = 1;
    129: op1_04_inv04 = 1;
    default: op1_04_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in05 = imem00_in[15:12];
    55: op1_04_in05 = reg_0245;
    53: op1_04_in05 = reg_1098;
    73: op1_04_in05 = reg_0333;
    86: op1_04_in05 = reg_1082;
    49: op1_04_in05 = reg_0139;
    61: op1_04_in05 = reg_1230;
    69: op1_04_in05 = reg_0533;
    102: op1_04_in05 = reg_0533;
    54: op1_04_in05 = reg_0663;
    50: op1_04_in05 = reg_0930;
    71: op1_04_in05 = reg_0804;
    63: op1_04_in05 = reg_0804;
    68: op1_04_in05 = reg_0506;
    74: op1_04_in05 = reg_0806;
    75: op1_04_in05 = reg_1053;
    87: op1_04_in05 = reg_1001;
    56: op1_04_in05 = reg_0892;
    46: op1_04_in05 = reg_0010;
    70: op1_04_in05 = reg_0010;
    60: op1_04_in05 = reg_0462;
    76: op1_04_in05 = reg_0350;
    48: op1_04_in05 = reg_0487;
    33: op1_04_in05 = reg_0051;
    57: op1_04_in05 = reg_0271;
    77: op1_04_in05 = reg_0061;
    52: op1_04_in05 = reg_1052;
    58: op1_04_in05 = reg_1083;
    78: op1_04_in05 = reg_0632;
    88: op1_04_in05 = reg_1448;
    51: op1_04_in05 = reg_0067;
    79: op1_04_in05 = reg_0206;
    59: op1_04_in05 = reg_0011;
    80: op1_04_in05 = reg_1453;
    62: op1_04_in05 = reg_0196;
    37: op1_04_in05 = reg_0028;
    44: op1_04_in05 = reg_0837;
    81: op1_04_in05 = reg_1231;
    22: op1_04_in05 = reg_0053;
    34: op1_04_in05 = reg_0518;
    82: op1_04_in05 = reg_0613;
    89: op1_04_in05 = reg_0128;
    83: op1_04_in05 = reg_0373;
    47: op1_04_in05 = reg_0212;
    64: op1_04_in05 = reg_1212;
    84: op1_04_in05 = reg_0795;
    40: op1_04_in05 = reg_0366;
    127: op1_04_in05 = reg_0366;
    65: op1_04_in05 = reg_0436;
    85: op1_04_in05 = reg_0332;
    90: op1_04_in05 = reg_0987;
    66: op1_04_in05 = reg_0523;
    91: op1_04_in05 = reg_0154;
    42: op1_04_in05 = reg_0637;
    67: op1_04_in05 = reg_1257;
    92: op1_04_in05 = reg_0590;
    93: op1_04_in05 = reg_0360;
    94: op1_04_in05 = reg_0961;
    126: op1_04_in05 = reg_0961;
    95: op1_04_in05 = reg_1401;
    96: op1_04_in05 = reg_1487;
    97: op1_04_in05 = reg_0805;
    98: op1_04_in05 = reg_0940;
    99: op1_04_in05 = reg_0731;
    100: op1_04_in05 = reg_0284;
    101: op1_04_in05 = reg_0404;
    103: op1_04_in05 = reg_0000;
    104: op1_04_in05 = reg_1169;
    105: op1_04_in05 = reg_0250;
    106: op1_04_in05 = reg_1279;
    107: op1_04_in05 = reg_0025;
    108: op1_04_in05 = imem03_in[15:12];
    109: op1_04_in05 = reg_0276;
    110: op1_04_in05 = reg_0461;
    111: op1_04_in05 = reg_1139;
    112: op1_04_in05 = reg_0415;
    113: op1_04_in05 = reg_0113;
    114: op1_04_in05 = reg_0868;
    115: op1_04_in05 = reg_1346;
    116: op1_04_in05 = reg_0018;
    117: op1_04_in05 = reg_0045;
    118: op1_04_in05 = reg_0870;
    119: op1_04_in05 = reg_1508;
    120: op1_04_in05 = reg_0638;
    121: op1_04_in05 = reg_0041;
    122: op1_04_in05 = reg_0375;
    29: op1_04_in05 = reg_0003;
    123: op1_04_in05 = imem02_in[15:12];
    124: op1_04_in05 = reg_0501;
    125: op1_04_in05 = reg_0753;
    128: op1_04_in05 = reg_1060;
    129: op1_04_in05 = reg_0349;
    130: op1_04_in05 = reg_0793;
    131: op1_04_in05 = reg_1091;
    default: op1_04_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_04_inv05 = 1;
    53: op1_04_inv05 = 1;
    73: op1_04_inv05 = 1;
    86: op1_04_inv05 = 1;
    61: op1_04_inv05 = 1;
    69: op1_04_inv05 = 1;
    50: op1_04_inv05 = 1;
    74: op1_04_inv05 = 1;
    75: op1_04_inv05 = 1;
    56: op1_04_inv05 = 1;
    57: op1_04_inv05 = 1;
    77: op1_04_inv05 = 1;
    70: op1_04_inv05 = 1;
    58: op1_04_inv05 = 1;
    78: op1_04_inv05 = 1;
    88: op1_04_inv05 = 1;
    79: op1_04_inv05 = 1;
    59: op1_04_inv05 = 1;
    62: op1_04_inv05 = 1;
    44: op1_04_inv05 = 1;
    34: op1_04_inv05 = 1;
    82: op1_04_inv05 = 1;
    47: op1_04_inv05 = 1;
    84: op1_04_inv05 = 1;
    65: op1_04_inv05 = 1;
    85: op1_04_inv05 = 1;
    91: op1_04_inv05 = 1;
    67: op1_04_inv05 = 1;
    92: op1_04_inv05 = 1;
    93: op1_04_inv05 = 1;
    94: op1_04_inv05 = 1;
    96: op1_04_inv05 = 1;
    98: op1_04_inv05 = 1;
    99: op1_04_inv05 = 1;
    100: op1_04_inv05 = 1;
    102: op1_04_inv05 = 1;
    103: op1_04_inv05 = 1;
    107: op1_04_inv05 = 1;
    108: op1_04_inv05 = 1;
    109: op1_04_inv05 = 1;
    110: op1_04_inv05 = 1;
    111: op1_04_inv05 = 1;
    116: op1_04_inv05 = 1;
    118: op1_04_inv05 = 1;
    121: op1_04_inv05 = 1;
    123: op1_04_inv05 = 1;
    124: op1_04_inv05 = 1;
    125: op1_04_inv05 = 1;
    127: op1_04_inv05 = 1;
    128: op1_04_inv05 = 1;
    130: op1_04_inv05 = 1;
    default: op1_04_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in06 = reg_0804;
    124: op1_04_in06 = reg_0804;
    55: op1_04_in06 = reg_0867;
    56: op1_04_in06 = reg_0867;
    53: op1_04_in06 = reg_0133;
    73: op1_04_in06 = reg_0131;
    86: op1_04_in06 = reg_1147;
    49: op1_04_in06 = reg_0140;
    61: op1_04_in06 = reg_1206;
    69: op1_04_in06 = reg_1018;
    54: op1_04_in06 = reg_0413;
    101: op1_04_in06 = reg_0413;
    50: op1_04_in06 = reg_0149;
    71: op1_04_in06 = reg_0803;
    74: op1_04_in06 = reg_0803;
    63: op1_04_in06 = reg_0803;
    68: op1_04_in06 = reg_0481;
    75: op1_04_in06 = reg_1027;
    52: op1_04_in06 = reg_1027;
    66: op1_04_in06 = reg_1027;
    105: op1_04_in06 = reg_1027;
    87: op1_04_in06 = reg_0707;
    46: op1_04_in06 = reg_0013;
    59: op1_04_in06 = reg_0013;
    60: op1_04_in06 = reg_1214;
    76: op1_04_in06 = reg_0805;
    48: op1_04_in06 = reg_0368;
    33: op1_04_in06 = reg_0084;
    57: op1_04_in06 = reg_0023;
    77: op1_04_in06 = reg_0304;
    70: op1_04_in06 = reg_1140;
    58: op1_04_in06 = reg_0904;
    78: op1_04_in06 = reg_0801;
    88: op1_04_in06 = reg_0177;
    51: op1_04_in06 = reg_0152;
    79: op1_04_in06 = reg_0037;
    80: op1_04_in06 = reg_0987;
    62: op1_04_in06 = reg_0864;
    37: op1_04_in06 = reg_0050;
    44: op1_04_in06 = reg_0094;
    81: op1_04_in06 = reg_0885;
    82: op1_04_in06 = reg_0250;
    89: op1_04_in06 = reg_0112;
    83: op1_04_in06 = reg_0586;
    119: op1_04_in06 = reg_0586;
    47: op1_04_in06 = reg_0215;
    64: op1_04_in06 = reg_0318;
    84: op1_04_in06 = reg_0906;
    40: op1_04_in06 = reg_0100;
    65: op1_04_in06 = reg_0778;
    85: op1_04_in06 = reg_0530;
    90: op1_04_in06 = reg_0961;
    91: op1_04_in06 = reg_0573;
    42: op1_04_in06 = reg_0617;
    67: op1_04_in06 = reg_1216;
    92: op1_04_in06 = reg_0824;
    93: op1_04_in06 = reg_0363;
    94: op1_04_in06 = reg_0155;
    95: op1_04_in06 = reg_0938;
    98: op1_04_in06 = reg_0938;
    96: op1_04_in06 = reg_1053;
    97: op1_04_in06 = reg_0523;
    99: op1_04_in06 = reg_1083;
    100: op1_04_in06 = reg_0415;
    102: op1_04_in06 = reg_0499;
    103: op1_04_in06 = reg_0789;
    104: op1_04_in06 = reg_1514;
    106: op1_04_in06 = reg_0501;
    107: op1_04_in06 = reg_0790;
    108: op1_04_in06 = reg_0328;
    109: op1_04_in06 = reg_0561;
    110: op1_04_in06 = reg_1415;
    111: op1_04_in06 = reg_1280;
    112: op1_04_in06 = reg_0593;
    113: op1_04_in06 = reg_0104;
    114: op1_04_in06 = reg_1511;
    115: op1_04_in06 = reg_0589;
    116: op1_04_in06 = imem07_in[7:4];
    117: op1_04_in06 = reg_0167;
    118: op1_04_in06 = reg_1209;
    120: op1_04_in06 = reg_0843;
    121: op1_04_in06 = reg_0012;
    122: op1_04_in06 = reg_1184;
    29: op1_04_in06 = imem07_in[15:12];
    123: op1_04_in06 = reg_0475;
    125: op1_04_in06 = reg_0264;
    126: op1_04_in06 = reg_1432;
    127: op1_04_in06 = reg_0437;
    128: op1_04_in06 = reg_0298;
    129: op1_04_in06 = reg_0962;
    130: op1_04_in06 = reg_0391;
    131: op1_04_in06 = reg_0227;
    default: op1_04_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv06 = 1;
    55: op1_04_inv06 = 1;
    53: op1_04_inv06 = 1;
    86: op1_04_inv06 = 1;
    49: op1_04_inv06 = 1;
    61: op1_04_inv06 = 1;
    69: op1_04_inv06 = 1;
    54: op1_04_inv06 = 1;
    50: op1_04_inv06 = 1;
    71: op1_04_inv06 = 1;
    68: op1_04_inv06 = 1;
    87: op1_04_inv06 = 1;
    56: op1_04_inv06 = 1;
    60: op1_04_inv06 = 1;
    76: op1_04_inv06 = 1;
    48: op1_04_inv06 = 1;
    33: op1_04_inv06 = 1;
    57: op1_04_inv06 = 1;
    77: op1_04_inv06 = 1;
    70: op1_04_inv06 = 1;
    78: op1_04_inv06 = 1;
    47: op1_04_inv06 = 1;
    84: op1_04_inv06 = 1;
    40: op1_04_inv06 = 1;
    90: op1_04_inv06 = 1;
    91: op1_04_inv06 = 1;
    42: op1_04_inv06 = 1;
    67: op1_04_inv06 = 1;
    92: op1_04_inv06 = 1;
    94: op1_04_inv06 = 1;
    97: op1_04_inv06 = 1;
    98: op1_04_inv06 = 1;
    99: op1_04_inv06 = 1;
    100: op1_04_inv06 = 1;
    101: op1_04_inv06 = 1;
    102: op1_04_inv06 = 1;
    103: op1_04_inv06 = 1;
    104: op1_04_inv06 = 1;
    106: op1_04_inv06 = 1;
    108: op1_04_inv06 = 1;
    109: op1_04_inv06 = 1;
    112: op1_04_inv06 = 1;
    113: op1_04_inv06 = 1;
    114: op1_04_inv06 = 1;
    119: op1_04_inv06 = 1;
    122: op1_04_inv06 = 1;
    124: op1_04_inv06 = 1;
    126: op1_04_inv06 = 1;
    130: op1_04_inv06 = 1;
    default: op1_04_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in07 = reg_0218;
    74: op1_04_in07 = reg_0218;
    55: op1_04_in07 = reg_0489;
    53: op1_04_in07 = reg_0922;
    73: op1_04_in07 = reg_1181;
    86: op1_04_in07 = reg_0421;
    49: op1_04_in07 = reg_0777;
    61: op1_04_in07 = reg_0725;
    69: op1_04_in07 = reg_0475;
    54: op1_04_in07 = reg_0621;
    50: op1_04_in07 = reg_0146;
    71: op1_04_in07 = imem00_in[15:12];
    68: op1_04_in07 = imem03_in[11:8];
    75: op1_04_in07 = reg_1454;
    87: op1_04_in07 = reg_0143;
    56: op1_04_in07 = reg_0298;
    46: op1_04_in07 = reg_0254;
    60: op1_04_in07 = reg_1203;
    67: op1_04_in07 = reg_1203;
    76: op1_04_in07 = reg_0523;
    48: op1_04_in07 = reg_0836;
    33: op1_04_in07 = reg_0087;
    57: op1_04_in07 = reg_0214;
    77: op1_04_in07 = reg_0262;
    70: op1_04_in07 = reg_0399;
    52: op1_04_in07 = reg_0249;
    58: op1_04_in07 = reg_0719;
    78: op1_04_in07 = reg_0800;
    88: op1_04_in07 = reg_0180;
    51: op1_04_in07 = reg_0215;
    79: op1_04_in07 = reg_0038;
    59: op1_04_in07 = reg_1103;
    80: op1_04_in07 = reg_0460;
    62: op1_04_in07 = imem05_in[15:12];
    37: op1_04_in07 = reg_0004;
    44: op1_04_in07 = reg_0096;
    81: op1_04_in07 = reg_0882;
    63: op1_04_in07 = reg_1052;
    82: op1_04_in07 = reg_0987;
    89: op1_04_in07 = reg_1433;
    83: op1_04_in07 = reg_0619;
    47: op1_04_in07 = reg_0213;
    64: op1_04_in07 = reg_0450;
    84: op1_04_in07 = reg_0905;
    40: op1_04_in07 = reg_0051;
    65: op1_04_in07 = reg_0973;
    85: op1_04_in07 = reg_0138;
    90: op1_04_in07 = reg_1432;
    96: op1_04_in07 = reg_1432;
    66: op1_04_in07 = reg_0155;
    91: op1_04_in07 = reg_0709;
    42: op1_04_in07 = reg_0585;
    92: op1_04_in07 = imem02_in[3:0];
    93: op1_04_in07 = reg_0292;
    94: op1_04_in07 = reg_0524;
    95: op1_04_in07 = reg_0418;
    97: op1_04_in07 = reg_1459;
    98: op1_04_in07 = reg_0937;
    99: op1_04_in07 = reg_1215;
    100: op1_04_in07 = reg_0618;
    101: op1_04_in07 = reg_0100;
    102: op1_04_in07 = reg_0668;
    103: op1_04_in07 = reg_1495;
    104: op1_04_in07 = reg_0873;
    105: op1_04_in07 = reg_0887;
    106: op1_04_in07 = reg_0804;
    120: op1_04_in07 = reg_0804;
    107: op1_04_in07 = reg_1280;
    108: op1_04_in07 = reg_0177;
    109: op1_04_in07 = reg_0532;
    110: op1_04_in07 = reg_0994;
    111: op1_04_in07 = reg_1339;
    112: op1_04_in07 = reg_0137;
    113: op1_04_in07 = reg_0880;
    114: op1_04_in07 = reg_0360;
    115: op1_04_in07 = reg_0864;
    116: op1_04_in07 = reg_1010;
    117: op1_04_in07 = reg_0334;
    118: op1_04_in07 = reg_0960;
    119: op1_04_in07 = reg_0571;
    121: op1_04_in07 = reg_1071;
    122: op1_04_in07 = reg_0070;
    29: op1_04_in07 = reg_0484;
    123: op1_04_in07 = reg_0889;
    124: op1_04_in07 = reg_0613;
    125: op1_04_in07 = reg_0929;
    126: op1_04_in07 = reg_0229;
    127: op1_04_in07 = reg_0623;
    128: op1_04_in07 = reg_1056;
    129: op1_04_in07 = reg_0178;
    130: op1_04_in07 = reg_0701;
    131: op1_04_in07 = reg_0563;
    default: op1_04_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_04_inv07 = 1;
    49: op1_04_inv07 = 1;
    69: op1_04_inv07 = 1;
    50: op1_04_inv07 = 1;
    71: op1_04_inv07 = 1;
    75: op1_04_inv07 = 1;
    87: op1_04_inv07 = 1;
    46: op1_04_inv07 = 1;
    60: op1_04_inv07 = 1;
    48: op1_04_inv07 = 1;
    77: op1_04_inv07 = 1;
    88: op1_04_inv07 = 1;
    51: op1_04_inv07 = 1;
    62: op1_04_inv07 = 1;
    37: op1_04_inv07 = 1;
    44: op1_04_inv07 = 1;
    81: op1_04_inv07 = 1;
    89: op1_04_inv07 = 1;
    83: op1_04_inv07 = 1;
    47: op1_04_inv07 = 1;
    64: op1_04_inv07 = 1;
    66: op1_04_inv07 = 1;
    91: op1_04_inv07 = 1;
    42: op1_04_inv07 = 1;
    92: op1_04_inv07 = 1;
    93: op1_04_inv07 = 1;
    94: op1_04_inv07 = 1;
    95: op1_04_inv07 = 1;
    98: op1_04_inv07 = 1;
    99: op1_04_inv07 = 1;
    101: op1_04_inv07 = 1;
    102: op1_04_inv07 = 1;
    105: op1_04_inv07 = 1;
    113: op1_04_inv07 = 1;
    115: op1_04_inv07 = 1;
    116: op1_04_inv07 = 1;
    117: op1_04_inv07 = 1;
    118: op1_04_inv07 = 1;
    119: op1_04_inv07 = 1;
    120: op1_04_inv07 = 1;
    121: op1_04_inv07 = 1;
    122: op1_04_inv07 = 1;
    29: op1_04_inv07 = 1;
    123: op1_04_inv07 = 1;
    126: op1_04_inv07 = 1;
    127: op1_04_inv07 = 1;
    128: op1_04_inv07 = 1;
    129: op1_04_inv07 = 1;
    130: op1_04_inv07 = 1;
    131: op1_04_inv07 = 1;
    default: op1_04_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in08 = reg_0250;
    55: op1_04_in08 = reg_0442;
    53: op1_04_in08 = reg_1029;
    73: op1_04_in08 = reg_1402;
    86: op1_04_in08 = reg_0471;
    49: op1_04_in08 = reg_0774;
    61: op1_04_in08 = reg_0641;
    69: op1_04_in08 = reg_0474;
    54: op1_04_in08 = reg_0618;
    50: op1_04_in08 = reg_0365;
    71: op1_04_in08 = reg_0353;
    68: op1_04_in08 = reg_0790;
    74: op1_04_in08 = reg_0221;
    75: op1_04_in08 = reg_1459;
    87: op1_04_in08 = reg_0891;
    56: op1_04_in08 = reg_0157;
    46: op1_04_in08 = reg_0631;
    60: op1_04_in08 = reg_0420;
    76: op1_04_in08 = reg_0293;
    48: op1_04_in08 = reg_0336;
    33: op1_04_in08 = reg_0521;
    57: op1_04_in08 = reg_0017;
    77: op1_04_in08 = reg_0097;
    70: op1_04_in08 = reg_0563;
    52: op1_04_in08 = reg_0203;
    58: op1_04_in08 = reg_0236;
    78: op1_04_in08 = reg_0281;
    88: op1_04_in08 = reg_0142;
    51: op1_04_in08 = reg_0018;
    79: op1_04_in08 = reg_0261;
    59: op1_04_in08 = reg_0607;
    80: op1_04_in08 = reg_0887;
    62: op1_04_in08 = reg_1035;
    37: op1_04_in08 = reg_0052;
    44: op1_04_in08 = reg_0237;
    81: op1_04_in08 = reg_0479;
    63: op1_04_in08 = reg_1201;
    82: op1_04_in08 = reg_1417;
    126: op1_04_in08 = reg_1417;
    89: op1_04_in08 = reg_1031;
    83: op1_04_in08 = reg_0132;
    47: op1_04_in08 = reg_0015;
    64: op1_04_in08 = reg_0300;
    95: op1_04_in08 = reg_0300;
    84: op1_04_in08 = reg_1426;
    40: op1_04_in08 = reg_0004;
    65: op1_04_in08 = reg_0935;
    85: op1_04_in08 = reg_0276;
    90: op1_04_in08 = reg_0524;
    66: op1_04_in08 = reg_0459;
    91: op1_04_in08 = reg_0330;
    42: op1_04_in08 = reg_0529;
    67: op1_04_in08 = reg_1198;
    92: op1_04_in08 = reg_0530;
    93: op1_04_in08 = reg_0724;
    94: op1_04_in08 = reg_0881;
    96: op1_04_in08 = reg_0476;
    97: op1_04_in08 = reg_0249;
    98: op1_04_in08 = reg_0090;
    99: op1_04_in08 = reg_0796;
    100: op1_04_in08 = reg_0001;
    101: op1_04_in08 = reg_0028;
    102: op1_04_in08 = reg_1235;
    103: op1_04_in08 = reg_0070;
    104: op1_04_in08 = reg_0601;
    105: op1_04_in08 = reg_0886;
    106: op1_04_in08 = reg_0580;
    107: op1_04_in08 = reg_0348;
    108: op1_04_in08 = reg_0312;
    109: op1_04_in08 = reg_0436;
    110: op1_04_in08 = reg_0894;
    111: op1_04_in08 = reg_0467;
    112: op1_04_in08 = reg_0102;
    113: op1_04_in08 = reg_0541;
    114: op1_04_in08 = reg_0901;
    115: op1_04_in08 = reg_0828;
    116: op1_04_in08 = reg_0892;
    117: op1_04_in08 = reg_0697;
    118: op1_04_in08 = reg_0316;
    119: op1_04_in08 = reg_0570;
    120: op1_04_in08 = reg_0841;
    121: op1_04_in08 = imem02_in[11:8];
    122: op1_04_in08 = reg_1518;
    123: op1_04_in08 = reg_0322;
    124: op1_04_in08 = reg_0961;
    125: op1_04_in08 = reg_0192;
    127: op1_04_in08 = reg_0591;
    128: op1_04_in08 = reg_0140;
    129: op1_04_in08 = reg_0291;
    130: op1_04_in08 = reg_0045;
    131: op1_04_in08 = imem03_in[11:8];
    default: op1_04_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv08 = 1;
    53: op1_04_inv08 = 1;
    73: op1_04_inv08 = 1;
    49: op1_04_inv08 = 1;
    54: op1_04_inv08 = 1;
    50: op1_04_inv08 = 1;
    74: op1_04_inv08 = 1;
    87: op1_04_inv08 = 1;
    60: op1_04_inv08 = 1;
    76: op1_04_inv08 = 1;
    33: op1_04_inv08 = 1;
    77: op1_04_inv08 = 1;
    52: op1_04_inv08 = 1;
    79: op1_04_inv08 = 1;
    62: op1_04_inv08 = 1;
    81: op1_04_inv08 = 1;
    63: op1_04_inv08 = 1;
    40: op1_04_inv08 = 1;
    91: op1_04_inv08 = 1;
    67: op1_04_inv08 = 1;
    95: op1_04_inv08 = 1;
    97: op1_04_inv08 = 1;
    98: op1_04_inv08 = 1;
    102: op1_04_inv08 = 1;
    105: op1_04_inv08 = 1;
    106: op1_04_inv08 = 1;
    107: op1_04_inv08 = 1;
    110: op1_04_inv08 = 1;
    111: op1_04_inv08 = 1;
    114: op1_04_inv08 = 1;
    115: op1_04_inv08 = 1;
    116: op1_04_inv08 = 1;
    121: op1_04_inv08 = 1;
    123: op1_04_inv08 = 1;
    124: op1_04_inv08 = 1;
    127: op1_04_inv08 = 1;
    128: op1_04_inv08 = 1;
    129: op1_04_inv08 = 1;
    131: op1_04_inv08 = 1;
    default: op1_04_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in09 = reg_1027;
    55: op1_04_in09 = reg_0103;
    53: op1_04_in09 = reg_0562;
    73: op1_04_in09 = reg_0873;
    86: op1_04_in09 = reg_0451;
    49: op1_04_in09 = reg_0029;
    61: op1_04_in09 = reg_0638;
    69: op1_04_in09 = reg_0472;
    54: op1_04_in09 = reg_0100;
    50: op1_04_in09 = reg_0047;
    71: op1_04_in09 = reg_0005;
    68: op1_04_in09 = reg_1280;
    129: op1_04_in09 = reg_1280;
    74: op1_04_in09 = reg_1201;
    75: op1_04_in09 = reg_1406;
    87: op1_04_in09 = reg_1314;
    122: op1_04_in09 = reg_1314;
    56: op1_04_in09 = reg_0489;
    46: op1_04_in09 = reg_0563;
    60: op1_04_in09 = reg_0414;
    76: op1_04_in09 = reg_1227;
    48: op1_04_in09 = reg_0097;
    33: op1_04_in09 = reg_0123;
    57: op1_04_in09 = reg_1170;
    77: op1_04_in09 = reg_1502;
    70: op1_04_in09 = reg_0233;
    52: op1_04_in09 = reg_0958;
    63: op1_04_in09 = reg_0958;
    66: op1_04_in09 = reg_0958;
    58: op1_04_in09 = reg_0181;
    81: op1_04_in09 = reg_0181;
    78: op1_04_in09 = reg_1515;
    88: op1_04_in09 = reg_0314;
    51: op1_04_in09 = reg_0191;
    79: op1_04_in09 = reg_0906;
    59: op1_04_in09 = reg_0253;
    80: op1_04_in09 = reg_0202;
    90: op1_04_in09 = reg_0202;
    62: op1_04_in09 = reg_0780;
    44: op1_04_in09 = reg_0211;
    82: op1_04_in09 = reg_1418;
    126: op1_04_in09 = reg_1418;
    89: op1_04_in09 = reg_0802;
    83: op1_04_in09 = reg_0046;
    47: op1_04_in09 = reg_0017;
    64: op1_04_in09 = reg_0301;
    95: op1_04_in09 = reg_0301;
    84: op1_04_in09 = reg_1420;
    40: op1_04_in09 = reg_0520;
    65: op1_04_in09 = reg_0106;
    85: op1_04_in09 = reg_1343;
    91: op1_04_in09 = reg_1448;
    42: op1_04_in09 = reg_0132;
    67: op1_04_in09 = reg_1065;
    92: op1_04_in09 = reg_0607;
    93: op1_04_in09 = imem02_in[3:0];
    94: op1_04_in09 = reg_0886;
    96: op1_04_in09 = reg_0881;
    97: op1_04_in09 = reg_0460;
    98: op1_04_in09 = reg_0318;
    99: op1_04_in09 = reg_0406;
    100: op1_04_in09 = reg_0002;
    101: op1_04_in09 = reg_0361;
    102: op1_04_in09 = reg_0561;
    103: op1_04_in09 = reg_0048;
    104: op1_04_in09 = reg_0196;
    105: op1_04_in09 = reg_0722;
    106: op1_04_in09 = reg_0523;
    107: op1_04_in09 = reg_0426;
    131: op1_04_in09 = reg_0426;
    108: op1_04_in09 = reg_0000;
    109: op1_04_in09 = reg_0054;
    110: op1_04_in09 = reg_0140;
    111: op1_04_in09 = reg_0032;
    112: op1_04_in09 = reg_0001;
    113: op1_04_in09 = reg_0025;
    114: op1_04_in09 = reg_0595;
    115: op1_04_in09 = reg_0207;
    116: op1_04_in09 = reg_0786;
    117: op1_04_in09 = reg_1403;
    118: op1_04_in09 = reg_0782;
    119: op1_04_in09 = reg_0295;
    120: op1_04_in09 = reg_0250;
    121: op1_04_in09 = reg_0877;
    123: op1_04_in09 = reg_0879;
    124: op1_04_in09 = reg_0927;
    125: op1_04_in09 = reg_0827;
    127: op1_04_in09 = reg_0053;
    128: op1_04_in09 = reg_0309;
    130: op1_04_in09 = reg_0131;
    default: op1_04_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_04_inv09 = 1;
    71: op1_04_inv09 = 1;
    68: op1_04_inv09 = 1;
    74: op1_04_inv09 = 1;
    60: op1_04_inv09 = 1;
    48: op1_04_inv09 = 1;
    33: op1_04_inv09 = 1;
    57: op1_04_inv09 = 1;
    77: op1_04_inv09 = 1;
    70: op1_04_inv09 = 1;
    52: op1_04_inv09 = 1;
    58: op1_04_inv09 = 1;
    88: op1_04_inv09 = 1;
    59: op1_04_inv09 = 1;
    62: op1_04_inv09 = 1;
    44: op1_04_inv09 = 1;
    81: op1_04_inv09 = 1;
    82: op1_04_inv09 = 1;
    89: op1_04_inv09 = 1;
    47: op1_04_inv09 = 1;
    84: op1_04_inv09 = 1;
    65: op1_04_inv09 = 1;
    85: op1_04_inv09 = 1;
    90: op1_04_inv09 = 1;
    66: op1_04_inv09 = 1;
    91: op1_04_inv09 = 1;
    67: op1_04_inv09 = 1;
    92: op1_04_inv09 = 1;
    93: op1_04_inv09 = 1;
    94: op1_04_inv09 = 1;
    96: op1_04_inv09 = 1;
    102: op1_04_inv09 = 1;
    104: op1_04_inv09 = 1;
    105: op1_04_inv09 = 1;
    106: op1_04_inv09 = 1;
    109: op1_04_inv09 = 1;
    110: op1_04_inv09 = 1;
    117: op1_04_inv09 = 1;
    118: op1_04_inv09 = 1;
    119: op1_04_inv09 = 1;
    121: op1_04_inv09 = 1;
    122: op1_04_inv09 = 1;
    124: op1_04_inv09 = 1;
    125: op1_04_inv09 = 1;
    128: op1_04_inv09 = 1;
    default: op1_04_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in10 = reg_0221;
    55: op1_04_in10 = reg_0100;
    53: op1_04_in10 = reg_0531;
    73: op1_04_in10 = reg_0318;
    86: op1_04_in10 = reg_0452;
    49: op1_04_in10 = reg_0738;
    61: op1_04_in10 = reg_0642;
    69: op1_04_in10 = reg_0494;
    54: op1_04_in10 = reg_0050;
    50: op1_04_in10 = reg_0899;
    71: op1_04_in10 = reg_0785;
    68: op1_04_in10 = reg_1339;
    74: op1_04_in10 = reg_0961;
    75: op1_04_in10 = reg_1393;
    124: op1_04_in10 = reg_1393;
    87: op1_04_in10 = reg_1313;
    56: op1_04_in10 = reg_0031;
    46: op1_04_in10 = reg_0560;
    60: op1_04_in10 = reg_0412;
    76: op1_04_in10 = reg_0249;
    48: op1_04_in10 = reg_0094;
    57: op1_04_in10 = reg_0191;
    77: op1_04_in10 = reg_0016;
    70: op1_04_in10 = reg_0495;
    52: op1_04_in10 = reg_0928;
    58: op1_04_in10 = reg_0150;
    78: op1_04_in10 = reg_1132;
    88: op1_04_in10 = reg_0627;
    51: op1_04_in10 = reg_0135;
    63: op1_04_in10 = reg_0135;
    47: op1_04_in10 = reg_0135;
    79: op1_04_in10 = reg_0264;
    59: op1_04_in10 = reg_0456;
    80: op1_04_in10 = reg_0416;
    62: op1_04_in10 = reg_0784;
    44: op1_04_in10 = reg_0061;
    81: op1_04_in10 = reg_1214;
    82: op1_04_in10 = reg_1405;
    89: op1_04_in10 = reg_0294;
    83: op1_04_in10 = reg_0152;
    64: op1_04_in10 = reg_0873;
    84: op1_04_in10 = reg_1323;
    65: op1_04_in10 = reg_0379;
    85: op1_04_in10 = reg_0981;
    90: op1_04_in10 = reg_0435;
    66: op1_04_in10 = reg_0351;
    91: op1_04_in10 = reg_0177;
    42: op1_04_in10 = reg_0171;
    67: op1_04_in10 = reg_0396;
    92: op1_04_in10 = reg_0588;
    93: op1_04_in10 = reg_0608;
    94: op1_04_in10 = reg_0202;
    96: op1_04_in10 = reg_0202;
    95: op1_04_in10 = reg_1486;
    97: op1_04_in10 = reg_0459;
    126: op1_04_in10 = reg_0459;
    98: op1_04_in10 = reg_0197;
    99: op1_04_in10 = reg_0454;
    100: op1_04_in10 = reg_1182;
    101: op1_04_in10 = reg_0003;
    102: op1_04_in10 = imem02_in[3:0];
    103: op1_04_in10 = reg_1093;
    104: op1_04_in10 = reg_0240;
    105: op1_04_in10 = reg_0410;
    106: op1_04_in10 = reg_1229;
    107: op1_04_in10 = reg_0898;
    108: op1_04_in10 = reg_0314;
    109: op1_04_in10 = reg_1451;
    110: op1_04_in10 = reg_0457;
    111: op1_04_in10 = reg_0181;
    112: op1_04_in10 = reg_0086;
    113: op1_04_in10 = reg_0313;
    114: op1_04_in10 = reg_0292;
    115: op1_04_in10 = reg_0670;
    116: op1_04_in10 = reg_0703;
    117: op1_04_in10 = reg_0940;
    118: op1_04_in10 = reg_0860;
    119: op1_04_in10 = reg_0244;
    120: op1_04_in10 = reg_1027;
    121: op1_04_in10 = reg_0846;
    122: op1_04_in10 = reg_0957;
    123: op1_04_in10 = reg_1018;
    125: op1_04_in10 = reg_1504;
    127: op1_04_in10 = reg_0226;
    128: op1_04_in10 = reg_0158;
    129: op1_04_in10 = reg_0368;
    130: op1_04_in10 = reg_1404;
    131: op1_04_in10 = reg_0185;
    default: op1_04_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    49: op1_04_inv10 = 1;
    74: op1_04_inv10 = 1;
    75: op1_04_inv10 = 1;
    87: op1_04_inv10 = 1;
    60: op1_04_inv10 = 1;
    76: op1_04_inv10 = 1;
    48: op1_04_inv10 = 1;
    57: op1_04_inv10 = 1;
    77: op1_04_inv10 = 1;
    52: op1_04_inv10 = 1;
    51: op1_04_inv10 = 1;
    79: op1_04_inv10 = 1;
    62: op1_04_inv10 = 1;
    81: op1_04_inv10 = 1;
    83: op1_04_inv10 = 1;
    47: op1_04_inv10 = 1;
    64: op1_04_inv10 = 1;
    84: op1_04_inv10 = 1;
    66: op1_04_inv10 = 1;
    91: op1_04_inv10 = 1;
    42: op1_04_inv10 = 1;
    92: op1_04_inv10 = 1;
    93: op1_04_inv10 = 1;
    94: op1_04_inv10 = 1;
    95: op1_04_inv10 = 1;
    97: op1_04_inv10 = 1;
    98: op1_04_inv10 = 1;
    99: op1_04_inv10 = 1;
    100: op1_04_inv10 = 1;
    101: op1_04_inv10 = 1;
    103: op1_04_inv10 = 1;
    105: op1_04_inv10 = 1;
    107: op1_04_inv10 = 1;
    108: op1_04_inv10 = 1;
    109: op1_04_inv10 = 1;
    110: op1_04_inv10 = 1;
    111: op1_04_inv10 = 1;
    112: op1_04_inv10 = 1;
    113: op1_04_inv10 = 1;
    114: op1_04_inv10 = 1;
    115: op1_04_inv10 = 1;
    121: op1_04_inv10 = 1;
    122: op1_04_inv10 = 1;
    124: op1_04_inv10 = 1;
    125: op1_04_inv10 = 1;
    127: op1_04_inv10 = 1;
    129: op1_04_inv10 = 1;
    130: op1_04_inv10 = 1;
    131: op1_04_inv10 = 1;
    default: op1_04_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in11 = reg_1417;
    55: op1_04_in11 = reg_0228;
    53: op1_04_in11 = imem02_in[3:0];
    70: op1_04_in11 = imem02_in[3:0];
    73: op1_04_in11 = imem05_in[3:0];
    86: op1_04_in11 = reg_1419;
    49: op1_04_in11 = reg_0102;
    61: op1_04_in11 = reg_0201;
    94: op1_04_in11 = reg_0201;
    124: op1_04_in11 = reg_0201;
    69: op1_04_in11 = reg_0432;
    54: op1_04_in11 = reg_0003;
    50: op1_04_in11 = reg_0871;
    71: op1_04_in11 = reg_0611;
    68: op1_04_in11 = reg_1338;
    74: op1_04_in11 = reg_0821;
    75: op1_04_in11 = reg_0134;
    87: op1_04_in11 = reg_0220;
    56: op1_04_in11 = reg_0665;
    46: op1_04_in11 = reg_0533;
    60: op1_04_in11 = reg_0598;
    67: op1_04_in11 = reg_0598;
    76: op1_04_in11 = reg_0987;
    106: op1_04_in11 = reg_0987;
    48: op1_04_in11 = reg_0095;
    57: op1_04_in11 = reg_0490;
    77: op1_04_in11 = reg_0470;
    52: op1_04_in11 = reg_0638;
    58: op1_04_in11 = reg_0016;
    78: op1_04_in11 = reg_0312;
    88: op1_04_in11 = reg_0952;
    51: op1_04_in11 = reg_0162;
    79: op1_04_in11 = reg_0669;
    59: op1_04_in11 = reg_1018;
    80: op1_04_in11 = reg_0410;
    62: op1_04_in11 = imem06_in[15:12];
    115: op1_04_in11 = imem06_in[15:12];
    44: op1_04_in11 = reg_0033;
    81: op1_04_in11 = reg_1198;
    63: op1_04_in11 = reg_0926;
    82: op1_04_in11 = reg_0202;
    89: op1_04_in11 = reg_0848;
    83: op1_04_in11 = imem07_in[11:8];
    47: op1_04_in11 = imem07_in[15:12];
    64: op1_04_in11 = reg_0118;
    98: op1_04_in11 = reg_0118;
    84: op1_04_in11 = reg_0827;
    65: op1_04_in11 = reg_0712;
    85: op1_04_in11 = reg_0532;
    90: op1_04_in11 = reg_0405;
    96: op1_04_in11 = reg_0405;
    66: op1_04_in11 = reg_0189;
    91: op1_04_in11 = reg_0191;
    42: op1_04_in11 = reg_0419;
    92: op1_04_in11 = reg_1207;
    93: op1_04_in11 = reg_1344;
    95: op1_04_in11 = reg_0196;
    97: op1_04_in11 = reg_0440;
    99: op1_04_in11 = reg_0342;
    101: op1_04_in11 = reg_0052;
    102: op1_04_in11 = imem02_in[11:8];
    103: op1_04_in11 = reg_1226;
    104: op1_04_in11 = reg_0344;
    105: op1_04_in11 = reg_0071;
    107: op1_04_in11 = reg_1372;
    108: op1_04_in11 = reg_1313;
    109: op1_04_in11 = reg_0105;
    110: op1_04_in11 = reg_0156;
    111: op1_04_in11 = reg_1367;
    112: op1_04_in11 = reg_0123;
    113: op1_04_in11 = reg_0288;
    114: op1_04_in11 = reg_0080;
    116: op1_04_in11 = reg_0851;
    117: op1_04_in11 = reg_0792;
    118: op1_04_in11 = reg_0752;
    119: op1_04_in11 = reg_0583;
    120: op1_04_in11 = reg_0221;
    121: op1_04_in11 = reg_0138;
    122: op1_04_in11 = reg_1231;
    123: op1_04_in11 = reg_0056;
    125: op1_04_in11 = reg_0109;
    126: op1_04_in11 = reg_0524;
    128: op1_04_in11 = reg_0921;
    129: op1_04_in11 = reg_0252;
    130: op1_04_in11 = reg_1070;
    131: op1_04_in11 = reg_0177;
    default: op1_04_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_04_inv11 = 1;
    86: op1_04_inv11 = 1;
    61: op1_04_inv11 = 1;
    69: op1_04_inv11 = 1;
    54: op1_04_inv11 = 1;
    74: op1_04_inv11 = 1;
    87: op1_04_inv11 = 1;
    56: op1_04_inv11 = 1;
    46: op1_04_inv11 = 1;
    76: op1_04_inv11 = 1;
    57: op1_04_inv11 = 1;
    52: op1_04_inv11 = 1;
    58: op1_04_inv11 = 1;
    88: op1_04_inv11 = 1;
    51: op1_04_inv11 = 1;
    59: op1_04_inv11 = 1;
    62: op1_04_inv11 = 1;
    82: op1_04_inv11 = 1;
    84: op1_04_inv11 = 1;
    65: op1_04_inv11 = 1;
    90: op1_04_inv11 = 1;
    91: op1_04_inv11 = 1;
    96: op1_04_inv11 = 1;
    97: op1_04_inv11 = 1;
    98: op1_04_inv11 = 1;
    101: op1_04_inv11 = 1;
    102: op1_04_inv11 = 1;
    105: op1_04_inv11 = 1;
    106: op1_04_inv11 = 1;
    108: op1_04_inv11 = 1;
    109: op1_04_inv11 = 1;
    111: op1_04_inv11 = 1;
    112: op1_04_inv11 = 1;
    113: op1_04_inv11 = 1;
    115: op1_04_inv11 = 1;
    121: op1_04_inv11 = 1;
    122: op1_04_inv11 = 1;
    130: op1_04_inv11 = 1;
    default: op1_04_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in12 = reg_1406;
    126: op1_04_in12 = reg_1406;
    55: op1_04_in12 = reg_0051;
    53: op1_04_in12 = reg_0429;
    73: op1_04_in12 = imem05_in[11:8];
    86: op1_04_in12 = reg_0262;
    49: op1_04_in12 = reg_0100;
    61: op1_04_in12 = reg_0189;
    94: op1_04_in12 = reg_0189;
    69: op1_04_in12 = reg_0973;
    54: op1_04_in12 = reg_0085;
    101: op1_04_in12 = reg_0085;
    50: op1_04_in12 = reg_0080;
    71: op1_04_in12 = reg_0930;
    68: op1_04_in12 = reg_1065;
    74: op1_04_in12 = reg_1405;
    75: op1_04_in12 = reg_0071;
    96: op1_04_in12 = reg_0071;
    87: op1_04_in12 = reg_1301;
    56: op1_04_in12 = reg_0287;
    46: op1_04_in12 = reg_0473;
    60: op1_04_in12 = reg_0969;
    76: op1_04_in12 = reg_0229;
    48: op1_04_in12 = reg_0237;
    57: op1_04_in12 = reg_0225;
    77: op1_04_in12 = reg_0370;
    70: op1_04_in12 = reg_0106;
    52: op1_04_in12 = reg_0722;
    58: op1_04_in12 = reg_0033;
    78: op1_04_in12 = reg_0313;
    88: op1_04_in12 = reg_0220;
    51: op1_04_in12 = imem07_in[3:0];
    79: op1_04_in12 = reg_0115;
    59: op1_04_in12 = reg_0256;
    80: op1_04_in12 = reg_0060;
    62: op1_04_in12 = reg_0109;
    44: op1_04_in12 = reg_0034;
    81: op1_04_in12 = reg_0598;
    63: op1_04_in12 = reg_0641;
    82: op1_04_in12 = reg_0352;
    89: op1_04_in12 = reg_1078;
    83: op1_04_in12 = reg_0673;
    47: op1_04_in12 = reg_0703;
    64: op1_04_in12 = reg_0575;
    84: op1_04_in12 = reg_0110;
    65: op1_04_in12 = reg_0153;
    85: op1_04_in12 = reg_0390;
    90: op1_04_in12 = reg_0134;
    66: op1_04_in12 = reg_0428;
    124: op1_04_in12 = reg_0428;
    91: op1_04_in12 = reg_0144;
    42: op1_04_in12 = reg_0308;
    67: op1_04_in12 = reg_0452;
    92: op1_04_in12 = reg_0054;
    93: op1_04_in12 = reg_0254;
    95: op1_04_in12 = reg_0243;
    97: op1_04_in12 = reg_0435;
    98: op1_04_in12 = reg_0014;
    99: op1_04_in12 = reg_0232;
    102: op1_04_in12 = reg_0712;
    103: op1_04_in12 = reg_0108;
    104: op1_04_in12 = imem06_in[3:0];
    105: op1_04_in12 = reg_0058;
    106: op1_04_in12 = reg_1201;
    107: op1_04_in12 = reg_0181;
    108: op1_04_in12 = reg_0048;
    109: op1_04_in12 = reg_0629;
    110: op1_04_in12 = reg_0158;
    111: op1_04_in12 = reg_0493;
    113: op1_04_in12 = reg_1280;
    114: op1_04_in12 = reg_0078;
    115: op1_04_in12 = reg_0316;
    116: op1_04_in12 = reg_1350;
    117: op1_04_in12 = reg_1163;
    118: op1_04_in12 = reg_1505;
    119: op1_04_in12 = reg_0152;
    120: op1_04_in12 = reg_1459;
    121: op1_04_in12 = reg_0934;
    123: op1_04_in12 = reg_0934;
    122: op1_04_in12 = reg_1092;
    125: op1_04_in12 = reg_1302;
    128: op1_04_in12 = reg_0923;
    129: op1_04_in12 = reg_0721;
    130: op1_04_in12 = reg_1169;
    131: op1_04_in12 = reg_0847;
    default: op1_04_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_04_inv12 = 1;
    73: op1_04_inv12 = 1;
    49: op1_04_inv12 = 1;
    61: op1_04_inv12 = 1;
    54: op1_04_inv12 = 1;
    87: op1_04_inv12 = 1;
    56: op1_04_inv12 = 1;
    60: op1_04_inv12 = 1;
    48: op1_04_inv12 = 1;
    77: op1_04_inv12 = 1;
    52: op1_04_inv12 = 1;
    58: op1_04_inv12 = 1;
    78: op1_04_inv12 = 1;
    88: op1_04_inv12 = 1;
    80: op1_04_inv12 = 1;
    62: op1_04_inv12 = 1;
    81: op1_04_inv12 = 1;
    89: op1_04_inv12 = 1;
    64: op1_04_inv12 = 1;
    65: op1_04_inv12 = 1;
    85: op1_04_inv12 = 1;
    90: op1_04_inv12 = 1;
    42: op1_04_inv12 = 1;
    67: op1_04_inv12 = 1;
    92: op1_04_inv12 = 1;
    93: op1_04_inv12 = 1;
    96: op1_04_inv12 = 1;
    98: op1_04_inv12 = 1;
    101: op1_04_inv12 = 1;
    102: op1_04_inv12 = 1;
    103: op1_04_inv12 = 1;
    105: op1_04_inv12 = 1;
    106: op1_04_inv12 = 1;
    107: op1_04_inv12 = 1;
    109: op1_04_inv12 = 1;
    110: op1_04_inv12 = 1;
    114: op1_04_inv12 = 1;
    115: op1_04_inv12 = 1;
    119: op1_04_inv12 = 1;
    121: op1_04_inv12 = 1;
    122: op1_04_inv12 = 1;
    123: op1_04_inv12 = 1;
    130: op1_04_inv12 = 1;
    131: op1_04_inv12 = 1;
    default: op1_04_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in13 = reg_0821;
    55: op1_04_in13 = reg_0052;
    53: op1_04_in13 = reg_0326;
    73: op1_04_in13 = reg_0275;
    86: op1_04_in13 = reg_0835;
    49: op1_04_in13 = reg_0003;
    61: op1_04_in13 = reg_0134;
    69: op1_04_in13 = reg_0626;
    77: op1_04_in13 = reg_0626;
    54: op1_04_in13 = reg_0087;
    101: op1_04_in13 = reg_0087;
    50: op1_04_in13 = reg_0290;
    71: op1_04_in13 = reg_0259;
    68: op1_04_in13 = reg_1147;
    74: op1_04_in13 = reg_0928;
    75: op1_04_in13 = reg_1321;
    87: op1_04_in13 = reg_1208;
    56: op1_04_in13 = reg_0442;
    46: op1_04_in13 = reg_0456;
    60: op1_04_in13 = reg_0599;
    76: op1_04_in13 = reg_0155;
    48: op1_04_in13 = reg_0032;
    57: op1_04_in13 = reg_0310;
    70: op1_04_in13 = reg_0105;
    52: op1_04_in13 = reg_0189;
    58: op1_04_in13 = reg_0035;
    78: op1_04_in13 = reg_0191;
    88: op1_04_in13 = reg_0246;
    51: op1_04_in13 = imem07_in[7:4];
    79: op1_04_in13 = reg_0109;
    59: op1_04_in13 = reg_0889;
    80: op1_04_in13 = reg_1324;
    62: op1_04_in13 = reg_0619;
    125: op1_04_in13 = reg_0619;
    44: op1_04_in13 = reg_0792;
    81: op1_04_in13 = reg_0969;
    63: op1_04_in13 = reg_0642;
    82: op1_04_in13 = reg_0440;
    89: op1_04_in13 = reg_0279;
    83: op1_04_in13 = reg_0489;
    110: op1_04_in13 = reg_0489;
    47: op1_04_in13 = reg_0892;
    64: op1_04_in13 = reg_1346;
    84: op1_04_in13 = reg_0717;
    65: op1_04_in13 = reg_0848;
    85: op1_04_in13 = reg_0666;
    90: op1_04_in13 = reg_0073;
    66: op1_04_in13 = reg_0410;
    91: op1_04_in13 = reg_1517;
    42: op1_04_in13 = reg_0289;
    67: op1_04_in13 = reg_0721;
    92: op1_04_in13 = reg_1451;
    93: op1_04_in13 = reg_0839;
    94: op1_04_in13 = reg_0075;
    95: op1_04_in13 = reg_0602;
    96: op1_04_in13 = reg_0072;
    97: op1_04_in13 = reg_0416;
    98: op1_04_in13 = reg_0784;
    104: op1_04_in13 = reg_0784;
    99: op1_04_in13 = reg_1143;
    102: op1_04_in13 = reg_0744;
    103: op1_04_in13 = reg_0107;
    105: op1_04_in13 = reg_0267;
    106: op1_04_in13 = reg_0961;
    107: op1_04_in13 = reg_1367;
    108: op1_04_in13 = reg_0104;
    109: op1_04_in13 = reg_0307;
    111: op1_04_in13 = reg_1258;
    113: op1_04_in13 = reg_0425;
    114: op1_04_in13 = reg_0042;
    115: op1_04_in13 = reg_1323;
    116: op1_04_in13 = reg_1349;
    117: op1_04_in13 = reg_0418;
    118: op1_04_in13 = reg_1504;
    119: op1_04_in13 = reg_0215;
    120: op1_04_in13 = reg_0249;
    121: op1_04_in13 = reg_0900;
    122: op1_04_in13 = reg_0880;
    123: op1_04_in13 = reg_0533;
    124: op1_04_in13 = reg_0388;
    126: op1_04_in13 = reg_0201;
    128: op1_04_in13 = reg_0031;
    129: op1_04_in13 = reg_0731;
    130: op1_04_in13 = reg_1514;
    131: op1_04_in13 = reg_1001;
    default: op1_04_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv13 = 1;
    53: op1_04_inv13 = 1;
    73: op1_04_inv13 = 1;
    86: op1_04_inv13 = 1;
    49: op1_04_inv13 = 1;
    61: op1_04_inv13 = 1;
    71: op1_04_inv13 = 1;
    75: op1_04_inv13 = 1;
    87: op1_04_inv13 = 1;
    46: op1_04_inv13 = 1;
    76: op1_04_inv13 = 1;
    48: op1_04_inv13 = 1;
    57: op1_04_inv13 = 1;
    77: op1_04_inv13 = 1;
    59: op1_04_inv13 = 1;
    80: op1_04_inv13 = 1;
    62: op1_04_inv13 = 1;
    63: op1_04_inv13 = 1;
    83: op1_04_inv13 = 1;
    47: op1_04_inv13 = 1;
    64: op1_04_inv13 = 1;
    65: op1_04_inv13 = 1;
    90: op1_04_inv13 = 1;
    66: op1_04_inv13 = 1;
    42: op1_04_inv13 = 1;
    67: op1_04_inv13 = 1;
    92: op1_04_inv13 = 1;
    93: op1_04_inv13 = 1;
    95: op1_04_inv13 = 1;
    97: op1_04_inv13 = 1;
    101: op1_04_inv13 = 1;
    104: op1_04_inv13 = 1;
    106: op1_04_inv13 = 1;
    108: op1_04_inv13 = 1;
    109: op1_04_inv13 = 1;
    110: op1_04_inv13 = 1;
    114: op1_04_inv13 = 1;
    118: op1_04_inv13 = 1;
    119: op1_04_inv13 = 1;
    126: op1_04_inv13 = 1;
    129: op1_04_inv13 = 1;
    default: op1_04_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in14 = reg_1393;
    53: op1_04_in14 = reg_0971;
    73: op1_04_in14 = reg_0118;
    86: op1_04_in14 = reg_0117;
    49: op1_04_in14 = reg_0084;
    61: op1_04_in14 = reg_0388;
    69: op1_04_in14 = reg_0125;
    54: op1_04_in14 = reg_0123;
    50: op1_04_in14 = reg_0278;
    71: op1_04_in14 = reg_0547;
    68: op1_04_in14 = reg_0795;
    60: op1_04_in14 = reg_0795;
    74: op1_04_in14 = reg_0722;
    63: op1_04_in14 = reg_0722;
    75: op1_04_in14 = reg_0122;
    97: op1_04_in14 = reg_0122;
    87: op1_04_in14 = reg_0481;
    56: op1_04_in14 = reg_0103;
    46: op1_04_in14 = reg_0455;
    76: op1_04_in14 = reg_0409;
    48: op1_04_in14 = reg_0035;
    57: op1_04_in14 = reg_0298;
    77: op1_04_in14 = reg_0587;
    70: op1_04_in14 = reg_0382;
    52: op1_04_in14 = reg_0428;
    58: op1_04_in14 = reg_0735;
    78: op1_04_in14 = reg_0328;
    88: op1_04_in14 = reg_0048;
    51: op1_04_in14 = reg_1056;
    79: op1_04_in14 = reg_0716;
    59: op1_04_in14 = reg_0433;
    80: op1_04_in14 = reg_0005;
    62: op1_04_in14 = reg_0617;
    44: op1_04_in14 = reg_0794;
    81: op1_04_in14 = reg_0599;
    82: op1_04_in14 = reg_1321;
    89: op1_04_in14 = reg_0227;
    83: op1_04_in14 = reg_0663;
    47: op1_04_in14 = reg_0867;
    64: op1_04_in14 = reg_0828;
    84: op1_04_in14 = reg_0141;
    65: op1_04_in14 = reg_0839;
    85: op1_04_in14 = reg_0494;
    102: op1_04_in14 = reg_0494;
    90: op1_04_in14 = reg_1322;
    66: op1_04_in14 = reg_0405;
    91: op1_04_in14 = reg_1313;
    42: op1_04_in14 = reg_0458;
    108: op1_04_in14 = reg_0458;
    67: op1_04_in14 = reg_0596;
    92: op1_04_in14 = reg_1450;
    93: op1_04_in14 = reg_0778;
    94: op1_04_in14 = reg_0057;
    95: op1_04_in14 = reg_0206;
    96: op1_04_in14 = reg_0089;
    98: op1_04_in14 = reg_0908;
    99: op1_04_in14 = reg_0338;
    101: op1_04_in14 = reg_0520;
    103: op1_04_in14 = reg_0707;
    104: op1_04_in14 = reg_1058;
    105: op1_04_in14 = reg_0723;
    106: op1_04_in14 = reg_1432;
    107: op1_04_in14 = reg_0978;
    109: op1_04_in14 = reg_0829;
    110: op1_04_in14 = reg_0664;
    111: op1_04_in14 = reg_1215;
    113: op1_04_in14 = reg_0577;
    114: op1_04_in14 = imem01_in[7:4];
    115: op1_04_in14 = reg_0714;
    116: op1_04_in14 = reg_0924;
    117: op1_04_in14 = reg_0303;
    130: op1_04_in14 = reg_0303;
    118: op1_04_in14 = reg_0116;
    119: op1_04_in14 = reg_0214;
    120: op1_04_in14 = reg_0229;
    121: op1_04_in14 = reg_0054;
    122: op1_04_in14 = reg_0350;
    123: op1_04_in14 = reg_1207;
    124: op1_04_in14 = reg_0203;
    125: op1_04_in14 = reg_0527;
    126: op1_04_in14 = reg_0189;
    128: op1_04_in14 = reg_0286;
    129: op1_04_in14 = reg_0552;
    131: op1_04_in14 = reg_0311;
    default: op1_04_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_04_inv14 = 1;
    73: op1_04_inv14 = 1;
    86: op1_04_inv14 = 1;
    49: op1_04_inv14 = 1;
    61: op1_04_inv14 = 1;
    69: op1_04_inv14 = 1;
    54: op1_04_inv14 = 1;
    71: op1_04_inv14 = 1;
    68: op1_04_inv14 = 1;
    74: op1_04_inv14 = 1;
    75: op1_04_inv14 = 1;
    70: op1_04_inv14 = 1;
    52: op1_04_inv14 = 1;
    58: op1_04_inv14 = 1;
    78: op1_04_inv14 = 1;
    59: op1_04_inv14 = 1;
    62: op1_04_inv14 = 1;
    44: op1_04_inv14 = 1;
    81: op1_04_inv14 = 1;
    63: op1_04_inv14 = 1;
    89: op1_04_inv14 = 1;
    47: op1_04_inv14 = 1;
    67: op1_04_inv14 = 1;
    93: op1_04_inv14 = 1;
    96: op1_04_inv14 = 1;
    97: op1_04_inv14 = 1;
    105: op1_04_inv14 = 1;
    106: op1_04_inv14 = 1;
    107: op1_04_inv14 = 1;
    117: op1_04_inv14 = 1;
    120: op1_04_inv14 = 1;
    122: op1_04_inv14 = 1;
    123: op1_04_inv14 = 1;
    124: op1_04_inv14 = 1;
    126: op1_04_inv14 = 1;
    129: op1_04_inv14 = 1;
    131: op1_04_inv14 = 1;
    default: op1_04_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in15 = reg_0883;
    53: op1_04_in15 = reg_0126;
    73: op1_04_in15 = reg_0631;
    86: op1_04_in15 = reg_0210;
    61: op1_04_in15 = reg_0073;
    76: op1_04_in15 = reg_0073;
    69: op1_04_in15 = reg_0106;
    93: op1_04_in15 = reg_0106;
    54: op1_04_in15 = imem07_in[3:0];
    50: op1_04_in15 = reg_0043;
    71: op1_04_in15 = reg_0241;
    68: op1_04_in15 = reg_0936;
    74: op1_04_in15 = reg_0189;
    63: op1_04_in15 = reg_0189;
    75: op1_04_in15 = reg_0026;
    87: op1_04_in15 = reg_0443;
    56: op1_04_in15 = reg_0321;
    46: op1_04_in15 = reg_0433;
    60: op1_04_in15 = reg_0164;
    48: op1_04_in15 = reg_0799;
    57: op1_04_in15 = reg_0309;
    77: op1_04_in15 = reg_0204;
    70: op1_04_in15 = reg_0138;
    52: op1_04_in15 = reg_0431;
    58: op1_04_in15 = reg_0832;
    78: op1_04_in15 = reg_0216;
    88: op1_04_in15 = reg_0329;
    51: op1_04_in15 = reg_1060;
    79: op1_04_in15 = reg_0718;
    59: op1_04_in15 = reg_0971;
    80: op1_04_in15 = reg_0917;
    96: op1_04_in15 = reg_0917;
    62: op1_04_in15 = reg_0526;
    44: op1_04_in15 = reg_0578;
    81: op1_04_in15 = reg_0454;
    82: op1_04_in15 = reg_1322;
    89: op1_04_in15 = reg_0840;
    83: op1_04_in15 = reg_0437;
    110: op1_04_in15 = reg_0437;
    47: op1_04_in15 = reg_0187;
    64: op1_04_in15 = reg_1105;
    84: op1_04_in15 = reg_0622;
    65: op1_04_in15 = reg_0009;
    85: op1_04_in15 = reg_0432;
    90: op1_04_in15 = imem01_in[15:12];
    66: op1_04_in15 = reg_0134;
    91: op1_04_in15 = reg_0108;
    42: op1_04_in15 = reg_0023;
    67: op1_04_in15 = reg_0837;
    92: op1_04_in15 = reg_1455;
    94: op1_04_in15 = reg_0089;
    95: op1_04_in15 = reg_0037;
    97: op1_04_in15 = reg_1291;
    98: op1_04_in15 = reg_0397;
    99: op1_04_in15 = reg_0065;
    102: op1_04_in15 = reg_0054;
    103: op1_04_in15 = reg_0291;
    104: op1_04_in15 = reg_0270;
    105: op1_04_in15 = reg_0355;
    106: op1_04_in15 = reg_0927;
    107: op1_04_in15 = reg_0531;
    108: op1_04_in15 = reg_1282;
    109: op1_04_in15 = reg_0801;
    111: op1_04_in15 = reg_0281;
    113: op1_04_in15 = reg_0088;
    114: op1_04_in15 = reg_0561;
    115: op1_04_in15 = reg_1302;
    116: op1_04_in15 = reg_0779;
    117: op1_04_in15 = reg_0300;
    118: op1_04_in15 = reg_0717;
    119: op1_04_in15 = reg_0213;
    120: op1_04_in15 = reg_1417;
    121: op1_04_in15 = reg_0973;
    122: op1_04_in15 = reg_0707;
    123: op1_04_in15 = reg_0494;
    124: op1_04_in15 = reg_0060;
    125: op1_04_in15 = reg_0522;
    126: op1_04_in15 = reg_0416;
    128: op1_04_in15 = reg_0366;
    129: op1_04_in15 = reg_1200;
    130: op1_04_in15 = reg_0302;
    131: op1_04_in15 = reg_0180;
    default: op1_04_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv15 = 1;
    69: op1_04_inv15 = 1;
    50: op1_04_inv15 = 1;
    71: op1_04_inv15 = 1;
    68: op1_04_inv15 = 1;
    74: op1_04_inv15 = 1;
    46: op1_04_inv15 = 1;
    60: op1_04_inv15 = 1;
    48: op1_04_inv15 = 1;
    57: op1_04_inv15 = 1;
    70: op1_04_inv15 = 1;
    52: op1_04_inv15 = 1;
    58: op1_04_inv15 = 1;
    88: op1_04_inv15 = 1;
    51: op1_04_inv15 = 1;
    79: op1_04_inv15 = 1;
    44: op1_04_inv15 = 1;
    81: op1_04_inv15 = 1;
    82: op1_04_inv15 = 1;
    89: op1_04_inv15 = 1;
    84: op1_04_inv15 = 1;
    90: op1_04_inv15 = 1;
    66: op1_04_inv15 = 1;
    94: op1_04_inv15 = 1;
    95: op1_04_inv15 = 1;
    102: op1_04_inv15 = 1;
    103: op1_04_inv15 = 1;
    105: op1_04_inv15 = 1;
    106: op1_04_inv15 = 1;
    108: op1_04_inv15 = 1;
    109: op1_04_inv15 = 1;
    110: op1_04_inv15 = 1;
    111: op1_04_inv15 = 1;
    114: op1_04_inv15 = 1;
    117: op1_04_inv15 = 1;
    118: op1_04_inv15 = 1;
    119: op1_04_inv15 = 1;
    120: op1_04_inv15 = 1;
    121: op1_04_inv15 = 1;
    122: op1_04_inv15 = 1;
    125: op1_04_inv15 = 1;
    131: op1_04_inv15 = 1;
    default: op1_04_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in16 = reg_0410;
    53: op1_04_in16 = reg_0381;
    73: op1_04_in16 = reg_0864;
    86: op1_04_in16 = reg_0370;
    61: op1_04_in16 = imem01_in[7:4];
    69: op1_04_in16 = reg_0105;
    50: op1_04_in16 = reg_0041;
    71: op1_04_in16 = reg_0438;
    68: op1_04_in16 = reg_0451;
    74: op1_04_in16 = reg_0071;
    66: op1_04_in16 = reg_0071;
    75: op1_04_in16 = reg_0917;
    87: op1_04_in16 = reg_0263;
    56: op1_04_in16 = reg_0028;
    110: op1_04_in16 = reg_0028;
    46: op1_04_in16 = reg_0054;
    60: op1_04_in16 = reg_0181;
    76: op1_04_in16 = reg_0058;
    48: op1_04_in16 = reg_0749;
    57: op1_04_in16 = reg_0672;
    77: op1_04_in16 = reg_1430;
    70: op1_04_in16 = reg_0380;
    52: op1_04_in16 = reg_0416;
    58: op1_04_in16 = imem05_in[3:0];
    78: op1_04_in16 = reg_0557;
    88: op1_04_in16 = reg_0558;
    51: op1_04_in16 = reg_0324;
    79: op1_04_in16 = reg_0585;
    59: op1_04_in16 = reg_0933;
    80: op1_04_in16 = reg_1255;
    62: op1_04_in16 = reg_0527;
    44: op1_04_in16 = reg_0576;
    81: op1_04_in16 = reg_0304;
    63: op1_04_in16 = reg_0440;
    82: op1_04_in16 = reg_0267;
    89: op1_04_in16 = reg_0889;
    83: op1_04_in16 = reg_0739;
    47: op1_04_in16 = reg_0170;
    64: op1_04_in16 = imem06_in[3:0];
    84: op1_04_in16 = reg_0270;
    65: op1_04_in16 = imem02_in[15:12];
    85: op1_04_in16 = reg_1455;
    90: op1_04_in16 = reg_0653;
    91: op1_04_in16 = reg_0882;
    42: op1_04_in16 = reg_0046;
    67: op1_04_in16 = reg_0337;
    92: op1_04_in16 = reg_0106;
    93: op1_04_in16 = reg_1433;
    94: op1_04_in16 = reg_1032;
    95: op1_04_in16 = reg_1468;
    96: op1_04_in16 = reg_0166;
    97: op1_04_in16 = reg_0282;
    98: op1_04_in16 = reg_1326;
    99: op1_04_in16 = reg_1503;
    102: op1_04_in16 = reg_0126;
    103: op1_04_in16 = reg_0427;
    104: op1_04_in16 = reg_0161;
    105: op1_04_in16 = reg_0874;
    106: op1_04_in16 = reg_0881;
    107: op1_04_in16 = reg_0297;
    108: op1_04_in16 = reg_0348;
    109: op1_04_in16 = reg_0253;
    111: op1_04_in16 = reg_1419;
    113: op1_04_in16 = reg_0264;
    114: op1_04_in16 = reg_0455;
    115: op1_04_in16 = reg_1303;
    116: op1_04_in16 = reg_0029;
    117: op1_04_in16 = reg_0794;
    118: op1_04_in16 = reg_0637;
    119: op1_04_in16 = reg_1415;
    120: op1_04_in16 = reg_0524;
    121: op1_04_in16 = reg_0496;
    122: op1_04_in16 = reg_0378;
    123: op1_04_in16 = reg_0436;
    124: op1_04_in16 = reg_0788;
    125: op1_04_in16 = reg_0132;
    126: op1_04_in16 = reg_0060;
    128: op1_04_in16 = reg_0741;
    129: op1_04_in16 = reg_1004;
    130: op1_04_in16 = reg_0090;
    131: op1_04_in16 = reg_0891;
    default: op1_04_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv16 = 1;
    73: op1_04_inv16 = 1;
    86: op1_04_inv16 = 1;
    50: op1_04_inv16 = 1;
    71: op1_04_inv16 = 1;
    75: op1_04_inv16 = 1;
    87: op1_04_inv16 = 1;
    56: op1_04_inv16 = 1;
    60: op1_04_inv16 = 1;
    57: op1_04_inv16 = 1;
    52: op1_04_inv16 = 1;
    58: op1_04_inv16 = 1;
    78: op1_04_inv16 = 1;
    88: op1_04_inv16 = 1;
    51: op1_04_inv16 = 1;
    79: op1_04_inv16 = 1;
    44: op1_04_inv16 = 1;
    63: op1_04_inv16 = 1;
    82: op1_04_inv16 = 1;
    83: op1_04_inv16 = 1;
    64: op1_04_inv16 = 1;
    85: op1_04_inv16 = 1;
    66: op1_04_inv16 = 1;
    42: op1_04_inv16 = 1;
    67: op1_04_inv16 = 1;
    92: op1_04_inv16 = 1;
    95: op1_04_inv16 = 1;
    96: op1_04_inv16 = 1;
    97: op1_04_inv16 = 1;
    99: op1_04_inv16 = 1;
    102: op1_04_inv16 = 1;
    105: op1_04_inv16 = 1;
    107: op1_04_inv16 = 1;
    109: op1_04_inv16 = 1;
    111: op1_04_inv16 = 1;
    113: op1_04_inv16 = 1;
    118: op1_04_inv16 = 1;
    121: op1_04_inv16 = 1;
    122: op1_04_inv16 = 1;
    124: op1_04_inv16 = 1;
    125: op1_04_inv16 = 1;
    126: op1_04_inv16 = 1;
    130: op1_04_inv16 = 1;
    131: op1_04_inv16 = 1;
    default: op1_04_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in17 = reg_0134;
    53: op1_04_in17 = reg_0897;
    73: op1_04_in17 = reg_0207;
    86: op1_04_in17 = reg_0750;
    61: op1_04_in17 = reg_1253;
    69: op1_04_in17 = imem02_in[15:12];
    46: op1_04_in17 = imem02_in[15:12];
    50: op1_04_in17 = reg_0486;
    71: op1_04_in17 = reg_0726;
    68: op1_04_in17 = reg_0320;
    74: op1_04_in17 = reg_1321;
    75: op1_04_in17 = reg_1070;
    87: op1_04_in17 = reg_1369;
    56: op1_04_in17 = reg_0228;
    60: op1_04_in17 = reg_0129;
    76: op1_04_in17 = reg_0785;
    48: op1_04_in17 = imem05_in[3:0];
    57: op1_04_in17 = reg_0140;
    77: op1_04_in17 = reg_1431;
    70: op1_04_in17 = reg_0381;
    52: op1_04_in17 = reg_0075;
    58: op1_04_in17 = reg_1164;
    78: op1_04_in17 = reg_0710;
    88: op1_04_in17 = reg_1231;
    51: op1_04_in17 = reg_0894;
    79: op1_04_in17 = reg_0586;
    115: op1_04_in17 = reg_0586;
    59: op1_04_in17 = reg_0125;
    80: op1_04_in17 = reg_0277;
    62: op1_04_in17 = reg_1228;
    44: op1_04_in17 = reg_0346;
    81: op1_04_in17 = reg_0319;
    63: op1_04_in17 = reg_0388;
    82: op1_04_in17 = imem01_in[7:4];
    126: op1_04_in17 = imem01_in[7:4];
    89: op1_04_in17 = reg_0235;
    83: op1_04_in17 = reg_0738;
    47: op1_04_in17 = reg_0851;
    64: op1_04_in17 = reg_0859;
    84: op1_04_in17 = reg_0269;
    65: op1_04_in17 = reg_0276;
    85: op1_04_in17 = reg_0106;
    90: op1_04_in17 = reg_0754;
    66: op1_04_in17 = reg_0203;
    91: op1_04_in17 = reg_0707;
    42: op1_04_in17 = reg_0213;
    67: op1_04_in17 = reg_0094;
    92: op1_04_in17 = reg_1091;
    93: op1_04_in17 = reg_1140;
    94: op1_04_in17 = reg_1254;
    95: op1_04_in17 = reg_0397;
    96: op1_04_in17 = reg_1291;
    97: op1_04_in17 = reg_0355;
    98: op1_04_in17 = reg_0751;
    99: op1_04_in17 = reg_0210;
    102: op1_04_in17 = reg_0631;
    103: op1_04_in17 = imem04_in[7:4];
    104: op1_04_in17 = reg_0730;
    105: op1_04_in17 = reg_0902;
    106: op1_04_in17 = reg_0883;
    107: op1_04_in17 = reg_0574;
    108: op1_04_in17 = reg_1383;
    109: op1_04_in17 = reg_0007;
    110: op1_04_in17 = reg_0361;
    111: op1_04_in17 = reg_0369;
    113: op1_04_in17 = reg_0797;
    114: op1_04_in17 = reg_0133;
    116: op1_04_in17 = reg_0665;
    117: op1_04_in17 = reg_0602;
    118: op1_04_in17 = reg_0529;
    119: op1_04_in17 = reg_1057;
    120: op1_04_in17 = reg_1405;
    121: op1_04_in17 = reg_0380;
    122: op1_04_in17 = reg_0218;
    123: op1_04_in17 = reg_0778;
    124: op1_04_in17 = reg_0331;
    125: op1_04_in17 = reg_0296;
    128: op1_04_in17 = reg_0408;
    129: op1_04_in17 = reg_0061;
    130: op1_04_in17 = reg_0736;
    131: op1_04_in17 = reg_0070;
    default: op1_04_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv17 = 1;
    86: op1_04_inv17 = 1;
    61: op1_04_inv17 = 1;
    50: op1_04_inv17 = 1;
    68: op1_04_inv17 = 1;
    74: op1_04_inv17 = 1;
    87: op1_04_inv17 = 1;
    56: op1_04_inv17 = 1;
    46: op1_04_inv17 = 1;
    60: op1_04_inv17 = 1;
    76: op1_04_inv17 = 1;
    48: op1_04_inv17 = 1;
    57: op1_04_inv17 = 1;
    77: op1_04_inv17 = 1;
    58: op1_04_inv17 = 1;
    78: op1_04_inv17 = 1;
    79: op1_04_inv17 = 1;
    62: op1_04_inv17 = 1;
    44: op1_04_inv17 = 1;
    63: op1_04_inv17 = 1;
    82: op1_04_inv17 = 1;
    83: op1_04_inv17 = 1;
    47: op1_04_inv17 = 1;
    84: op1_04_inv17 = 1;
    90: op1_04_inv17 = 1;
    66: op1_04_inv17 = 1;
    91: op1_04_inv17 = 1;
    42: op1_04_inv17 = 1;
    93: op1_04_inv17 = 1;
    94: op1_04_inv17 = 1;
    95: op1_04_inv17 = 1;
    96: op1_04_inv17 = 1;
    97: op1_04_inv17 = 1;
    98: op1_04_inv17 = 1;
    104: op1_04_inv17 = 1;
    107: op1_04_inv17 = 1;
    110: op1_04_inv17 = 1;
    114: op1_04_inv17 = 1;
    118: op1_04_inv17 = 1;
    123: op1_04_inv17 = 1;
    125: op1_04_inv17 = 1;
    126: op1_04_inv17 = 1;
    128: op1_04_inv17 = 1;
    129: op1_04_inv17 = 1;
    130: op1_04_inv17 = 1;
    131: op1_04_inv17 = 1;
    default: op1_04_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in18 = reg_0073;
    53: op1_04_in18 = reg_0898;
    73: op1_04_in18 = reg_0037;
    86: op1_04_in18 = reg_1431;
    61: op1_04_in18 = reg_1256;
    69: op1_04_in18 = reg_0379;
    59: op1_04_in18 = reg_0379;
    50: op1_04_in18 = imem02_in[15:12];
    71: op1_04_in18 = reg_0092;
    68: op1_04_in18 = reg_0342;
    74: op1_04_in18 = reg_0122;
    75: op1_04_in18 = reg_1069;
    87: op1_04_in18 = reg_1368;
    56: op1_04_in18 = reg_0051;
    46: op1_04_in18 = reg_0934;
    60: op1_04_in18 = reg_0016;
    76: op1_04_in18 = reg_0448;
    48: op1_04_in18 = reg_0646;
    57: op1_04_in18 = reg_0285;
    77: op1_04_in18 = reg_0879;
    70: op1_04_in18 = reg_0708;
    52: op1_04_in18 = reg_0057;
    58: op1_04_in18 = reg_1169;
    78: op1_04_in18 = reg_0199;
    88: op1_04_in18 = reg_1199;
    51: op1_04_in18 = reg_0170;
    79: op1_04_in18 = reg_0571;
    80: op1_04_in18 = reg_0963;
    62: op1_04_in18 = reg_0171;
    44: op1_04_in18 = reg_0828;
    81: op1_04_in18 = reg_0487;
    63: op1_04_in18 = reg_0352;
    106: op1_04_in18 = reg_0352;
    120: op1_04_in18 = reg_0352;
    82: op1_04_in18 = imem01_in[11:8];
    89: op1_04_in18 = reg_0185;
    83: op1_04_in18 = reg_0408;
    47: op1_04_in18 = reg_0672;
    64: op1_04_in18 = reg_0752;
    84: op1_04_in18 = reg_0213;
    65: op1_04_in18 = reg_1132;
    85: op1_04_in18 = reg_0824;
    90: op1_04_in18 = reg_0610;
    66: op1_04_in18 = reg_1322;
    91: op1_04_in18 = reg_0378;
    42: op1_04_in18 = reg_0230;
    67: op1_04_in18 = reg_0164;
    92: op1_04_in18 = reg_0024;
    93: op1_04_in18 = reg_0473;
    94: op1_04_in18 = reg_0754;
    95: op1_04_in18 = reg_0960;
    96: op1_04_in18 = reg_1032;
    97: op1_04_in18 = reg_0258;
    98: op1_04_in18 = reg_0109;
    99: op1_04_in18 = reg_1164;
    102: op1_04_in18 = reg_0897;
    103: op1_04_in18 = reg_1383;
    104: op1_04_in18 = reg_0984;
    105: op1_04_in18 = reg_0093;
    107: op1_04_in18 = reg_0406;
    108: op1_04_in18 = reg_0731;
    109: op1_04_in18 = reg_1078;
    110: op1_04_in18 = reg_0228;
    111: op1_04_in18 = reg_0268;
    113: op1_04_in18 = reg_0462;
    114: op1_04_in18 = reg_0839;
    115: op1_04_in18 = reg_0617;
    116: op1_04_in18 = reg_0663;
    117: op1_04_in18 = reg_0589;
    118: op1_04_in18 = reg_0568;
    119: op1_04_in18 = reg_0993;
    121: op1_04_in18 = reg_0381;
    122: op1_04_in18 = reg_0313;
    123: op1_04_in18 = reg_0128;
    124: op1_04_in18 = reg_0968;
    125: op1_04_in18 = reg_0977;
    126: op1_04_in18 = reg_0548;
    128: op1_04_in18 = reg_0620;
    129: op1_04_in18 = reg_0369;
    130: op1_04_in18 = reg_0450;
    131: op1_04_in18 = reg_1518;
    default: op1_04_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv18 = 1;
    53: op1_04_inv18 = 1;
    61: op1_04_inv18 = 1;
    71: op1_04_inv18 = 1;
    74: op1_04_inv18 = 1;
    75: op1_04_inv18 = 1;
    87: op1_04_inv18 = 1;
    48: op1_04_inv18 = 1;
    70: op1_04_inv18 = 1;
    58: op1_04_inv18 = 1;
    78: op1_04_inv18 = 1;
    88: op1_04_inv18 = 1;
    51: op1_04_inv18 = 1;
    59: op1_04_inv18 = 1;
    62: op1_04_inv18 = 1;
    47: op1_04_inv18 = 1;
    64: op1_04_inv18 = 1;
    66: op1_04_inv18 = 1;
    91: op1_04_inv18 = 1;
    67: op1_04_inv18 = 1;
    92: op1_04_inv18 = 1;
    94: op1_04_inv18 = 1;
    96: op1_04_inv18 = 1;
    99: op1_04_inv18 = 1;
    102: op1_04_inv18 = 1;
    103: op1_04_inv18 = 1;
    105: op1_04_inv18 = 1;
    107: op1_04_inv18 = 1;
    109: op1_04_inv18 = 1;
    110: op1_04_inv18 = 1;
    111: op1_04_inv18 = 1;
    113: op1_04_inv18 = 1;
    115: op1_04_inv18 = 1;
    116: op1_04_inv18 = 1;
    117: op1_04_inv18 = 1;
    119: op1_04_inv18 = 1;
    122: op1_04_inv18 = 1;
    124: op1_04_inv18 = 1;
    125: op1_04_inv18 = 1;
    126: op1_04_inv18 = 1;
    128: op1_04_inv18 = 1;
    default: op1_04_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in19 = reg_0060;
    53: op1_04_in19 = reg_0708;
    73: op1_04_in19 = reg_0038;
    86: op1_04_in19 = reg_0272;
    61: op1_04_in19 = reg_1034;
    69: op1_04_in19 = reg_0848;
    50: op1_04_in19 = reg_1029;
    71: op1_04_in19 = reg_0874;
    68: op1_04_in19 = reg_0721;
    74: op1_04_in19 = reg_0026;
    75: op1_04_in19 = imem01_in[15:12];
    87: op1_04_in19 = reg_0493;
    56: op1_04_in19 = reg_0004;
    46: op1_04_in19 = reg_0105;
    60: op1_04_in19 = reg_0032;
    103: op1_04_in19 = reg_0032;
    76: op1_04_in19 = reg_1255;
    48: op1_04_in19 = reg_0997;
    57: op1_04_in19 = reg_0366;
    77: op1_04_in19 = reg_1168;
    70: op1_04_in19 = reg_0379;
    52: op1_04_in19 = reg_0267;
    58: op1_04_in19 = reg_0996;
    99: op1_04_in19 = reg_0996;
    78: op1_04_in19 = reg_1033;
    88: op1_04_in19 = reg_0448;
    51: op1_04_in19 = reg_0309;
    79: op1_04_in19 = reg_1225;
    59: op1_04_in19 = reg_0390;
    80: op1_04_in19 = reg_0798;
    62: op1_04_in19 = reg_0269;
    44: op1_04_in19 = reg_0701;
    81: op1_04_in19 = reg_0368;
    63: op1_04_in19 = reg_0122;
    82: op1_04_in19 = reg_1290;
    89: op1_04_in19 = reg_0823;
    83: op1_04_in19 = reg_0618;
    47: op1_04_in19 = reg_0159;
    64: op1_04_in19 = reg_0133;
    84: op1_04_in19 = reg_0034;
    65: op1_04_in19 = reg_0227;
    85: op1_04_in19 = imem02_in[11:8];
    90: op1_04_in19 = reg_0609;
    66: op1_04_in19 = reg_0089;
    91: op1_04_in19 = reg_0247;
    42: op1_04_in19 = reg_0231;
    67: op1_04_in19 = reg_0035;
    92: op1_04_in19 = imem03_in[11:8];
    93: op1_04_in19 = reg_0801;
    94: op1_04_in19 = reg_0549;
    95: op1_04_in19 = reg_0751;
    96: op1_04_in19 = reg_0930;
    97: op1_04_in19 = reg_0550;
    98: op1_04_in19 = reg_0714;
    102: op1_04_in19 = reg_1098;
    104: op1_04_in19 = reg_0585;
    105: op1_04_in19 = reg_0463;
    106: op1_04_in19 = reg_0201;
    107: op1_04_in19 = reg_0471;
    108: op1_04_in19 = reg_0694;
    109: op1_04_in19 = reg_0069;
    110: op1_04_in19 = reg_0051;
    111: op1_04_in19 = reg_0862;
    113: op1_04_in19 = reg_1083;
    114: op1_04_in19 = reg_0533;
    115: op1_04_in19 = reg_0345;
    116: op1_04_in19 = reg_0741;
    117: op1_04_in19 = reg_0449;
    118: op1_04_in19 = reg_0583;
    119: op1_04_in19 = reg_1056;
    120: op1_04_in19 = reg_0189;
    121: op1_04_in19 = reg_0307;
    122: op1_04_in19 = reg_0425;
    123: op1_04_in19 = reg_0382;
    124: op1_04_in19 = reg_0819;
    125: op1_04_in19 = reg_0214;
    126: op1_04_in19 = reg_0260;
    128: op1_04_in19 = reg_0593;
    129: op1_04_in19 = reg_0836;
    130: op1_04_in19 = reg_0066;
    131: op1_04_in19 = reg_1314;
    default: op1_04_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv19 = 1;
    73: op1_04_inv19 = 1;
    71: op1_04_inv19 = 1;
    74: op1_04_inv19 = 1;
    75: op1_04_inv19 = 1;
    46: op1_04_inv19 = 1;
    70: op1_04_inv19 = 1;
    78: op1_04_inv19 = 1;
    59: op1_04_inv19 = 1;
    62: op1_04_inv19 = 1;
    44: op1_04_inv19 = 1;
    89: op1_04_inv19 = 1;
    64: op1_04_inv19 = 1;
    65: op1_04_inv19 = 1;
    91: op1_04_inv19 = 1;
    67: op1_04_inv19 = 1;
    92: op1_04_inv19 = 1;
    93: op1_04_inv19 = 1;
    94: op1_04_inv19 = 1;
    95: op1_04_inv19 = 1;
    97: op1_04_inv19 = 1;
    98: op1_04_inv19 = 1;
    102: op1_04_inv19 = 1;
    105: op1_04_inv19 = 1;
    113: op1_04_inv19 = 1;
    114: op1_04_inv19 = 1;
    116: op1_04_inv19 = 1;
    118: op1_04_inv19 = 1;
    119: op1_04_inv19 = 1;
    123: op1_04_inv19 = 1;
    126: op1_04_inv19 = 1;
    128: op1_04_inv19 = 1;
    130: op1_04_inv19 = 1;
    default: op1_04_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in20 = reg_1321;
    53: op1_04_in20 = reg_0009;
    73: op1_04_in20 = reg_0040;
    86: op1_04_in20 = reg_0700;
    61: op1_04_in20 = reg_0984;
    69: op1_04_in20 = reg_0327;
    50: op1_04_in20 = reg_0456;
    71: op1_04_in20 = reg_0079;
    68: op1_04_in20 = reg_0837;
    81: op1_04_in20 = reg_0837;
    74: op1_04_in20 = reg_1100;
    75: op1_04_in20 = reg_0047;
    87: op1_04_in20 = reg_0264;
    56: op1_04_in20 = reg_0002;
    46: op1_04_in20 = reg_0381;
    123: op1_04_in20 = reg_0381;
    60: op1_04_in20 = reg_0631;
    76: op1_04_in20 = reg_1253;
    48: op1_04_in20 = reg_0332;
    57: op1_04_in20 = reg_0739;
    77: op1_04_in20 = reg_1169;
    70: op1_04_in20 = reg_0695;
    52: op1_04_in20 = reg_0723;
    58: op1_04_in20 = reg_1212;
    78: op1_04_in20 = reg_0376;
    88: op1_04_in20 = reg_0458;
    51: op1_04_in20 = reg_0672;
    79: op1_04_in20 = reg_0419;
    59: op1_04_in20 = reg_0900;
    80: op1_04_in20 = reg_1474;
    62: op1_04_in20 = reg_0215;
    44: op1_04_in20 = reg_0250;
    63: op1_04_in20 = reg_0089;
    82: op1_04_in20 = reg_0549;
    105: op1_04_in20 = reg_0549;
    89: op1_04_in20 = reg_1184;
    83: op1_04_in20 = reg_0593;
    47: op1_04_in20 = reg_0157;
    64: op1_04_in20 = reg_0316;
    84: op1_04_in20 = imem07_in[11:8];
    65: op1_04_in20 = reg_0707;
    85: op1_04_in20 = reg_0294;
    90: op1_04_in20 = reg_0239;
    66: op1_04_in20 = reg_0026;
    91: op1_04_in20 = reg_0263;
    103: op1_04_in20 = reg_0263;
    42: op1_04_in20 = reg_0246;
    67: op1_04_in20 = reg_0793;
    92: op1_04_in20 = reg_0504;
    93: op1_04_in20 = reg_0006;
    94: op1_04_in20 = reg_0609;
    97: op1_04_in20 = reg_0609;
    95: op1_04_in20 = reg_0860;
    96: op1_04_in20 = reg_0163;
    98: op1_04_in20 = reg_0194;
    99: op1_04_in20 = reg_0992;
    102: op1_04_in20 = reg_0235;
    104: op1_04_in20 = reg_0295;
    106: op1_04_in20 = reg_0416;
    107: op1_04_in20 = reg_0061;
    108: op1_04_in20 = reg_0297;
    109: op1_04_in20 = reg_0710;
    111: op1_04_in20 = reg_0835;
    113: op1_04_in20 = reg_1200;
    114: op1_04_in20 = reg_1207;
    115: op1_04_in20 = reg_0308;
    116: op1_04_in20 = reg_0408;
    117: op1_04_in20 = reg_0929;
    118: op1_04_in20 = reg_0195;
    119: op1_04_in20 = reg_0309;
    120: op1_04_in20 = reg_0405;
    121: op1_04_in20 = reg_0473;
    122: op1_04_in20 = imem04_in[11:8];
    124: op1_04_in20 = reg_0439;
    125: op1_04_in20 = reg_0169;
    126: op1_04_in20 = reg_0820;
    128: op1_04_in20 = reg_0321;
    129: op1_04_in20 = imem04_in[3:0];
    130: op1_04_in20 = reg_0347;
    131: op1_04_in20 = reg_1092;
    default: op1_04_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv20 = 1;
    53: op1_04_inv20 = 1;
    50: op1_04_inv20 = 1;
    71: op1_04_inv20 = 1;
    68: op1_04_inv20 = 1;
    46: op1_04_inv20 = 1;
    70: op1_04_inv20 = 1;
    78: op1_04_inv20 = 1;
    80: op1_04_inv20 = 1;
    62: op1_04_inv20 = 1;
    63: op1_04_inv20 = 1;
    82: op1_04_inv20 = 1;
    89: op1_04_inv20 = 1;
    85: op1_04_inv20 = 1;
    42: op1_04_inv20 = 1;
    67: op1_04_inv20 = 1;
    92: op1_04_inv20 = 1;
    93: op1_04_inv20 = 1;
    94: op1_04_inv20 = 1;
    95: op1_04_inv20 = 1;
    96: op1_04_inv20 = 1;
    102: op1_04_inv20 = 1;
    103: op1_04_inv20 = 1;
    105: op1_04_inv20 = 1;
    106: op1_04_inv20 = 1;
    107: op1_04_inv20 = 1;
    108: op1_04_inv20 = 1;
    113: op1_04_inv20 = 1;
    117: op1_04_inv20 = 1;
    118: op1_04_inv20 = 1;
    119: op1_04_inv20 = 1;
    120: op1_04_inv20 = 1;
    121: op1_04_inv20 = 1;
    122: op1_04_inv20 = 1;
    124: op1_04_inv20 = 1;
    125: op1_04_inv20 = 1;
    126: op1_04_inv20 = 1;
    128: op1_04_inv20 = 1;
    129: op1_04_inv20 = 1;
    130: op1_04_inv20 = 1;
    default: op1_04_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in21 = reg_0057;
    53: op1_04_in21 = reg_0024;
    73: op1_04_in21 = reg_0039;
    86: op1_04_in21 = reg_0648;
    61: op1_04_in21 = reg_1151;
    111: op1_04_in21 = reg_1151;
    69: op1_04_in21 = reg_0820;
    50: op1_04_in21 = reg_0588;
    71: op1_04_in21 = reg_0283;
    68: op1_04_in21 = reg_0117;
    74: op1_04_in21 = reg_0372;
    75: op1_04_in21 = reg_0258;
    87: op1_04_in21 = reg_1338;
    56: op1_04_in21 = reg_0053;
    46: op1_04_in21 = reg_0390;
    60: op1_04_in21 = reg_0346;
    76: op1_04_in21 = imem01_in[3:0];
    124: op1_04_in21 = imem01_in[3:0];
    48: op1_04_in21 = reg_0450;
    57: op1_04_in21 = reg_0741;
    77: op1_04_in21 = reg_0174;
    70: op1_04_in21 = reg_0756;
    52: op1_04_in21 = reg_1090;
    58: op1_04_in21 = reg_0565;
    78: op1_04_in21 = imem03_in[11:8];
    109: op1_04_in21 = imem03_in[11:8];
    88: op1_04_in21 = reg_1139;
    51: op1_04_in21 = reg_0924;
    79: op1_04_in21 = reg_0289;
    115: op1_04_in21 = reg_0289;
    59: op1_04_in21 = reg_0708;
    80: op1_04_in21 = reg_0469;
    97: op1_04_in21 = reg_0469;
    62: op1_04_in21 = reg_1170;
    44: op1_04_in21 = reg_0649;
    81: op1_04_in21 = reg_0719;
    63: op1_04_in21 = reg_0027;
    82: op1_04_in21 = reg_0222;
    89: op1_04_in21 = reg_0964;
    83: op1_04_in21 = reg_0050;
    47: op1_04_in21 = reg_0139;
    64: op1_04_in21 = reg_0194;
    84: op1_04_in21 = imem07_in[15:12];
    65: op1_04_in21 = reg_0375;
    85: op1_04_in21 = reg_0068;
    90: op1_04_in21 = reg_0468;
    66: op1_04_in21 = reg_0267;
    91: op1_04_in21 = reg_0088;
    103: op1_04_in21 = reg_0088;
    42: op1_04_in21 = reg_0324;
    67: op1_04_in21 = reg_0391;
    92: op1_04_in21 = reg_0889;
    93: op1_04_in21 = reg_0758;
    94: op1_04_in21 = reg_0239;
    95: op1_04_in21 = reg_1504;
    96: op1_04_in21 = reg_0547;
    98: op1_04_in21 = reg_0398;
    99: op1_04_in21 = reg_0604;
    102: op1_04_in21 = reg_0505;
    104: op1_04_in21 = reg_0308;
    105: op1_04_in21 = reg_0966;
    106: op1_04_in21 = reg_0409;
    107: op1_04_in21 = reg_0062;
    108: op1_04_in21 = reg_1082;
    113: op1_04_in21 = reg_0281;
    114: op1_04_in21 = reg_0436;
    116: op1_04_in21 = reg_0028;
    128: op1_04_in21 = reg_0028;
    117: op1_04_in21 = reg_0669;
    118: op1_04_in21 = reg_0067;
    119: op1_04_in21 = reg_0851;
    120: op1_04_in21 = reg_0387;
    121: op1_04_in21 = reg_0802;
    122: op1_04_in21 = reg_1339;
    123: op1_04_in21 = reg_0306;
    125: op1_04_in21 = reg_0087;
    126: op1_04_in21 = reg_0742;
    129: op1_04_in21 = reg_0095;
    130: op1_04_in21 = reg_0601;
    131: op1_04_in21 = reg_1208;
    default: op1_04_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_04_inv21 = 1;
    50: op1_04_inv21 = 1;
    71: op1_04_inv21 = 1;
    68: op1_04_inv21 = 1;
    74: op1_04_inv21 = 1;
    75: op1_04_inv21 = 1;
    87: op1_04_inv21 = 1;
    56: op1_04_inv21 = 1;
    46: op1_04_inv21 = 1;
    60: op1_04_inv21 = 1;
    76: op1_04_inv21 = 1;
    48: op1_04_inv21 = 1;
    78: op1_04_inv21 = 1;
    88: op1_04_inv21 = 1;
    51: op1_04_inv21 = 1;
    79: op1_04_inv21 = 1;
    59: op1_04_inv21 = 1;
    62: op1_04_inv21 = 1;
    44: op1_04_inv21 = 1;
    81: op1_04_inv21 = 1;
    63: op1_04_inv21 = 1;
    82: op1_04_inv21 = 1;
    47: op1_04_inv21 = 1;
    85: op1_04_inv21 = 1;
    90: op1_04_inv21 = 1;
    66: op1_04_inv21 = 1;
    91: op1_04_inv21 = 1;
    92: op1_04_inv21 = 1;
    94: op1_04_inv21 = 1;
    95: op1_04_inv21 = 1;
    96: op1_04_inv21 = 1;
    98: op1_04_inv21 = 1;
    99: op1_04_inv21 = 1;
    106: op1_04_inv21 = 1;
    107: op1_04_inv21 = 1;
    108: op1_04_inv21 = 1;
    109: op1_04_inv21 = 1;
    111: op1_04_inv21 = 1;
    113: op1_04_inv21 = 1;
    114: op1_04_inv21 = 1;
    115: op1_04_inv21 = 1;
    117: op1_04_inv21 = 1;
    120: op1_04_inv21 = 1;
    122: op1_04_inv21 = 1;
    123: op1_04_inv21 = 1;
    125: op1_04_inv21 = 1;
    126: op1_04_inv21 = 1;
    128: op1_04_inv21 = 1;
    130: op1_04_inv21 = 1;
    131: op1_04_inv21 = 1;
    default: op1_04_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in22 = reg_0122;
    53: op1_04_in22 = reg_0802;
    73: op1_04_in22 = reg_0195;
    86: op1_04_in22 = reg_0649;
    61: op1_04_in22 = reg_0982;
    69: op1_04_in22 = reg_0801;
    50: op1_04_in22 = reg_0562;
    99: op1_04_in22 = reg_0562;
    71: op1_04_in22 = reg_0043;
    68: op1_04_in22 = reg_0210;
    74: op1_04_in22 = reg_1290;
    66: op1_04_in22 = reg_1290;
    75: op1_04_in22 = reg_0549;
    96: op1_04_in22 = reg_0549;
    87: op1_04_in22 = reg_0531;
    56: op1_04_in22 = reg_1182;
    116: op1_04_in22 = reg_1182;
    46: op1_04_in22 = reg_0055;
    60: op1_04_in22 = reg_0174;
    76: op1_04_in22 = reg_0331;
    48: op1_04_in22 = reg_0168;
    57: op1_04_in22 = reg_0592;
    77: op1_04_in22 = imem05_in[15:12];
    70: op1_04_in22 = reg_0732;
    52: op1_04_in22 = reg_1070;
    58: op1_04_in22 = reg_0564;
    78: op1_04_in22 = imem03_in[15:12];
    88: op1_04_in22 = reg_1325;
    51: op1_04_in22 = reg_0139;
    79: op1_04_in22 = reg_0165;
    59: op1_04_in22 = reg_0705;
    80: op1_04_in22 = reg_0966;
    62: op1_04_in22 = reg_0230;
    44: op1_04_in22 = reg_0604;
    81: op1_04_in22 = reg_0096;
    63: op1_04_in22 = reg_0822;
    82: op1_04_in22 = reg_0238;
    89: op1_04_in22 = reg_0478;
    83: op1_04_in22 = reg_0519;
    47: op1_04_in22 = reg_0404;
    64: op1_04_in22 = reg_0585;
    84: op1_04_in22 = reg_0186;
    65: op1_04_in22 = reg_0640;
    85: op1_04_in22 = reg_0217;
    90: op1_04_in22 = reg_0430;
    91: op1_04_in22 = reg_0034;
    42: op1_04_in22 = reg_0191;
    67: op1_04_in22 = reg_0750;
    92: op1_04_in22 = reg_0559;
    93: op1_04_in22 = reg_0759;
    94: op1_04_in22 = reg_0830;
    95: op1_04_in22 = reg_0372;
    97: op1_04_in22 = reg_0968;
    98: op1_04_in22 = reg_0584;
    102: op1_04_in22 = reg_0840;
    103: op1_04_in22 = reg_0731;
    104: op1_04_in22 = reg_0119;
    105: op1_04_in22 = reg_0147;
    106: op1_04_in22 = reg_0075;
    107: op1_04_in22 = reg_0338;
    108: op1_04_in22 = reg_1147;
    109: op1_04_in22 = reg_0706;
    111: op1_04_in22 = reg_0209;
    113: op1_04_in22 = reg_0796;
    114: op1_04_in22 = reg_1450;
    115: op1_04_in22 = reg_0583;
    117: op1_04_in22 = reg_0397;
    118: op1_04_in22 = reg_0015;
    119: op1_04_in22 = reg_0779;
    120: op1_04_in22 = reg_0071;
    121: op1_04_in22 = reg_0227;
    122: op1_04_in22 = reg_0252;
    123: op1_04_in22 = reg_0897;
    124: op1_04_in22 = imem01_in[15:12];
    125: op1_04_in22 = reg_0498;
    126: op1_04_in22 = reg_1475;
    128: op1_04_in22 = reg_0053;
    129: op1_04_in22 = reg_0021;
    130: op1_04_in22 = reg_0130;
    131: op1_04_in22 = reg_0885;
    default: op1_04_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_04_inv22 = 1;
    61: op1_04_inv22 = 1;
    50: op1_04_inv22 = 1;
    71: op1_04_inv22 = 1;
    68: op1_04_inv22 = 1;
    74: op1_04_inv22 = 1;
    75: op1_04_inv22 = 1;
    87: op1_04_inv22 = 1;
    56: op1_04_inv22 = 1;
    46: op1_04_inv22 = 1;
    70: op1_04_inv22 = 1;
    88: op1_04_inv22 = 1;
    51: op1_04_inv22 = 1;
    59: op1_04_inv22 = 1;
    80: op1_04_inv22 = 1;
    62: op1_04_inv22 = 1;
    44: op1_04_inv22 = 1;
    82: op1_04_inv22 = 1;
    83: op1_04_inv22 = 1;
    84: op1_04_inv22 = 1;
    65: op1_04_inv22 = 1;
    91: op1_04_inv22 = 1;
    42: op1_04_inv22 = 1;
    92: op1_04_inv22 = 1;
    94: op1_04_inv22 = 1;
    95: op1_04_inv22 = 1;
    97: op1_04_inv22 = 1;
    98: op1_04_inv22 = 1;
    102: op1_04_inv22 = 1;
    103: op1_04_inv22 = 1;
    104: op1_04_inv22 = 1;
    105: op1_04_inv22 = 1;
    106: op1_04_inv22 = 1;
    108: op1_04_inv22 = 1;
    114: op1_04_inv22 = 1;
    115: op1_04_inv22 = 1;
    117: op1_04_inv22 = 1;
    123: op1_04_inv22 = 1;
    124: op1_04_inv22 = 1;
    125: op1_04_inv22 = 1;
    129: op1_04_inv22 = 1;
    130: op1_04_inv22 = 1;
    131: op1_04_inv22 = 1;
    default: op1_04_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in23 = reg_0089;
    53: op1_04_in23 = reg_0281;
    73: op1_04_in23 = reg_0261;
    86: op1_04_in23 = reg_0391;
    61: op1_04_in23 = reg_0430;
    80: op1_04_in23 = reg_0430;
    69: op1_04_in23 = reg_1132;
    50: op1_04_in23 = reg_0561;
    71: op1_04_in23 = reg_0010;
    68: op1_04_in23 = reg_0033;
    74: op1_04_in23 = reg_0788;
    75: op1_04_in23 = reg_0819;
    97: op1_04_in23 = reg_0819;
    87: op1_04_in23 = reg_0552;
    46: op1_04_in23 = reg_0903;
    60: op1_04_in23 = reg_0648;
    76: op1_04_in23 = reg_0260;
    48: op1_04_in23 = reg_0196;
    57: op1_04_in23 = reg_0321;
    77: op1_04_in23 = reg_0937;
    70: op1_04_in23 = reg_0288;
    52: op1_04_in23 = reg_1033;
    58: op1_04_in23 = reg_0745;
    78: op1_04_in23 = reg_0377;
    88: op1_04_in23 = reg_1282;
    51: op1_04_in23 = reg_0284;
    79: op1_04_in23 = reg_0371;
    104: op1_04_in23 = reg_0371;
    59: op1_04_in23 = reg_0154;
    62: op1_04_in23 = reg_1150;
    44: op1_04_in23 = reg_0602;
    81: op1_04_in23 = reg_1488;
    63: op1_04_in23 = reg_0175;
    124: op1_04_in23 = reg_0175;
    82: op1_04_in23 = reg_0820;
    89: op1_04_in23 = reg_0425;
    83: op1_04_in23 = reg_0520;
    47: op1_04_in23 = reg_0415;
    64: op1_04_in23 = reg_0527;
    84: op1_04_in23 = reg_0922;
    65: op1_04_in23 = reg_0638;
    85: op1_04_in23 = reg_0069;
    90: op1_04_in23 = reg_0438;
    66: op1_04_in23 = reg_1291;
    91: op1_04_in23 = reg_1258;
    42: op1_04_in23 = reg_0190;
    67: op1_04_in23 = reg_1269;
    92: op1_04_in23 = reg_0699;
    93: op1_04_in23 = reg_1447;
    94: op1_04_in23 = reg_0468;
    95: op1_04_in23 = reg_0585;
    96: op1_04_in23 = reg_0746;
    98: op1_04_in23 = reg_0571;
    99: op1_04_in23 = reg_0491;
    102: op1_04_in23 = reg_0573;
    103: op1_04_in23 = reg_1083;
    105: op1_04_in23 = reg_0360;
    106: op1_04_in23 = reg_0026;
    107: op1_04_in23 = reg_0339;
    108: op1_04_in23 = reg_0406;
    109: op1_04_in23 = reg_0216;
    111: op1_04_in23 = reg_0063;
    113: op1_04_in23 = reg_0471;
    114: op1_04_in23 = reg_0128;
    115: op1_04_in23 = reg_0977;
    117: op1_04_in23 = reg_0925;
    118: op1_04_in23 = reg_0498;
    119: op1_04_in23 = reg_0774;
    120: op1_04_in23 = reg_0058;
    121: op1_04_in23 = reg_0255;
    122: op1_04_in23 = reg_0181;
    123: op1_04_in23 = reg_0802;
    125: op1_04_in23 = reg_1057;
    126: op1_04_in23 = reg_1474;
    128: op1_04_in23 = reg_0004;
    129: op1_04_in23 = reg_0020;
    130: op1_04_in23 = reg_0118;
    131: op1_04_in23 = reg_1149;
    default: op1_04_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv23 = 1;
    53: op1_04_inv23 = 1;
    86: op1_04_inv23 = 1;
    71: op1_04_inv23 = 1;
    68: op1_04_inv23 = 1;
    74: op1_04_inv23 = 1;
    75: op1_04_inv23 = 1;
    60: op1_04_inv23 = 1;
    57: op1_04_inv23 = 1;
    77: op1_04_inv23 = 1;
    58: op1_04_inv23 = 1;
    88: op1_04_inv23 = 1;
    51: op1_04_inv23 = 1;
    79: op1_04_inv23 = 1;
    59: op1_04_inv23 = 1;
    89: op1_04_inv23 = 1;
    83: op1_04_inv23 = 1;
    47: op1_04_inv23 = 1;
    84: op1_04_inv23 = 1;
    67: op1_04_inv23 = 1;
    92: op1_04_inv23 = 1;
    93: op1_04_inv23 = 1;
    95: op1_04_inv23 = 1;
    96: op1_04_inv23 = 1;
    97: op1_04_inv23 = 1;
    98: op1_04_inv23 = 1;
    103: op1_04_inv23 = 1;
    106: op1_04_inv23 = 1;
    107: op1_04_inv23 = 1;
    108: op1_04_inv23 = 1;
    113: op1_04_inv23 = 1;
    114: op1_04_inv23 = 1;
    118: op1_04_inv23 = 1;
    119: op1_04_inv23 = 1;
    120: op1_04_inv23 = 1;
    122: op1_04_inv23 = 1;
    123: op1_04_inv23 = 1;
    124: op1_04_inv23 = 1;
    125: op1_04_inv23 = 1;
    131: op1_04_inv23 = 1;
    default: op1_04_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in24 = reg_0267;
    53: op1_04_in24 = reg_0276;
    73: op1_04_in24 = reg_1467;
    86: op1_04_in24 = reg_1181;
    61: op1_04_in24 = reg_0726;
    90: op1_04_in24 = reg_0726;
    69: op1_04_in24 = reg_0311;
    50: op1_04_in24 = reg_0495;
    71: op1_04_in24 = reg_0013;
    68: op1_04_in24 = reg_0793;
    74: op1_04_in24 = reg_1253;
    75: op1_04_in24 = reg_1457;
    87: op1_04_in24 = reg_0796;
    46: op1_04_in24 = reg_0708;
    60: op1_04_in24 = reg_0066;
    76: op1_04_in24 = reg_0966;
    48: op1_04_in24 = reg_0118;
    57: op1_04_in24 = reg_0519;
    77: op1_04_in24 = reg_1485;
    70: op1_04_in24 = reg_0707;
    52: op1_04_in24 = reg_0549;
    58: op1_04_in24 = reg_0317;
    78: op1_04_in24 = reg_1003;
    88: op1_04_in24 = reg_1280;
    51: op1_04_in24 = reg_0408;
    79: op1_04_in24 = reg_0067;
    115: op1_04_in24 = reg_0067;
    59: op1_04_in24 = reg_0279;
    80: op1_04_in24 = reg_0434;
    62: op1_04_in24 = reg_0461;
    44: op1_04_in24 = reg_0603;
    81: op1_04_in24 = reg_0370;
    63: op1_04_in24 = reg_0448;
    82: op1_04_in24 = reg_0468;
    89: op1_04_in24 = imem04_in[11:8];
    47: op1_04_in24 = reg_0413;
    64: op1_04_in24 = reg_0568;
    84: op1_04_in24 = reg_0225;
    65: op1_04_in24 = reg_0891;
    85: op1_04_in24 = reg_1515;
    121: op1_04_in24 = reg_1515;
    66: op1_04_in24 = reg_1255;
    91: op1_04_in24 = reg_0297;
    42: op1_04_in24 = imem07_in[15:12];
    67: op1_04_in24 = reg_0832;
    92: op1_04_in24 = reg_0154;
    93: op1_04_in24 = reg_0049;
    94: op1_04_in24 = reg_0146;
    95: op1_04_in24 = reg_0617;
    96: op1_04_in24 = reg_0612;
    97: op1_04_in24 = reg_0430;
    98: op1_04_in24 = reg_0979;
    99: op1_04_in24 = reg_1401;
    102: op1_04_in24 = reg_1033;
    103: op1_04_in24 = reg_1198;
    104: op1_04_in24 = reg_0215;
    105: op1_04_in24 = reg_0092;
    106: op1_04_in24 = reg_0005;
    107: op1_04_in24 = reg_1151;
    108: op1_04_in24 = reg_1065;
    109: op1_04_in24 = reg_0144;
    111: op1_04_in24 = reg_0065;
    113: op1_04_in24 = reg_0199;
    114: op1_04_in24 = reg_0876;
    117: op1_04_in24 = reg_1420;
    118: op1_04_in24 = reg_1095;
    119: op1_04_in24 = reg_0031;
    120: op1_04_in24 = reg_1322;
    122: op1_04_in24 = reg_1367;
    123: op1_04_in24 = reg_0801;
    124: op1_04_in24 = reg_0078;
    125: op1_04_in24 = reg_0457;
    126: op1_04_in24 = reg_0147;
    129: op1_04_in24 = reg_0210;
    130: op1_04_in24 = reg_1348;
    131: op1_04_in24 = reg_0559;
    default: op1_04_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_04_inv24 = 1;
    73: op1_04_inv24 = 1;
    86: op1_04_inv24 = 1;
    61: op1_04_inv24 = 1;
    50: op1_04_inv24 = 1;
    68: op1_04_inv24 = 1;
    75: op1_04_inv24 = 1;
    60: op1_04_inv24 = 1;
    48: op1_04_inv24 = 1;
    57: op1_04_inv24 = 1;
    58: op1_04_inv24 = 1;
    78: op1_04_inv24 = 1;
    59: op1_04_inv24 = 1;
    62: op1_04_inv24 = 1;
    81: op1_04_inv24 = 1;
    63: op1_04_inv24 = 1;
    47: op1_04_inv24 = 1;
    64: op1_04_inv24 = 1;
    65: op1_04_inv24 = 1;
    90: op1_04_inv24 = 1;
    66: op1_04_inv24 = 1;
    91: op1_04_inv24 = 1;
    42: op1_04_inv24 = 1;
    92: op1_04_inv24 = 1;
    94: op1_04_inv24 = 1;
    97: op1_04_inv24 = 1;
    98: op1_04_inv24 = 1;
    99: op1_04_inv24 = 1;
    104: op1_04_inv24 = 1;
    106: op1_04_inv24 = 1;
    109: op1_04_inv24 = 1;
    114: op1_04_inv24 = 1;
    119: op1_04_inv24 = 1;
    120: op1_04_inv24 = 1;
    122: op1_04_inv24 = 1;
    124: op1_04_inv24 = 1;
    130: op1_04_inv24 = 1;
    default: op1_04_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in25 = reg_1291;
    63: op1_04_in25 = reg_1291;
    53: op1_04_in25 = reg_0313;
    69: op1_04_in25 = reg_0313;
    73: op1_04_in25 = reg_1420;
    86: op1_04_in25 = reg_0794;
    61: op1_04_in25 = reg_0147;
    80: op1_04_in25 = reg_0147;
    50: op1_04_in25 = reg_0989;
    71: op1_04_in25 = reg_0457;
    68: op1_04_in25 = reg_0578;
    74: op1_04_in25 = reg_1254;
    75: op1_04_in25 = reg_0726;
    87: op1_04_in25 = reg_1147;
    46: op1_04_in25 = reg_0153;
    60: op1_04_in25 = reg_1181;
    76: op1_04_in25 = reg_0434;
    97: op1_04_in25 = reg_0434;
    48: op1_04_in25 = reg_0272;
    57: op1_04_in25 = reg_0521;
    77: op1_04_in25 = reg_0576;
    70: op1_04_in25 = imem03_in[3:0];
    52: op1_04_in25 = reg_0166;
    58: op1_04_in25 = reg_0367;
    78: op1_04_in25 = reg_0964;
    88: op1_04_in25 = reg_0427;
    51: op1_04_in25 = reg_0137;
    79: op1_04_in25 = reg_0023;
    59: op1_04_in25 = reg_0755;
    62: op1_04_in25 = imem07_in[3:0];
    44: op1_04_in25 = imem05_in[15:12];
    81: op1_04_in25 = reg_0708;
    82: op1_04_in25 = reg_0430;
    89: op1_04_in25 = reg_1312;
    47: op1_04_in25 = reg_0623;
    64: op1_04_in25 = reg_0571;
    84: op1_04_in25 = reg_0309;
    65: op1_04_in25 = reg_1001;
    85: op1_04_in25 = reg_1132;
    90: op1_04_in25 = reg_0383;
    66: op1_04_in25 = reg_0241;
    91: op1_04_in25 = reg_0552;
    42: op1_04_in25 = reg_0674;
    67: op1_04_in25 = reg_1212;
    92: op1_04_in25 = reg_1447;
    93: op1_04_in25 = reg_0261;
    94: op1_04_in25 = reg_0092;
    95: op1_04_in25 = reg_0215;
    96: op1_04_in25 = reg_0715;
    98: op1_04_in25 = reg_1228;
    99: op1_04_in25 = reg_0183;
    102: op1_04_in25 = reg_0198;
    103: op1_04_in25 = reg_0574;
    104: op1_04_in25 = reg_0213;
    105: op1_04_in25 = reg_0901;
    106: op1_04_in25 = reg_0980;
    107: op1_04_in25 = reg_0236;
    108: op1_04_in25 = reg_0097;
    109: op1_04_in25 = reg_0000;
    111: op1_04_in25 = reg_0370;
    113: op1_04_in25 = reg_1065;
    114: op1_04_in25 = reg_0829;
    115: op1_04_in25 = reg_0015;
    117: op1_04_in25 = reg_1437;
    118: op1_04_in25 = reg_0140;
    119: op1_04_in25 = reg_0404;
    120: op1_04_in25 = reg_0089;
    121: op1_04_in25 = reg_0480;
    122: op1_04_in25 = reg_0531;
    123: op1_04_in25 = reg_0255;
    124: op1_04_in25 = reg_0043;
    125: op1_04_in25 = reg_1350;
    126: op1_04_in25 = reg_0365;
    129: op1_04_in25 = imem05_in[3:0];
    130: op1_04_in25 = reg_0151;
    131: op1_04_in25 = reg_0218;
    default: op1_04_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv25 = 1;
    53: op1_04_inv25 = 1;
    73: op1_04_inv25 = 1;
    86: op1_04_inv25 = 1;
    68: op1_04_inv25 = 1;
    74: op1_04_inv25 = 1;
    87: op1_04_inv25 = 1;
    46: op1_04_inv25 = 1;
    60: op1_04_inv25 = 1;
    76: op1_04_inv25 = 1;
    77: op1_04_inv25 = 1;
    52: op1_04_inv25 = 1;
    78: op1_04_inv25 = 1;
    51: op1_04_inv25 = 1;
    81: op1_04_inv25 = 1;
    63: op1_04_inv25 = 1;
    89: op1_04_inv25 = 1;
    47: op1_04_inv25 = 1;
    64: op1_04_inv25 = 1;
    85: op1_04_inv25 = 1;
    66: op1_04_inv25 = 1;
    42: op1_04_inv25 = 1;
    67: op1_04_inv25 = 1;
    92: op1_04_inv25 = 1;
    95: op1_04_inv25 = 1;
    96: op1_04_inv25 = 1;
    98: op1_04_inv25 = 1;
    103: op1_04_inv25 = 1;
    104: op1_04_inv25 = 1;
    107: op1_04_inv25 = 1;
    108: op1_04_inv25 = 1;
    109: op1_04_inv25 = 1;
    115: op1_04_inv25 = 1;
    118: op1_04_inv25 = 1;
    120: op1_04_inv25 = 1;
    121: op1_04_inv25 = 1;
    123: op1_04_inv25 = 1;
    126: op1_04_inv25 = 1;
    131: op1_04_inv25 = 1;
    default: op1_04_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in26 = reg_1255;
    63: op1_04_in26 = reg_1255;
    53: op1_04_in26 = reg_0757;
    73: op1_04_in26 = reg_0160;
    86: op1_04_in26 = reg_0183;
    61: op1_04_in26 = reg_0360;
    69: op1_04_in26 = reg_0218;
    50: op1_04_in26 = reg_0971;
    71: op1_04_in26 = reg_1343;
    68: op1_04_in26 = reg_0315;
    74: op1_04_in26 = reg_0743;
    52: op1_04_in26 = reg_0743;
    75: op1_04_in26 = reg_0149;
    87: op1_04_in26 = reg_0421;
    46: op1_04_in26 = reg_0878;
    60: op1_04_in26 = reg_0697;
    76: op1_04_in26 = reg_0438;
    48: op1_04_in26 = imem06_in[15:12];
    77: op1_04_in26 = reg_0197;
    70: op1_04_in26 = reg_0704;
    58: op1_04_in26 = reg_0303;
    78: op1_04_in26 = reg_1517;
    88: op1_04_in26 = reg_1383;
    51: op1_04_in26 = reg_0103;
    79: op1_04_in26 = reg_0213;
    59: op1_04_in26 = reg_0678;
    80: op1_04_in26 = reg_0400;
    82: op1_04_in26 = reg_0400;
    105: op1_04_in26 = reg_0400;
    62: op1_04_in26 = reg_0894;
    44: op1_04_in26 = reg_0367;
    81: op1_04_in26 = reg_0175;
    89: op1_04_in26 = reg_0208;
    47: op1_04_in26 = reg_0591;
    64: op1_04_in26 = reg_0295;
    84: op1_04_in26 = reg_0489;
    65: op1_04_in26 = reg_0999;
    85: op1_04_in26 = reg_0312;
    90: op1_04_in26 = reg_0363;
    126: op1_04_in26 = reg_0363;
    66: op1_04_in26 = reg_0439;
    91: op1_04_in26 = reg_1215;
    42: op1_04_in26 = reg_0157;
    67: op1_04_in26 = reg_0745;
    92: op1_04_in26 = reg_0216;
    93: op1_04_in26 = reg_1063;
    94: op1_04_in26 = reg_0901;
    95: op1_04_in26 = reg_0214;
    96: op1_04_in26 = reg_0469;
    97: op1_04_in26 = reg_0868;
    98: op1_04_in26 = reg_0171;
    99: op1_04_in26 = reg_0302;
    102: op1_04_in26 = reg_1001;
    103: op1_04_in26 = reg_1200;
    104: op1_04_in26 = reg_1057;
    106: op1_04_in26 = reg_0282;
    107: op1_04_in26 = reg_0117;
    108: op1_04_in26 = reg_0698;
    109: op1_04_in26 = reg_0180;
    111: op1_04_in26 = reg_0708;
    113: op1_04_in26 = reg_0232;
    114: op1_04_in26 = reg_0294;
    115: op1_04_in26 = reg_0017;
    117: op1_04_in26 = reg_0718;
    118: op1_04_in26 = reg_0457;
    119: op1_04_in26 = reg_0592;
    120: op1_04_in26 = reg_1100;
    121: op1_04_in26 = reg_0179;
    122: op1_04_in26 = reg_0488;
    123: op1_04_in26 = reg_0840;
    124: op1_04_in26 = reg_0012;
    125: op1_04_in26 = reg_0139;
    129: op1_04_in26 = imem05_in[11:8];
    130: op1_04_in26 = reg_1431;
    131: op1_04_in26 = reg_0291;
    default: op1_04_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_04_inv26 = 1;
    86: op1_04_inv26 = 1;
    61: op1_04_inv26 = 1;
    69: op1_04_inv26 = 1;
    50: op1_04_inv26 = 1;
    71: op1_04_inv26 = 1;
    75: op1_04_inv26 = 1;
    87: op1_04_inv26 = 1;
    60: op1_04_inv26 = 1;
    70: op1_04_inv26 = 1;
    78: op1_04_inv26 = 1;
    51: op1_04_inv26 = 1;
    79: op1_04_inv26 = 1;
    59: op1_04_inv26 = 1;
    80: op1_04_inv26 = 1;
    62: op1_04_inv26 = 1;
    81: op1_04_inv26 = 1;
    84: op1_04_inv26 = 1;
    85: op1_04_inv26 = 1;
    90: op1_04_inv26 = 1;
    66: op1_04_inv26 = 1;
    67: op1_04_inv26 = 1;
    93: op1_04_inv26 = 1;
    94: op1_04_inv26 = 1;
    96: op1_04_inv26 = 1;
    97: op1_04_inv26 = 1;
    103: op1_04_inv26 = 1;
    104: op1_04_inv26 = 1;
    106: op1_04_inv26 = 1;
    108: op1_04_inv26 = 1;
    109: op1_04_inv26 = 1;
    111: op1_04_inv26 = 1;
    113: op1_04_inv26 = 1;
    114: op1_04_inv26 = 1;
    115: op1_04_inv26 = 1;
    118: op1_04_inv26 = 1;
    120: op1_04_inv26 = 1;
    124: op1_04_inv26 = 1;
    125: op1_04_inv26 = 1;
    131: op1_04_inv26 = 1;
    default: op1_04_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in27 = reg_1031;
    53: op1_04_in27 = reg_0756;
    73: op1_04_in27 = reg_0860;
    86: op1_04_in27 = reg_0300;
    99: op1_04_in27 = reg_0300;
    61: op1_04_in27 = reg_0899;
    97: op1_04_in27 = reg_0899;
    69: op1_04_in27 = reg_0198;
    50: op1_04_in27 = reg_0127;
    71: op1_04_in27 = reg_0497;
    68: op1_04_in27 = reg_0736;
    74: op1_04_in27 = reg_0609;
    75: op1_04_in27 = reg_0402;
    87: op1_04_in27 = reg_0412;
    46: op1_04_in27 = reg_0009;
    60: op1_04_in27 = reg_0317;
    76: op1_04_in27 = reg_0149;
    48: op1_04_in27 = reg_0960;
    77: op1_04_in27 = reg_0243;
    70: op1_04_in27 = reg_0185;
    52: op1_04_in27 = reg_0572;
    58: op1_04_in27 = reg_0251;
    78: op1_04_in27 = reg_1300;
    88: op1_04_in27 = reg_0032;
    51: op1_04_in27 = reg_0050;
    79: op1_04_in27 = reg_0022;
    59: op1_04_in27 = reg_0707;
    80: op1_04_in27 = reg_0363;
    62: op1_04_in27 = reg_0140;
    44: op1_04_in27 = reg_0090;
    81: op1_04_in27 = reg_0578;
    63: op1_04_in27 = reg_1034;
    82: op1_04_in27 = reg_0091;
    126: op1_04_in27 = reg_0091;
    89: op1_04_in27 = reg_0181;
    47: op1_04_in27 = reg_0002;
    64: op1_04_in27 = reg_1179;
    84: op1_04_in27 = reg_0777;
    65: op1_04_in27 = reg_0329;
    85: op1_04_in27 = reg_1494;
    90: op1_04_in27 = reg_0875;
    66: op1_04_in27 = reg_0434;
    91: op1_04_in27 = reg_1233;
    42: op1_04_in27 = reg_0169;
    67: op1_04_in27 = reg_0940;
    92: op1_04_in27 = reg_0312;
    102: op1_04_in27 = reg_0312;
    93: op1_04_in27 = reg_1033;
    94: op1_04_in27 = reg_0464;
    95: op1_04_in27 = reg_1170;
    115: op1_04_in27 = reg_1170;
    96: op1_04_in27 = reg_0438;
    98: op1_04_in27 = reg_0017;
    103: op1_04_in27 = reg_0281;
    104: op1_04_in27 = reg_0993;
    105: op1_04_in27 = reg_0042;
    106: op1_04_in27 = reg_1255;
    107: op1_04_in27 = reg_0209;
    108: op1_04_in27 = reg_0487;
    109: op1_04_in27 = reg_1495;
    111: op1_04_in27 = reg_0793;
    113: op1_04_in27 = reg_1312;
    114: op1_04_in27 = reg_0007;
    117: op1_04_in27 = reg_1303;
    118: op1_04_in27 = reg_0224;
    119: op1_04_in27 = imem07_in[15:12];
    120: op1_04_in27 = reg_1512;
    121: op1_04_in27 = reg_0177;
    122: op1_04_in27 = reg_0796;
    123: op1_04_in27 = reg_0989;
    124: op1_04_in27 = reg_0011;
    125: op1_04_in27 = reg_0029;
    129: op1_04_in27 = reg_0174;
    130: op1_04_in27 = reg_0475;
    131: op1_04_in27 = reg_0673;
    default: op1_04_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv27 = 1;
    53: op1_04_inv27 = 1;
    73: op1_04_inv27 = 1;
    61: op1_04_inv27 = 1;
    50: op1_04_inv27 = 1;
    71: op1_04_inv27 = 1;
    75: op1_04_inv27 = 1;
    46: op1_04_inv27 = 1;
    76: op1_04_inv27 = 1;
    52: op1_04_inv27 = 1;
    78: op1_04_inv27 = 1;
    88: op1_04_inv27 = 1;
    51: op1_04_inv27 = 1;
    79: op1_04_inv27 = 1;
    59: op1_04_inv27 = 1;
    62: op1_04_inv27 = 1;
    44: op1_04_inv27 = 1;
    81: op1_04_inv27 = 1;
    82: op1_04_inv27 = 1;
    84: op1_04_inv27 = 1;
    91: op1_04_inv27 = 1;
    93: op1_04_inv27 = 1;
    98: op1_04_inv27 = 1;
    104: op1_04_inv27 = 1;
    106: op1_04_inv27 = 1;
    113: op1_04_inv27 = 1;
    118: op1_04_inv27 = 1;
    121: op1_04_inv27 = 1;
    122: op1_04_inv27 = 1;
    123: op1_04_inv27 = 1;
    124: op1_04_inv27 = 1;
    125: op1_04_inv27 = 1;
    126: op1_04_inv27 = 1;
    129: op1_04_inv27 = 1;
    130: op1_04_inv27 = 1;
    default: op1_04_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in28 = reg_0547;
    53: op1_04_in28 = reg_0677;
    73: op1_04_in28 = imem06_in[7:4];
    86: op1_04_in28 = reg_0301;
    61: op1_04_in28 = reg_0077;
    69: op1_04_in28 = reg_0177;
    50: op1_04_in28 = reg_0898;
    71: op1_04_in28 = reg_0474;
    68: op1_04_in28 = reg_0735;
    74: op1_04_in28 = reg_0742;
    75: op1_04_in28 = reg_0403;
    87: op1_04_in28 = reg_0406;
    46: op1_04_in28 = reg_0801;
    60: op1_04_in28 = reg_0541;
    76: op1_04_in28 = reg_0384;
    48: op1_04_in28 = reg_0866;
    77: op1_04_in28 = reg_0631;
    70: op1_04_in28 = reg_1425;
    52: op1_04_in28 = reg_0727;
    58: op1_04_in28 = reg_0275;
    78: op1_04_in28 = reg_1231;
    88: op1_04_in28 = reg_1368;
    51: op1_04_in28 = reg_0052;
    79: op1_04_in28 = imem07_in[7:4];
    104: op1_04_in28 = imem07_in[7:4];
    59: op1_04_in28 = reg_1145;
    80: op1_04_in28 = reg_0088;
    62: op1_04_in28 = reg_0924;
    44: op1_04_in28 = reg_0872;
    81: op1_04_in28 = reg_0251;
    63: op1_04_in28 = reg_0549;
    82: op1_04_in28 = reg_0874;
    89: op1_04_in28 = reg_0034;
    47: op1_04_in28 = reg_0053;
    64: op1_04_in28 = reg_0046;
    84: op1_04_in28 = reg_0741;
    65: op1_04_in28 = reg_1226;
    85: op1_04_in28 = reg_0559;
    90: op1_04_in28 = reg_0464;
    66: op1_04_in28 = reg_0930;
    91: op1_04_in28 = reg_0796;
    103: op1_04_in28 = reg_0796;
    42: op1_04_in28 = reg_0779;
    118: op1_04_in28 = reg_0779;
    67: op1_04_in28 = reg_0937;
    92: op1_04_in28 = reg_0180;
    93: op1_04_in28 = reg_0600;
    94: op1_04_in28 = reg_0079;
    95: op1_04_in28 = reg_0230;
    96: op1_04_in28 = reg_0091;
    97: op1_04_in28 = reg_0901;
    126: op1_04_in28 = reg_0901;
    98: op1_04_in28 = imem07_in[3:0];
    99: op1_04_in28 = reg_0090;
    102: op1_04_in28 = reg_0144;
    105: op1_04_in28 = reg_0447;
    106: op1_04_in28 = reg_1253;
    107: op1_04_in28 = reg_0065;
    108: op1_04_in28 = reg_0835;
    109: op1_04_in28 = reg_1184;
    111: op1_04_in28 = reg_0832;
    113: op1_04_in28 = reg_1340;
    114: op1_04_in28 = reg_0217;
    115: op1_04_in28 = reg_1056;
    117: op1_04_in28 = reg_0374;
    120: op1_04_in28 = reg_1031;
    121: op1_04_in28 = reg_0000;
    122: op1_04_in28 = reg_1041;
    123: op1_04_in28 = reg_0233;
    124: op1_04_in28 = reg_0889;
    125: op1_04_in28 = reg_0030;
    129: op1_04_in28 = reg_0332;
    130: op1_04_in28 = reg_0974;
    131: op1_04_in28 = reg_0288;
    default: op1_04_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_04_inv28 = 1;
    86: op1_04_inv28 = 1;
    75: op1_04_inv28 = 1;
    46: op1_04_inv28 = 1;
    60: op1_04_inv28 = 1;
    76: op1_04_inv28 = 1;
    70: op1_04_inv28 = 1;
    52: op1_04_inv28 = 1;
    58: op1_04_inv28 = 1;
    78: op1_04_inv28 = 1;
    51: op1_04_inv28 = 1;
    59: op1_04_inv28 = 1;
    44: op1_04_inv28 = 1;
    89: op1_04_inv28 = 1;
    47: op1_04_inv28 = 1;
    85: op1_04_inv28 = 1;
    42: op1_04_inv28 = 1;
    67: op1_04_inv28 = 1;
    92: op1_04_inv28 = 1;
    97: op1_04_inv28 = 1;
    98: op1_04_inv28 = 1;
    99: op1_04_inv28 = 1;
    102: op1_04_inv28 = 1;
    105: op1_04_inv28 = 1;
    107: op1_04_inv28 = 1;
    109: op1_04_inv28 = 1;
    114: op1_04_inv28 = 1;
    118: op1_04_inv28 = 1;
    122: op1_04_inv28 = 1;
    124: op1_04_inv28 = 1;
    125: op1_04_inv28 = 1;
    131: op1_04_inv28 = 1;
    default: op1_04_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in29 = reg_0548;
    53: op1_04_in29 = reg_0288;
    73: op1_04_in29 = imem06_in[11:8];
    86: op1_04_in29 = reg_0197;
    44: op1_04_in29 = reg_0197;
    61: op1_04_in29 = reg_0277;
    69: op1_04_in29 = imem03_in[3:0];
    50: op1_04_in29 = reg_0900;
    71: op1_04_in29 = reg_0494;
    68: op1_04_in29 = reg_1269;
    74: op1_04_in29 = reg_0967;
    75: op1_04_in29 = reg_0385;
    87: op1_04_in29 = reg_1004;
    46: op1_04_in29 = reg_0279;
    60: op1_04_in29 = reg_0939;
    76: op1_04_in29 = reg_0360;
    52: op1_04_in29 = reg_0360;
    48: op1_04_in29 = reg_0373;
    77: op1_04_in29 = reg_0014;
    70: op1_04_in29 = reg_0640;
    58: op1_04_in29 = reg_1036;
    78: op1_04_in29 = reg_1208;
    65: op1_04_in29 = reg_1208;
    88: op1_04_in29 = reg_0034;
    51: op1_04_in29 = reg_0085;
    79: op1_04_in29 = reg_1440;
    59: op1_04_in29 = reg_0234;
    80: op1_04_in29 = reg_0278;
    111: op1_04_in29 = reg_0278;
    62: op1_04_in29 = reg_0224;
    81: op1_04_in29 = reg_1268;
    63: op1_04_in29 = reg_0746;
    82: op1_04_in29 = reg_0042;
    89: op1_04_in29 = reg_1257;
    47: op1_04_in29 = reg_0084;
    64: op1_04_in29 = reg_0212;
    84: op1_04_in29 = reg_0593;
    85: op1_04_in29 = reg_0185;
    90: op1_04_in29 = reg_0292;
    66: op1_04_in29 = reg_0726;
    91: op1_04_in29 = reg_1041;
    42: op1_04_in29 = reg_0774;
    67: op1_04_in29 = reg_0938;
    92: op1_04_in29 = reg_1003;
    93: op1_04_in29 = reg_0145;
    94: op1_04_in29 = reg_0257;
    95: op1_04_in29 = reg_0509;
    96: op1_04_in29 = reg_0092;
    97: op1_04_in29 = reg_0335;
    98: op1_04_in29 = reg_0324;
    99: op1_04_in29 = reg_0826;
    102: op1_04_in29 = reg_0965;
    103: op1_04_in29 = reg_0407;
    104: op1_04_in29 = imem07_in[15:12];
    105: op1_04_in29 = imem02_in[7:4];
    106: op1_04_in29 = reg_0576;
    107: op1_04_in29 = reg_0016;
    108: op1_04_in29 = reg_1189;
    109: op1_04_in29 = reg_1516;
    113: op1_04_in29 = reg_1151;
    114: op1_04_in29 = reg_0563;
    115: op1_04_in29 = reg_0225;
    117: op1_04_in29 = reg_0586;
    118: op1_04_in29 = reg_0030;
    120: op1_04_in29 = reg_0238;
    121: op1_04_in29 = reg_0891;
    122: op1_04_in29 = reg_0199;
    123: op1_04_in29 = reg_0557;
    124: op1_04_in29 = reg_0588;
    125: op1_04_in29 = reg_0739;
    126: op1_04_in29 = reg_0875;
    129: op1_04_in29 = reg_0346;
    130: op1_04_in29 = reg_0863;
    131: op1_04_in29 = reg_0790;
    default: op1_04_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_04_inv29 = 1;
    53: op1_04_inv29 = 1;
    86: op1_04_inv29 = 1;
    69: op1_04_inv29 = 1;
    50: op1_04_inv29 = 1;
    71: op1_04_inv29 = 1;
    68: op1_04_inv29 = 1;
    74: op1_04_inv29 = 1;
    87: op1_04_inv29 = 1;
    60: op1_04_inv29 = 1;
    48: op1_04_inv29 = 1;
    52: op1_04_inv29 = 1;
    58: op1_04_inv29 = 1;
    51: op1_04_inv29 = 1;
    79: op1_04_inv29 = 1;
    59: op1_04_inv29 = 1;
    80: op1_04_inv29 = 1;
    62: op1_04_inv29 = 1;
    44: op1_04_inv29 = 1;
    63: op1_04_inv29 = 1;
    47: op1_04_inv29 = 1;
    64: op1_04_inv29 = 1;
    65: op1_04_inv29 = 1;
    91: op1_04_inv29 = 1;
    42: op1_04_inv29 = 1;
    92: op1_04_inv29 = 1;
    94: op1_04_inv29 = 1;
    95: op1_04_inv29 = 1;
    96: op1_04_inv29 = 1;
    97: op1_04_inv29 = 1;
    104: op1_04_inv29 = 1;
    105: op1_04_inv29 = 1;
    108: op1_04_inv29 = 1;
    109: op1_04_inv29 = 1;
    111: op1_04_inv29 = 1;
    113: op1_04_inv29 = 1;
    115: op1_04_inv29 = 1;
    120: op1_04_inv29 = 1;
    122: op1_04_inv29 = 1;
    123: op1_04_inv29 = 1;
    125: op1_04_inv29 = 1;
    default: op1_04_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_04_in30 = reg_0787;
    53: op1_04_in30 = reg_1092;
    73: op1_04_in30 = reg_0116;
    86: op1_04_in30 = reg_0118;
    61: op1_04_in30 = reg_0446;
    69: op1_04_in30 = imem03_in[7:4];
    50: op1_04_in30 = reg_0879;
    71: op1_04_in30 = reg_0776;
    68: op1_04_in30 = imem05_in[11:8];
    74: op1_04_in30 = reg_0968;
    75: op1_04_in30 = reg_0365;
    87: op1_04_in30 = reg_0097;
    46: op1_04_in30 = reg_0276;
    60: op1_04_in30 = reg_0418;
    76: op1_04_in30 = reg_0091;
    48: op1_04_in30 = reg_0822;
    77: op1_04_in30 = reg_1168;
    70: op1_04_in30 = reg_1139;
    52: op1_04_in30 = reg_0868;
    58: op1_04_in30 = reg_0729;
    78: op1_04_in30 = reg_0113;
    88: op1_04_in30 = reg_0462;
    51: op1_04_in30 = reg_0084;
    79: op1_04_in30 = reg_0490;
    59: op1_04_in30 = reg_0000;
    80: op1_04_in30 = reg_0043;
    62: op1_04_in30 = reg_0779;
    44: op1_04_in30 = reg_0243;
    81: op1_04_in30 = reg_1163;
    63: op1_04_in30 = reg_0610;
    82: op1_04_in30 = reg_0662;
    89: op1_04_in30 = reg_1258;
    64: op1_04_in30 = reg_0191;
    84: op1_04_in30 = reg_0051;
    65: op1_04_in30 = reg_0107;
    85: op1_04_in30 = reg_0179;
    90: op1_04_in30 = reg_0162;
    66: op1_04_in30 = reg_0363;
    91: op1_04_in30 = reg_1065;
    42: op1_04_in30 = reg_0285;
    67: op1_04_in30 = reg_0575;
    92: op1_04_in30 = reg_0965;
    93: op1_04_in30 = reg_0180;
    94: op1_04_in30 = reg_0041;
    95: op1_04_in30 = imem07_in[3:0];
    96: op1_04_in30 = reg_0175;
    97: op1_04_in30 = reg_0724;
    98: op1_04_in30 = reg_0498;
    99: op1_04_in30 = reg_0784;
    102: op1_04_in30 = reg_0952;
    103: op1_04_in30 = reg_0471;
    104: op1_04_in30 = reg_0893;
    105: op1_04_in30 = imem02_in[11:8];
    106: op1_04_in30 = reg_0902;
    107: op1_04_in30 = reg_0035;
    108: op1_04_in30 = reg_0236;
    109: op1_04_in30 = reg_0190;
    111: op1_04_in30 = reg_0184;
    113: op1_04_in30 = reg_0932;
    114: op1_04_in30 = reg_0632;
    115: op1_04_in30 = reg_0457;
    117: op1_04_in30 = reg_0526;
    118: op1_04_in30 = reg_0284;
    120: op1_04_in30 = reg_0820;
    121: op1_04_in30 = reg_0556;
    122: op1_04_in30 = reg_0342;
    123: op1_04_in30 = reg_0783;
    124: op1_04_in30 = reg_0390;
    125: op1_04_in30 = reg_0404;
    126: op1_04_in30 = reg_0080;
    129: op1_04_in30 = reg_1059;
    130: op1_04_in30 = reg_0827;
    131: op1_04_in30 = reg_0348;
    default: op1_04_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_04_inv30 = 1;
    61: op1_04_inv30 = 1;
    50: op1_04_inv30 = 1;
    68: op1_04_inv30 = 1;
    74: op1_04_inv30 = 1;
    75: op1_04_inv30 = 1;
    87: op1_04_inv30 = 1;
    60: op1_04_inv30 = 1;
    76: op1_04_inv30 = 1;
    48: op1_04_inv30 = 1;
    58: op1_04_inv30 = 1;
    78: op1_04_inv30 = 1;
    79: op1_04_inv30 = 1;
    59: op1_04_inv30 = 1;
    80: op1_04_inv30 = 1;
    62: op1_04_inv30 = 1;
    81: op1_04_inv30 = 1;
    82: op1_04_inv30 = 1;
    89: op1_04_inv30 = 1;
    64: op1_04_inv30 = 1;
    90: op1_04_inv30 = 1;
    42: op1_04_inv30 = 1;
    67: op1_04_inv30 = 1;
    93: op1_04_inv30 = 1;
    95: op1_04_inv30 = 1;
    96: op1_04_inv30 = 1;
    98: op1_04_inv30 = 1;
    99: op1_04_inv30 = 1;
    102: op1_04_inv30 = 1;
    103: op1_04_inv30 = 1;
    107: op1_04_inv30 = 1;
    108: op1_04_inv30 = 1;
    109: op1_04_inv30 = 1;
    113: op1_04_inv30 = 1;
    114: op1_04_inv30 = 1;
    115: op1_04_inv30 = 1;
    121: op1_04_inv30 = 1;
    122: op1_04_inv30 = 1;
    123: op1_04_inv30 = 1;
    125: op1_04_inv30 = 1;
    131: op1_04_inv30 = 1;
    default: op1_04_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_04_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#4の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_04_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in00 = reg_0733;
    55: op1_05_in00 = reg_0022;
    53: op1_05_in00 = reg_0092;
    86: op1_05_in00 = reg_1301;
    80: op1_05_in00 = reg_1301;
    69: op1_05_in00 = reg_0403;
    73: op1_05_in00 = reg_0541;
    61: op1_05_in00 = reg_0748;
    85: op1_05_in00 = reg_0748;
    49: op1_05_in00 = reg_0998;
    50: op1_05_in00 = reg_0826;
    71: op1_05_in00 = reg_0555;
    54: op1_05_in00 = reg_0966;
    68: op1_05_in00 = reg_1325;
    74: op1_05_in00 = reg_0236;
    75: op1_05_in00 = reg_0370;
    56: op1_05_in00 = reg_0430;
    87: op1_05_in00 = reg_0710;
    76: op1_05_in00 = reg_1151;
    60: op1_05_in00 = reg_0480;
    46: op1_05_in00 = imem04_in[15:12];
    57: op1_05_in00 = reg_0374;
    77: op1_05_in00 = reg_1281;
    48: op1_05_in00 = reg_0596;
    33: op1_05_in00 = imem07_in[11:8];
    70: op1_05_in00 = reg_0896;
    58: op1_05_in00 = reg_0049;
    78: op1_05_in00 = reg_0347;
    88: op1_05_in00 = reg_1314;
    51: op1_05_in00 = reg_0930;
    79: op1_05_in00 = reg_1279;
    59: op1_05_in00 = reg_0308;
    28: op1_05_in00 = reg_0219;
    62: op1_05_in00 = reg_0669;
    52: op1_05_in00 = reg_0436;
    37: op1_05_in00 = reg_0158;
    81: op1_05_in00 = reg_1242;
    63: op1_05_in00 = reg_0148;
    82: op1_05_in00 = reg_0869;
    89: op1_05_in00 = reg_1149;
    22: op1_05_in00 = reg_0103;
    83: op1_05_in00 = reg_0907;
    64: op1_05_in00 = reg_1055;
    84: op1_05_in00 = reg_0616;
    47: op1_05_in00 = reg_0527;
    65: op1_05_in00 = reg_0627;
    40: op1_05_in00 = reg_0225;
    90: op1_05_in00 = reg_0048;
    66: op1_05_in00 = reg_0277;
    44: op1_05_in00 = reg_0421;
    91: op1_05_in00 = reg_0342;
    67: op1_05_in00 = reg_0151;
    92: op1_05_in00 = reg_0791;
    34: op1_05_in00 = reg_0223;
    93: op1_05_in00 = imem03_in[3:0];
    42: op1_05_in00 = reg_0201;
    94: op1_05_in00 = reg_0011;
    95: op1_05_in00 = reg_0922;
    96: op1_05_in00 = reg_0400;
    97: op1_05_in00 = reg_0257;
    98: op1_05_in00 = reg_0461;
    99: op1_05_in00 = reg_0192;
    100: op1_05_in00 = reg_0638;
    101: op1_05_in00 = reg_1469;
    102: op1_05_in00 = reg_1300;
    103: op1_05_in00 = reg_0599;
    104: op1_05_in00 = reg_0394;
    105: op1_05_in00 = imem02_in[15:12];
    106: op1_05_in00 = reg_0787;
    107: op1_05_in00 = reg_0213;
    108: op1_05_in00 = reg_0065;
    109: op1_05_in00 = reg_0378;
    110: op1_05_in00 = reg_0958;
    128: op1_05_in00 = reg_0958;
    111: op1_05_in00 = reg_0395;
    112: op1_05_in00 = reg_1277;
    113: op1_05_in00 = reg_0117;
    38: op1_05_in00 = reg_0159;
    114: op1_05_in00 = reg_0479;
    115: op1_05_in00 = reg_1347;
    116: op1_05_in00 = imem00_in[7:4];
    117: op1_05_in00 = reg_0528;
    118: op1_05_in00 = imem00_in[3:0];
    119: op1_05_in00 = imem00_in[15:12];
    120: op1_05_in00 = reg_1473;
    121: op1_05_in00 = reg_0964;
    122: op1_05_in00 = reg_1419;
    123: op1_05_in00 = reg_0823;
    124: op1_05_in00 = reg_0900;
    125: op1_05_in00 = reg_1243;
    126: op1_05_in00 = reg_0077;
    127: op1_05_in00 = reg_1490;
    129: op1_05_in00 = reg_0649;
    130: op1_05_in00 = reg_1179;
    29: op1_05_in00 = reg_0124;
    131: op1_05_in00 = reg_0443;
    default: op1_05_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_05_inv00 = 1;
    69: op1_05_inv00 = 1;
    73: op1_05_inv00 = 1;
    49: op1_05_inv00 = 1;
    71: op1_05_inv00 = 1;
    75: op1_05_inv00 = 1;
    56: op1_05_inv00 = 1;
    87: op1_05_inv00 = 1;
    76: op1_05_inv00 = 1;
    60: op1_05_inv00 = 1;
    33: op1_05_inv00 = 1;
    78: op1_05_inv00 = 1;
    88: op1_05_inv00 = 1;
    51: op1_05_inv00 = 1;
    28: op1_05_inv00 = 1;
    62: op1_05_inv00 = 1;
    52: op1_05_inv00 = 1;
    63: op1_05_inv00 = 1;
    82: op1_05_inv00 = 1;
    22: op1_05_inv00 = 1;
    64: op1_05_inv00 = 1;
    47: op1_05_inv00 = 1;
    85: op1_05_inv00 = 1;
    66: op1_05_inv00 = 1;
    44: op1_05_inv00 = 1;
    91: op1_05_inv00 = 1;
    34: op1_05_inv00 = 1;
    94: op1_05_inv00 = 1;
    95: op1_05_inv00 = 1;
    100: op1_05_inv00 = 1;
    104: op1_05_inv00 = 1;
    106: op1_05_inv00 = 1;
    107: op1_05_inv00 = 1;
    112: op1_05_inv00 = 1;
    38: op1_05_inv00 = 1;
    114: op1_05_inv00 = 1;
    117: op1_05_inv00 = 1;
    119: op1_05_inv00 = 1;
    120: op1_05_inv00 = 1;
    121: op1_05_inv00 = 1;
    122: op1_05_inv00 = 1;
    123: op1_05_inv00 = 1;
    125: op1_05_inv00 = 1;
    127: op1_05_inv00 = 1;
    128: op1_05_inv00 = 1;
    129: op1_05_inv00 = 1;
    130: op1_05_inv00 = 1;
    29: op1_05_inv00 = 1;
    default: op1_05_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in01 = reg_1163;
    55: op1_05_in01 = reg_0491;
    53: op1_05_in01 = reg_0093;
    86: op1_05_in01 = reg_1231;
    69: op1_05_in01 = reg_0401;
    73: op1_05_in01 = reg_0090;
    61: op1_05_in01 = reg_1277;
    49: op1_05_in01 = reg_0704;
    50: op1_05_in01 = reg_0825;
    57: op1_05_in01 = reg_0825;
    71: op1_05_in01 = reg_0580;
    54: op1_05_in01 = reg_0968;
    68: op1_05_in01 = reg_0145;
    74: op1_05_in01 = reg_0117;
    75: op1_05_in01 = reg_0750;
    56: op1_05_in01 = reg_0726;
    87: op1_05_in01 = reg_0444;
    76: op1_05_in01 = reg_1419;
    60: op1_05_in01 = reg_0790;
    46: op1_05_in01 = reg_0451;
    77: op1_05_in01 = reg_1079;
    48: op1_05_in01 = reg_0340;
    33: op1_05_in01 = imem07_in[15:12];
    70: op1_05_in01 = reg_0874;
    58: op1_05_in01 = reg_0232;
    78: op1_05_in01 = reg_1259;
    88: op1_05_in01 = reg_1313;
    51: op1_05_in01 = reg_0047;
    79: op1_05_in01 = reg_0218;
    59: op1_05_in01 = reg_0212;
    28: op1_05_in01 = reg_0084;
    80: op1_05_in01 = reg_1226;
    62: op1_05_in01 = reg_0842;
    52: op1_05_in01 = reg_0626;
    37: op1_05_in01 = reg_0029;
    22: op1_05_in01 = reg_0029;
    81: op1_05_in01 = reg_0615;
    100: op1_05_in01 = reg_0615;
    63: op1_05_in01 = reg_0386;
    82: op1_05_in01 = reg_0752;
    89: op1_05_in01 = reg_0480;
    83: op1_05_in01 = reg_1279;
    112: op1_05_in01 = reg_1279;
    64: op1_05_in01 = reg_0629;
    84: op1_05_in01 = reg_0907;
    127: op1_05_in01 = reg_0907;
    47: op1_05_in01 = reg_0308;
    65: op1_05_in01 = reg_0885;
    40: op1_05_in01 = reg_0190;
    85: op1_05_in01 = reg_0579;
    90: op1_05_in01 = reg_0104;
    66: op1_05_in01 = reg_0283;
    44: op1_05_in01 = reg_0796;
    91: op1_05_in01 = reg_0369;
    67: op1_05_in01 = reg_0861;
    92: op1_05_in01 = reg_1510;
    34: op1_05_in01 = reg_0324;
    93: op1_05_in01 = imem03_in[11:8];
    42: op1_05_in01 = imem00_in[11:8];
    94: op1_05_in01 = reg_1068;
    95: op1_05_in01 = reg_0892;
    96: op1_05_in01 = reg_0335;
    97: op1_05_in01 = reg_0896;
    98: op1_05_in01 = reg_0921;
    99: op1_05_in01 = reg_1420;
    101: op1_05_in01 = reg_1281;
    118: op1_05_in01 = reg_1281;
    102: op1_05_in01 = reg_0558;
    103: op1_05_in01 = reg_0452;
    104: op1_05_in01 = reg_0461;
    105: op1_05_in01 = reg_0169;
    106: op1_05_in01 = reg_0260;
    107: op1_05_in01 = reg_0015;
    108: op1_05_in01 = reg_0019;
    109: op1_05_in01 = reg_0025;
    110: op1_05_in01 = reg_0866;
    111: op1_05_in01 = reg_0251;
    113: op1_05_in01 = reg_0063;
    38: op1_05_in01 = reg_0158;
    114: op1_05_in01 = imem03_in[3:0];
    115: op1_05_in01 = reg_0159;
    116: op1_05_in01 = reg_1242;
    117: op1_05_in01 = reg_0529;
    119: op1_05_in01 = reg_1244;
    120: op1_05_in01 = reg_1474;
    121: op1_05_in01 = reg_0349;
    122: op1_05_in01 = reg_0837;
    123: op1_05_in01 = reg_0964;
    124: op1_05_in01 = reg_0495;
    125: op1_05_in01 = reg_0926;
    126: op1_05_in01 = reg_0079;
    128: op1_05_in01 = reg_0841;
    129: op1_05_in01 = reg_0300;
    130: op1_05_in01 = reg_0780;
    131: op1_05_in01 = reg_0411;
    default: op1_05_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv01 = 1;
    55: op1_05_inv01 = 1;
    53: op1_05_inv01 = 1;
    49: op1_05_inv01 = 1;
    71: op1_05_inv01 = 1;
    68: op1_05_inv01 = 1;
    74: op1_05_inv01 = 1;
    75: op1_05_inv01 = 1;
    46: op1_05_inv01 = 1;
    57: op1_05_inv01 = 1;
    77: op1_05_inv01 = 1;
    33: op1_05_inv01 = 1;
    88: op1_05_inv01 = 1;
    51: op1_05_inv01 = 1;
    59: op1_05_inv01 = 1;
    62: op1_05_inv01 = 1;
    52: op1_05_inv01 = 1;
    81: op1_05_inv01 = 1;
    63: op1_05_inv01 = 1;
    82: op1_05_inv01 = 1;
    89: op1_05_inv01 = 1;
    22: op1_05_inv01 = 1;
    83: op1_05_inv01 = 1;
    64: op1_05_inv01 = 1;
    47: op1_05_inv01 = 1;
    90: op1_05_inv01 = 1;
    91: op1_05_inv01 = 1;
    34: op1_05_inv01 = 1;
    42: op1_05_inv01 = 1;
    97: op1_05_inv01 = 1;
    98: op1_05_inv01 = 1;
    99: op1_05_inv01 = 1;
    100: op1_05_inv01 = 1;
    102: op1_05_inv01 = 1;
    103: op1_05_inv01 = 1;
    104: op1_05_inv01 = 1;
    105: op1_05_inv01 = 1;
    108: op1_05_inv01 = 1;
    109: op1_05_inv01 = 1;
    110: op1_05_inv01 = 1;
    111: op1_05_inv01 = 1;
    115: op1_05_inv01 = 1;
    116: op1_05_inv01 = 1;
    119: op1_05_inv01 = 1;
    122: op1_05_inv01 = 1;
    123: op1_05_inv01 = 1;
    124: op1_05_inv01 = 1;
    125: op1_05_inv01 = 1;
    126: op1_05_inv01 = 1;
    127: op1_05_inv01 = 1;
    128: op1_05_inv01 = 1;
    130: op1_05_inv01 = 1;
    default: op1_05_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in02 = reg_0996;
    55: op1_05_in02 = imem07_in[15:12];
    53: op1_05_in02 = reg_0724;
    86: op1_05_in02 = reg_1226;
    69: op1_05_in02 = reg_0360;
    73: op1_05_in02 = reg_0275;
    61: op1_05_in02 = reg_1079;
    49: op1_05_in02 = reg_0157;
    50: op1_05_in02 = reg_0716;
    71: op1_05_in02 = reg_0701;
    54: op1_05_in02 = reg_0819;
    68: op1_05_in02 = reg_0597;
    74: op1_05_in02 = imem04_in[7:4];
    75: op1_05_in02 = reg_1298;
    108: op1_05_in02 = reg_1298;
    56: op1_05_in02 = reg_0146;
    87: op1_05_in02 = reg_0706;
    76: op1_05_in02 = reg_0719;
    60: op1_05_in02 = reg_0426;
    46: op1_05_in02 = reg_0835;
    57: op1_05_in02 = reg_0718;
    77: op1_05_in02 = reg_1080;
    48: op1_05_in02 = reg_0305;
    33: op1_05_in02 = reg_0103;
    70: op1_05_in02 = reg_0283;
    58: op1_05_in02 = imem03_in[15:12];
    78: op1_05_in02 = reg_0176;
    88: op1_05_in02 = reg_1301;
    51: op1_05_in02 = reg_0871;
    79: op1_05_in02 = reg_1028;
    62: op1_05_in02 = reg_1028;
    59: op1_05_in02 = reg_0214;
    28: op1_05_in02 = reg_0053;
    80: op1_05_in02 = reg_0104;
    52: op1_05_in02 = reg_0934;
    37: op1_05_in02 = reg_0665;
    81: op1_05_in02 = reg_0485;
    63: op1_05_in02 = reg_0091;
    82: op1_05_in02 = reg_0780;
    89: op1_05_in02 = reg_1139;
    22: op1_05_in02 = imem07_in[3:0];
    83: op1_05_in02 = reg_1489;
    118: op1_05_in02 = reg_1489;
    64: op1_05_in02 = reg_0298;
    84: op1_05_in02 = reg_0640;
    47: op1_05_in02 = reg_0215;
    65: op1_05_in02 = reg_0505;
    40: op1_05_in02 = reg_0672;
    85: op1_05_in02 = reg_0833;
    90: op1_05_in02 = reg_0880;
    66: op1_05_in02 = reg_0041;
    44: op1_05_in02 = reg_0599;
    91: op1_05_in02 = reg_0698;
    67: op1_05_in02 = reg_0207;
    92: op1_05_in02 = reg_1487;
    34: op1_05_in02 = reg_0140;
    93: op1_05_in02 = reg_1516;
    42: op1_05_in02 = reg_0611;
    94: op1_05_in02 = reg_0666;
    95: op1_05_in02 = reg_0309;
    96: op1_05_in02 = reg_0078;
    97: op1_05_in02 = imem01_in[3:0];
    98: op1_05_in02 = reg_0924;
    99: op1_05_in02 = reg_0860;
    100: op1_05_in02 = reg_0153;
    101: op1_05_in02 = reg_1099;
    102: op1_05_in02 = reg_0107;
    103: op1_05_in02 = reg_1143;
    104: op1_05_in02 = reg_1415;
    105: op1_05_in02 = reg_0056;
    106: op1_05_in02 = reg_1475;
    107: op1_05_in02 = reg_0017;
    109: op1_05_in02 = reg_0673;
    110: op1_05_in02 = reg_1141;
    111: op1_05_in02 = reg_0831;
    112: op1_05_in02 = reg_0748;
    113: op1_05_in02 = reg_1502;
    38: op1_05_in02 = imem07_in[7:4];
    114: op1_05_in02 = imem03_in[7:4];
    115: op1_05_in02 = reg_0921;
    116: op1_05_in02 = reg_0843;
    117: op1_05_in02 = reg_0568;
    119: op1_05_in02 = reg_0248;
    120: op1_05_in02 = reg_1457;
    121: op1_05_in02 = reg_1313;
    122: op1_05_in02 = reg_1312;
    123: op1_05_in02 = reg_0558;
    124: op1_05_in02 = reg_0433;
    125: op1_05_in02 = reg_0806;
    128: op1_05_in02 = reg_0806;
    126: op1_05_in02 = reg_1071;
    127: op1_05_in02 = reg_1102;
    129: op1_05_in02 = reg_0333;
    130: op1_05_in02 = reg_0115;
    131: op1_05_in02 = reg_0016;
    default: op1_05_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_05_inv02 = 1;
    86: op1_05_inv02 = 1;
    73: op1_05_inv02 = 1;
    61: op1_05_inv02 = 1;
    54: op1_05_inv02 = 1;
    68: op1_05_inv02 = 1;
    76: op1_05_inv02 = 1;
    46: op1_05_inv02 = 1;
    57: op1_05_inv02 = 1;
    33: op1_05_inv02 = 1;
    70: op1_05_inv02 = 1;
    58: op1_05_inv02 = 1;
    78: op1_05_inv02 = 1;
    88: op1_05_inv02 = 1;
    79: op1_05_inv02 = 1;
    59: op1_05_inv02 = 1;
    80: op1_05_inv02 = 1;
    63: op1_05_inv02 = 1;
    89: op1_05_inv02 = 1;
    83: op1_05_inv02 = 1;
    64: op1_05_inv02 = 1;
    44: op1_05_inv02 = 1;
    67: op1_05_inv02 = 1;
    42: op1_05_inv02 = 1;
    94: op1_05_inv02 = 1;
    95: op1_05_inv02 = 1;
    96: op1_05_inv02 = 1;
    98: op1_05_inv02 = 1;
    99: op1_05_inv02 = 1;
    101: op1_05_inv02 = 1;
    102: op1_05_inv02 = 1;
    105: op1_05_inv02 = 1;
    106: op1_05_inv02 = 1;
    108: op1_05_inv02 = 1;
    109: op1_05_inv02 = 1;
    111: op1_05_inv02 = 1;
    113: op1_05_inv02 = 1;
    114: op1_05_inv02 = 1;
    115: op1_05_inv02 = 1;
    116: op1_05_inv02 = 1;
    118: op1_05_inv02 = 1;
    119: op1_05_inv02 = 1;
    121: op1_05_inv02 = 1;
    124: op1_05_inv02 = 1;
    125: op1_05_inv02 = 1;
    128: op1_05_inv02 = 1;
    default: op1_05_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in03 = reg_1180;
    55: op1_05_in03 = reg_0224;
    53: op1_05_in03 = reg_0899;
    86: op1_05_in03 = reg_0178;
    123: op1_05_in03 = reg_0178;
    69: op1_05_in03 = reg_0365;
    73: op1_05_in03 = reg_1346;
    61: op1_05_in03 = reg_0843;
    49: op1_05_in03 = imem07_in[15:12];
    28: op1_05_in03 = imem07_in[15:12];
    50: op1_05_in03 = reg_0714;
    71: op1_05_in03 = reg_0445;
    84: op1_05_in03 = reg_0445;
    54: op1_05_in03 = reg_0430;
    68: op1_05_in03 = reg_1301;
    74: op1_05_in03 = reg_0370;
    75: op1_05_in03 = reg_0136;
    56: op1_05_in03 = reg_0401;
    87: op1_05_in03 = reg_0378;
    76: op1_05_in03 = reg_0337;
    60: op1_05_in03 = reg_0247;
    46: op1_05_in03 = reg_0339;
    57: op1_05_in03 = reg_0635;
    77: op1_05_in03 = reg_0552;
    48: op1_05_in03 = reg_0862;
    33: op1_05_in03 = reg_0028;
    70: op1_05_in03 = reg_0222;
    58: op1_05_in03 = reg_0999;
    78: op1_05_in03 = reg_0174;
    88: op1_05_in03 = reg_1208;
    51: op1_05_in03 = reg_0042;
    79: op1_05_in03 = reg_1459;
    59: op1_05_in03 = reg_0185;
    80: op1_05_in03 = reg_0480;
    62: op1_05_in03 = reg_0492;
    52: op1_05_in03 = reg_0105;
    37: op1_05_in03 = reg_0661;
    81: op1_05_in03 = reg_0249;
    63: op1_05_in03 = reg_0724;
    82: op1_05_in03 = reg_0115;
    89: op1_05_in03 = reg_1280;
    22: op1_05_in03 = reg_0003;
    83: op1_05_in03 = reg_1491;
    64: op1_05_in03 = reg_1350;
    47: op1_05_in03 = reg_0213;
    65: op1_05_in03 = reg_0478;
    40: op1_05_in03 = imem07_in[11:8];
    85: op1_05_in03 = reg_1164;
    90: op1_05_in03 = imem03_in[7:4];
    66: op1_05_in03 = reg_0012;
    44: op1_05_in03 = imem04_in[11:8];
    91: op1_05_in03 = reg_0304;
    67: op1_05_in03 = reg_0206;
    92: op1_05_in03 = reg_0186;
    34: op1_05_in03 = reg_0465;
    93: op1_05_in03 = reg_1518;
    42: op1_05_in03 = reg_0612;
    94: op1_05_in03 = reg_0669;
    95: op1_05_in03 = reg_0489;
    96: op1_05_in03 = reg_0447;
    97: op1_05_in03 = imem01_in[11:8];
    120: op1_05_in03 = imem01_in[11:8];
    98: op1_05_in03 = reg_0923;
    99: op1_05_in03 = reg_0869;
    100: op1_05_in03 = reg_0486;
    101: op1_05_in03 = reg_1489;
    110: op1_05_in03 = reg_1489;
    102: op1_05_in03 = reg_0113;
    103: op1_05_in03 = reg_0837;
    104: op1_05_in03 = reg_0219;
    105: op1_05_in03 = reg_0608;
    106: op1_05_in03 = reg_0439;
    107: op1_05_in03 = imem07_in[7:4];
    108: op1_05_in03 = imem05_in[3:0];
    109: op1_05_in03 = reg_0288;
    111: op1_05_in03 = reg_0648;
    112: op1_05_in03 = reg_0907;
    118: op1_05_in03 = reg_0907;
    113: op1_05_in03 = reg_0470;
    38: op1_05_in03 = reg_0031;
    114: op1_05_in03 = reg_0732;
    115: op1_05_in03 = reg_0223;
    116: op1_05_in03 = reg_1279;
    117: op1_05_in03 = reg_0570;
    119: op1_05_in03 = reg_0638;
    121: op1_05_in03 = reg_0957;
    122: op1_05_in03 = reg_0256;
    124: op1_05_in03 = reg_0436;
    125: op1_05_in03 = reg_0615;
    126: op1_05_in03 = reg_0138;
    127: op1_05_in03 = reg_0523;
    128: op1_05_in03 = reg_0153;
    129: op1_05_in03 = reg_0601;
    130: op1_05_in03 = reg_0716;
    131: op1_05_in03 = reg_1338;
    default: op1_05_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_05_inv03 = 1;
    86: op1_05_inv03 = 1;
    69: op1_05_inv03 = 1;
    73: op1_05_inv03 = 1;
    61: op1_05_inv03 = 1;
    49: op1_05_inv03 = 1;
    50: op1_05_inv03 = 1;
    54: op1_05_inv03 = 1;
    68: op1_05_inv03 = 1;
    74: op1_05_inv03 = 1;
    75: op1_05_inv03 = 1;
    87: op1_05_inv03 = 1;
    76: op1_05_inv03 = 1;
    57: op1_05_inv03 = 1;
    77: op1_05_inv03 = 1;
    48: op1_05_inv03 = 1;
    70: op1_05_inv03 = 1;
    78: op1_05_inv03 = 1;
    79: op1_05_inv03 = 1;
    28: op1_05_inv03 = 1;
    62: op1_05_inv03 = 1;
    52: op1_05_inv03 = 1;
    63: op1_05_inv03 = 1;
    82: op1_05_inv03 = 1;
    89: op1_05_inv03 = 1;
    84: op1_05_inv03 = 1;
    65: op1_05_inv03 = 1;
    40: op1_05_inv03 = 1;
    85: op1_05_inv03 = 1;
    90: op1_05_inv03 = 1;
    66: op1_05_inv03 = 1;
    44: op1_05_inv03 = 1;
    67: op1_05_inv03 = 1;
    92: op1_05_inv03 = 1;
    34: op1_05_inv03 = 1;
    97: op1_05_inv03 = 1;
    98: op1_05_inv03 = 1;
    101: op1_05_inv03 = 1;
    105: op1_05_inv03 = 1;
    106: op1_05_inv03 = 1;
    109: op1_05_inv03 = 1;
    111: op1_05_inv03 = 1;
    112: op1_05_inv03 = 1;
    38: op1_05_inv03 = 1;
    115: op1_05_inv03 = 1;
    118: op1_05_inv03 = 1;
    119: op1_05_inv03 = 1;
    122: op1_05_inv03 = 1;
    126: op1_05_inv03 = 1;
    129: op1_05_inv03 = 1;
    131: op1_05_inv03 = 1;
    default: op1_05_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in04 = reg_0697;
    55: op1_05_in04 = reg_0703;
    53: op1_05_in04 = reg_0871;
    86: op1_05_in04 = reg_1208;
    123: op1_05_in04 = reg_1208;
    69: op1_05_in04 = reg_0091;
    73: op1_05_in04 = reg_0828;
    61: op1_05_in04 = reg_0803;
    49: op1_05_in04 = reg_0287;
    50: op1_05_in04 = reg_0635;
    71: op1_05_in04 = reg_1278;
    54: op1_05_in04 = reg_0726;
    68: op1_05_in04 = reg_1093;
    74: op1_05_in04 = reg_0578;
    75: op1_05_in04 = reg_0347;
    56: op1_05_in04 = reg_0092;
    87: op1_05_in04 = reg_0246;
    76: op1_05_in04 = imem04_in[3:0];
    60: op1_05_in04 = reg_0582;
    46: op1_05_in04 = reg_0336;
    57: op1_05_in04 = reg_0637;
    77: op1_05_in04 = reg_0562;
    48: op1_05_in04 = reg_0719;
    33: op1_05_in04 = reg_0050;
    70: op1_05_in04 = reg_0662;
    58: op1_05_in04 = reg_0963;
    78: op1_05_in04 = reg_0650;
    88: op1_05_in04 = reg_0113;
    51: op1_05_in04 = reg_0666;
    79: op1_05_in04 = reg_1227;
    59: op1_05_in04 = reg_0496;
    80: op1_05_in04 = reg_0481;
    62: op1_05_in04 = reg_0959;
    52: op1_05_in04 = reg_0900;
    37: op1_05_in04 = reg_0663;
    81: op1_05_in04 = reg_1206;
    63: op1_05_in04 = reg_0088;
    82: op1_05_in04 = reg_0109;
    89: op1_05_in04 = imem04_in[7:4];
    22: op1_05_in04 = reg_0085;
    83: op1_05_in04 = reg_0841;
    101: op1_05_in04 = reg_0841;
    64: op1_05_in04 = reg_0921;
    84: op1_05_in04 = reg_1489;
    47: op1_05_in04 = reg_0017;
    65: op1_05_in04 = reg_1280;
    40: op1_05_in04 = reg_0465;
    85: op1_05_in04 = reg_0701;
    90: op1_05_in04 = reg_0268;
    66: op1_05_in04 = reg_0013;
    44: op1_05_in04 = reg_0319;
    91: op1_05_in04 = reg_0319;
    67: op1_05_in04 = reg_0931;
    92: op1_05_in04 = reg_1053;
    128: op1_05_in04 = reg_1053;
    34: op1_05_in04 = reg_0030;
    93: op1_05_in04 = reg_1313;
    42: op1_05_in04 = reg_0695;
    94: op1_05_in04 = reg_0668;
    95: op1_05_in04 = reg_1094;
    98: op1_05_in04 = reg_1094;
    96: op1_05_in04 = reg_0475;
    97: op1_05_in04 = reg_0041;
    99: op1_05_in04 = reg_1505;
    100: op1_05_in04 = reg_0640;
    102: op1_05_in04 = reg_0378;
    103: op1_05_in04 = reg_0338;
    104: op1_05_in04 = reg_1440;
    105: op1_05_in04 = reg_0975;
    106: op1_05_in04 = reg_0868;
    107: op1_05_in04 = reg_1097;
    108: op1_05_in04 = reg_1431;
    109: op1_05_in04 = reg_0443;
    110: op1_05_in04 = reg_0613;
    112: op1_05_in04 = reg_0613;
    111: op1_05_in04 = reg_0066;
    113: op1_05_in04 = imem05_in[3:0];
    38: op1_05_in04 = reg_0665;
    114: op1_05_in04 = reg_0179;
    115: op1_05_in04 = reg_0779;
    116: op1_05_in04 = reg_0805;
    117: op1_05_in04 = reg_1228;
    118: op1_05_in04 = reg_0186;
    119: op1_05_in04 = reg_0748;
    120: op1_05_in04 = reg_0257;
    121: op1_05_in04 = reg_1447;
    122: op1_05_in04 = reg_1151;
    124: op1_05_in04 = reg_0054;
    125: op1_05_in04 = reg_0554;
    126: op1_05_in04 = reg_0497;
    127: op1_05_in04 = reg_0221;
    129: op1_05_in04 = reg_0393;
    130: op1_05_in04 = reg_0717;
    131: op1_05_in04 = reg_0236;
    default: op1_05_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv04 = 1;
    55: op1_05_inv04 = 1;
    53: op1_05_inv04 = 1;
    69: op1_05_inv04 = 1;
    73: op1_05_inv04 = 1;
    50: op1_05_inv04 = 1;
    75: op1_05_inv04 = 1;
    48: op1_05_inv04 = 1;
    78: op1_05_inv04 = 1;
    88: op1_05_inv04 = 1;
    51: op1_05_inv04 = 1;
    79: op1_05_inv04 = 1;
    59: op1_05_inv04 = 1;
    80: op1_05_inv04 = 1;
    62: op1_05_inv04 = 1;
    89: op1_05_inv04 = 1;
    22: op1_05_inv04 = 1;
    83: op1_05_inv04 = 1;
    64: op1_05_inv04 = 1;
    84: op1_05_inv04 = 1;
    66: op1_05_inv04 = 1;
    44: op1_05_inv04 = 1;
    91: op1_05_inv04 = 1;
    92: op1_05_inv04 = 1;
    34: op1_05_inv04 = 1;
    93: op1_05_inv04 = 1;
    94: op1_05_inv04 = 1;
    97: op1_05_inv04 = 1;
    99: op1_05_inv04 = 1;
    100: op1_05_inv04 = 1;
    101: op1_05_inv04 = 1;
    102: op1_05_inv04 = 1;
    104: op1_05_inv04 = 1;
    110: op1_05_inv04 = 1;
    115: op1_05_inv04 = 1;
    118: op1_05_inv04 = 1;
    119: op1_05_inv04 = 1;
    120: op1_05_inv04 = 1;
    121: op1_05_inv04 = 1;
    123: op1_05_inv04 = 1;
    124: op1_05_inv04 = 1;
    128: op1_05_inv04 = 1;
    129: op1_05_inv04 = 1;
    130: op1_05_inv04 = 1;
    131: op1_05_inv04 = 1;
    default: op1_05_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in05 = reg_0937;
    55: op1_05_in05 = reg_0892;
    53: op1_05_in05 = reg_0874;
    86: op1_05_in05 = reg_0108;
    69: op1_05_in05 = reg_0092;
    73: op1_05_in05 = reg_0206;
    61: op1_05_in05 = reg_1230;
    49: op1_05_in05 = reg_0285;
    50: op1_05_in05 = reg_0264;
    71: op1_05_in05 = imem00_in[15:12];
    54: op1_05_in05 = reg_0402;
    68: op1_05_in05 = reg_0107;
    74: op1_05_in05 = reg_1431;
    75: op1_05_in05 = reg_1168;
    56: op1_05_in05 = reg_0093;
    87: op1_05_in05 = reg_1208;
    76: op1_05_in05 = imem04_in[15:12];
    60: op1_05_in05 = reg_1146;
    46: op1_05_in05 = reg_0164;
    57: op1_05_in05 = reg_0323;
    77: op1_05_in05 = reg_0805;
    48: op1_05_in05 = reg_0339;
    33: op1_05_in05 = reg_0053;
    70: op1_05_in05 = reg_0744;
    58: op1_05_in05 = reg_0964;
    78: op1_05_in05 = reg_0333;
    88: op1_05_in05 = reg_0481;
    51: op1_05_in05 = reg_0256;
    79: op1_05_in05 = reg_1417;
    59: op1_05_in05 = reg_0461;
    80: op1_05_in05 = reg_0831;
    62: op1_05_in05 = reg_1148;
    52: op1_05_in05 = reg_0712;
    37: op1_05_in05 = reg_0664;
    38: op1_05_in05 = reg_0664;
    81: op1_05_in05 = reg_0351;
    63: op1_05_in05 = reg_0292;
    82: op1_05_in05 = reg_1302;
    89: op1_05_in05 = reg_0694;
    90: op1_05_in05 = reg_0694;
    22: op1_05_in05 = reg_0087;
    83: op1_05_in05 = reg_0615;
    64: op1_05_in05 = reg_0223;
    84: op1_05_in05 = reg_1487;
    47: op1_05_in05 = reg_0191;
    65: op1_05_in05 = reg_0247;
    40: op1_05_in05 = reg_0366;
    85: op1_05_in05 = reg_1181;
    66: op1_05_in05 = reg_0662;
    44: op1_05_in05 = reg_0262;
    91: op1_05_in05 = reg_0862;
    67: op1_05_in05 = reg_0860;
    92: op1_05_in05 = reg_0293;
    34: op1_05_in05 = imem07_in[7:4];
    93: op1_05_in05 = reg_0954;
    42: op1_05_in05 = reg_0819;
    94: op1_05_in05 = reg_0530;
    95: op1_05_in05 = reg_0740;
    96: op1_05_in05 = reg_0626;
    97: op1_05_in05 = reg_1068;
    98: op1_05_in05 = reg_0286;
    99: op1_05_in05 = reg_0372;
    100: op1_05_in05 = reg_1053;
    101: op1_05_in05 = reg_0640;
    110: op1_05_in05 = reg_0640;
    102: op1_05_in05 = reg_0025;
    103: op1_05_in05 = reg_0117;
    104: op1_05_in05 = reg_0225;
    105: op1_05_in05 = reg_0455;
    106: op1_05_in05 = reg_0360;
    107: op1_05_in05 = reg_0226;
    108: op1_05_in05 = reg_0466;
    109: op1_05_in05 = reg_0411;
    111: op1_05_in05 = reg_0566;
    112: op1_05_in05 = reg_0186;
    125: op1_05_in05 = reg_0186;
    113: op1_05_in05 = reg_0708;
    114: op1_05_in05 = reg_0709;
    115: op1_05_in05 = reg_0774;
    116: op1_05_in05 = reg_0486;
    117: op1_05_in05 = reg_0583;
    118: op1_05_in05 = reg_1027;
    128: op1_05_in05 = reg_1027;
    119: op1_05_in05 = reg_1099;
    120: op1_05_in05 = reg_0042;
    121: op1_05_in05 = imem03_in[11:8];
    122: op1_05_in05 = reg_1189;
    123: op1_05_in05 = reg_0113;
    124: op1_05_in05 = reg_0307;
    126: op1_05_in05 = reg_0898;
    127: op1_05_in05 = reg_1454;
    129: op1_05_in05 = reg_0344;
    130: op1_05_in05 = reg_0622;
    131: op1_05_in05 = reg_1258;
    default: op1_05_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_05_inv05 = 1;
    69: op1_05_inv05 = 1;
    73: op1_05_inv05 = 1;
    49: op1_05_inv05 = 1;
    71: op1_05_inv05 = 1;
    54: op1_05_inv05 = 1;
    75: op1_05_inv05 = 1;
    87: op1_05_inv05 = 1;
    76: op1_05_inv05 = 1;
    60: op1_05_inv05 = 1;
    70: op1_05_inv05 = 1;
    78: op1_05_inv05 = 1;
    88: op1_05_inv05 = 1;
    79: op1_05_inv05 = 1;
    80: op1_05_inv05 = 1;
    62: op1_05_inv05 = 1;
    81: op1_05_inv05 = 1;
    22: op1_05_inv05 = 1;
    83: op1_05_inv05 = 1;
    64: op1_05_inv05 = 1;
    84: op1_05_inv05 = 1;
    47: op1_05_inv05 = 1;
    40: op1_05_inv05 = 1;
    85: op1_05_inv05 = 1;
    66: op1_05_inv05 = 1;
    91: op1_05_inv05 = 1;
    67: op1_05_inv05 = 1;
    92: op1_05_inv05 = 1;
    94: op1_05_inv05 = 1;
    95: op1_05_inv05 = 1;
    96: op1_05_inv05 = 1;
    98: op1_05_inv05 = 1;
    99: op1_05_inv05 = 1;
    104: op1_05_inv05 = 1;
    105: op1_05_inv05 = 1;
    106: op1_05_inv05 = 1;
    107: op1_05_inv05 = 1;
    108: op1_05_inv05 = 1;
    109: op1_05_inv05 = 1;
    110: op1_05_inv05 = 1;
    111: op1_05_inv05 = 1;
    117: op1_05_inv05 = 1;
    118: op1_05_inv05 = 1;
    120: op1_05_inv05 = 1;
    121: op1_05_inv05 = 1;
    122: op1_05_inv05 = 1;
    123: op1_05_inv05 = 1;
    126: op1_05_inv05 = 1;
    127: op1_05_inv05 = 1;
    131: op1_05_inv05 = 1;
    default: op1_05_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in06 = reg_0167;
    55: op1_05_in06 = reg_0924;
    53: op1_05_in06 = reg_0080;
    86: op1_05_in06 = reg_0885;
    69: op1_05_in06 = reg_0896;
    73: op1_05_in06 = reg_1468;
    61: op1_05_in06 = reg_0202;
    49: op1_05_in06 = reg_0286;
    50: op1_05_in06 = reg_0528;
    71: op1_05_in06 = reg_0221;
    128: op1_05_in06 = reg_0221;
    54: op1_05_in06 = reg_0365;
    68: op1_05_in06 = reg_0113;
    74: op1_05_in06 = reg_0702;
    75: op1_05_in06 = reg_1164;
    56: op1_05_in06 = reg_0901;
    87: op1_05_in06 = reg_0104;
    123: op1_05_in06 = reg_0104;
    76: op1_05_in06 = reg_0065;
    46: op1_05_in06 = reg_0065;
    60: op1_05_in06 = imem04_in[15:12];
    57: op1_05_in06 = reg_0295;
    77: op1_05_in06 = reg_1053;
    48: op1_05_in06 = reg_0095;
    33: op1_05_in06 = reg_0085;
    70: op1_05_in06 = reg_1029;
    58: op1_05_in06 = reg_0952;
    93: op1_05_in06 = reg_0952;
    78: op1_05_in06 = reg_0567;
    88: op1_05_in06 = reg_0025;
    121: op1_05_in06 = reg_0025;
    51: op1_05_in06 = reg_0975;
    79: op1_05_in06 = reg_0524;
    59: op1_05_in06 = reg_0667;
    80: op1_05_in06 = reg_0734;
    62: op1_05_in06 = reg_0926;
    52: op1_05_in06 = reg_0876;
    37: op1_05_in06 = reg_0287;
    34: op1_05_in06 = reg_0287;
    81: op1_05_in06 = reg_0188;
    63: op1_05_in06 = reg_0043;
    82: op1_05_in06 = reg_0568;
    89: op1_05_in06 = reg_0341;
    83: op1_05_in06 = reg_0806;
    64: op1_05_in06 = reg_0777;
    84: op1_05_in06 = reg_0613;
    119: op1_05_in06 = reg_0613;
    47: op1_05_in06 = reg_0491;
    65: op1_05_in06 = reg_0534;
    40: op1_05_in06 = reg_0413;
    85: op1_05_in06 = reg_1403;
    90: op1_05_in06 = reg_0181;
    66: op1_05_in06 = reg_1103;
    44: op1_05_in06 = reg_0117;
    91: op1_05_in06 = reg_1189;
    67: op1_05_in06 = reg_0863;
    92: op1_05_in06 = reg_0821;
    42: op1_05_in06 = reg_0786;
    94: op1_05_in06 = reg_0169;
    95: op1_05_in06 = reg_0621;
    96: op1_05_in06 = reg_0399;
    97: op1_05_in06 = reg_0475;
    98: op1_05_in06 = reg_0441;
    99: op1_05_in06 = reg_0115;
    100: op1_05_in06 = reg_1459;
    101: op1_05_in06 = reg_0523;
    102: op1_05_in06 = reg_1325;
    103: op1_05_in06 = reg_0016;
    104: op1_05_in06 = reg_1349;
    105: op1_05_in06 = reg_0972;
    106: op1_05_in06 = reg_0363;
    107: op1_05_in06 = reg_0867;
    108: op1_05_in06 = reg_0332;
    109: op1_05_in06 = imem04_in[7:4];
    110: op1_05_in06 = reg_1028;
    112: op1_05_in06 = reg_1028;
    111: op1_05_in06 = reg_0697;
    113: op1_05_in06 = reg_0579;
    38: op1_05_in06 = reg_0284;
    114: op1_05_in06 = reg_0330;
    115: op1_05_in06 = reg_0285;
    116: op1_05_in06 = reg_0555;
    117: op1_05_in06 = reg_0022;
    118: op1_05_in06 = reg_1453;
    120: op1_05_in06 = reg_0010;
    122: op1_05_in06 = reg_0904;
    124: op1_05_in06 = reg_0829;
    125: op1_05_in06 = reg_0293;
    126: op1_05_in06 = reg_1458;
    127: op1_05_in06 = reg_1393;
    129: op1_05_in06 = reg_0861;
    130: op1_05_in06 = reg_0529;
    131: op1_05_in06 = reg_0978;
    default: op1_05_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_05_inv06 = 1;
    73: op1_05_inv06 = 1;
    61: op1_05_inv06 = 1;
    50: op1_05_inv06 = 1;
    75: op1_05_inv06 = 1;
    56: op1_05_inv06 = 1;
    76: op1_05_inv06 = 1;
    48: op1_05_inv06 = 1;
    78: op1_05_inv06 = 1;
    51: op1_05_inv06 = 1;
    79: op1_05_inv06 = 1;
    80: op1_05_inv06 = 1;
    52: op1_05_inv06 = 1;
    81: op1_05_inv06 = 1;
    63: op1_05_inv06 = 1;
    82: op1_05_inv06 = 1;
    89: op1_05_inv06 = 1;
    83: op1_05_inv06 = 1;
    64: op1_05_inv06 = 1;
    84: op1_05_inv06 = 1;
    90: op1_05_inv06 = 1;
    66: op1_05_inv06 = 1;
    91: op1_05_inv06 = 1;
    92: op1_05_inv06 = 1;
    93: op1_05_inv06 = 1;
    95: op1_05_inv06 = 1;
    97: op1_05_inv06 = 1;
    99: op1_05_inv06 = 1;
    100: op1_05_inv06 = 1;
    101: op1_05_inv06 = 1;
    102: op1_05_inv06 = 1;
    104: op1_05_inv06 = 1;
    105: op1_05_inv06 = 1;
    106: op1_05_inv06 = 1;
    108: op1_05_inv06 = 1;
    110: op1_05_inv06 = 1;
    111: op1_05_inv06 = 1;
    112: op1_05_inv06 = 1;
    115: op1_05_inv06 = 1;
    116: op1_05_inv06 = 1;
    117: op1_05_inv06 = 1;
    118: op1_05_inv06 = 1;
    119: op1_05_inv06 = 1;
    120: op1_05_inv06 = 1;
    124: op1_05_inv06 = 1;
    default: op1_05_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in07 = reg_0302;
    55: op1_05_in07 = reg_0284;
    37: op1_05_in07 = reg_0284;
    53: op1_05_in07 = reg_0290;
    86: op1_05_in07 = reg_0880;
    69: op1_05_in07 = reg_0277;
    73: op1_05_in07 = reg_1467;
    61: op1_05_in07 = reg_0492;
    49: op1_05_in07 = reg_0366;
    98: op1_05_in07 = reg_0366;
    50: op1_05_in07 = reg_0152;
    71: op1_05_in07 = reg_1227;
    100: op1_05_in07 = reg_1227;
    116: op1_05_in07 = reg_1227;
    54: op1_05_in07 = reg_0047;
    68: op1_05_in07 = reg_0882;
    74: op1_05_in07 = reg_0992;
    75: op1_05_in07 = reg_0346;
    56: op1_05_in07 = reg_0078;
    87: op1_05_in07 = reg_0479;
    76: op1_05_in07 = reg_1431;
    60: op1_05_in07 = reg_1203;
    46: op1_05_in07 = reg_0062;
    57: op1_05_in07 = reg_1204;
    77: op1_05_in07 = reg_0293;
    48: op1_05_in07 = reg_0164;
    70: op1_05_in07 = reg_0589;
    58: op1_05_in07 = reg_0448;
    78: op1_05_in07 = reg_1403;
    111: op1_05_in07 = reg_1403;
    88: op1_05_in07 = reg_1325;
    51: op1_05_in07 = reg_1029;
    66: op1_05_in07 = reg_1029;
    79: op1_05_in07 = reg_0821;
    110: op1_05_in07 = reg_0821;
    59: op1_05_in07 = reg_0668;
    80: op1_05_in07 = reg_0573;
    62: op1_05_in07 = reg_0435;
    52: op1_05_in07 = reg_0007;
    81: op1_05_in07 = reg_0722;
    63: op1_05_in07 = reg_0976;
    82: op1_05_in07 = reg_0569;
    89: op1_05_in07 = reg_1367;
    83: op1_05_in07 = reg_0805;
    64: op1_05_in07 = reg_0031;
    84: op1_05_in07 = reg_0580;
    47: op1_05_in07 = reg_0489;
    65: op1_05_in07 = imem04_in[7:4];
    102: op1_05_in07 = imem04_in[7:4];
    40: op1_05_in07 = reg_0102;
    85: op1_05_in07 = reg_1402;
    90: op1_05_in07 = reg_1368;
    44: op1_05_in07 = reg_0065;
    91: op1_05_in07 = reg_0932;
    122: op1_05_in07 = reg_0932;
    67: op1_05_in07 = reg_0133;
    92: op1_05_in07 = reg_0201;
    34: op1_05_in07 = reg_0413;
    93: op1_05_in07 = reg_0190;
    42: op1_05_in07 = reg_0549;
    94: op1_05_in07 = reg_0846;
    96: op1_05_in07 = reg_0846;
    95: op1_05_in07 = reg_0593;
    97: op1_05_in07 = reg_1260;
    99: op1_05_in07 = reg_0718;
    101: op1_05_in07 = reg_0987;
    118: op1_05_in07 = reg_0987;
    103: op1_05_in07 = reg_0877;
    104: op1_05_in07 = reg_0924;
    105: op1_05_in07 = reg_1451;
    106: op1_05_in07 = reg_0899;
    107: op1_05_in07 = reg_0994;
    108: op1_05_in07 = reg_0272;
    109: op1_05_in07 = reg_0181;
    112: op1_05_in07 = reg_0221;
    113: op1_05_in07 = reg_0183;
    38: op1_05_in07 = reg_0739;
    114: op1_05_in07 = reg_0198;
    115: op1_05_in07 = reg_0740;
    117: op1_05_in07 = reg_1170;
    119: op1_05_in07 = reg_0486;
    120: op1_05_in07 = reg_1068;
    121: op1_05_in07 = reg_0032;
    123: op1_05_in07 = reg_0885;
    124: op1_05_in07 = reg_0903;
    125: op1_05_in07 = reg_0485;
    126: op1_05_in07 = reg_1450;
    127: op1_05_in07 = reg_0886;
    128: op1_05_in07 = reg_0249;
    129: op1_05_in07 = reg_0565;
    130: op1_05_in07 = reg_0345;
    131: op1_05_in07 = reg_1083;
    default: op1_05_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_05_inv07 = 1;
    61: op1_05_inv07 = 1;
    49: op1_05_inv07 = 1;
    50: op1_05_inv07 = 1;
    71: op1_05_inv07 = 1;
    54: op1_05_inv07 = 1;
    74: op1_05_inv07 = 1;
    56: op1_05_inv07 = 1;
    76: op1_05_inv07 = 1;
    57: op1_05_inv07 = 1;
    58: op1_05_inv07 = 1;
    51: op1_05_inv07 = 1;
    79: op1_05_inv07 = 1;
    59: op1_05_inv07 = 1;
    37: op1_05_inv07 = 1;
    81: op1_05_inv07 = 1;
    82: op1_05_inv07 = 1;
    89: op1_05_inv07 = 1;
    65: op1_05_inv07 = 1;
    40: op1_05_inv07 = 1;
    90: op1_05_inv07 = 1;
    66: op1_05_inv07 = 1;
    44: op1_05_inv07 = 1;
    67: op1_05_inv07 = 1;
    34: op1_05_inv07 = 1;
    93: op1_05_inv07 = 1;
    94: op1_05_inv07 = 1;
    96: op1_05_inv07 = 1;
    97: op1_05_inv07 = 1;
    98: op1_05_inv07 = 1;
    102: op1_05_inv07 = 1;
    104: op1_05_inv07 = 1;
    106: op1_05_inv07 = 1;
    108: op1_05_inv07 = 1;
    109: op1_05_inv07 = 1;
    110: op1_05_inv07 = 1;
    111: op1_05_inv07 = 1;
    113: op1_05_inv07 = 1;
    38: op1_05_inv07 = 1;
    115: op1_05_inv07 = 1;
    117: op1_05_inv07 = 1;
    119: op1_05_inv07 = 1;
    120: op1_05_inv07 = 1;
    123: op1_05_inv07 = 1;
    126: op1_05_inv07 = 1;
    128: op1_05_inv07 = 1;
    129: op1_05_inv07 = 1;
    130: op1_05_inv07 = 1;
    131: op1_05_inv07 = 1;
    default: op1_05_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in08 = reg_0301;
    55: op1_05_in08 = reg_0285;
    53: op1_05_in08 = reg_0292;
    86: op1_05_in08 = reg_0505;
    69: op1_05_in08 = reg_0043;
    73: op1_05_in08 = reg_0795;
    61: op1_05_in08 = reg_1148;
    49: op1_05_in08 = reg_0415;
    115: op1_05_in08 = reg_0415;
    50: op1_05_in08 = reg_0213;
    71: op1_05_in08 = reg_0249;
    54: op1_05_in08 = reg_0724;
    68: op1_05_in08 = reg_0481;
    58: op1_05_in08 = reg_0481;
    74: op1_05_in08 = reg_0173;
    75: op1_05_in08 = reg_0303;
    56: op1_05_in08 = reg_0077;
    87: op1_05_in08 = reg_0313;
    76: op1_05_in08 = reg_1268;
    60: op1_05_in08 = reg_0574;
    46: op1_05_in08 = reg_0799;
    57: op1_05_in08 = reg_0583;
    77: op1_05_in08 = reg_1027;
    48: op1_05_in08 = reg_0211;
    70: op1_05_in08 = reg_0562;
    78: op1_05_in08 = reg_0939;
    88: op1_05_in08 = reg_1282;
    51: op1_05_in08 = reg_0455;
    79: op1_05_in08 = reg_0886;
    59: op1_05_in08 = reg_0673;
    80: op1_05_in08 = reg_0330;
    62: op1_05_in08 = reg_0405;
    52: op1_05_in08 = reg_0276;
    94: op1_05_in08 = reg_0276;
    37: op1_05_in08 = reg_0366;
    81: op1_05_in08 = reg_0388;
    63: op1_05_in08 = reg_0530;
    66: op1_05_in08 = reg_0530;
    82: op1_05_in08 = reg_0165;
    89: op1_05_in08 = reg_0264;
    67: op1_05_in08 = reg_0264;
    83: op1_05_in08 = reg_0218;
    64: op1_05_in08 = reg_0441;
    84: op1_05_in08 = reg_1469;
    47: op1_05_in08 = imem07_in[11:8];
    65: op1_05_in08 = reg_1338;
    40: op1_05_in08 = reg_0100;
    85: op1_05_in08 = reg_1401;
    90: op1_05_in08 = reg_0493;
    121: op1_05_in08 = reg_0493;
    44: op1_05_in08 = reg_0150;
    91: op1_05_in08 = reg_0063;
    92: op1_05_in08 = reg_0189;
    34: op1_05_in08 = reg_0623;
    38: op1_05_in08 = reg_0623;
    93: op1_05_in08 = reg_1199;
    42: op1_05_in08 = reg_0726;
    95: op1_05_in08 = reg_0591;
    96: op1_05_in08 = reg_0608;
    97: op1_05_in08 = reg_0472;
    98: op1_05_in08 = reg_0408;
    99: op1_05_in08 = reg_0717;
    100: op1_05_in08 = reg_1206;
    101: op1_05_in08 = reg_1432;
    102: op1_05_in08 = imem04_in[11:8];
    103: op1_05_in08 = reg_0579;
    104: op1_05_in08 = reg_0663;
    105: op1_05_in08 = reg_0111;
    106: op1_05_in08 = reg_0901;
    107: op1_05_in08 = reg_0667;
    108: op1_05_in08 = reg_0992;
    109: op1_05_in08 = reg_1367;
    110: op1_05_in08 = reg_0428;
    111: op1_05_in08 = reg_0266;
    112: op1_05_in08 = reg_1230;
    113: op1_05_in08 = reg_0793;
    114: op1_05_in08 = reg_0556;
    116: op1_05_in08 = reg_0987;
    117: op1_05_in08 = reg_1096;
    118: op1_05_in08 = reg_1418;
    119: op1_05_in08 = reg_1053;
    120: op1_05_in08 = reg_1071;
    122: op1_05_in08 = reg_0117;
    123: op1_05_in08 = reg_0025;
    124: op1_05_in08 = reg_1078;
    125: op1_05_in08 = reg_0821;
    126: op1_05_in08 = reg_0106;
    127: op1_05_in08 = reg_0353;
    128: op1_05_in08 = reg_0460;
    129: op1_05_in08 = reg_1299;
    130: op1_05_in08 = reg_0295;
    131: op1_05_in08 = reg_1215;
    default: op1_05_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_05_inv08 = 1;
    69: op1_05_inv08 = 1;
    73: op1_05_inv08 = 1;
    49: op1_05_inv08 = 1;
    50: op1_05_inv08 = 1;
    68: op1_05_inv08 = 1;
    74: op1_05_inv08 = 1;
    75: op1_05_inv08 = 1;
    56: op1_05_inv08 = 1;
    87: op1_05_inv08 = 1;
    46: op1_05_inv08 = 1;
    48: op1_05_inv08 = 1;
    58: op1_05_inv08 = 1;
    59: op1_05_inv08 = 1;
    80: op1_05_inv08 = 1;
    62: op1_05_inv08 = 1;
    52: op1_05_inv08 = 1;
    63: op1_05_inv08 = 1;
    82: op1_05_inv08 = 1;
    89: op1_05_inv08 = 1;
    90: op1_05_inv08 = 1;
    66: op1_05_inv08 = 1;
    91: op1_05_inv08 = 1;
    92: op1_05_inv08 = 1;
    34: op1_05_inv08 = 1;
    93: op1_05_inv08 = 1;
    95: op1_05_inv08 = 1;
    96: op1_05_inv08 = 1;
    97: op1_05_inv08 = 1;
    99: op1_05_inv08 = 1;
    101: op1_05_inv08 = 1;
    102: op1_05_inv08 = 1;
    103: op1_05_inv08 = 1;
    105: op1_05_inv08 = 1;
    107: op1_05_inv08 = 1;
    109: op1_05_inv08 = 1;
    38: op1_05_inv08 = 1;
    115: op1_05_inv08 = 1;
    118: op1_05_inv08 = 1;
    119: op1_05_inv08 = 1;
    121: op1_05_inv08 = 1;
    122: op1_05_inv08 = 1;
    125: op1_05_inv08 = 1;
    128: op1_05_inv08 = 1;
    130: op1_05_inv08 = 1;
    default: op1_05_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in09 = reg_0492;
    55: op1_05_in09 = reg_0441;
    53: op1_05_in09 = reg_0282;
    86: op1_05_in09 = reg_0507;
    69: op1_05_in09 = reg_0011;
    73: op1_05_in09 = reg_0908;
    61: op1_05_in09 = reg_0640;
    49: op1_05_in09 = reg_0618;
    115: op1_05_in09 = reg_0618;
    50: op1_05_in09 = reg_0017;
    71: op1_05_in09 = reg_1418;
    54: op1_05_in09 = reg_0868;
    68: op1_05_in09 = reg_0478;
    58: op1_05_in09 = reg_0478;
    74: op1_05_in09 = reg_0174;
    75: op1_05_in09 = reg_0274;
    56: op1_05_in09 = reg_0292;
    106: op1_05_in09 = reg_0292;
    87: op1_05_in09 = reg_1139;
    76: op1_05_in09 = reg_1169;
    60: op1_05_in09 = reg_0466;
    46: op1_05_in09 = reg_0575;
    57: op1_05_in09 = reg_1170;
    77: op1_05_in09 = reg_1453;
    48: op1_05_in09 = reg_0033;
    70: op1_05_in09 = reg_0473;
    78: op1_05_in09 = reg_0938;
    88: op1_05_in09 = reg_0426;
    51: op1_05_in09 = reg_0588;
    79: op1_05_in09 = reg_0188;
    59: op1_05_in09 = reg_0924;
    80: op1_05_in09 = reg_1280;
    62: op1_05_in09 = reg_0786;
    52: op1_05_in09 = imem03_in[7:4];
    37: op1_05_in09 = imem07_in[3:0];
    81: op1_05_in09 = reg_1068;
    63: op1_05_in09 = reg_0456;
    82: op1_05_in09 = reg_0583;
    89: op1_05_in09 = reg_1257;
    65: op1_05_in09 = reg_1257;
    83: op1_05_in09 = reg_0523;
    64: op1_05_in09 = reg_0740;
    84: op1_05_in09 = reg_0221;
    119: op1_05_in09 = reg_0221;
    47: op1_05_in09 = reg_0703;
    40: op1_05_in09 = reg_0228;
    85: op1_05_in09 = reg_1486;
    90: op1_05_in09 = reg_0535;
    66: op1_05_in09 = reg_0589;
    44: op1_05_in09 = reg_0210;
    91: op1_05_in09 = reg_1503;
    67: op1_05_in09 = reg_0116;
    92: op1_05_in09 = reg_0409;
    34: op1_05_in09 = reg_0593;
    93: op1_05_in09 = reg_1208;
    42: op1_05_in09 = reg_0715;
    94: op1_05_in09 = reg_1344;
    95: op1_05_in09 = reg_0103;
    96: op1_05_in09 = reg_0532;
    97: op1_05_in09 = reg_0971;
    98: op1_05_in09 = reg_0591;
    99: op1_05_in09 = reg_0528;
    100: op1_05_in09 = reg_0524;
    101: op1_05_in09 = reg_1417;
    102: op1_05_in09 = imem04_in[15:12];
    103: op1_05_in09 = reg_0347;
    104: op1_05_in09 = reg_0286;
    105: op1_05_in09 = reg_0629;
    107: op1_05_in09 = reg_0663;
    108: op1_05_in09 = reg_0066;
    109: op1_05_in09 = reg_0731;
    110: op1_05_in09 = reg_0431;
    111: op1_05_in09 = reg_1163;
    112: op1_05_in09 = reg_0881;
    113: op1_05_in09 = reg_0338;
    38: op1_05_in09 = reg_0321;
    114: op1_05_in09 = reg_0965;
    116: op1_05_in09 = reg_1201;
    117: op1_05_in09 = reg_0867;
    118: op1_05_in09 = reg_1405;
    120: op1_05_in09 = reg_0662;
    121: op1_05_in09 = reg_0264;
    122: op1_05_in09 = reg_0536;
    123: op1_05_in09 = reg_0218;
    124: op1_05_in09 = reg_1006;
    125: op1_05_in09 = reg_0883;
    126: op1_05_in09 = reg_0631;
    127: op1_05_in09 = reg_0352;
    128: op1_05_in09 = reg_0229;
    129: op1_05_in09 = reg_0172;
    130: op1_05_in09 = reg_0244;
    131: op1_05_in09 = reg_0500;
    default: op1_05_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_05_inv09 = 1;
    61: op1_05_inv09 = 1;
    71: op1_05_inv09 = 1;
    54: op1_05_inv09 = 1;
    74: op1_05_inv09 = 1;
    75: op1_05_inv09 = 1;
    56: op1_05_inv09 = 1;
    46: op1_05_inv09 = 1;
    57: op1_05_inv09 = 1;
    48: op1_05_inv09 = 1;
    78: op1_05_inv09 = 1;
    88: op1_05_inv09 = 1;
    79: op1_05_inv09 = 1;
    62: op1_05_inv09 = 1;
    81: op1_05_inv09 = 1;
    63: op1_05_inv09 = 1;
    82: op1_05_inv09 = 1;
    89: op1_05_inv09 = 1;
    84: op1_05_inv09 = 1;
    65: op1_05_inv09 = 1;
    40: op1_05_inv09 = 1;
    85: op1_05_inv09 = 1;
    90: op1_05_inv09 = 1;
    42: op1_05_inv09 = 1;
    95: op1_05_inv09 = 1;
    98: op1_05_inv09 = 1;
    99: op1_05_inv09 = 1;
    100: op1_05_inv09 = 1;
    104: op1_05_inv09 = 1;
    105: op1_05_inv09 = 1;
    107: op1_05_inv09 = 1;
    109: op1_05_inv09 = 1;
    110: op1_05_inv09 = 1;
    112: op1_05_inv09 = 1;
    113: op1_05_inv09 = 1;
    38: op1_05_inv09 = 1;
    117: op1_05_inv09 = 1;
    118: op1_05_inv09 = 1;
    119: op1_05_inv09 = 1;
    120: op1_05_inv09 = 1;
    121: op1_05_inv09 = 1;
    123: op1_05_inv09 = 1;
    127: op1_05_inv09 = 1;
    128: op1_05_inv09 = 1;
    130: op1_05_inv09 = 1;
    default: op1_05_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in10 = imem05_in[15:12];
    55: op1_05_in10 = reg_0437;
    53: op1_05_in10 = reg_0278;
    86: op1_05_in10 = reg_0481;
    69: op1_05_in10 = reg_0662;
    73: op1_05_in10 = reg_0925;
    61: op1_05_in10 = reg_0352;
    49: op1_05_in10 = reg_0591;
    64: op1_05_in10 = reg_0591;
    50: op1_05_in10 = reg_0393;
    71: op1_05_in10 = reg_0351;
    112: op1_05_in10 = reg_0351;
    54: op1_05_in10 = reg_0078;
    68: op1_05_in10 = imem03_in[15:12];
    74: op1_05_in10 = reg_0333;
    75: op1_05_in10 = reg_0118;
    56: op1_05_in10 = reg_0043;
    87: op1_05_in10 = reg_0288;
    76: op1_05_in10 = reg_0700;
    60: op1_05_in10 = reg_0412;
    46: op1_05_in10 = reg_0576;
    85: op1_05_in10 = reg_0576;
    57: op1_05_in10 = reg_1150;
    77: op1_05_in10 = reg_1230;
    48: op1_05_in10 = reg_0578;
    70: op1_05_in10 = imem02_in[15:12];
    58: op1_05_in10 = reg_0328;
    78: op1_05_in10 = reg_0275;
    88: op1_05_in10 = reg_0443;
    51: op1_05_in10 = reg_0589;
    79: op1_05_in10 = reg_0201;
    59: op1_05_in10 = reg_0774;
    80: op1_05_in10 = reg_1372;
    62: op1_05_in10 = reg_0822;
    52: op1_05_in10 = reg_0121;
    37: op1_05_in10 = imem07_in[15:12];
    81: op1_05_in10 = reg_0446;
    63: op1_05_in10 = imem02_in[3:0];
    82: op1_05_in10 = reg_0067;
    89: op1_05_in10 = reg_1233;
    83: op1_05_in10 = reg_0250;
    84: op1_05_in10 = reg_1229;
    47: op1_05_in10 = reg_0298;
    65: op1_05_in10 = reg_1258;
    109: op1_05_in10 = reg_1258;
    40: op1_05_in10 = reg_0051;
    90: op1_05_in10 = reg_0252;
    66: op1_05_in10 = reg_0587;
    44: op1_05_in10 = reg_0020;
    91: op1_05_in10 = reg_0347;
    67: op1_05_in10 = reg_0714;
    92: op1_05_in10 = reg_0073;
    34: op1_05_in10 = reg_0321;
    93: op1_05_in10 = reg_0218;
    42: op1_05_in10 = reg_0469;
    94: op1_05_in10 = reg_0497;
    96: op1_05_in10 = reg_0497;
    95: op1_05_in10 = reg_0084;
    97: op1_05_in10 = reg_0972;
    98: op1_05_in10 = reg_0519;
    99: op1_05_in10 = reg_0527;
    100: op1_05_in10 = reg_0821;
    101: op1_05_in10 = reg_0887;
    102: op1_05_in10 = reg_1340;
    103: op1_05_in10 = reg_0272;
    104: op1_05_in10 = reg_0621;
    105: op1_05_in10 = reg_0307;
    106: op1_05_in10 = imem01_in[7:4];
    107: op1_05_in10 = reg_0441;
    108: op1_05_in10 = reg_0392;
    110: op1_05_in10 = reg_0057;
    111: op1_05_in10 = reg_0301;
    113: op1_05_in10 = reg_1431;
    38: op1_05_in10 = reg_0050;
    114: op1_05_in10 = reg_0142;
    115: op1_05_in10 = reg_0102;
    116: op1_05_in10 = reg_1417;
    117: op1_05_in10 = reg_1183;
    118: op1_05_in10 = reg_0927;
    119: op1_05_in10 = reg_0485;
    120: op1_05_in10 = reg_0588;
    121: op1_05_in10 = reg_0731;
    122: op1_05_in10 = reg_1503;
    123: op1_05_in10 = reg_0208;
    124: op1_05_in10 = reg_0009;
    125: op1_05_in10 = reg_0886;
    126: op1_05_in10 = reg_0473;
    127: op1_05_in10 = reg_0188;
    128: op1_05_in10 = reg_1406;
    129: op1_05_in10 = imem06_in[3:0];
    130: op1_05_in10 = reg_1202;
    131: op1_05_in10 = reg_1082;
    default: op1_05_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv10 = 1;
    53: op1_05_inv10 = 1;
    86: op1_05_inv10 = 1;
    69: op1_05_inv10 = 1;
    61: op1_05_inv10 = 1;
    71: op1_05_inv10 = 1;
    54: op1_05_inv10 = 1;
    68: op1_05_inv10 = 1;
    74: op1_05_inv10 = 1;
    75: op1_05_inv10 = 1;
    76: op1_05_inv10 = 1;
    60: op1_05_inv10 = 1;
    46: op1_05_inv10 = 1;
    57: op1_05_inv10 = 1;
    77: op1_05_inv10 = 1;
    48: op1_05_inv10 = 1;
    78: op1_05_inv10 = 1;
    88: op1_05_inv10 = 1;
    51: op1_05_inv10 = 1;
    80: op1_05_inv10 = 1;
    52: op1_05_inv10 = 1;
    37: op1_05_inv10 = 1;
    81: op1_05_inv10 = 1;
    82: op1_05_inv10 = 1;
    89: op1_05_inv10 = 1;
    64: op1_05_inv10 = 1;
    84: op1_05_inv10 = 1;
    47: op1_05_inv10 = 1;
    65: op1_05_inv10 = 1;
    40: op1_05_inv10 = 1;
    85: op1_05_inv10 = 1;
    44: op1_05_inv10 = 1;
    91: op1_05_inv10 = 1;
    42: op1_05_inv10 = 1;
    94: op1_05_inv10 = 1;
    96: op1_05_inv10 = 1;
    98: op1_05_inv10 = 1;
    99: op1_05_inv10 = 1;
    100: op1_05_inv10 = 1;
    103: op1_05_inv10 = 1;
    106: op1_05_inv10 = 1;
    107: op1_05_inv10 = 1;
    108: op1_05_inv10 = 1;
    111: op1_05_inv10 = 1;
    112: op1_05_inv10 = 1;
    113: op1_05_inv10 = 1;
    38: op1_05_inv10 = 1;
    115: op1_05_inv10 = 1;
    118: op1_05_inv10 = 1;
    119: op1_05_inv10 = 1;
    124: op1_05_inv10 = 1;
    128: op1_05_inv10 = 1;
    129: op1_05_inv10 = 1;
    131: op1_05_inv10 = 1;
    default: op1_05_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in11 = reg_0206;
    55: op1_05_in11 = reg_0738;
    53: op1_05_in11 = reg_0043;
    86: op1_05_in11 = imem03_in[11:8];
    69: op1_05_in11 = reg_0976;
    73: op1_05_in11 = reg_0860;
    61: op1_05_in11 = reg_0122;
    49: op1_05_in11 = reg_0102;
    50: op1_05_in11 = reg_0135;
    71: op1_05_in11 = reg_0352;
    54: op1_05_in11 = reg_0077;
    68: op1_05_in11 = reg_0840;
    58: op1_05_in11 = reg_0840;
    74: op1_05_in11 = reg_0567;
    75: op1_05_in11 = reg_0631;
    56: op1_05_in11 = reg_0679;
    87: op1_05_in11 = reg_0443;
    76: op1_05_in11 = reg_0650;
    60: op1_05_in11 = reg_0406;
    46: op1_05_in11 = reg_0748;
    57: op1_05_in11 = reg_1097;
    77: op1_05_in11 = reg_1229;
    48: op1_05_in11 = imem05_in[11:8];
    70: op1_05_in11 = reg_0820;
    78: op1_05_in11 = reg_1373;
    88: op1_05_in11 = reg_0088;
    51: op1_05_in11 = reg_0531;
    79: op1_05_in11 = reg_0189;
    59: op1_05_in11 = reg_0665;
    80: op1_05_in11 = reg_0493;
    62: op1_05_in11 = reg_0785;
    52: op1_05_in11 = reg_0630;
    37: op1_05_in11 = reg_0408;
    81: op1_05_in11 = reg_0963;
    63: op1_05_in11 = imem02_in[11:8];
    82: op1_05_in11 = reg_0214;
    89: op1_05_in11 = reg_1214;
    83: op1_05_in11 = reg_0293;
    84: op1_05_in11 = reg_1206;
    47: op1_05_in11 = reg_0158;
    65: op1_05_in11 = reg_1203;
    85: op1_05_in11 = reg_0492;
    90: op1_05_in11 = reg_1338;
    66: op1_05_in11 = reg_0255;
    44: op1_05_in11 = reg_0579;
    91: op1_05_in11 = reg_1169;
    67: op1_05_in11 = reg_1302;
    92: op1_05_in11 = reg_0057;
    34: op1_05_in11 = reg_0087;
    93: op1_05_in11 = reg_0313;
    42: op1_05_in11 = reg_0572;
    94: op1_05_in11 = reg_0495;
    95: op1_05_in11 = reg_0520;
    96: op1_05_in11 = reg_0472;
    97: op1_05_in11 = reg_0629;
    99: op1_05_in11 = reg_0345;
    100: op1_05_in11 = reg_1405;
    101: op1_05_in11 = reg_0351;
    102: op1_05_in11 = reg_0467;
    103: op1_05_in11 = reg_0251;
    104: op1_05_in11 = reg_0592;
    105: op1_05_in11 = reg_0473;
    106: op1_05_in11 = reg_0900;
    107: op1_05_in11 = reg_0739;
    108: op1_05_in11 = reg_0491;
    109: op1_05_in11 = reg_0462;
    110: op1_05_in11 = imem01_in[11:8];
    111: op1_05_in11 = reg_0888;
    112: op1_05_in11 = reg_0722;
    113: op1_05_in11 = reg_0136;
    38: op1_05_in11 = reg_0003;
    114: op1_05_in11 = reg_1313;
    115: op1_05_in11 = reg_0103;
    116: op1_05_in11 = reg_0155;
    117: op1_05_in11 = reg_1010;
    118: op1_05_in11 = reg_0887;
    119: op1_05_in11 = reg_1230;
    120: op1_05_in11 = reg_0712;
    121: op1_05_in11 = reg_0797;
    122: op1_05_in11 = reg_0016;
    123: op1_05_in11 = reg_0164;
    124: op1_05_in11 = reg_0049;
    125: op1_05_in11 = reg_0071;
    126: op1_05_in11 = reg_1091;
    127: op1_05_in11 = reg_0073;
    128: op1_05_in11 = reg_0821;
    129: op1_05_in11 = reg_0475;
    130: op1_05_in11 = reg_0754;
    131: op1_05_in11 = reg_0412;
    default: op1_05_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv11 = 1;
    55: op1_05_inv11 = 1;
    53: op1_05_inv11 = 1;
    69: op1_05_inv11 = 1;
    73: op1_05_inv11 = 1;
    61: op1_05_inv11 = 1;
    49: op1_05_inv11 = 1;
    50: op1_05_inv11 = 1;
    71: op1_05_inv11 = 1;
    54: op1_05_inv11 = 1;
    68: op1_05_inv11 = 1;
    74: op1_05_inv11 = 1;
    75: op1_05_inv11 = 1;
    56: op1_05_inv11 = 1;
    60: op1_05_inv11 = 1;
    46: op1_05_inv11 = 1;
    77: op1_05_inv11 = 1;
    70: op1_05_inv11 = 1;
    78: op1_05_inv11 = 1;
    88: op1_05_inv11 = 1;
    79: op1_05_inv11 = 1;
    59: op1_05_inv11 = 1;
    80: op1_05_inv11 = 1;
    62: op1_05_inv11 = 1;
    81: op1_05_inv11 = 1;
    63: op1_05_inv11 = 1;
    82: op1_05_inv11 = 1;
    89: op1_05_inv11 = 1;
    84: op1_05_inv11 = 1;
    85: op1_05_inv11 = 1;
    44: op1_05_inv11 = 1;
    91: op1_05_inv11 = 1;
    67: op1_05_inv11 = 1;
    34: op1_05_inv11 = 1;
    94: op1_05_inv11 = 1;
    95: op1_05_inv11 = 1;
    96: op1_05_inv11 = 1;
    97: op1_05_inv11 = 1;
    102: op1_05_inv11 = 1;
    103: op1_05_inv11 = 1;
    104: op1_05_inv11 = 1;
    105: op1_05_inv11 = 1;
    106: op1_05_inv11 = 1;
    38: op1_05_inv11 = 1;
    114: op1_05_inv11 = 1;
    115: op1_05_inv11 = 1;
    117: op1_05_inv11 = 1;
    119: op1_05_inv11 = 1;
    121: op1_05_inv11 = 1;
    122: op1_05_inv11 = 1;
    124: op1_05_inv11 = 1;
    126: op1_05_inv11 = 1;
    128: op1_05_inv11 = 1;
    129: op1_05_inv11 = 1;
    default: op1_05_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in12 = reg_0039;
    78: op1_05_in12 = reg_0039;
    55: op1_05_in12 = reg_0413;
    53: op1_05_in12 = reg_0041;
    86: op1_05_in12 = reg_1139;
    69: op1_05_in12 = reg_0605;
    73: op1_05_in12 = imem06_in[15:12];
    61: op1_05_in12 = reg_0026;
    49: op1_05_in12 = reg_0321;
    50: op1_05_in12 = imem07_in[3:0];
    82: op1_05_in12 = imem07_in[3:0];
    71: op1_05_in12 = reg_0387;
    54: op1_05_in12 = reg_0282;
    68: op1_05_in12 = reg_0330;
    74: op1_05_in12 = reg_0566;
    75: op1_05_in12 = reg_0589;
    56: op1_05_in12 = reg_0606;
    87: op1_05_in12 = reg_0411;
    76: op1_05_in12 = reg_0565;
    60: op1_05_in12 = reg_0795;
    46: op1_05_in12 = reg_0345;
    57: op1_05_in12 = reg_1094;
    77: op1_05_in12 = reg_1406;
    48: op1_05_in12 = reg_0649;
    70: op1_05_in12 = reg_0068;
    58: op1_05_in12 = reg_0048;
    88: op1_05_in12 = reg_1340;
    51: op1_05_in12 = reg_0496;
    97: op1_05_in12 = reg_0496;
    79: op1_05_in12 = reg_0405;
    59: op1_05_in12 = reg_0661;
    80: op1_05_in12 = reg_1257;
    121: op1_05_in12 = reg_1257;
    62: op1_05_in12 = reg_0335;
    52: op1_05_in12 = reg_1092;
    37: op1_05_in12 = reg_0618;
    81: op1_05_in12 = reg_0258;
    63: op1_05_in12 = reg_0472;
    89: op1_05_in12 = reg_0406;
    83: op1_05_in12 = reg_1227;
    84: op1_05_in12 = reg_0961;
    47: op1_05_in12 = reg_0169;
    65: op1_05_in12 = reg_1198;
    109: op1_05_in12 = reg_1198;
    85: op1_05_in12 = reg_0393;
    90: op1_05_in12 = reg_1203;
    66: op1_05_in12 = reg_0497;
    44: op1_05_in12 = reg_0391;
    91: op1_05_in12 = reg_0831;
    67: op1_05_in12 = reg_0636;
    92: op1_05_in12 = reg_0723;
    34: op1_05_in12 = reg_0519;
    93: op1_05_in12 = reg_1282;
    42: op1_05_in12 = reg_0430;
    94: op1_05_in12 = reg_0971;
    95: op1_05_in12 = reg_0483;
    96: op1_05_in12 = reg_0970;
    99: op1_05_in12 = reg_1225;
    100: op1_05_in12 = reg_0928;
    101: op1_05_in12 = reg_0352;
    102: op1_05_in12 = reg_1368;
    103: op1_05_in12 = reg_0648;
    104: op1_05_in12 = reg_0102;
    105: op1_05_in12 = reg_0379;
    106: op1_05_in12 = reg_0607;
    107: op1_05_in12 = reg_0100;
    108: op1_05_in12 = reg_0167;
    110: op1_05_in12 = reg_0635;
    111: op1_05_in12 = reg_0130;
    112: op1_05_in12 = reg_0440;
    113: op1_05_in12 = reg_0733;
    38: op1_05_in12 = reg_0001;
    114: op1_05_in12 = reg_0954;
    115: op1_05_in12 = reg_0114;
    116: op1_05_in12 = reg_0459;
    117: op1_05_in12 = reg_1315;
    118: op1_05_in12 = reg_0202;
    119: op1_05_in12 = reg_0460;
    120: op1_05_in12 = reg_0390;
    122: op1_05_in12 = reg_1298;
    123: op1_05_in12 = reg_0032;
    124: op1_05_in12 = reg_1003;
    125: op1_05_in12 = reg_0073;
    126: op1_05_in12 = imem03_in[15:12];
    127: op1_05_in12 = reg_0075;
    128: op1_05_in12 = reg_0881;
    129: op1_05_in12 = reg_0397;
    130: op1_05_in12 = reg_0067;
    131: op1_05_in12 = reg_0471;
    default: op1_05_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv12 = 1;
    55: op1_05_inv12 = 1;
    53: op1_05_inv12 = 1;
    86: op1_05_inv12 = 1;
    73: op1_05_inv12 = 1;
    50: op1_05_inv12 = 1;
    54: op1_05_inv12 = 1;
    75: op1_05_inv12 = 1;
    56: op1_05_inv12 = 1;
    46: op1_05_inv12 = 1;
    70: op1_05_inv12 = 1;
    78: op1_05_inv12 = 1;
    51: op1_05_inv12 = 1;
    52: op1_05_inv12 = 1;
    89: op1_05_inv12 = 1;
    83: op1_05_inv12 = 1;
    47: op1_05_inv12 = 1;
    85: op1_05_inv12 = 1;
    44: op1_05_inv12 = 1;
    91: op1_05_inv12 = 1;
    67: op1_05_inv12 = 1;
    34: op1_05_inv12 = 1;
    42: op1_05_inv12 = 1;
    94: op1_05_inv12 = 1;
    97: op1_05_inv12 = 1;
    99: op1_05_inv12 = 1;
    103: op1_05_inv12 = 1;
    104: op1_05_inv12 = 1;
    105: op1_05_inv12 = 1;
    108: op1_05_inv12 = 1;
    110: op1_05_inv12 = 1;
    111: op1_05_inv12 = 1;
    112: op1_05_inv12 = 1;
    114: op1_05_inv12 = 1;
    118: op1_05_inv12 = 1;
    120: op1_05_inv12 = 1;
    122: op1_05_inv12 = 1;
    123: op1_05_inv12 = 1;
    125: op1_05_inv12 = 1;
    126: op1_05_inv12 = 1;
    127: op1_05_inv12 = 1;
    130: op1_05_inv12 = 1;
    default: op1_05_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in13 = reg_0754;
    55: op1_05_in13 = reg_0623;
    53: op1_05_in13 = reg_0011;
    86: op1_05_in13 = reg_0673;
    69: op1_05_in13 = reg_0608;
    56: op1_05_in13 = reg_0608;
    73: op1_05_in13 = reg_0115;
    61: op1_05_in13 = reg_0027;
    50: op1_05_in13 = imem07_in[15:12];
    71: op1_05_in13 = reg_0389;
    54: op1_05_in13 = reg_0446;
    68: op1_05_in13 = reg_0790;
    74: op1_05_in13 = reg_0272;
    75: op1_05_in13 = reg_0864;
    87: op1_05_in13 = reg_0208;
    76: op1_05_in13 = reg_1181;
    60: op1_05_in13 = reg_0304;
    46: op1_05_in13 = reg_0833;
    57: op1_05_in13 = imem07_in[7:4];
    77: op1_05_in13 = reg_0881;
    119: op1_05_in13 = reg_0881;
    48: op1_05_in13 = reg_0996;
    70: op1_05_in13 = reg_0280;
    58: op1_05_in13 = reg_0411;
    78: op1_05_in13 = reg_1064;
    88: op1_05_in13 = reg_0252;
    51: op1_05_in13 = reg_0981;
    79: op1_05_in13 = reg_0072;
    125: op1_05_in13 = reg_0072;
    59: op1_05_in13 = reg_0664;
    80: op1_05_in13 = reg_1258;
    121: op1_05_in13 = reg_1258;
    62: op1_05_in13 = reg_0166;
    52: op1_05_in13 = reg_1093;
    37: op1_05_in13 = reg_0123;
    81: op1_05_in13 = reg_0609;
    63: op1_05_in13 = reg_0128;
    82: op1_05_in13 = reg_0298;
    89: op1_05_in13 = reg_1040;
    83: op1_05_in13 = reg_1230;
    84: op1_05_in13 = reg_0155;
    47: op1_05_in13 = reg_0140;
    65: op1_05_in13 = reg_0552;
    85: op1_05_in13 = reg_1348;
    90: op1_05_in13 = reg_0796;
    66: op1_05_in13 = reg_0889;
    44: op1_05_in13 = reg_0393;
    91: op1_05_in13 = reg_0066;
    67: op1_05_in13 = reg_0570;
    92: op1_05_in13 = reg_0611;
    93: op1_05_in13 = reg_0443;
    42: op1_05_in13 = reg_0161;
    94: op1_05_in13 = reg_0105;
    95: op1_05_in13 = reg_0124;
    115: op1_05_in13 = reg_0124;
    96: op1_05_in13 = reg_0127;
    97: op1_05_in13 = reg_0802;
    99: op1_05_in13 = reg_0296;
    100: op1_05_in13 = reg_0886;
    101: op1_05_in13 = reg_0188;
    102: op1_05_in13 = reg_0531;
    123: op1_05_in13 = reg_0531;
    103: op1_05_in13 = reg_0562;
    104: op1_05_in13 = reg_0103;
    105: op1_05_in13 = reg_0800;
    106: op1_05_in13 = reg_0845;
    107: op1_05_in13 = reg_0050;
    108: op1_05_in13 = reg_0564;
    109: op1_05_in13 = reg_0574;
    110: op1_05_in13 = reg_0871;
    111: op1_05_in13 = imem06_in[11:8];
    112: op1_05_in13 = reg_0409;
    113: op1_05_in13 = reg_1268;
    38: op1_05_in13 = reg_0084;
    114: op1_05_in13 = reg_0957;
    116: op1_05_in13 = reg_0927;
    117: op1_05_in13 = reg_0156;
    118: op1_05_in13 = reg_0387;
    120: op1_05_in13 = reg_0497;
    122: op1_05_in13 = reg_0315;
    124: op1_05_in13 = reg_0573;
    126: op1_05_in13 = reg_1009;
    127: op1_05_in13 = reg_1321;
    128: op1_05_in13 = reg_0089;
    129: op1_05_in13 = reg_0870;
    130: op1_05_in13 = reg_0215;
    131: op1_05_in13 = reg_1041;
    default: op1_05_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_05_inv13 = 1;
    86: op1_05_inv13 = 1;
    69: op1_05_inv13 = 1;
    73: op1_05_inv13 = 1;
    61: op1_05_inv13 = 1;
    50: op1_05_inv13 = 1;
    71: op1_05_inv13 = 1;
    54: op1_05_inv13 = 1;
    68: op1_05_inv13 = 1;
    74: op1_05_inv13 = 1;
    75: op1_05_inv13 = 1;
    56: op1_05_inv13 = 1;
    87: op1_05_inv13 = 1;
    76: op1_05_inv13 = 1;
    60: op1_05_inv13 = 1;
    57: op1_05_inv13 = 1;
    77: op1_05_inv13 = 1;
    48: op1_05_inv13 = 1;
    70: op1_05_inv13 = 1;
    78: op1_05_inv13 = 1;
    88: op1_05_inv13 = 1;
    51: op1_05_inv13 = 1;
    79: op1_05_inv13 = 1;
    80: op1_05_inv13 = 1;
    52: op1_05_inv13 = 1;
    63: op1_05_inv13 = 1;
    89: op1_05_inv13 = 1;
    65: op1_05_inv13 = 1;
    92: op1_05_inv13 = 1;
    93: op1_05_inv13 = 1;
    96: op1_05_inv13 = 1;
    97: op1_05_inv13 = 1;
    100: op1_05_inv13 = 1;
    105: op1_05_inv13 = 1;
    106: op1_05_inv13 = 1;
    109: op1_05_inv13 = 1;
    110: op1_05_inv13 = 1;
    111: op1_05_inv13 = 1;
    119: op1_05_inv13 = 1;
    120: op1_05_inv13 = 1;
    123: op1_05_inv13 = 1;
    125: op1_05_inv13 = 1;
    126: op1_05_inv13 = 1;
    127: op1_05_inv13 = 1;
    129: op1_05_inv13 = 1;
    default: op1_05_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in14 = reg_0751;
    55: op1_05_in14 = reg_0321;
    53: op1_05_in14 = reg_0222;
    86: op1_05_in14 = reg_1325;
    69: op1_05_in14 = reg_1344;
    73: op1_05_in14 = reg_0110;
    61: op1_05_in14 = imem01_in[3:0];
    50: op1_05_in14 = reg_0226;
    71: op1_05_in14 = reg_0917;
    116: op1_05_in14 = reg_0917;
    54: op1_05_in14 = reg_0254;
    68: op1_05_in14 = reg_0425;
    74: op1_05_in14 = reg_0697;
    75: op1_05_in14 = reg_0151;
    56: op1_05_in14 = reg_0588;
    87: op1_05_in14 = reg_1368;
    76: op1_05_in14 = reg_1404;
    60: op1_05_in14 = reg_0338;
    46: op1_05_in14 = reg_0702;
    57: op1_05_in14 = imem07_in[15:12];
    77: op1_05_in14 = reg_0886;
    48: op1_05_in14 = reg_0565;
    70: op1_05_in14 = reg_0732;
    58: op1_05_in14 = reg_0595;
    78: op1_05_in14 = reg_0192;
    88: op1_05_in14 = reg_0531;
    51: op1_05_in14 = reg_0973;
    79: op1_05_in14 = reg_0057;
    59: op1_05_in14 = reg_0366;
    80: op1_05_in14 = reg_0462;
    62: op1_05_in14 = reg_1290;
    52: op1_05_in14 = reg_1091;
    81: op1_05_in14 = reg_0715;
    63: op1_05_in14 = reg_0111;
    82: op1_05_in14 = reg_0894;
    89: op1_05_in14 = reg_0451;
    83: op1_05_in14 = reg_1229;
    84: op1_05_in14 = reg_0202;
    47: op1_05_in14 = reg_0779;
    65: op1_05_in14 = reg_0464;
    85: op1_05_in14 = reg_0828;
    90: op1_05_in14 = reg_1077;
    66: op1_05_in14 = reg_0475;
    44: op1_05_in14 = reg_0736;
    91: op1_05_in14 = reg_0604;
    67: op1_05_in14 = reg_0345;
    92: op1_05_in14 = reg_1253;
    93: op1_05_in14 = imem04_in[3:0];
    42: op1_05_in14 = reg_0162;
    94: op1_05_in14 = reg_0629;
    95: op1_05_in14 = reg_1182;
    115: op1_05_in14 = reg_1182;
    96: op1_05_in14 = reg_0382;
    97: op1_05_in14 = reg_0695;
    99: op1_05_in14 = reg_0419;
    100: op1_05_in14 = reg_0352;
    101: op1_05_in14 = reg_0201;
    102: op1_05_in14 = reg_0796;
    103: op1_05_in14 = reg_0173;
    104: op1_05_in14 = reg_0004;
    105: op1_05_in14 = reg_0294;
    106: op1_05_in14 = reg_0608;
    107: op1_05_in14 = reg_0003;
    108: op1_05_in14 = reg_0300;
    109: op1_05_in14 = reg_1215;
    110: op1_05_in14 = reg_0902;
    111: op1_05_in14 = reg_1064;
    112: op1_05_in14 = reg_0134;
    113: op1_05_in14 = reg_0176;
    38: op1_05_in14 = reg_0521;
    114: op1_05_in14 = reg_0952;
    117: op1_05_in14 = reg_0489;
    118: op1_05_in14 = reg_0723;
    119: op1_05_in14 = reg_0405;
    120: op1_05_in14 = reg_0898;
    121: op1_05_in14 = reg_0297;
    122: op1_05_in14 = reg_0735;
    123: op1_05_in14 = reg_1200;
    124: op1_05_in14 = reg_0597;
    125: op1_05_in14 = reg_0005;
    126: op1_05_in14 = reg_1145;
    127: op1_05_in14 = reg_1324;
    128: op1_05_in14 = reg_0386;
    129: op1_05_in14 = reg_0960;
    130: op1_05_in14 = reg_0214;
    131: op1_05_in14 = reg_1040;
    default: op1_05_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv14 = 1;
    55: op1_05_inv14 = 1;
    53: op1_05_inv14 = 1;
    86: op1_05_inv14 = 1;
    69: op1_05_inv14 = 1;
    73: op1_05_inv14 = 1;
    61: op1_05_inv14 = 1;
    50: op1_05_inv14 = 1;
    54: op1_05_inv14 = 1;
    68: op1_05_inv14 = 1;
    75: op1_05_inv14 = 1;
    56: op1_05_inv14 = 1;
    46: op1_05_inv14 = 1;
    77: op1_05_inv14 = 1;
    70: op1_05_inv14 = 1;
    51: op1_05_inv14 = 1;
    59: op1_05_inv14 = 1;
    80: op1_05_inv14 = 1;
    52: op1_05_inv14 = 1;
    82: op1_05_inv14 = 1;
    83: op1_05_inv14 = 1;
    85: op1_05_inv14 = 1;
    94: op1_05_inv14 = 1;
    97: op1_05_inv14 = 1;
    100: op1_05_inv14 = 1;
    101: op1_05_inv14 = 1;
    103: op1_05_inv14 = 1;
    107: op1_05_inv14 = 1;
    111: op1_05_inv14 = 1;
    114: op1_05_inv14 = 1;
    117: op1_05_inv14 = 1;
    119: op1_05_inv14 = 1;
    120: op1_05_inv14 = 1;
    123: op1_05_inv14 = 1;
    125: op1_05_inv14 = 1;
    128: op1_05_inv14 = 1;
    129: op1_05_inv14 = 1;
    130: op1_05_inv14 = 1;
    default: op1_05_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in15 = imem06_in[15:12];
    53: op1_05_in15 = reg_0666;
    86: op1_05_in15 = reg_1280;
    69: op1_05_in15 = reg_1260;
    73: op1_05_in15 = reg_0109;
    61: op1_05_in15 = imem01_in[11:8];
    125: op1_05_in15 = imem01_in[11:8];
    50: op1_05_in15 = reg_0892;
    71: op1_05_in15 = reg_0822;
    54: op1_05_in15 = reg_0629;
    68: op1_05_in15 = reg_0208;
    74: op1_05_in15 = reg_1404;
    75: op1_05_in15 = reg_1105;
    56: op1_05_in15 = reg_0590;
    87: op1_05_in15 = reg_1367;
    76: op1_05_in15 = reg_0541;
    60: op1_05_in15 = reg_0236;
    46: op1_05_in15 = reg_0646;
    57: op1_05_in15 = reg_0600;
    77: op1_05_in15 = reg_0188;
    84: op1_05_in15 = reg_0188;
    100: op1_05_in15 = reg_0188;
    48: op1_05_in15 = reg_0066;
    70: op1_05_in15 = reg_0191;
    58: op1_05_in15 = reg_0268;
    78: op1_05_in15 = reg_1209;
    88: op1_05_in15 = reg_0297;
    51: op1_05_in15 = reg_0125;
    79: op1_05_in15 = reg_1322;
    59: op1_05_in15 = reg_0442;
    80: op1_05_in15 = reg_1082;
    62: op1_05_in15 = reg_1070;
    52: op1_05_in15 = reg_0709;
    81: op1_05_in15 = reg_0968;
    63: op1_05_in15 = reg_0106;
    82: op1_05_in15 = reg_0135;
    89: op1_05_in15 = reg_0033;
    83: op1_05_in15 = reg_0460;
    47: op1_05_in15 = reg_0775;
    65: op1_05_in15 = reg_0451;
    85: op1_05_in15 = reg_0458;
    90: op1_05_in15 = reg_0698;
    66: op1_05_in15 = reg_0474;
    44: op1_05_in15 = reg_0345;
    91: op1_05_in15 = reg_0391;
    67: op1_05_in15 = reg_0132;
    92: op1_05_in15 = reg_0277;
    93: op1_05_in15 = imem04_in[7:4];
    42: op1_05_in15 = reg_0365;
    94: op1_05_in15 = reg_0496;
    96: op1_05_in15 = reg_0876;
    97: op1_05_in15 = reg_0009;
    99: op1_05_in15 = reg_0244;
    101: op1_05_in15 = reg_0410;
    102: op1_05_in15 = reg_0412;
    103: op1_05_in15 = reg_0182;
    104: op1_05_in15 = reg_0003;
    105: op1_05_in15 = reg_1078;
    106: op1_05_in15 = reg_0839;
    107: op1_05_in15 = reg_0001;
    108: op1_05_in15 = reg_0492;
    109: op1_05_in15 = reg_0407;
    110: op1_05_in15 = reg_0463;
    111: op1_05_in15 = reg_1334;
    112: op1_05_in15 = reg_0388;
    113: op1_05_in15 = reg_0992;
    114: op1_05_in15 = reg_1092;
    116: op1_05_in15 = reg_1100;
    118: op1_05_in15 = reg_1100;
    117: op1_05_in15 = reg_0224;
    119: op1_05_in15 = reg_0060;
    120: op1_05_in15 = reg_0472;
    121: op1_05_in15 = reg_1083;
    122: op1_05_in15 = reg_1168;
    123: op1_05_in15 = reg_0969;
    124: op1_05_in15 = reg_0261;
    126: op1_05_in15 = reg_0154;
    127: op1_05_in15 = reg_0026;
    128: op1_05_in15 = reg_0547;
    129: op1_05_in15 = reg_0696;
    130: op1_05_in15 = reg_0022;
    131: op1_05_in15 = reg_0452;
    default: op1_05_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv15 = 1;
    86: op1_05_inv15 = 1;
    68: op1_05_inv15 = 1;
    74: op1_05_inv15 = 1;
    75: op1_05_inv15 = 1;
    76: op1_05_inv15 = 1;
    46: op1_05_inv15 = 1;
    57: op1_05_inv15 = 1;
    77: op1_05_inv15 = 1;
    70: op1_05_inv15 = 1;
    58: op1_05_inv15 = 1;
    78: op1_05_inv15 = 1;
    88: op1_05_inv15 = 1;
    51: op1_05_inv15 = 1;
    79: op1_05_inv15 = 1;
    59: op1_05_inv15 = 1;
    52: op1_05_inv15 = 1;
    81: op1_05_inv15 = 1;
    89: op1_05_inv15 = 1;
    83: op1_05_inv15 = 1;
    47: op1_05_inv15 = 1;
    85: op1_05_inv15 = 1;
    90: op1_05_inv15 = 1;
    91: op1_05_inv15 = 1;
    92: op1_05_inv15 = 1;
    42: op1_05_inv15 = 1;
    96: op1_05_inv15 = 1;
    99: op1_05_inv15 = 1;
    100: op1_05_inv15 = 1;
    102: op1_05_inv15 = 1;
    105: op1_05_inv15 = 1;
    106: op1_05_inv15 = 1;
    108: op1_05_inv15 = 1;
    110: op1_05_inv15 = 1;
    111: op1_05_inv15 = 1;
    112: op1_05_inv15 = 1;
    113: op1_05_inv15 = 1;
    117: op1_05_inv15 = 1;
    119: op1_05_inv15 = 1;
    123: op1_05_inv15 = 1;
    125: op1_05_inv15 = 1;
    129: op1_05_inv15 = 1;
    130: op1_05_inv15 = 1;
    131: op1_05_inv15 = 1;
    default: op1_05_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in16 = reg_1436;
    53: op1_05_in16 = reg_0820;
    86: op1_05_in16 = reg_0443;
    69: op1_05_in16 = reg_0332;
    73: op1_05_in16 = reg_0374;
    129: op1_05_in16 = reg_0374;
    61: op1_05_in16 = reg_1290;
    50: op1_05_in16 = reg_0851;
    71: op1_05_in16 = reg_0335;
    54: op1_05_in16 = reg_0590;
    68: op1_05_in16 = reg_0181;
    74: op1_05_in16 = reg_0541;
    75: op1_05_in16 = reg_0780;
    56: op1_05_in16 = reg_0563;
    87: op1_05_in16 = reg_0088;
    76: op1_05_in16 = imem05_in[11:8];
    60: op1_05_in16 = reg_0237;
    46: op1_05_in16 = reg_0602;
    57: op1_05_in16 = reg_0667;
    77: op1_05_in16 = reg_0435;
    48: op1_05_in16 = reg_0045;
    103: op1_05_in16 = reg_0045;
    70: op1_05_in16 = reg_0216;
    58: op1_05_in16 = imem04_in[15:12];
    93: op1_05_in16 = imem04_in[15:12];
    78: op1_05_in16 = reg_0974;
    88: op1_05_in16 = reg_1083;
    51: op1_05_in16 = reg_0105;
    79: op1_05_in16 = reg_0122;
    59: op1_05_in16 = reg_0741;
    80: op1_05_in16 = reg_0464;
    62: op1_05_in16 = reg_0549;
    52: op1_05_in16 = reg_0235;
    81: op1_05_in16 = reg_0146;
    63: op1_05_in16 = reg_0382;
    82: op1_05_in16 = reg_1345;
    89: op1_05_in16 = reg_0487;
    83: op1_05_in16 = reg_1405;
    84: op1_05_in16 = reg_0201;
    47: op1_05_in16 = reg_0031;
    65: op1_05_in16 = reg_0320;
    85: op1_05_in16 = reg_0133;
    90: op1_05_in16 = reg_0262;
    66: op1_05_in16 = reg_0934;
    44: op1_05_in16 = reg_0700;
    91: op1_05_in16 = reg_0303;
    67: op1_05_in16 = reg_0119;
    92: op1_05_in16 = reg_0754;
    42: op1_05_in16 = reg_0363;
    94: op1_05_in16 = reg_0560;
    96: op1_05_in16 = reg_0473;
    97: op1_05_in16 = imem03_in[3:0];
    99: op1_05_in16 = reg_0977;
    100: op1_05_in16 = reg_0388;
    101: op1_05_in16 = reg_0405;
    102: op1_05_in16 = reg_0407;
    104: op1_05_in16 = reg_0001;
    105: op1_05_in16 = reg_0068;
    106: op1_05_in16 = reg_0744;
    107: op1_05_in16 = reg_0123;
    108: op1_05_in16 = reg_1373;
    109: op1_05_in16 = reg_0061;
    110: op1_05_in16 = reg_0163;
    111: op1_05_in16 = reg_0751;
    112: op1_05_in16 = reg_0071;
    113: op1_05_in16 = reg_0562;
    114: op1_05_in16 = reg_0108;
    116: op1_05_in16 = reg_0282;
    118: op1_05_in16 = reg_0282;
    117: op1_05_in16 = reg_0775;
    119: op1_05_in16 = reg_1321;
    120: op1_05_in16 = reg_0433;
    121: op1_05_in16 = reg_0412;
    122: op1_05_in16 = reg_0445;
    123: op1_05_in16 = reg_1077;
    124: op1_05_in16 = reg_0557;
    125: op1_05_in16 = reg_0120;
    126: op1_05_in16 = reg_0444;
    127: op1_05_in16 = reg_0917;
    128: op1_05_in16 = reg_0372;
    130: op1_05_in16 = reg_1170;
    131: op1_05_in16 = reg_0062;
    default: op1_05_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_05_inv16 = 1;
    69: op1_05_inv16 = 1;
    73: op1_05_inv16 = 1;
    61: op1_05_inv16 = 1;
    68: op1_05_inv16 = 1;
    76: op1_05_inv16 = 1;
    46: op1_05_inv16 = 1;
    57: op1_05_inv16 = 1;
    48: op1_05_inv16 = 1;
    79: op1_05_inv16 = 1;
    59: op1_05_inv16 = 1;
    62: op1_05_inv16 = 1;
    83: op1_05_inv16 = 1;
    84: op1_05_inv16 = 1;
    47: op1_05_inv16 = 1;
    90: op1_05_inv16 = 1;
    44: op1_05_inv16 = 1;
    91: op1_05_inv16 = 1;
    67: op1_05_inv16 = 1;
    93: op1_05_inv16 = 1;
    42: op1_05_inv16 = 1;
    101: op1_05_inv16 = 1;
    103: op1_05_inv16 = 1;
    108: op1_05_inv16 = 1;
    112: op1_05_inv16 = 1;
    114: op1_05_inv16 = 1;
    116: op1_05_inv16 = 1;
    119: op1_05_inv16 = 1;
    121: op1_05_inv16 = 1;
    122: op1_05_inv16 = 1;
    130: op1_05_inv16 = 1;
    131: op1_05_inv16 = 1;
    default: op1_05_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in17 = reg_0905;
    53: op1_05_in17 = reg_0632;
    86: op1_05_in17 = reg_0411;
    69: op1_05_in17 = reg_0475;
    73: op1_05_in17 = reg_1225;
    61: op1_05_in17 = reg_1254;
    50: op1_05_in17 = reg_0159;
    71: op1_05_in17 = reg_1253;
    54: op1_05_in17 = reg_0589;
    68: op1_05_in17 = reg_1338;
    74: op1_05_in17 = imem05_in[3:0];
    75: op1_05_in17 = reg_0261;
    56: op1_05_in17 = reg_0530;
    87: op1_05_in17 = reg_0264;
    76: op1_05_in17 = imem05_in[15:12];
    60: op1_05_in17 = reg_0181;
    46: op1_05_in17 = reg_0567;
    57: op1_05_in17 = reg_0223;
    82: op1_05_in17 = reg_0223;
    77: op1_05_in17 = reg_0409;
    48: op1_05_in17 = reg_0315;
    70: op1_05_in17 = imem03_in[7:4];
    58: op1_05_in17 = reg_1258;
    78: op1_05_in17 = reg_1420;
    88: op1_05_in17 = reg_1203;
    51: op1_05_in17 = reg_0138;
    79: op1_05_in17 = reg_1068;
    59: op1_05_in17 = reg_0114;
    80: op1_05_in17 = reg_1147;
    62: op1_05_in17 = reg_0550;
    52: op1_05_in17 = reg_1064;
    81: op1_05_in17 = reg_0383;
    63: op1_05_in17 = reg_0306;
    89: op1_05_in17 = reg_0837;
    90: op1_05_in17 = reg_0837;
    83: op1_05_in17 = reg_0928;
    84: op1_05_in17 = reg_0431;
    47: op1_05_in17 = reg_0664;
    65: op1_05_in17 = reg_0342;
    85: op1_05_in17 = imem06_in[11:8];
    66: op1_05_in17 = reg_0382;
    44: op1_05_in17 = reg_0701;
    91: op1_05_in17 = reg_0873;
    67: op1_05_in17 = reg_0270;
    92: op1_05_in17 = reg_0093;
    93: op1_05_in17 = reg_0032;
    42: op1_05_in17 = reg_0183;
    128: op1_05_in17 = reg_0183;
    94: op1_05_in17 = reg_1392;
    96: op1_05_in17 = reg_0829;
    97: op1_05_in17 = reg_0505;
    99: op1_05_in17 = reg_0023;
    100: op1_05_in17 = reg_0060;
    101: op1_05_in17 = reg_0060;
    102: op1_05_in17 = reg_0199;
    103: op1_05_in17 = reg_0564;
    104: op1_05_in17 = reg_0521;
    105: op1_05_in17 = reg_0168;
    106: op1_05_in17 = reg_0532;
    107: op1_05_in17 = reg_0124;
    108: op1_05_in17 = reg_0864;
    109: op1_05_in17 = reg_0862;
    110: op1_05_in17 = reg_0747;
    111: op1_05_in17 = reg_0860;
    112: op1_05_in17 = reg_0072;
    113: op1_05_in17 = reg_0630;
    114: op1_05_in17 = reg_0882;
    116: op1_05_in17 = reg_0871;
    127: op1_05_in17 = reg_0871;
    117: op1_05_in17 = reg_0774;
    118: op1_05_in17 = reg_0734;
    119: op1_05_in17 = reg_0057;
    120: op1_05_in17 = reg_0776;
    121: op1_05_in17 = reg_0471;
    122: op1_05_in17 = reg_0251;
    123: op1_05_in17 = reg_0454;
    124: op1_05_in17 = reg_0783;
    125: op1_05_in17 = reg_0874;
    126: op1_05_in17 = reg_0709;
    129: op1_05_in17 = reg_0585;
    130: op1_05_in17 = reg_0087;
    131: op1_05_in17 = reg_0487;
    default: op1_05_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv17 = 1;
    53: op1_05_inv17 = 1;
    86: op1_05_inv17 = 1;
    50: op1_05_inv17 = 1;
    71: op1_05_inv17 = 1;
    74: op1_05_inv17 = 1;
    56: op1_05_inv17 = 1;
    60: op1_05_inv17 = 1;
    57: op1_05_inv17 = 1;
    77: op1_05_inv17 = 1;
    48: op1_05_inv17 = 1;
    70: op1_05_inv17 = 1;
    78: op1_05_inv17 = 1;
    88: op1_05_inv17 = 1;
    51: op1_05_inv17 = 1;
    79: op1_05_inv17 = 1;
    80: op1_05_inv17 = 1;
    62: op1_05_inv17 = 1;
    81: op1_05_inv17 = 1;
    63: op1_05_inv17 = 1;
    82: op1_05_inv17 = 1;
    89: op1_05_inv17 = 1;
    47: op1_05_inv17 = 1;
    65: op1_05_inv17 = 1;
    85: op1_05_inv17 = 1;
    91: op1_05_inv17 = 1;
    92: op1_05_inv17 = 1;
    42: op1_05_inv17 = 1;
    96: op1_05_inv17 = 1;
    97: op1_05_inv17 = 1;
    101: op1_05_inv17 = 1;
    104: op1_05_inv17 = 1;
    106: op1_05_inv17 = 1;
    109: op1_05_inv17 = 1;
    112: op1_05_inv17 = 1;
    117: op1_05_inv17 = 1;
    118: op1_05_inv17 = 1;
    120: op1_05_inv17 = 1;
    124: op1_05_inv17 = 1;
    125: op1_05_inv17 = 1;
    128: op1_05_inv17 = 1;
    129: op1_05_inv17 = 1;
    130: op1_05_inv17 = 1;
    default: op1_05_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in18 = reg_0870;
    53: op1_05_in18 = reg_0629;
    86: op1_05_in18 = reg_0493;
    69: op1_05_in18 = reg_0436;
    73: op1_05_in18 = reg_0323;
    61: op1_05_in18 = reg_1032;
    50: op1_05_in18 = reg_0923;
    71: op1_05_in18 = reg_0728;
    54: op1_05_in18 = reg_0561;
    68: op1_05_in18 = reg_1083;
    74: op1_05_in18 = reg_0318;
    48: op1_05_in18 = reg_0318;
    75: op1_05_in18 = reg_0466;
    56: op1_05_in18 = reg_0531;
    87: op1_05_in18 = reg_0034;
    76: op1_05_in18 = reg_0477;
    60: op1_05_in18 = reg_0129;
    46: op1_05_in18 = reg_0565;
    57: op1_05_in18 = reg_0892;
    77: op1_05_in18 = reg_0071;
    70: op1_05_in18 = reg_1149;
    58: op1_05_in18 = reg_0462;
    78: op1_05_in18 = reg_0133;
    88: op1_05_in18 = reg_1198;
    51: op1_05_in18 = reg_0708;
    79: op1_05_in18 = reg_1256;
    59: op1_05_in18 = reg_0520;
    80: op1_05_in18 = reg_0796;
    62: op1_05_in18 = reg_0468;
    52: op1_05_in18 = reg_0375;
    81: op1_05_in18 = reg_0092;
    63: op1_05_in18 = reg_0848;
    82: op1_05_in18 = reg_0663;
    89: op1_05_in18 = reg_1151;
    83: op1_05_in18 = reg_0883;
    84: op1_05_in18 = reg_0416;
    47: op1_05_in18 = reg_0285;
    65: op1_05_in18 = reg_0470;
    85: op1_05_in18 = reg_0860;
    90: op1_05_in18 = reg_0336;
    66: op1_05_in18 = reg_0903;
    44: op1_05_in18 = reg_0523;
    91: op1_05_in18 = reg_0872;
    67: op1_05_in18 = reg_0229;
    92: op1_05_in18 = reg_0331;
    93: op1_05_in18 = reg_1372;
    42: op1_05_in18 = reg_0077;
    94: op1_05_in18 = imem03_in[11:8];
    96: op1_05_in18 = reg_0695;
    97: op1_05_in18 = reg_0999;
    105: op1_05_in18 = reg_0999;
    99: op1_05_in18 = imem07_in[3:0];
    100: op1_05_in18 = reg_0026;
    101: op1_05_in18 = reg_0734;
    102: op1_05_in18 = reg_1004;
    103: op1_05_in18 = reg_0131;
    106: op1_05_in18 = reg_0433;
    108: op1_05_in18 = reg_0449;
    109: op1_05_in18 = reg_0836;
    110: op1_05_in18 = reg_0222;
    111: op1_05_in18 = reg_0863;
    112: op1_05_in18 = reg_0059;
    113: op1_05_in18 = reg_1181;
    114: op1_05_in18 = reg_0448;
    116: op1_05_in18 = reg_0401;
    117: op1_05_in18 = reg_0441;
    118: op1_05_in18 = reg_0463;
    119: op1_05_in18 = reg_0122;
    120: op1_05_in18 = reg_1450;
    121: op1_05_in18 = reg_1077;
    122: op1_05_in18 = reg_0066;
    123: op1_05_in18 = reg_0061;
    124: op1_05_in18 = reg_0145;
    125: op1_05_in18 = reg_0930;
    126: op1_05_in18 = reg_0965;
    127: op1_05_in18 = reg_0550;
    128: op1_05_in18 = reg_0902;
    129: op1_05_in18 = reg_0624;
    130: op1_05_in18 = reg_1060;
    131: op1_05_in18 = reg_0719;
    default: op1_05_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv18 = 1;
    53: op1_05_inv18 = 1;
    86: op1_05_inv18 = 1;
    69: op1_05_inv18 = 1;
    50: op1_05_inv18 = 1;
    87: op1_05_inv18 = 1;
    60: op1_05_inv18 = 1;
    46: op1_05_inv18 = 1;
    48: op1_05_inv18 = 1;
    88: op1_05_inv18 = 1;
    51: op1_05_inv18 = 1;
    59: op1_05_inv18 = 1;
    80: op1_05_inv18 = 1;
    52: op1_05_inv18 = 1;
    63: op1_05_inv18 = 1;
    83: op1_05_inv18 = 1;
    85: op1_05_inv18 = 1;
    44: op1_05_inv18 = 1;
    92: op1_05_inv18 = 1;
    96: op1_05_inv18 = 1;
    97: op1_05_inv18 = 1;
    99: op1_05_inv18 = 1;
    100: op1_05_inv18 = 1;
    103: op1_05_inv18 = 1;
    108: op1_05_inv18 = 1;
    109: op1_05_inv18 = 1;
    117: op1_05_inv18 = 1;
    119: op1_05_inv18 = 1;
    123: op1_05_inv18 = 1;
    124: op1_05_inv18 = 1;
    125: op1_05_inv18 = 1;
    126: op1_05_inv18 = 1;
    default: op1_05_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in19 = reg_1323;
    111: op1_05_in19 = reg_1323;
    53: op1_05_in19 = reg_0607;
    86: op1_05_in19 = imem04_in[7:4];
    69: op1_05_in19 = reg_0128;
    73: op1_05_in19 = reg_0371;
    61: op1_05_in19 = reg_0372;
    50: op1_05_in19 = reg_0029;
    71: op1_05_in19 = reg_1031;
    54: op1_05_in19 = reg_1140;
    68: op1_05_in19 = reg_1147;
    74: op1_05_in19 = reg_1485;
    75: op1_05_in19 = reg_0316;
    56: op1_05_in19 = reg_0256;
    87: op1_05_in19 = reg_0252;
    76: op1_05_in19 = reg_1514;
    60: op1_05_in19 = reg_0063;
    46: op1_05_in19 = reg_0183;
    57: op1_05_in19 = reg_0893;
    77: op1_05_in19 = reg_0060;
    48: op1_05_in19 = reg_0938;
    70: op1_05_in19 = reg_0376;
    58: op1_05_in19 = reg_1215;
    88: op1_05_in19 = reg_1215;
    78: op1_05_in19 = reg_0860;
    51: op1_05_in19 = reg_0711;
    79: op1_05_in19 = reg_0277;
    59: op1_05_in19 = reg_0124;
    80: op1_05_in19 = reg_0033;
    62: op1_05_in19 = reg_0430;
    52: op1_05_in19 = reg_1003;
    81: op1_05_in19 = reg_0257;
    63: op1_05_in19 = reg_0008;
    96: op1_05_in19 = reg_0008;
    82: op1_05_in19 = reg_0664;
    89: op1_05_in19 = reg_1189;
    83: op1_05_in19 = reg_0886;
    84: op1_05_in19 = reg_0388;
    47: op1_05_in19 = reg_0741;
    65: op1_05_in19 = reg_0488;
    85: op1_05_in19 = reg_0720;
    90: op1_05_in19 = reg_0932;
    66: op1_05_in19 = reg_0876;
    44: op1_05_in19 = reg_0445;
    91: op1_05_in19 = reg_0575;
    67: op1_05_in19 = reg_0185;
    92: op1_05_in19 = reg_0260;
    93: op1_05_in19 = reg_0264;
    42: op1_05_in19 = reg_0044;
    94: op1_05_in19 = reg_0121;
    97: op1_05_in19 = reg_0573;
    99: op1_05_in19 = imem07_in[11:8];
    100: op1_05_in19 = reg_0267;
    101: op1_05_in19 = imem01_in[3:0];
    102: op1_05_in19 = reg_0452;
    103: op1_05_in19 = imem05_in[3:0];
    105: op1_05_in19 = reg_1448;
    106: op1_05_in19 = reg_0429;
    108: op1_05_in19 = reg_0828;
    109: op1_05_in19 = reg_1151;
    110: op1_05_in19 = reg_0241;
    118: op1_05_in19 = reg_0241;
    112: op1_05_in19 = reg_1322;
    113: op1_05_in19 = reg_1070;
    114: op1_05_in19 = reg_0707;
    116: op1_05_in19 = reg_0787;
    117: op1_05_in19 = reg_0739;
    119: op1_05_in19 = reg_1512;
    120: op1_05_in19 = reg_1455;
    121: op1_05_in19 = reg_1065;
    122: op1_05_in19 = reg_0562;
    123: op1_05_in19 = reg_0862;
    124: op1_05_in19 = reg_1314;
    125: op1_05_in19 = reg_0547;
    126: op1_05_in19 = reg_0954;
    127: op1_05_in19 = reg_0548;
    128: op1_05_in19 = reg_1255;
    129: op1_05_in19 = reg_0132;
    130: op1_05_in19 = reg_0231;
    131: op1_05_in19 = reg_0594;
    default: op1_05_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv19 = 1;
    53: op1_05_inv19 = 1;
    86: op1_05_inv19 = 1;
    61: op1_05_inv19 = 1;
    50: op1_05_inv19 = 1;
    71: op1_05_inv19 = 1;
    54: op1_05_inv19 = 1;
    74: op1_05_inv19 = 1;
    75: op1_05_inv19 = 1;
    56: op1_05_inv19 = 1;
    87: op1_05_inv19 = 1;
    76: op1_05_inv19 = 1;
    60: op1_05_inv19 = 1;
    77: op1_05_inv19 = 1;
    48: op1_05_inv19 = 1;
    70: op1_05_inv19 = 1;
    78: op1_05_inv19 = 1;
    51: op1_05_inv19 = 1;
    79: op1_05_inv19 = 1;
    80: op1_05_inv19 = 1;
    52: op1_05_inv19 = 1;
    63: op1_05_inv19 = 1;
    89: op1_05_inv19 = 1;
    83: op1_05_inv19 = 1;
    84: op1_05_inv19 = 1;
    65: op1_05_inv19 = 1;
    85: op1_05_inv19 = 1;
    91: op1_05_inv19 = 1;
    67: op1_05_inv19 = 1;
    42: op1_05_inv19 = 1;
    96: op1_05_inv19 = 1;
    101: op1_05_inv19 = 1;
    102: op1_05_inv19 = 1;
    108: op1_05_inv19 = 1;
    109: op1_05_inv19 = 1;
    110: op1_05_inv19 = 1;
    111: op1_05_inv19 = 1;
    112: op1_05_inv19 = 1;
    113: op1_05_inv19 = 1;
    119: op1_05_inv19 = 1;
    122: op1_05_inv19 = 1;
    123: op1_05_inv19 = 1;
    126: op1_05_inv19 = 1;
    127: op1_05_inv19 = 1;
    128: op1_05_inv19 = 1;
    131: op1_05_inv19 = 1;
    default: op1_05_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in20 = reg_0752;
    53: op1_05_in20 = reg_0590;
    86: op1_05_in20 = reg_1338;
    69: op1_05_in20 = reg_0876;
    73: op1_05_in20 = reg_0269;
    61: op1_05_in20 = reg_0634;
    50: op1_05_in20 = reg_0661;
    71: op1_05_in20 = reg_0610;
    54: op1_05_in20 = reg_0474;
    68: op1_05_in20 = reg_0454;
    74: op1_05_in20 = reg_0576;
    119: op1_05_in20 = reg_0576;
    75: op1_05_in20 = reg_0296;
    56: op1_05_in20 = reg_0497;
    87: op1_05_in20 = reg_1215;
    76: op1_05_in20 = reg_0300;
    60: op1_05_in20 = reg_0331;
    46: op1_05_in20 = reg_0301;
    57: op1_05_in20 = reg_0310;
    77: op1_05_in20 = reg_0175;
    48: op1_05_in20 = reg_0418;
    70: op1_05_in20 = reg_0350;
    58: op1_05_in20 = reg_1203;
    78: op1_05_in20 = reg_0859;
    88: op1_05_in20 = reg_0681;
    51: op1_05_in20 = reg_0008;
    79: op1_05_in20 = reg_1512;
    80: op1_05_in20 = reg_0340;
    62: op1_05_in20 = reg_0727;
    81: op1_05_in20 = reg_0727;
    52: op1_05_in20 = reg_0218;
    63: op1_05_in20 = reg_0006;
    82: op1_05_in20 = reg_0286;
    89: op1_05_in20 = reg_0209;
    123: op1_05_in20 = reg_0209;
    83: op1_05_in20 = reg_0722;
    84: op1_05_in20 = reg_0073;
    47: op1_05_in20 = reg_0740;
    65: op1_05_in20 = reg_0305;
    85: op1_05_in20 = reg_0780;
    90: op1_05_in20 = reg_0063;
    66: op1_05_in20 = reg_0879;
    44: op1_05_in20 = reg_0650;
    91: op1_05_in20 = imem05_in[15:12];
    67: op1_05_in20 = reg_0230;
    92: op1_05_in20 = reg_0242;
    93: op1_05_in20 = reg_1258;
    42: op1_05_in20 = reg_0012;
    94: op1_05_in20 = reg_0049;
    96: op1_05_in20 = reg_0227;
    97: op1_05_in20 = reg_0709;
    99: op1_05_in20 = reg_1183;
    100: op1_05_in20 = reg_0723;
    101: op1_05_in20 = reg_0282;
    102: op1_05_in20 = reg_0232;
    103: op1_05_in20 = reg_0303;
    105: op1_05_in20 = reg_0198;
    106: op1_05_in20 = reg_0972;
    108: op1_05_in20 = reg_0317;
    109: op1_05_in20 = reg_1503;
    110: op1_05_in20 = reg_0438;
    111: op1_05_in20 = reg_1179;
    112: op1_05_in20 = reg_0011;
    113: op1_05_in20 = reg_0318;
    114: op1_05_in20 = reg_0025;
    116: op1_05_in20 = reg_0609;
    117: op1_05_in20 = reg_0413;
    118: op1_05_in20 = reg_0430;
    120: op1_05_in20 = reg_0382;
    121: op1_05_in20 = reg_0342;
    122: op1_05_in20 = reg_0173;
    124: op1_05_in20 = reg_0957;
    125: op1_05_in20 = reg_0239;
    126: op1_05_in20 = reg_0962;
    127: op1_05_in20 = reg_0787;
    128: op1_05_in20 = reg_0013;
    129: op1_05_in20 = reg_0308;
    130: op1_05_in20 = reg_0309;
    131: op1_05_in20 = reg_0117;
    default: op1_05_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_05_inv20 = 1;
    86: op1_05_inv20 = 1;
    73: op1_05_inv20 = 1;
    71: op1_05_inv20 = 1;
    74: op1_05_inv20 = 1;
    56: op1_05_inv20 = 1;
    87: op1_05_inv20 = 1;
    76: op1_05_inv20 = 1;
    60: op1_05_inv20 = 1;
    46: op1_05_inv20 = 1;
    77: op1_05_inv20 = 1;
    58: op1_05_inv20 = 1;
    88: op1_05_inv20 = 1;
    80: op1_05_inv20 = 1;
    52: op1_05_inv20 = 1;
    81: op1_05_inv20 = 1;
    63: op1_05_inv20 = 1;
    82: op1_05_inv20 = 1;
    83: op1_05_inv20 = 1;
    84: op1_05_inv20 = 1;
    47: op1_05_inv20 = 1;
    65: op1_05_inv20 = 1;
    85: op1_05_inv20 = 1;
    42: op1_05_inv20 = 1;
    96: op1_05_inv20 = 1;
    97: op1_05_inv20 = 1;
    99: op1_05_inv20 = 1;
    103: op1_05_inv20 = 1;
    105: op1_05_inv20 = 1;
    106: op1_05_inv20 = 1;
    108: op1_05_inv20 = 1;
    109: op1_05_inv20 = 1;
    111: op1_05_inv20 = 1;
    113: op1_05_inv20 = 1;
    114: op1_05_inv20 = 1;
    116: op1_05_inv20 = 1;
    117: op1_05_inv20 = 1;
    121: op1_05_inv20 = 1;
    122: op1_05_inv20 = 1;
    123: op1_05_inv20 = 1;
    125: op1_05_inv20 = 1;
    128: op1_05_inv20 = 1;
    129: op1_05_inv20 = 1;
    130: op1_05_inv20 = 1;
    default: op1_05_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in21 = reg_0264;
    53: op1_05_in21 = reg_0562;
    86: op1_05_in21 = reg_0297;
    69: op1_05_in21 = reg_0381;
    73: op1_05_in21 = reg_0212;
    61: op1_05_in21 = reg_0602;
    103: op1_05_in21 = reg_0602;
    50: op1_05_in21 = reg_0664;
    71: op1_05_in21 = reg_0420;
    54: op1_05_in21 = reg_0433;
    68: op1_05_in21 = reg_0094;
    87: op1_05_in21 = reg_0094;
    74: op1_05_in21 = reg_0197;
    75: op1_05_in21 = reg_0419;
    56: op1_05_in21 = reg_0494;
    76: op1_05_in21 = reg_1484;
    60: op1_05_in21 = imem05_in[7:4];
    46: op1_05_in21 = reg_0090;
    57: op1_05_in21 = reg_0309;
    77: op1_05_in21 = reg_1254;
    48: op1_05_in21 = reg_0300;
    70: op1_05_in21 = reg_0144;
    58: op1_05_in21 = reg_1198;
    78: op1_05_in21 = reg_1323;
    88: op1_05_in21 = reg_1082;
    51: op1_05_in21 = reg_0279;
    79: op1_05_in21 = reg_0550;
    80: op1_05_in21 = reg_0211;
    62: op1_05_in21 = reg_0360;
    52: op1_05_in21 = reg_0557;
    81: op1_05_in21 = reg_0895;
    63: op1_05_in21 = reg_0732;
    82: op1_05_in21 = reg_0741;
    89: op1_05_in21 = reg_0064;
    83: op1_05_in21 = reg_0405;
    84: op1_05_in21 = reg_0059;
    47: op1_05_in21 = reg_0404;
    65: op1_05_in21 = reg_0862;
    85: op1_05_in21 = reg_0116;
    90: op1_05_in21 = reg_0065;
    66: op1_05_in21 = imem02_in[3:0];
    44: op1_05_in21 = reg_0604;
    91: op1_05_in21 = reg_0864;
    67: op1_05_in21 = reg_0378;
    92: op1_05_in21 = reg_0820;
    116: op1_05_in21 = reg_0820;
    93: op1_05_in21 = reg_0531;
    42: op1_05_in21 = reg_0679;
    94: op1_05_in21 = reg_0261;
    96: op1_05_in21 = reg_0168;
    97: op1_05_in21 = reg_0706;
    99: op1_05_in21 = reg_1416;
    100: op1_05_in21 = reg_0871;
    101: op1_05_in21 = reg_1290;
    102: op1_05_in21 = reg_0836;
    105: op1_05_in21 = reg_0783;
    106: op1_05_in21 = reg_1458;
    108: op1_05_in21 = reg_0206;
    109: op1_05_in21 = reg_0470;
    110: op1_05_in21 = reg_0875;
    111: op1_05_in21 = reg_0637;
    112: op1_05_in21 = imem01_in[11:8];
    113: op1_05_in21 = reg_0492;
    114: op1_05_in21 = reg_0291;
    117: op1_05_in21 = reg_0618;
    118: op1_05_in21 = reg_0726;
    119: op1_05_in21 = reg_1474;
    120: op1_05_in21 = reg_0496;
    121: op1_05_in21 = reg_0268;
    122: op1_05_in21 = reg_0701;
    123: op1_05_in21 = reg_0540;
    124: op1_05_in21 = reg_0505;
    125: op1_05_in21 = reg_0830;
    126: op1_05_in21 = reg_0376;
    127: op1_05_in21 = reg_0572;
    128: op1_05_in21 = reg_0258;
    129: op1_05_in21 = reg_0195;
    130: op1_05_in21 = reg_1349;
    131: op1_05_in21 = reg_0210;
    default: op1_05_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_05_inv21 = 1;
    73: op1_05_inv21 = 1;
    61: op1_05_inv21 = 1;
    50: op1_05_inv21 = 1;
    71: op1_05_inv21 = 1;
    74: op1_05_inv21 = 1;
    75: op1_05_inv21 = 1;
    87: op1_05_inv21 = 1;
    76: op1_05_inv21 = 1;
    60: op1_05_inv21 = 1;
    46: op1_05_inv21 = 1;
    77: op1_05_inv21 = 1;
    48: op1_05_inv21 = 1;
    58: op1_05_inv21 = 1;
    79: op1_05_inv21 = 1;
    52: op1_05_inv21 = 1;
    81: op1_05_inv21 = 1;
    82: op1_05_inv21 = 1;
    89: op1_05_inv21 = 1;
    83: op1_05_inv21 = 1;
    65: op1_05_inv21 = 1;
    66: op1_05_inv21 = 1;
    67: op1_05_inv21 = 1;
    94: op1_05_inv21 = 1;
    96: op1_05_inv21 = 1;
    97: op1_05_inv21 = 1;
    99: op1_05_inv21 = 1;
    100: op1_05_inv21 = 1;
    101: op1_05_inv21 = 1;
    103: op1_05_inv21 = 1;
    106: op1_05_inv21 = 1;
    109: op1_05_inv21 = 1;
    110: op1_05_inv21 = 1;
    112: op1_05_inv21 = 1;
    114: op1_05_inv21 = 1;
    116: op1_05_inv21 = 1;
    118: op1_05_inv21 = 1;
    119: op1_05_inv21 = 1;
    124: op1_05_inv21 = 1;
    126: op1_05_inv21 = 1;
    127: op1_05_inv21 = 1;
    128: op1_05_inv21 = 1;
    129: op1_05_inv21 = 1;
    default: op1_05_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in22 = reg_0115;
    53: op1_05_in22 = imem02_in[3:0];
    86: op1_05_in22 = reg_1083;
    69: op1_05_in22 = reg_0024;
    73: op1_05_in22 = reg_0215;
    61: op1_05_in22 = reg_0575;
    50: op1_05_in22 = reg_0284;
    71: op1_05_in22 = imem01_in[7:4];
    54: op1_05_in22 = reg_0972;
    68: op1_05_in22 = reg_0164;
    74: op1_05_in22 = reg_0196;
    75: op1_05_in22 = reg_0165;
    56: op1_05_in22 = reg_0432;
    87: op1_05_in22 = reg_0451;
    76: op1_05_in22 = reg_0130;
    60: op1_05_in22 = reg_0831;
    46: op1_05_in22 = reg_0275;
    57: op1_05_in22 = reg_0489;
    77: op1_05_in22 = reg_1256;
    48: op1_05_in22 = reg_0273;
    70: op1_05_in22 = reg_0559;
    58: op1_05_in22 = reg_1082;
    78: op1_05_in22 = reg_0172;
    88: op1_05_in22 = reg_0599;
    51: op1_05_in22 = reg_0525;
    79: op1_05_in22 = reg_0610;
    80: op1_05_in22 = reg_0065;
    62: op1_05_in22 = reg_0078;
    52: op1_05_in22 = reg_0556;
    81: op1_05_in22 = reg_0874;
    63: op1_05_in22 = reg_0675;
    82: op1_05_in22 = reg_0623;
    89: op1_05_in22 = reg_0021;
    83: op1_05_in22 = reg_0387;
    84: op1_05_in22 = reg_0058;
    47: op1_05_in22 = reg_0592;
    65: op1_05_in22 = reg_0836;
    85: op1_05_in22 = reg_0110;
    90: op1_05_in22 = reg_0095;
    66: op1_05_in22 = reg_0281;
    44: op1_05_in22 = reg_0564;
    91: op1_05_in22 = reg_0828;
    67: op1_05_in22 = reg_0629;
    92: op1_05_in22 = reg_0819;
    93: op1_05_in22 = reg_0471;
    42: op1_05_in22 = reg_0666;
    94: op1_05_in22 = reg_1063;
    96: op1_05_in22 = reg_0507;
    97: op1_05_in22 = reg_0198;
    99: op1_05_in22 = reg_0478;
    100: op1_05_in22 = imem01_in[11:8];
    101: op1_05_in22 = reg_0553;
    102: op1_05_in22 = reg_0835;
    103: op1_05_in22 = reg_0861;
    105: op1_05_in22 = reg_0600;
    106: op1_05_in22 = reg_0380;
    108: op1_05_in22 = reg_0038;
    109: op1_05_in22 = reg_0204;
    110: op1_05_in22 = reg_0402;
    111: op1_05_in22 = reg_0526;
    112: op1_05_in22 = reg_0747;
    113: op1_05_in22 = reg_1348;
    114: op1_05_in22 = reg_1339;
    116: op1_05_in22 = reg_1473;
    125: op1_05_in22 = reg_1473;
    117: op1_05_in22 = reg_0591;
    118: op1_05_in22 = reg_0146;
    119: op1_05_in22 = reg_0726;
    120: op1_05_in22 = reg_0631;
    121: op1_05_in22 = reg_0262;
    122: op1_05_in22 = reg_0566;
    123: op1_05_in22 = imem05_in[7:4];
    124: op1_05_in22 = reg_1199;
    126: op1_05_in22 = reg_0558;
    127: op1_05_in22 = reg_1511;
    128: op1_05_in22 = reg_0548;
    129: op1_05_in22 = reg_0519;
    130: op1_05_in22 = reg_0921;
    131: op1_05_in22 = reg_0832;
    default: op1_05_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv22 = 1;
    53: op1_05_inv22 = 1;
    73: op1_05_inv22 = 1;
    61: op1_05_inv22 = 1;
    50: op1_05_inv22 = 1;
    54: op1_05_inv22 = 1;
    75: op1_05_inv22 = 1;
    56: op1_05_inv22 = 1;
    87: op1_05_inv22 = 1;
    60: op1_05_inv22 = 1;
    57: op1_05_inv22 = 1;
    77: op1_05_inv22 = 1;
    48: op1_05_inv22 = 1;
    70: op1_05_inv22 = 1;
    78: op1_05_inv22 = 1;
    79: op1_05_inv22 = 1;
    80: op1_05_inv22 = 1;
    62: op1_05_inv22 = 1;
    63: op1_05_inv22 = 1;
    84: op1_05_inv22 = 1;
    91: op1_05_inv22 = 1;
    42: op1_05_inv22 = 1;
    94: op1_05_inv22 = 1;
    96: op1_05_inv22 = 1;
    97: op1_05_inv22 = 1;
    99: op1_05_inv22 = 1;
    100: op1_05_inv22 = 1;
    101: op1_05_inv22 = 1;
    103: op1_05_inv22 = 1;
    116: op1_05_inv22 = 1;
    123: op1_05_inv22 = 1;
    124: op1_05_inv22 = 1;
    125: op1_05_inv22 = 1;
    126: op1_05_inv22 = 1;
    129: op1_05_inv22 = 1;
    130: op1_05_inv22 = 1;
    default: op1_05_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in23 = reg_1302;
    53: op1_05_in23 = imem02_in[11:8];
    86: op1_05_in23 = reg_1198;
    69: op1_05_in23 = reg_0280;
    73: op1_05_in23 = reg_0490;
    61: op1_05_in23 = reg_0438;
    50: op1_05_in23 = reg_0285;
    71: op1_05_in23 = reg_0572;
    116: op1_05_in23 = reg_0572;
    54: op1_05_in23 = reg_0127;
    68: op1_05_in23 = reg_0236;
    74: op1_05_in23 = reg_0602;
    75: op1_05_in23 = reg_0371;
    56: op1_05_in23 = reg_0778;
    87: op1_05_in23 = reg_0487;
    76: op1_05_in23 = reg_1346;
    60: op1_05_in23 = reg_0832;
    46: op1_05_in23 = reg_0207;
    103: op1_05_in23 = reg_0207;
    57: op1_05_in23 = reg_0030;
    77: op1_05_in23 = reg_0163;
    48: op1_05_in23 = reg_0272;
    70: op1_05_in23 = reg_1001;
    58: op1_05_in23 = reg_0797;
    78: op1_05_in23 = reg_0161;
    88: op1_05_in23 = reg_1041;
    51: op1_05_in23 = reg_0675;
    79: op1_05_in23 = reg_0715;
    80: op1_05_in23 = reg_0021;
    62: op1_05_in23 = reg_0077;
    52: op1_05_in23 = reg_0108;
    81: op1_05_in23 = reg_0290;
    63: op1_05_in23 = reg_1149;
    82: op1_05_in23 = reg_0591;
    89: op1_05_in23 = reg_0470;
    83: op1_05_in23 = reg_0611;
    84: op1_05_in23 = reg_0267;
    47: op1_05_in23 = reg_0028;
    65: op1_05_in23 = reg_0094;
    85: op1_05_in23 = reg_0109;
    90: op1_05_in23 = reg_1298;
    66: op1_05_in23 = reg_0276;
    44: op1_05_in23 = reg_0182;
    91: op1_05_in23 = reg_0206;
    67: op1_05_in23 = reg_0673;
    92: op1_05_in23 = reg_0434;
    93: op1_05_in23 = reg_0320;
    42: op1_05_in23 = reg_0256;
    94: op1_05_in23 = reg_0177;
    96: op1_05_in23 = reg_1000;
    97: op1_05_in23 = reg_0145;
    99: op1_05_in23 = reg_0310;
    100: op1_05_in23 = reg_0902;
    101: op1_05_in23 = reg_0093;
    102: op1_05_in23 = reg_0211;
    105: op1_05_in23 = reg_1314;
    106: op1_05_in23 = reg_0800;
    108: op1_05_in23 = reg_0475;
    109: op1_05_in23 = reg_1430;
    110: op1_05_in23 = reg_1392;
    111: op1_05_in23 = reg_0345;
    112: op1_05_in23 = reg_0241;
    113: op1_05_in23 = reg_0040;
    114: op1_05_in23 = reg_0577;
    117: op1_05_in23 = reg_0137;
    118: op1_05_in23 = reg_0383;
    119: op1_05_in23 = reg_1456;
    120: op1_05_in23 = reg_0897;
    121: op1_05_in23 = reg_0836;
    122: op1_05_in23 = reg_0131;
    123: op1_05_in23 = imem05_in[15:12];
    124: op1_05_in23 = reg_1208;
    125: op1_05_in23 = reg_0469;
    126: op1_05_in23 = reg_1093;
    127: op1_05_in23 = reg_0679;
    128: op1_05_in23 = reg_1473;
    129: op1_05_in23 = reg_0135;
    130: op1_05_in23 = reg_0139;
    131: op1_05_in23 = reg_0833;
    default: op1_05_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv23 = 1;
    86: op1_05_inv23 = 1;
    73: op1_05_inv23 = 1;
    61: op1_05_inv23 = 1;
    50: op1_05_inv23 = 1;
    71: op1_05_inv23 = 1;
    68: op1_05_inv23 = 1;
    74: op1_05_inv23 = 1;
    56: op1_05_inv23 = 1;
    87: op1_05_inv23 = 1;
    76: op1_05_inv23 = 1;
    60: op1_05_inv23 = 1;
    46: op1_05_inv23 = 1;
    57: op1_05_inv23 = 1;
    77: op1_05_inv23 = 1;
    78: op1_05_inv23 = 1;
    88: op1_05_inv23 = 1;
    79: op1_05_inv23 = 1;
    62: op1_05_inv23 = 1;
    82: op1_05_inv23 = 1;
    65: op1_05_inv23 = 1;
    85: op1_05_inv23 = 1;
    67: op1_05_inv23 = 1;
    92: op1_05_inv23 = 1;
    93: op1_05_inv23 = 1;
    42: op1_05_inv23 = 1;
    94: op1_05_inv23 = 1;
    97: op1_05_inv23 = 1;
    102: op1_05_inv23 = 1;
    108: op1_05_inv23 = 1;
    110: op1_05_inv23 = 1;
    111: op1_05_inv23 = 1;
    112: op1_05_inv23 = 1;
    121: op1_05_inv23 = 1;
    124: op1_05_inv23 = 1;
    126: op1_05_inv23 = 1;
    127: op1_05_inv23 = 1;
    128: op1_05_inv23 = 1;
    131: op1_05_inv23 = 1;
    default: op1_05_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in24 = reg_0194;
    53: op1_05_in24 = reg_0496;
    86: op1_05_in24 = reg_0281;
    69: op1_05_in24 = reg_1132;
    73: op1_05_in24 = reg_0186;
    61: op1_05_in24 = reg_0728;
    50: op1_05_in24 = reg_0321;
    71: op1_05_in24 = reg_0819;
    54: op1_05_in24 = reg_0111;
    68: op1_05_in24 = reg_0129;
    74: op1_05_in24 = reg_0449;
    75: op1_05_in24 = reg_0018;
    56: op1_05_in24 = reg_0379;
    87: op1_05_in24 = reg_0837;
    76: op1_05_in24 = reg_0631;
    60: op1_05_in24 = reg_0395;
    46: op1_05_in24 = reg_0040;
    57: op1_05_in24 = reg_0366;
    77: op1_05_in24 = reg_0548;
    100: op1_05_in24 = reg_0548;
    48: op1_05_in24 = reg_0205;
    70: op1_05_in24 = reg_0965;
    58: op1_05_in24 = reg_0795;
    78: op1_05_in24 = reg_0115;
    88: op1_05_in24 = reg_1040;
    51: op1_05_in24 = imem03_in[7:4];
    79: op1_05_in24 = reg_0967;
    80: op1_05_in24 = reg_0470;
    62: op1_05_in24 = reg_1103;
    52: op1_05_in24 = reg_0107;
    81: op1_05_in24 = reg_0088;
    63: op1_05_in24 = reg_0177;
    82: op1_05_in24 = reg_0592;
    117: op1_05_in24 = reg_0592;
    89: op1_05_in24 = imem05_in[7:4];
    83: op1_05_in24 = reg_0448;
    84: op1_05_in24 = reg_0788;
    47: op1_05_in24 = reg_0228;
    65: op1_05_in24 = reg_0164;
    85: op1_05_in24 = reg_0584;
    90: op1_05_in24 = reg_0251;
    66: op1_05_in24 = reg_0311;
    44: op1_05_in24 = reg_0131;
    91: op1_05_in24 = reg_0038;
    67: op1_05_in24 = reg_1315;
    92: op1_05_in24 = reg_0147;
    93: op1_05_in24 = reg_1419;
    42: op1_05_in24 = reg_0563;
    94: op1_05_in24 = reg_0847;
    96: op1_05_in24 = reg_0840;
    97: op1_05_in24 = reg_0000;
    99: op1_05_in24 = reg_0170;
    101: op1_05_in24 = reg_0550;
    102: op1_05_in24 = reg_0021;
    103: op1_05_in24 = reg_0206;
    105: op1_05_in24 = reg_0954;
    106: op1_05_in24 = reg_0327;
    108: op1_05_in24 = reg_0905;
    109: op1_05_in24 = reg_0466;
    110: op1_05_in24 = imem02_in[11:8];
    111: op1_05_in24 = reg_0419;
    112: op1_05_in24 = reg_1473;
    113: op1_05_in24 = imem06_in[3:0];
    114: op1_05_in24 = reg_0731;
    116: op1_05_in24 = reg_0434;
    118: op1_05_in24 = reg_0091;
    119: op1_05_in24 = reg_0384;
    120: op1_05_in24 = reg_0801;
    121: op1_05_in24 = reg_0536;
    122: op1_05_in24 = reg_0697;
    123: op1_05_in24 = reg_0538;
    124: op1_05_in24 = reg_0104;
    125: op1_05_in24 = reg_0430;
    126: op1_05_in24 = reg_1092;
    127: op1_05_in24 = reg_0362;
    128: op1_05_in24 = reg_0715;
    129: op1_05_in24 = reg_0993;
    130: op1_05_in24 = reg_0777;
    131: op1_05_in24 = reg_0735;
    default: op1_05_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv24 = 1;
    53: op1_05_inv24 = 1;
    86: op1_05_inv24 = 1;
    73: op1_05_inv24 = 1;
    61: op1_05_inv24 = 1;
    74: op1_05_inv24 = 1;
    56: op1_05_inv24 = 1;
    60: op1_05_inv24 = 1;
    46: op1_05_inv24 = 1;
    57: op1_05_inv24 = 1;
    77: op1_05_inv24 = 1;
    48: op1_05_inv24 = 1;
    88: op1_05_inv24 = 1;
    51: op1_05_inv24 = 1;
    79: op1_05_inv24 = 1;
    80: op1_05_inv24 = 1;
    62: op1_05_inv24 = 1;
    52: op1_05_inv24 = 1;
    81: op1_05_inv24 = 1;
    82: op1_05_inv24 = 1;
    89: op1_05_inv24 = 1;
    83: op1_05_inv24 = 1;
    85: op1_05_inv24 = 1;
    66: op1_05_inv24 = 1;
    44: op1_05_inv24 = 1;
    91: op1_05_inv24 = 1;
    67: op1_05_inv24 = 1;
    92: op1_05_inv24 = 1;
    93: op1_05_inv24 = 1;
    101: op1_05_inv24 = 1;
    103: op1_05_inv24 = 1;
    106: op1_05_inv24 = 1;
    108: op1_05_inv24 = 1;
    109: op1_05_inv24 = 1;
    110: op1_05_inv24 = 1;
    112: op1_05_inv24 = 1;
    114: op1_05_inv24 = 1;
    120: op1_05_inv24 = 1;
    123: op1_05_inv24 = 1;
    124: op1_05_inv24 = 1;
    125: op1_05_inv24 = 1;
    126: op1_05_inv24 = 1;
    129: op1_05_inv24 = 1;
    130: op1_05_inv24 = 1;
    131: op1_05_inv24 = 1;
    default: op1_05_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in25 = reg_0584;
    53: op1_05_in25 = reg_0472;
    86: op1_05_in25 = reg_0500;
    69: op1_05_in25 = reg_0235;
    73: op1_05_in25 = reg_0298;
    61: op1_05_in25 = reg_0091;
    50: op1_05_in25 = reg_0228;
    117: op1_05_in25 = reg_0228;
    71: op1_05_in25 = reg_0439;
    54: op1_05_in25 = reg_0105;
    68: op1_05_in25 = reg_0016;
    74: op1_05_in25 = reg_0206;
    75: op1_05_in25 = imem07_in[15:12];
    56: op1_05_in25 = reg_0903;
    87: op1_05_in25 = reg_1151;
    76: op1_05_in25 = reg_0151;
    60: op1_05_in25 = reg_0700;
    46: op1_05_in25 = reg_0784;
    57: op1_05_in25 = reg_0740;
    77: op1_05_in25 = reg_0743;
    48: op1_05_in25 = reg_0014;
    70: op1_05_in25 = reg_0314;
    58: op1_05_in25 = reg_0488;
    78: op1_05_in25 = reg_0116;
    88: op1_05_in25 = reg_0451;
    51: op1_05_in25 = reg_0444;
    79: op1_05_in25 = reg_0968;
    80: op1_05_in25 = reg_0737;
    62: op1_05_in25 = reg_0606;
    52: op1_05_in25 = reg_0479;
    81: op1_05_in25 = reg_0291;
    63: op1_05_in25 = reg_0142;
    82: op1_05_in25 = reg_0100;
    89: op1_05_in25 = reg_0205;
    83: op1_05_in25 = reg_1253;
    84: op1_05_in25 = reg_0754;
    47: op1_05_in25 = reg_0003;
    65: op1_05_in25 = reg_0150;
    85: op1_05_in25 = reg_0526;
    90: op1_05_in25 = reg_1431;
    66: op1_05_in25 = reg_0573;
    44: op1_05_in25 = reg_0333;
    91: op1_05_in25 = reg_0040;
    67: op1_05_in25 = reg_0667;
    92: op1_05_in25 = reg_0149;
    93: op1_05_in25 = reg_0236;
    42: op1_05_in25 = reg_0562;
    94: op1_05_in25 = reg_0234;
    96: op1_05_in25 = reg_0889;
    97: op1_05_in25 = reg_0375;
    99: op1_05_in25 = reg_0923;
    100: op1_05_in25 = reg_0746;
    101: op1_05_in25 = reg_0548;
    102: op1_05_in25 = reg_1488;
    103: op1_05_in25 = reg_0039;
    105: op1_05_in25 = reg_0957;
    106: op1_05_in25 = reg_0848;
    120: op1_05_in25 = reg_0848;
    108: op1_05_in25 = reg_0870;
    109: op1_05_in25 = reg_0346;
    110: op1_05_in25 = reg_0845;
    111: op1_05_in25 = reg_0308;
    112: op1_05_in25 = reg_0572;
    113: op1_05_in25 = reg_0670;
    114: op1_05_in25 = reg_0797;
    116: op1_05_in25 = reg_0384;
    118: op1_05_in25 = reg_0634;
    119: op1_05_in25 = reg_0383;
    121: op1_05_in25 = reg_0470;
    122: op1_05_in25 = reg_0938;
    123: op1_05_in25 = reg_0890;
    124: op1_05_in25 = reg_0350;
    125: op1_05_in25 = reg_1032;
    128: op1_05_in25 = reg_1032;
    126: op1_05_in25 = reg_0108;
    127: op1_05_in25 = reg_0365;
    129: op1_05_in25 = reg_1315;
    130: op1_05_in25 = reg_0031;
    131: op1_05_in25 = reg_0733;
    default: op1_05_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_05_inv25 = 1;
    73: op1_05_inv25 = 1;
    61: op1_05_inv25 = 1;
    71: op1_05_inv25 = 1;
    54: op1_05_inv25 = 1;
    76: op1_05_inv25 = 1;
    46: op1_05_inv25 = 1;
    57: op1_05_inv25 = 1;
    48: op1_05_inv25 = 1;
    51: op1_05_inv25 = 1;
    79: op1_05_inv25 = 1;
    62: op1_05_inv25 = 1;
    81: op1_05_inv25 = 1;
    63: op1_05_inv25 = 1;
    89: op1_05_inv25 = 1;
    83: op1_05_inv25 = 1;
    84: op1_05_inv25 = 1;
    47: op1_05_inv25 = 1;
    65: op1_05_inv25 = 1;
    92: op1_05_inv25 = 1;
    93: op1_05_inv25 = 1;
    42: op1_05_inv25 = 1;
    96: op1_05_inv25 = 1;
    99: op1_05_inv25 = 1;
    100: op1_05_inv25 = 1;
    101: op1_05_inv25 = 1;
    102: op1_05_inv25 = 1;
    105: op1_05_inv25 = 1;
    108: op1_05_inv25 = 1;
    110: op1_05_inv25 = 1;
    114: op1_05_inv25 = 1;
    116: op1_05_inv25 = 1;
    117: op1_05_inv25 = 1;
    120: op1_05_inv25 = 1;
    121: op1_05_inv25 = 1;
    122: op1_05_inv25 = 1;
    123: op1_05_inv25 = 1;
    125: op1_05_inv25 = 1;
    127: op1_05_inv25 = 1;
    128: op1_05_inv25 = 1;
    130: op1_05_inv25 = 1;
    default: op1_05_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in26 = reg_0619;
    53: op1_05_in26 = reg_0474;
    86: op1_05_in26 = reg_0796;
    69: op1_05_in26 = reg_0177;
    73: op1_05_in26 = reg_0667;
    61: op1_05_in26 = reg_0011;
    50: op1_05_in26 = reg_0051;
    71: op1_05_in26 = reg_0149;
    54: op1_05_in26 = reg_0056;
    68: op1_05_in26 = reg_0792;
    74: op1_05_in26 = reg_0754;
    111: op1_05_in26 = reg_0754;
    75: op1_05_in26 = reg_0461;
    56: op1_05_in26 = reg_0900;
    87: op1_05_in26 = reg_0236;
    76: op1_05_in26 = reg_0828;
    60: op1_05_in26 = reg_0646;
    46: op1_05_in26 = reg_0160;
    57: op1_05_in26 = reg_0738;
    77: op1_05_in26 = reg_0242;
    48: op1_05_in26 = reg_0194;
    70: op1_05_in26 = reg_0952;
    58: op1_05_in26 = reg_0596;
    78: op1_05_in26 = reg_0585;
    88: op1_05_in26 = reg_0097;
    51: op1_05_in26 = reg_0185;
    79: op1_05_in26 = reg_0439;
    80: op1_05_in26 = reg_0176;
    62: op1_05_in26 = reg_0532;
    42: op1_05_in26 = reg_0532;
    52: op1_05_in26 = reg_0330;
    81: op1_05_in26 = reg_0043;
    118: op1_05_in26 = reg_0043;
    63: op1_05_in26 = reg_1001;
    82: op1_05_in26 = reg_0321;
    89: op1_05_in26 = reg_1431;
    83: op1_05_in26 = reg_0549;
    84: op1_05_in26 = reg_0166;
    47: op1_05_in26 = reg_0518;
    65: op1_05_in26 = reg_0211;
    85: op1_05_in26 = reg_0528;
    90: op1_05_in26 = reg_0332;
    66: op1_05_in26 = reg_0677;
    44: op1_05_in26 = reg_0541;
    91: op1_05_in26 = reg_0039;
    67: op1_05_in26 = reg_0245;
    92: op1_05_in26 = reg_0148;
    93: op1_05_in26 = reg_1107;
    94: op1_05_in26 = reg_1494;
    96: op1_05_in26 = reg_0328;
    97: op1_05_in26 = reg_0142;
    99: op1_05_in26 = reg_1094;
    100: op1_05_in26 = reg_0610;
    101: op1_05_in26 = reg_0610;
    102: op1_05_in26 = reg_0877;
    103: op1_05_in26 = imem06_in[15:12];
    105: op1_05_in26 = reg_1301;
    106: op1_05_in26 = reg_0068;
    108: op1_05_in26 = reg_1209;
    109: op1_05_in26 = reg_0173;
    110: op1_05_in26 = reg_0561;
    112: op1_05_in26 = reg_0430;
    113: op1_05_in26 = reg_0729;
    114: op1_05_in26 = reg_0531;
    116: op1_05_in26 = reg_0363;
    128: op1_05_in26 = reg_0363;
    117: op1_05_in26 = reg_0004;
    119: op1_05_in26 = reg_0362;
    120: op1_05_in26 = reg_0217;
    121: op1_05_in26 = reg_0650;
    122: op1_05_in26 = reg_1514;
    123: op1_05_in26 = reg_0272;
    124: op1_05_in26 = reg_1149;
    125: op1_05_in26 = reg_0092;
    126: op1_05_in26 = reg_0790;
    127: op1_05_in26 = reg_0901;
    129: op1_05_in26 = reg_0457;
    130: op1_05_in26 = reg_0740;
    131: op1_05_in26 = reg_0340;
    default: op1_05_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv26 = 1;
    53: op1_05_inv26 = 1;
    86: op1_05_inv26 = 1;
    69: op1_05_inv26 = 1;
    61: op1_05_inv26 = 1;
    74: op1_05_inv26 = 1;
    75: op1_05_inv26 = 1;
    87: op1_05_inv26 = 1;
    60: op1_05_inv26 = 1;
    57: op1_05_inv26 = 1;
    77: op1_05_inv26 = 1;
    48: op1_05_inv26 = 1;
    58: op1_05_inv26 = 1;
    79: op1_05_inv26 = 1;
    62: op1_05_inv26 = 1;
    81: op1_05_inv26 = 1;
    63: op1_05_inv26 = 1;
    65: op1_05_inv26 = 1;
    85: op1_05_inv26 = 1;
    44: op1_05_inv26 = 1;
    67: op1_05_inv26 = 1;
    92: op1_05_inv26 = 1;
    96: op1_05_inv26 = 1;
    100: op1_05_inv26 = 1;
    103: op1_05_inv26 = 1;
    108: op1_05_inv26 = 1;
    109: op1_05_inv26 = 1;
    113: op1_05_inv26 = 1;
    117: op1_05_inv26 = 1;
    118: op1_05_inv26 = 1;
    121: op1_05_inv26 = 1;
    123: op1_05_inv26 = 1;
    126: op1_05_inv26 = 1;
    128: op1_05_inv26 = 1;
    131: op1_05_inv26 = 1;
    default: op1_05_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in27 = reg_1228;
    53: op1_05_in27 = reg_0990;
    86: op1_05_in27 = reg_1147;
    69: op1_05_in27 = imem03_in[7:4];
    73: op1_05_in27 = reg_0892;
    61: op1_05_in27 = reg_0010;
    50: op1_05_in27 = reg_0003;
    71: op1_05_in27 = reg_0146;
    54: op1_05_in27 = reg_0390;
    68: op1_05_in27 = reg_0315;
    74: op1_05_in27 = reg_0466;
    75: op1_05_in27 = reg_0158;
    129: op1_05_in27 = reg_0158;
    56: op1_05_in27 = reg_0153;
    87: op1_05_in27 = reg_1107;
    76: op1_05_in27 = reg_0040;
    60: op1_05_in27 = reg_0567;
    46: op1_05_in27 = reg_0906;
    57: op1_05_in27 = reg_0623;
    77: op1_05_in27 = reg_0742;
    48: op1_05_in27 = reg_0193;
    70: op1_05_in27 = reg_1199;
    58: op1_05_in27 = reg_0368;
    78: op1_05_in27 = reg_0584;
    88: op1_05_in27 = reg_0061;
    51: op1_05_in27 = reg_0179;
    79: op1_05_in27 = reg_1456;
    80: op1_05_in27 = reg_0648;
    62: op1_05_in27 = reg_0253;
    52: op1_05_in27 = reg_0329;
    81: op1_05_in27 = reg_0042;
    63: op1_05_in27 = reg_0965;
    94: op1_05_in27 = reg_0965;
    82: op1_05_in27 = reg_0361;
    89: op1_05_in27 = reg_0136;
    83: op1_05_in27 = reg_0548;
    84: op1_05_in27 = reg_0930;
    47: op1_05_in27 = reg_0520;
    65: op1_05_in27 = reg_0034;
    85: op1_05_in27 = reg_0569;
    90: op1_05_in27 = reg_0604;
    66: op1_05_in27 = reg_0216;
    44: op1_05_in27 = reg_0539;
    91: op1_05_in27 = reg_0014;
    67: op1_05_in27 = reg_0225;
    92: op1_05_in27 = reg_0092;
    128: op1_05_in27 = reg_0092;
    93: op1_05_in27 = reg_0209;
    42: op1_05_in27 = reg_0530;
    96: op1_05_in27 = reg_0709;
    97: op1_05_in27 = reg_0190;
    99: op1_05_in27 = reg_0779;
    100: op1_05_in27 = reg_0242;
    101: op1_05_in27 = reg_0222;
    102: op1_05_in27 = reg_0204;
    103: op1_05_in27 = reg_0931;
    105: op1_05_in27 = reg_1208;
    106: op1_05_in27 = reg_0009;
    120: op1_05_in27 = reg_0009;
    108: op1_05_in27 = reg_0271;
    109: op1_05_in27 = reg_0045;
    110: op1_05_in27 = reg_0254;
    111: op1_05_in27 = reg_0195;
    112: op1_05_in27 = reg_0434;
    113: op1_05_in27 = reg_0784;
    114: op1_05_in27 = reg_0297;
    116: op1_05_in27 = reg_0335;
    117: op1_05_in27 = reg_0085;
    118: op1_05_in27 = reg_0327;
    119: op1_05_in27 = reg_0899;
    121: op1_05_in27 = imem05_in[11:8];
    122: op1_05_in27 = reg_0300;
    123: op1_05_in27 = reg_0992;
    124: op1_05_in27 = reg_1139;
    125: op1_05_in27 = reg_0595;
    126: op1_05_in27 = imem04_in[3:0];
    127: op1_05_in27 = reg_0175;
    130: op1_05_in27 = reg_0592;
    131: op1_05_in27 = reg_0793;
    default: op1_05_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_05_inv27 = 1;
    86: op1_05_inv27 = 1;
    69: op1_05_inv27 = 1;
    73: op1_05_inv27 = 1;
    50: op1_05_inv27 = 1;
    71: op1_05_inv27 = 1;
    54: op1_05_inv27 = 1;
    68: op1_05_inv27 = 1;
    74: op1_05_inv27 = 1;
    56: op1_05_inv27 = 1;
    76: op1_05_inv27 = 1;
    60: op1_05_inv27 = 1;
    46: op1_05_inv27 = 1;
    57: op1_05_inv27 = 1;
    48: op1_05_inv27 = 1;
    58: op1_05_inv27 = 1;
    78: op1_05_inv27 = 1;
    51: op1_05_inv27 = 1;
    62: op1_05_inv27 = 1;
    52: op1_05_inv27 = 1;
    65: op1_05_inv27 = 1;
    85: op1_05_inv27 = 1;
    90: op1_05_inv27 = 1;
    66: op1_05_inv27 = 1;
    42: op1_05_inv27 = 1;
    94: op1_05_inv27 = 1;
    99: op1_05_inv27 = 1;
    105: op1_05_inv27 = 1;
    106: op1_05_inv27 = 1;
    108: op1_05_inv27 = 1;
    112: op1_05_inv27 = 1;
    114: op1_05_inv27 = 1;
    118: op1_05_inv27 = 1;
    121: op1_05_inv27 = 1;
    123: op1_05_inv27 = 1;
    125: op1_05_inv27 = 1;
    127: op1_05_inv27 = 1;
    129: op1_05_inv27 = 1;
    default: op1_05_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in28 = reg_1204;
    53: op1_05_in28 = reg_0991;
    86: op1_05_in28 = reg_1041;
    69: op1_05_in28 = reg_0261;
    73: op1_05_in28 = reg_0310;
    61: op1_05_in28 = reg_0222;
    50: op1_05_in28 = reg_0084;
    71: op1_05_in28 = reg_0402;
    54: op1_05_in28 = reg_0897;
    68: op1_05_in28 = reg_0168;
    120: op1_05_in28 = reg_0168;
    74: op1_05_in28 = reg_0377;
    75: op1_05_in28 = reg_0157;
    56: op1_05_in28 = reg_0878;
    87: op1_05_in28 = reg_0209;
    76: op1_05_in28 = reg_0754;
    60: op1_05_in28 = reg_0566;
    46: op1_05_in28 = imem06_in[7:4];
    57: op1_05_in28 = reg_0618;
    77: op1_05_in28 = reg_0715;
    48: op1_05_in28 = reg_0192;
    113: op1_05_in28 = reg_0192;
    70: op1_05_in28 = reg_1092;
    58: op1_05_in28 = reg_0836;
    78: op1_05_in28 = reg_0619;
    88: op1_05_in28 = reg_0837;
    51: op1_05_in28 = reg_0957;
    79: op1_05_in28 = reg_0149;
    80: op1_05_in28 = reg_1181;
    62: op1_05_in28 = reg_0589;
    52: op1_05_in28 = reg_0426;
    81: op1_05_in28 = reg_0011;
    63: op1_05_in28 = reg_0962;
    82: op1_05_in28 = reg_0085;
    89: op1_05_in28 = reg_0702;
    83: op1_05_in28 = reg_0747;
    84: op1_05_in28 = reg_0547;
    47: op1_05_in28 = reg_0483;
    65: op1_05_in28 = reg_0792;
    85: op1_05_in28 = reg_0295;
    90: op1_05_in28 = reg_0562;
    66: op1_05_in28 = reg_0227;
    44: op1_05_in28 = imem05_in[15:12];
    91: op1_05_in28 = imem06_in[15:12];
    67: op1_05_in28 = reg_0309;
    92: op1_05_in28 = reg_0595;
    93: op1_05_in28 = reg_0536;
    42: op1_05_in28 = reg_0533;
    94: op1_05_in28 = reg_0349;
    96: op1_05_in28 = reg_0330;
    97: op1_05_in28 = reg_1300;
    99: op1_05_in28 = reg_0774;
    100: op1_05_in28 = reg_0820;
    101: op1_05_in28 = reg_0830;
    102: op1_05_in28 = reg_0986;
    121: op1_05_in28 = reg_0986;
    103: op1_05_in28 = reg_0906;
    105: op1_05_in28 = reg_0107;
    106: op1_05_in28 = imem03_in[11:8];
    108: op1_05_in28 = reg_0720;
    109: op1_05_in28 = reg_1180;
    110: op1_05_in28 = reg_0133;
    111: op1_05_in28 = reg_0215;
    112: op1_05_in28 = reg_0438;
    114: op1_05_in28 = reg_1200;
    116: op1_05_in28 = reg_0080;
    117: op1_05_in28 = reg_0123;
    118: op1_05_in28 = reg_0889;
    119: op1_05_in28 = reg_0175;
    128: op1_05_in28 = reg_0175;
    122: op1_05_in28 = reg_0090;
    123: op1_05_in28 = reg_0649;
    124: op1_05_in28 = reg_0348;
    125: op1_05_in28 = reg_0012;
    126: op1_05_in28 = reg_1384;
    127: op1_05_in28 = reg_0464;
    129: op1_05_in28 = reg_0489;
    130: op1_05_in28 = reg_0001;
    131: op1_05_in28 = reg_0045;
    default: op1_05_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv28 = 1;
    86: op1_05_inv28 = 1;
    69: op1_05_inv28 = 1;
    61: op1_05_inv28 = 1;
    71: op1_05_inv28 = 1;
    54: op1_05_inv28 = 1;
    68: op1_05_inv28 = 1;
    74: op1_05_inv28 = 1;
    75: op1_05_inv28 = 1;
    56: op1_05_inv28 = 1;
    87: op1_05_inv28 = 1;
    46: op1_05_inv28 = 1;
    77: op1_05_inv28 = 1;
    70: op1_05_inv28 = 1;
    58: op1_05_inv28 = 1;
    88: op1_05_inv28 = 1;
    79: op1_05_inv28 = 1;
    89: op1_05_inv28 = 1;
    83: op1_05_inv28 = 1;
    84: op1_05_inv28 = 1;
    85: op1_05_inv28 = 1;
    90: op1_05_inv28 = 1;
    66: op1_05_inv28 = 1;
    91: op1_05_inv28 = 1;
    67: op1_05_inv28 = 1;
    93: op1_05_inv28 = 1;
    94: op1_05_inv28 = 1;
    96: op1_05_inv28 = 1;
    97: op1_05_inv28 = 1;
    99: op1_05_inv28 = 1;
    105: op1_05_inv28 = 1;
    106: op1_05_inv28 = 1;
    113: op1_05_inv28 = 1;
    114: op1_05_inv28 = 1;
    117: op1_05_inv28 = 1;
    119: op1_05_inv28 = 1;
    120: op1_05_inv28 = 1;
    122: op1_05_inv28 = 1;
    123: op1_05_inv28 = 1;
    127: op1_05_inv28 = 1;
    129: op1_05_inv28 = 1;
    130: op1_05_inv28 = 1;
    131: op1_05_inv28 = 1;
    default: op1_05_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in29 = reg_0213;
    53: op1_05_in29 = reg_0125;
    86: op1_05_in29 = reg_1040;
    69: op1_05_in29 = reg_1233;
    73: op1_05_in29 = reg_0703;
    61: op1_05_in29 = reg_0457;
    50: op1_05_in29 = reg_0087;
    71: op1_05_in29 = reg_0384;
    79: op1_05_in29 = reg_0384;
    54: op1_05_in29 = reg_0839;
    68: op1_05_in29 = reg_0173;
    74: op1_05_in29 = reg_0399;
    62: op1_05_in29 = reg_0399;
    75: op1_05_in29 = reg_0923;
    56: op1_05_in29 = reg_0007;
    87: op1_05_in29 = reg_0063;
    93: op1_05_in29 = reg_0063;
    76: op1_05_in29 = reg_0466;
    60: op1_05_in29 = reg_0745;
    46: op1_05_in29 = reg_0870;
    57: op1_05_in29 = reg_0050;
    77: op1_05_in29 = reg_0968;
    48: op1_05_in29 = imem06_in[3:0];
    70: op1_05_in29 = reg_0831;
    58: op1_05_in29 = reg_0164;
    78: op1_05_in29 = reg_0571;
    88: op1_05_in29 = reg_0117;
    51: op1_05_in29 = reg_0597;
    80: op1_05_in29 = reg_0697;
    90: op1_05_in29 = reg_0697;
    109: op1_05_in29 = reg_0697;
    131: op1_05_in29 = reg_0697;
    52: op1_05_in29 = reg_0582;
    81: op1_05_in29 = reg_1493;
    63: op1_05_in29 = reg_0246;
    82: op1_05_in29 = reg_0084;
    89: op1_05_in29 = reg_0174;
    83: op1_05_in29 = reg_0242;
    84: op1_05_in29 = reg_0610;
    65: op1_05_in29 = reg_0794;
    85: op1_05_in29 = reg_0289;
    66: op1_05_in29 = reg_0710;
    44: op1_05_in29 = reg_0477;
    91: op1_05_in29 = reg_0396;
    67: op1_05_in29 = reg_0924;
    92: op1_05_in29 = reg_0464;
    128: op1_05_in29 = reg_0464;
    42: op1_05_in29 = reg_0473;
    94: op1_05_in29 = reg_1313;
    96: op1_05_in29 = reg_0198;
    97: op1_05_in29 = reg_0178;
    99: op1_05_in29 = reg_0030;
    100: op1_05_in29 = reg_1475;
    101: op1_05_in29 = reg_0798;
    102: op1_05_in29 = reg_0735;
    121: op1_05_in29 = reg_0735;
    103: op1_05_in29 = reg_1467;
    105: op1_05_in29 = reg_0104;
    106: op1_05_in29 = reg_0377;
    108: op1_05_in29 = reg_1179;
    110: op1_05_in29 = reg_0900;
    111: op1_05_in29 = reg_0017;
    112: op1_05_in29 = reg_0149;
    113: op1_05_in29 = reg_0696;
    114: op1_05_in29 = reg_0500;
    116: op1_05_in29 = reg_0042;
    117: op1_05_in29 = reg_1182;
    118: op1_05_in29 = imem02_in[3:0];
    119: op1_05_in29 = reg_0727;
    120: op1_05_in29 = reg_0632;
    122: op1_05_in29 = reg_0873;
    123: op1_05_in29 = reg_1104;
    124: op1_05_in29 = reg_0425;
    125: op1_05_in29 = reg_0011;
    126: op1_05_in29 = reg_0016;
    127: op1_05_in29 = reg_0080;
    129: op1_05_in29 = reg_0224;
    130: op1_05_in29 = reg_0404;
    default: op1_05_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv29 = 1;
    53: op1_05_inv29 = 1;
    86: op1_05_inv29 = 1;
    69: op1_05_inv29 = 1;
    71: op1_05_inv29 = 1;
    68: op1_05_inv29 = 1;
    74: op1_05_inv29 = 1;
    75: op1_05_inv29 = 1;
    56: op1_05_inv29 = 1;
    76: op1_05_inv29 = 1;
    48: op1_05_inv29 = 1;
    78: op1_05_inv29 = 1;
    88: op1_05_inv29 = 1;
    51: op1_05_inv29 = 1;
    80: op1_05_inv29 = 1;
    62: op1_05_inv29 = 1;
    81: op1_05_inv29 = 1;
    82: op1_05_inv29 = 1;
    89: op1_05_inv29 = 1;
    65: op1_05_inv29 = 1;
    90: op1_05_inv29 = 1;
    44: op1_05_inv29 = 1;
    42: op1_05_inv29 = 1;
    96: op1_05_inv29 = 1;
    99: op1_05_inv29 = 1;
    100: op1_05_inv29 = 1;
    102: op1_05_inv29 = 1;
    106: op1_05_inv29 = 1;
    109: op1_05_inv29 = 1;
    111: op1_05_inv29 = 1;
    112: op1_05_inv29 = 1;
    117: op1_05_inv29 = 1;
    119: op1_05_inv29 = 1;
    120: op1_05_inv29 = 1;
    121: op1_05_inv29 = 1;
    123: op1_05_inv29 = 1;
    125: op1_05_inv29 = 1;
    127: op1_05_inv29 = 1;
    129: op1_05_inv29 = 1;
    131: op1_05_inv29 = 1;
    default: op1_05_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_05_in30 = imem07_in[3:0];
    111: op1_05_in30 = imem07_in[3:0];
    53: op1_05_in30 = reg_0105;
    86: op1_05_in30 = reg_0199;
    69: op1_05_in30 = reg_1231;
    73: op1_05_in30 = reg_0170;
    61: op1_05_in30 = reg_0255;
    50: op1_05_in30 = reg_0124;
    71: op1_05_in30 = reg_0360;
    54: op1_05_in30 = reg_0009;
    68: op1_05_in30 = reg_0346;
    74: op1_05_in30 = reg_0541;
    75: op1_05_in30 = reg_0774;
    56: op1_05_in30 = reg_0121;
    87: op1_05_in30 = reg_1502;
    76: op1_05_in30 = reg_1436;
    60: op1_05_in30 = reg_0697;
    46: op1_05_in30 = reg_0396;
    57: op1_05_in30 = reg_0484;
    77: op1_05_in30 = reg_0439;
    100: op1_05_in30 = reg_0439;
    48: op1_05_in30 = imem06_in[7:4];
    70: op1_05_in30 = reg_0525;
    58: op1_05_in30 = reg_0032;
    78: op1_05_in30 = reg_1228;
    88: op1_05_in30 = reg_0063;
    51: op1_05_in30 = reg_0246;
    79: op1_05_in30 = reg_0899;
    80: op1_05_in30 = reg_1403;
    62: op1_05_in30 = reg_0612;
    52: op1_05_in30 = reg_0744;
    81: op1_05_in30 = reg_0744;
    63: op1_05_in30 = reg_1199;
    82: op1_05_in30 = reg_0087;
    89: op1_05_in30 = reg_0066;
    83: op1_05_in30 = reg_0241;
    84: op1_05_in30 = reg_0798;
    65: op1_05_in30 = reg_0347;
    85: op1_05_in30 = reg_1202;
    90: op1_05_in30 = reg_1401;
    66: op1_05_in30 = reg_1063;
    44: op1_05_in30 = reg_0895;
    91: op1_05_in30 = reg_1030;
    67: op1_05_in30 = reg_0223;
    92: op1_05_in30 = reg_0077;
    93: op1_05_in30 = reg_0019;
    42: op1_05_in30 = reg_0475;
    94: op1_05_in30 = reg_0884;
    96: op1_05_in30 = reg_0847;
    97: op1_05_in30 = reg_0885;
    105: op1_05_in30 = reg_0885;
    99: op1_05_in30 = reg_0442;
    101: op1_05_in30 = reg_0572;
    102: op1_05_in30 = reg_1430;
    103: op1_05_in30 = reg_0860;
    106: op1_05_in30 = reg_0699;
    108: op1_05_in30 = reg_0780;
    109: op1_05_in30 = reg_1402;
    110: op1_05_in30 = reg_0495;
    112: op1_05_in30 = reg_0146;
    113: op1_05_in30 = reg_0271;
    114: op1_05_in30 = reg_0407;
    116: op1_05_in30 = reg_1071;
    118: op1_05_in30 = reg_1235;
    119: op1_05_in30 = reg_0257;
    120: op1_05_in30 = reg_0999;
    121: op1_05_in30 = reg_0136;
    122: op1_05_in30 = reg_0736;
    123: op1_05_in30 = reg_1181;
    124: op1_05_in30 = reg_0411;
    125: op1_05_in30 = reg_0668;
    126: op1_05_in30 = reg_1216;
    127: op1_05_in30 = reg_0403;
    128: op1_05_in30 = reg_0335;
    129: op1_05_in30 = reg_0777;
    130: op1_05_in30 = reg_0483;
    131: op1_05_in30 = reg_0939;
    default: op1_05_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_05_inv30 = 1;
    86: op1_05_inv30 = 1;
    69: op1_05_inv30 = 1;
    73: op1_05_inv30 = 1;
    61: op1_05_inv30 = 1;
    71: op1_05_inv30 = 1;
    54: op1_05_inv30 = 1;
    87: op1_05_inv30 = 1;
    76: op1_05_inv30 = 1;
    57: op1_05_inv30 = 1;
    48: op1_05_inv30 = 1;
    58: op1_05_inv30 = 1;
    78: op1_05_inv30 = 1;
    88: op1_05_inv30 = 1;
    62: op1_05_inv30 = 1;
    81: op1_05_inv30 = 1;
    63: op1_05_inv30 = 1;
    82: op1_05_inv30 = 1;
    89: op1_05_inv30 = 1;
    83: op1_05_inv30 = 1;
    84: op1_05_inv30 = 1;
    65: op1_05_inv30 = 1;
    90: op1_05_inv30 = 1;
    44: op1_05_inv30 = 1;
    91: op1_05_inv30 = 1;
    67: op1_05_inv30 = 1;
    92: op1_05_inv30 = 1;
    93: op1_05_inv30 = 1;
    42: op1_05_inv30 = 1;
    94: op1_05_inv30 = 1;
    97: op1_05_inv30 = 1;
    100: op1_05_inv30 = 1;
    102: op1_05_inv30 = 1;
    105: op1_05_inv30 = 1;
    109: op1_05_inv30 = 1;
    112: op1_05_inv30 = 1;
    113: op1_05_inv30 = 1;
    118: op1_05_inv30 = 1;
    119: op1_05_inv30 = 1;
    121: op1_05_inv30 = 1;
    122: op1_05_inv30 = 1;
    125: op1_05_inv30 = 1;
    127: op1_05_inv30 = 1;
    128: op1_05_inv30 = 1;
    130: op1_05_inv30 = 1;
    131: op1_05_inv30 = 1;
    default: op1_05_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_05_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#5の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_05_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in00 = reg_1281;
    82: op1_06_in00 = reg_1281;
    53: op1_06_in00 = reg_0932;
    55: op1_06_in00 = reg_0399;
    86: op1_06_in00 = reg_1425;
    73: op1_06_in00 = reg_0631;
    69: op1_06_in00 = reg_0222;
    49: op1_06_in00 = reg_0297;
    71: op1_06_in00 = reg_0824;
    95: op1_06_in00 = reg_0824;
    50: op1_06_in00 = reg_0271;
    54: op1_06_in00 = reg_0968;
    74: op1_06_in00 = reg_0580;
    68: op1_06_in00 = reg_0997;
    61: op1_06_in00 = reg_0614;
    75: op1_06_in00 = reg_0219;
    87: op1_06_in00 = reg_0375;
    56: op1_06_in00 = reg_0940;
    76: op1_06_in00 = reg_0613;
    60: op1_06_in00 = reg_0000;
    57: op1_06_in00 = reg_0960;
    77: op1_06_in00 = reg_0983;
    98: op1_06_in00 = reg_0983;
    33: op1_06_in00 = reg_0170;
    70: op1_06_in00 = reg_0699;
    124: op1_06_in00 = reg_0699;
    58: op1_06_in00 = reg_0171;
    48: op1_06_in00 = reg_0750;
    78: op1_06_in00 = imem06_in[11:8];
    46: op1_06_in00 = reg_0823;
    88: op1_06_in00 = reg_1314;
    51: op1_06_in00 = reg_0245;
    79: op1_06_in00 = reg_0347;
    59: op1_06_in00 = reg_0149;
    28: op1_06_in00 = imem07_in[3:0];
    40: op1_06_in00 = imem07_in[3:0];
    80: op1_06_in00 = reg_1384;
    62: op1_06_in00 = reg_0874;
    52: op1_06_in00 = reg_0899;
    81: op1_06_in00 = reg_0590;
    63: op1_06_in00 = reg_0345;
    89: op1_06_in00 = reg_0233;
    120: op1_06_in00 = reg_0233;
    83: op1_06_in00 = reg_0209;
    64: op1_06_in00 = reg_0042;
    127: op1_06_in00 = reg_0042;
    22: op1_06_in00 = imem07_in[15:12];
    34: op1_06_in00 = imem07_in[15:12];
    111: op1_06_in00 = imem07_in[15:12];
    37: op1_06_in00 = reg_0441;
    84: op1_06_in00 = reg_1474;
    47: op1_06_in00 = imem07_in[7:4];
    65: op1_06_in00 = reg_0488;
    85: op1_06_in00 = reg_0791;
    90: op1_06_in00 = reg_0078;
    66: op1_06_in00 = reg_0046;
    91: op1_06_in00 = reg_1244;
    44: op1_06_in00 = reg_0795;
    67: op1_06_in00 = reg_1001;
    92: op1_06_in00 = reg_1068;
    93: op1_06_in00 = reg_0370;
    94: op1_06_in00 = reg_0707;
    96: op1_06_in00 = reg_0311;
    42: op1_06_in00 = reg_0746;
    97: op1_06_in00 = reg_0882;
    99: op1_06_in00 = reg_1079;
    100: op1_06_in00 = reg_0595;
    101: op1_06_in00 = reg_1456;
    102: op1_06_in00 = reg_0833;
    103: op1_06_in00 = reg_0863;
    104: op1_06_in00 = reg_0121;
    105: op1_06_in00 = reg_0541;
    106: op1_06_in00 = reg_0154;
    107: op1_06_in00 = reg_1081;
    108: op1_06_in00 = reg_0716;
    109: op1_06_in00 = reg_0274;
    110: op1_06_in00 = reg_0432;
    112: op1_06_in00 = reg_0384;
    113: op1_06_in00 = reg_1326;
    114: op1_06_in00 = reg_0471;
    115: op1_06_in00 = imem00_in[3:0];
    116: op1_06_in00 = reg_0606;
    38: op1_06_in00 = reg_0672;
    117: op1_06_in00 = imem00_in[11:8];
    118: op1_06_in00 = reg_0588;
    119: op1_06_in00 = reg_0162;
    121: op1_06_in00 = reg_0272;
    122: op1_06_in00 = reg_0197;
    123: op1_06_in00 = reg_0697;
    125: op1_06_in00 = imem02_in[3:0];
    126: op1_06_in00 = reg_0032;
    128: op1_06_in00 = reg_0079;
    129: op1_06_in00 = reg_0287;
    130: op1_06_in00 = imem00_in[15:12];
    131: op1_06_in00 = reg_1163;
    default: op1_06_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv00 = 1;
    86: op1_06_inv00 = 1;
    73: op1_06_inv00 = 1;
    69: op1_06_inv00 = 1;
    71: op1_06_inv00 = 1;
    54: op1_06_inv00 = 1;
    74: op1_06_inv00 = 1;
    61: op1_06_inv00 = 1;
    87: op1_06_inv00 = 1;
    56: op1_06_inv00 = 1;
    76: op1_06_inv00 = 1;
    60: op1_06_inv00 = 1;
    77: op1_06_inv00 = 1;
    58: op1_06_inv00 = 1;
    51: op1_06_inv00 = 1;
    79: op1_06_inv00 = 1;
    28: op1_06_inv00 = 1;
    80: op1_06_inv00 = 1;
    81: op1_06_inv00 = 1;
    63: op1_06_inv00 = 1;
    82: op1_06_inv00 = 1;
    89: op1_06_inv00 = 1;
    47: op1_06_inv00 = 1;
    65: op1_06_inv00 = 1;
    90: op1_06_inv00 = 1;
    91: op1_06_inv00 = 1;
    44: op1_06_inv00 = 1;
    67: op1_06_inv00 = 1;
    94: op1_06_inv00 = 1;
    96: op1_06_inv00 = 1;
    42: op1_06_inv00 = 1;
    98: op1_06_inv00 = 1;
    99: op1_06_inv00 = 1;
    101: op1_06_inv00 = 1;
    102: op1_06_inv00 = 1;
    103: op1_06_inv00 = 1;
    34: op1_06_inv00 = 1;
    106: op1_06_inv00 = 1;
    107: op1_06_inv00 = 1;
    108: op1_06_inv00 = 1;
    109: op1_06_inv00 = 1;
    111: op1_06_inv00 = 1;
    112: op1_06_inv00 = 1;
    113: op1_06_inv00 = 1;
    115: op1_06_inv00 = 1;
    116: op1_06_inv00 = 1;
    38: op1_06_inv00 = 1;
    117: op1_06_inv00 = 1;
    118: op1_06_inv00 = 1;
    119: op1_06_inv00 = 1;
    121: op1_06_inv00 = 1;
    122: op1_06_inv00 = 1;
    123: op1_06_inv00 = 1;
    124: op1_06_inv00 = 1;
    127: op1_06_inv00 = 1;
    129: op1_06_inv00 = 1;
    default: op1_06_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in01 = imem00_in[11:8];
    53: op1_06_in01 = reg_0320;
    114: op1_06_in01 = reg_0320;
    55: op1_06_in01 = reg_0720;
    86: op1_06_in01 = reg_0707;
    73: op1_06_in01 = reg_0040;
    69: op1_06_in01 = reg_0679;
    49: op1_06_in01 = reg_0674;
    71: op1_06_in01 = reg_1279;
    50: op1_06_in01 = reg_0023;
    54: op1_06_in01 = reg_0727;
    74: op1_06_in01 = reg_0614;
    68: op1_06_in01 = reg_0169;
    61: op1_06_in01 = reg_0701;
    75: op1_06_in01 = reg_0121;
    87: op1_06_in01 = reg_0377;
    56: op1_06_in01 = reg_0890;
    76: op1_06_in01 = reg_1241;
    60: op1_06_in01 = reg_0559;
    57: op1_06_in01 = reg_0396;
    77: op1_06_in01 = reg_1278;
    82: op1_06_in01 = reg_1278;
    33: op1_06_in01 = reg_0297;
    70: op1_06_in01 = reg_0742;
    58: op1_06_in01 = reg_1204;
    48: op1_06_in01 = reg_0733;
    78: op1_06_in01 = reg_0906;
    46: op1_06_in01 = reg_0443;
    88: op1_06_in01 = reg_0957;
    51: op1_06_in01 = reg_0298;
    79: op1_06_in01 = reg_1168;
    59: op1_06_in01 = reg_0088;
    80: op1_06_in01 = reg_0341;
    62: op1_06_in01 = reg_0010;
    64: op1_06_in01 = reg_0010;
    52: op1_06_in01 = reg_0871;
    81: op1_06_in01 = reg_0276;
    63: op1_06_in01 = reg_0171;
    89: op1_06_in01 = reg_0185;
    83: op1_06_in01 = reg_0832;
    22: op1_06_in01 = reg_0004;
    37: op1_06_in01 = imem07_in[15:12];
    84: op1_06_in01 = reg_0715;
    47: op1_06_in01 = reg_0223;
    65: op1_06_in01 = reg_0262;
    85: op1_06_in01 = reg_1510;
    91: op1_06_in01 = reg_1510;
    90: op1_06_in01 = reg_0042;
    66: op1_06_in01 = reg_0017;
    44: op1_06_in01 = imem04_in[11:8];
    67: op1_06_in01 = reg_1003;
    92: op1_06_in01 = reg_1071;
    93: op1_06_in01 = reg_0266;
    40: op1_06_in01 = imem07_in[11:8];
    38: op1_06_in01 = imem07_in[11:8];
    94: op1_06_in01 = reg_0025;
    95: op1_06_in01 = imem00_in[3:0];
    107: op1_06_in01 = imem00_in[3:0];
    96: op1_06_in01 = reg_0180;
    42: op1_06_in01 = reg_0747;
    97: op1_06_in01 = reg_0884;
    98: op1_06_in01 = reg_0445;
    99: op1_06_in01 = reg_0672;
    100: op1_06_in01 = reg_0077;
    101: op1_06_in01 = reg_0148;
    102: op1_06_in01 = reg_0333;
    103: op1_06_in01 = reg_1504;
    104: op1_06_in01 = imem00_in[7:4];
    34: op1_06_in01 = reg_0593;
    105: op1_06_in01 = reg_1009;
    106: op1_06_in01 = reg_0216;
    108: op1_06_in01 = reg_1303;
    109: op1_06_in01 = reg_0393;
    110: op1_06_in01 = reg_0433;
    111: op1_06_in01 = reg_0461;
    112: op1_06_in01 = reg_0386;
    113: op1_06_in01 = reg_0860;
    115: op1_06_in01 = imem00_in[15:12];
    116: op1_06_in01 = reg_0934;
    117: op1_06_in01 = reg_0841;
    118: op1_06_in01 = reg_0975;
    119: op1_06_in01 = reg_0728;
    120: op1_06_in01 = reg_0177;
    121: op1_06_in01 = reg_0205;
    122: op1_06_in01 = reg_0601;
    123: op1_06_in01 = reg_1404;
    124: op1_06_in01 = reg_0534;
    125: op1_06_in01 = reg_0879;
    126: op1_06_in01 = reg_0164;
    127: op1_06_in01 = reg_0041;
    128: op1_06_in01 = reg_0634;
    129: op1_06_in01 = reg_0442;
    130: op1_06_in01 = reg_0153;
    131: op1_06_in01 = reg_0418;
    default: op1_06_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv01 = 1;
    53: op1_06_inv01 = 1;
    55: op1_06_inv01 = 1;
    86: op1_06_inv01 = 1;
    73: op1_06_inv01 = 1;
    50: op1_06_inv01 = 1;
    74: op1_06_inv01 = 1;
    87: op1_06_inv01 = 1;
    57: op1_06_inv01 = 1;
    77: op1_06_inv01 = 1;
    48: op1_06_inv01 = 1;
    51: op1_06_inv01 = 1;
    80: op1_06_inv01 = 1;
    62: op1_06_inv01 = 1;
    83: op1_06_inv01 = 1;
    22: op1_06_inv01 = 1;
    37: op1_06_inv01 = 1;
    84: op1_06_inv01 = 1;
    47: op1_06_inv01 = 1;
    85: op1_06_inv01 = 1;
    90: op1_06_inv01 = 1;
    66: op1_06_inv01 = 1;
    91: op1_06_inv01 = 1;
    40: op1_06_inv01 = 1;
    95: op1_06_inv01 = 1;
    96: op1_06_inv01 = 1;
    42: op1_06_inv01 = 1;
    98: op1_06_inv01 = 1;
    100: op1_06_inv01 = 1;
    101: op1_06_inv01 = 1;
    102: op1_06_inv01 = 1;
    103: op1_06_inv01 = 1;
    106: op1_06_inv01 = 1;
    108: op1_06_inv01 = 1;
    109: op1_06_inv01 = 1;
    110: op1_06_inv01 = 1;
    111: op1_06_inv01 = 1;
    114: op1_06_inv01 = 1;
    117: op1_06_inv01 = 1;
    118: op1_06_inv01 = 1;
    120: op1_06_inv01 = 1;
    121: op1_06_inv01 = 1;
    122: op1_06_inv01 = 1;
    126: op1_06_inv01 = 1;
    128: op1_06_inv01 = 1;
    129: op1_06_inv01 = 1;
    130: op1_06_inv01 = 1;
    default: op1_06_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in02 = reg_1470;
    53: op1_06_in02 = reg_0488;
    55: op1_06_in02 = reg_0863;
    86: op1_06_in02 = reg_0989;
    73: op1_06_in02 = reg_1105;
    69: op1_06_in02 = reg_1140;
    49: op1_06_in02 = imem07_in[15:12];
    71: op1_06_in02 = reg_1079;
    98: op1_06_in02 = reg_1079;
    50: op1_06_in02 = reg_0015;
    54: op1_06_in02 = reg_0148;
    74: op1_06_in02 = reg_0748;
    68: op1_06_in02 = reg_0456;
    61: op1_06_in02 = reg_0824;
    75: op1_06_in02 = reg_0805;
    130: op1_06_in02 = reg_0805;
    87: op1_06_in02 = reg_0965;
    56: op1_06_in02 = reg_0168;
    76: op1_06_in02 = reg_0121;
    60: op1_06_in02 = reg_1233;
    57: op1_06_in02 = reg_0860;
    77: op1_06_in02 = reg_1490;
    33: op1_06_in02 = reg_0156;
    70: op1_06_in02 = reg_0744;
    58: op1_06_in02 = reg_0371;
    48: op1_06_in02 = reg_0828;
    78: op1_06_in02 = reg_0870;
    46: op1_06_in02 = reg_0537;
    88: op1_06_in02 = reg_0952;
    51: op1_06_in02 = reg_0299;
    79: op1_06_in02 = reg_0173;
    59: op1_06_in02 = reg_0291;
    80: op1_06_in02 = reg_0462;
    124: op1_06_in02 = reg_0462;
    62: op1_06_in02 = reg_1029;
    52: op1_06_in02 = reg_0868;
    81: op1_06_in02 = reg_0608;
    63: op1_06_in02 = reg_0308;
    82: op1_06_in02 = reg_1487;
    89: op1_06_in02 = reg_0709;
    83: op1_06_in02 = reg_0395;
    64: op1_06_in02 = reg_0457;
    22: op1_06_in02 = reg_0003;
    37: op1_06_in02 = reg_0408;
    84: op1_06_in02 = reg_0401;
    47: op1_06_in02 = reg_0297;
    65: op1_06_in02 = reg_0337;
    85: op1_06_in02 = reg_1281;
    90: op1_06_in02 = reg_0012;
    128: op1_06_in02 = reg_0012;
    66: op1_06_in02 = reg_1055;
    91: op1_06_in02 = reg_1278;
    44: op1_06_in02 = reg_0262;
    67: op1_06_in02 = reg_0597;
    92: op1_06_in02 = imem02_in[3:0];
    93: op1_06_in02 = reg_0367;
    40: op1_06_in02 = reg_0169;
    94: op1_06_in02 = reg_0425;
    95: op1_06_in02 = reg_1279;
    96: op1_06_in02 = reg_1184;
    120: op1_06_in02 = reg_1184;
    42: op1_06_in02 = reg_0742;
    97: op1_06_in02 = reg_0707;
    99: op1_06_in02 = reg_0486;
    100: op1_06_in02 = reg_0079;
    101: op1_06_in02 = reg_0091;
    102: op1_06_in02 = reg_0205;
    103: op1_06_in02 = reg_1179;
    104: op1_06_in02 = reg_0638;
    34: op1_06_in02 = reg_0228;
    105: op1_06_in02 = reg_0426;
    106: op1_06_in02 = reg_0600;
    107: op1_06_in02 = reg_0501;
    108: op1_06_in02 = reg_0295;
    109: op1_06_in02 = reg_0589;
    110: op1_06_in02 = reg_0776;
    111: op1_06_in02 = reg_0298;
    112: op1_06_in02 = reg_0362;
    113: op1_06_in02 = reg_1323;
    114: op1_06_in02 = reg_0342;
    115: op1_06_in02 = reg_1101;
    116: op1_06_in02 = reg_0390;
    38: op1_06_in02 = reg_0030;
    117: op1_06_in02 = reg_0153;
    118: op1_06_in02 = reg_0455;
    119: op1_06_in02 = reg_0042;
    121: op1_06_in02 = reg_1268;
    122: op1_06_in02 = reg_0196;
    123: op1_06_in02 = reg_0939;
    125: op1_06_in02 = reg_0055;
    126: op1_06_in02 = reg_0328;
    127: op1_06_in02 = reg_0011;
    129: op1_06_in02 = reg_0321;
    131: op1_06_in02 = reg_0303;
    default: op1_06_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_06_inv02 = 1;
    73: op1_06_inv02 = 1;
    69: op1_06_inv02 = 1;
    68: op1_06_inv02 = 1;
    75: op1_06_inv02 = 1;
    87: op1_06_inv02 = 1;
    56: op1_06_inv02 = 1;
    76: op1_06_inv02 = 1;
    57: op1_06_inv02 = 1;
    70: op1_06_inv02 = 1;
    78: op1_06_inv02 = 1;
    52: op1_06_inv02 = 1;
    82: op1_06_inv02 = 1;
    22: op1_06_inv02 = 1;
    47: op1_06_inv02 = 1;
    65: op1_06_inv02 = 1;
    66: op1_06_inv02 = 1;
    67: op1_06_inv02 = 1;
    92: op1_06_inv02 = 1;
    93: op1_06_inv02 = 1;
    40: op1_06_inv02 = 1;
    95: op1_06_inv02 = 1;
    42: op1_06_inv02 = 1;
    97: op1_06_inv02 = 1;
    98: op1_06_inv02 = 1;
    99: op1_06_inv02 = 1;
    105: op1_06_inv02 = 1;
    108: op1_06_inv02 = 1;
    109: op1_06_inv02 = 1;
    110: op1_06_inv02 = 1;
    112: op1_06_inv02 = 1;
    115: op1_06_inv02 = 1;
    116: op1_06_inv02 = 1;
    117: op1_06_inv02 = 1;
    119: op1_06_inv02 = 1;
    123: op1_06_inv02 = 1;
    124: op1_06_inv02 = 1;
    126: op1_06_inv02 = 1;
    128: op1_06_inv02 = 1;
    129: op1_06_inv02 = 1;
    130: op1_06_inv02 = 1;
    131: op1_06_inv02 = 1;
    default: op1_06_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in03 = reg_1053;
    53: op1_06_in03 = reg_0340;
    55: op1_06_in03 = reg_0859;
    86: op1_06_in03 = reg_1003;
    73: op1_06_in03 = reg_1437;
    69: op1_06_in03 = reg_0981;
    49: op1_06_in03 = reg_0029;
    71: op1_06_in03 = reg_1081;
    50: op1_06_in03 = reg_0018;
    54: op1_06_in03 = reg_0386;
    74: op1_06_in03 = reg_1079;
    85: op1_06_in03 = reg_1079;
    95: op1_06_in03 = reg_1079;
    68: op1_06_in03 = reg_0561;
    61: op1_06_in03 = reg_1279;
    75: op1_06_in03 = reg_1471;
    87: op1_06_in03 = reg_1517;
    56: op1_06_in03 = reg_0196;
    76: op1_06_in03 = reg_0552;
    60: op1_06_in03 = reg_0145;
    57: op1_06_in03 = reg_0863;
    77: op1_06_in03 = reg_1242;
    33: op1_06_in03 = reg_0140;
    70: op1_06_in03 = reg_0606;
    58: op1_06_in03 = reg_0152;
    48: op1_06_in03 = reg_0175;
    78: op1_06_in03 = reg_0960;
    46: op1_06_in03 = reg_0536;
    88: op1_06_in03 = reg_0220;
    51: op1_06_in03 = reg_0309;
    79: op1_06_in03 = reg_0174;
    59: op1_06_in03 = reg_0277;
    80: op1_06_in03 = reg_1083;
    62: op1_06_in03 = reg_0605;
    52: op1_06_in03 = reg_0874;
    81: op1_06_in03 = reg_0256;
    63: op1_06_in03 = reg_0371;
    82: op1_06_in03 = reg_0805;
    117: op1_06_in03 = reg_0805;
    89: op1_06_in03 = reg_1448;
    83: op1_06_in03 = reg_0347;
    64: op1_06_in03 = reg_0744;
    22: op1_06_in03 = reg_0085;
    37: op1_06_in03 = reg_0413;
    84: op1_06_in03 = reg_0365;
    47: op1_06_in03 = reg_0159;
    65: op1_06_in03 = reg_0097;
    90: op1_06_in03 = reg_0011;
    66: op1_06_in03 = reg_0496;
    91: op1_06_in03 = reg_0153;
    44: op1_06_in03 = reg_0837;
    67: op1_06_in03 = reg_0048;
    92: op1_06_in03 = imem02_in[11:8];
    93: op1_06_in03 = imem05_in[7:4];
    40: op1_06_in03 = reg_0779;
    94: op1_06_in03 = reg_0181;
    96: op1_06_in03 = reg_0246;
    42: op1_06_in03 = reg_0727;
    97: op1_06_in03 = reg_0025;
    98: op1_06_in03 = reg_1487;
    99: op1_06_in03 = reg_0249;
    100: op1_06_in03 = reg_0724;
    101: op1_06_in03 = reg_0724;
    102: op1_06_in03 = reg_0649;
    103: op1_06_in03 = reg_0714;
    104: op1_06_in03 = reg_0501;
    34: op1_06_in03 = reg_0050;
    105: op1_06_in03 = imem04_in[11:8];
    106: op1_06_in03 = reg_0311;
    107: op1_06_in03 = reg_0907;
    108: op1_06_in03 = reg_0165;
    109: op1_06_in03 = reg_1334;
    110: op1_06_in03 = reg_0112;
    111: op1_06_in03 = reg_0703;
    112: op1_06_in03 = reg_0899;
    113: op1_06_in03 = reg_0115;
    114: op1_06_in03 = reg_1419;
    115: op1_06_in03 = reg_0843;
    116: op1_06_in03 = reg_0054;
    38: op1_06_in03 = reg_0661;
    118: op1_06_in03 = reg_1074;
    119: op1_06_in03 = reg_0041;
    120: op1_06_in03 = reg_1313;
    121: op1_06_in03 = reg_0251;
    122: op1_06_in03 = reg_0603;
    123: op1_06_in03 = reg_0792;
    124: op1_06_in03 = reg_1203;
    125: op1_06_in03 = reg_0254;
    126: op1_06_in03 = reg_1147;
    127: op1_06_in03 = imem02_in[15:12];
    128: op1_06_in03 = reg_0662;
    129: op1_06_in03 = reg_0361;
    130: op1_06_in03 = reg_0554;
    131: op1_06_in03 = reg_0873;
    default: op1_06_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv03 = 1;
    53: op1_06_inv03 = 1;
    55: op1_06_inv03 = 1;
    86: op1_06_inv03 = 1;
    54: op1_06_inv03 = 1;
    68: op1_06_inv03 = 1;
    61: op1_06_inv03 = 1;
    75: op1_06_inv03 = 1;
    87: op1_06_inv03 = 1;
    76: op1_06_inv03 = 1;
    77: op1_06_inv03 = 1;
    33: op1_06_inv03 = 1;
    70: op1_06_inv03 = 1;
    58: op1_06_inv03 = 1;
    78: op1_06_inv03 = 1;
    46: op1_06_inv03 = 1;
    80: op1_06_inv03 = 1;
    52: op1_06_inv03 = 1;
    81: op1_06_inv03 = 1;
    63: op1_06_inv03 = 1;
    82: op1_06_inv03 = 1;
    89: op1_06_inv03 = 1;
    64: op1_06_inv03 = 1;
    37: op1_06_inv03 = 1;
    84: op1_06_inv03 = 1;
    65: op1_06_inv03 = 1;
    44: op1_06_inv03 = 1;
    92: op1_06_inv03 = 1;
    40: op1_06_inv03 = 1;
    95: op1_06_inv03 = 1;
    98: op1_06_inv03 = 1;
    99: op1_06_inv03 = 1;
    100: op1_06_inv03 = 1;
    101: op1_06_inv03 = 1;
    104: op1_06_inv03 = 1;
    109: op1_06_inv03 = 1;
    111: op1_06_inv03 = 1;
    112: op1_06_inv03 = 1;
    113: op1_06_inv03 = 1;
    114: op1_06_inv03 = 1;
    115: op1_06_inv03 = 1;
    38: op1_06_inv03 = 1;
    119: op1_06_inv03 = 1;
    120: op1_06_inv03 = 1;
    123: op1_06_inv03 = 1;
    125: op1_06_inv03 = 1;
    126: op1_06_inv03 = 1;
    129: op1_06_inv03 = 1;
    131: op1_06_inv03 = 1;
    default: op1_06_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in04 = reg_1052;
    53: op1_06_in04 = reg_0262;
    55: op1_06_in04 = reg_0373;
    86: op1_06_in04 = reg_0952;
    73: op1_06_in04 = reg_0925;
    69: op1_06_in04 = reg_0256;
    49: op1_06_in04 = reg_0665;
    71: op1_06_in04 = reg_0842;
    50: op1_06_in04 = reg_0457;
    54: op1_06_in04 = reg_0724;
    74: op1_06_in04 = reg_0121;
    68: op1_06_in04 = reg_0560;
    61: op1_06_in04 = reg_1080;
    75: op1_06_in04 = reg_0987;
    87: op1_06_in04 = reg_0190;
    56: op1_06_in04 = reg_0205;
    76: op1_06_in04 = reg_0806;
    104: op1_06_in04 = reg_0806;
    60: op1_06_in04 = reg_0143;
    57: op1_06_in04 = reg_0826;
    77: op1_06_in04 = reg_0552;
    33: op1_06_in04 = reg_0029;
    70: op1_06_in04 = reg_0530;
    58: op1_06_in04 = reg_0212;
    48: op1_06_in04 = reg_0176;
    78: op1_06_in04 = reg_1065;
    46: op1_06_in04 = reg_0493;
    88: op1_06_in04 = reg_0178;
    51: op1_06_in04 = reg_0674;
    79: op1_06_in04 = reg_0567;
    59: op1_06_in04 = reg_0282;
    80: op1_06_in04 = reg_0407;
    62: op1_06_in04 = reg_0607;
    52: op1_06_in04 = reg_0077;
    81: op1_06_in04 = reg_0474;
    63: op1_06_in04 = reg_0046;
    82: op1_06_in04 = reg_1469;
    89: op1_06_in04 = reg_1001;
    83: op1_06_in04 = reg_1259;
    64: op1_06_in04 = imem02_in[15:12];
    22: op1_06_in04 = reg_0052;
    37: op1_06_in04 = reg_0618;
    84: op1_06_in04 = reg_0875;
    47: op1_06_in04 = reg_0157;
    65: op1_06_in04 = reg_0065;
    85: op1_06_in04 = reg_1244;
    90: op1_06_in04 = reg_0590;
    66: op1_06_in04 = reg_0673;
    91: op1_06_in04 = reg_0616;
    44: op1_06_in04 = reg_0096;
    67: op1_06_in04 = reg_0882;
    92: op1_06_in04 = reg_0626;
    93: op1_06_in04 = imem05_in[11:8];
    40: op1_06_in04 = reg_0465;
    94: op1_06_in04 = reg_1367;
    95: op1_06_in04 = reg_0445;
    96: op1_06_in04 = reg_0113;
    42: op1_06_in04 = reg_0451;
    97: op1_06_in04 = reg_1139;
    98: op1_06_in04 = reg_0804;
    99: op1_06_in04 = reg_0229;
    100: op1_06_in04 = reg_0896;
    101: op1_06_in04 = reg_0896;
    102: op1_06_in04 = reg_1180;
    103: op1_06_in04 = reg_0636;
    34: op1_06_in04 = reg_0053;
    105: op1_06_in04 = reg_1144;
    106: op1_06_in04 = reg_0312;
    107: op1_06_in04 = reg_0841;
    108: op1_06_in04 = reg_0195;
    109: op1_06_in04 = reg_1209;
    110: op1_06_in04 = reg_1433;
    111: op1_06_in04 = reg_0158;
    112: op1_06_in04 = reg_0078;
    113: op1_06_in04 = reg_1303;
    114: op1_06_in04 = reg_0487;
    115: op1_06_in04 = reg_1277;
    116: op1_06_in04 = reg_0776;
    38: op1_06_in04 = reg_0740;
    117: op1_06_in04 = reg_0486;
    118: op1_06_in04 = reg_0126;
    119: op1_06_in04 = reg_0012;
    120: op1_06_in04 = reg_1208;
    121: op1_06_in04 = reg_0174;
    122: op1_06_in04 = reg_0449;
    123: op1_06_in04 = reg_0303;
    124: op1_06_in04 = reg_1215;
    125: op1_06_in04 = reg_0712;
    126: op1_06_in04 = reg_0406;
    127: op1_06_in04 = reg_0495;
    128: op1_06_in04 = imem02_in[11:8];
    129: op1_06_in04 = reg_0998;
    130: op1_06_in04 = reg_0555;
    131: op1_06_in04 = reg_0066;
    default: op1_06_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_06_inv04 = 1;
    55: op1_06_inv04 = 1;
    86: op1_06_inv04 = 1;
    73: op1_06_inv04 = 1;
    50: op1_06_inv04 = 1;
    54: op1_06_inv04 = 1;
    74: op1_06_inv04 = 1;
    68: op1_06_inv04 = 1;
    61: op1_06_inv04 = 1;
    75: op1_06_inv04 = 1;
    56: op1_06_inv04 = 1;
    77: op1_06_inv04 = 1;
    33: op1_06_inv04 = 1;
    70: op1_06_inv04 = 1;
    46: op1_06_inv04 = 1;
    79: op1_06_inv04 = 1;
    59: op1_06_inv04 = 1;
    80: op1_06_inv04 = 1;
    52: op1_06_inv04 = 1;
    63: op1_06_inv04 = 1;
    89: op1_06_inv04 = 1;
    83: op1_06_inv04 = 1;
    64: op1_06_inv04 = 1;
    22: op1_06_inv04 = 1;
    84: op1_06_inv04 = 1;
    65: op1_06_inv04 = 1;
    85: op1_06_inv04 = 1;
    90: op1_06_inv04 = 1;
    66: op1_06_inv04 = 1;
    91: op1_06_inv04 = 1;
    44: op1_06_inv04 = 1;
    42: op1_06_inv04 = 1;
    97: op1_06_inv04 = 1;
    99: op1_06_inv04 = 1;
    100: op1_06_inv04 = 1;
    102: op1_06_inv04 = 1;
    105: op1_06_inv04 = 1;
    107: op1_06_inv04 = 1;
    109: op1_06_inv04 = 1;
    110: op1_06_inv04 = 1;
    112: op1_06_inv04 = 1;
    113: op1_06_inv04 = 1;
    114: op1_06_inv04 = 1;
    116: op1_06_inv04 = 1;
    117: op1_06_inv04 = 1;
    120: op1_06_inv04 = 1;
    121: op1_06_inv04 = 1;
    122: op1_06_inv04 = 1;
    124: op1_06_inv04 = 1;
    125: op1_06_inv04 = 1;
    127: op1_06_inv04 = 1;
    128: op1_06_inv04 = 1;
    129: op1_06_inv04 = 1;
    130: op1_06_inv04 = 1;
    default: op1_06_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in05 = reg_1028;
    117: op1_06_in05 = reg_1028;
    53: op1_06_in05 = reg_0862;
    55: op1_06_in05 = reg_0374;
    86: op1_06_in05 = reg_0329;
    73: op1_06_in05 = reg_0536;
    69: op1_06_in05 = reg_0473;
    49: op1_06_in05 = reg_0663;
    71: op1_06_in05 = imem00_in[3:0];
    50: op1_06_in05 = imem07_in[3:0];
    54: op1_06_in05 = reg_0079;
    74: op1_06_in05 = reg_0804;
    104: op1_06_in05 = reg_0804;
    68: op1_06_in05 = reg_0255;
    61: op1_06_in05 = reg_0842;
    75: op1_06_in05 = reg_1206;
    87: op1_06_in05 = reg_0246;
    56: op1_06_in05 = reg_0039;
    76: op1_06_in05 = reg_0803;
    60: op1_06_in05 = reg_1208;
    57: op1_06_in05 = reg_0825;
    77: op1_06_in05 = reg_1053;
    130: op1_06_in05 = reg_1053;
    33: op1_06_in05 = reg_0030;
    70: op1_06_in05 = reg_0590;
    58: op1_06_in05 = reg_1150;
    48: op1_06_in05 = imem05_in[11:8];
    78: op1_06_in05 = reg_0109;
    46: op1_06_in05 = reg_0681;
    88: op1_06_in05 = reg_0108;
    51: op1_06_in05 = reg_0159;
    79: op1_06_in05 = reg_0566;
    59: op1_06_in05 = reg_0699;
    80: op1_06_in05 = reg_0094;
    62: op1_06_in05 = reg_0588;
    52: op1_06_in05 = reg_0222;
    81: op1_06_in05 = reg_0494;
    63: op1_06_in05 = reg_0015;
    82: op1_06_in05 = reg_0293;
    89: op1_06_in05 = reg_0144;
    83: op1_06_in05 = reg_1169;
    64: op1_06_in05 = reg_0981;
    37: op1_06_in05 = reg_0593;
    84: op1_06_in05 = reg_0595;
    47: op1_06_in05 = reg_0139;
    65: op1_06_in05 = reg_0209;
    85: op1_06_in05 = reg_0615;
    90: op1_06_in05 = reg_0666;
    66: op1_06_in05 = reg_1351;
    91: op1_06_in05 = reg_0186;
    115: op1_06_in05 = reg_0186;
    44: op1_06_in05 = reg_0237;
    67: op1_06_in05 = reg_0884;
    120: op1_06_in05 = reg_0884;
    92: op1_06_in05 = reg_0253;
    93: op1_06_in05 = reg_0702;
    40: op1_06_in05 = reg_0661;
    94: op1_06_in05 = reg_1083;
    95: op1_06_in05 = reg_1487;
    96: op1_06_in05 = reg_0707;
    42: op1_06_in05 = reg_0160;
    97: op1_06_in05 = reg_0443;
    98: op1_06_in05 = reg_0555;
    99: op1_06_in05 = reg_1417;
    100: op1_06_in05 = reg_0162;
    101: op1_06_in05 = reg_0042;
    102: op1_06_in05 = reg_1401;
    103: op1_06_in05 = reg_0398;
    34: op1_06_in05 = reg_0519;
    105: op1_06_in05 = reg_0208;
    106: op1_06_in05 = reg_0143;
    107: op1_06_in05 = reg_0580;
    108: op1_06_in05 = reg_0212;
    109: op1_06_in05 = reg_1179;
    110: op1_06_in05 = reg_0307;
    111: op1_06_in05 = reg_0664;
    112: op1_06_in05 = reg_0012;
    113: op1_06_in05 = reg_0636;
    114: op1_06_in05 = reg_0096;
    116: op1_06_in05 = reg_1455;
    38: op1_06_in05 = reg_0623;
    118: op1_06_in05 = reg_0111;
    119: op1_06_in05 = reg_0662;
    121: op1_06_in05 = reg_0173;
    122: op1_06_in05 = reg_0317;
    123: op1_06_in05 = reg_0301;
    124: op1_06_in05 = reg_1041;
    125: op1_06_in05 = reg_1493;
    126: op1_06_in05 = reg_0969;
    127: op1_06_in05 = reg_1235;
    128: op1_06_in05 = reg_0495;
    129: op1_06_in05 = reg_0052;
    131: op1_06_in05 = reg_0575;
    default: op1_06_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv05 = 1;
    53: op1_06_inv05 = 1;
    55: op1_06_inv05 = 1;
    73: op1_06_inv05 = 1;
    69: op1_06_inv05 = 1;
    49: op1_06_inv05 = 1;
    74: op1_06_inv05 = 1;
    68: op1_06_inv05 = 1;
    61: op1_06_inv05 = 1;
    60: op1_06_inv05 = 1;
    57: op1_06_inv05 = 1;
    77: op1_06_inv05 = 1;
    58: op1_06_inv05 = 1;
    48: op1_06_inv05 = 1;
    78: op1_06_inv05 = 1;
    46: op1_06_inv05 = 1;
    88: op1_06_inv05 = 1;
    79: op1_06_inv05 = 1;
    81: op1_06_inv05 = 1;
    89: op1_06_inv05 = 1;
    64: op1_06_inv05 = 1;
    84: op1_06_inv05 = 1;
    47: op1_06_inv05 = 1;
    65: op1_06_inv05 = 1;
    90: op1_06_inv05 = 1;
    66: op1_06_inv05 = 1;
    44: op1_06_inv05 = 1;
    67: op1_06_inv05 = 1;
    97: op1_06_inv05 = 1;
    100: op1_06_inv05 = 1;
    102: op1_06_inv05 = 1;
    34: op1_06_inv05 = 1;
    105: op1_06_inv05 = 1;
    106: op1_06_inv05 = 1;
    111: op1_06_inv05 = 1;
    112: op1_06_inv05 = 1;
    115: op1_06_inv05 = 1;
    116: op1_06_inv05 = 1;
    119: op1_06_inv05 = 1;
    120: op1_06_inv05 = 1;
    124: op1_06_inv05 = 1;
    125: op1_06_inv05 = 1;
    127: op1_06_inv05 = 1;
    default: op1_06_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in06 = reg_1454;
    53: op1_06_in06 = reg_0836;
    55: op1_06_in06 = reg_0822;
    86: op1_06_in06 = reg_1301;
    87: op1_06_in06 = reg_1301;
    73: op1_06_in06 = reg_0720;
    69: op1_06_in06 = reg_1207;
    49: op1_06_in06 = reg_0286;
    33: op1_06_in06 = reg_0286;
    71: op1_06_in06 = imem00_in[15:12];
    50: op1_06_in06 = reg_0995;
    54: op1_06_in06 = reg_0282;
    74: op1_06_in06 = reg_0803;
    61: op1_06_in06 = reg_0803;
    68: op1_06_in06 = reg_0128;
    75: op1_06_in06 = reg_0961;
    117: op1_06_in06 = reg_0961;
    56: op1_06_in06 = reg_1036;
    76: op1_06_in06 = reg_1052;
    60: op1_06_in06 = reg_0884;
    57: op1_06_in06 = reg_0116;
    77: op1_06_in06 = reg_0523;
    70: op1_06_in06 = reg_0255;
    58: op1_06_in06 = reg_0491;
    48: op1_06_in06 = reg_0648;
    78: op1_06_in06 = reg_0717;
    46: op1_06_in06 = reg_0552;
    88: op1_06_in06 = reg_0882;
    51: op1_06_in06 = reg_0923;
    79: op1_06_in06 = reg_0045;
    59: op1_06_in06 = reg_1103;
    80: op1_06_in06 = reg_0837;
    62: op1_06_in06 = reg_0587;
    52: op1_06_in06 = reg_0667;
    81: op1_06_in06 = reg_0970;
    63: op1_06_in06 = reg_0821;
    82: op1_06_in06 = reg_1227;
    89: op1_06_in06 = reg_0349;
    83: op1_06_in06 = reg_1104;
    64: op1_06_in06 = reg_0256;
    37: op1_06_in06 = reg_0137;
    84: op1_06_in06 = reg_0077;
    47: op1_06_in06 = reg_0777;
    65: op1_06_in06 = reg_0016;
    85: op1_06_in06 = reg_0804;
    90: op1_06_in06 = reg_0456;
    66: op1_06_in06 = reg_0703;
    91: op1_06_in06 = reg_0640;
    98: op1_06_in06 = reg_0640;
    44: op1_06_in06 = reg_0181;
    105: op1_06_in06 = reg_0181;
    67: op1_06_in06 = reg_0504;
    92: op1_06_in06 = reg_0588;
    93: op1_06_in06 = reg_0466;
    40: op1_06_in06 = reg_0739;
    94: op1_06_in06 = reg_1214;
    95: op1_06_in06 = reg_0806;
    96: op1_06_in06 = reg_0378;
    42: op1_06_in06 = reg_0163;
    97: op1_06_in06 = reg_1146;
    99: op1_06_in06 = reg_0155;
    100: op1_06_in06 = reg_1068;
    101: op1_06_in06 = reg_1068;
    102: op1_06_in06 = reg_0939;
    103: op1_06_in06 = reg_0617;
    104: op1_06_in06 = reg_0841;
    106: op1_06_in06 = reg_1184;
    107: op1_06_in06 = reg_0186;
    108: op1_06_in06 = reg_0018;
    109: op1_06_in06 = reg_0110;
    110: op1_06_in06 = reg_0473;
    111: op1_06_in06 = reg_0740;
    112: op1_06_in06 = reg_0662;
    113: op1_06_in06 = reg_0637;
    114: op1_06_in06 = reg_1189;
    115: op1_06_in06 = reg_0555;
    116: op1_06_in06 = reg_1140;
    38: op1_06_in06 = reg_0618;
    118: op1_06_in06 = reg_0105;
    119: op1_06_in06 = imem02_in[11:8];
    120: op1_06_in06 = reg_1144;
    121: op1_06_in06 = reg_0697;
    122: op1_06_in06 = reg_0206;
    123: op1_06_in06 = reg_0450;
    124: op1_06_in06 = reg_1040;
    125: op1_06_in06 = reg_0054;
    126: op1_06_in06 = reg_0199;
    127: op1_06_in06 = reg_0276;
    128: op1_06_in06 = reg_0008;
    129: op1_06_in06 = reg_0086;
    130: op1_06_in06 = reg_0293;
    131: op1_06_in06 = reg_0151;
    default: op1_06_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv06 = 1;
    49: op1_06_inv06 = 1;
    50: op1_06_inv06 = 1;
    74: op1_06_inv06 = 1;
    75: op1_06_inv06 = 1;
    56: op1_06_inv06 = 1;
    60: op1_06_inv06 = 1;
    77: op1_06_inv06 = 1;
    33: op1_06_inv06 = 1;
    70: op1_06_inv06 = 1;
    58: op1_06_inv06 = 1;
    48: op1_06_inv06 = 1;
    88: op1_06_inv06 = 1;
    79: op1_06_inv06 = 1;
    59: op1_06_inv06 = 1;
    80: op1_06_inv06 = 1;
    62: op1_06_inv06 = 1;
    52: op1_06_inv06 = 1;
    82: op1_06_inv06 = 1;
    64: op1_06_inv06 = 1;
    47: op1_06_inv06 = 1;
    65: op1_06_inv06 = 1;
    85: op1_06_inv06 = 1;
    90: op1_06_inv06 = 1;
    66: op1_06_inv06 = 1;
    95: op1_06_inv06 = 1;
    96: op1_06_inv06 = 1;
    42: op1_06_inv06 = 1;
    97: op1_06_inv06 = 1;
    98: op1_06_inv06 = 1;
    101: op1_06_inv06 = 1;
    103: op1_06_inv06 = 1;
    105: op1_06_inv06 = 1;
    107: op1_06_inv06 = 1;
    108: op1_06_inv06 = 1;
    110: op1_06_inv06 = 1;
    120: op1_06_inv06 = 1;
    123: op1_06_inv06 = 1;
    125: op1_06_inv06 = 1;
    126: op1_06_inv06 = 1;
    127: op1_06_inv06 = 1;
    128: op1_06_inv06 = 1;
    129: op1_06_inv06 = 1;
    130: op1_06_inv06 = 1;
    131: op1_06_inv06 = 1;
    default: op1_06_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in07 = reg_1453;
    130: op1_06_in07 = reg_1453;
    53: op1_06_in07 = reg_0237;
    55: op1_06_in07 = reg_0718;
    86: op1_06_in07 = reg_0108;
    73: op1_06_in07 = imem06_in[3:0];
    69: op1_06_in07 = reg_0626;
    49: op1_06_in07 = reg_0441;
    71: op1_06_in07 = reg_0221;
    77: op1_06_in07 = reg_0221;
    50: op1_06_in07 = reg_0223;
    54: op1_06_in07 = reg_0044;
    74: op1_06_in07 = reg_1053;
    98: op1_06_in07 = reg_1053;
    68: op1_06_in07 = reg_0125;
    61: op1_06_in07 = reg_0249;
    75: op1_06_in07 = reg_0524;
    87: op1_06_in07 = reg_1226;
    56: op1_06_in07 = reg_0753;
    76: op1_06_in07 = reg_1028;
    60: op1_06_in07 = reg_0478;
    57: op1_06_in07 = reg_0671;
    33: op1_06_in07 = reg_0437;
    70: op1_06_in07 = reg_0631;
    58: op1_06_in07 = imem07_in[7:4];
    48: op1_06_in07 = reg_0992;
    78: op1_06_in07 = reg_1302;
    46: op1_06_in07 = reg_0467;
    88: op1_06_in07 = reg_0458;
    51: op1_06_in07 = reg_0029;
    79: op1_06_in07 = reg_1181;
    59: op1_06_in07 = reg_0975;
    80: op1_06_in07 = reg_0337;
    62: op1_06_in07 = reg_1140;
    52: op1_06_in07 = imem02_in[3:0];
    81: op1_06_in07 = reg_1455;
    63: op1_06_in07 = reg_1055;
    82: op1_06_in07 = reg_1230;
    89: op1_06_in07 = reg_0954;
    83: op1_06_in07 = reg_0566;
    64: op1_06_in07 = reg_0473;
    37: op1_06_in07 = reg_0103;
    84: op1_06_in07 = reg_0079;
    47: op1_06_in07 = reg_0661;
    65: op1_06_in07 = reg_0750;
    85: op1_06_in07 = reg_1471;
    90: op1_06_in07 = reg_1018;
    112: op1_06_in07 = reg_1018;
    66: op1_06_in07 = reg_0140;
    91: op1_06_in07 = reg_0293;
    44: op1_06_in07 = reg_0117;
    67: op1_06_in07 = reg_0840;
    92: op1_06_in07 = reg_0532;
    93: op1_06_in07 = reg_0184;
    40: op1_06_in07 = reg_0623;
    94: op1_06_in07 = reg_1082;
    95: op1_06_in07 = reg_0613;
    96: op1_06_in07 = reg_0541;
    42: op1_06_in07 = reg_0146;
    97: op1_06_in07 = reg_1383;
    99: op1_06_in07 = reg_0883;
    100: op1_06_in07 = reg_0662;
    101: op1_06_in07 = reg_0322;
    102: op1_06_in07 = reg_0937;
    103: op1_06_in07 = reg_0528;
    104: op1_06_in07 = reg_0153;
    105: op1_06_in07 = reg_0493;
    106: op1_06_in07 = reg_1517;
    107: op1_06_in07 = reg_1227;
    108: op1_06_in07 = imem07_in[3:0];
    109: op1_06_in07 = reg_0716;
    110: op1_06_in07 = reg_0829;
    111: op1_06_in07 = reg_0102;
    113: op1_06_in07 = reg_0374;
    114: op1_06_in07 = reg_0211;
    115: op1_06_in07 = reg_0640;
    116: op1_06_in07 = reg_0628;
    38: op1_06_in07 = reg_0591;
    117: op1_06_in07 = reg_0459;
    118: op1_06_in07 = reg_0382;
    119: op1_06_in07 = reg_0659;
    120: op1_06_in07 = reg_1257;
    121: op1_06_in07 = reg_1401;
    122: op1_06_in07 = reg_0461;
    123: op1_06_in07 = reg_0601;
    124: op1_06_in07 = reg_0232;
    125: op1_06_in07 = reg_0971;
    126: op1_06_in07 = reg_0454;
    127: op1_06_in07 = reg_0839;
    128: op1_06_in07 = reg_0666;
    129: op1_06_in07 = reg_0483;
    131: op1_06_in07 = reg_0014;
    default: op1_06_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_06_inv07 = 1;
    54: op1_06_inv07 = 1;
    68: op1_06_inv07 = 1;
    75: op1_06_inv07 = 1;
    57: op1_06_inv07 = 1;
    77: op1_06_inv07 = 1;
    48: op1_06_inv07 = 1;
    78: op1_06_inv07 = 1;
    46: op1_06_inv07 = 1;
    88: op1_06_inv07 = 1;
    51: op1_06_inv07 = 1;
    82: op1_06_inv07 = 1;
    89: op1_06_inv07 = 1;
    37: op1_06_inv07 = 1;
    84: op1_06_inv07 = 1;
    65: op1_06_inv07 = 1;
    44: op1_06_inv07 = 1;
    67: op1_06_inv07 = 1;
    92: op1_06_inv07 = 1;
    93: op1_06_inv07 = 1;
    95: op1_06_inv07 = 1;
    42: op1_06_inv07 = 1;
    98: op1_06_inv07 = 1;
    101: op1_06_inv07 = 1;
    103: op1_06_inv07 = 1;
    104: op1_06_inv07 = 1;
    105: op1_06_inv07 = 1;
    106: op1_06_inv07 = 1;
    107: op1_06_inv07 = 1;
    108: op1_06_inv07 = 1;
    109: op1_06_inv07 = 1;
    110: op1_06_inv07 = 1;
    112: op1_06_inv07 = 1;
    114: op1_06_inv07 = 1;
    117: op1_06_inv07 = 1;
    120: op1_06_inv07 = 1;
    121: op1_06_inv07 = 1;
    122: op1_06_inv07 = 1;
    125: op1_06_inv07 = 1;
    127: op1_06_inv07 = 1;
    128: op1_06_inv07 = 1;
    129: op1_06_inv07 = 1;
    130: op1_06_inv07 = 1;
    default: op1_06_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in08 = reg_0476;
    53: op1_06_in08 = reg_0210;
    55: op1_06_in08 = reg_0669;
    86: op1_06_in08 = imem03_in[3:0];
    73: op1_06_in08 = imem06_in[11:8];
    122: op1_06_in08 = imem06_in[11:8];
    69: op1_06_in08 = reg_0933;
    49: op1_06_in08 = reg_0618;
    71: op1_06_in08 = reg_1453;
    50: op1_06_in08 = reg_0224;
    54: op1_06_in08 = reg_0011;
    74: op1_06_in08 = reg_1201;
    68: op1_06_in08 = reg_0055;
    61: op1_06_in08 = reg_1230;
    75: op1_06_in08 = reg_0928;
    87: op1_06_in08 = reg_0880;
    56: op1_06_in08 = reg_0752;
    76: op1_06_in08 = reg_1027;
    60: op1_06_in08 = reg_0425;
    57: op1_06_in08 = reg_0637;
    77: op1_06_in08 = reg_0485;
    33: op1_06_in08 = imem07_in[3:0];
    70: op1_06_in08 = reg_0474;
    58: op1_06_in08 = imem07_in[15:12];
    108: op1_06_in08 = imem07_in[15:12];
    48: op1_06_in08 = reg_0565;
    78: op1_06_in08 = reg_0570;
    103: op1_06_in08 = reg_0570;
    46: op1_06_in08 = reg_0421;
    88: op1_06_in08 = reg_0218;
    51: op1_06_in08 = reg_0661;
    79: op1_06_in08 = reg_1403;
    59: op1_06_in08 = reg_0922;
    80: op1_06_in08 = reg_0336;
    62: op1_06_in08 = reg_0497;
    52: op1_06_in08 = reg_0563;
    81: op1_06_in08 = reg_0496;
    63: op1_06_in08 = reg_0998;
    82: op1_06_in08 = reg_1229;
    130: op1_06_in08 = reg_1229;
    89: op1_06_in08 = reg_0957;
    83: op1_06_in08 = reg_0630;
    64: op1_06_in08 = reg_0475;
    37: op1_06_in08 = reg_0100;
    38: op1_06_in08 = reg_0100;
    84: op1_06_in08 = reg_0088;
    47: op1_06_in08 = reg_0285;
    65: op1_06_in08 = reg_0251;
    85: op1_06_in08 = reg_1470;
    90: op1_06_in08 = reg_0495;
    66: op1_06_in08 = reg_0156;
    91: op1_06_in08 = reg_0221;
    98: op1_06_in08 = reg_0221;
    44: op1_06_in08 = reg_0129;
    67: op1_06_in08 = reg_0330;
    92: op1_06_in08 = reg_0776;
    93: op1_06_in08 = reg_1268;
    40: op1_06_in08 = reg_0621;
    94: op1_06_in08 = reg_1147;
    95: op1_06_in08 = reg_0486;
    104: op1_06_in08 = reg_0486;
    96: op1_06_in08 = reg_1009;
    42: op1_06_in08 = reg_0402;
    97: op1_06_in08 = reg_1368;
    99: op1_06_in08 = reg_0352;
    100: op1_06_in08 = reg_0590;
    101: op1_06_in08 = reg_0533;
    102: op1_06_in08 = reg_0303;
    105: op1_06_in08 = reg_1257;
    106: op1_06_in08 = reg_0246;
    107: op1_06_in08 = reg_1205;
    109: op1_06_in08 = reg_0586;
    110: op1_06_in08 = reg_0745;
    111: op1_06_in08 = reg_0028;
    112: op1_06_in08 = reg_0588;
    113: op1_06_in08 = reg_0619;
    114: op1_06_in08 = reg_0470;
    115: op1_06_in08 = reg_1052;
    116: op1_06_in08 = reg_0876;
    117: op1_06_in08 = reg_0524;
    118: op1_06_in08 = reg_0631;
    119: op1_06_in08 = reg_0184;
    120: op1_06_in08 = reg_0094;
    121: op1_06_in08 = reg_0477;
    123: op1_06_in08 = reg_0274;
    124: op1_06_in08 = reg_1143;
    125: op1_06_in08 = reg_0127;
    126: op1_06_in08 = reg_0033;
    127: op1_06_in08 = reg_0900;
    128: op1_06_in08 = reg_0879;
    129: op1_06_in08 = reg_1182;
    131: op1_06_in08 = imem06_in[3:0];
    default: op1_06_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv08 = 1;
    55: op1_06_inv08 = 1;
    49: op1_06_inv08 = 1;
    61: op1_06_inv08 = 1;
    76: op1_06_inv08 = 1;
    46: op1_06_inv08 = 1;
    59: op1_06_inv08 = 1;
    80: op1_06_inv08 = 1;
    81: op1_06_inv08 = 1;
    63: op1_06_inv08 = 1;
    89: op1_06_inv08 = 1;
    65: op1_06_inv08 = 1;
    85: op1_06_inv08 = 1;
    66: op1_06_inv08 = 1;
    67: op1_06_inv08 = 1;
    93: op1_06_inv08 = 1;
    96: op1_06_inv08 = 1;
    42: op1_06_inv08 = 1;
    98: op1_06_inv08 = 1;
    100: op1_06_inv08 = 1;
    101: op1_06_inv08 = 1;
    104: op1_06_inv08 = 1;
    106: op1_06_inv08 = 1;
    109: op1_06_inv08 = 1;
    111: op1_06_inv08 = 1;
    113: op1_06_inv08 = 1;
    114: op1_06_inv08 = 1;
    116: op1_06_inv08 = 1;
    38: op1_06_inv08 = 1;
    120: op1_06_inv08 = 1;
    121: op1_06_inv08 = 1;
    124: op1_06_inv08 = 1;
    126: op1_06_inv08 = 1;
    129: op1_06_inv08 = 1;
    130: op1_06_inv08 = 1;
    default: op1_06_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in09 = reg_0928;
    53: op1_06_in09 = reg_0209;
    55: op1_06_in09 = reg_0636;
    86: op1_06_in09 = imem03_in[7:4];
    87: op1_06_in09 = imem03_in[7:4];
    73: op1_06_in09 = reg_0110;
    69: op1_06_in09 = reg_0712;
    68: op1_06_in09 = reg_0712;
    49: op1_06_in09 = reg_0103;
    71: op1_06_in09 = reg_0459;
    50: op1_06_in09 = reg_0309;
    54: op1_06_in09 = imem02_in[3:0];
    74: op1_06_in09 = reg_0961;
    61: op1_06_in09 = reg_1229;
    75: op1_06_in09 = reg_0202;
    56: op1_06_in09 = reg_1058;
    76: op1_06_in09 = reg_0485;
    60: op1_06_in09 = reg_0582;
    57: op1_06_in09 = reg_0295;
    77: op1_06_in09 = reg_1227;
    33: op1_06_in09 = reg_0591;
    70: op1_06_in09 = reg_0432;
    58: op1_06_in09 = reg_0461;
    48: op1_06_in09 = reg_0066;
    78: op1_06_in09 = reg_0132;
    103: op1_06_in09 = reg_0132;
    46: op1_06_in09 = imem04_in[7:4];
    88: op1_06_in09 = reg_0426;
    51: op1_06_in09 = reg_0285;
    79: op1_06_in09 = reg_0940;
    59: op1_06_in09 = reg_0976;
    80: op1_06_in09 = reg_0211;
    62: op1_06_in09 = imem02_in[15:12];
    52: op1_06_in09 = reg_0560;
    110: op1_06_in09 = reg_0560;
    81: op1_06_in09 = reg_0878;
    63: op1_06_in09 = reg_0496;
    82: op1_06_in09 = reg_1417;
    89: op1_06_in09 = reg_0220;
    83: op1_06_in09 = reg_1181;
    64: op1_06_in09 = reg_0494;
    37: op1_06_in09 = reg_0050;
    84: op1_06_in09 = reg_0044;
    47: op1_06_in09 = reg_0441;
    65: op1_06_in09 = reg_0737;
    85: op1_06_in09 = reg_0523;
    90: op1_06_in09 = reg_1207;
    66: op1_06_in09 = reg_0921;
    91: op1_06_in09 = reg_1454;
    44: op1_06_in09 = reg_0575;
    67: op1_06_in09 = reg_1312;
    92: op1_06_in09 = reg_0380;
    93: op1_06_in09 = reg_0604;
    40: op1_06_in09 = reg_0618;
    94: op1_06_in09 = reg_0414;
    95: op1_06_in09 = reg_0293;
    96: op1_06_in09 = reg_0313;
    42: op1_06_in09 = reg_0384;
    97: op1_06_in09 = reg_0264;
    98: op1_06_in09 = reg_1459;
    99: op1_06_in09 = reg_0428;
    100: op1_06_in09 = reg_0845;
    101: op1_06_in09 = reg_0475;
    102: op1_06_in09 = reg_0872;
    104: op1_06_in09 = reg_0250;
    105: op1_06_in09 = reg_0978;
    106: op1_06_in09 = reg_0884;
    107: op1_06_in09 = reg_0476;
    108: op1_06_in09 = reg_0963;
    109: op1_06_in09 = reg_0979;
    111: op1_06_in09 = reg_0228;
    112: op1_06_in09 = reg_0822;
    113: op1_06_in09 = reg_0624;
    114: op1_06_in09 = reg_0038;
    115: op1_06_in09 = reg_0221;
    116: op1_06_in09 = reg_0381;
    127: op1_06_in09 = reg_0381;
    38: op1_06_in09 = reg_0001;
    117: op1_06_in09 = reg_0821;
    118: op1_06_in09 = reg_0473;
    119: op1_06_in09 = reg_0877;
    120: op1_06_in09 = reg_0421;
    121: op1_06_in09 = reg_0937;
    122: op1_06_in09 = reg_0397;
    123: op1_06_in09 = reg_0240;
    124: op1_06_in09 = reg_0062;
    125: op1_06_in09 = reg_0125;
    126: op1_06_in09 = reg_0698;
    128: op1_06_in09 = reg_0138;
    130: op1_06_in09 = reg_0987;
    131: op1_06_in09 = reg_0289;
    default: op1_06_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_06_inv09 = 1;
    69: op1_06_inv09 = 1;
    49: op1_06_inv09 = 1;
    54: op1_06_inv09 = 1;
    74: op1_06_inv09 = 1;
    68: op1_06_inv09 = 1;
    61: op1_06_inv09 = 1;
    75: op1_06_inv09 = 1;
    60: op1_06_inv09 = 1;
    57: op1_06_inv09 = 1;
    70: op1_06_inv09 = 1;
    78: op1_06_inv09 = 1;
    46: op1_06_inv09 = 1;
    88: op1_06_inv09 = 1;
    51: op1_06_inv09 = 1;
    79: op1_06_inv09 = 1;
    62: op1_06_inv09 = 1;
    52: op1_06_inv09 = 1;
    81: op1_06_inv09 = 1;
    89: op1_06_inv09 = 1;
    47: op1_06_inv09 = 1;
    90: op1_06_inv09 = 1;
    66: op1_06_inv09 = 1;
    44: op1_06_inv09 = 1;
    67: op1_06_inv09 = 1;
    93: op1_06_inv09 = 1;
    40: op1_06_inv09 = 1;
    94: op1_06_inv09 = 1;
    95: op1_06_inv09 = 1;
    42: op1_06_inv09 = 1;
    97: op1_06_inv09 = 1;
    98: op1_06_inv09 = 1;
    99: op1_06_inv09 = 1;
    100: op1_06_inv09 = 1;
    102: op1_06_inv09 = 1;
    104: op1_06_inv09 = 1;
    109: op1_06_inv09 = 1;
    112: op1_06_inv09 = 1;
    113: op1_06_inv09 = 1;
    115: op1_06_inv09 = 1;
    116: op1_06_inv09 = 1;
    38: op1_06_inv09 = 1;
    117: op1_06_inv09 = 1;
    118: op1_06_inv09 = 1;
    119: op1_06_inv09 = 1;
    121: op1_06_inv09 = 1;
    126: op1_06_inv09 = 1;
    127: op1_06_inv09 = 1;
    128: op1_06_inv09 = 1;
    131: op1_06_inv09 = 1;
    default: op1_06_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in10 = reg_0188;
    82: op1_06_in10 = reg_0188;
    53: op1_06_in10 = reg_0208;
    55: op1_06_in10 = reg_0264;
    86: op1_06_in10 = imem03_in[11:8];
    73: op1_06_in10 = reg_0717;
    69: op1_06_in10 = reg_0705;
    49: op1_06_in10 = reg_0050;
    71: op1_06_in10 = reg_0928;
    115: op1_06_in10 = reg_0928;
    50: op1_06_in10 = reg_0159;
    54: op1_06_in10 = reg_1098;
    92: op1_06_in10 = reg_1098;
    74: op1_06_in10 = reg_1417;
    76: op1_06_in10 = reg_1417;
    68: op1_06_in10 = reg_0708;
    61: op1_06_in10 = reg_0959;
    75: op1_06_in10 = reg_0351;
    87: op1_06_in10 = reg_0480;
    89: op1_06_in10 = reg_0480;
    56: op1_06_in10 = reg_0863;
    60: op1_06_in10 = imem04_in[11:8];
    57: op1_06_in10 = reg_1179;
    77: op1_06_in10 = reg_0961;
    33: op1_06_in10 = reg_0100;
    70: op1_06_in10 = reg_0778;
    58: op1_06_in10 = reg_0703;
    48: op1_06_in10 = reg_0045;
    78: op1_06_in10 = reg_0308;
    46: op1_06_in10 = reg_0798;
    88: op1_06_in10 = reg_0534;
    67: op1_06_in10 = reg_0534;
    51: op1_06_in10 = reg_0441;
    79: op1_06_in10 = reg_1514;
    59: op1_06_in10 = reg_0456;
    80: op1_06_in10 = reg_1502;
    62: op1_06_in10 = reg_0472;
    52: op1_06_in10 = reg_0495;
    81: op1_06_in10 = reg_0307;
    63: op1_06_in10 = reg_0673;
    96: op1_06_in10 = reg_0673;
    83: op1_06_in10 = reg_1404;
    64: op1_06_in10 = reg_0433;
    37: op1_06_in10 = reg_0521;
    84: op1_06_in10 = reg_0846;
    100: op1_06_in10 = reg_0846;
    47: op1_06_in10 = reg_0740;
    65: op1_06_in10 = reg_0735;
    85: op1_06_in10 = reg_0250;
    90: op1_06_in10 = reg_0432;
    66: op1_06_in10 = reg_0923;
    91: op1_06_in10 = reg_1230;
    95: op1_06_in10 = reg_1230;
    44: op1_06_in10 = reg_0578;
    93: op1_06_in10 = reg_0562;
    40: op1_06_in10 = reg_0002;
    94: op1_06_in10 = reg_0412;
    42: op1_06_in10 = reg_0386;
    97: op1_06_in10 = reg_1257;
    98: op1_06_in10 = reg_1227;
    99: op1_06_in10 = reg_0440;
    101: op1_06_in10 = imem02_in[7:4];
    102: op1_06_in10 = imem05_in[11:8];
    103: op1_06_in10 = reg_0419;
    104: op1_06_in10 = reg_1027;
    105: op1_06_in10 = reg_0488;
    106: op1_06_in10 = reg_0448;
    107: op1_06_in10 = reg_0387;
    108: op1_06_in10 = reg_0498;
    109: op1_06_in10 = reg_1225;
    110: op1_06_in10 = reg_1492;
    111: op1_06_in10 = reg_0086;
    112: op1_06_in10 = reg_0533;
    113: op1_06_in10 = reg_0977;
    114: op1_06_in10 = reg_0183;
    116: op1_06_in10 = reg_0829;
    118: op1_06_in10 = reg_0829;
    38: op1_06_in10 = reg_0087;
    117: op1_06_in10 = reg_1393;
    119: op1_06_in10 = reg_0276;
    120: op1_06_in10 = reg_0406;
    121: op1_06_in10 = reg_0303;
    122: op1_06_in10 = reg_0192;
    123: op1_06_in10 = reg_0014;
    124: op1_06_in10 = reg_1312;
    125: op1_06_in10 = reg_0126;
    126: op1_06_in10 = reg_0487;
    127: op1_06_in10 = reg_0802;
    128: op1_06_in10 = reg_0934;
    130: op1_06_in10 = reg_1201;
    131: op1_06_in10 = reg_0316;
    default: op1_06_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_06_inv10 = 1;
    86: op1_06_inv10 = 1;
    71: op1_06_inv10 = 1;
    50: op1_06_inv10 = 1;
    54: op1_06_inv10 = 1;
    75: op1_06_inv10 = 1;
    56: op1_06_inv10 = 1;
    60: op1_06_inv10 = 1;
    57: op1_06_inv10 = 1;
    33: op1_06_inv10 = 1;
    70: op1_06_inv10 = 1;
    78: op1_06_inv10 = 1;
    46: op1_06_inv10 = 1;
    59: op1_06_inv10 = 1;
    80: op1_06_inv10 = 1;
    62: op1_06_inv10 = 1;
    52: op1_06_inv10 = 1;
    82: op1_06_inv10 = 1;
    89: op1_06_inv10 = 1;
    64: op1_06_inv10 = 1;
    37: op1_06_inv10 = 1;
    47: op1_06_inv10 = 1;
    85: op1_06_inv10 = 1;
    90: op1_06_inv10 = 1;
    67: op1_06_inv10 = 1;
    92: op1_06_inv10 = 1;
    94: op1_06_inv10 = 1;
    95: op1_06_inv10 = 1;
    96: op1_06_inv10 = 1;
    42: op1_06_inv10 = 1;
    98: op1_06_inv10 = 1;
    100: op1_06_inv10 = 1;
    101: op1_06_inv10 = 1;
    102: op1_06_inv10 = 1;
    104: op1_06_inv10 = 1;
    106: op1_06_inv10 = 1;
    107: op1_06_inv10 = 1;
    108: op1_06_inv10 = 1;
    109: op1_06_inv10 = 1;
    111: op1_06_inv10 = 1;
    113: op1_06_inv10 = 1;
    124: op1_06_inv10 = 1;
    128: op1_06_inv10 = 1;
    130: op1_06_inv10 = 1;
    131: op1_06_inv10 = 1;
    default: op1_06_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in11 = reg_0428;
    53: op1_06_in11 = reg_0061;
    55: op1_06_in11 = reg_0622;
    86: op1_06_in11 = imem03_in[15:12];
    73: op1_06_in11 = reg_0527;
    69: op1_06_in11 = reg_0531;
    49: op1_06_in11 = reg_0051;
    71: op1_06_in11 = reg_0886;
    50: op1_06_in11 = reg_0156;
    54: op1_06_in11 = reg_0587;
    74: op1_06_in11 = reg_0155;
    68: op1_06_in11 = reg_0820;
    61: op1_06_in11 = reg_0725;
    75: op1_06_in11 = reg_0201;
    87: op1_06_in11 = reg_0291;
    89: op1_06_in11 = reg_0291;
    56: op1_06_in11 = reg_0373;
    76: op1_06_in11 = reg_0524;
    60: op1_06_in11 = reg_0463;
    57: op1_06_in11 = reg_0046;
    77: op1_06_in11 = reg_0459;
    33: op1_06_in11 = reg_0228;
    70: op1_06_in11 = imem02_in[7:4];
    58: op1_06_in11 = reg_0893;
    48: op1_06_in11 = reg_0334;
    78: op1_06_in11 = reg_0289;
    103: op1_06_in11 = reg_0289;
    46: op1_06_in11 = reg_0719;
    88: op1_06_in11 = reg_0694;
    51: op1_06_in11 = reg_0618;
    79: op1_06_in11 = reg_0492;
    59: op1_06_in11 = reg_1018;
    80: op1_06_in11 = reg_0370;
    62: op1_06_in11 = reg_0429;
    52: op1_06_in11 = reg_0494;
    81: op1_06_in11 = reg_0306;
    63: op1_06_in11 = reg_1315;
    82: op1_06_in11 = reg_0409;
    83: op1_06_in11 = reg_0939;
    64: op1_06_in11 = reg_0436;
    90: op1_06_in11 = reg_0436;
    84: op1_06_in11 = reg_0934;
    47: op1_06_in11 = reg_0413;
    65: op1_06_in11 = reg_1269;
    85: op1_06_in11 = reg_1459;
    66: op1_06_in11 = reg_0139;
    91: op1_06_in11 = reg_1432;
    95: op1_06_in11 = reg_1432;
    130: op1_06_in11 = reg_1432;
    44: op1_06_in11 = reg_0750;
    67: op1_06_in11 = reg_0181;
    92: op1_06_in11 = reg_1392;
    93: op1_06_in11 = reg_0173;
    40: op1_06_in11 = reg_0087;
    94: op1_06_in11 = reg_0407;
    96: op1_06_in11 = reg_1280;
    42: op1_06_in11 = reg_0385;
    97: op1_06_in11 = reg_1258;
    98: op1_06_in11 = reg_1230;
    104: op1_06_in11 = reg_1230;
    99: op1_06_in11 = reg_0416;
    100: op1_06_in11 = reg_0588;
    101: op1_06_in11 = reg_0276;
    102: op1_06_in11 = reg_0130;
    105: op1_06_in11 = reg_1233;
    106: op1_06_in11 = reg_0378;
    107: op1_06_in11 = reg_0075;
    108: op1_06_in11 = reg_0667;
    109: op1_06_in11 = reg_0132;
    110: op1_06_in11 = reg_0800;
    111: op1_06_in11 = reg_0518;
    112: op1_06_in11 = reg_1207;
    113: op1_06_in11 = reg_0214;
    114: op1_06_in11 = reg_1059;
    115: op1_06_in11 = reg_0351;
    116: op1_06_in11 = reg_0802;
    117: op1_06_in11 = reg_0202;
    118: op1_06_in11 = reg_0563;
    119: op1_06_in11 = reg_0561;
    120: op1_06_in11 = reg_0537;
    121: op1_06_in11 = reg_0240;
    122: op1_06_in11 = reg_0870;
    123: op1_06_in11 = reg_0908;
    124: op1_06_in11 = reg_0932;
    125: op1_06_in11 = reg_0628;
    126: op1_06_in11 = reg_0837;
    127: op1_06_in11 = reg_0711;
    128: op1_06_in11 = reg_0254;
    131: op1_06_in11 = reg_0263;
    default: op1_06_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv11 = 1;
    53: op1_06_inv11 = 1;
    86: op1_06_inv11 = 1;
    69: op1_06_inv11 = 1;
    49: op1_06_inv11 = 1;
    71: op1_06_inv11 = 1;
    68: op1_06_inv11 = 1;
    76: op1_06_inv11 = 1;
    57: op1_06_inv11 = 1;
    77: op1_06_inv11 = 1;
    70: op1_06_inv11 = 1;
    88: op1_06_inv11 = 1;
    79: op1_06_inv11 = 1;
    80: op1_06_inv11 = 1;
    62: op1_06_inv11 = 1;
    81: op1_06_inv11 = 1;
    83: op1_06_inv11 = 1;
    65: op1_06_inv11 = 1;
    85: op1_06_inv11 = 1;
    90: op1_06_inv11 = 1;
    66: op1_06_inv11 = 1;
    91: op1_06_inv11 = 1;
    44: op1_06_inv11 = 1;
    67: op1_06_inv11 = 1;
    92: op1_06_inv11 = 1;
    93: op1_06_inv11 = 1;
    94: op1_06_inv11 = 1;
    42: op1_06_inv11 = 1;
    98: op1_06_inv11 = 1;
    99: op1_06_inv11 = 1;
    101: op1_06_inv11 = 1;
    102: op1_06_inv11 = 1;
    103: op1_06_inv11 = 1;
    104: op1_06_inv11 = 1;
    105: op1_06_inv11 = 1;
    106: op1_06_inv11 = 1;
    111: op1_06_inv11 = 1;
    114: op1_06_inv11 = 1;
    116: op1_06_inv11 = 1;
    117: op1_06_inv11 = 1;
    118: op1_06_inv11 = 1;
    121: op1_06_inv11 = 1;
    124: op1_06_inv11 = 1;
    125: op1_06_inv11 = 1;
    126: op1_06_inv11 = 1;
    127: op1_06_inv11 = 1;
    default: op1_06_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in12 = reg_0387;
    53: op1_06_in12 = reg_0794;
    55: op1_06_in12 = reg_0624;
    86: op1_06_in12 = reg_1325;
    73: op1_06_in12 = reg_0571;
    69: op1_06_in12 = reg_0802;
    49: op1_06_in12 = reg_0086;
    71: op1_06_in12 = reg_0416;
    50: op1_06_in12 = reg_0169;
    54: op1_06_in12 = reg_0561;
    74: op1_06_in12 = reg_1418;
    68: op1_06_in12 = reg_0695;
    61: op1_06_in12 = reg_0201;
    117: op1_06_in12 = reg_0201;
    75: op1_06_in12 = reg_0440;
    87: op1_06_in12 = reg_0694;
    56: op1_06_in12 = reg_0109;
    76: op1_06_in12 = reg_1405;
    60: op1_06_in12 = reg_0252;
    57: op1_06_in12 = reg_1094;
    77: op1_06_in12 = reg_0927;
    91: op1_06_in12 = reg_0927;
    33: op1_06_in12 = reg_0003;
    70: op1_06_in12 = reg_0629;
    58: op1_06_in12 = reg_0187;
    48: op1_06_in12 = reg_0315;
    78: op1_06_in12 = reg_1202;
    46: op1_06_in12 = reg_0129;
    88: op1_06_in12 = reg_1383;
    51: op1_06_in12 = reg_0620;
    79: op1_06_in12 = reg_0799;
    59: op1_06_in12 = imem02_in[3:0];
    80: op1_06_in12 = reg_0175;
    62: op1_06_in12 = reg_0380;
    52: op1_06_in12 = reg_0472;
    81: op1_06_in12 = reg_0009;
    63: op1_06_in12 = reg_0298;
    82: op1_06_in12 = reg_0134;
    99: op1_06_in12 = reg_0134;
    89: op1_06_in12 = reg_0411;
    96: op1_06_in12 = reg_0411;
    83: op1_06_in12 = reg_0938;
    64: op1_06_in12 = reg_0326;
    84: op1_06_in12 = reg_0055;
    47: op1_06_in12 = reg_0100;
    65: op1_06_in12 = reg_1259;
    85: op1_06_in12 = reg_0821;
    90: op1_06_in12 = reg_0776;
    66: op1_06_in12 = reg_0777;
    44: op1_06_in12 = reg_0737;
    67: op1_06_in12 = reg_1367;
    92: op1_06_in12 = imem03_in[7:4];
    93: op1_06_in12 = reg_0701;
    40: op1_06_in12 = reg_0519;
    94: op1_06_in12 = reg_0471;
    95: op1_06_in12 = reg_0476;
    42: op1_06_in12 = reg_0362;
    97: op1_06_in12 = reg_1083;
    98: op1_06_in12 = reg_0987;
    100: op1_06_in12 = reg_0712;
    101: op1_06_in12 = reg_0744;
    119: op1_06_in12 = reg_0744;
    102: op1_06_in12 = reg_0118;
    103: op1_06_in12 = reg_0754;
    104: op1_06_in12 = reg_0460;
    105: op1_06_in12 = reg_1214;
    106: op1_06_in12 = reg_0288;
    107: op1_06_in12 = reg_1321;
    108: op1_06_in12 = reg_1440;
    109: op1_06_in12 = reg_0419;
    110: op1_06_in12 = reg_0563;
    111: op1_06_in12 = reg_0484;
    112: op1_06_in12 = reg_0494;
    113: op1_06_in12 = reg_0015;
    114: op1_06_in12 = reg_0793;
    115: op1_06_in12 = reg_0428;
    116: op1_06_in12 = reg_0800;
    118: op1_06_in12 = reg_0168;
    120: op1_06_in12 = reg_1065;
    121: op1_06_in12 = reg_0589;
    122: op1_06_in12 = reg_1209;
    123: op1_06_in12 = reg_0729;
    124: op1_06_in12 = reg_0065;
    125: op1_06_in12 = reg_0381;
    126: op1_06_in12 = reg_0420;
    127: op1_06_in12 = reg_0255;
    128: op1_06_in12 = reg_0455;
    130: op1_06_in12 = reg_0883;
    131: op1_06_in12 = reg_0120;
    default: op1_06_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv12 = 1;
    53: op1_06_inv12 = 1;
    86: op1_06_inv12 = 1;
    73: op1_06_inv12 = 1;
    69: op1_06_inv12 = 1;
    71: op1_06_inv12 = 1;
    61: op1_06_inv12 = 1;
    75: op1_06_inv12 = 1;
    87: op1_06_inv12 = 1;
    56: op1_06_inv12 = 1;
    60: op1_06_inv12 = 1;
    57: op1_06_inv12 = 1;
    77: op1_06_inv12 = 1;
    48: op1_06_inv12 = 1;
    88: op1_06_inv12 = 1;
    79: op1_06_inv12 = 1;
    80: op1_06_inv12 = 1;
    52: op1_06_inv12 = 1;
    64: op1_06_inv12 = 1;
    84: op1_06_inv12 = 1;
    90: op1_06_inv12 = 1;
    91: op1_06_inv12 = 1;
    92: op1_06_inv12 = 1;
    93: op1_06_inv12 = 1;
    94: op1_06_inv12 = 1;
    96: op1_06_inv12 = 1;
    42: op1_06_inv12 = 1;
    102: op1_06_inv12 = 1;
    103: op1_06_inv12 = 1;
    110: op1_06_inv12 = 1;
    111: op1_06_inv12 = 1;
    112: op1_06_inv12 = 1;
    114: op1_06_inv12 = 1;
    115: op1_06_inv12 = 1;
    117: op1_06_inv12 = 1;
    118: op1_06_inv12 = 1;
    120: op1_06_inv12 = 1;
    121: op1_06_inv12 = 1;
    122: op1_06_inv12 = 1;
    123: op1_06_inv12 = 1;
    124: op1_06_inv12 = 1;
    128: op1_06_inv12 = 1;
    130: op1_06_inv12 = 1;
    default: op1_06_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in13 = reg_0073;
    53: op1_06_in13 = reg_0579;
    55: op1_06_in13 = reg_0585;
    86: op1_06_in13 = reg_0427;
    73: op1_06_in13 = reg_0345;
    69: op1_06_in13 = reg_0757;
    49: op1_06_in13 = reg_0520;
    71: op1_06_in13 = reg_0058;
    50: op1_06_in13 = reg_0777;
    54: op1_06_in13 = reg_0560;
    74: op1_06_in13 = reg_0459;
    68: op1_06_in13 = reg_0802;
    61: op1_06_in13 = reg_0416;
    75: op1_06_in13 = reg_0122;
    87: op1_06_in13 = reg_0032;
    56: op1_06_in13 = reg_0670;
    76: op1_06_in13 = reg_0353;
    60: op1_06_in13 = reg_0978;
    57: op1_06_in13 = imem07_in[7:4];
    77: op1_06_in13 = reg_0886;
    91: op1_06_in13 = reg_0886;
    130: op1_06_in13 = reg_0886;
    33: op1_06_in13 = reg_0086;
    70: op1_06_in13 = reg_0496;
    58: op1_06_in13 = reg_0851;
    48: op1_06_in13 = reg_0938;
    78: op1_06_in13 = reg_0018;
    46: op1_06_in13 = reg_0211;
    88: op1_06_in13 = reg_1372;
    51: op1_06_in13 = reg_0114;
    79: op1_06_in13 = reg_0449;
    59: op1_06_in13 = imem02_in[7:4];
    80: op1_06_in13 = reg_0272;
    62: op1_06_in13 = reg_0898;
    52: op1_06_in13 = reg_0473;
    125: op1_06_in13 = reg_0473;
    81: op1_06_in13 = reg_0379;
    63: op1_06_in13 = reg_0893;
    82: op1_06_in13 = reg_0387;
    89: op1_06_in13 = reg_0534;
    83: op1_06_in13 = reg_0477;
    64: op1_06_in13 = reg_0971;
    84: op1_06_in13 = reg_0474;
    47: op1_06_in13 = reg_0051;
    65: op1_06_in13 = reg_1163;
    85: op1_06_in13 = reg_1405;
    90: op1_06_in13 = reg_0326;
    66: op1_06_in13 = reg_0779;
    44: op1_06_in13 = reg_0346;
    67: op1_06_in13 = reg_1338;
    92: op1_06_in13 = imem03_in[15:12];
    93: op1_06_in13 = reg_0630;
    94: op1_06_in13 = reg_0454;
    95: op1_06_in13 = reg_0928;
    96: op1_06_in13 = reg_0252;
    113: op1_06_in13 = reg_0252;
    42: op1_06_in13 = reg_0320;
    97: op1_06_in13 = reg_0681;
    98: op1_06_in13 = reg_1201;
    99: op1_06_in13 = reg_0203;
    100: op1_06_in13 = reg_0532;
    101: op1_06_in13 = reg_1002;
    102: op1_06_in13 = reg_0240;
    103: op1_06_in13 = reg_0023;
    104: op1_06_in13 = reg_1418;
    105: op1_06_in13 = reg_0414;
    106: op1_06_in13 = reg_0411;
    107: op1_06_in13 = reg_0057;
    108: op1_06_in13 = reg_0703;
    109: op1_06_in13 = reg_0215;
    110: op1_06_in13 = reg_0632;
    118: op1_06_in13 = reg_0632;
    112: op1_06_in13 = reg_0432;
    114: op1_06_in13 = reg_0445;
    115: op1_06_in13 = reg_0440;
    116: op1_06_in13 = reg_0253;
    117: op1_06_in13 = reg_0059;
    119: op1_06_in13 = reg_0822;
    120: op1_06_in13 = reg_0836;
    121: op1_06_in13 = reg_0603;
    122: op1_06_in13 = reg_1420;
    123: op1_06_in13 = reg_0925;
    124: op1_06_in13 = reg_0095;
    126: op1_06_in13 = reg_0633;
    127: op1_06_in13 = reg_0952;
    128: op1_06_in13 = reg_0839;
    131: op1_06_in13 = reg_0960;
    default: op1_06_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_06_inv13 = 1;
    69: op1_06_inv13 = 1;
    71: op1_06_inv13 = 1;
    50: op1_06_inv13 = 1;
    74: op1_06_inv13 = 1;
    68: op1_06_inv13 = 1;
    56: op1_06_inv13 = 1;
    60: op1_06_inv13 = 1;
    33: op1_06_inv13 = 1;
    70: op1_06_inv13 = 1;
    48: op1_06_inv13 = 1;
    78: op1_06_inv13 = 1;
    59: op1_06_inv13 = 1;
    52: op1_06_inv13 = 1;
    63: op1_06_inv13 = 1;
    82: op1_06_inv13 = 1;
    89: op1_06_inv13 = 1;
    83: op1_06_inv13 = 1;
    64: op1_06_inv13 = 1;
    85: op1_06_inv13 = 1;
    90: op1_06_inv13 = 1;
    66: op1_06_inv13 = 1;
    91: op1_06_inv13 = 1;
    67: op1_06_inv13 = 1;
    92: op1_06_inv13 = 1;
    93: op1_06_inv13 = 1;
    94: op1_06_inv13 = 1;
    96: op1_06_inv13 = 1;
    98: op1_06_inv13 = 1;
    105: op1_06_inv13 = 1;
    107: op1_06_inv13 = 1;
    110: op1_06_inv13 = 1;
    112: op1_06_inv13 = 1;
    115: op1_06_inv13 = 1;
    120: op1_06_inv13 = 1;
    124: op1_06_inv13 = 1;
    125: op1_06_inv13 = 1;
    128: op1_06_inv13 = 1;
    130: op1_06_inv13 = 1;
    131: op1_06_inv13 = 1;
    default: op1_06_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in14 = reg_0026;
    53: op1_06_in14 = reg_0745;
    55: op1_06_in14 = reg_0586;
    86: op1_06_in14 = reg_0411;
    73: op1_06_in14 = reg_0165;
    69: op1_06_in14 = reg_0121;
    49: op1_06_in14 = reg_0123;
    71: op1_06_in14 = reg_1253;
    50: op1_06_in14 = reg_0775;
    54: op1_06_in14 = reg_1139;
    74: op1_06_in14 = reg_0886;
    95: op1_06_in14 = reg_0886;
    68: op1_06_in14 = reg_0800;
    61: op1_06_in14 = reg_0409;
    75: op1_06_in14 = reg_0089;
    87: op1_06_in14 = reg_0535;
    88: op1_06_in14 = reg_0535;
    56: op1_06_in14 = reg_0634;
    76: op1_06_in14 = reg_0722;
    60: op1_06_in14 = reg_0577;
    57: op1_06_in14 = imem07_in[11:8];
    109: op1_06_in14 = imem07_in[11:8];
    77: op1_06_in14 = reg_0202;
    91: op1_06_in14 = reg_0202;
    33: op1_06_in14 = reg_0084;
    70: op1_06_in14 = reg_0138;
    58: op1_06_in14 = reg_0673;
    48: op1_06_in14 = reg_0477;
    78: op1_06_in14 = reg_0022;
    46: op1_06_in14 = reg_0063;
    51: op1_06_in14 = reg_0002;
    47: op1_06_in14 = reg_0002;
    79: op1_06_in14 = reg_0151;
    59: op1_06_in14 = reg_0497;
    80: op1_06_in14 = reg_0578;
    62: op1_06_in14 = reg_0708;
    52: op1_06_in14 = reg_0436;
    81: op1_06_in14 = reg_0801;
    63: op1_06_in14 = reg_0297;
    82: op1_06_in14 = reg_0075;
    89: op1_06_in14 = reg_0694;
    83: op1_06_in14 = reg_0302;
    64: op1_06_in14 = reg_0128;
    84: op1_06_in14 = reg_0054;
    65: op1_06_in14 = reg_0648;
    85: op1_06_in14 = reg_0881;
    90: op1_06_in14 = reg_0971;
    66: op1_06_in14 = reg_0029;
    44: op1_06_in14 = reg_0832;
    67: op1_06_in14 = reg_1198;
    92: op1_06_in14 = reg_0328;
    118: op1_06_in14 = reg_0328;
    93: op1_06_in14 = reg_0418;
    94: op1_06_in14 = reg_0061;
    96: op1_06_in14 = imem04_in[15:12];
    42: op1_06_in14 = reg_0093;
    97: op1_06_in14 = reg_0599;
    98: op1_06_in14 = reg_0460;
    99: op1_06_in14 = reg_1324;
    100: op1_06_in14 = reg_1002;
    101: op1_06_in14 = reg_0495;
    102: op1_06_in14 = reg_1348;
    103: op1_06_in14 = reg_0215;
    104: op1_06_in14 = reg_0524;
    105: op1_06_in14 = reg_0969;
    106: op1_06_in14 = imem04_in[7:4];
    107: op1_06_in14 = reg_0005;
    108: op1_06_in14 = reg_1350;
    110: op1_06_in14 = reg_0006;
    112: op1_06_in14 = reg_0112;
    113: op1_06_in14 = reg_0190;
    114: op1_06_in14 = reg_0702;
    115: op1_06_in14 = reg_0073;
    116: op1_06_in14 = reg_1515;
    117: op1_06_in14 = reg_1321;
    119: op1_06_in14 = reg_0900;
    120: op1_06_in14 = reg_0096;
    121: op1_06_in14 = reg_0864;
    122: op1_06_in14 = reg_0782;
    123: op1_06_in14 = reg_0751;
    124: op1_06_in14 = reg_0019;
    125: op1_06_in14 = reg_1492;
    126: op1_06_in14 = reg_0021;
    127: op1_06_in14 = reg_1009;
    128: op1_06_in14 = reg_0744;
    130: op1_06_in14 = reg_0743;
    131: op1_06_in14 = reg_0869;
    default: op1_06_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_06_inv14 = 1;
    73: op1_06_inv14 = 1;
    69: op1_06_inv14 = 1;
    71: op1_06_inv14 = 1;
    74: op1_06_inv14 = 1;
    68: op1_06_inv14 = 1;
    56: op1_06_inv14 = 1;
    76: op1_06_inv14 = 1;
    60: op1_06_inv14 = 1;
    57: op1_06_inv14 = 1;
    70: op1_06_inv14 = 1;
    58: op1_06_inv14 = 1;
    48: op1_06_inv14 = 1;
    78: op1_06_inv14 = 1;
    46: op1_06_inv14 = 1;
    80: op1_06_inv14 = 1;
    63: op1_06_inv14 = 1;
    82: op1_06_inv14 = 1;
    65: op1_06_inv14 = 1;
    85: op1_06_inv14 = 1;
    91: op1_06_inv14 = 1;
    67: op1_06_inv14 = 1;
    93: op1_06_inv14 = 1;
    94: op1_06_inv14 = 1;
    97: op1_06_inv14 = 1;
    99: op1_06_inv14 = 1;
    100: op1_06_inv14 = 1;
    103: op1_06_inv14 = 1;
    105: op1_06_inv14 = 1;
    107: op1_06_inv14 = 1;
    108: op1_06_inv14 = 1;
    110: op1_06_inv14 = 1;
    112: op1_06_inv14 = 1;
    115: op1_06_inv14 = 1;
    116: op1_06_inv14 = 1;
    117: op1_06_inv14 = 1;
    118: op1_06_inv14 = 1;
    121: op1_06_inv14 = 1;
    123: op1_06_inv14 = 1;
    127: op1_06_inv14 = 1;
    128: op1_06_inv14 = 1;
    130: op1_06_inv14 = 1;
    131: op1_06_inv14 = 1;
    default: op1_06_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in15 = reg_0027;
    53: op1_06_in15 = reg_0749;
    55: op1_06_in15 = reg_0584;
    86: op1_06_in15 = reg_0898;
    73: op1_06_in15 = imem07_in[11:8];
    69: op1_06_in15 = reg_0154;
    71: op1_06_in15 = reg_1256;
    107: op1_06_in15 = reg_1256;
    50: op1_06_in15 = reg_0465;
    54: op1_06_in15 = reg_0473;
    74: op1_06_in15 = reg_0202;
    68: op1_06_in15 = reg_0279;
    61: op1_06_in15 = reg_0073;
    75: op1_06_in15 = reg_0026;
    87: op1_06_in15 = reg_0599;
    56: op1_06_in15 = reg_0568;
    76: op1_06_in15 = reg_0189;
    60: op1_06_in15 = reg_0574;
    67: op1_06_in15 = reg_0574;
    57: op1_06_in15 = reg_0496;
    77: op1_06_in15 = reg_0428;
    33: op1_06_in15 = reg_0087;
    70: op1_06_in15 = reg_0705;
    58: op1_06_in15 = reg_0158;
    48: op1_06_in15 = reg_0896;
    78: op1_06_in15 = reg_0706;
    46: op1_06_in15 = reg_0035;
    88: op1_06_in15 = reg_0297;
    51: op1_06_in15 = reg_0052;
    79: op1_06_in15 = reg_0206;
    59: op1_06_in15 = reg_0474;
    80: op1_06_in15 = reg_0315;
    62: op1_06_in15 = reg_0007;
    52: op1_06_in15 = reg_0973;
    81: op1_06_in15 = reg_0327;
    63: op1_06_in15 = imem07_in[3:0];
    82: op1_06_in15 = reg_0060;
    115: op1_06_in15 = reg_0060;
    89: op1_06_in15 = reg_0032;
    83: op1_06_in15 = reg_0300;
    64: op1_06_in15 = reg_0382;
    84: op1_06_in15 = reg_1451;
    47: op1_06_in15 = reg_0053;
    65: op1_06_in15 = reg_0538;
    85: op1_06_in15 = reg_0887;
    90: op1_06_in15 = reg_1455;
    66: op1_06_in15 = reg_0739;
    91: op1_06_in15 = reg_0351;
    44: op1_06_in15 = reg_0702;
    92: op1_06_in15 = reg_0573;
    93: op1_06_in15 = reg_0301;
    94: op1_06_in15 = reg_0698;
    95: op1_06_in15 = reg_0188;
    96: op1_06_in15 = reg_1383;
    42: op1_06_in15 = imem01_in[3:0];
    97: op1_06_in15 = reg_1041;
    105: op1_06_in15 = reg_1041;
    98: op1_06_in15 = reg_1405;
    104: op1_06_in15 = reg_1405;
    99: op1_06_in15 = reg_0089;
    100: op1_06_in15 = reg_1450;
    101: op1_06_in15 = reg_0433;
    102: op1_06_in15 = reg_0344;
    103: op1_06_in15 = reg_0015;
    106: op1_06_in15 = imem04_in[15:12];
    108: op1_06_in15 = reg_0489;
    109: op1_06_in15 = reg_0998;
    110: op1_06_in15 = reg_0989;
    112: op1_06_in15 = reg_0684;
    113: op1_06_in15 = reg_0394;
    114: op1_06_in15 = reg_0184;
    116: op1_06_in15 = reg_0235;
    117: op1_06_in15 = reg_1324;
    118: op1_06_in15 = reg_0750;
    119: op1_06_in15 = reg_0472;
    120: op1_06_in15 = reg_1189;
    121: op1_06_in15 = reg_0207;
    122: op1_06_in15 = reg_0696;
    123: op1_06_in15 = reg_0752;
    124: op1_06_in15 = imem05_in[3:0];
    125: op1_06_in15 = reg_0801;
    126: op1_06_in15 = reg_0470;
    127: op1_06_in15 = imem03_in[11:8];
    128: op1_06_in15 = reg_0106;
    130: op1_06_in15 = reg_0830;
    131: op1_06_in15 = reg_1504;
    default: op1_06_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv15 = 1;
    55: op1_06_inv15 = 1;
    86: op1_06_inv15 = 1;
    71: op1_06_inv15 = 1;
    74: op1_06_inv15 = 1;
    68: op1_06_inv15 = 1;
    75: op1_06_inv15 = 1;
    87: op1_06_inv15 = 1;
    60: op1_06_inv15 = 1;
    57: op1_06_inv15 = 1;
    77: op1_06_inv15 = 1;
    33: op1_06_inv15 = 1;
    46: op1_06_inv15 = 1;
    51: op1_06_inv15 = 1;
    59: op1_06_inv15 = 1;
    80: op1_06_inv15 = 1;
    62: op1_06_inv15 = 1;
    52: op1_06_inv15 = 1;
    81: op1_06_inv15 = 1;
    63: op1_06_inv15 = 1;
    83: op1_06_inv15 = 1;
    64: op1_06_inv15 = 1;
    85: op1_06_inv15 = 1;
    90: op1_06_inv15 = 1;
    66: op1_06_inv15 = 1;
    91: op1_06_inv15 = 1;
    44: op1_06_inv15 = 1;
    93: op1_06_inv15 = 1;
    94: op1_06_inv15 = 1;
    95: op1_06_inv15 = 1;
    96: op1_06_inv15 = 1;
    97: op1_06_inv15 = 1;
    101: op1_06_inv15 = 1;
    104: op1_06_inv15 = 1;
    105: op1_06_inv15 = 1;
    108: op1_06_inv15 = 1;
    110: op1_06_inv15 = 1;
    112: op1_06_inv15 = 1;
    115: op1_06_inv15 = 1;
    116: op1_06_inv15 = 1;
    117: op1_06_inv15 = 1;
    120: op1_06_inv15 = 1;
    124: op1_06_inv15 = 1;
    126: op1_06_inv15 = 1;
    128: op1_06_inv15 = 1;
    default: op1_06_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in16 = reg_0786;
    53: op1_06_in16 = reg_0750;
    55: op1_06_in16 = reg_0529;
    86: op1_06_in16 = reg_0696;
    73: op1_06_in16 = reg_1439;
    69: op1_06_in16 = reg_0707;
    71: op1_06_in16 = reg_0576;
    50: op1_06_in16 = reg_0664;
    54: op1_06_in16 = reg_0326;
    74: op1_06_in16 = reg_0352;
    68: op1_06_in16 = reg_0311;
    61: op1_06_in16 = reg_0075;
    75: op1_06_in16 = reg_1100;
    87: op1_06_in16 = reg_1065;
    56: op1_06_in16 = reg_1204;
    76: op1_06_in16 = reg_0440;
    60: op1_06_in16 = reg_1083;
    88: op1_06_in16 = reg_1083;
    67: op1_06_in16 = reg_1083;
    57: op1_06_in16 = reg_1183;
    77: op1_06_in16 = reg_0203;
    33: op1_06_in16 = reg_0519;
    70: op1_06_in16 = reg_0007;
    58: op1_06_in16 = reg_0923;
    48: op1_06_in16 = reg_0302;
    78: op1_06_in16 = reg_1440;
    46: op1_06_in16 = reg_0391;
    51: op1_06_in16 = reg_0085;
    79: op1_06_in16 = reg_0037;
    59: op1_06_in16 = reg_0971;
    80: op1_06_in16 = reg_0702;
    62: op1_06_in16 = reg_0008;
    52: op1_06_in16 = reg_0935;
    81: op1_06_in16 = reg_1392;
    63: op1_06_in16 = reg_0159;
    82: op1_06_in16 = reg_0057;
    89: op1_06_in16 = reg_1368;
    83: op1_06_in16 = reg_0090;
    93: op1_06_in16 = reg_0090;
    64: op1_06_in16 = reg_0379;
    84: op1_06_in16 = reg_0125;
    90: op1_06_in16 = reg_0125;
    47: op1_06_in16 = reg_0086;
    65: op1_06_in16 = reg_0167;
    85: op1_06_in16 = reg_0883;
    66: op1_06_in16 = reg_0028;
    91: op1_06_in16 = reg_0188;
    44: op1_06_in16 = reg_0173;
    92: op1_06_in16 = reg_0179;
    94: op1_06_in16 = reg_0582;
    95: op1_06_in16 = reg_0201;
    96: op1_06_in16 = reg_0535;
    42: op1_06_in16 = imem01_in[15:12];
    97: op1_06_in16 = reg_1077;
    98: op1_06_in16 = reg_0351;
    99: op1_06_in16 = reg_0026;
    100: op1_06_in16 = reg_0382;
    101: op1_06_in16 = reg_0429;
    102: op1_06_in16 = reg_0828;
    103: op1_06_in16 = reg_0022;
    104: op1_06_in16 = reg_0476;
    105: op1_06_in16 = reg_0537;
    106: op1_06_in16 = reg_0208;
    107: op1_06_in16 = reg_1290;
    108: op1_06_in16 = reg_0223;
    109: op1_06_in16 = reg_0893;
    110: op1_06_in16 = reg_0479;
    118: op1_06_in16 = reg_0479;
    112: op1_06_in16 = reg_0628;
    113: op1_06_in16 = reg_1095;
    114: op1_06_in16 = reg_0346;
    115: op1_06_in16 = reg_1321;
    116: op1_06_in16 = reg_0677;
    117: op1_06_in16 = reg_1322;
    119: op1_06_in16 = reg_1207;
    120: op1_06_in16 = reg_0932;
    121: op1_06_in16 = reg_0565;
    122: op1_06_in16 = reg_0271;
    123: op1_06_in16 = reg_1501;
    124: op1_06_in16 = reg_0735;
    125: op1_06_in16 = reg_0294;
    126: op1_06_in16 = imem05_in[7:4];
    127: op1_06_in16 = reg_0597;
    128: op1_06_in16 = reg_0105;
    130: op1_06_in16 = reg_0798;
    131: op1_06_in16 = reg_1508;
    default: op1_06_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv16 = 1;
    55: op1_06_inv16 = 1;
    86: op1_06_inv16 = 1;
    73: op1_06_inv16 = 1;
    50: op1_06_inv16 = 1;
    54: op1_06_inv16 = 1;
    68: op1_06_inv16 = 1;
    61: op1_06_inv16 = 1;
    75: op1_06_inv16 = 1;
    77: op1_06_inv16 = 1;
    33: op1_06_inv16 = 1;
    70: op1_06_inv16 = 1;
    78: op1_06_inv16 = 1;
    46: op1_06_inv16 = 1;
    88: op1_06_inv16 = 1;
    51: op1_06_inv16 = 1;
    79: op1_06_inv16 = 1;
    59: op1_06_inv16 = 1;
    80: op1_06_inv16 = 1;
    62: op1_06_inv16 = 1;
    63: op1_06_inv16 = 1;
    47: op1_06_inv16 = 1;
    65: op1_06_inv16 = 1;
    85: op1_06_inv16 = 1;
    90: op1_06_inv16 = 1;
    66: op1_06_inv16 = 1;
    92: op1_06_inv16 = 1;
    93: op1_06_inv16 = 1;
    95: op1_06_inv16 = 1;
    96: op1_06_inv16 = 1;
    42: op1_06_inv16 = 1;
    97: op1_06_inv16 = 1;
    100: op1_06_inv16 = 1;
    103: op1_06_inv16 = 1;
    104: op1_06_inv16 = 1;
    105: op1_06_inv16 = 1;
    108: op1_06_inv16 = 1;
    115: op1_06_inv16 = 1;
    119: op1_06_inv16 = 1;
    120: op1_06_inv16 = 1;
    121: op1_06_inv16 = 1;
    122: op1_06_inv16 = 1;
    123: op1_06_inv16 = 1;
    124: op1_06_inv16 = 1;
    126: op1_06_inv16 = 1;
    127: op1_06_inv16 = 1;
    default: op1_06_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in17 = reg_0372;
    53: op1_06_in17 = reg_0733;
    114: op1_06_in17 = reg_0733;
    55: op1_06_in17 = reg_0171;
    86: op1_06_in17 = reg_1368;
    73: op1_06_in17 = reg_0490;
    69: op1_06_in17 = imem03_in[7:4];
    71: op1_06_in17 = reg_0260;
    50: op1_06_in17 = reg_0286;
    54: op1_06_in17 = reg_0935;
    74: op1_06_in17 = reg_0440;
    68: op1_06_in17 = reg_0198;
    92: op1_06_in17 = reg_0198;
    61: op1_06_in17 = reg_0060;
    75: op1_06_in17 = reg_1068;
    87: op1_06_in17 = reg_1004;
    97: op1_06_in17 = reg_1004;
    56: op1_06_in17 = reg_1202;
    76: op1_06_in17 = reg_1034;
    60: op1_06_in17 = reg_0406;
    57: op1_06_in17 = reg_0668;
    77: op1_06_in17 = reg_0089;
    33: op1_06_in17 = reg_0518;
    70: op1_06_in17 = reg_0820;
    58: op1_06_in17 = reg_0791;
    48: op1_06_in17 = reg_0090;
    78: op1_06_in17 = reg_0922;
    46: op1_06_in17 = reg_0750;
    88: op1_06_in17 = reg_1203;
    51: op1_06_in17 = reg_0084;
    79: op1_06_in17 = imem06_in[7:4];
    59: op1_06_in17 = reg_0972;
    80: op1_06_in17 = reg_0877;
    62: op1_06_in17 = reg_0068;
    52: op1_06_in17 = reg_0307;
    81: op1_06_in17 = imem02_in[3:0];
    63: op1_06_in17 = reg_0924;
    82: op1_06_in17 = reg_0122;
    89: op1_06_in17 = reg_0264;
    83: op1_06_in17 = reg_0576;
    107: op1_06_in17 = reg_0576;
    64: op1_06_in17 = reg_0900;
    84: op1_06_in17 = reg_0105;
    47: op1_06_in17 = reg_0484;
    65: op1_06_in17 = reg_0163;
    85: op1_06_in17 = reg_0410;
    90: op1_06_in17 = reg_0126;
    66: op1_06_in17 = reg_0361;
    91: op1_06_in17 = reg_0409;
    44: op1_06_in17 = reg_0523;
    67: op1_06_in17 = reg_0681;
    96: op1_06_in17 = reg_0681;
    93: op1_06_in17 = reg_0275;
    94: op1_06_in17 = reg_0368;
    95: op1_06_in17 = reg_0416;
    42: op1_06_in17 = reg_0277;
    98: op1_06_in17 = reg_0201;
    99: op1_06_in17 = reg_0282;
    100: op1_06_in17 = reg_0745;
    101: op1_06_in17 = reg_0970;
    102: op1_06_in17 = imem06_in[11:8];
    103: op1_06_in17 = reg_0394;
    104: op1_06_in17 = reg_0351;
    105: op1_06_in17 = reg_0836;
    106: op1_06_in17 = reg_0032;
    108: op1_06_in17 = reg_0774;
    109: op1_06_in17 = reg_1183;
    110: op1_06_in17 = imem03_in[11:8];
    112: op1_06_in17 = reg_0829;
    113: op1_06_in17 = imem07_in[3:0];
    115: op1_06_in17 = reg_0057;
    116: op1_06_in17 = reg_0185;
    117: op1_06_in17 = reg_0723;
    118: op1_06_in17 = reg_0376;
    119: op1_06_in17 = reg_0494;
    120: op1_06_in17 = reg_0117;
    121: op1_06_in17 = reg_1299;
    122: op1_06_in17 = reg_1326;
    123: op1_06_in17 = reg_1179;
    124: op1_06_in17 = reg_0395;
    125: op1_06_in17 = reg_0007;
    126: op1_06_in17 = reg_0579;
    127: op1_06_in17 = reg_0220;
    128: op1_06_in17 = reg_0629;
    130: op1_06_in17 = reg_0715;
    131: op1_06_in17 = reg_0110;
    default: op1_06_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_06_inv17 = 1;
    73: op1_06_inv17 = 1;
    71: op1_06_inv17 = 1;
    54: op1_06_inv17 = 1;
    74: op1_06_inv17 = 1;
    68: op1_06_inv17 = 1;
    61: op1_06_inv17 = 1;
    75: op1_06_inv17 = 1;
    87: op1_06_inv17 = 1;
    56: op1_06_inv17 = 1;
    76: op1_06_inv17 = 1;
    77: op1_06_inv17 = 1;
    48: op1_06_inv17 = 1;
    46: op1_06_inv17 = 1;
    88: op1_06_inv17 = 1;
    59: op1_06_inv17 = 1;
    80: op1_06_inv17 = 1;
    62: op1_06_inv17 = 1;
    52: op1_06_inv17 = 1;
    81: op1_06_inv17 = 1;
    82: op1_06_inv17 = 1;
    89: op1_06_inv17 = 1;
    64: op1_06_inv17 = 1;
    84: op1_06_inv17 = 1;
    47: op1_06_inv17 = 1;
    65: op1_06_inv17 = 1;
    90: op1_06_inv17 = 1;
    93: op1_06_inv17 = 1;
    94: op1_06_inv17 = 1;
    95: op1_06_inv17 = 1;
    96: op1_06_inv17 = 1;
    98: op1_06_inv17 = 1;
    102: op1_06_inv17 = 1;
    105: op1_06_inv17 = 1;
    106: op1_06_inv17 = 1;
    107: op1_06_inv17 = 1;
    108: op1_06_inv17 = 1;
    109: op1_06_inv17 = 1;
    110: op1_06_inv17 = 1;
    116: op1_06_inv17 = 1;
    121: op1_06_inv17 = 1;
    122: op1_06_inv17 = 1;
    123: op1_06_inv17 = 1;
    124: op1_06_inv17 = 1;
    125: op1_06_inv17 = 1;
    130: op1_06_inv17 = 1;
    131: op1_06_inv17 = 1;
    default: op1_06_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in18 = reg_0788;
    76: op1_06_in18 = reg_0788;
    53: op1_06_in18 = reg_1059;
    55: op1_06_in18 = reg_0165;
    86: op1_06_in18 = reg_0493;
    73: op1_06_in18 = reg_0162;
    69: op1_06_in18 = reg_0963;
    71: op1_06_in18 = reg_0550;
    50: op1_06_in18 = reg_0437;
    54: op1_06_in18 = reg_0125;
    74: op1_06_in18 = reg_0416;
    68: op1_06_in18 = reg_0232;
    61: op1_06_in18 = imem01_in[7:4];
    115: op1_06_in18 = imem01_in[7:4];
    75: op1_06_in18 = imem01_in[3:0];
    117: op1_06_in18 = imem01_in[3:0];
    87: op1_06_in18 = reg_0342;
    56: op1_06_in18 = reg_0046;
    60: op1_06_in18 = reg_0370;
    57: op1_06_in18 = reg_0894;
    77: op1_06_in18 = reg_0917;
    70: op1_06_in18 = reg_0801;
    58: op1_06_in18 = reg_0287;
    48: op1_06_in18 = reg_0873;
    78: op1_06_in18 = reg_0310;
    46: op1_06_in18 = reg_0347;
    80: op1_06_in18 = reg_0347;
    88: op1_06_in18 = reg_0488;
    79: op1_06_in18 = reg_0261;
    59: op1_06_in18 = reg_0154;
    62: op1_06_in18 = reg_0557;
    52: op1_06_in18 = reg_0878;
    81: op1_06_in18 = imem02_in[7:4];
    63: op1_06_in18 = reg_0777;
    82: op1_06_in18 = reg_0089;
    89: op1_06_in18 = reg_0252;
    83: op1_06_in18 = reg_0038;
    64: op1_06_in18 = reg_0307;
    84: op1_06_in18 = reg_0496;
    65: op1_06_in18 = reg_0367;
    85: op1_06_in18 = reg_0026;
    90: op1_06_in18 = reg_0745;
    66: op1_06_in18 = reg_0003;
    91: op1_06_in18 = reg_0075;
    44: op1_06_in18 = reg_0604;
    67: op1_06_in18 = reg_0552;
    92: op1_06_in18 = reg_0191;
    93: op1_06_in18 = reg_1346;
    94: op1_06_in18 = reg_0837;
    95: op1_06_in18 = reg_0058;
    96: op1_06_in18 = reg_0421;
    42: op1_06_in18 = reg_0282;
    97: op1_06_in18 = reg_1419;
    98: op1_06_in18 = reg_0409;
    99: op1_06_in18 = reg_1031;
    100: op1_06_in18 = reg_0802;
    101: op1_06_in18 = reg_0972;
    102: op1_06_in18 = reg_1030;
    103: op1_06_in18 = reg_1010;
    104: op1_06_in18 = reg_0435;
    105: op1_06_in18 = reg_0835;
    106: op1_06_in18 = reg_1369;
    107: op1_06_in18 = reg_0609;
    108: op1_06_in18 = reg_0465;
    109: op1_06_in18 = reg_0461;
    110: op1_06_in18 = reg_0559;
    112: op1_06_in18 = reg_0897;
    113: op1_06_in18 = reg_1055;
    114: op1_06_in18 = reg_1164;
    116: op1_06_in18 = reg_0179;
    118: op1_06_in18 = imem03_in[3:0];
    119: op1_06_in18 = reg_1451;
    120: op1_06_in18 = reg_0065;
    121: op1_06_in18 = reg_0270;
    122: op1_06_in18 = reg_0720;
    123: op1_06_in18 = reg_1508;
    124: op1_06_in18 = reg_0251;
    125: op1_06_in18 = reg_1006;
    126: op1_06_in18 = reg_0832;
    127: op1_06_in18 = reg_1001;
    128: op1_06_in18 = reg_1433;
    130: op1_06_in18 = reg_0726;
    131: op1_06_in18 = reg_1303;
    default: op1_06_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_06_inv18 = 1;
    73: op1_06_inv18 = 1;
    50: op1_06_inv18 = 1;
    75: op1_06_inv18 = 1;
    60: op1_06_inv18 = 1;
    57: op1_06_inv18 = 1;
    77: op1_06_inv18 = 1;
    58: op1_06_inv18 = 1;
    46: op1_06_inv18 = 1;
    88: op1_06_inv18 = 1;
    79: op1_06_inv18 = 1;
    80: op1_06_inv18 = 1;
    62: op1_06_inv18 = 1;
    81: op1_06_inv18 = 1;
    63: op1_06_inv18 = 1;
    89: op1_06_inv18 = 1;
    64: op1_06_inv18 = 1;
    91: op1_06_inv18 = 1;
    44: op1_06_inv18 = 1;
    93: op1_06_inv18 = 1;
    94: op1_06_inv18 = 1;
    96: op1_06_inv18 = 1;
    42: op1_06_inv18 = 1;
    97: op1_06_inv18 = 1;
    98: op1_06_inv18 = 1;
    99: op1_06_inv18 = 1;
    100: op1_06_inv18 = 1;
    105: op1_06_inv18 = 1;
    107: op1_06_inv18 = 1;
    109: op1_06_inv18 = 1;
    112: op1_06_inv18 = 1;
    117: op1_06_inv18 = 1;
    122: op1_06_inv18 = 1;
    123: op1_06_inv18 = 1;
    125: op1_06_inv18 = 1;
    127: op1_06_inv18 = 1;
    128: op1_06_inv18 = 1;
    131: op1_06_inv18 = 1;
    default: op1_06_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in19 = reg_1032;
    84: op1_06_in19 = reg_1032;
    53: op1_06_in19 = reg_0702;
    55: op1_06_in19 = reg_1179;
    86: op1_06_in19 = imem04_in[7:4];
    73: op1_06_in19 = reg_0298;
    69: op1_06_in19 = reg_1314;
    71: op1_06_in19 = reg_0161;
    50: op1_06_in19 = reg_0741;
    54: op1_06_in19 = reg_0126;
    119: op1_06_in19 = reg_0126;
    74: op1_06_in19 = reg_0405;
    68: op1_06_in19 = reg_0375;
    61: op1_06_in19 = imem01_in[11:8];
    115: op1_06_in19 = imem01_in[11:8];
    75: op1_06_in19 = reg_0258;
    87: op1_06_in19 = reg_0698;
    56: op1_06_in19 = reg_0022;
    76: op1_06_in19 = reg_1256;
    60: op1_06_in19 = reg_0320;
    57: op1_06_in19 = reg_0310;
    77: op1_06_in19 = reg_1100;
    85: op1_06_in19 = reg_1100;
    70: op1_06_in19 = reg_0280;
    58: op1_06_in19 = reg_0413;
    48: op1_06_in19 = reg_0206;
    78: op1_06_in19 = reg_0158;
    46: op1_06_in19 = reg_0445;
    88: op1_06_in19 = reg_0681;
    79: op1_06_in19 = reg_0795;
    59: op1_06_in19 = reg_0802;
    80: op1_06_in19 = reg_0992;
    62: op1_06_in19 = reg_0709;
    52: op1_06_in19 = reg_0846;
    81: op1_06_in19 = imem02_in[11:8];
    63: op1_06_in19 = reg_0774;
    82: op1_06_in19 = reg_0026;
    89: op1_06_in19 = reg_0531;
    83: op1_06_in19 = reg_0039;
    64: op1_06_in19 = reg_0306;
    65: op1_06_in19 = imem05_in[11:8];
    90: op1_06_in19 = reg_0897;
    66: op1_06_in19 = reg_0521;
    91: op1_06_in19 = reg_0027;
    44: op1_06_in19 = reg_0565;
    67: op1_06_in19 = reg_0406;
    92: op1_06_in19 = reg_0143;
    93: op1_06_in19 = reg_0603;
    94: op1_06_in19 = reg_0336;
    95: op1_06_in19 = reg_1324;
    96: op1_06_in19 = reg_1065;
    42: op1_06_in19 = reg_0278;
    97: op1_06_in19 = reg_0340;
    98: op1_06_in19 = reg_0410;
    99: op1_06_in19 = reg_0902;
    100: op1_06_in19 = reg_0800;
    101: op1_06_in19 = reg_1455;
    102: op1_06_in19 = reg_0755;
    103: op1_06_in19 = reg_1414;
    104: op1_06_in19 = reg_0060;
    105: op1_06_in19 = reg_0211;
    106: op1_06_in19 = reg_0535;
    107: op1_06_in19 = reg_0798;
    108: op1_06_in19 = reg_0030;
    109: op1_06_in19 = reg_0135;
    110: op1_06_in19 = reg_0706;
    112: op1_06_in19 = reg_0560;
    113: op1_06_in19 = reg_0478;
    114: op1_06_in19 = reg_0334;
    116: op1_06_in19 = reg_0330;
    117: op1_06_in19 = imem01_in[7:4];
    118: op1_06_in19 = imem03_in[7:4];
    120: op1_06_in19 = reg_0420;
    121: op1_06_in19 = reg_0825;
    122: op1_06_in19 = reg_0859;
    123: op1_06_in19 = reg_0398;
    124: op1_06_in19 = reg_0996;
    125: op1_06_in19 = reg_0069;
    126: op1_06_in19 = reg_1168;
    127: op1_06_in19 = reg_0145;
    128: op1_06_in19 = reg_0631;
    130: op1_06_in19 = reg_1253;
    131: op1_06_in19 = reg_0624;
    default: op1_06_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_06_inv19 = 1;
    69: op1_06_inv19 = 1;
    71: op1_06_inv19 = 1;
    54: op1_06_inv19 = 1;
    68: op1_06_inv19 = 1;
    76: op1_06_inv19 = 1;
    60: op1_06_inv19 = 1;
    57: op1_06_inv19 = 1;
    58: op1_06_inv19 = 1;
    48: op1_06_inv19 = 1;
    78: op1_06_inv19 = 1;
    88: op1_06_inv19 = 1;
    80: op1_06_inv19 = 1;
    81: op1_06_inv19 = 1;
    63: op1_06_inv19 = 1;
    82: op1_06_inv19 = 1;
    90: op1_06_inv19 = 1;
    66: op1_06_inv19 = 1;
    93: op1_06_inv19 = 1;
    95: op1_06_inv19 = 1;
    97: op1_06_inv19 = 1;
    99: op1_06_inv19 = 1;
    100: op1_06_inv19 = 1;
    101: op1_06_inv19 = 1;
    104: op1_06_inv19 = 1;
    105: op1_06_inv19 = 1;
    110: op1_06_inv19 = 1;
    115: op1_06_inv19 = 1;
    118: op1_06_inv19 = 1;
    120: op1_06_inv19 = 1;
    122: op1_06_inv19 = 1;
    123: op1_06_inv19 = 1;
    124: op1_06_inv19 = 1;
    125: op1_06_inv19 = 1;
    126: op1_06_inv19 = 1;
    127: op1_06_inv19 = 1;
    128: op1_06_inv19 = 1;
    130: op1_06_inv19 = 1;
    131: op1_06_inv19 = 1;
    default: op1_06_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in20 = reg_1031;
    53: op1_06_in20 = imem05_in[11:8];
    55: op1_06_in20 = reg_0270;
    86: op1_06_in20 = imem04_in[11:8];
    73: op1_06_in20 = reg_0156;
    69: op1_06_in20 = reg_0220;
    71: op1_06_in20 = reg_0609;
    50: op1_06_in20 = reg_0415;
    54: op1_06_in20 = reg_0390;
    74: op1_06_in20 = reg_0071;
    68: op1_06_in20 = reg_0145;
    61: op1_06_in20 = reg_0788;
    85: op1_06_in20 = reg_0788;
    75: op1_06_in20 = reg_0549;
    87: op1_06_in20 = reg_0340;
    56: op1_06_in20 = reg_1170;
    76: op1_06_in20 = reg_0047;
    60: op1_06_in20 = reg_0596;
    57: op1_06_in20 = reg_0851;
    77: op1_06_in20 = reg_1254;
    70: op1_06_in20 = reg_0757;
    58: op1_06_in20 = reg_0623;
    48: op1_06_in20 = reg_0784;
    78: op1_06_in20 = reg_0924;
    46: op1_06_in20 = reg_0648;
    88: op1_06_in20 = reg_0796;
    79: op1_06_in20 = reg_0869;
    59: op1_06_in20 = reg_0313;
    80: op1_06_in20 = reg_0173;
    62: op1_06_in20 = reg_0710;
    52: op1_06_in20 = reg_0024;
    81: op1_06_in20 = imem02_in[15:12];
    63: op1_06_in20 = reg_0465;
    82: op1_06_in20 = reg_1255;
    89: op1_06_in20 = reg_0297;
    83: op1_06_in20 = reg_0195;
    64: op1_06_in20 = reg_0877;
    84: op1_06_in20 = reg_0824;
    65: op1_06_in20 = reg_0601;
    90: op1_06_in20 = reg_0695;
    66: op1_06_in20 = reg_0484;
    91: op1_06_in20 = imem01_in[3:0];
    44: op1_06_in20 = reg_0564;
    67: op1_06_in20 = reg_0969;
    92: op1_06_in20 = reg_0891;
    93: op1_06_in20 = reg_0864;
    94: op1_06_in20 = reg_0932;
    95: op1_06_in20 = reg_0917;
    96: op1_06_in20 = reg_0232;
    42: op1_06_in20 = reg_0042;
    97: op1_06_in20 = reg_0862;
    98: op1_06_in20 = reg_0060;
    99: op1_06_in20 = reg_0331;
    100: op1_06_in20 = reg_0007;
    101: op1_06_in20 = reg_0128;
    102: op1_06_in20 = reg_1058;
    121: op1_06_in20 = reg_1058;
    103: op1_06_in20 = reg_0461;
    104: op1_06_in20 = reg_0277;
    105: op1_06_in20 = reg_0904;
    106: op1_06_in20 = reg_0034;
    107: op1_06_in20 = reg_1475;
    108: op1_06_in20 = reg_0618;
    109: op1_06_in20 = reg_0309;
    110: op1_06_in20 = reg_0840;
    112: op1_06_in20 = reg_0802;
    113: op1_06_in20 = reg_0298;
    114: op1_06_in20 = reg_1403;
    115: op1_06_in20 = imem01_in[15:12];
    116: op1_06_in20 = reg_0597;
    117: op1_06_in20 = reg_1090;
    118: op1_06_in20 = reg_1145;
    119: op1_06_in20 = reg_0112;
    120: op1_06_in20 = reg_1488;
    122: op1_06_in20 = reg_1323;
    123: op1_06_in20 = reg_0374;
    124: op1_06_in20 = reg_1059;
    125: op1_06_in20 = imem03_in[7:4];
    126: op1_06_in20 = reg_0566;
    127: op1_06_in20 = reg_0143;
    128: op1_06_in20 = reg_0876;
    130: op1_06_in20 = reg_0875;
    131: op1_06_in20 = reg_0345;
    default: op1_06_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv20 = 1;
    53: op1_06_inv20 = 1;
    73: op1_06_inv20 = 1;
    69: op1_06_inv20 = 1;
    71: op1_06_inv20 = 1;
    74: op1_06_inv20 = 1;
    61: op1_06_inv20 = 1;
    75: op1_06_inv20 = 1;
    56: op1_06_inv20 = 1;
    76: op1_06_inv20 = 1;
    60: op1_06_inv20 = 1;
    77: op1_06_inv20 = 1;
    70: op1_06_inv20 = 1;
    58: op1_06_inv20 = 1;
    48: op1_06_inv20 = 1;
    80: op1_06_inv20 = 1;
    52: op1_06_inv20 = 1;
    81: op1_06_inv20 = 1;
    63: op1_06_inv20 = 1;
    89: op1_06_inv20 = 1;
    83: op1_06_inv20 = 1;
    67: op1_06_inv20 = 1;
    94: op1_06_inv20 = 1;
    96: op1_06_inv20 = 1;
    97: op1_06_inv20 = 1;
    98: op1_06_inv20 = 1;
    101: op1_06_inv20 = 1;
    102: op1_06_inv20 = 1;
    105: op1_06_inv20 = 1;
    106: op1_06_inv20 = 1;
    109: op1_06_inv20 = 1;
    114: op1_06_inv20 = 1;
    116: op1_06_inv20 = 1;
    117: op1_06_inv20 = 1;
    119: op1_06_inv20 = 1;
    120: op1_06_inv20 = 1;
    122: op1_06_inv20 = 1;
    123: op1_06_inv20 = 1;
    125: op1_06_inv20 = 1;
    126: op1_06_inv20 = 1;
    127: op1_06_inv20 = 1;
    128: op1_06_inv20 = 1;
    default: op1_06_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in21 = reg_0239;
    53: op1_06_in21 = imem05_in[15:12];
    55: op1_06_in21 = reg_0152;
    86: op1_06_in21 = reg_0252;
    73: op1_06_in21 = reg_0777;
    69: op1_06_in21 = reg_1226;
    71: op1_06_in21 = imem01_in[3:0];
    50: op1_06_in21 = reg_0413;
    54: op1_06_in21 = reg_0878;
    74: op1_06_in21 = reg_0203;
    68: op1_06_in21 = reg_1003;
    92: op1_06_in21 = reg_1003;
    61: op1_06_in21 = reg_1291;
    85: op1_06_in21 = reg_1291;
    75: op1_06_in21 = reg_0609;
    87: op1_06_in21 = reg_0420;
    56: op1_06_in21 = reg_0821;
    76: op1_06_in21 = reg_0553;
    60: op1_06_in21 = reg_0368;
    57: op1_06_in21 = reg_0157;
    77: op1_06_in21 = reg_0611;
    70: op1_06_in21 = reg_0756;
    58: op1_06_in21 = reg_0592;
    48: op1_06_in21 = imem06_in[11:8];
    78: op1_06_in21 = reg_0223;
    46: op1_06_in21 = reg_0566;
    88: op1_06_in21 = reg_1040;
    79: op1_06_in21 = reg_1505;
    59: op1_06_in21 = reg_0757;
    80: op1_06_in21 = reg_0567;
    62: op1_06_in21 = reg_0375;
    52: op1_06_in21 = reg_0217;
    81: op1_06_in21 = reg_1494;
    127: op1_06_in21 = reg_1494;
    63: op1_06_in21 = reg_0437;
    82: op1_06_in21 = reg_0463;
    89: op1_06_in21 = reg_1083;
    83: op1_06_in21 = imem06_in[15:12];
    64: op1_06_in21 = reg_0009;
    84: op1_06_in21 = reg_0381;
    65: op1_06_in21 = reg_0274;
    90: op1_06_in21 = reg_0327;
    91: op1_06_in21 = reg_1290;
    44: op1_06_in21 = reg_0182;
    67: op1_06_in21 = reg_0342;
    93: op1_06_in21 = reg_0828;
    94: op1_06_in21 = reg_0063;
    95: op1_06_in21 = reg_0355;
    96: op1_06_in21 = reg_0337;
    42: op1_06_in21 = reg_0013;
    97: op1_06_in21 = reg_0719;
    98: op1_06_in21 = reg_1322;
    99: op1_06_in21 = reg_0787;
    100: op1_06_in21 = reg_0999;
    101: op1_06_in21 = reg_0876;
    102: op1_06_in21 = reg_0906;
    103: op1_06_in21 = reg_1416;
    104: op1_06_in21 = reg_0788;
    117: op1_06_in21 = reg_0788;
    105: op1_06_in21 = reg_0117;
    106: op1_06_in21 = reg_0797;
    107: op1_06_in21 = reg_0966;
    108: op1_06_in21 = reg_0137;
    109: op1_06_in21 = reg_1350;
    110: op1_06_in21 = reg_0216;
    112: op1_06_in21 = reg_1098;
    113: op1_06_in21 = reg_0667;
    114: op1_06_in21 = reg_0940;
    115: op1_06_in21 = reg_0982;
    116: op1_06_in21 = reg_0198;
    118: op1_06_in21 = reg_0049;
    119: op1_06_in21 = reg_0106;
    120: op1_06_in21 = reg_0470;
    121: op1_06_in21 = reg_1035;
    122: op1_06_in21 = reg_0780;
    123: op1_06_in21 = reg_0585;
    124: op1_06_in21 = reg_0793;
    125: op1_06_in21 = reg_1145;
    126: op1_06_in21 = reg_0564;
    128: op1_06_in21 = reg_0745;
    130: op1_06_in21 = reg_0080;
    131: op1_06_in21 = reg_1228;
    default: op1_06_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv21 = 1;
    53: op1_06_inv21 = 1;
    69: op1_06_inv21 = 1;
    71: op1_06_inv21 = 1;
    50: op1_06_inv21 = 1;
    54: op1_06_inv21 = 1;
    74: op1_06_inv21 = 1;
    75: op1_06_inv21 = 1;
    87: op1_06_inv21 = 1;
    57: op1_06_inv21 = 1;
    77: op1_06_inv21 = 1;
    58: op1_06_inv21 = 1;
    48: op1_06_inv21 = 1;
    59: op1_06_inv21 = 1;
    52: op1_06_inv21 = 1;
    63: op1_06_inv21 = 1;
    82: op1_06_inv21 = 1;
    83: op1_06_inv21 = 1;
    64: op1_06_inv21 = 1;
    84: op1_06_inv21 = 1;
    90: op1_06_inv21 = 1;
    44: op1_06_inv21 = 1;
    93: op1_06_inv21 = 1;
    94: op1_06_inv21 = 1;
    95: op1_06_inv21 = 1;
    97: op1_06_inv21 = 1;
    100: op1_06_inv21 = 1;
    101: op1_06_inv21 = 1;
    103: op1_06_inv21 = 1;
    104: op1_06_inv21 = 1;
    105: op1_06_inv21 = 1;
    106: op1_06_inv21 = 1;
    107: op1_06_inv21 = 1;
    108: op1_06_inv21 = 1;
    109: op1_06_inv21 = 1;
    112: op1_06_inv21 = 1;
    113: op1_06_inv21 = 1;
    115: op1_06_inv21 = 1;
    116: op1_06_inv21 = 1;
    120: op1_06_inv21 = 1;
    122: op1_06_inv21 = 1;
    128: op1_06_inv21 = 1;
    default: op1_06_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in22 = reg_0241;
    75: op1_06_in22 = reg_0241;
    53: op1_06_in22 = reg_0333;
    44: op1_06_in22 = reg_0333;
    55: op1_06_in22 = reg_0213;
    86: op1_06_in22 = reg_0552;
    73: op1_06_in22 = reg_0029;
    78: op1_06_in22 = reg_0029;
    69: op1_06_in22 = reg_0885;
    71: op1_06_in22 = imem01_in[15:12];
    50: op1_06_in22 = reg_0103;
    54: op1_06_in22 = reg_0069;
    74: op1_06_in22 = reg_0122;
    68: op1_06_in22 = reg_0965;
    61: op1_06_in22 = reg_1255;
    87: op1_06_in22 = reg_1502;
    56: op1_06_in22 = reg_1096;
    76: op1_06_in22 = reg_0547;
    82: op1_06_in22 = reg_0547;
    60: op1_06_in22 = reg_0837;
    57: op1_06_in22 = reg_0621;
    77: op1_06_in22 = reg_0728;
    130: op1_06_in22 = reg_0728;
    70: op1_06_in22 = reg_0191;
    110: op1_06_in22 = reg_0191;
    58: op1_06_in22 = reg_0114;
    48: op1_06_in22 = reg_0908;
    46: op1_06_in22 = reg_0450;
    88: op1_06_in22 = reg_0452;
    79: op1_06_in22 = reg_1501;
    59: op1_06_in22 = reg_0734;
    80: op1_06_in22 = reg_1404;
    62: op1_06_in22 = reg_0177;
    52: op1_06_in22 = reg_0801;
    81: op1_06_in22 = reg_0233;
    63: op1_06_in22 = reg_0593;
    89: op1_06_in22 = reg_1215;
    83: op1_06_in22 = reg_0925;
    64: op1_06_in22 = reg_0830;
    84: op1_06_in22 = imem02_in[3:0];
    65: op1_06_in22 = reg_0575;
    114: op1_06_in22 = reg_0575;
    85: op1_06_in22 = reg_0277;
    90: op1_06_in22 = reg_0848;
    91: op1_06_in22 = reg_1291;
    67: op1_06_in22 = reg_0721;
    92: op1_06_in22 = reg_0957;
    93: op1_06_in22 = reg_0206;
    94: op1_06_in22 = reg_0095;
    95: op1_06_in22 = reg_1253;
    96: op1_06_in22 = reg_0211;
    42: op1_06_in22 = reg_0662;
    97: op1_06_in22 = reg_0016;
    98: op1_06_in22 = imem01_in[3:0];
    104: op1_06_in22 = imem01_in[3:0];
    99: op1_06_in22 = reg_0260;
    100: op1_06_in22 = reg_0699;
    101: op1_06_in22 = reg_0380;
    102: op1_06_in22 = reg_0397;
    103: op1_06_in22 = reg_0994;
    105: op1_06_in22 = reg_0209;
    106: op1_06_in22 = reg_1257;
    107: op1_06_in22 = reg_0147;
    108: op1_06_in22 = reg_0051;
    109: op1_06_in22 = reg_0157;
    112: op1_06_in22 = reg_0711;
    113: op1_06_in22 = reg_0894;
    115: op1_06_in22 = reg_0871;
    116: op1_06_in22 = reg_0847;
    117: op1_06_in22 = reg_1034;
    118: op1_06_in22 = reg_0444;
    119: op1_06_in22 = reg_0876;
    120: op1_06_in22 = reg_0370;
    121: op1_06_in22 = reg_0730;
    122: op1_06_in22 = reg_0109;
    123: op1_06_in22 = reg_0617;
    124: op1_06_in22 = reg_0045;
    125: op1_06_in22 = reg_0185;
    126: op1_06_in22 = reg_0697;
    127: op1_06_in22 = reg_0070;
    128: op1_06_in22 = reg_0897;
    131: op1_06_in22 = reg_0295;
    default: op1_06_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_06_inv22 = 1;
    50: op1_06_inv22 = 1;
    54: op1_06_inv22 = 1;
    68: op1_06_inv22 = 1;
    61: op1_06_inv22 = 1;
    75: op1_06_inv22 = 1;
    87: op1_06_inv22 = 1;
    56: op1_06_inv22 = 1;
    76: op1_06_inv22 = 1;
    57: op1_06_inv22 = 1;
    77: op1_06_inv22 = 1;
    46: op1_06_inv22 = 1;
    88: op1_06_inv22 = 1;
    80: op1_06_inv22 = 1;
    52: op1_06_inv22 = 1;
    81: op1_06_inv22 = 1;
    63: op1_06_inv22 = 1;
    89: op1_06_inv22 = 1;
    65: op1_06_inv22 = 1;
    44: op1_06_inv22 = 1;
    67: op1_06_inv22 = 1;
    94: op1_06_inv22 = 1;
    96: op1_06_inv22 = 1;
    97: op1_06_inv22 = 1;
    98: op1_06_inv22 = 1;
    99: op1_06_inv22 = 1;
    101: op1_06_inv22 = 1;
    102: op1_06_inv22 = 1;
    104: op1_06_inv22 = 1;
    109: op1_06_inv22 = 1;
    112: op1_06_inv22 = 1;
    114: op1_06_inv22 = 1;
    115: op1_06_inv22 = 1;
    116: op1_06_inv22 = 1;
    117: op1_06_inv22 = 1;
    121: op1_06_inv22 = 1;
    122: op1_06_inv22 = 1;
    123: op1_06_inv22 = 1;
    124: op1_06_inv22 = 1;
    125: op1_06_inv22 = 1;
    128: op1_06_inv22 = 1;
    130: op1_06_inv22 = 1;
    131: op1_06_inv22 = 1;
    default: op1_06_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in23 = reg_1473;
    53: op1_06_in23 = reg_0445;
    55: op1_06_in23 = reg_0017;
    86: op1_06_in23 = reg_1203;
    106: op1_06_in23 = reg_1203;
    73: op1_06_in23 = reg_0661;
    69: op1_06_in23 = reg_0573;
    100: op1_06_in23 = reg_0573;
    71: op1_06_in23 = reg_0469;
    50: op1_06_in23 = reg_0003;
    54: op1_06_in23 = reg_0801;
    128: op1_06_in23 = reg_0801;
    74: op1_06_in23 = reg_0005;
    68: op1_06_in23 = reg_0190;
    61: op1_06_in23 = reg_1256;
    75: op1_06_in23 = reg_0468;
    87: op1_06_in23 = reg_0832;
    56: op1_06_in23 = reg_0394;
    76: op1_06_in23 = reg_0222;
    77: op1_06_in23 = reg_0222;
    60: op1_06_in23 = reg_0097;
    57: op1_06_in23 = reg_0620;
    70: op1_06_in23 = reg_0830;
    58: op1_06_in23 = reg_0085;
    48: op1_06_in23 = reg_0905;
    78: op1_06_in23 = reg_0665;
    46: op1_06_in23 = reg_0070;
    88: op1_06_in23 = reg_1419;
    79: op1_06_in23 = reg_0115;
    59: op1_06_in23 = reg_0678;
    80: op1_06_in23 = reg_0794;
    62: op1_06_in23 = imem03_in[7:4];
    52: op1_06_in23 = reg_0800;
    84: op1_06_in23 = reg_0800;
    81: op1_06_in23 = reg_0154;
    63: op1_06_in23 = reg_0103;
    82: op1_06_in23 = reg_0260;
    89: op1_06_in23 = reg_1082;
    83: op1_06_in23 = reg_0974;
    64: op1_06_in23 = reg_0802;
    65: op1_06_in23 = reg_0602;
    85: op1_06_in23 = reg_1512;
    90: op1_06_in23 = reg_1091;
    91: op1_06_in23 = reg_0549;
    117: op1_06_in23 = reg_0549;
    44: op1_06_in23 = reg_0331;
    67: op1_06_in23 = reg_0470;
    92: op1_06_in23 = reg_1300;
    93: op1_06_in23 = reg_0038;
    94: op1_06_in23 = reg_0019;
    95: op1_06_in23 = reg_0785;
    96: op1_06_in23 = reg_0236;
    42: op1_06_in23 = reg_0256;
    97: op1_06_in23 = reg_0020;
    98: op1_06_in23 = reg_1031;
    99: op1_06_in23 = reg_0242;
    101: op1_06_in23 = reg_0306;
    102: op1_06_in23 = reg_0161;
    103: op1_06_in23 = reg_0135;
    113: op1_06_in23 = reg_0135;
    104: op1_06_in23 = imem01_in[15:12];
    105: op1_06_in23 = reg_0016;
    107: op1_06_in23 = reg_0386;
    108: op1_06_in23 = reg_0002;
    109: op1_06_in23 = reg_1094;
    110: op1_06_in23 = reg_0964;
    112: op1_06_in23 = reg_0294;
    114: op1_06_in23 = reg_0864;
    115: op1_06_in23 = reg_0985;
    116: op1_06_in23 = reg_0783;
    118: op1_06_in23 = reg_0261;
    119: op1_06_in23 = reg_0380;
    120: op1_06_in23 = imem05_in[15:12];
    121: op1_06_in23 = reg_0984;
    122: op1_06_in23 = reg_0716;
    123: op1_06_in23 = reg_0528;
    124: op1_06_in23 = reg_0697;
    125: op1_06_in23 = reg_0444;
    126: op1_06_in23 = reg_1403;
    127: op1_06_in23 = reg_1314;
    130: op1_06_in23 = reg_0043;
    131: op1_06_in23 = reg_0308;
    default: op1_06_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_06_inv23 = 1;
    71: op1_06_inv23 = 1;
    50: op1_06_inv23 = 1;
    54: op1_06_inv23 = 1;
    68: op1_06_inv23 = 1;
    61: op1_06_inv23 = 1;
    56: op1_06_inv23 = 1;
    76: op1_06_inv23 = 1;
    60: op1_06_inv23 = 1;
    57: op1_06_inv23 = 1;
    58: op1_06_inv23 = 1;
    78: op1_06_inv23 = 1;
    46: op1_06_inv23 = 1;
    59: op1_06_inv23 = 1;
    80: op1_06_inv23 = 1;
    62: op1_06_inv23 = 1;
    52: op1_06_inv23 = 1;
    81: op1_06_inv23 = 1;
    63: op1_06_inv23 = 1;
    89: op1_06_inv23 = 1;
    83: op1_06_inv23 = 1;
    64: op1_06_inv23 = 1;
    85: op1_06_inv23 = 1;
    44: op1_06_inv23 = 1;
    92: op1_06_inv23 = 1;
    93: op1_06_inv23 = 1;
    94: op1_06_inv23 = 1;
    95: op1_06_inv23 = 1;
    97: op1_06_inv23 = 1;
    100: op1_06_inv23 = 1;
    102: op1_06_inv23 = 1;
    103: op1_06_inv23 = 1;
    104: op1_06_inv23 = 1;
    105: op1_06_inv23 = 1;
    107: op1_06_inv23 = 1;
    109: op1_06_inv23 = 1;
    115: op1_06_inv23 = 1;
    123: op1_06_inv23 = 1;
    125: op1_06_inv23 = 1;
    126: op1_06_inv23 = 1;
    128: op1_06_inv23 = 1;
    130: op1_06_inv23 = 1;
    default: op1_06_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in24 = reg_0819;
    53: op1_06_in24 = reg_0173;
    55: op1_06_in24 = reg_0230;
    86: op1_06_in24 = reg_0281;
    64: op1_06_in24 = reg_0281;
    73: op1_06_in24 = reg_0366;
    78: op1_06_in24 = reg_0366;
    69: op1_06_in24 = reg_0426;
    71: op1_06_in24 = reg_0438;
    50: op1_06_in24 = reg_0052;
    54: op1_06_in24 = reg_0802;
    74: op1_06_in24 = reg_1290;
    68: op1_06_in24 = reg_0597;
    61: op1_06_in24 = reg_0549;
    75: op1_06_in24 = reg_0967;
    87: op1_06_in24 = imem05_in[3:0];
    56: op1_06_in24 = reg_0225;
    76: op1_06_in24 = reg_0609;
    60: op1_06_in24 = reg_0096;
    57: op1_06_in24 = reg_0103;
    77: op1_06_in24 = reg_1474;
    70: op1_06_in24 = reg_0377;
    58: op1_06_in24 = reg_1182;
    48: op1_06_in24 = reg_0960;
    46: op1_06_in24 = reg_0418;
    88: op1_06_in24 = reg_0368;
    79: op1_06_in24 = reg_0110;
    59: op1_06_in24 = reg_0121;
    80: op1_06_in24 = reg_1373;
    62: op1_06_in24 = reg_0180;
    52: op1_06_in24 = imem03_in[7:4];
    81: op1_06_in24 = reg_1447;
    63: op1_06_in24 = reg_0085;
    82: op1_06_in24 = reg_0830;
    89: op1_06_in24 = reg_0421;
    83: op1_06_in24 = reg_0397;
    84: op1_06_in24 = reg_0068;
    65: op1_06_in24 = reg_0151;
    85: op1_06_in24 = reg_0047;
    90: op1_06_in24 = reg_0217;
    91: op1_06_in24 = reg_0548;
    44: op1_06_in24 = reg_0541;
    67: op1_06_in24 = reg_0199;
    92: op1_06_in24 = reg_0048;
    93: op1_06_in24 = reg_0039;
    94: op1_06_in24 = reg_0470;
    95: op1_06_in24 = reg_0930;
    96: op1_06_in24 = reg_0095;
    42: op1_06_in24 = reg_0561;
    97: op1_06_in24 = reg_0204;
    98: op1_06_in24 = reg_1253;
    99: op1_06_in24 = reg_0239;
    100: op1_06_in24 = reg_0706;
    101: op1_06_in24 = reg_0560;
    102: op1_06_in24 = reg_0925;
    103: op1_06_in24 = reg_0703;
    104: op1_06_in24 = reg_0874;
    115: op1_06_in24 = reg_0874;
    105: op1_06_in24 = reg_1488;
    106: op1_06_in24 = reg_0574;
    107: op1_06_in24 = reg_0363;
    108: op1_06_in24 = reg_0087;
    109: op1_06_in24 = reg_0779;
    110: op1_06_in24 = reg_0142;
    112: op1_06_in24 = reg_1078;
    113: op1_06_in24 = reg_0309;
    114: op1_06_in24 = reg_0317;
    116: op1_06_in24 = reg_1517;
    117: op1_06_in24 = reg_0242;
    118: op1_06_in24 = reg_1425;
    119: op1_06_in24 = reg_0897;
    120: op1_06_in24 = reg_0538;
    121: op1_06_in24 = reg_0863;
    122: op1_06_in24 = reg_0714;
    123: op1_06_in24 = reg_0213;
    124: op1_06_in24 = reg_1070;
    125: op1_06_in24 = reg_0709;
    126: op1_06_in24 = reg_1401;
    127: op1_06_in24 = reg_0756;
    128: op1_06_in24 = reg_0253;
    130: op1_06_in24 = reg_0447;
    131: op1_06_in24 = reg_0371;
    default: op1_06_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_06_inv24 = 1;
    73: op1_06_inv24 = 1;
    74: op1_06_inv24 = 1;
    56: op1_06_inv24 = 1;
    76: op1_06_inv24 = 1;
    57: op1_06_inv24 = 1;
    77: op1_06_inv24 = 1;
    70: op1_06_inv24 = 1;
    58: op1_06_inv24 = 1;
    88: op1_06_inv24 = 1;
    52: op1_06_inv24 = 1;
    63: op1_06_inv24 = 1;
    82: op1_06_inv24 = 1;
    64: op1_06_inv24 = 1;
    84: op1_06_inv24 = 1;
    65: op1_06_inv24 = 1;
    85: op1_06_inv24 = 1;
    67: op1_06_inv24 = 1;
    92: op1_06_inv24 = 1;
    93: op1_06_inv24 = 1;
    95: op1_06_inv24 = 1;
    99: op1_06_inv24 = 1;
    101: op1_06_inv24 = 1;
    103: op1_06_inv24 = 1;
    104: op1_06_inv24 = 1;
    105: op1_06_inv24 = 1;
    106: op1_06_inv24 = 1;
    110: op1_06_inv24 = 1;
    113: op1_06_inv24 = 1;
    114: op1_06_inv24 = 1;
    115: op1_06_inv24 = 1;
    117: op1_06_inv24 = 1;
    118: op1_06_inv24 = 1;
    121: op1_06_inv24 = 1;
    122: op1_06_inv24 = 1;
    123: op1_06_inv24 = 1;
    125: op1_06_inv24 = 1;
    127: op1_06_inv24 = 1;
    128: op1_06_inv24 = 1;
    131: op1_06_inv24 = 1;
    default: op1_06_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in25 = reg_1456;
    53: op1_06_in25 = reg_0346;
    55: op1_06_in25 = reg_0491;
    86: op1_06_in25 = reg_1147;
    73: op1_06_in25 = reg_0740;
    78: op1_06_in25 = reg_0740;
    69: op1_06_in25 = reg_0427;
    71: op1_06_in25 = reg_1452;
    54: op1_06_in25 = reg_0758;
    74: op1_06_in25 = reg_0448;
    68: op1_06_in25 = reg_0048;
    61: op1_06_in25 = reg_0610;
    75: op1_06_in25 = reg_0968;
    87: op1_06_in25 = reg_0733;
    56: op1_06_in25 = reg_0224;
    76: op1_06_in25 = reg_0242;
    60: op1_06_in25 = reg_0095;
    57: op1_06_in25 = reg_0321;
    77: op1_06_in25 = reg_0715;
    70: op1_06_in25 = imem03_in[3:0];
    48: op1_06_in25 = reg_0866;
    46: op1_06_in25 = reg_0303;
    88: op1_06_in25 = reg_0836;
    79: op1_06_in25 = reg_0716;
    59: op1_06_in25 = reg_0378;
    80: op1_06_in25 = reg_0602;
    62: op1_06_in25 = reg_1000;
    90: op1_06_in25 = reg_1000;
    52: op1_06_in25 = imem03_in[11:8];
    81: op1_06_in25 = reg_0198;
    63: op1_06_in25 = reg_0086;
    82: op1_06_in25 = reg_0612;
    89: op1_06_in25 = reg_0412;
    83: op1_06_in25 = reg_1334;
    64: op1_06_in25 = reg_0276;
    130: op1_06_in25 = reg_0276;
    84: op1_06_in25 = reg_0311;
    65: op1_06_in25 = reg_1036;
    85: op1_06_in25 = reg_0093;
    95: op1_06_in25 = reg_0093;
    91: op1_06_in25 = reg_0609;
    44: op1_06_in25 = imem05_in[7:4];
    94: op1_06_in25 = imem05_in[7:4];
    67: op1_06_in25 = reg_0305;
    92: op1_06_in25 = reg_1199;
    93: op1_06_in25 = reg_1508;
    96: op1_06_in25 = reg_0016;
    42: op1_06_in25 = reg_0496;
    97: op1_06_in25 = reg_0315;
    98: op1_06_in25 = reg_0553;
    99: op1_06_in25 = reg_0238;
    117: op1_06_in25 = reg_0238;
    100: op1_06_in25 = reg_0330;
    101: op1_06_in25 = reg_0007;
    102: op1_06_in25 = reg_1420;
    103: op1_06_in25 = reg_0299;
    104: op1_06_in25 = reg_1290;
    105: op1_06_in25 = reg_0136;
    106: op1_06_in25 = reg_0681;
    107: op1_06_in25 = reg_0901;
    108: op1_06_in25 = reg_0483;
    109: op1_06_in25 = reg_0285;
    110: op1_06_in25 = reg_0957;
    112: op1_06_in25 = reg_0255;
    113: op1_06_in25 = reg_1347;
    114: op1_06_in25 = reg_0206;
    115: op1_06_in25 = reg_0576;
    116: op1_06_in25 = reg_0627;
    118: op1_06_in25 = reg_1033;
    119: op1_06_in25 = reg_0560;
    120: op1_06_in25 = reg_0832;
    121: op1_06_in25 = reg_1323;
    122: op1_06_in25 = reg_0373;
    123: op1_06_in25 = reg_0050;
    124: op1_06_in25 = reg_0302;
    125: op1_06_in25 = reg_0706;
    126: op1_06_in25 = reg_1404;
    127: op1_06_in25 = reg_0290;
    128: op1_06_in25 = reg_0217;
    131: op1_06_in25 = reg_0195;
    default: op1_06_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_06_inv25 = 1;
    73: op1_06_inv25 = 1;
    69: op1_06_inv25 = 1;
    54: op1_06_inv25 = 1;
    61: op1_06_inv25 = 1;
    75: op1_06_inv25 = 1;
    87: op1_06_inv25 = 1;
    76: op1_06_inv25 = 1;
    60: op1_06_inv25 = 1;
    57: op1_06_inv25 = 1;
    78: op1_06_inv25 = 1;
    88: op1_06_inv25 = 1;
    80: op1_06_inv25 = 1;
    52: op1_06_inv25 = 1;
    63: op1_06_inv25 = 1;
    82: op1_06_inv25 = 1;
    89: op1_06_inv25 = 1;
    65: op1_06_inv25 = 1;
    90: op1_06_inv25 = 1;
    91: op1_06_inv25 = 1;
    67: op1_06_inv25 = 1;
    93: op1_06_inv25 = 1;
    94: op1_06_inv25 = 1;
    95: op1_06_inv25 = 1;
    96: op1_06_inv25 = 1;
    97: op1_06_inv25 = 1;
    100: op1_06_inv25 = 1;
    103: op1_06_inv25 = 1;
    106: op1_06_inv25 = 1;
    107: op1_06_inv25 = 1;
    108: op1_06_inv25 = 1;
    110: op1_06_inv25 = 1;
    112: op1_06_inv25 = 1;
    114: op1_06_inv25 = 1;
    119: op1_06_inv25 = 1;
    121: op1_06_inv25 = 1;
    122: op1_06_inv25 = 1;
    123: op1_06_inv25 = 1;
    124: op1_06_inv25 = 1;
    125: op1_06_inv25 = 1;
    128: op1_06_inv25 = 1;
    130: op1_06_inv25 = 1;
    131: op1_06_inv25 = 1;
    default: op1_06_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in26 = reg_0385;
    53: op1_06_in26 = reg_0650;
    55: op1_06_in26 = reg_0821;
    86: op1_06_in26 = reg_0598;
    73: op1_06_in26 = reg_0738;
    78: op1_06_in26 = reg_0738;
    69: op1_06_in26 = reg_0247;
    71: op1_06_in26 = reg_0726;
    54: op1_06_in26 = reg_0757;
    74: op1_06_in26 = reg_1255;
    68: op1_06_in26 = reg_0885;
    61: op1_06_in26 = reg_0242;
    75: op1_06_in26 = reg_0401;
    104: op1_06_in26 = reg_0401;
    87: op1_06_in26 = reg_0648;
    56: op1_06_in26 = reg_0226;
    76: op1_06_in26 = reg_0966;
    60: op1_06_in26 = reg_0236;
    57: op1_06_in26 = reg_0085;
    77: op1_06_in26 = reg_0434;
    70: op1_06_in26 = reg_0177;
    48: op1_06_in26 = reg_0863;
    46: op1_06_in26 = reg_0301;
    88: op1_06_in26 = reg_0719;
    79: op1_06_in26 = reg_0714;
    59: op1_06_in26 = reg_0376;
    80: op1_06_in26 = reg_0449;
    62: op1_06_in26 = reg_0999;
    84: op1_06_in26 = reg_0999;
    52: op1_06_in26 = reg_0525;
    81: op1_06_in26 = reg_0378;
    63: op1_06_in26 = reg_0484;
    82: op1_06_in26 = reg_0468;
    89: op1_06_in26 = reg_1041;
    83: op1_06_in26 = reg_1505;
    64: op1_06_in26 = reg_1132;
    65: op1_06_in26 = reg_0754;
    85: op1_06_in26 = reg_0548;
    90: op1_06_in26 = reg_0759;
    91: op1_06_in26 = reg_0239;
    44: op1_06_in26 = reg_0367;
    120: op1_06_in26 = reg_0367;
    67: op1_06_in26 = reg_0835;
    92: op1_06_in26 = reg_1092;
    93: op1_06_in26 = reg_0931;
    94: op1_06_in26 = imem05_in[11:8];
    95: op1_06_in26 = reg_0746;
    96: op1_06_in26 = reg_0210;
    42: op1_06_in26 = reg_0475;
    97: op1_06_in26 = reg_0793;
    98: op1_06_in26 = reg_0093;
    99: op1_06_in26 = reg_1473;
    100: op1_06_in26 = reg_1447;
    101: op1_06_in26 = reg_0217;
    102: op1_06_in26 = reg_0782;
    103: op1_06_in26 = reg_0457;
    105: op1_06_in26 = reg_0332;
    106: op1_06_in26 = reg_0500;
    107: op1_06_in26 = reg_0875;
    108: op1_06_in26 = reg_0124;
    109: op1_06_in26 = reg_0739;
    110: op1_06_in26 = reg_0190;
    112: op1_06_in26 = reg_0632;
    113: op1_06_in26 = reg_0159;
    114: op1_06_in26 = reg_0825;
    115: op1_06_in26 = reg_0258;
    116: op1_06_in26 = reg_0558;
    117: op1_06_in26 = reg_0968;
    118: op1_06_in26 = reg_0198;
    119: op1_06_in26 = reg_0802;
    121: op1_06_in26 = reg_1179;
    122: op1_06_in26 = reg_0586;
    123: op1_06_in26 = reg_0169;
    124: op1_06_in26 = reg_0197;
    125: op1_06_in26 = reg_1033;
    126: op1_06_in26 = reg_0266;
    127: op1_06_in26 = reg_1208;
    128: op1_06_in26 = reg_0006;
    130: op1_06_in26 = imem02_in[11:8];
    131: op1_06_in26 = reg_0977;
    default: op1_06_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_06_inv26 = 1;
    55: op1_06_inv26 = 1;
    86: op1_06_inv26 = 1;
    73: op1_06_inv26 = 1;
    69: op1_06_inv26 = 1;
    71: op1_06_inv26 = 1;
    74: op1_06_inv26 = 1;
    75: op1_06_inv26 = 1;
    76: op1_06_inv26 = 1;
    77: op1_06_inv26 = 1;
    70: op1_06_inv26 = 1;
    48: op1_06_inv26 = 1;
    46: op1_06_inv26 = 1;
    79: op1_06_inv26 = 1;
    80: op1_06_inv26 = 1;
    62: op1_06_inv26 = 1;
    81: op1_06_inv26 = 1;
    89: op1_06_inv26 = 1;
    83: op1_06_inv26 = 1;
    64: op1_06_inv26 = 1;
    65: op1_06_inv26 = 1;
    67: op1_06_inv26 = 1;
    92: op1_06_inv26 = 1;
    95: op1_06_inv26 = 1;
    97: op1_06_inv26 = 1;
    98: op1_06_inv26 = 1;
    103: op1_06_inv26 = 1;
    105: op1_06_inv26 = 1;
    106: op1_06_inv26 = 1;
    108: op1_06_inv26 = 1;
    116: op1_06_inv26 = 1;
    118: op1_06_inv26 = 1;
    119: op1_06_inv26 = 1;
    120: op1_06_inv26 = 1;
    121: op1_06_inv26 = 1;
    122: op1_06_inv26 = 1;
    123: op1_06_inv26 = 1;
    125: op1_06_inv26 = 1;
    128: op1_06_inv26 = 1;
    130: op1_06_inv26 = 1;
    default: op1_06_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in27 = reg_0896;
    53: op1_06_in27 = reg_0996;
    55: op1_06_in27 = reg_1096;
    86: op1_06_in27 = reg_0599;
    73: op1_06_in27 = reg_0408;
    69: op1_06_in27 = reg_1339;
    71: op1_06_in27 = reg_0147;
    54: op1_06_in27 = reg_0710;
    74: op1_06_in27 = reg_1070;
    68: op1_06_in27 = reg_0507;
    61: op1_06_in27 = reg_0609;
    75: op1_06_in27 = reg_0595;
    87: op1_06_in27 = reg_0066;
    56: op1_06_in27 = reg_0245;
    76: op1_06_in27 = reg_1456;
    60: op1_06_in27 = reg_0209;
    57: op1_06_in27 = reg_0086;
    77: op1_06_in27 = reg_1452;
    70: op1_06_in27 = reg_0185;
    48: op1_06_in27 = reg_0671;
    78: op1_06_in27 = reg_0593;
    46: op1_06_in27 = reg_0873;
    88: op1_06_in27 = reg_0338;
    79: op1_06_in27 = reg_0637;
    59: op1_06_in27 = reg_0314;
    80: op1_06_in27 = reg_0206;
    62: op1_06_in27 = reg_0964;
    52: op1_06_in27 = reg_0216;
    81: op1_06_in27 = reg_0000;
    82: op1_06_in27 = reg_0149;
    89: op1_06_in27 = reg_0199;
    83: op1_06_in27 = reg_1504;
    64: op1_06_in27 = reg_0311;
    84: op1_06_in27 = reg_0559;
    65: op1_06_in27 = reg_0977;
    85: op1_06_in27 = reg_0742;
    90: op1_06_in27 = reg_0049;
    112: op1_06_in27 = reg_0049;
    91: op1_06_in27 = reg_0798;
    44: op1_06_in27 = reg_0888;
    67: op1_06_in27 = reg_0117;
    92: op1_06_in27 = reg_0178;
    93: op1_06_in27 = reg_0193;
    94: op1_06_in27 = reg_1430;
    95: op1_06_in27 = reg_0747;
    96: op1_06_in27 = reg_0035;
    42: op1_06_in27 = reg_0452;
    97: op1_06_in27 = reg_0347;
    98: op1_06_in27 = reg_0163;
    99: op1_06_in27 = reg_0430;
    100: op1_06_in27 = reg_1448;
    101: op1_06_in27 = reg_0009;
    102: op1_06_in27 = reg_0271;
    103: op1_06_in27 = reg_1350;
    104: op1_06_in27 = reg_0222;
    105: op1_06_in27 = reg_0272;
    106: op1_06_in27 = reg_1214;
    107: op1_06_in27 = reg_0727;
    109: op1_06_in27 = reg_0415;
    110: op1_06_in27 = reg_0448;
    113: op1_06_in27 = reg_0661;
    114: op1_06_in27 = imem06_in[15:12];
    115: op1_06_in27 = reg_0550;
    116: op1_06_in27 = reg_1226;
    117: op1_06_in27 = reg_0438;
    118: op1_06_in27 = reg_0600;
    119: op1_06_in27 = reg_1098;
    120: op1_06_in27 = reg_0466;
    121: op1_06_in27 = reg_0265;
    122: op1_06_in27 = reg_0619;
    123: op1_06_in27 = reg_0087;
    124: op1_06_in27 = reg_0799;
    125: op1_06_in27 = reg_0180;
    126: op1_06_in27 = reg_0418;
    127: op1_06_in27 = reg_0107;
    128: op1_06_in27 = reg_0378;
    130: op1_06_in27 = reg_0877;
    131: op1_06_in27 = reg_0046;
    default: op1_06_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_06_inv27 = 1;
    69: op1_06_inv27 = 1;
    54: op1_06_inv27 = 1;
    74: op1_06_inv27 = 1;
    61: op1_06_inv27 = 1;
    75: op1_06_inv27 = 1;
    87: op1_06_inv27 = 1;
    56: op1_06_inv27 = 1;
    76: op1_06_inv27 = 1;
    77: op1_06_inv27 = 1;
    70: op1_06_inv27 = 1;
    48: op1_06_inv27 = 1;
    78: op1_06_inv27 = 1;
    46: op1_06_inv27 = 1;
    59: op1_06_inv27 = 1;
    52: op1_06_inv27 = 1;
    82: op1_06_inv27 = 1;
    89: op1_06_inv27 = 1;
    84: op1_06_inv27 = 1;
    85: op1_06_inv27 = 1;
    44: op1_06_inv27 = 1;
    67: op1_06_inv27 = 1;
    93: op1_06_inv27 = 1;
    94: op1_06_inv27 = 1;
    95: op1_06_inv27 = 1;
    96: op1_06_inv27 = 1;
    97: op1_06_inv27 = 1;
    98: op1_06_inv27 = 1;
    101: op1_06_inv27 = 1;
    103: op1_06_inv27 = 1;
    106: op1_06_inv27 = 1;
    112: op1_06_inv27 = 1;
    114: op1_06_inv27 = 1;
    115: op1_06_inv27 = 1;
    119: op1_06_inv27 = 1;
    121: op1_06_inv27 = 1;
    123: op1_06_inv27 = 1;
    125: op1_06_inv27 = 1;
    126: op1_06_inv27 = 1;
    127: op1_06_inv27 = 1;
    128: op1_06_inv27 = 1;
    131: op1_06_inv27 = 1;
    default: op1_06_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in28 = reg_0080;
    53: op1_06_in28 = reg_0997;
    55: op1_06_in28 = reg_1056;
    86: op1_06_in28 = reg_1041;
    73: op1_06_in28 = reg_0004;
    69: op1_06_in28 = reg_0577;
    71: op1_06_in28 = reg_0402;
    54: op1_06_in28 = reg_0444;
    112: op1_06_in28 = reg_0444;
    74: op1_06_in28 = reg_1031;
    68: op1_06_in28 = imem03_in[11:8];
    61: op1_06_in28 = reg_0439;
    75: op1_06_in28 = reg_0457;
    87: op1_06_in28 = reg_0392;
    56: op1_06_in28 = reg_0893;
    76: op1_06_in28 = reg_0365;
    60: op1_06_in28 = reg_0062;
    57: op1_06_in28 = reg_0484;
    77: op1_06_in28 = reg_0146;
    70: op1_06_in28 = reg_0378;
    48: op1_06_in28 = reg_0617;
    78: op1_06_in28 = reg_0102;
    109: op1_06_in28 = reg_0102;
    46: op1_06_in28 = reg_0168;
    88: op1_06_in28 = reg_0336;
    79: op1_06_in28 = reg_0619;
    59: op1_06_in28 = reg_1149;
    80: op1_06_in28 = reg_0039;
    62: op1_06_in28 = reg_0113;
    127: op1_06_in28 = reg_0113;
    52: op1_06_in28 = reg_0198;
    81: op1_06_in28 = reg_0891;
    125: op1_06_in28 = reg_0891;
    82: op1_06_in28 = reg_0148;
    89: op1_06_in28 = reg_0033;
    83: op1_06_in28 = reg_1035;
    64: op1_06_in28 = reg_0227;
    84: op1_06_in28 = reg_0330;
    65: op1_06_in28 = imem06_in[15:12];
    85: op1_06_in28 = reg_1473;
    90: op1_06_in28 = reg_0557;
    91: op1_06_in28 = reg_0384;
    44: op1_06_in28 = reg_0090;
    67: op1_06_in28 = reg_0211;
    92: op1_06_in28 = reg_0025;
    93: op1_06_in28 = reg_0730;
    94: op1_06_in28 = reg_0347;
    95: op1_06_in28 = reg_0610;
    96: op1_06_in28 = reg_1169;
    42: op1_06_in28 = reg_0138;
    97: op1_06_in28 = reg_0733;
    98: op1_06_in28 = reg_0548;
    99: op1_06_in28 = reg_1452;
    100: op1_06_in28 = reg_1063;
    101: op1_06_in28 = reg_0279;
    102: op1_06_in28 = reg_1504;
    103: op1_06_in28 = reg_0224;
    104: op1_06_in28 = reg_0798;
    105: op1_06_in28 = reg_0205;
    106: op1_06_in28 = reg_0796;
    107: op1_06_in28 = reg_0335;
    110: op1_06_in28 = reg_0291;
    113: op1_06_in28 = reg_0663;
    114: op1_06_in28 = reg_1334;
    115: op1_06_in28 = reg_0787;
    116: op1_06_in28 = reg_1199;
    117: op1_06_in28 = reg_0403;
    118: op1_06_in28 = reg_0191;
    119: op1_06_in28 = reg_0800;
    120: op1_06_in28 = reg_0332;
    121: op1_06_in28 = reg_0780;
    122: op1_06_in28 = reg_0624;
    123: op1_06_in28 = reg_0157;
    124: op1_06_in28 = reg_0603;
    126: op1_06_in28 = reg_0872;
    128: op1_06_in28 = imem03_in[7:4];
    130: op1_06_in28 = reg_0423;
    131: op1_06_in28 = reg_0152;
    default: op1_06_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_06_inv28 = 1;
    55: op1_06_inv28 = 1;
    71: op1_06_inv28 = 1;
    54: op1_06_inv28 = 1;
    74: op1_06_inv28 = 1;
    75: op1_06_inv28 = 1;
    76: op1_06_inv28 = 1;
    70: op1_06_inv28 = 1;
    48: op1_06_inv28 = 1;
    78: op1_06_inv28 = 1;
    46: op1_06_inv28 = 1;
    88: op1_06_inv28 = 1;
    59: op1_06_inv28 = 1;
    64: op1_06_inv28 = 1;
    85: op1_06_inv28 = 1;
    91: op1_06_inv28 = 1;
    44: op1_06_inv28 = 1;
    93: op1_06_inv28 = 1;
    94: op1_06_inv28 = 1;
    96: op1_06_inv28 = 1;
    97: op1_06_inv28 = 1;
    98: op1_06_inv28 = 1;
    99: op1_06_inv28 = 1;
    101: op1_06_inv28 = 1;
    103: op1_06_inv28 = 1;
    104: op1_06_inv28 = 1;
    106: op1_06_inv28 = 1;
    107: op1_06_inv28 = 1;
    110: op1_06_inv28 = 1;
    112: op1_06_inv28 = 1;
    113: op1_06_inv28 = 1;
    114: op1_06_inv28 = 1;
    116: op1_06_inv28 = 1;
    118: op1_06_inv28 = 1;
    119: op1_06_inv28 = 1;
    120: op1_06_inv28 = 1;
    121: op1_06_inv28 = 1;
    124: op1_06_inv28 = 1;
    126: op1_06_inv28 = 1;
    130: op1_06_inv28 = 1;
    131: op1_06_inv28 = 1;
    default: op1_06_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in29 = reg_0079;
    107: op1_06_in29 = reg_0079;
    53: op1_06_in29 = reg_0567;
    55: op1_06_in29 = imem07_in[3:0];
    86: op1_06_in29 = reg_1004;
    73: op1_06_in29 = reg_0003;
    69: op1_06_in29 = reg_1065;
    71: op1_06_in29 = reg_0403;
    54: op1_06_in29 = reg_0377;
    74: op1_06_in29 = reg_0930;
    68: op1_06_in29 = imem03_in[15:12];
    61: op1_06_in29 = reg_0430;
    75: op1_06_in29 = reg_1103;
    87: op1_06_in29 = reg_0491;
    56: op1_06_in29 = reg_0170;
    76: op1_06_in29 = reg_0091;
    60: op1_06_in29 = reg_0016;
    57: op1_06_in29 = reg_0123;
    77: op1_06_in29 = reg_0899;
    70: op1_06_in29 = reg_1033;
    84: op1_06_in29 = reg_1033;
    48: op1_06_in29 = reg_0569;
    78: op1_06_in29 = reg_0361;
    46: op1_06_in29 = reg_0118;
    88: op1_06_in29 = reg_0633;
    79: op1_06_in29 = reg_0571;
    59: op1_06_in29 = reg_0349;
    80: op1_06_in29 = reg_0458;
    127: op1_06_in29 = reg_0458;
    62: op1_06_in29 = reg_0840;
    52: op1_06_in29 = reg_1091;
    81: op1_06_in29 = reg_0989;
    82: op1_06_in29 = reg_0400;
    89: op1_06_in29 = reg_0061;
    83: op1_06_in29 = reg_1228;
    64: op1_06_in29 = reg_0709;
    65: op1_06_in29 = reg_0730;
    85: op1_06_in29 = reg_1475;
    90: op1_06_in29 = reg_0198;
    112: op1_06_in29 = reg_0198;
    91: op1_06_in29 = reg_0362;
    44: op1_06_in29 = reg_0872;
    67: op1_06_in29 = reg_0064;
    92: op1_06_in29 = reg_0291;
    93: op1_06_in29 = imem06_in[11:8];
    94: op1_06_in29 = reg_0184;
    95: op1_06_in29 = reg_1474;
    104: op1_06_in29 = reg_1474;
    96: op1_06_in29 = reg_0986;
    42: op1_06_in29 = reg_0380;
    97: op1_06_in29 = reg_0176;
    98: op1_06_in29 = reg_0746;
    99: op1_06_in29 = reg_1456;
    100: op1_06_in29 = reg_0177;
    101: op1_06_in29 = reg_0006;
    102: op1_06_in29 = reg_0109;
    103: op1_06_in29 = reg_1094;
    105: op1_06_in29 = reg_0648;
    106: op1_06_in29 = reg_0471;
    109: op1_06_in29 = reg_0028;
    110: op1_06_in29 = reg_1282;
    113: op1_06_in29 = reg_0441;
    114: op1_06_in29 = reg_0960;
    115: op1_06_in29 = reg_0742;
    116: op1_06_in29 = reg_0541;
    117: op1_06_in29 = reg_0043;
    118: op1_06_in29 = reg_0556;
    119: op1_06_in29 = reg_0253;
    120: op1_06_in29 = reg_0392;
    121: op1_06_in29 = reg_1508;
    122: op1_06_in29 = reg_0528;
    123: op1_06_in29 = reg_0921;
    124: op1_06_in29 = reg_0565;
    125: op1_06_in29 = reg_1184;
    126: op1_06_in29 = reg_0318;
    128: op1_06_in29 = imem03_in[11:8];
    130: op1_06_in29 = reg_0588;
    131: op1_06_in29 = reg_0214;
    default: op1_06_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_06_inv29 = 1;
    86: op1_06_inv29 = 1;
    73: op1_06_inv29 = 1;
    71: op1_06_inv29 = 1;
    75: op1_06_inv29 = 1;
    87: op1_06_inv29 = 1;
    56: op1_06_inv29 = 1;
    60: op1_06_inv29 = 1;
    57: op1_06_inv29 = 1;
    70: op1_06_inv29 = 1;
    78: op1_06_inv29 = 1;
    46: op1_06_inv29 = 1;
    79: op1_06_inv29 = 1;
    59: op1_06_inv29 = 1;
    62: op1_06_inv29 = 1;
    81: op1_06_inv29 = 1;
    82: op1_06_inv29 = 1;
    64: op1_06_inv29 = 1;
    65: op1_06_inv29 = 1;
    91: op1_06_inv29 = 1;
    92: op1_06_inv29 = 1;
    94: op1_06_inv29 = 1;
    95: op1_06_inv29 = 1;
    96: op1_06_inv29 = 1;
    97: op1_06_inv29 = 1;
    98: op1_06_inv29 = 1;
    99: op1_06_inv29 = 1;
    100: op1_06_inv29 = 1;
    101: op1_06_inv29 = 1;
    102: op1_06_inv29 = 1;
    103: op1_06_inv29 = 1;
    104: op1_06_inv29 = 1;
    105: op1_06_inv29 = 1;
    107: op1_06_inv29 = 1;
    109: op1_06_inv29 = 1;
    110: op1_06_inv29 = 1;
    113: op1_06_inv29 = 1;
    114: op1_06_inv29 = 1;
    116: op1_06_inv29 = 1;
    117: op1_06_inv29 = 1;
    118: op1_06_inv29 = 1;
    119: op1_06_inv29 = 1;
    120: op1_06_inv29 = 1;
    121: op1_06_inv29 = 1;
    122: op1_06_inv29 = 1;
    123: op1_06_inv29 = 1;
    125: op1_06_inv29 = 1;
    126: op1_06_inv29 = 1;
    128: op1_06_inv29 = 1;
    130: op1_06_inv29 = 1;
    131: op1_06_inv29 = 1;
    default: op1_06_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_06_in30 = reg_0041;
    53: op1_06_in30 = reg_0565;
    55: op1_06_in30 = reg_0867;
    86: op1_06_in30 = reg_0342;
    73: op1_06_in30 = reg_0087;
    69: op1_06_in30 = reg_0396;
    71: op1_06_in30 = reg_0384;
    54: op1_06_in30 = reg_0025;
    74: op1_06_in30 = imem01_in[7:4];
    68: op1_06_in30 = reg_0840;
    61: op1_06_in30 = reg_0438;
    75: op1_06_in30 = reg_0532;
    87: op1_06_in30 = reg_0131;
    56: op1_06_in30 = reg_0921;
    76: op1_06_in30 = reg_0874;
    60: op1_06_in30 = reg_0034;
    77: op1_06_in30 = reg_0901;
    70: op1_06_in30 = reg_0640;
    48: op1_06_in30 = reg_0570;
    122: op1_06_in30 = reg_0570;
    78: op1_06_in30 = reg_0228;
    46: op1_06_in30 = reg_0240;
    88: op1_06_in30 = reg_0021;
    79: op1_06_in30 = reg_1225;
    59: op1_06_in30 = reg_0233;
    80: op1_06_in30 = reg_0751;
    62: op1_06_in30 = reg_0411;
    52: op1_06_in30 = reg_1064;
    81: op1_06_in30 = reg_0964;
    125: op1_06_in30 = reg_0964;
    82: op1_06_in30 = reg_0724;
    89: op1_06_in30 = reg_0698;
    83: op1_06_in30 = reg_0171;
    64: op1_06_in30 = reg_0235;
    84: op1_06_in30 = reg_0707;
    65: op1_06_in30 = reg_0172;
    85: op1_06_in30 = reg_0572;
    104: op1_06_in30 = reg_0572;
    90: op1_06_in30 = reg_1001;
    91: op1_06_in30 = reg_0365;
    44: op1_06_in30 = reg_0038;
    67: op1_06_in30 = reg_0019;
    92: op1_06_in30 = reg_0313;
    93: op1_06_in30 = reg_1467;
    94: op1_06_in30 = reg_0251;
    95: op1_06_in30 = reg_0715;
    96: op1_06_in30 = reg_1268;
    42: op1_06_in30 = reg_0343;
    97: op1_06_in30 = reg_0648;
    98: op1_06_in30 = reg_0787;
    99: op1_06_in30 = reg_0147;
    100: op1_06_in30 = reg_0198;
    101: op1_06_in30 = reg_1515;
    102: op1_06_in30 = reg_0714;
    121: op1_06_in30 = reg_0714;
    103: op1_06_in30 = reg_0665;
    105: op1_06_in30 = reg_0649;
    106: op1_06_in30 = reg_0537;
    107: op1_06_in30 = reg_0257;
    109: op1_06_in30 = reg_0002;
    110: op1_06_in30 = reg_0348;
    112: op1_06_in30 = reg_0078;
    113: op1_06_in30 = reg_0741;
    114: op1_06_in30 = reg_0271;
    115: op1_06_in30 = reg_1475;
    116: op1_06_in30 = reg_0218;
    117: op1_06_in30 = reg_0099;
    118: op1_06_in30 = reg_0965;
    119: op1_06_in30 = reg_1078;
    120: op1_06_in30 = reg_0566;
    123: op1_06_in30 = reg_1094;
    124: op1_06_in30 = reg_0270;
    126: op1_06_in30 = reg_0794;
    127: op1_06_in30 = reg_0427;
    128: op1_06_in30 = imem03_in[15:12];
    130: op1_06_in30 = reg_0934;
    131: op1_06_in30 = reg_0213;
    default: op1_06_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_06_inv30 = 1;
    69: op1_06_inv30 = 1;
    71: op1_06_inv30 = 1;
    54: op1_06_inv30 = 1;
    68: op1_06_inv30 = 1;
    75: op1_06_inv30 = 1;
    87: op1_06_inv30 = 1;
    56: op1_06_inv30 = 1;
    60: op1_06_inv30 = 1;
    77: op1_06_inv30 = 1;
    70: op1_06_inv30 = 1;
    78: op1_06_inv30 = 1;
    46: op1_06_inv30 = 1;
    59: op1_06_inv30 = 1;
    62: op1_06_inv30 = 1;
    81: op1_06_inv30 = 1;
    89: op1_06_inv30 = 1;
    83: op1_06_inv30 = 1;
    44: op1_06_inv30 = 1;
    67: op1_06_inv30 = 1;
    92: op1_06_inv30 = 1;
    93: op1_06_inv30 = 1;
    94: op1_06_inv30 = 1;
    95: op1_06_inv30 = 1;
    101: op1_06_inv30 = 1;
    103: op1_06_inv30 = 1;
    104: op1_06_inv30 = 1;
    106: op1_06_inv30 = 1;
    107: op1_06_inv30 = 1;
    110: op1_06_inv30 = 1;
    112: op1_06_inv30 = 1;
    115: op1_06_inv30 = 1;
    119: op1_06_inv30 = 1;
    120: op1_06_inv30 = 1;
    121: op1_06_inv30 = 1;
    122: op1_06_inv30 = 1;
    124: op1_06_inv30 = 1;
    125: op1_06_inv30 = 1;
    131: op1_06_inv30 = 1;
    default: op1_06_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_06_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#6の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_06_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in00 = reg_0613;
    53: op1_07_in00 = reg_0717;
    55: op1_07_in00 = reg_0207;
    86: op1_07_in00 = imem02_in[15:12];
    69: op1_07_in00 = reg_1064;
    73: op1_07_in00 = reg_0862;
    49: op1_07_in00 = reg_0298;
    50: op1_07_in00 = reg_0615;
    54: op1_07_in00 = reg_0819;
    71: op1_07_in00 = reg_0555;
    74: op1_07_in00 = reg_0183;
    68: op1_07_in00 = reg_0000;
    84: op1_07_in00 = reg_0000;
    75: op1_07_in00 = reg_1485;
    61: op1_07_in00 = reg_0616;
    56: op1_07_in00 = reg_0554;
    87: op1_07_in00 = reg_0480;
    76: op1_07_in00 = reg_0567;
    57: op1_07_in00 = reg_0438;
    77: op1_07_in00 = reg_1503;
    33: op1_07_in00 = imem07_in[3:0];
    40: op1_07_in00 = imem07_in[3:0];
    60: op1_07_in00 = reg_0876;
    58: op1_07_in00 = reg_1202;
    78: op1_07_in00 = reg_1502;
    70: op1_07_in00 = reg_0831;
    46: op1_07_in00 = reg_0563;
    51: op1_07_in00 = reg_0135;
    88: op1_07_in00 = reg_1078;
    91: op1_07_in00 = reg_1078;
    79: op1_07_in00 = reg_0095;
    59: op1_07_in00 = reg_0585;
    48: op1_07_in00 = reg_0932;
    80: op1_07_in00 = reg_0960;
    62: op1_07_in00 = reg_0240;
    52: op1_07_in00 = reg_0192;
    81: op1_07_in00 = reg_1404;
    63: op1_07_in00 = reg_1065;
    82: op1_07_in00 = reg_0290;
    89: op1_07_in00 = reg_0198;
    28: op1_07_in00 = imem07_in[15:12];
    22: op1_07_in00 = imem07_in[15:12];
    83: op1_07_in00 = reg_1490;
    123: op1_07_in00 = reg_1490;
    64: op1_07_in00 = reg_0378;
    65: op1_07_in00 = reg_0215;
    85: op1_07_in00 = reg_1488;
    37: op1_07_in00 = reg_0529;
    121: op1_07_in00 = reg_0529;
    90: op1_07_in00 = reg_0783;
    66: op1_07_in00 = reg_0249;
    47: op1_07_in00 = reg_0924;
    67: op1_07_in00 = reg_0374;
    92: op1_07_in00 = reg_0541;
    93: op1_07_in00 = reg_0720;
    94: op1_07_in00 = reg_0700;
    95: op1_07_in00 = reg_0149;
    44: op1_07_in00 = reg_0337;
    96: op1_07_in00 = reg_0604;
    97: op1_07_in00 = reg_0392;
    98: op1_07_in00 = reg_0609;
    99: op1_07_in00 = reg_0146;
    100: op1_07_in00 = reg_1184;
    101: op1_07_in00 = imem03_in[11:8];
    102: op1_07_in00 = reg_1302;
    103: op1_07_in00 = imem00_in[7:4];
    104: op1_07_in00 = reg_0968;
    105: op1_07_in00 = reg_0319;
    111: op1_07_in00 = reg_0319;
    106: op1_07_in00 = reg_0320;
    107: op1_07_in00 = reg_0447;
    108: op1_07_in00 = reg_1243;
    109: op1_07_in00 = reg_0843;
    110: op1_07_in00 = imem04_in[15:12];
    112: op1_07_in00 = reg_0600;
    34: op1_07_in00 = reg_0404;
    113: op1_07_in00 = reg_1242;
    114: op1_07_in00 = reg_0984;
    115: op1_07_in00 = reg_0434;
    116: op1_07_in00 = reg_0673;
    38: op1_07_in00 = reg_0740;
    117: op1_07_in00 = reg_0933;
    118: op1_07_in00 = reg_0142;
    119: op1_07_in00 = reg_0963;
    42: op1_07_in00 = reg_0238;
    120: op1_07_in00 = reg_0926;
    122: op1_07_in00 = reg_0345;
    124: op1_07_in00 = reg_0133;
    125: op1_07_in00 = reg_1516;
    126: op1_07_in00 = reg_0888;
    127: op1_07_in00 = reg_0181;
    128: op1_07_in00 = reg_0233;
    129: op1_07_in00 = imem00_in[15:12];
    130: op1_07_in00 = reg_0390;
    131: op1_07_in00 = reg_0051;
    default: op1_07_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_07_inv00 = 1;
    73: op1_07_inv00 = 1;
    50: op1_07_inv00 = 1;
    71: op1_07_inv00 = 1;
    74: op1_07_inv00 = 1;
    75: op1_07_inv00 = 1;
    57: op1_07_inv00 = 1;
    77: op1_07_inv00 = 1;
    60: op1_07_inv00 = 1;
    79: op1_07_inv00 = 1;
    59: op1_07_inv00 = 1;
    80: op1_07_inv00 = 1;
    62: op1_07_inv00 = 1;
    52: op1_07_inv00 = 1;
    81: op1_07_inv00 = 1;
    89: op1_07_inv00 = 1;
    64: op1_07_inv00 = 1;
    85: op1_07_inv00 = 1;
    90: op1_07_inv00 = 1;
    47: op1_07_inv00 = 1;
    92: op1_07_inv00 = 1;
    93: op1_07_inv00 = 1;
    94: op1_07_inv00 = 1;
    95: op1_07_inv00 = 1;
    44: op1_07_inv00 = 1;
    96: op1_07_inv00 = 1;
    97: op1_07_inv00 = 1;
    100: op1_07_inv00 = 1;
    101: op1_07_inv00 = 1;
    102: op1_07_inv00 = 1;
    103: op1_07_inv00 = 1;
    104: op1_07_inv00 = 1;
    106: op1_07_inv00 = 1;
    111: op1_07_inv00 = 1;
    112: op1_07_inv00 = 1;
    34: op1_07_inv00 = 1;
    113: op1_07_inv00 = 1;
    114: op1_07_inv00 = 1;
    115: op1_07_inv00 = 1;
    116: op1_07_inv00 = 1;
    38: op1_07_inv00 = 1;
    119: op1_07_inv00 = 1;
    42: op1_07_inv00 = 1;
    120: op1_07_inv00 = 1;
    122: op1_07_inv00 = 1;
    123: op1_07_inv00 = 1;
    124: op1_07_inv00 = 1;
    126: op1_07_inv00 = 1;
    127: op1_07_inv00 = 1;
    129: op1_07_inv00 = 1;
    131: op1_07_inv00 = 1;
    default: op1_07_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in01 = reg_0866;
    53: op1_07_in01 = reg_0634;
    55: op1_07_in01 = reg_1030;
    86: op1_07_in01 = reg_0745;
    69: op1_07_in01 = imem03_in[11:8];
    73: op1_07_in01 = reg_0835;
    49: op1_07_in01 = reg_0309;
    50: op1_07_in01 = reg_0219;
    54: op1_07_in01 = reg_0728;
    71: op1_07_in01 = reg_0842;
    74: op1_07_in01 = reg_0240;
    68: op1_07_in01 = reg_0891;
    84: op1_07_in01 = reg_0891;
    75: op1_07_in01 = reg_0449;
    61: op1_07_in01 = reg_0791;
    56: op1_07_in01 = reg_1099;
    87: op1_07_in01 = reg_0025;
    76: op1_07_in01 = reg_0697;
    57: op1_07_in01 = reg_0149;
    77: op1_07_in01 = reg_0019;
    79: op1_07_in01 = reg_0019;
    33: op1_07_in01 = imem07_in[15:12];
    60: op1_07_in01 = reg_0154;
    58: op1_07_in01 = reg_0271;
    78: op1_07_in01 = reg_0630;
    70: op1_07_in01 = reg_0694;
    46: op1_07_in01 = reg_0561;
    51: op1_07_in01 = reg_0998;
    88: op1_07_in01 = reg_0279;
    59: op1_07_in01 = reg_0569;
    48: op1_07_in01 = reg_0452;
    80: op1_07_in01 = reg_1326;
    62: op1_07_in01 = reg_0274;
    52: op1_07_in01 = reg_0730;
    81: op1_07_in01 = reg_0986;
    63: op1_07_in01 = reg_0406;
    82: op1_07_in01 = reg_0042;
    89: op1_07_in01 = reg_1001;
    83: op1_07_in01 = reg_1244;
    64: op1_07_in01 = reg_0377;
    65: op1_07_in01 = reg_0018;
    85: op1_07_in01 = reg_0470;
    37: op1_07_in01 = reg_0527;
    121: op1_07_in01 = reg_0527;
    90: op1_07_in01 = reg_0823;
    66: op1_07_in01 = reg_1230;
    91: op1_07_in01 = reg_1006;
    47: op1_07_in01 = reg_0490;
    67: op1_07_in01 = reg_0619;
    92: op1_07_in01 = reg_1009;
    93: op1_07_in01 = reg_0859;
    94: op1_07_in01 = reg_0992;
    40: op1_07_in01 = reg_0140;
    95: op1_07_in01 = reg_0148;
    44: op1_07_in01 = reg_0094;
    96: op1_07_in01 = reg_0391;
    97: op1_07_in01 = reg_0564;
    98: op1_07_in01 = reg_0612;
    99: op1_07_in01 = reg_0868;
    100: op1_07_in01 = reg_0070;
    101: op1_07_in01 = reg_0699;
    102: op1_07_in01 = reg_0141;
    103: op1_07_in01 = reg_0824;
    104: op1_07_in01 = reg_0439;
    105: op1_07_in01 = reg_1281;
    106: op1_07_in01 = reg_0698;
    107: op1_07_in01 = reg_0530;
    108: op1_07_in01 = reg_0983;
    109: op1_07_in01 = reg_1278;
    110: op1_07_in01 = reg_0507;
    111: op1_07_in01 = reg_0672;
    112: op1_07_in01 = reg_0311;
    34: op1_07_in01 = reg_0623;
    113: op1_07_in01 = reg_0725;
    120: op1_07_in01 = reg_0725;
    114: op1_07_in01 = reg_1467;
    115: op1_07_in01 = reg_0386;
    116: op1_07_in01 = reg_1282;
    38: op1_07_in01 = reg_0618;
    22: op1_07_in01 = reg_0001;
    117: op1_07_in01 = imem02_in[15:12];
    118: op1_07_in01 = reg_0349;
    119: op1_07_in01 = reg_0376;
    42: op1_07_in01 = reg_0727;
    122: op1_07_in01 = reg_1225;
    123: op1_07_in01 = reg_0554;
    124: op1_07_in01 = reg_0974;
    125: op1_07_in01 = reg_1518;
    126: op1_07_in01 = reg_0197;
    127: op1_07_in01 = reg_1339;
    128: op1_07_in01 = reg_0479;
    129: op1_07_in01 = reg_1081;
    130: op1_07_in01 = reg_0497;
    131: op1_07_in01 = reg_0156;
    default: op1_07_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_07_inv01 = 1;
    55: op1_07_inv01 = 1;
    86: op1_07_inv01 = 1;
    69: op1_07_inv01 = 1;
    50: op1_07_inv01 = 1;
    54: op1_07_inv01 = 1;
    68: op1_07_inv01 = 1;
    87: op1_07_inv01 = 1;
    76: op1_07_inv01 = 1;
    57: op1_07_inv01 = 1;
    77: op1_07_inv01 = 1;
    58: op1_07_inv01 = 1;
    78: op1_07_inv01 = 1;
    70: op1_07_inv01 = 1;
    51: op1_07_inv01 = 1;
    88: op1_07_inv01 = 1;
    62: op1_07_inv01 = 1;
    52: op1_07_inv01 = 1;
    81: op1_07_inv01 = 1;
    63: op1_07_inv01 = 1;
    82: op1_07_inv01 = 1;
    89: op1_07_inv01 = 1;
    83: op1_07_inv01 = 1;
    65: op1_07_inv01 = 1;
    85: op1_07_inv01 = 1;
    90: op1_07_inv01 = 1;
    67: op1_07_inv01 = 1;
    92: op1_07_inv01 = 1;
    93: op1_07_inv01 = 1;
    40: op1_07_inv01 = 1;
    95: op1_07_inv01 = 1;
    44: op1_07_inv01 = 1;
    96: op1_07_inv01 = 1;
    97: op1_07_inv01 = 1;
    99: op1_07_inv01 = 1;
    101: op1_07_inv01 = 1;
    102: op1_07_inv01 = 1;
    105: op1_07_inv01 = 1;
    106: op1_07_inv01 = 1;
    107: op1_07_inv01 = 1;
    110: op1_07_inv01 = 1;
    111: op1_07_inv01 = 1;
    34: op1_07_inv01 = 1;
    113: op1_07_inv01 = 1;
    22: op1_07_inv01 = 1;
    117: op1_07_inv01 = 1;
    122: op1_07_inv01 = 1;
    125: op1_07_inv01 = 1;
    126: op1_07_inv01 = 1;
    127: op1_07_inv01 = 1;
    129: op1_07_inv01 = 1;
    131: op1_07_inv01 = 1;
    default: op1_07_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in02 = reg_1277;
    53: op1_07_in02 = reg_0635;
    55: op1_07_in02 = reg_1036;
    86: op1_07_in02 = reg_0897;
    69: op1_07_in02 = reg_0261;
    73: op1_07_in02 = reg_0095;
    49: op1_07_in02 = imem07_in[3:0];
    47: op1_07_in02 = imem07_in[3:0];
    50: op1_07_in02 = reg_0580;
    54: op1_07_in02 = reg_0148;
    71: op1_07_in02 = reg_1243;
    74: op1_07_in02 = reg_1348;
    68: op1_07_in02 = reg_1003;
    128: op1_07_in02 = reg_1003;
    75: op1_07_in02 = reg_0151;
    61: op1_07_in02 = reg_1081;
    56: op1_07_in02 = reg_1080;
    87: op1_07_in02 = reg_1325;
    76: op1_07_in02 = reg_1401;
    57: op1_07_in02 = reg_0384;
    77: op1_07_in02 = reg_0578;
    33: op1_07_in02 = reg_0593;
    60: op1_07_in02 = reg_0830;
    58: op1_07_in02 = reg_0023;
    78: op1_07_in02 = reg_0736;
    70: op1_07_in02 = reg_1384;
    46: op1_07_in02 = reg_0531;
    51: op1_07_in02 = reg_0223;
    88: op1_07_in02 = imem03_in[11:8];
    79: op1_07_in02 = imem05_in[15:12];
    59: op1_07_in02 = reg_0570;
    48: op1_07_in02 = reg_0904;
    80: op1_07_in02 = reg_0160;
    62: op1_07_in02 = reg_0275;
    52: op1_07_in02 = reg_0866;
    81: op1_07_in02 = reg_0318;
    63: op1_07_in02 = reg_0407;
    82: op1_07_in02 = reg_0456;
    89: op1_07_in02 = reg_0000;
    83: op1_07_in02 = reg_1241;
    64: op1_07_in02 = reg_0143;
    84: op1_07_in02 = reg_0989;
    65: op1_07_in02 = reg_0191;
    90: op1_07_in02 = reg_0191;
    85: op1_07_in02 = reg_0735;
    37: op1_07_in02 = reg_0171;
    66: op1_07_in02 = reg_0987;
    91: op1_07_in02 = reg_1091;
    67: op1_07_in02 = reg_0528;
    92: op1_07_in02 = reg_1139;
    93: op1_07_in02 = reg_0752;
    94: op1_07_in02 = reg_0391;
    40: op1_07_in02 = reg_0621;
    34: op1_07_in02 = reg_0621;
    95: op1_07_in02 = reg_0402;
    44: op1_07_in02 = reg_0236;
    96: op1_07_in02 = reg_1104;
    97: op1_07_in02 = reg_0334;
    98: op1_07_in02 = reg_1474;
    99: op1_07_in02 = reg_0383;
    100: op1_07_in02 = reg_1313;
    101: op1_07_in02 = reg_0706;
    102: op1_07_in02 = reg_1228;
    103: op1_07_in02 = reg_0486;
    104: op1_07_in02 = reg_1457;
    105: op1_07_in02 = reg_1141;
    106: op1_07_in02 = reg_1143;
    107: op1_07_in02 = reg_0138;
    108: op1_07_in02 = reg_0638;
    109: op1_07_in02 = reg_0841;
    110: op1_07_in02 = reg_0252;
    111: op1_07_in02 = reg_1099;
    112: op1_07_in02 = reg_0234;
    113: op1_07_in02 = reg_1281;
    114: op1_07_in02 = reg_0859;
    115: op1_07_in02 = reg_0091;
    116: op1_07_in02 = reg_0348;
    38: op1_07_in02 = reg_0620;
    22: op1_07_in02 = reg_0004;
    117: op1_07_in02 = reg_0455;
    118: op1_07_in02 = reg_0954;
    119: op1_07_in02 = imem03_in[7:4];
    42: op1_07_in02 = reg_0453;
    120: op1_07_in02 = reg_1052;
    121: op1_07_in02 = reg_0295;
    122: op1_07_in02 = reg_0296;
    123: op1_07_in02 = reg_0523;
    124: op1_07_in02 = reg_0782;
    125: op1_07_in02 = reg_0505;
    126: op1_07_in02 = reg_1373;
    127: op1_07_in02 = imem04_in[7:4];
    129: op1_07_in02 = reg_0983;
    130: op1_07_in02 = reg_0326;
    131: op1_07_in02 = reg_0298;
    default: op1_07_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv02 = 1;
    86: op1_07_inv02 = 1;
    69: op1_07_inv02 = 1;
    73: op1_07_inv02 = 1;
    54: op1_07_inv02 = 1;
    75: op1_07_inv02 = 1;
    61: op1_07_inv02 = 1;
    87: op1_07_inv02 = 1;
    76: op1_07_inv02 = 1;
    33: op1_07_inv02 = 1;
    58: op1_07_inv02 = 1;
    78: op1_07_inv02 = 1;
    70: op1_07_inv02 = 1;
    80: op1_07_inv02 = 1;
    63: op1_07_inv02 = 1;
    82: op1_07_inv02 = 1;
    89: op1_07_inv02 = 1;
    84: op1_07_inv02 = 1;
    65: op1_07_inv02 = 1;
    85: op1_07_inv02 = 1;
    37: op1_07_inv02 = 1;
    90: op1_07_inv02 = 1;
    67: op1_07_inv02 = 1;
    92: op1_07_inv02 = 1;
    93: op1_07_inv02 = 1;
    94: op1_07_inv02 = 1;
    40: op1_07_inv02 = 1;
    97: op1_07_inv02 = 1;
    98: op1_07_inv02 = 1;
    101: op1_07_inv02 = 1;
    104: op1_07_inv02 = 1;
    105: op1_07_inv02 = 1;
    107: op1_07_inv02 = 1;
    109: op1_07_inv02 = 1;
    110: op1_07_inv02 = 1;
    111: op1_07_inv02 = 1;
    114: op1_07_inv02 = 1;
    115: op1_07_inv02 = 1;
    116: op1_07_inv02 = 1;
    38: op1_07_inv02 = 1;
    118: op1_07_inv02 = 1;
    119: op1_07_inv02 = 1;
    120: op1_07_inv02 = 1;
    124: op1_07_inv02 = 1;
    126: op1_07_inv02 = 1;
    129: op1_07_inv02 = 1;
    131: op1_07_inv02 = 1;
    default: op1_07_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in03 = reg_1279;
    53: op1_07_in03 = reg_0636;
    55: op1_07_in03 = reg_0974;
    86: op1_07_in03 = reg_0802;
    69: op1_07_in03 = reg_0964;
    64: op1_07_in03 = reg_0964;
    73: op1_07_in03 = reg_0117;
    49: op1_07_in03 = reg_0169;
    50: op1_07_in03 = reg_0554;
    54: op1_07_in03 = reg_0146;
    71: op1_07_in03 = imem00_in[7:4];
    74: op1_07_in03 = reg_0602;
    68: op1_07_in03 = reg_0963;
    75: op1_07_in03 = reg_0207;
    61: op1_07_in03 = reg_1052;
    56: op1_07_in03 = reg_0824;
    87: op1_07_in03 = reg_0425;
    76: op1_07_in03 = reg_0540;
    57: op1_07_in03 = reg_0385;
    77: op1_07_in03 = reg_0750;
    33: op1_07_in03 = reg_0592;
    40: op1_07_in03 = reg_0592;
    60: op1_07_in03 = reg_0573;
    58: op1_07_in03 = reg_1170;
    78: op1_07_in03 = reg_0735;
    70: op1_07_in03 = reg_1339;
    46: op1_07_in03 = reg_0496;
    51: op1_07_in03 = reg_0298;
    88: op1_07_in03 = reg_0328;
    79: op1_07_in03 = reg_1298;
    59: op1_07_in03 = reg_0323;
    48: op1_07_in03 = reg_0470;
    80: op1_07_in03 = imem06_in[7:4];
    62: op1_07_in03 = reg_0151;
    52: op1_07_in03 = reg_0398;
    81: op1_07_in03 = reg_0275;
    63: op1_07_in03 = reg_0797;
    82: op1_07_in03 = reg_0608;
    89: op1_07_in03 = reg_0180;
    83: op1_07_in03 = reg_0613;
    84: op1_07_in03 = reg_1516;
    65: op1_07_in03 = reg_0229;
    85: op1_07_in03 = reg_1299;
    37: op1_07_in03 = reg_0289;
    90: op1_07_in03 = reg_0145;
    66: op1_07_in03 = reg_0460;
    91: op1_07_in03 = reg_0632;
    47: op1_07_in03 = reg_0223;
    67: op1_07_in03 = reg_0568;
    92: op1_07_in03 = reg_1325;
    93: op1_07_in03 = reg_1505;
    94: op1_07_in03 = reg_0045;
    95: op1_07_in03 = reg_0384;
    44: op1_07_in03 = reg_0181;
    96: op1_07_in03 = reg_0940;
    97: op1_07_in03 = reg_0697;
    98: op1_07_in03 = reg_0468;
    99: op1_07_in03 = reg_0292;
    100: op1_07_in03 = reg_0627;
    101: op1_07_in03 = reg_0557;
    128: op1_07_in03 = reg_0557;
    102: op1_07_in03 = reg_0522;
    103: op1_07_in03 = reg_0186;
    104: op1_07_in03 = reg_0726;
    105: op1_07_in03 = reg_1489;
    106: op1_07_in03 = reg_0719;
    107: op1_07_in03 = reg_0975;
    108: op1_07_in03 = reg_0843;
    109: op1_07_in03 = reg_0615;
    110: op1_07_in03 = reg_1372;
    111: op1_07_in03 = reg_0806;
    112: op1_07_in03 = reg_0789;
    34: op1_07_in03 = reg_0618;
    113: op1_07_in03 = reg_1277;
    114: op1_07_in03 = reg_0869;
    115: op1_07_in03 = reg_0901;
    116: op1_07_in03 = reg_0443;
    38: op1_07_in03 = reg_0593;
    22: op1_07_in03 = reg_0087;
    117: op1_07_in03 = reg_0390;
    118: op1_07_in03 = reg_1447;
    119: op1_07_in03 = reg_0049;
    42: op1_07_in03 = reg_0438;
    120: op1_07_in03 = reg_1028;
    121: op1_07_in03 = reg_1204;
    122: op1_07_in03 = reg_0295;
    123: op1_07_in03 = reg_0249;
    124: op1_07_in03 = reg_0271;
    125: op1_07_in03 = reg_1199;
    126: op1_07_in03 = reg_0393;
    127: op1_07_in03 = imem04_in[15:12];
    129: op1_07_in03 = reg_0059;
    130: op1_07_in03 = reg_1455;
    131: op1_07_in03 = reg_0667;
    default: op1_07_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv03 = 1;
    53: op1_07_inv03 = 1;
    55: op1_07_inv03 = 1;
    50: op1_07_inv03 = 1;
    56: op1_07_inv03 = 1;
    87: op1_07_inv03 = 1;
    60: op1_07_inv03 = 1;
    58: op1_07_inv03 = 1;
    51: op1_07_inv03 = 1;
    79: op1_07_inv03 = 1;
    59: op1_07_inv03 = 1;
    48: op1_07_inv03 = 1;
    81: op1_07_inv03 = 1;
    89: op1_07_inv03 = 1;
    64: op1_07_inv03 = 1;
    37: op1_07_inv03 = 1;
    66: op1_07_inv03 = 1;
    44: op1_07_inv03 = 1;
    96: op1_07_inv03 = 1;
    99: op1_07_inv03 = 1;
    100: op1_07_inv03 = 1;
    103: op1_07_inv03 = 1;
    104: op1_07_inv03 = 1;
    105: op1_07_inv03 = 1;
    112: op1_07_inv03 = 1;
    113: op1_07_inv03 = 1;
    115: op1_07_inv03 = 1;
    117: op1_07_inv03 = 1;
    42: op1_07_inv03 = 1;
    120: op1_07_inv03 = 1;
    126: op1_07_inv03 = 1;
    127: op1_07_inv03 = 1;
    130: op1_07_inv03 = 1;
    131: op1_07_inv03 = 1;
    default: op1_07_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in04 = reg_0843;
    53: op1_07_in04 = reg_0637;
    55: op1_07_in04 = reg_0931;
    86: op1_07_in04 = reg_1098;
    69: op1_07_in04 = reg_0952;
    73: op1_07_in04 = reg_0063;
    49: op1_07_in04 = reg_0029;
    50: op1_07_in04 = reg_0555;
    129: op1_07_in04 = reg_0555;
    54: op1_07_in04 = reg_0402;
    71: op1_07_in04 = reg_1027;
    74: op1_07_in04 = reg_0861;
    68: op1_07_in04 = reg_1093;
    75: op1_07_in04 = reg_0458;
    61: op1_07_in04 = reg_0221;
    56: op1_07_in04 = reg_0804;
    87: op1_07_in04 = reg_0411;
    76: op1_07_in04 = reg_0418;
    57: op1_07_in04 = reg_0362;
    77: op1_07_in04 = reg_1298;
    78: op1_07_in04 = reg_1298;
    33: op1_07_in04 = reg_0004;
    60: op1_07_in04 = reg_0709;
    58: op1_07_in04 = imem07_in[15:12];
    70: op1_07_in04 = reg_0319;
    48: op1_07_in04 = reg_0319;
    46: op1_07_in04 = reg_0474;
    51: op1_07_in04 = reg_0297;
    88: op1_07_in04 = reg_0759;
    79: op1_07_in04 = reg_0832;
    85: op1_07_in04 = reg_0832;
    59: op1_07_in04 = reg_0270;
    80: op1_07_in04 = reg_0116;
    62: op1_07_in04 = imem05_in[3:0];
    52: op1_07_in04 = reg_0859;
    81: op1_07_in04 = reg_0799;
    63: op1_07_in04 = reg_0370;
    82: op1_07_in04 = reg_0055;
    89: op1_07_in04 = reg_0789;
    83: op1_07_in04 = reg_0250;
    64: op1_07_in04 = reg_0314;
    84: op1_07_in04 = reg_1517;
    65: op1_07_in04 = reg_0600;
    101: op1_07_in04 = reg_0600;
    37: op1_07_in04 = reg_0459;
    90: op1_07_in04 = reg_0142;
    66: op1_07_in04 = reg_0959;
    91: op1_07_in04 = reg_0006;
    47: op1_07_in04 = reg_0324;
    67: op1_07_in04 = reg_0979;
    92: op1_07_in04 = imem04_in[3:0];
    116: op1_07_in04 = imem04_in[3:0];
    93: op1_07_in04 = reg_1504;
    94: op1_07_in04 = reg_1402;
    95: op1_07_in04 = reg_0385;
    44: op1_07_in04 = reg_0150;
    96: op1_07_in04 = reg_1070;
    97: op1_07_in04 = reg_0794;
    98: op1_07_in04 = reg_0430;
    99: op1_07_in04 = reg_0077;
    100: op1_07_in04 = reg_0048;
    102: op1_07_in04 = reg_0171;
    122: op1_07_in04 = reg_0171;
    103: op1_07_in04 = reg_1453;
    104: op1_07_in04 = reg_0148;
    105: op1_07_in04 = reg_1487;
    106: op1_07_in04 = reg_0065;
    107: op1_07_in04 = reg_0712;
    108: op1_07_in04 = reg_1281;
    109: op1_07_in04 = reg_0486;
    110: op1_07_in04 = reg_0034;
    111: op1_07_in04 = reg_0613;
    112: op1_07_in04 = reg_0375;
    34: op1_07_in04 = reg_0103;
    113: op1_07_in04 = reg_0806;
    114: op1_07_in04 = reg_0752;
    115: op1_07_in04 = reg_0080;
    38: op1_07_in04 = reg_0053;
    22: op1_07_in04 = reg_0050;
    117: op1_07_in04 = reg_0326;
    118: op1_07_in04 = reg_0962;
    119: op1_07_in04 = reg_0444;
    42: op1_07_in04 = reg_0161;
    120: op1_07_in04 = reg_0485;
    121: op1_07_in04 = reg_0396;
    123: op1_07_in04 = reg_1405;
    124: op1_07_in04 = reg_1326;
    125: op1_07_in04 = reg_0178;
    126: op1_07_in04 = reg_0828;
    127: op1_07_in04 = reg_1200;
    128: op1_07_in04 = reg_1314;
    130: op1_07_in04 = reg_0112;
    131: op1_07_in04 = reg_1350;
    default: op1_07_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_07_inv04 = 1;
    73: op1_07_inv04 = 1;
    50: op1_07_inv04 = 1;
    71: op1_07_inv04 = 1;
    74: op1_07_inv04 = 1;
    61: op1_07_inv04 = 1;
    56: op1_07_inv04 = 1;
    76: op1_07_inv04 = 1;
    58: op1_07_inv04 = 1;
    79: op1_07_inv04 = 1;
    59: op1_07_inv04 = 1;
    48: op1_07_inv04 = 1;
    62: op1_07_inv04 = 1;
    52: op1_07_inv04 = 1;
    81: op1_07_inv04 = 1;
    63: op1_07_inv04 = 1;
    89: op1_07_inv04 = 1;
    83: op1_07_inv04 = 1;
    85: op1_07_inv04 = 1;
    37: op1_07_inv04 = 1;
    66: op1_07_inv04 = 1;
    47: op1_07_inv04 = 1;
    67: op1_07_inv04 = 1;
    93: op1_07_inv04 = 1;
    97: op1_07_inv04 = 1;
    98: op1_07_inv04 = 1;
    100: op1_07_inv04 = 1;
    103: op1_07_inv04 = 1;
    104: op1_07_inv04 = 1;
    105: op1_07_inv04 = 1;
    106: op1_07_inv04 = 1;
    110: op1_07_inv04 = 1;
    112: op1_07_inv04 = 1;
    113: op1_07_inv04 = 1;
    115: op1_07_inv04 = 1;
    116: op1_07_inv04 = 1;
    38: op1_07_inv04 = 1;
    42: op1_07_inv04 = 1;
    121: op1_07_inv04 = 1;
    123: op1_07_inv04 = 1;
    127: op1_07_inv04 = 1;
    129: op1_07_inv04 = 1;
    130: op1_07_inv04 = 1;
    131: op1_07_inv04 = 1;
    default: op1_07_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in05 = reg_1243;
    53: op1_07_in05 = reg_0261;
    55: op1_07_in05 = reg_0783;
    86: op1_07_in05 = reg_0255;
    69: op1_07_in05 = reg_1092;
    73: op1_07_in05 = reg_0675;
    49: op1_07_in05 = reg_0741;
    50: op1_07_in05 = reg_0229;
    54: op1_07_in05 = reg_0383;
    71: op1_07_in05 = reg_1453;
    83: op1_07_in05 = reg_1453;
    74: op1_07_in05 = reg_0828;
    68: op1_07_in05 = reg_0108;
    75: op1_07_in05 = reg_0780;
    61: op1_07_in05 = reg_0476;
    56: op1_07_in05 = reg_0805;
    113: op1_07_in05 = reg_0805;
    87: op1_07_in05 = imem04_in[11:8];
    76: op1_07_in05 = reg_0872;
    57: op1_07_in05 = reg_0093;
    77: op1_07_in05 = reg_0168;
    60: op1_07_in05 = reg_0706;
    119: op1_07_in05 = reg_0706;
    58: op1_07_in05 = reg_0629;
    78: op1_07_in05 = reg_1431;
    126: op1_07_in05 = reg_1431;
    70: op1_07_in05 = reg_0862;
    46: op1_07_in05 = reg_0457;
    51: op1_07_in05 = reg_0923;
    88: op1_07_in05 = reg_0154;
    79: op1_07_in05 = reg_0733;
    59: op1_07_in05 = reg_0269;
    48: op1_07_in05 = reg_0338;
    80: op1_07_in05 = reg_0716;
    62: op1_07_in05 = reg_1035;
    52: op1_07_in05 = reg_0371;
    81: op1_07_in05 = reg_0207;
    63: op1_07_in05 = reg_0904;
    82: op1_07_in05 = reg_0256;
    89: op1_07_in05 = reg_0989;
    64: op1_07_in05 = reg_1314;
    84: op1_07_in05 = reg_0627;
    65: op1_07_in05 = imem07_in[7:4];
    85: op1_07_in05 = reg_0877;
    37: op1_07_in05 = reg_0271;
    90: op1_07_in05 = reg_1518;
    66: op1_07_in05 = imem00_in[3:0];
    91: op1_07_in05 = reg_0840;
    47: op1_07_in05 = reg_0299;
    67: op1_07_in05 = reg_0522;
    92: op1_07_in05 = imem04_in[15:12];
    93: op1_07_in05 = reg_0585;
    94: op1_07_in05 = reg_0183;
    95: op1_07_in05 = reg_0078;
    44: op1_07_in05 = reg_0575;
    96: op1_07_in05 = reg_0090;
    97: op1_07_in05 = reg_0937;
    98: op1_07_in05 = reg_0438;
    99: op1_07_in05 = reg_0896;
    100: op1_07_in05 = reg_0880;
    101: op1_07_in05 = reg_0349;
    102: op1_07_in05 = reg_0419;
    103: op1_07_in05 = reg_1201;
    104: op1_07_in05 = reg_0290;
    105: op1_07_in05 = reg_0806;
    106: op1_07_in05 = reg_0445;
    107: op1_07_in05 = reg_0495;
    108: op1_07_in05 = reg_1277;
    109: op1_07_in05 = reg_0523;
    110: op1_07_in05 = reg_0574;
    111: op1_07_in05 = reg_0555;
    112: op1_07_in05 = reg_0556;
    34: op1_07_in05 = reg_0114;
    114: op1_07_in05 = reg_1501;
    115: op1_07_in05 = reg_0041;
    116: op1_07_in05 = reg_0656;
    38: op1_07_in05 = reg_0087;
    117: op1_07_in05 = reg_1451;
    118: op1_07_in05 = reg_1093;
    42: op1_07_in05 = reg_0162;
    120: op1_07_in05 = reg_0459;
    121: op1_07_in05 = reg_0977;
    122: op1_07_in05 = reg_0119;
    123: op1_07_in05 = reg_1393;
    124: op1_07_in05 = reg_0859;
    125: op1_07_in05 = reg_0107;
    127: op1_07_in05 = reg_0681;
    128: op1_07_in05 = reg_0957;
    129: op1_07_in05 = reg_1052;
    130: op1_07_in05 = reg_0628;
    131: op1_07_in05 = reg_1349;
    default: op1_07_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_07_inv05 = 1;
    69: op1_07_inv05 = 1;
    73: op1_07_inv05 = 1;
    50: op1_07_inv05 = 1;
    71: op1_07_inv05 = 1;
    74: op1_07_inv05 = 1;
    57: op1_07_inv05 = 1;
    60: op1_07_inv05 = 1;
    46: op1_07_inv05 = 1;
    59: op1_07_inv05 = 1;
    48: op1_07_inv05 = 1;
    62: op1_07_inv05 = 1;
    89: op1_07_inv05 = 1;
    83: op1_07_inv05 = 1;
    64: op1_07_inv05 = 1;
    65: op1_07_inv05 = 1;
    85: op1_07_inv05 = 1;
    37: op1_07_inv05 = 1;
    90: op1_07_inv05 = 1;
    66: op1_07_inv05 = 1;
    91: op1_07_inv05 = 1;
    92: op1_07_inv05 = 1;
    93: op1_07_inv05 = 1;
    94: op1_07_inv05 = 1;
    44: op1_07_inv05 = 1;
    97: op1_07_inv05 = 1;
    98: op1_07_inv05 = 1;
    102: op1_07_inv05 = 1;
    105: op1_07_inv05 = 1;
    108: op1_07_inv05 = 1;
    111: op1_07_inv05 = 1;
    112: op1_07_inv05 = 1;
    113: op1_07_inv05 = 1;
    115: op1_07_inv05 = 1;
    116: op1_07_inv05 = 1;
    38: op1_07_inv05 = 1;
    117: op1_07_inv05 = 1;
    119: op1_07_inv05 = 1;
    42: op1_07_inv05 = 1;
    120: op1_07_inv05 = 1;
    122: op1_07_inv05 = 1;
    130: op1_07_inv05 = 1;
    default: op1_07_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in06 = imem00_in[7:4];
    53: op1_07_in06 = reg_0583;
    55: op1_07_in06 = reg_0141;
    86: op1_07_in06 = reg_0632;
    69: op1_07_in06 = reg_0478;
    73: op1_07_in06 = reg_0204;
    49: op1_07_in06 = reg_0740;
    50: op1_07_in06 = imem00_in[3:0];
    54: op1_07_in06 = reg_0362;
    71: op1_07_in06 = reg_1229;
    74: op1_07_in06 = reg_0206;
    68: op1_07_in06 = reg_0505;
    75: op1_07_in06 = reg_1436;
    61: op1_07_in06 = reg_1206;
    56: op1_07_in06 = imem00_in[11:8];
    87: op1_07_in06 = reg_0975;
    76: op1_07_in06 = reg_0318;
    57: op1_07_in06 = reg_0079;
    77: op1_07_in06 = reg_1259;
    60: op1_07_in06 = reg_0710;
    58: op1_07_in06 = reg_1183;
    78: op1_07_in06 = reg_0395;
    70: op1_07_in06 = imem05_in[3:0];
    46: op1_07_in06 = reg_0776;
    107: op1_07_in06 = reg_0776;
    51: op1_07_in06 = reg_0140;
    88: op1_07_in06 = reg_0573;
    79: op1_07_in06 = reg_0168;
    59: op1_07_in06 = reg_0461;
    48: op1_07_in06 = reg_0020;
    80: op1_07_in06 = reg_0194;
    62: op1_07_in06 = reg_0925;
    52: op1_07_in06 = reg_0822;
    81: op1_07_in06 = imem06_in[15:12];
    63: op1_07_in06 = reg_0470;
    82: op1_07_in06 = reg_1260;
    89: op1_07_in06 = reg_0070;
    83: op1_07_in06 = reg_1230;
    64: op1_07_in06 = reg_0329;
    84: op1_07_in06 = reg_0220;
    65: op1_07_in06 = reg_1351;
    85: op1_07_in06 = imem05_in[11:8];
    37: op1_07_in06 = reg_0213;
    90: op1_07_in06 = reg_1517;
    66: op1_07_in06 = reg_0353;
    91: op1_07_in06 = reg_0699;
    47: op1_07_in06 = reg_0157;
    67: op1_07_in06 = reg_0323;
    92: op1_07_in06 = reg_0297;
    93: op1_07_in06 = reg_0529;
    94: op1_07_in06 = reg_0090;
    95: op1_07_in06 = reg_0257;
    44: op1_07_in06 = reg_0736;
    96: op1_07_in06 = reg_0275;
    97: op1_07_in06 = reg_0418;
    98: op1_07_in06 = reg_0290;
    99: op1_07_in06 = reg_1068;
    100: op1_07_in06 = reg_1149;
    128: op1_07_in06 = reg_1149;
    101: op1_07_in06 = reg_0954;
    102: op1_07_in06 = reg_0023;
    103: op1_07_in06 = reg_1205;
    104: op1_07_in06 = reg_0360;
    105: op1_07_in06 = reg_0613;
    106: op1_07_in06 = reg_0579;
    108: op1_07_in06 = reg_1491;
    109: op1_07_in06 = reg_0293;
    110: op1_07_in06 = reg_0488;
    111: op1_07_in06 = reg_1052;
    112: op1_07_in06 = reg_1314;
    34: op1_07_in06 = reg_0228;
    113: op1_07_in06 = reg_0486;
    114: op1_07_in06 = reg_1504;
    115: op1_07_in06 = reg_0011;
    116: op1_07_in06 = reg_1383;
    117: op1_07_in06 = reg_0126;
    118: op1_07_in06 = reg_0252;
    119: op1_07_in06 = reg_1063;
    42: op1_07_in06 = reg_0146;
    120: op1_07_in06 = reg_0927;
    121: op1_07_in06 = reg_0015;
    122: op1_07_in06 = reg_1202;
    123: op1_07_in06 = reg_0202;
    124: op1_07_in06 = reg_0752;
    125: op1_07_in06 = reg_0104;
    126: op1_07_in06 = reg_0039;
    127: op1_07_in06 = reg_1082;
    129: op1_07_in06 = reg_0523;
    130: op1_07_in06 = reg_0379;
    131: op1_07_in06 = reg_0159;
    default: op1_07_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv06 = 1;
    50: op1_07_inv06 = 1;
    68: op1_07_inv06 = 1;
    61: op1_07_inv06 = 1;
    87: op1_07_inv06 = 1;
    76: op1_07_inv06 = 1;
    57: op1_07_inv06 = 1;
    60: op1_07_inv06 = 1;
    78: op1_07_inv06 = 1;
    70: op1_07_inv06 = 1;
    51: op1_07_inv06 = 1;
    59: op1_07_inv06 = 1;
    62: op1_07_inv06 = 1;
    52: op1_07_inv06 = 1;
    81: op1_07_inv06 = 1;
    89: op1_07_inv06 = 1;
    83: op1_07_inv06 = 1;
    84: op1_07_inv06 = 1;
    37: op1_07_inv06 = 1;
    66: op1_07_inv06 = 1;
    91: op1_07_inv06 = 1;
    47: op1_07_inv06 = 1;
    67: op1_07_inv06 = 1;
    92: op1_07_inv06 = 1;
    93: op1_07_inv06 = 1;
    94: op1_07_inv06 = 1;
    44: op1_07_inv06 = 1;
    96: op1_07_inv06 = 1;
    99: op1_07_inv06 = 1;
    101: op1_07_inv06 = 1;
    105: op1_07_inv06 = 1;
    106: op1_07_inv06 = 1;
    107: op1_07_inv06 = 1;
    109: op1_07_inv06 = 1;
    113: op1_07_inv06 = 1;
    117: op1_07_inv06 = 1;
    118: op1_07_inv06 = 1;
    119: op1_07_inv06 = 1;
    121: op1_07_inv06 = 1;
    124: op1_07_inv06 = 1;
    127: op1_07_inv06 = 1;
    128: op1_07_inv06 = 1;
    default: op1_07_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in07 = imem00_in[11:8];
    53: op1_07_in07 = reg_0586;
    55: op1_07_in07 = reg_0397;
    86: op1_07_in07 = reg_0006;
    69: op1_07_in07 = reg_0831;
    73: op1_07_in07 = reg_1269;
    70: op1_07_in07 = reg_1269;
    49: op1_07_in07 = reg_0137;
    50: op1_07_in07 = reg_0820;
    54: op1_07_in07 = reg_0047;
    71: op1_07_in07 = reg_0459;
    61: op1_07_in07 = reg_0459;
    74: op1_07_in07 = reg_0038;
    68: op1_07_in07 = imem03_in[3:0];
    75: op1_07_in07 = reg_1435;
    56: op1_07_in07 = reg_1201;
    83: op1_07_in07 = reg_1201;
    87: op1_07_in07 = reg_0534;
    76: op1_07_in07 = reg_1373;
    96: op1_07_in07 = reg_1373;
    57: op1_07_in07 = reg_0088;
    77: op1_07_in07 = reg_0346;
    60: op1_07_in07 = reg_0444;
    58: op1_07_in07 = reg_0245;
    78: op1_07_in07 = reg_1168;
    46: op1_07_in07 = imem02_in[7:4];
    51: op1_07_in07 = reg_0030;
    88: op1_07_in07 = reg_0049;
    79: op1_07_in07 = reg_0646;
    59: op1_07_in07 = reg_0667;
    48: op1_07_in07 = reg_0794;
    80: op1_07_in07 = reg_0527;
    62: op1_07_in07 = reg_1105;
    52: op1_07_in07 = reg_0718;
    81: op1_07_in07 = reg_1437;
    63: op1_07_in07 = reg_0097;
    82: op1_07_in07 = reg_0474;
    89: op1_07_in07 = reg_1313;
    64: op1_07_in07 = reg_1301;
    112: op1_07_in07 = reg_1301;
    84: op1_07_in07 = reg_0558;
    65: op1_07_in07 = reg_0225;
    85: op1_07_in07 = reg_1164;
    37: op1_07_in07 = reg_0230;
    90: op1_07_in07 = reg_1208;
    66: op1_07_in07 = reg_0189;
    91: op1_07_in07 = reg_0235;
    47: op1_07_in07 = reg_0169;
    67: op1_07_in07 = reg_0296;
    92: op1_07_in07 = reg_1203;
    93: op1_07_in07 = reg_0979;
    94: op1_07_in07 = reg_0492;
    95: op1_07_in07 = reg_0662;
    44: op1_07_in07 = reg_0733;
    97: op1_07_in07 = reg_0302;
    98: op1_07_in07 = reg_0362;
    99: op1_07_in07 = imem02_in[3:0];
    100: op1_07_in07 = reg_0291;
    128: op1_07_in07 = reg_0291;
    101: op1_07_in07 = reg_0957;
    102: op1_07_in07 = imem07_in[15:12];
    103: op1_07_in07 = reg_0155;
    104: op1_07_in07 = reg_0365;
    105: op1_07_in07 = reg_1227;
    106: op1_07_in07 = reg_0735;
    107: op1_07_in07 = reg_1455;
    108: op1_07_in07 = reg_0580;
    109: op1_07_in07 = reg_1027;
    110: op1_07_in07 = reg_1215;
    111: op1_07_in07 = reg_1229;
    34: op1_07_in07 = reg_0084;
    113: op1_07_in07 = reg_0523;
    114: op1_07_in07 = reg_0116;
    115: op1_07_in07 = reg_1068;
    116: op1_07_in07 = reg_1368;
    117: op1_07_in07 = reg_0106;
    118: op1_07_in07 = reg_1216;
    119: op1_07_in07 = reg_0216;
    42: op1_07_in07 = reg_0402;
    120: op1_07_in07 = reg_0435;
    121: op1_07_in07 = reg_0017;
    122: op1_07_in07 = reg_0754;
    123: op1_07_in07 = reg_0353;
    124: op1_07_in07 = reg_1508;
    125: op1_07_in07 = reg_0458;
    126: op1_07_in07 = reg_0784;
    127: op1_07_in07 = reg_1041;
    129: op1_07_in07 = reg_0293;
    130: op1_07_in07 = reg_0007;
    131: op1_07_in07 = reg_0921;
    default: op1_07_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_07_inv07 = 1;
    55: op1_07_inv07 = 1;
    69: op1_07_inv07 = 1;
    73: op1_07_inv07 = 1;
    50: op1_07_inv07 = 1;
    68: op1_07_inv07 = 1;
    87: op1_07_inv07 = 1;
    60: op1_07_inv07 = 1;
    58: op1_07_inv07 = 1;
    78: op1_07_inv07 = 1;
    70: op1_07_inv07 = 1;
    46: op1_07_inv07 = 1;
    79: op1_07_inv07 = 1;
    48: op1_07_inv07 = 1;
    81: op1_07_inv07 = 1;
    82: op1_07_inv07 = 1;
    64: op1_07_inv07 = 1;
    84: op1_07_inv07 = 1;
    90: op1_07_inv07 = 1;
    91: op1_07_inv07 = 1;
    92: op1_07_inv07 = 1;
    93: op1_07_inv07 = 1;
    95: op1_07_inv07 = 1;
    96: op1_07_inv07 = 1;
    97: op1_07_inv07 = 1;
    100: op1_07_inv07 = 1;
    104: op1_07_inv07 = 1;
    107: op1_07_inv07 = 1;
    116: op1_07_inv07 = 1;
    117: op1_07_inv07 = 1;
    118: op1_07_inv07 = 1;
    42: op1_07_inv07 = 1;
    120: op1_07_inv07 = 1;
    123: op1_07_inv07 = 1;
    124: op1_07_inv07 = 1;
    125: op1_07_inv07 = 1;
    127: op1_07_inv07 = 1;
    128: op1_07_inv07 = 1;
    129: op1_07_inv07 = 1;
    default: op1_07_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in08 = imem00_in[15:12];
    53: op1_07_in08 = reg_0584;
    55: op1_07_in08 = reg_0374;
    86: op1_07_in08 = reg_0191;
    69: op1_07_in08 = reg_0734;
    73: op1_07_in08 = reg_0136;
    49: op1_07_in08 = reg_0228;
    50: op1_07_in08 = reg_0293;
    54: op1_07_in08 = reg_0899;
    104: op1_07_in08 = reg_0899;
    71: op1_07_in08 = reg_0201;
    74: op1_07_in08 = reg_0039;
    68: op1_07_in08 = imem03_in[7:4];
    75: op1_07_in08 = reg_0268;
    81: op1_07_in08 = reg_0268;
    61: op1_07_in08 = reg_0959;
    56: op1_07_in08 = reg_1205;
    87: op1_07_in08 = reg_1369;
    76: op1_07_in08 = reg_0601;
    57: op1_07_in08 = reg_0043;
    77: op1_07_in08 = reg_0567;
    60: op1_07_in08 = reg_0177;
    58: op1_07_in08 = reg_0187;
    78: op1_07_in08 = reg_0996;
    70: op1_07_in08 = reg_0333;
    46: op1_07_in08 = reg_0934;
    51: op1_07_in08 = reg_0661;
    88: op1_07_in08 = reg_1448;
    79: op1_07_in08 = reg_0649;
    59: op1_07_in08 = reg_0668;
    48: op1_07_in08 = reg_0799;
    80: op1_07_in08 = reg_0571;
    62: op1_07_in08 = reg_0193;
    52: op1_07_in08 = reg_0670;
    63: op1_07_in08 = reg_0032;
    82: op1_07_in08 = reg_0494;
    89: op1_07_in08 = reg_0627;
    83: op1_07_in08 = reg_1418;
    64: op1_07_in08 = reg_0505;
    84: op1_07_in08 = reg_1208;
    65: op1_07_in08 = reg_1345;
    85: op1_07_in08 = reg_0648;
    37: op1_07_in08 = reg_0169;
    90: op1_07_in08 = reg_0104;
    66: op1_07_in08 = reg_0428;
    91: op1_07_in08 = reg_0185;
    47: op1_07_in08 = reg_0665;
    67: op1_07_in08 = reg_0295;
    92: op1_07_in08 = reg_0574;
    93: op1_07_in08 = reg_1225;
    94: op1_07_in08 = reg_0864;
    95: op1_07_in08 = reg_0989;
    44: op1_07_in08 = reg_0735;
    96: op1_07_in08 = reg_0344;
    97: op1_07_in08 = reg_1486;
    98: op1_07_in08 = reg_0092;
    99: op1_07_in08 = reg_0475;
    100: op1_07_in08 = reg_0673;
    101: op1_07_in08 = reg_0597;
    102: op1_07_in08 = reg_0135;
    103: op1_07_in08 = reg_0821;
    105: op1_07_in08 = reg_1393;
    106: op1_07_in08 = reg_1431;
    107: op1_07_in08 = reg_0106;
    108: op1_07_in08 = reg_0805;
    109: op1_07_in08 = reg_0221;
    110: op1_07_in08 = reg_1041;
    111: op1_07_in08 = reg_1417;
    112: op1_07_in08 = reg_1093;
    113: op1_07_in08 = reg_0485;
    114: op1_07_in08 = reg_1303;
    115: op1_07_in08 = reg_0895;
    116: op1_07_in08 = reg_0337;
    117: op1_07_in08 = reg_0629;
    118: op1_07_in08 = reg_0656;
    119: op1_07_in08 = reg_1001;
    42: op1_07_in08 = reg_0403;
    120: op1_07_in08 = reg_0387;
    121: op1_07_in08 = imem07_in[11:8];
    122: op1_07_in08 = reg_0195;
    123: op1_07_in08 = reg_0188;
    124: op1_07_in08 = reg_1302;
    125: op1_07_in08 = reg_0750;
    126: op1_07_in08 = reg_0826;
    127: op1_07_in08 = reg_0097;
    128: op1_07_in08 = reg_0288;
    129: op1_07_in08 = reg_1027;
    130: op1_07_in08 = reg_0903;
    131: op1_07_in08 = reg_0139;
    default: op1_07_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_07_inv08 = 1;
    55: op1_07_inv08 = 1;
    69: op1_07_inv08 = 1;
    73: op1_07_inv08 = 1;
    50: op1_07_inv08 = 1;
    54: op1_07_inv08 = 1;
    71: op1_07_inv08 = 1;
    75: op1_07_inv08 = 1;
    87: op1_07_inv08 = 1;
    76: op1_07_inv08 = 1;
    77: op1_07_inv08 = 1;
    58: op1_07_inv08 = 1;
    70: op1_07_inv08 = 1;
    46: op1_07_inv08 = 1;
    51: op1_07_inv08 = 1;
    48: op1_07_inv08 = 1;
    80: op1_07_inv08 = 1;
    62: op1_07_inv08 = 1;
    81: op1_07_inv08 = 1;
    82: op1_07_inv08 = 1;
    89: op1_07_inv08 = 1;
    64: op1_07_inv08 = 1;
    65: op1_07_inv08 = 1;
    85: op1_07_inv08 = 1;
    37: op1_07_inv08 = 1;
    90: op1_07_inv08 = 1;
    91: op1_07_inv08 = 1;
    67: op1_07_inv08 = 1;
    92: op1_07_inv08 = 1;
    93: op1_07_inv08 = 1;
    94: op1_07_inv08 = 1;
    95: op1_07_inv08 = 1;
    97: op1_07_inv08 = 1;
    98: op1_07_inv08 = 1;
    103: op1_07_inv08 = 1;
    106: op1_07_inv08 = 1;
    109: op1_07_inv08 = 1;
    110: op1_07_inv08 = 1;
    113: op1_07_inv08 = 1;
    114: op1_07_inv08 = 1;
    118: op1_07_inv08 = 1;
    119: op1_07_inv08 = 1;
    42: op1_07_inv08 = 1;
    121: op1_07_inv08 = 1;
    124: op1_07_inv08 = 1;
    131: op1_07_inv08 = 1;
    default: op1_07_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in09 = reg_0218;
    53: op1_07_in09 = reg_0570;
    55: op1_07_in09 = reg_0825;
    86: op1_07_in09 = reg_0233;
    60: op1_07_in09 = reg_0233;
    69: op1_07_in09 = reg_0573;
    91: op1_07_in09 = reg_0573;
    73: op1_07_in09 = reg_0700;
    49: op1_07_in09 = reg_0004;
    50: op1_07_in09 = reg_0221;
    129: op1_07_in09 = reg_0221;
    54: op1_07_in09 = reg_0902;
    71: op1_07_in09 = reg_0440;
    74: op1_07_in09 = reg_0458;
    68: op1_07_in09 = reg_1282;
    75: op1_07_in09 = reg_0908;
    61: op1_07_in09 = reg_1148;
    56: op1_07_in09 = reg_0459;
    87: op1_07_in09 = reg_1367;
    76: op1_07_in09 = reg_0631;
    57: op1_07_in09 = reg_0041;
    77: op1_07_in09 = reg_0565;
    58: op1_07_in09 = reg_0297;
    78: op1_07_in09 = reg_0174;
    70: op1_07_in09 = reg_0564;
    46: op1_07_in09 = reg_0935;
    51: op1_07_in09 = reg_0285;
    88: op1_07_in09 = reg_0143;
    79: op1_07_in09 = reg_0333;
    59: op1_07_in09 = reg_0324;
    48: op1_07_in09 = reg_0579;
    80: op1_07_in09 = reg_0569;
    124: op1_07_in09 = reg_0569;
    62: op1_07_in09 = reg_0696;
    52: op1_07_in09 = reg_0264;
    81: op1_07_in09 = reg_1508;
    63: op1_07_in09 = reg_1164;
    82: op1_07_in09 = reg_0429;
    89: op1_07_in09 = reg_0952;
    83: op1_07_in09 = reg_0928;
    64: op1_07_in09 = reg_0507;
    84: op1_07_in09 = reg_0113;
    65: op1_07_in09 = reg_0489;
    85: op1_07_in09 = reg_0391;
    37: op1_07_in09 = reg_0185;
    90: op1_07_in09 = reg_1280;
    66: op1_07_in09 = reg_0416;
    47: op1_07_in09 = reg_0661;
    67: op1_07_in09 = reg_0244;
    92: op1_07_in09 = reg_1215;
    93: op1_07_in09 = reg_0323;
    94: op1_07_in09 = reg_0396;
    95: op1_07_in09 = reg_0975;
    44: op1_07_in09 = reg_0346;
    96: op1_07_in09 = reg_0589;
    97: op1_07_in09 = reg_0275;
    98: op1_07_in09 = reg_0901;
    99: op1_07_in09 = reg_0626;
    100: op1_07_in09 = reg_0427;
    101: op1_07_in09 = reg_1300;
    102: op1_07_in09 = reg_0310;
    103: op1_07_in09 = reg_0927;
    104: op1_07_in09 = reg_0595;
    105: op1_07_in09 = reg_0886;
    106: op1_07_in09 = reg_0702;
    107: op1_07_in09 = reg_0802;
    108: op1_07_in09 = reg_1028;
    109: op1_07_in09 = reg_1230;
    110: op1_07_in09 = reg_0199;
    111: op1_07_in09 = reg_1405;
    112: op1_07_in09 = reg_1208;
    113: op1_07_in09 = reg_0987;
    114: op1_07_in09 = reg_0194;
    115: op1_07_in09 = reg_0475;
    116: op1_07_in09 = reg_0694;
    117: op1_07_in09 = reg_1140;
    118: op1_07_in09 = imem04_in[11:8];
    119: op1_07_in09 = reg_1494;
    42: op1_07_in09 = reg_0384;
    120: op1_07_in09 = reg_1254;
    121: op1_07_in09 = reg_0498;
    122: op1_07_in09 = reg_0152;
    123: op1_07_in09 = reg_0410;
    125: op1_07_in09 = reg_0288;
    126: op1_07_in09 = reg_0730;
    127: op1_07_in09 = reg_1151;
    128: op1_07_in09 = reg_0790;
    130: op1_07_in09 = reg_0563;
    131: op1_07_in09 = reg_0779;
    default: op1_07_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_07_inv09 = 1;
    49: op1_07_inv09 = 1;
    50: op1_07_inv09 = 1;
    54: op1_07_inv09 = 1;
    75: op1_07_inv09 = 1;
    87: op1_07_inv09 = 1;
    57: op1_07_inv09 = 1;
    77: op1_07_inv09 = 1;
    60: op1_07_inv09 = 1;
    58: op1_07_inv09 = 1;
    78: op1_07_inv09 = 1;
    70: op1_07_inv09 = 1;
    88: op1_07_inv09 = 1;
    59: op1_07_inv09 = 1;
    80: op1_07_inv09 = 1;
    52: op1_07_inv09 = 1;
    81: op1_07_inv09 = 1;
    64: op1_07_inv09 = 1;
    37: op1_07_inv09 = 1;
    47: op1_07_inv09 = 1;
    93: op1_07_inv09 = 1;
    96: op1_07_inv09 = 1;
    97: op1_07_inv09 = 1;
    98: op1_07_inv09 = 1;
    101: op1_07_inv09 = 1;
    105: op1_07_inv09 = 1;
    106: op1_07_inv09 = 1;
    110: op1_07_inv09 = 1;
    111: op1_07_inv09 = 1;
    112: op1_07_inv09 = 1;
    114: op1_07_inv09 = 1;
    116: op1_07_inv09 = 1;
    118: op1_07_inv09 = 1;
    119: op1_07_inv09 = 1;
    42: op1_07_inv09 = 1;
    120: op1_07_inv09 = 1;
    121: op1_07_inv09 = 1;
    131: op1_07_inv09 = 1;
    default: op1_07_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in10 = reg_1052;
    53: op1_07_in10 = reg_0529;
    55: op1_07_in10 = reg_0827;
    86: op1_07_in10 = reg_0330;
    69: op1_07_in10 = reg_0790;
    73: op1_07_in10 = reg_0173;
    63: op1_07_in10 = reg_0173;
    49: op1_07_in10 = reg_0124;
    50: op1_07_in10 = reg_0172;
    54: op1_07_in10 = reg_0077;
    71: op1_07_in10 = reg_0410;
    74: op1_07_in10 = reg_0399;
    115: op1_07_in10 = reg_0399;
    68: op1_07_in10 = reg_1280;
    75: op1_07_in10 = reg_0984;
    61: op1_07_in10 = reg_0883;
    83: op1_07_in10 = reg_0883;
    103: op1_07_in10 = reg_0883;
    56: op1_07_in10 = reg_0959;
    87: op1_07_in10 = reg_0264;
    76: op1_07_in10 = reg_0589;
    97: op1_07_in10 = reg_0589;
    57: op1_07_in10 = reg_0446;
    77: op1_07_in10 = reg_1181;
    60: op1_07_in10 = reg_0261;
    58: op1_07_in10 = reg_0674;
    78: op1_07_in10 = reg_0648;
    70: op1_07_in10 = reg_0745;
    46: op1_07_in10 = reg_0382;
    51: op1_07_in10 = reg_0366;
    88: op1_07_in10 = reg_0891;
    79: op1_07_in10 = reg_0182;
    59: op1_07_in10 = reg_0310;
    48: op1_07_in10 = reg_0736;
    80: op1_07_in10 = reg_0419;
    62: op1_07_in10 = reg_0870;
    52: op1_07_in10 = reg_0585;
    81: op1_07_in10 = reg_0869;
    82: op1_07_in10 = reg_0326;
    89: op1_07_in10 = reg_0246;
    64: op1_07_in10 = reg_0478;
    84: op1_07_in10 = reg_0505;
    65: op1_07_in10 = reg_0777;
    85: op1_07_in10 = reg_0939;
    37: op1_07_in10 = reg_0187;
    90: op1_07_in10 = reg_0427;
    66: op1_07_in10 = reg_0387;
    91: op1_07_in10 = reg_0179;
    47: op1_07_in10 = reg_0663;
    67: op1_07_in10 = reg_0165;
    92: op1_07_in10 = reg_1214;
    93: op1_07_in10 = reg_0270;
    94: op1_07_in10 = reg_1030;
    95: op1_07_in10 = reg_0530;
    44: op1_07_in10 = reg_0700;
    96: op1_07_in10 = reg_0864;
    98: op1_07_in10 = reg_0464;
    99: op1_07_in10 = reg_0138;
    100: op1_07_in10 = imem04_in[7:4];
    101: op1_07_in10 = reg_0329;
    102: op1_07_in10 = reg_1440;
    104: op1_07_in10 = reg_0727;
    105: op1_07_in10 = reg_0189;
    106: op1_07_in10 = reg_0347;
    107: op1_07_in10 = reg_1098;
    108: op1_07_in10 = reg_0485;
    109: op1_07_in10 = reg_0987;
    110: op1_07_in10 = reg_0033;
    111: op1_07_in10 = reg_1393;
    112: op1_07_in10 = reg_0884;
    113: op1_07_in10 = reg_0460;
    114: op1_07_in10 = reg_0374;
    116: op1_07_in10 = reg_0297;
    117: op1_07_in10 = reg_0631;
    118: op1_07_in10 = reg_0493;
    119: op1_07_in10 = reg_1495;
    42: op1_07_in10 = reg_0386;
    120: op1_07_in10 = reg_0982;
    121: op1_07_in10 = reg_0668;
    122: op1_07_in10 = reg_0215;
    123: op1_07_in10 = reg_0060;
    124: op1_07_in10 = reg_0979;
    125: op1_07_in10 = reg_0531;
    126: op1_07_in10 = reg_0974;
    127: op1_07_in10 = reg_1503;
    128: op1_07_in10 = reg_0411;
    129: op1_07_in10 = reg_1227;
    130: op1_07_in10 = reg_1515;
    131: op1_07_in10 = reg_0031;
    default: op1_07_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_07_inv10 = 1;
    73: op1_07_inv10 = 1;
    49: op1_07_inv10 = 1;
    50: op1_07_inv10 = 1;
    54: op1_07_inv10 = 1;
    68: op1_07_inv10 = 1;
    75: op1_07_inv10 = 1;
    87: op1_07_inv10 = 1;
    76: op1_07_inv10 = 1;
    77: op1_07_inv10 = 1;
    58: op1_07_inv10 = 1;
    78: op1_07_inv10 = 1;
    46: op1_07_inv10 = 1;
    88: op1_07_inv10 = 1;
    59: op1_07_inv10 = 1;
    62: op1_07_inv10 = 1;
    82: op1_07_inv10 = 1;
    89: op1_07_inv10 = 1;
    83: op1_07_inv10 = 1;
    64: op1_07_inv10 = 1;
    65: op1_07_inv10 = 1;
    85: op1_07_inv10 = 1;
    37: op1_07_inv10 = 1;
    91: op1_07_inv10 = 1;
    47: op1_07_inv10 = 1;
    44: op1_07_inv10 = 1;
    97: op1_07_inv10 = 1;
    98: op1_07_inv10 = 1;
    102: op1_07_inv10 = 1;
    105: op1_07_inv10 = 1;
    106: op1_07_inv10 = 1;
    107: op1_07_inv10 = 1;
    109: op1_07_inv10 = 1;
    114: op1_07_inv10 = 1;
    116: op1_07_inv10 = 1;
    118: op1_07_inv10 = 1;
    119: op1_07_inv10 = 1;
    42: op1_07_inv10 = 1;
    120: op1_07_inv10 = 1;
    123: op1_07_inv10 = 1;
    124: op1_07_inv10 = 1;
    125: op1_07_inv10 = 1;
    127: op1_07_inv10 = 1;
    129: op1_07_inv10 = 1;
    130: op1_07_inv10 = 1;
    default: op1_07_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in11 = reg_1454;
    53: op1_07_in11 = reg_0527;
    55: op1_07_in11 = reg_0115;
    86: op1_07_in11 = reg_1063;
    69: op1_07_in11 = reg_0425;
    68: op1_07_in11 = reg_0425;
    73: op1_07_in11 = reg_0646;
    50: op1_07_in11 = reg_0136;
    54: op1_07_in11 = reg_0290;
    71: op1_07_in11 = reg_0203;
    74: op1_07_in11 = reg_0730;
    75: op1_07_in11 = reg_0161;
    61: op1_07_in11 = reg_0188;
    56: op1_07_in11 = reg_0958;
    87: op1_07_in11 = reg_1203;
    76: op1_07_in11 = reg_0151;
    57: op1_07_in11 = reg_0662;
    77: op1_07_in11 = reg_0794;
    85: op1_07_in11 = reg_0794;
    60: op1_07_in11 = reg_1092;
    58: op1_07_in11 = reg_0186;
    78: op1_07_in11 = reg_0650;
    127: op1_07_in11 = reg_0650;
    70: op1_07_in11 = reg_0045;
    46: op1_07_in11 = reg_0379;
    51: op1_07_in11 = reg_0408;
    88: op1_07_in11 = reg_0989;
    79: op1_07_in11 = reg_0986;
    59: op1_07_in11 = reg_0674;
    48: op1_07_in11 = reg_0176;
    80: op1_07_in11 = reg_0583;
    62: op1_07_in11 = imem06_in[7:4];
    52: op1_07_in11 = reg_0584;
    81: op1_07_in11 = reg_0635;
    63: op1_07_in11 = reg_0392;
    82: op1_07_in11 = reg_0105;
    89: op1_07_in11 = reg_1149;
    83: op1_07_in11 = reg_0189;
    64: op1_07_in11 = reg_0328;
    84: op1_07_in11 = reg_0504;
    65: op1_07_in11 = reg_0779;
    37: op1_07_in11 = reg_0170;
    90: op1_07_in11 = reg_0467;
    100: op1_07_in11 = reg_0467;
    66: op1_07_in11 = reg_0075;
    91: op1_07_in11 = reg_0709;
    47: op1_07_in11 = reg_0413;
    67: op1_07_in11 = reg_0269;
    92: op1_07_in11 = reg_0421;
    93: op1_07_in11 = reg_0067;
    94: op1_07_in11 = reg_0193;
    95: op1_07_in11 = reg_0607;
    44: op1_07_in11 = reg_0701;
    96: op1_07_in11 = reg_0449;
    97: op1_07_in11 = reg_0861;
    98: op1_07_in11 = reg_0257;
    99: op1_07_in11 = reg_1260;
    101: op1_07_in11 = reg_0885;
    102: op1_07_in11 = reg_0921;
    103: op1_07_in11 = reg_0722;
    104: op1_07_in11 = reg_0292;
    105: op1_07_in11 = reg_0431;
    106: op1_07_in11 = reg_0184;
    107: op1_07_in11 = reg_0801;
    108: op1_07_in11 = reg_1230;
    109: op1_07_in11 = reg_1201;
    110: op1_07_in11 = reg_0368;
    111: op1_07_in11 = reg_0353;
    112: op1_07_in11 = reg_0350;
    113: op1_07_in11 = reg_0459;
    114: op1_07_in11 = reg_0571;
    115: op1_07_in11 = reg_0845;
    116: op1_07_in11 = reg_0598;
    117: op1_07_in11 = reg_0306;
    118: op1_07_in11 = reg_0297;
    119: op1_07_in11 = reg_1226;
    42: op1_07_in11 = reg_0183;
    120: op1_07_in11 = reg_0163;
    121: op1_07_in11 = reg_0394;
    122: op1_07_in11 = reg_0214;
    123: op1_07_in11 = reg_0072;
    124: op1_07_in11 = reg_1228;
    125: op1_07_in11 = reg_0406;
    126: op1_07_in11 = reg_0860;
    128: op1_07_in11 = reg_1384;
    129: op1_07_in11 = reg_1229;
    130: op1_07_in11 = reg_0330;
    131: op1_07_in11 = reg_0663;
    default: op1_07_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_07_inv11 = 1;
    50: op1_07_inv11 = 1;
    71: op1_07_inv11 = 1;
    61: op1_07_inv11 = 1;
    87: op1_07_inv11 = 1;
    57: op1_07_inv11 = 1;
    60: op1_07_inv11 = 1;
    58: op1_07_inv11 = 1;
    78: op1_07_inv11 = 1;
    46: op1_07_inv11 = 1;
    51: op1_07_inv11 = 1;
    59: op1_07_inv11 = 1;
    48: op1_07_inv11 = 1;
    80: op1_07_inv11 = 1;
    62: op1_07_inv11 = 1;
    81: op1_07_inv11 = 1;
    63: op1_07_inv11 = 1;
    82: op1_07_inv11 = 1;
    89: op1_07_inv11 = 1;
    85: op1_07_inv11 = 1;
    37: op1_07_inv11 = 1;
    66: op1_07_inv11 = 1;
    67: op1_07_inv11 = 1;
    92: op1_07_inv11 = 1;
    95: op1_07_inv11 = 1;
    44: op1_07_inv11 = 1;
    98: op1_07_inv11 = 1;
    99: op1_07_inv11 = 1;
    104: op1_07_inv11 = 1;
    106: op1_07_inv11 = 1;
    115: op1_07_inv11 = 1;
    117: op1_07_inv11 = 1;
    118: op1_07_inv11 = 1;
    119: op1_07_inv11 = 1;
    120: op1_07_inv11 = 1;
    121: op1_07_inv11 = 1;
    122: op1_07_inv11 = 1;
    124: op1_07_inv11 = 1;
    125: op1_07_inv11 = 1;
    126: op1_07_inv11 = 1;
    default: op1_07_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in12 = reg_1230;
    53: op1_07_in12 = reg_0522;
    55: op1_07_in12 = reg_0634;
    86: op1_07_in12 = reg_0177;
    69: op1_07_in12 = reg_0426;
    73: op1_07_in12 = reg_1212;
    50: op1_07_in12 = reg_0492;
    54: op1_07_in12 = reg_0088;
    71: op1_07_in12 = reg_1324;
    123: op1_07_in12 = reg_1324;
    74: op1_07_in12 = reg_0870;
    68: op1_07_in12 = reg_0488;
    75: op1_07_in12 = reg_0716;
    81: op1_07_in12 = reg_0716;
    61: op1_07_in12 = reg_0428;
    56: op1_07_in12 = reg_0524;
    87: op1_07_in12 = reg_1215;
    76: op1_07_in12 = reg_0206;
    57: op1_07_in12 = reg_0742;
    77: op1_07_in12 = reg_0183;
    60: op1_07_in12 = reg_0458;
    58: op1_07_in12 = reg_0169;
    78: op1_07_in12 = reg_0333;
    70: op1_07_in12 = reg_0697;
    44: op1_07_in12 = reg_0697;
    46: op1_07_in12 = reg_0138;
    115: op1_07_in12 = reg_0138;
    51: op1_07_in12 = reg_0413;
    88: op1_07_in12 = reg_0964;
    79: op1_07_in12 = reg_0303;
    59: op1_07_in12 = reg_0156;
    48: op1_07_in12 = reg_0650;
    80: op1_07_in12 = reg_0270;
    62: op1_07_in12 = imem06_in[15:12];
    52: op1_07_in12 = reg_0570;
    114: op1_07_in12 = reg_0570;
    63: op1_07_in12 = reg_0646;
    82: op1_07_in12 = reg_1433;
    89: op1_07_in12 = reg_0481;
    84: op1_07_in12 = reg_0481;
    83: op1_07_in12 = reg_0072;
    64: op1_07_in12 = reg_0330;
    65: op1_07_in12 = reg_0366;
    85: op1_07_in12 = reg_0300;
    37: op1_07_in12 = reg_0310;
    90: op1_07_in12 = reg_0268;
    66: op1_07_in12 = reg_0060;
    91: op1_07_in12 = reg_1425;
    47: op1_07_in12 = reg_0621;
    67: op1_07_in12 = reg_0046;
    92: op1_07_in12 = reg_0412;
    93: op1_07_in12 = reg_0212;
    94: op1_07_in12 = reg_0977;
    95: op1_07_in12 = reg_1235;
    96: op1_07_in12 = reg_0040;
    97: op1_07_in12 = reg_0040;
    98: op1_07_in12 = reg_0402;
    99: op1_07_in12 = reg_0326;
    100: op1_07_in12 = reg_0032;
    101: op1_07_in12 = reg_0443;
    102: op1_07_in12 = reg_0739;
    103: op1_07_in12 = reg_0435;
    104: op1_07_in12 = reg_0335;
    105: op1_07_in12 = reg_0059;
    106: op1_07_in12 = reg_0392;
    107: op1_07_in12 = reg_0069;
    108: op1_07_in12 = reg_0987;
    109: op1_07_in12 = reg_0155;
    110: op1_07_in12 = reg_0065;
    111: op1_07_in12 = reg_0189;
    112: op1_07_in12 = reg_1282;
    113: op1_07_in12 = reg_1406;
    116: op1_07_in12 = reg_1040;
    117: op1_07_in12 = reg_0379;
    118: op1_07_in12 = reg_0281;
    119: op1_07_in12 = reg_1208;
    42: op1_07_in12 = reg_0320;
    120: op1_07_in12 = reg_0241;
    121: op1_07_in12 = reg_1057;
    122: op1_07_in12 = reg_0213;
    124: op1_07_in12 = reg_0296;
    125: op1_07_in12 = reg_0407;
    126: op1_07_in12 = reg_1323;
    127: op1_07_in12 = reg_0579;
    128: op1_07_in12 = reg_0936;
    129: op1_07_in12 = reg_1418;
    130: op1_07_in12 = reg_0444;
    131: op1_07_in12 = reg_0664;
    default: op1_07_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_07_inv12 = 1;
    73: op1_07_inv12 = 1;
    50: op1_07_inv12 = 1;
    54: op1_07_inv12 = 1;
    71: op1_07_inv12 = 1;
    61: op1_07_inv12 = 1;
    87: op1_07_inv12 = 1;
    76: op1_07_inv12 = 1;
    77: op1_07_inv12 = 1;
    60: op1_07_inv12 = 1;
    78: op1_07_inv12 = 1;
    46: op1_07_inv12 = 1;
    79: op1_07_inv12 = 1;
    59: op1_07_inv12 = 1;
    48: op1_07_inv12 = 1;
    62: op1_07_inv12 = 1;
    63: op1_07_inv12 = 1;
    82: op1_07_inv12 = 1;
    89: op1_07_inv12 = 1;
    85: op1_07_inv12 = 1;
    90: op1_07_inv12 = 1;
    91: op1_07_inv12 = 1;
    47: op1_07_inv12 = 1;
    67: op1_07_inv12 = 1;
    94: op1_07_inv12 = 1;
    95: op1_07_inv12 = 1;
    96: op1_07_inv12 = 1;
    98: op1_07_inv12 = 1;
    99: op1_07_inv12 = 1;
    100: op1_07_inv12 = 1;
    103: op1_07_inv12 = 1;
    106: op1_07_inv12 = 1;
    109: op1_07_inv12 = 1;
    112: op1_07_inv12 = 1;
    116: op1_07_inv12 = 1;
    118: op1_07_inv12 = 1;
    120: op1_07_inv12 = 1;
    121: op1_07_inv12 = 1;
    124: op1_07_inv12 = 1;
    125: op1_07_inv12 = 1;
    128: op1_07_inv12 = 1;
    130: op1_07_inv12 = 1;
    default: op1_07_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in13 = reg_0881;
    53: op1_07_in13 = reg_0419;
    55: op1_07_in13 = reg_0636;
    86: op1_07_in13 = reg_0823;
    69: op1_07_in13 = reg_0534;
    64: op1_07_in13 = reg_0534;
    73: op1_07_in13 = reg_0745;
    50: op1_07_in13 = reg_0928;
    54: op1_07_in13 = reg_0291;
    71: op1_07_in13 = reg_0089;
    74: op1_07_in13 = reg_0536;
    68: op1_07_in13 = reg_1367;
    128: op1_07_in13 = reg_1367;
    75: op1_07_in13 = reg_0714;
    81: op1_07_in13 = reg_0714;
    61: op1_07_in13 = reg_0058;
    56: op1_07_in13 = reg_1148;
    87: op1_07_in13 = reg_1082;
    76: op1_07_in13 = reg_0261;
    57: op1_07_in13 = reg_0632;
    77: op1_07_in13 = reg_0477;
    60: op1_07_in13 = reg_1144;
    58: op1_07_in13 = reg_0777;
    78: op1_07_in13 = reg_0565;
    70: op1_07_in13 = reg_0939;
    46: op1_07_in13 = reg_0055;
    51: op1_07_in13 = reg_0100;
    88: op1_07_in13 = reg_0349;
    79: op1_07_in13 = reg_0301;
    59: op1_07_in13 = imem07_in[15:12];
    48: op1_07_in13 = reg_0992;
    80: op1_07_in13 = reg_0152;
    62: op1_07_in13 = reg_0264;
    52: op1_07_in13 = reg_0526;
    63: op1_07_in13 = reg_0066;
    82: op1_07_in13 = reg_0217;
    89: op1_07_in13 = reg_0673;
    83: op1_07_in13 = reg_0057;
    84: op1_07_in13 = reg_0525;
    65: op1_07_in13 = reg_0413;
    85: op1_07_in13 = reg_0872;
    37: op1_07_in13 = reg_0299;
    90: op1_07_in13 = reg_1312;
    66: op1_07_in13 = reg_0059;
    91: op1_07_in13 = reg_0198;
    47: op1_07_in13 = reg_0620;
    67: op1_07_in13 = reg_0537;
    92: op1_07_in13 = reg_0451;
    93: op1_07_in13 = imem07_in[7:4];
    94: op1_07_in13 = reg_0906;
    95: op1_07_in13 = reg_0845;
    44: op1_07_in13 = reg_0175;
    96: op1_07_in13 = reg_0014;
    97: op1_07_in13 = reg_0014;
    98: op1_07_in13 = reg_0728;
    104: op1_07_in13 = reg_0728;
    99: op1_07_in13 = reg_1458;
    100: op1_07_in13 = reg_1369;
    101: op1_07_in13 = reg_0319;
    102: op1_07_in13 = reg_0741;
    103: op1_07_in13 = reg_0071;
    105: op1_07_in13 = reg_0122;
    106: op1_07_in13 = reg_0391;
    107: op1_07_in13 = reg_0006;
    108: op1_07_in13 = reg_0524;
    109: op1_07_in13 = reg_0459;
    110: op1_07_in13 = reg_0346;
    111: op1_07_in13 = reg_0409;
    112: op1_07_in13 = reg_0790;
    113: op1_07_in13 = reg_0927;
    114: op1_07_in13 = reg_0119;
    115: op1_07_in13 = reg_0744;
    116: op1_07_in13 = reg_1143;
    117: op1_07_in13 = reg_0800;
    118: op1_07_in13 = reg_0796;
    119: op1_07_in13 = reg_0707;
    42: op1_07_in13 = reg_0092;
    120: op1_07_in13 = reg_0742;
    121: op1_07_in13 = reg_1055;
    122: op1_07_in13 = reg_0017;
    123: op1_07_in13 = reg_0026;
    124: op1_07_in13 = reg_0977;
    125: op1_07_in13 = reg_0471;
    126: op1_07_in13 = reg_1504;
    127: op1_07_in13 = reg_0332;
    129: op1_07_in13 = reg_0352;
    130: op1_07_in13 = reg_1425;
    131: op1_07_in13 = reg_0740;
    default: op1_07_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_07_inv13 = 1;
    73: op1_07_inv13 = 1;
    50: op1_07_inv13 = 1;
    54: op1_07_inv13 = 1;
    71: op1_07_inv13 = 1;
    74: op1_07_inv13 = 1;
    75: op1_07_inv13 = 1;
    56: op1_07_inv13 = 1;
    87: op1_07_inv13 = 1;
    76: op1_07_inv13 = 1;
    57: op1_07_inv13 = 1;
    77: op1_07_inv13 = 1;
    58: op1_07_inv13 = 1;
    46: op1_07_inv13 = 1;
    51: op1_07_inv13 = 1;
    79: op1_07_inv13 = 1;
    59: op1_07_inv13 = 1;
    48: op1_07_inv13 = 1;
    80: op1_07_inv13 = 1;
    81: op1_07_inv13 = 1;
    83: op1_07_inv13 = 1;
    37: op1_07_inv13 = 1;
    66: op1_07_inv13 = 1;
    47: op1_07_inv13 = 1;
    92: op1_07_inv13 = 1;
    93: op1_07_inv13 = 1;
    95: op1_07_inv13 = 1;
    44: op1_07_inv13 = 1;
    97: op1_07_inv13 = 1;
    101: op1_07_inv13 = 1;
    103: op1_07_inv13 = 1;
    105: op1_07_inv13 = 1;
    110: op1_07_inv13 = 1;
    118: op1_07_inv13 = 1;
    119: op1_07_inv13 = 1;
    120: op1_07_inv13 = 1;
    121: op1_07_inv13 = 1;
    129: op1_07_inv13 = 1;
    130: op1_07_inv13 = 1;
    default: op1_07_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in14 = reg_0267;
    53: op1_07_in14 = reg_0067;
    55: op1_07_in14 = reg_0261;
    86: op1_07_in14 = reg_0707;
    69: op1_07_in14 = reg_0032;
    101: op1_07_in14 = reg_0032;
    73: op1_07_in14 = reg_1181;
    50: op1_07_in14 = reg_0926;
    54: op1_07_in14 = reg_0012;
    71: op1_07_in14 = reg_0372;
    74: op1_07_in14 = reg_0669;
    68: op1_07_in14 = reg_1339;
    75: op1_07_in14 = reg_1302;
    81: op1_07_in14 = reg_1302;
    61: op1_07_in14 = reg_0027;
    56: op1_07_in14 = reg_0928;
    87: op1_07_in14 = reg_0969;
    118: op1_07_in14 = reg_0969;
    76: op1_07_in14 = reg_0399;
    57: op1_07_in14 = reg_0561;
    77: op1_07_in14 = reg_1514;
    60: op1_07_in14 = reg_1147;
    58: op1_07_in14 = reg_0029;
    78: op1_07_in14 = reg_0564;
    70: op1_07_in14 = reg_0302;
    46: op1_07_in14 = reg_0307;
    51: op1_07_in14 = reg_0052;
    88: op1_07_in14 = reg_1314;
    79: op1_07_in14 = reg_0873;
    59: op1_07_in14 = reg_0774;
    48: op1_07_in14 = reg_0045;
    80: op1_07_in14 = reg_0672;
    62: op1_07_in14 = reg_0109;
    52: op1_07_in14 = reg_0528;
    63: op1_07_in14 = reg_0272;
    82: op1_07_in14 = imem02_in[3:0];
    89: op1_07_in14 = reg_0288;
    83: op1_07_in14 = reg_1322;
    64: op1_07_in14 = reg_0531;
    84: op1_07_in14 = reg_0694;
    65: op1_07_in14 = reg_0103;
    85: op1_07_in14 = reg_0274;
    37: op1_07_in14 = reg_0297;
    90: op1_07_in14 = reg_0975;
    66: op1_07_in14 = reg_0786;
    91: op1_07_in14 = reg_1001;
    47: op1_07_in14 = reg_0084;
    67: op1_07_in14 = reg_0496;
    92: op1_07_in14 = reg_0061;
    93: op1_07_in14 = reg_1439;
    94: op1_07_in14 = reg_0397;
    95: op1_07_in14 = reg_0056;
    44: op1_07_in14 = reg_0523;
    96: op1_07_in14 = imem06_in[11:8];
    97: op1_07_in14 = reg_1468;
    98: op1_07_in14 = reg_0042;
    99: op1_07_in14 = reg_1450;
    100: op1_07_in14 = reg_1368;
    102: op1_07_in14 = reg_0620;
    103: op1_07_in14 = reg_0203;
    104: op1_07_in14 = reg_0011;
    105: op1_07_in14 = reg_0277;
    106: op1_07_in14 = reg_1104;
    107: op1_07_in14 = reg_1515;
    108: op1_07_in14 = reg_1406;
    109: op1_07_in14 = reg_0476;
    110: op1_07_in14 = reg_0173;
    111: op1_07_in14 = reg_0410;
    112: op1_07_in14 = reg_1338;
    113: op1_07_in14 = reg_0722;
    129: op1_07_in14 = reg_0722;
    114: op1_07_in14 = reg_0023;
    115: op1_07_in14 = reg_0054;
    116: op1_07_in14 = reg_0268;
    117: op1_07_in14 = reg_0903;
    119: op1_07_in14 = reg_0291;
    42: op1_07_in14 = imem01_in[15:12];
    120: op1_07_in14 = reg_0715;
    121: op1_07_in14 = reg_1315;
    122: op1_07_in14 = reg_0050;
    123: op1_07_in14 = reg_1100;
    124: op1_07_in14 = reg_0046;
    125: op1_07_in14 = reg_0537;
    126: op1_07_in14 = reg_1179;
    127: op1_07_in14 = reg_0604;
    128: op1_07_in14 = reg_0535;
    130: op1_07_in14 = reg_0847;
    131: op1_07_in14 = reg_0415;
    default: op1_07_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_07_inv14 = 1;
    50: op1_07_inv14 = 1;
    74: op1_07_inv14 = 1;
    68: op1_07_inv14 = 1;
    75: op1_07_inv14 = 1;
    61: op1_07_inv14 = 1;
    56: op1_07_inv14 = 1;
    76: op1_07_inv14 = 1;
    57: op1_07_inv14 = 1;
    60: op1_07_inv14 = 1;
    70: op1_07_inv14 = 1;
    59: op1_07_inv14 = 1;
    52: op1_07_inv14 = 1;
    82: op1_07_inv14 = 1;
    83: op1_07_inv14 = 1;
    84: op1_07_inv14 = 1;
    65: op1_07_inv14 = 1;
    37: op1_07_inv14 = 1;
    91: op1_07_inv14 = 1;
    93: op1_07_inv14 = 1;
    94: op1_07_inv14 = 1;
    96: op1_07_inv14 = 1;
    97: op1_07_inv14 = 1;
    98: op1_07_inv14 = 1;
    100: op1_07_inv14 = 1;
    107: op1_07_inv14 = 1;
    112: op1_07_inv14 = 1;
    115: op1_07_inv14 = 1;
    117: op1_07_inv14 = 1;
    42: op1_07_inv14 = 1;
    121: op1_07_inv14 = 1;
    125: op1_07_inv14 = 1;
    128: op1_07_inv14 = 1;
    131: op1_07_inv14 = 1;
    default: op1_07_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in15 = reg_0917;
    53: op1_07_in15 = reg_0023;
    55: op1_07_in15 = reg_0264;
    86: op1_07_in15 = reg_0891;
    69: op1_07_in15 = reg_0252;
    73: op1_07_in15 = reg_0183;
    50: op1_07_in15 = reg_0389;
    54: op1_07_in15 = reg_0662;
    71: op1_07_in15 = reg_0258;
    74: op1_07_in15 = reg_0115;
    68: op1_07_in15 = reg_1215;
    75: op1_07_in15 = reg_0398;
    61: op1_07_in15 = imem00_in[3:0];
    56: op1_07_in15 = reg_0638;
    87: op1_07_in15 = reg_1004;
    76: op1_07_in15 = reg_0316;
    57: op1_07_in15 = reg_0530;
    77: op1_07_in15 = reg_0300;
    60: op1_07_in15 = imem04_in[11:8];
    58: op1_07_in15 = reg_0285;
    78: op1_07_in15 = imem05_in[3:0];
    70: op1_07_in15 = reg_0601;
    46: op1_07_in15 = reg_0006;
    51: op1_07_in15 = reg_0087;
    88: op1_07_in15 = reg_0957;
    79: op1_07_in15 = reg_0631;
    59: op1_07_in15 = reg_0030;
    48: op1_07_in15 = reg_0541;
    80: op1_07_in15 = reg_0491;
    62: op1_07_in15 = reg_0586;
    52: op1_07_in15 = reg_0527;
    81: op1_07_in15 = reg_1303;
    63: op1_07_in15 = reg_0318;
    82: op1_07_in15 = reg_1000;
    89: op1_07_in15 = reg_0348;
    83: op1_07_in15 = reg_0122;
    64: op1_07_in15 = imem04_in[3:0];
    84: op1_07_in15 = reg_0263;
    65: op1_07_in15 = reg_0114;
    85: op1_07_in15 = reg_0240;
    37: op1_07_in15 = reg_0465;
    90: op1_07_in15 = imem04_in[7:4];
    66: op1_07_in15 = reg_0175;
    91: op1_07_in15 = reg_0312;
    47: op1_07_in15 = reg_0519;
    67: op1_07_in15 = reg_1183;
    92: op1_07_in15 = reg_0305;
    93: op1_07_in15 = reg_0394;
    94: op1_07_in15 = reg_0730;
    95: op1_07_in15 = reg_0839;
    44: op1_07_in15 = reg_0221;
    96: op1_07_in15 = reg_0977;
    97: op1_07_in15 = reg_0782;
    98: op1_07_in15 = reg_0041;
    99: op1_07_in15 = reg_0112;
    100: op1_07_in15 = reg_0034;
    101: op1_07_in15 = reg_1369;
    102: op1_07_in15 = reg_0591;
    103: op1_07_in15 = reg_0060;
    104: op1_07_in15 = reg_0013;
    105: op1_07_in15 = reg_0166;
    106: op1_07_in15 = reg_0045;
    107: op1_07_in15 = imem03_in[11:8];
    108: op1_07_in15 = reg_0202;
    109: op1_07_in15 = reg_0881;
    110: op1_07_in15 = reg_0630;
    111: op1_07_in15 = reg_1032;
    112: op1_07_in15 = reg_1383;
    113: op1_07_in15 = reg_0405;
    114: op1_07_in15 = reg_0212;
    115: op1_07_in15 = reg_0970;
    116: op1_07_in15 = reg_0836;
    117: op1_07_in15 = imem03_in[7:4];
    118: op1_07_in15 = reg_0451;
    119: op1_07_in15 = reg_1282;
    42: op1_07_in15 = reg_0088;
    120: op1_07_in15 = reg_1456;
    121: op1_07_in15 = reg_0892;
    122: op1_07_in15 = imem07_in[3:0];
    123: op1_07_in15 = reg_0985;
    124: op1_07_in15 = reg_1170;
    125: op1_07_in15 = reg_1065;
    126: op1_07_in15 = reg_0717;
    127: op1_07_in15 = reg_0167;
    128: op1_07_in15 = reg_0462;
    129: op1_07_in15 = reg_0431;
    130: op1_07_in15 = reg_0556;
    131: op1_07_in15 = reg_0623;
    default: op1_07_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv15 = 1;
    55: op1_07_inv15 = 1;
    86: op1_07_inv15 = 1;
    54: op1_07_inv15 = 1;
    71: op1_07_inv15 = 1;
    75: op1_07_inv15 = 1;
    61: op1_07_inv15 = 1;
    57: op1_07_inv15 = 1;
    60: op1_07_inv15 = 1;
    58: op1_07_inv15 = 1;
    78: op1_07_inv15 = 1;
    80: op1_07_inv15 = 1;
    62: op1_07_inv15 = 1;
    63: op1_07_inv15 = 1;
    89: op1_07_inv15 = 1;
    65: op1_07_inv15 = 1;
    37: op1_07_inv15 = 1;
    47: op1_07_inv15 = 1;
    92: op1_07_inv15 = 1;
    93: op1_07_inv15 = 1;
    94: op1_07_inv15 = 1;
    95: op1_07_inv15 = 1;
    98: op1_07_inv15 = 1;
    102: op1_07_inv15 = 1;
    103: op1_07_inv15 = 1;
    104: op1_07_inv15 = 1;
    105: op1_07_inv15 = 1;
    106: op1_07_inv15 = 1;
    107: op1_07_inv15 = 1;
    108: op1_07_inv15 = 1;
    110: op1_07_inv15 = 1;
    111: op1_07_inv15 = 1;
    112: op1_07_inv15 = 1;
    113: op1_07_inv15 = 1;
    115: op1_07_inv15 = 1;
    42: op1_07_inv15 = 1;
    121: op1_07_inv15 = 1;
    125: op1_07_inv15 = 1;
    126: op1_07_inv15 = 1;
    default: op1_07_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in16 = reg_0175;
    53: op1_07_in16 = reg_0152;
    55: op1_07_in16 = reg_0624;
    86: op1_07_in16 = reg_0375;
    69: op1_07_in16 = reg_1214;
    73: op1_07_in16 = reg_0070;
    50: op1_07_in16 = reg_0351;
    108: op1_07_in16 = reg_0351;
    54: op1_07_in16 = reg_0255;
    71: op1_07_in16 = reg_0548;
    74: op1_07_in16 = reg_0109;
    68: op1_07_in16 = reg_1216;
    75: op1_07_in16 = reg_0141;
    61: op1_07_in16 = reg_0695;
    56: op1_07_in16 = reg_0188;
    109: op1_07_in16 = reg_0188;
    87: op1_07_in16 = reg_0719;
    76: op1_07_in16 = reg_0264;
    112: op1_07_in16 = reg_0264;
    57: op1_07_in16 = reg_0533;
    77: op1_07_in16 = reg_0090;
    60: op1_07_in16 = reg_0464;
    58: op1_07_in16 = reg_0738;
    78: op1_07_in16 = imem05_in[7:4];
    70: op1_07_in16 = reg_0130;
    46: op1_07_in16 = reg_0800;
    51: op1_07_in16 = reg_0519;
    88: op1_07_in16 = reg_0329;
    79: op1_07_in16 = reg_0449;
    59: op1_07_in16 = reg_0285;
    48: op1_07_in16 = reg_0539;
    80: op1_07_in16 = reg_1414;
    62: op1_07_in16 = reg_0527;
    52: op1_07_in16 = reg_0323;
    81: op1_07_in16 = reg_0194;
    63: op1_07_in16 = reg_0538;
    82: op1_07_in16 = reg_0999;
    89: op1_07_in16 = reg_0427;
    83: op1_07_in16 = reg_1100;
    64: op1_07_in16 = imem04_in[15:12];
    84: op1_07_in16 = reg_0181;
    65: op1_07_in16 = reg_0004;
    85: op1_07_in16 = reg_0799;
    37: op1_07_in16 = reg_0366;
    90: op1_07_in16 = reg_1368;
    66: op1_07_in16 = reg_0372;
    91: op1_07_in16 = reg_0142;
    47: op1_07_in16 = reg_0518;
    67: op1_07_in16 = reg_0225;
    121: op1_07_in16 = reg_0225;
    92: op1_07_in16 = reg_0862;
    93: op1_07_in16 = reg_1415;
    94: op1_07_in16 = reg_0316;
    95: op1_07_in16 = reg_0744;
    44: op1_07_in16 = reg_0445;
    96: op1_07_in16 = reg_0870;
    97: op1_07_in16 = reg_1437;
    98: op1_07_in16 = reg_0662;
    99: op1_07_in16 = reg_0382;
    100: op1_07_in16 = reg_0978;
    101: op1_07_in16 = reg_0034;
    102: op1_07_in16 = reg_0103;
    103: op1_07_in16 = reg_0059;
    104: op1_07_in16 = imem02_in[15:12];
    105: op1_07_in16 = reg_1290;
    106: op1_07_in16 = reg_1181;
    107: op1_07_in16 = reg_1145;
    110: op1_07_in16 = reg_1180;
    111: op1_07_in16 = reg_0635;
    113: op1_07_in16 = reg_0389;
    114: op1_07_in16 = reg_0213;
    115: op1_07_in16 = reg_0128;
    116: op1_07_in16 = reg_0835;
    117: op1_07_in16 = imem03_in[11:8];
    118: op1_07_in16 = reg_0452;
    119: op1_07_in16 = reg_0348;
    42: op1_07_in16 = reg_0283;
    120: op1_07_in16 = reg_0386;
    122: op1_07_in16 = imem07_in[7:4];
    123: op1_07_in16 = reg_0874;
    124: op1_07_in16 = reg_0087;
    125: op1_07_in16 = reg_0320;
    126: op1_07_in16 = reg_1302;
    127: op1_07_in16 = reg_1070;
    128: op1_07_in16 = reg_0531;
    129: op1_07_in16 = reg_0409;
    130: op1_07_in16 = reg_0178;
    131: op1_07_in16 = reg_0114;
    default: op1_07_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv16 = 1;
    53: op1_07_inv16 = 1;
    86: op1_07_inv16 = 1;
    69: op1_07_inv16 = 1;
    73: op1_07_inv16 = 1;
    50: op1_07_inv16 = 1;
    68: op1_07_inv16 = 1;
    75: op1_07_inv16 = 1;
    61: op1_07_inv16 = 1;
    87: op1_07_inv16 = 1;
    57: op1_07_inv16 = 1;
    60: op1_07_inv16 = 1;
    78: op1_07_inv16 = 1;
    51: op1_07_inv16 = 1;
    59: op1_07_inv16 = 1;
    48: op1_07_inv16 = 1;
    80: op1_07_inv16 = 1;
    62: op1_07_inv16 = 1;
    52: op1_07_inv16 = 1;
    81: op1_07_inv16 = 1;
    63: op1_07_inv16 = 1;
    82: op1_07_inv16 = 1;
    89: op1_07_inv16 = 1;
    65: op1_07_inv16 = 1;
    85: op1_07_inv16 = 1;
    90: op1_07_inv16 = 1;
    66: op1_07_inv16 = 1;
    94: op1_07_inv16 = 1;
    44: op1_07_inv16 = 1;
    96: op1_07_inv16 = 1;
    97: op1_07_inv16 = 1;
    98: op1_07_inv16 = 1;
    100: op1_07_inv16 = 1;
    106: op1_07_inv16 = 1;
    108: op1_07_inv16 = 1;
    110: op1_07_inv16 = 1;
    111: op1_07_inv16 = 1;
    117: op1_07_inv16 = 1;
    119: op1_07_inv16 = 1;
    121: op1_07_inv16 = 1;
    123: op1_07_inv16 = 1;
    124: op1_07_inv16 = 1;
    126: op1_07_inv16 = 1;
    127: op1_07_inv16 = 1;
    128: op1_07_inv16 = 1;
    130: op1_07_inv16 = 1;
    default: op1_07_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in17 = reg_0448;
    61: op1_07_in17 = reg_0448;
    53: op1_07_in17 = reg_0213;
    55: op1_07_in17 = reg_0526;
    86: op1_07_in17 = reg_0989;
    69: op1_07_in17 = reg_1077;
    73: op1_07_in17 = reg_0418;
    50: op1_07_in17 = reg_0352;
    54: op1_07_in17 = reg_0629;
    71: op1_07_in17 = reg_0787;
    74: op1_07_in17 = reg_0584;
    75: op1_07_in17 = reg_0584;
    68: op1_07_in17 = reg_1082;
    56: op1_07_in17 = reg_0189;
    87: op1_07_in17 = reg_0835;
    76: op1_07_in17 = reg_0859;
    57: op1_07_in17 = reg_1140;
    77: op1_07_in17 = reg_1486;
    60: op1_07_in17 = reg_0969;
    58: op1_07_in17 = reg_0593;
    78: op1_07_in17 = imem05_in[15:12];
    70: op1_07_in17 = reg_0243;
    46: op1_07_in17 = reg_0314;
    51: op1_07_in17 = reg_0484;
    88: op1_07_in17 = reg_1226;
    79: op1_07_in17 = reg_0861;
    59: op1_07_in17 = reg_0437;
    48: op1_07_in17 = reg_0938;
    80: op1_07_in17 = reg_1183;
    62: op1_07_in17 = reg_0568;
    52: op1_07_in17 = reg_0308;
    81: op1_07_in17 = reg_0617;
    63: op1_07_in17 = reg_0541;
    82: op1_07_in17 = imem03_in[7:4];
    89: op1_07_in17 = reg_1384;
    83: op1_07_in17 = reg_0464;
    64: op1_07_in17 = reg_0462;
    84: op1_07_in17 = reg_1369;
    65: op1_07_in17 = reg_0003;
    85: op1_07_in17 = reg_0864;
    37: op1_07_in17 = imem07_in[3:0];
    114: op1_07_in17 = imem07_in[3:0];
    90: op1_07_in17 = reg_0535;
    66: op1_07_in17 = reg_1253;
    91: op1_07_in17 = reg_1518;
    47: op1_07_in17 = reg_0123;
    67: op1_07_in17 = reg_0140;
    121: op1_07_in17 = reg_0140;
    92: op1_07_in17 = reg_1237;
    93: op1_07_in17 = reg_1096;
    94: op1_07_in17 = reg_0670;
    95: op1_07_in17 = reg_0054;
    44: op1_07_in17 = reg_0650;
    96: op1_07_in17 = reg_0860;
    97: op1_07_in17 = reg_0869;
    98: op1_07_in17 = reg_0590;
    99: op1_07_in17 = reg_1433;
    100: op1_07_in17 = reg_1233;
    101: op1_07_in17 = reg_1258;
    102: op1_07_in17 = reg_0114;
    103: op1_07_in17 = reg_0785;
    104: op1_07_in17 = reg_0879;
    105: op1_07_in17 = reg_0401;
    123: op1_07_in17 = reg_0401;
    106: op1_07_in17 = reg_1402;
    107: op1_07_in17 = reg_0198;
    108: op1_07_in17 = reg_0440;
    109: op1_07_in17 = reg_0201;
    110: op1_07_in17 = reg_1401;
    111: op1_07_in17 = reg_1152;
    112: op1_07_in17 = reg_0694;
    113: op1_07_in17 = reg_0057;
    115: op1_07_in17 = reg_0125;
    116: op1_07_in17 = reg_0117;
    117: op1_07_in17 = reg_0479;
    118: op1_07_in17 = reg_0698;
    119: op1_07_in17 = reg_0443;
    42: op1_07_in17 = reg_0042;
    120: op1_07_in17 = reg_0724;
    122: op1_07_in17 = reg_1095;
    124: op1_07_in17 = reg_0394;
    125: op1_07_in17 = reg_1143;
    126: op1_07_in17 = reg_1303;
    127: op1_07_in17 = reg_1169;
    128: op1_07_in17 = reg_0297;
    129: op1_07_in17 = reg_0089;
    130: op1_07_in17 = reg_0107;
    131: op1_07_in17 = reg_0028;
    default: op1_07_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_07_inv17 = 1;
    55: op1_07_inv17 = 1;
    69: op1_07_inv17 = 1;
    73: op1_07_inv17 = 1;
    54: op1_07_inv17 = 1;
    74: op1_07_inv17 = 1;
    76: op1_07_inv17 = 1;
    57: op1_07_inv17 = 1;
    77: op1_07_inv17 = 1;
    46: op1_07_inv17 = 1;
    79: op1_07_inv17 = 1;
    48: op1_07_inv17 = 1;
    62: op1_07_inv17 = 1;
    81: op1_07_inv17 = 1;
    82: op1_07_inv17 = 1;
    89: op1_07_inv17 = 1;
    84: op1_07_inv17 = 1;
    65: op1_07_inv17 = 1;
    85: op1_07_inv17 = 1;
    37: op1_07_inv17 = 1;
    90: op1_07_inv17 = 1;
    66: op1_07_inv17 = 1;
    92: op1_07_inv17 = 1;
    44: op1_07_inv17 = 1;
    96: op1_07_inv17 = 1;
    99: op1_07_inv17 = 1;
    101: op1_07_inv17 = 1;
    102: op1_07_inv17 = 1;
    106: op1_07_inv17 = 1;
    110: op1_07_inv17 = 1;
    111: op1_07_inv17 = 1;
    112: op1_07_inv17 = 1;
    113: op1_07_inv17 = 1;
    114: op1_07_inv17 = 1;
    118: op1_07_inv17 = 1;
    119: op1_07_inv17 = 1;
    120: op1_07_inv17 = 1;
    122: op1_07_inv17 = 1;
    123: op1_07_inv17 = 1;
    124: op1_07_inv17 = 1;
    125: op1_07_inv17 = 1;
    126: op1_07_inv17 = 1;
    129: op1_07_inv17 = 1;
    130: op1_07_inv17 = 1;
    131: op1_07_inv17 = 1;
    default: op1_07_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in18 = reg_1256;
    103: op1_07_in18 = reg_1256;
    53: op1_07_in18 = imem06_in[3:0];
    55: op1_07_in18 = imem06_in[7:4];
    86: op1_07_in18 = reg_0220;
    69: op1_07_in18 = reg_0676;
    73: op1_07_in18 = reg_0873;
    50: op1_07_in18 = reg_0089;
    54: op1_07_in18 = reg_0606;
    71: op1_07_in18 = reg_0420;
    74: op1_07_in18 = reg_0526;
    68: op1_07_in18 = reg_0598;
    75: op1_07_in18 = reg_0568;
    61: op1_07_in18 = reg_0260;
    56: op1_07_in18 = reg_0410;
    87: op1_07_in18 = reg_0339;
    76: op1_07_in18 = reg_0869;
    96: op1_07_in18 = reg_0869;
    57: op1_07_in18 = reg_1139;
    77: op1_07_in18 = reg_0275;
    60: op1_07_in18 = reg_0798;
    58: op1_07_in18 = reg_0592;
    78: op1_07_in18 = reg_1180;
    70: op1_07_in18 = reg_0118;
    46: op1_07_in18 = reg_0732;
    88: op1_07_in18 = reg_1208;
    79: op1_07_in18 = reg_0317;
    59: op1_07_in18 = reg_0002;
    48: op1_07_in18 = reg_0168;
    80: op1_07_in18 = reg_0140;
    62: op1_07_in18 = reg_1225;
    52: op1_07_in18 = reg_0271;
    81: op1_07_in18 = reg_0345;
    63: op1_07_in18 = reg_0539;
    82: op1_07_in18 = reg_0177;
    89: op1_07_in18 = reg_1383;
    83: op1_07_in18 = reg_1034;
    64: op1_07_in18 = reg_1077;
    84: op1_07_in18 = reg_0493;
    65: op1_07_in18 = reg_0052;
    85: op1_07_in18 = reg_0449;
    37: op1_07_in18 = reg_0404;
    90: op1_07_in18 = reg_0264;
    66: op1_07_in18 = reg_1254;
    91: op1_07_in18 = reg_0048;
    67: op1_07_in18 = reg_1350;
    92: op1_07_in18 = reg_0117;
    93: op1_07_in18 = reg_0922;
    94: op1_07_in18 = reg_0247;
    95: op1_07_in18 = reg_0125;
    44: op1_07_in18 = reg_0045;
    97: op1_07_in18 = reg_1504;
    98: op1_07_in18 = reg_0133;
    99: op1_07_in18 = reg_0684;
    100: op1_07_in18 = reg_1082;
    101: op1_07_in18 = reg_0531;
    112: op1_07_in18 = reg_0531;
    102: op1_07_in18 = reg_0051;
    104: op1_07_in18 = reg_0055;
    105: op1_07_in18 = reg_0548;
    106: op1_07_in18 = reg_1401;
    107: op1_07_in18 = reg_0783;
    108: op1_07_in18 = reg_0058;
    109: op1_07_in18 = reg_0405;
    110: op1_07_in18 = reg_0940;
    111: op1_07_in18 = reg_0985;
    113: op1_07_in18 = reg_0026;
    114: op1_07_in18 = imem07_in[11:8];
    115: op1_07_in18 = reg_0382;
    116: op1_07_in18 = reg_0633;
    117: op1_07_in18 = reg_0759;
    118: op1_07_in18 = reg_0835;
    119: op1_07_in18 = reg_0263;
    42: op1_07_in18 = reg_0044;
    120: op1_07_in18 = reg_0933;
    121: op1_07_in18 = reg_0661;
    122: op1_07_in18 = reg_0135;
    123: op1_07_in18 = reg_0163;
    124: op1_07_in18 = reg_0157;
    125: op1_07_in18 = reg_0256;
    126: op1_07_in18 = reg_0619;
    127: op1_07_in18 = reg_0477;
    128: op1_07_in18 = reg_1215;
    129: op1_07_in18 = reg_0384;
    130: op1_07_in18 = reg_0559;
    131: op1_07_in18 = reg_0235;
    default: op1_07_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv18 = 1;
    69: op1_07_inv18 = 1;
    54: op1_07_inv18 = 1;
    71: op1_07_inv18 = 1;
    68: op1_07_inv18 = 1;
    56: op1_07_inv18 = 1;
    87: op1_07_inv18 = 1;
    76: op1_07_inv18 = 1;
    77: op1_07_inv18 = 1;
    78: op1_07_inv18 = 1;
    70: op1_07_inv18 = 1;
    88: op1_07_inv18 = 1;
    79: op1_07_inv18 = 1;
    48: op1_07_inv18 = 1;
    62: op1_07_inv18 = 1;
    63: op1_07_inv18 = 1;
    82: op1_07_inv18 = 1;
    83: op1_07_inv18 = 1;
    64: op1_07_inv18 = 1;
    84: op1_07_inv18 = 1;
    66: op1_07_inv18 = 1;
    67: op1_07_inv18 = 1;
    94: op1_07_inv18 = 1;
    44: op1_07_inv18 = 1;
    96: op1_07_inv18 = 1;
    97: op1_07_inv18 = 1;
    98: op1_07_inv18 = 1;
    99: op1_07_inv18 = 1;
    100: op1_07_inv18 = 1;
    101: op1_07_inv18 = 1;
    102: op1_07_inv18 = 1;
    105: op1_07_inv18 = 1;
    106: op1_07_inv18 = 1;
    110: op1_07_inv18 = 1;
    111: op1_07_inv18 = 1;
    112: op1_07_inv18 = 1;
    113: op1_07_inv18 = 1;
    115: op1_07_inv18 = 1;
    117: op1_07_inv18 = 1;
    119: op1_07_inv18 = 1;
    42: op1_07_inv18 = 1;
    120: op1_07_inv18 = 1;
    123: op1_07_inv18 = 1;
    128: op1_07_inv18 = 1;
    129: op1_07_inv18 = 1;
    default: op1_07_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in19 = reg_1070;
    53: op1_07_in19 = imem07_in[7:4];
    55: op1_07_in19 = reg_0015;
    86: op1_07_in19 = reg_1231;
    69: op1_07_in19 = reg_0797;
    60: op1_07_in19 = reg_0797;
    73: op1_07_in19 = imem05_in[11:8];
    50: op1_07_in19 = reg_0609;
    54: op1_07_in19 = reg_0587;
    71: op1_07_in19 = reg_0468;
    74: op1_07_in19 = reg_0527;
    68: op1_07_in19 = reg_0471;
    64: op1_07_in19 = reg_0471;
    75: op1_07_in19 = reg_0295;
    61: op1_07_in19 = reg_0241;
    56: op1_07_in19 = reg_0134;
    87: op1_07_in19 = reg_1237;
    76: op1_07_in19 = reg_0116;
    57: op1_07_in19 = imem02_in[7:4];
    77: op1_07_in19 = reg_0274;
    58: op1_07_in19 = reg_0361;
    78: op1_07_in19 = reg_0938;
    70: op1_07_in19 = reg_0151;
    46: op1_07_in19 = reg_0675;
    88: op1_07_in19 = reg_0479;
    79: op1_07_in19 = reg_1435;
    59: op1_07_in19 = reg_0053;
    131: op1_07_in19 = reg_0053;
    48: op1_07_in19 = reg_0449;
    80: op1_07_in19 = reg_0309;
    62: op1_07_in19 = reg_0244;
    52: op1_07_in19 = reg_0046;
    81: op1_07_in19 = reg_0296;
    63: op1_07_in19 = reg_0243;
    82: op1_07_in19 = reg_0198;
    89: op1_07_in19 = reg_0181;
    83: op1_07_in19 = reg_0448;
    84: op1_07_in19 = reg_1216;
    65: op1_07_in19 = reg_0518;
    85: op1_07_in19 = reg_0206;
    37: op1_07_in19 = reg_0621;
    90: op1_07_in19 = reg_1198;
    66: op1_07_in19 = reg_1068;
    91: op1_07_in19 = reg_0880;
    67: op1_07_in19 = reg_0139;
    92: op1_07_in19 = reg_0209;
    125: op1_07_in19 = reg_0209;
    93: op1_07_in19 = reg_0894;
    94: op1_07_in19 = reg_0751;
    95: op1_07_in19 = reg_0105;
    44: op1_07_in19 = reg_0332;
    96: op1_07_in19 = reg_1505;
    97: op1_07_in19 = reg_0109;
    98: op1_07_in19 = imem02_in[11:8];
    99: op1_07_in19 = reg_0381;
    100: op1_07_in19 = reg_0796;
    101: op1_07_in19 = reg_0297;
    112: op1_07_in19 = reg_0297;
    102: op1_07_in19 = reg_0001;
    103: op1_07_in19 = reg_0902;
    104: op1_07_in19 = reg_0497;
    105: op1_07_in19 = reg_0610;
    106: op1_07_in19 = reg_0937;
    127: op1_07_in19 = reg_0937;
    107: op1_07_in19 = reg_0311;
    108: op1_07_in19 = imem01_in[11:8];
    109: op1_07_in19 = reg_0388;
    110: op1_07_in19 = reg_0266;
    111: op1_07_in19 = reg_0548;
    113: op1_07_in19 = reg_0917;
    114: op1_07_in19 = imem07_in[15:12];
    115: op1_07_in19 = reg_1433;
    116: op1_07_in19 = reg_0019;
    117: op1_07_in19 = reg_0154;
    118: op1_07_in19 = reg_1340;
    119: op1_07_in19 = reg_0338;
    42: op1_07_in19 = reg_0041;
    120: op1_07_in19 = reg_0606;
    121: op1_07_in19 = reg_0442;
    122: op1_07_in19 = reg_0310;
    123: op1_07_in19 = reg_0258;
    124: op1_07_in19 = reg_0924;
    126: op1_07_in19 = reg_0568;
    128: op1_07_in19 = reg_1214;
    129: op1_07_in19 = imem01_in[3:0];
    130: op1_07_in19 = reg_1282;
    default: op1_07_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv19 = 1;
    53: op1_07_inv19 = 1;
    55: op1_07_inv19 = 1;
    86: op1_07_inv19 = 1;
    73: op1_07_inv19 = 1;
    50: op1_07_inv19 = 1;
    54: op1_07_inv19 = 1;
    74: op1_07_inv19 = 1;
    56: op1_07_inv19 = 1;
    87: op1_07_inv19 = 1;
    76: op1_07_inv19 = 1;
    77: op1_07_inv19 = 1;
    78: op1_07_inv19 = 1;
    70: op1_07_inv19 = 1;
    59: op1_07_inv19 = 1;
    48: op1_07_inv19 = 1;
    62: op1_07_inv19 = 1;
    52: op1_07_inv19 = 1;
    81: op1_07_inv19 = 1;
    82: op1_07_inv19 = 1;
    89: op1_07_inv19 = 1;
    64: op1_07_inv19 = 1;
    65: op1_07_inv19 = 1;
    85: op1_07_inv19 = 1;
    37: op1_07_inv19 = 1;
    91: op1_07_inv19 = 1;
    92: op1_07_inv19 = 1;
    93: op1_07_inv19 = 1;
    94: op1_07_inv19 = 1;
    96: op1_07_inv19 = 1;
    98: op1_07_inv19 = 1;
    99: op1_07_inv19 = 1;
    101: op1_07_inv19 = 1;
    103: op1_07_inv19 = 1;
    106: op1_07_inv19 = 1;
    107: op1_07_inv19 = 1;
    108: op1_07_inv19 = 1;
    111: op1_07_inv19 = 1;
    113: op1_07_inv19 = 1;
    114: op1_07_inv19 = 1;
    116: op1_07_inv19 = 1;
    119: op1_07_inv19 = 1;
    122: op1_07_inv19 = 1;
    124: op1_07_inv19 = 1;
    125: op1_07_inv19 = 1;
    131: op1_07_inv19 = 1;
    default: op1_07_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in20 = reg_1069;
    53: op1_07_in20 = reg_1095;
    55: op1_07_in20 = reg_0017;
    86: op1_07_in20 = reg_0107;
    69: op1_07_in20 = reg_0936;
    73: op1_07_in20 = reg_0274;
    50: op1_07_in20 = imem01_in[11:8];
    113: op1_07_in20 = imem01_in[11:8];
    129: op1_07_in20 = imem01_in[11:8];
    54: op1_07_in20 = reg_0530;
    71: op1_07_in20 = reg_0715;
    74: op1_07_in20 = reg_0296;
    68: op1_07_in20 = reg_0796;
    75: op1_07_in20 = reg_0119;
    61: op1_07_in20 = reg_0469;
    56: op1_07_in20 = reg_0388;
    87: op1_07_in20 = reg_0211;
    76: op1_07_in20 = reg_0617;
    57: op1_07_in20 = reg_0666;
    77: op1_07_in20 = reg_0243;
    60: op1_07_in20 = reg_0369;
    58: op1_07_in20 = reg_0519;
    78: op1_07_in20 = reg_0183;
    70: op1_07_in20 = reg_0317;
    46: op1_07_in20 = reg_0216;
    88: op1_07_in20 = reg_0478;
    79: op1_07_in20 = reg_1064;
    59: op1_07_in20 = reg_0518;
    48: op1_07_in20 = reg_0040;
    80: op1_07_in20 = reg_0223;
    62: op1_07_in20 = reg_0270;
    52: op1_07_in20 = reg_0212;
    81: op1_07_in20 = reg_0295;
    63: op1_07_in20 = reg_0240;
    82: op1_07_in20 = reg_0145;
    89: op1_07_in20 = reg_1368;
    83: op1_07_in20 = reg_1255;
    64: op1_07_in20 = reg_0795;
    84: op1_07_in20 = reg_0574;
    65: op1_07_in20 = reg_0123;
    85: op1_07_in20 = reg_1105;
    37: op1_07_in20 = reg_0103;
    90: op1_07_in20 = reg_0281;
    66: op1_07_in20 = reg_0258;
    91: op1_07_in20 = reg_0884;
    67: op1_07_in20 = reg_0777;
    92: op1_07_in20 = reg_0065;
    93: op1_07_in20 = reg_1056;
    94: op1_07_in20 = reg_0720;
    95: op1_07_in20 = reg_0876;
    44: op1_07_in20 = reg_0316;
    96: op1_07_in20 = reg_1504;
    97: op1_07_in20 = reg_0716;
    98: op1_07_in20 = reg_0975;
    99: op1_07_in20 = reg_0306;
    100: op1_07_in20 = reg_0199;
    101: op1_07_in20 = reg_0552;
    102: op1_07_in20 = reg_0483;
    103: op1_07_in20 = reg_0401;
    104: op1_07_in20 = reg_1260;
    105: op1_07_in20 = reg_0239;
    106: op1_07_in20 = reg_0418;
    110: op1_07_in20 = reg_0418;
    107: op1_07_in20 = reg_0789;
    108: op1_07_in20 = reg_0871;
    109: op1_07_in20 = reg_0387;
    111: op1_07_in20 = reg_0242;
    112: op1_07_in20 = reg_1083;
    114: op1_07_in20 = reg_0394;
    115: op1_07_in20 = reg_0684;
    116: op1_07_in20 = reg_0021;
    117: op1_07_in20 = reg_0573;
    118: op1_07_in20 = reg_1151;
    119: op1_07_in20 = reg_0534;
    42: op1_07_in20 = reg_0012;
    120: op1_07_in20 = reg_1235;
    121: op1_07_in20 = reg_0437;
    122: op1_07_in20 = reg_0457;
    123: op1_07_in20 = reg_0747;
    124: op1_07_in20 = reg_0139;
    125: op1_07_in20 = reg_0538;
    126: op1_07_in20 = reg_0570;
    127: op1_07_in20 = reg_0318;
    128: op1_07_in20 = reg_0094;
    130: op1_07_in20 = reg_0348;
    131: op1_07_in20 = reg_0404;
    default: op1_07_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv20 = 1;
    73: op1_07_inv20 = 1;
    54: op1_07_inv20 = 1;
    71: op1_07_inv20 = 1;
    68: op1_07_inv20 = 1;
    75: op1_07_inv20 = 1;
    61: op1_07_inv20 = 1;
    56: op1_07_inv20 = 1;
    76: op1_07_inv20 = 1;
    77: op1_07_inv20 = 1;
    60: op1_07_inv20 = 1;
    78: op1_07_inv20 = 1;
    70: op1_07_inv20 = 1;
    46: op1_07_inv20 = 1;
    59: op1_07_inv20 = 1;
    80: op1_07_inv20 = 1;
    52: op1_07_inv20 = 1;
    63: op1_07_inv20 = 1;
    64: op1_07_inv20 = 1;
    90: op1_07_inv20 = 1;
    66: op1_07_inv20 = 1;
    91: op1_07_inv20 = 1;
    93: op1_07_inv20 = 1;
    98: op1_07_inv20 = 1;
    101: op1_07_inv20 = 1;
    104: op1_07_inv20 = 1;
    110: op1_07_inv20 = 1;
    112: op1_07_inv20 = 1;
    116: op1_07_inv20 = 1;
    118: op1_07_inv20 = 1;
    119: op1_07_inv20 = 1;
    42: op1_07_inv20 = 1;
    120: op1_07_inv20 = 1;
    124: op1_07_inv20 = 1;
    125: op1_07_inv20 = 1;
    130: op1_07_inv20 = 1;
    default: op1_07_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in21 = reg_0166;
    53: op1_07_in21 = reg_1057;
    55: op1_07_in21 = reg_1150;
    86: op1_07_in21 = reg_0504;
    69: op1_07_in21 = reg_0451;
    73: op1_07_in21 = reg_1348;
    127: op1_07_in21 = reg_1348;
    50: op1_07_in21 = reg_1032;
    54: op1_07_in21 = reg_0531;
    71: op1_07_in21 = reg_1457;
    74: op1_07_in21 = reg_0295;
    68: op1_07_in21 = reg_0452;
    75: op1_07_in21 = reg_0371;
    61: op1_07_in21 = reg_0430;
    56: op1_07_in21 = reg_0057;
    87: op1_07_in21 = reg_0210;
    116: op1_07_in21 = reg_0210;
    76: op1_07_in21 = reg_0569;
    57: op1_07_in21 = reg_0475;
    77: op1_07_in21 = reg_0602;
    60: op1_07_in21 = reg_0305;
    58: op1_07_in21 = reg_0520;
    59: op1_07_in21 = reg_0520;
    78: op1_07_in21 = reg_0090;
    70: op1_07_in21 = reg_0037;
    46: op1_07_in21 = reg_0288;
    88: op1_07_in21 = reg_0288;
    79: op1_07_in21 = reg_0730;
    48: op1_07_in21 = reg_0195;
    80: op1_07_in21 = reg_0775;
    62: op1_07_in21 = reg_0269;
    52: op1_07_in21 = reg_0213;
    81: op1_07_in21 = reg_1179;
    63: op1_07_in21 = imem05_in[7:4];
    82: op1_07_in21 = reg_0989;
    89: op1_07_in21 = reg_0264;
    83: op1_07_in21 = reg_0785;
    64: op1_07_in21 = reg_0904;
    84: op1_07_in21 = reg_0454;
    100: op1_07_in21 = reg_0454;
    85: op1_07_in21 = reg_0268;
    37: op1_07_in21 = reg_0361;
    90: op1_07_in21 = reg_1082;
    66: op1_07_in21 = reg_0420;
    92: op1_07_in21 = reg_0420;
    91: op1_07_in21 = reg_1149;
    67: op1_07_in21 = reg_0031;
    93: op1_07_in21 = reg_0170;
    94: op1_07_in21 = reg_0141;
    95: op1_07_in21 = reg_0878;
    115: op1_07_in21 = reg_0878;
    44: op1_07_in21 = reg_0539;
    96: op1_07_in21 = reg_0115;
    97: op1_07_in21 = reg_0636;
    98: op1_07_in21 = reg_0845;
    99: op1_07_in21 = reg_1098;
    101: op1_07_in21 = reg_1233;
    102: op1_07_in21 = reg_1182;
    103: op1_07_in21 = reg_0463;
    104: op1_07_in21 = reg_1207;
    105: op1_07_in21 = reg_0238;
    106: op1_07_in21 = reg_0302;
    107: op1_07_in21 = reg_0142;
    108: op1_07_in21 = reg_0985;
    113: op1_07_in21 = reg_0985;
    109: op1_07_in21 = reg_0027;
    110: op1_07_in21 = reg_0303;
    111: op1_07_in21 = reg_0468;
    112: op1_07_in21 = reg_1203;
    114: op1_07_in21 = reg_0478;
    117: op1_07_in21 = reg_0198;
    118: op1_07_in21 = reg_0209;
    119: op1_07_in21 = reg_1368;
    42: op1_07_in21 = reg_0662;
    120: op1_07_in21 = reg_0254;
    121: op1_07_in21 = reg_0591;
    122: op1_07_in21 = reg_1349;
    123: op1_07_in21 = reg_0743;
    124: op1_07_in21 = reg_0224;
    125: op1_07_in21 = reg_0367;
    126: op1_07_in21 = reg_1225;
    128: op1_07_in21 = reg_1147;
    129: op1_07_in21 = reg_0047;
    130: op1_07_in21 = reg_0443;
    131: op1_07_in21 = reg_0002;
    default: op1_07_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    54: op1_07_inv21 = 1;
    71: op1_07_inv21 = 1;
    68: op1_07_inv21 = 1;
    61: op1_07_inv21 = 1;
    57: op1_07_inv21 = 1;
    77: op1_07_inv21 = 1;
    60: op1_07_inv21 = 1;
    58: op1_07_inv21 = 1;
    78: op1_07_inv21 = 1;
    70: op1_07_inv21 = 1;
    46: op1_07_inv21 = 1;
    48: op1_07_inv21 = 1;
    80: op1_07_inv21 = 1;
    62: op1_07_inv21 = 1;
    81: op1_07_inv21 = 1;
    63: op1_07_inv21 = 1;
    82: op1_07_inv21 = 1;
    89: op1_07_inv21 = 1;
    83: op1_07_inv21 = 1;
    84: op1_07_inv21 = 1;
    85: op1_07_inv21 = 1;
    37: op1_07_inv21 = 1;
    90: op1_07_inv21 = 1;
    66: op1_07_inv21 = 1;
    91: op1_07_inv21 = 1;
    94: op1_07_inv21 = 1;
    44: op1_07_inv21 = 1;
    97: op1_07_inv21 = 1;
    99: op1_07_inv21 = 1;
    101: op1_07_inv21 = 1;
    102: op1_07_inv21 = 1;
    104: op1_07_inv21 = 1;
    106: op1_07_inv21 = 1;
    109: op1_07_inv21 = 1;
    110: op1_07_inv21 = 1;
    111: op1_07_inv21 = 1;
    114: op1_07_inv21 = 1;
    117: op1_07_inv21 = 1;
    120: op1_07_inv21 = 1;
    121: op1_07_inv21 = 1;
    123: op1_07_inv21 = 1;
    124: op1_07_inv21 = 1;
    125: op1_07_inv21 = 1;
    126: op1_07_inv21 = 1;
    130: op1_07_inv21 = 1;
    default: op1_07_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in22 = reg_0715;
    53: op1_07_in22 = reg_0998;
    55: op1_07_in22 = reg_1095;
    86: op1_07_in22 = reg_0507;
    69: op1_07_in22 = reg_0369;
    73: op1_07_in22 = reg_0828;
    77: op1_07_in22 = reg_0828;
    50: op1_07_in22 = reg_0788;
    54: op1_07_in22 = reg_0256;
    71: op1_07_in22 = reg_0384;
    74: op1_07_in22 = reg_0419;
    68: op1_07_in22 = reg_0305;
    75: op1_07_in22 = reg_0215;
    61: op1_07_in22 = reg_0438;
    56: op1_07_in22 = reg_0059;
    87: op1_07_in22 = reg_0748;
    76: op1_07_in22 = reg_0289;
    57: op1_07_in22 = reg_0433;
    60: op1_07_in22 = reg_0319;
    58: op1_07_in22 = reg_0123;
    78: op1_07_in22 = reg_0873;
    70: op1_07_in22 = reg_0780;
    46: op1_07_in22 = reg_0707;
    88: op1_07_in22 = reg_1325;
    79: op1_07_in22 = reg_1508;
    48: op1_07_in22 = reg_0931;
    80: op1_07_in22 = reg_0663;
    62: op1_07_in22 = reg_0213;
    52: op1_07_in22 = reg_0015;
    81: op1_07_in22 = imem07_in[15:12];
    63: op1_07_in22 = imem05_in[15:12];
    82: op1_07_in22 = reg_1003;
    89: op1_07_in22 = reg_0252;
    83: op1_07_in22 = reg_0258;
    64: op1_07_in22 = reg_0199;
    84: op1_07_in22 = reg_0451;
    100: op1_07_in22 = reg_0451;
    85: op1_07_in22 = reg_0192;
    37: op1_07_in22 = reg_0519;
    90: op1_07_in22 = reg_0471;
    66: op1_07_in22 = reg_0241;
    91: op1_07_in22 = reg_0458;
    67: op1_07_in22 = reg_0465;
    92: op1_07_in22 = reg_1503;
    93: op1_07_in22 = reg_0489;
    94: op1_07_in22 = reg_0526;
    95: op1_07_in22 = reg_0897;
    44: op1_07_in22 = reg_0492;
    96: op1_07_in22 = reg_0110;
    97: op1_07_in22 = reg_0141;
    98: op1_07_in22 = reg_0253;
    99: op1_07_in22 = reg_0024;
    101: op1_07_in22 = reg_0407;
    103: op1_07_in22 = reg_0242;
    104: op1_07_in22 = reg_0381;
    105: op1_07_in22 = reg_0612;
    106: op1_07_in22 = reg_0872;
    107: op1_07_in22 = reg_0349;
    108: op1_07_in22 = reg_0547;
    109: op1_07_in22 = reg_0874;
    110: op1_07_in22 = reg_0794;
    111: op1_07_in22 = reg_0469;
    112: op1_07_in22 = reg_1198;
    113: op1_07_in22 = reg_0463;
    114: op1_07_in22 = reg_1060;
    115: op1_07_in22 = reg_1492;
    116: op1_07_in22 = reg_0370;
    117: op1_07_in22 = reg_0823;
    118: op1_07_in22 = reg_0095;
    119: op1_07_in22 = reg_0493;
    42: op1_07_in22 = reg_0628;
    120: op1_07_in22 = reg_0533;
    121: op1_07_in22 = reg_0028;
    122: op1_07_in22 = reg_0923;
    123: op1_07_in22 = reg_0238;
    124: op1_07_in22 = reg_0777;
    125: op1_07_in22 = reg_0136;
    126: op1_07_in22 = reg_0522;
    127: op1_07_in22 = reg_0589;
    128: op1_07_in22 = reg_0414;
    129: op1_07_in22 = reg_0577;
    130: op1_07_in22 = reg_0129;
    131: op1_07_in22 = reg_0484;
    default: op1_07_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv22 = 1;
    53: op1_07_inv22 = 1;
    55: op1_07_inv22 = 1;
    86: op1_07_inv22 = 1;
    69: op1_07_inv22 = 1;
    50: op1_07_inv22 = 1;
    71: op1_07_inv22 = 1;
    74: op1_07_inv22 = 1;
    75: op1_07_inv22 = 1;
    56: op1_07_inv22 = 1;
    87: op1_07_inv22 = 1;
    76: op1_07_inv22 = 1;
    57: op1_07_inv22 = 1;
    77: op1_07_inv22 = 1;
    58: op1_07_inv22 = 1;
    78: op1_07_inv22 = 1;
    46: op1_07_inv22 = 1;
    88: op1_07_inv22 = 1;
    79: op1_07_inv22 = 1;
    48: op1_07_inv22 = 1;
    62: op1_07_inv22 = 1;
    52: op1_07_inv22 = 1;
    81: op1_07_inv22 = 1;
    89: op1_07_inv22 = 1;
    83: op1_07_inv22 = 1;
    64: op1_07_inv22 = 1;
    85: op1_07_inv22 = 1;
    90: op1_07_inv22 = 1;
    66: op1_07_inv22 = 1;
    91: op1_07_inv22 = 1;
    67: op1_07_inv22 = 1;
    92: op1_07_inv22 = 1;
    93: op1_07_inv22 = 1;
    94: op1_07_inv22 = 1;
    96: op1_07_inv22 = 1;
    97: op1_07_inv22 = 1;
    98: op1_07_inv22 = 1;
    99: op1_07_inv22 = 1;
    100: op1_07_inv22 = 1;
    103: op1_07_inv22 = 1;
    104: op1_07_inv22 = 1;
    105: op1_07_inv22 = 1;
    107: op1_07_inv22 = 1;
    110: op1_07_inv22 = 1;
    111: op1_07_inv22 = 1;
    117: op1_07_inv22 = 1;
    119: op1_07_inv22 = 1;
    121: op1_07_inv22 = 1;
    122: op1_07_inv22 = 1;
    124: op1_07_inv22 = 1;
    125: op1_07_inv22 = 1;
    127: op1_07_inv22 = 1;
    128: op1_07_inv22 = 1;
    129: op1_07_inv22 = 1;
    130: op1_07_inv22 = 1;
    default: op1_07_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in23 = reg_0572;
    53: op1_07_in23 = reg_0245;
    55: op1_07_in23 = reg_1055;
    86: op1_07_in23 = reg_0481;
    69: op1_07_in23 = reg_0698;
    73: op1_07_in23 = reg_0377;
    50: op1_07_in23 = reg_0785;
    54: op1_07_in23 = reg_1139;
    71: op1_07_in23 = reg_0360;
    74: op1_07_in23 = reg_0244;
    68: op1_07_in23 = reg_0837;
    60: op1_07_in23 = reg_0837;
    75: op1_07_in23 = reg_1170;
    62: op1_07_in23 = reg_1170;
    61: op1_07_in23 = reg_0363;
    56: op1_07_in23 = reg_0026;
    87: op1_07_in23 = reg_1430;
    76: op1_07_in23 = imem07_in[7:4];
    57: op1_07_in23 = reg_0429;
    77: op1_07_in23 = reg_0038;
    116: op1_07_in23 = reg_0038;
    58: op1_07_in23 = reg_1182;
    131: op1_07_in23 = reg_1182;
    78: op1_07_in23 = reg_0631;
    70: op1_07_in23 = reg_0906;
    46: op1_07_in23 = reg_0378;
    88: op1_07_in23 = reg_0425;
    79: op1_07_in23 = reg_0397;
    48: op1_07_in23 = imem06_in[3:0];
    80: op1_07_in23 = reg_0441;
    52: op1_07_in23 = reg_0018;
    81: op1_07_in23 = reg_0786;
    63: op1_07_in23 = reg_0039;
    82: op1_07_in23 = reg_0070;
    89: op1_07_in23 = reg_1338;
    83: op1_07_in23 = reg_0746;
    64: op1_07_in23 = reg_0340;
    84: op1_07_in23 = reg_0033;
    85: op1_07_in23 = reg_0925;
    37: op1_07_in23 = reg_0521;
    90: op1_07_in23 = reg_0342;
    66: op1_07_in23 = reg_0743;
    91: op1_07_in23 = reg_0707;
    67: op1_07_in23 = reg_0623;
    92: op1_07_in23 = reg_0020;
    93: op1_07_in23 = reg_0366;
    94: op1_07_in23 = reg_0527;
    95: op1_07_in23 = reg_1098;
    115: op1_07_in23 = reg_1098;
    44: op1_07_in23 = imem05_in[3:0];
    96: op1_07_in23 = reg_0617;
    97: op1_07_in23 = reg_0568;
    98: op1_07_in23 = reg_1344;
    99: op1_07_in23 = reg_0168;
    100: op1_07_in23 = reg_1419;
    101: op1_07_in23 = reg_0199;
    103: op1_07_in23 = reg_0830;
    104: op1_07_in23 = reg_0802;
    105: op1_07_in23 = reg_1457;
    106: op1_07_in23 = reg_0344;
    107: op1_07_in23 = reg_1313;
    108: op1_07_in23 = reg_0260;
    109: op1_07_in23 = reg_1290;
    110: op1_07_in23 = reg_0799;
    111: op1_07_in23 = reg_0430;
    112: op1_07_in23 = reg_1215;
    113: op1_07_in23 = reg_0163;
    114: op1_07_in23 = reg_1315;
    117: op1_07_in23 = reg_0311;
    118: op1_07_in23 = reg_1503;
    119: op1_07_in23 = reg_0088;
    42: op1_07_in23 = reg_0606;
    120: op1_07_in23 = reg_0436;
    121: op1_07_in23 = reg_0052;
    122: op1_07_in23 = reg_0777;
    123: op1_07_in23 = reg_0241;
    124: op1_07_in23 = reg_0030;
    125: op1_07_in23 = reg_0702;
    126: op1_07_in23 = reg_0022;
    127: op1_07_in23 = reg_0828;
    128: op1_07_in23 = reg_1004;
    129: op1_07_in23 = reg_0871;
    130: op1_07_in23 = reg_0795;
    default: op1_07_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_07_inv23 = 1;
    73: op1_07_inv23 = 1;
    71: op1_07_inv23 = 1;
    68: op1_07_inv23 = 1;
    76: op1_07_inv23 = 1;
    57: op1_07_inv23 = 1;
    77: op1_07_inv23 = 1;
    60: op1_07_inv23 = 1;
    58: op1_07_inv23 = 1;
    78: op1_07_inv23 = 1;
    46: op1_07_inv23 = 1;
    80: op1_07_inv23 = 1;
    81: op1_07_inv23 = 1;
    82: op1_07_inv23 = 1;
    84: op1_07_inv23 = 1;
    37: op1_07_inv23 = 1;
    67: op1_07_inv23 = 1;
    92: op1_07_inv23 = 1;
    94: op1_07_inv23 = 1;
    44: op1_07_inv23 = 1;
    96: op1_07_inv23 = 1;
    97: op1_07_inv23 = 1;
    98: op1_07_inv23 = 1;
    99: op1_07_inv23 = 1;
    101: op1_07_inv23 = 1;
    104: op1_07_inv23 = 1;
    105: op1_07_inv23 = 1;
    106: op1_07_inv23 = 1;
    109: op1_07_inv23 = 1;
    111: op1_07_inv23 = 1;
    112: op1_07_inv23 = 1;
    113: op1_07_inv23 = 1;
    115: op1_07_inv23 = 1;
    116: op1_07_inv23 = 1;
    117: op1_07_inv23 = 1;
    118: op1_07_inv23 = 1;
    119: op1_07_inv23 = 1;
    42: op1_07_inv23 = 1;
    120: op1_07_inv23 = 1;
    121: op1_07_inv23 = 1;
    122: op1_07_inv23 = 1;
    123: op1_07_inv23 = 1;
    124: op1_07_inv23 = 1;
    125: op1_07_inv23 = 1;
    126: op1_07_inv23 = 1;
    128: op1_07_inv23 = 1;
    130: op1_07_inv23 = 1;
    default: op1_07_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in24 = reg_0439;
    53: op1_07_in24 = reg_0310;
    55: op1_07_in24 = reg_0993;
    86: op1_07_in24 = reg_1139;
    69: op1_07_in24 = reg_0862;
    73: op1_07_in24 = reg_1468;
    50: op1_07_in24 = reg_0550;
    54: op1_07_in24 = reg_0475;
    71: op1_07_in24 = reg_0365;
    74: op1_07_in24 = reg_0269;
    68: op1_07_in24 = reg_0097;
    75: op1_07_in24 = reg_0034;
    61: op1_07_in24 = reg_0283;
    56: op1_07_in24 = reg_0160;
    87: op1_07_in24 = reg_1168;
    76: op1_07_in24 = reg_1351;
    57: op1_07_in24 = reg_0106;
    77: op1_07_in24 = reg_0014;
    60: op1_07_in24 = reg_0719;
    78: op1_07_in24 = reg_0449;
    70: op1_07_in24 = reg_0908;
    46: op1_07_in24 = reg_0377;
    88: op1_07_in24 = reg_0426;
    79: op1_07_in24 = reg_0869;
    48: op1_07_in24 = reg_0977;
    80: op1_07_in24 = reg_0366;
    62: op1_07_in24 = reg_0229;
    52: op1_07_in24 = imem07_in[11:8];
    81: op1_07_in24 = reg_0461;
    63: op1_07_in24 = reg_0974;
    82: op1_07_in24 = reg_1518;
    89: op1_07_in24 = reg_1200;
    83: op1_07_in24 = reg_0715;
    64: op1_07_in24 = reg_0305;
    84: op1_07_in24 = reg_0582;
    85: op1_07_in24 = imem06_in[7:4];
    90: op1_07_in24 = reg_0368;
    66: op1_07_in24 = reg_0609;
    91: op1_07_in24 = reg_1009;
    67: op1_07_in24 = reg_0591;
    92: op1_07_in24 = reg_1488;
    93: op1_07_in24 = reg_0741;
    94: op1_07_in24 = reg_0522;
    95: op1_07_in24 = reg_0008;
    44: op1_07_in24 = imem05_in[11:8];
    96: op1_07_in24 = reg_0526;
    97: op1_07_in24 = reg_0132;
    98: op1_07_in24 = reg_0712;
    99: op1_07_in24 = reg_0507;
    100: op1_07_in24 = reg_0835;
    101: op1_07_in24 = reg_0454;
    103: op1_07_in24 = reg_0966;
    104: op1_07_in24 = reg_0327;
    105: op1_07_in24 = reg_0901;
    106: op1_07_in24 = reg_0589;
    107: op1_07_in24 = reg_0957;
    108: op1_07_in24 = reg_0242;
    109: op1_07_in24 = reg_0548;
    110: op1_07_in24 = reg_0037;
    111: op1_07_in24 = reg_0434;
    112: op1_07_in24 = reg_0500;
    113: op1_07_in24 = reg_0547;
    114: op1_07_in24 = reg_0786;
    115: op1_07_in24 = reg_1091;
    116: op1_07_in24 = reg_0650;
    117: op1_07_in24 = reg_0312;
    118: op1_07_in24 = reg_0021;
    119: op1_07_in24 = reg_0264;
    42: op1_07_in24 = reg_0605;
    120: op1_07_in24 = reg_1433;
    121: op1_07_in24 = reg_0226;
    122: op1_07_in24 = reg_0775;
    123: op1_07_in24 = reg_1474;
    124: op1_07_in24 = reg_0664;
    125: op1_07_in24 = reg_0466;
    126: op1_07_in24 = imem07_in[15:12];
    127: op1_07_in24 = reg_0206;
    128: op1_07_in24 = reg_0342;
    129: op1_07_in24 = reg_0401;
    130: op1_07_in24 = reg_1372;
    default: op1_07_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv24 = 1;
    53: op1_07_inv24 = 1;
    55: op1_07_inv24 = 1;
    69: op1_07_inv24 = 1;
    73: op1_07_inv24 = 1;
    50: op1_07_inv24 = 1;
    54: op1_07_inv24 = 1;
    75: op1_07_inv24 = 1;
    61: op1_07_inv24 = 1;
    76: op1_07_inv24 = 1;
    77: op1_07_inv24 = 1;
    60: op1_07_inv24 = 1;
    78: op1_07_inv24 = 1;
    70: op1_07_inv24 = 1;
    79: op1_07_inv24 = 1;
    80: op1_07_inv24 = 1;
    52: op1_07_inv24 = 1;
    83: op1_07_inv24 = 1;
    84: op1_07_inv24 = 1;
    85: op1_07_inv24 = 1;
    66: op1_07_inv24 = 1;
    92: op1_07_inv24 = 1;
    97: op1_07_inv24 = 1;
    98: op1_07_inv24 = 1;
    100: op1_07_inv24 = 1;
    101: op1_07_inv24 = 1;
    103: op1_07_inv24 = 1;
    105: op1_07_inv24 = 1;
    107: op1_07_inv24 = 1;
    110: op1_07_inv24 = 1;
    114: op1_07_inv24 = 1;
    115: op1_07_inv24 = 1;
    116: op1_07_inv24 = 1;
    117: op1_07_inv24 = 1;
    118: op1_07_inv24 = 1;
    119: op1_07_inv24 = 1;
    42: op1_07_inv24 = 1;
    120: op1_07_inv24 = 1;
    122: op1_07_inv24 = 1;
    123: op1_07_inv24 = 1;
    125: op1_07_inv24 = 1;
    129: op1_07_inv24 = 1;
    default: op1_07_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in25 = reg_0875;
    53: op1_07_in25 = reg_0156;
    55: op1_07_in25 = imem07_in[15:12];
    52: op1_07_in25 = imem07_in[15:12];
    86: op1_07_in25 = reg_0425;
    69: op1_07_in25 = reg_0836;
    73: op1_07_in25 = reg_1064;
    50: op1_07_in25 = reg_0258;
    54: op1_07_in25 = reg_0326;
    71: op1_07_in25 = reg_0899;
    74: op1_07_in25 = reg_0868;
    68: op1_07_in25 = reg_0095;
    75: op1_07_in25 = reg_0672;
    61: op1_07_in25 = reg_0041;
    56: op1_07_in25 = reg_1070;
    87: op1_07_in25 = reg_1169;
    76: op1_07_in25 = reg_0674;
    57: op1_07_in25 = reg_0379;
    77: op1_07_in25 = reg_1334;
    60: op1_07_in25 = reg_0181;
    78: op1_07_in25 = reg_0861;
    70: op1_07_in25 = reg_0905;
    46: op1_07_in25 = reg_0235;
    88: op1_07_in25 = reg_0411;
    79: op1_07_in25 = reg_0752;
    48: op1_07_in25 = reg_0906;
    80: op1_07_in25 = reg_0739;
    62: op1_07_in25 = reg_0998;
    81: op1_07_in25 = reg_1415;
    63: op1_07_in25 = reg_0753;
    127: op1_07_in25 = reg_0753;
    82: op1_07_in25 = reg_1314;
    89: op1_07_in25 = reg_1215;
    83: op1_07_in25 = reg_0967;
    64: op1_07_in25 = reg_0719;
    84: op1_07_in25 = reg_0368;
    85: op1_07_in25 = reg_1501;
    90: op1_07_in25 = reg_0338;
    100: op1_07_in25 = reg_0338;
    66: op1_07_in25 = reg_0982;
    91: op1_07_in25 = reg_0291;
    67: op1_07_in25 = reg_0137;
    92: op1_07_in25 = reg_0470;
    93: op1_07_in25 = reg_0051;
    94: op1_07_in25 = reg_0583;
    97: op1_07_in25 = reg_0583;
    95: op1_07_in25 = reg_1091;
    44: op1_07_in25 = reg_0896;
    96: op1_07_in25 = reg_0529;
    98: op1_07_in25 = reg_0495;
    99: op1_07_in25 = reg_0699;
    101: op1_07_in25 = reg_0062;
    103: op1_07_in25 = reg_1452;
    104: op1_07_in25 = reg_0024;
    105: op1_07_in25 = reg_0078;
    106: op1_07_in25 = reg_0784;
    107: op1_07_in25 = reg_0220;
    108: op1_07_in25 = reg_0241;
    109: op1_07_in25 = reg_0787;
    110: op1_07_in25 = reg_0372;
    111: op1_07_in25 = reg_1457;
    112: op1_07_in25 = reg_1041;
    113: op1_07_in25 = reg_0747;
    114: op1_07_in25 = reg_1349;
    115: op1_07_in25 = reg_0279;
    116: op1_07_in25 = reg_0700;
    117: op1_07_in25 = reg_0191;
    118: op1_07_in25 = reg_0793;
    119: op1_07_in25 = reg_0797;
    42: op1_07_in25 = reg_0590;
    120: op1_07_in25 = reg_1140;
    122: op1_07_in25 = reg_0663;
    123: op1_07_in25 = reg_0468;
    124: op1_07_in25 = reg_0413;
    125: op1_07_in25 = reg_0332;
    126: op1_07_in25 = reg_0087;
    128: op1_07_in25 = reg_1419;
    129: op1_07_in25 = reg_0550;
    130: op1_07_in25 = imem04_in[3:0];
    default: op1_07_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_07_inv25 = 1;
    54: op1_07_inv25 = 1;
    71: op1_07_inv25 = 1;
    76: op1_07_inv25 = 1;
    57: op1_07_inv25 = 1;
    77: op1_07_inv25 = 1;
    60: op1_07_inv25 = 1;
    46: op1_07_inv25 = 1;
    88: op1_07_inv25 = 1;
    79: op1_07_inv25 = 1;
    80: op1_07_inv25 = 1;
    62: op1_07_inv25 = 1;
    52: op1_07_inv25 = 1;
    81: op1_07_inv25 = 1;
    82: op1_07_inv25 = 1;
    85: op1_07_inv25 = 1;
    90: op1_07_inv25 = 1;
    91: op1_07_inv25 = 1;
    92: op1_07_inv25 = 1;
    93: op1_07_inv25 = 1;
    94: op1_07_inv25 = 1;
    95: op1_07_inv25 = 1;
    44: op1_07_inv25 = 1;
    97: op1_07_inv25 = 1;
    99: op1_07_inv25 = 1;
    101: op1_07_inv25 = 1;
    103: op1_07_inv25 = 1;
    104: op1_07_inv25 = 1;
    106: op1_07_inv25 = 1;
    108: op1_07_inv25 = 1;
    109: op1_07_inv25 = 1;
    111: op1_07_inv25 = 1;
    114: op1_07_inv25 = 1;
    115: op1_07_inv25 = 1;
    117: op1_07_inv25 = 1;
    119: op1_07_inv25 = 1;
    42: op1_07_inv25 = 1;
    120: op1_07_inv25 = 1;
    122: op1_07_inv25 = 1;
    123: op1_07_inv25 = 1;
    124: op1_07_inv25 = 1;
    127: op1_07_inv25 = 1;
    default: op1_07_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in26 = reg_0744;
    53: op1_07_in26 = reg_0157;
    55: op1_07_in26 = reg_0309;
    86: op1_07_in26 = reg_0247;
    69: op1_07_in26 = reg_0835;
    73: op1_07_in26 = reg_0536;
    50: op1_07_in26 = reg_0242;
    54: op1_07_in26 = reg_0106;
    71: op1_07_in26 = reg_0875;
    74: op1_07_in26 = reg_1439;
    68: op1_07_in26 = reg_0129;
    60: op1_07_in26 = reg_0129;
    75: op1_07_in26 = reg_0997;
    61: op1_07_in26 = reg_0254;
    56: op1_07_in26 = reg_1069;
    87: op1_07_in26 = reg_0391;
    76: op1_07_in26 = reg_0156;
    57: op1_07_in26 = reg_0056;
    77: op1_07_in26 = reg_0720;
    78: op1_07_in26 = reg_0828;
    70: op1_07_in26 = reg_1420;
    46: op1_07_in26 = reg_0232;
    88: op1_07_in26 = reg_0032;
    79: op1_07_in26 = reg_1505;
    48: op1_07_in26 = reg_0730;
    80: op1_07_in26 = reg_0738;
    62: op1_07_in26 = reg_0298;
    52: op1_07_in26 = reg_1094;
    81: op1_07_in26 = reg_0673;
    63: op1_07_in26 = reg_0929;
    82: op1_07_in26 = reg_1231;
    89: op1_07_in26 = reg_0681;
    83: op1_07_in26 = reg_0439;
    64: op1_07_in26 = reg_0095;
    84: op1_07_in26 = reg_0337;
    85: op1_07_in26 = reg_0635;
    90: op1_07_in26 = reg_1237;
    66: op1_07_in26 = reg_0966;
    109: op1_07_in26 = reg_0966;
    91: op1_07_in26 = imem04_in[3:0];
    92: op1_07_in26 = reg_0370;
    93: op1_07_in26 = reg_0002;
    94: op1_07_in26 = reg_1202;
    95: op1_07_in26 = reg_0279;
    44: op1_07_in26 = reg_0888;
    96: op1_07_in26 = reg_0583;
    97: op1_07_in26 = reg_0023;
    98: op1_07_in26 = reg_0776;
    99: op1_07_in26 = reg_0185;
    100: op1_07_in26 = reg_0210;
    101: op1_07_in26 = reg_0487;
    103: op1_07_in26 = reg_0726;
    104: op1_07_in26 = reg_0009;
    105: op1_07_in26 = reg_0724;
    106: op1_07_in26 = reg_0906;
    107: op1_07_in26 = reg_0246;
    108: op1_07_in26 = reg_0798;
    113: op1_07_in26 = reg_0798;
    129: op1_07_in26 = reg_0798;
    110: op1_07_in26 = imem06_in[15:12];
    111: op1_07_in26 = reg_1456;
    123: op1_07_in26 = reg_1456;
    112: op1_07_in26 = reg_0097;
    114: op1_07_in26 = reg_0139;
    115: op1_07_in26 = reg_0255;
    116: op1_07_in26 = reg_0831;
    117: op1_07_in26 = reg_0145;
    118: op1_07_in26 = reg_0347;
    119: op1_07_in26 = reg_0462;
    42: op1_07_in26 = reg_0562;
    120: op1_07_in26 = reg_0628;
    122: op1_07_in26 = reg_0741;
    124: op1_07_in26 = reg_0618;
    125: op1_07_in26 = reg_0890;
    126: op1_07_in26 = reg_0051;
    127: op1_07_in26 = reg_0264;
    128: op1_07_in26 = reg_0063;
    130: op1_07_in26 = imem04_in[15:12];
    default: op1_07_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_07_inv26 = 1;
    69: op1_07_inv26 = 1;
    50: op1_07_inv26 = 1;
    75: op1_07_inv26 = 1;
    61: op1_07_inv26 = 1;
    87: op1_07_inv26 = 1;
    57: op1_07_inv26 = 1;
    77: op1_07_inv26 = 1;
    60: op1_07_inv26 = 1;
    78: op1_07_inv26 = 1;
    70: op1_07_inv26 = 1;
    48: op1_07_inv26 = 1;
    81: op1_07_inv26 = 1;
    82: op1_07_inv26 = 1;
    89: op1_07_inv26 = 1;
    93: op1_07_inv26 = 1;
    94: op1_07_inv26 = 1;
    95: op1_07_inv26 = 1;
    97: op1_07_inv26 = 1;
    100: op1_07_inv26 = 1;
    103: op1_07_inv26 = 1;
    105: op1_07_inv26 = 1;
    108: op1_07_inv26 = 1;
    109: op1_07_inv26 = 1;
    110: op1_07_inv26 = 1;
    111: op1_07_inv26 = 1;
    112: op1_07_inv26 = 1;
    116: op1_07_inv26 = 1;
    42: op1_07_inv26 = 1;
    122: op1_07_inv26 = 1;
    123: op1_07_inv26 = 1;
    125: op1_07_inv26 = 1;
    126: op1_07_inv26 = 1;
    127: op1_07_inv26 = 1;
    default: op1_07_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in27 = reg_0184;
    53: op1_07_in27 = reg_0924;
    76: op1_07_in27 = reg_0924;
    55: op1_07_in27 = reg_0169;
    86: op1_07_in27 = reg_1383;
    69: op1_07_in27 = reg_0337;
    101: op1_07_in27 = reg_0337;
    73: op1_07_in27 = reg_0264;
    50: op1_07_in27 = reg_0742;
    54: op1_07_in27 = reg_0105;
    71: op1_07_in27 = reg_0080;
    74: op1_07_in27 = reg_0391;
    68: op1_07_in27 = reg_0150;
    75: op1_07_in27 = reg_0324;
    61: op1_07_in27 = reg_0532;
    56: op1_07_in27 = reg_1034;
    87: op1_07_in27 = reg_0566;
    57: op1_07_in27 = reg_0390;
    77: op1_07_in27 = reg_0827;
    60: op1_07_in27 = reg_0210;
    78: op1_07_in27 = reg_0206;
    70: op1_07_in27 = reg_0870;
    46: op1_07_in27 = reg_0025;
    88: op1_07_in27 = reg_0263;
    127: op1_07_in27 = reg_0263;
    79: op1_07_in27 = reg_0110;
    48: op1_07_in27 = reg_0825;
    80: op1_07_in27 = reg_0408;
    62: op1_07_in27 = reg_0894;
    52: op1_07_in27 = reg_0673;
    81: op1_07_in27 = reg_0298;
    63: op1_07_in27 = reg_0193;
    82: op1_07_in27 = reg_1093;
    89: op1_07_in27 = reg_1233;
    83: op1_07_in27 = reg_0430;
    64: op1_07_in27 = reg_0117;
    84: op1_07_in27 = reg_0236;
    85: op1_07_in27 = reg_0115;
    90: op1_07_in27 = reg_0211;
    66: op1_07_in27 = reg_0438;
    91: op1_07_in27 = imem04_in[11:8];
    92: op1_07_in27 = reg_0579;
    93: op1_07_in27 = reg_0052;
    94: op1_07_in27 = reg_0371;
    95: op1_07_in27 = reg_0255;
    44: op1_07_in27 = reg_0873;
    96: op1_07_in27 = reg_1202;
    97: op1_07_in27 = imem07_in[7:4];
    98: op1_07_in27 = reg_0326;
    99: op1_07_in27 = reg_0154;
    100: op1_07_in27 = reg_0470;
    103: op1_07_in27 = reg_0386;
    104: op1_07_in27 = reg_0279;
    105: op1_07_in27 = reg_0634;
    106: op1_07_in27 = reg_0859;
    107: op1_07_in27 = reg_0558;
    108: op1_07_in27 = reg_0966;
    109: op1_07_in27 = reg_0967;
    110: op1_07_in27 = reg_0906;
    111: op1_07_in27 = reg_0147;
    123: op1_07_in27 = reg_0147;
    112: op1_07_in27 = reg_0369;
    113: op1_07_in27 = reg_1474;
    129: op1_07_in27 = reg_1474;
    114: op1_07_in27 = reg_0031;
    115: op1_07_in27 = reg_0006;
    116: op1_07_in27 = reg_0066;
    117: op1_07_in27 = reg_0000;
    118: op1_07_in27 = reg_1164;
    119: op1_07_in27 = reg_0531;
    42: op1_07_in27 = reg_0560;
    120: op1_07_in27 = reg_0745;
    122: op1_07_in27 = reg_0413;
    124: op1_07_in27 = reg_0591;
    125: op1_07_in27 = reg_0445;
    126: op1_07_in27 = reg_0851;
    128: op1_07_in27 = reg_0035;
    130: op1_07_in27 = reg_0936;
    default: op1_07_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_07_inv27 = 1;
    69: op1_07_inv27 = 1;
    73: op1_07_inv27 = 1;
    74: op1_07_inv27 = 1;
    75: op1_07_inv27 = 1;
    56: op1_07_inv27 = 1;
    57: op1_07_inv27 = 1;
    70: op1_07_inv27 = 1;
    46: op1_07_inv27 = 1;
    88: op1_07_inv27 = 1;
    79: op1_07_inv27 = 1;
    62: op1_07_inv27 = 1;
    52: op1_07_inv27 = 1;
    81: op1_07_inv27 = 1;
    84: op1_07_inv27 = 1;
    85: op1_07_inv27 = 1;
    90: op1_07_inv27 = 1;
    91: op1_07_inv27 = 1;
    92: op1_07_inv27 = 1;
    93: op1_07_inv27 = 1;
    94: op1_07_inv27 = 1;
    44: op1_07_inv27 = 1;
    96: op1_07_inv27 = 1;
    98: op1_07_inv27 = 1;
    103: op1_07_inv27 = 1;
    104: op1_07_inv27 = 1;
    105: op1_07_inv27 = 1;
    107: op1_07_inv27 = 1;
    108: op1_07_inv27 = 1;
    109: op1_07_inv27 = 1;
    113: op1_07_inv27 = 1;
    114: op1_07_inv27 = 1;
    118: op1_07_inv27 = 1;
    42: op1_07_inv27 = 1;
    120: op1_07_inv27 = 1;
    124: op1_07_inv27 = 1;
    125: op1_07_inv27 = 1;
    126: op1_07_inv27 = 1;
    127: op1_07_inv27 = 1;
    130: op1_07_inv27 = 1;
    default: op1_07_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in28 = reg_0253;
    120: op1_07_in28 = reg_0253;
    53: op1_07_in28 = reg_0777;
    55: op1_07_in28 = reg_0777;
    86: op1_07_in28 = reg_1372;
    69: op1_07_in28 = reg_0338;
    73: op1_07_in28 = imem06_in[11:8];
    50: op1_07_in28 = reg_0984;
    54: op1_07_in28 = reg_0380;
    71: op1_07_in28 = reg_0078;
    74: op1_07_in28 = reg_1440;
    68: op1_07_in28 = reg_0792;
    75: op1_07_in28 = reg_1414;
    61: op1_07_in28 = reg_0455;
    56: op1_07_in28 = imem01_in[3:0];
    87: op1_07_in28 = reg_0167;
    76: op1_07_in28 = reg_0139;
    57: op1_07_in28 = reg_0294;
    77: op1_07_in28 = reg_0161;
    60: op1_07_in28 = reg_0209;
    84: op1_07_in28 = reg_0209;
    78: op1_07_in28 = imem06_in[7:4];
    70: op1_07_in28 = reg_0264;
    46: op1_07_in28 = reg_0790;
    88: op1_07_in28 = reg_0493;
    79: op1_07_in28 = reg_0718;
    48: op1_07_in28 = reg_0109;
    80: op1_07_in28 = reg_0623;
    62: op1_07_in28 = reg_0225;
    52: op1_07_in28 = reg_0157;
    81: op1_07_in28 = reg_0667;
    63: op1_07_in28 = reg_0696;
    82: op1_07_in28 = reg_1208;
    89: op1_07_in28 = reg_0500;
    83: op1_07_in28 = reg_0434;
    64: op1_07_in28 = reg_0061;
    85: op1_07_in28 = reg_0194;
    90: op1_07_in28 = reg_0236;
    66: op1_07_in28 = reg_0930;
    91: op1_07_in28 = reg_1369;
    92: op1_07_in28 = reg_0735;
    93: op1_07_in28 = reg_0518;
    94: op1_07_in28 = reg_1179;
    96: op1_07_in28 = reg_1179;
    95: op1_07_in28 = reg_0632;
    104: op1_07_in28 = reg_0632;
    44: op1_07_in28 = reg_0196;
    97: op1_07_in28 = imem07_in[11:8];
    98: op1_07_in28 = reg_0971;
    99: op1_07_in28 = reg_1063;
    100: op1_07_in28 = imem05_in[3:0];
    101: op1_07_in28 = reg_0035;
    103: op1_07_in28 = reg_0091;
    105: op1_07_in28 = imem01_in[11:8];
    106: op1_07_in28 = reg_0827;
    107: op1_07_in28 = reg_1149;
    108: op1_07_in28 = reg_0968;
    109: op1_07_in28 = reg_0726;
    110: op1_07_in28 = reg_0192;
    111: op1_07_in28 = reg_0899;
    112: op1_07_in28 = reg_0835;
    113: op1_07_in28 = reg_0715;
    114: op1_07_in28 = reg_0413;
    115: op1_07_in28 = reg_0328;
    116: op1_07_in28 = reg_0491;
    117: op1_07_in28 = reg_0891;
    118: op1_07_in28 = reg_0649;
    119: op1_07_in28 = reg_0552;
    42: op1_07_in28 = reg_0530;
    122: op1_07_in28 = reg_0621;
    123: op1_07_in28 = reg_0146;
    124: op1_07_in28 = reg_0520;
    125: op1_07_in28 = reg_0733;
    126: op1_07_in28 = reg_0159;
    127: op1_07_in28 = reg_0960;
    128: op1_07_in28 = reg_0832;
    129: op1_07_in28 = reg_0572;
    130: op1_07_in28 = reg_0034;
    default: op1_07_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_07_inv28 = 1;
    73: op1_07_inv28 = 1;
    54: op1_07_inv28 = 1;
    74: op1_07_inv28 = 1;
    75: op1_07_inv28 = 1;
    87: op1_07_inv28 = 1;
    77: op1_07_inv28 = 1;
    78: op1_07_inv28 = 1;
    70: op1_07_inv28 = 1;
    88: op1_07_inv28 = 1;
    79: op1_07_inv28 = 1;
    48: op1_07_inv28 = 1;
    80: op1_07_inv28 = 1;
    63: op1_07_inv28 = 1;
    89: op1_07_inv28 = 1;
    84: op1_07_inv28 = 1;
    85: op1_07_inv28 = 1;
    90: op1_07_inv28 = 1;
    91: op1_07_inv28 = 1;
    93: op1_07_inv28 = 1;
    94: op1_07_inv28 = 1;
    95: op1_07_inv28 = 1;
    96: op1_07_inv28 = 1;
    99: op1_07_inv28 = 1;
    100: op1_07_inv28 = 1;
    101: op1_07_inv28 = 1;
    104: op1_07_inv28 = 1;
    107: op1_07_inv28 = 1;
    109: op1_07_inv28 = 1;
    111: op1_07_inv28 = 1;
    112: op1_07_inv28 = 1;
    113: op1_07_inv28 = 1;
    115: op1_07_inv28 = 1;
    117: op1_07_inv28 = 1;
    118: op1_07_inv28 = 1;
    119: op1_07_inv28 = 1;
    120: op1_07_inv28 = 1;
    122: op1_07_inv28 = 1;
    124: op1_07_inv28 = 1;
    125: op1_07_inv28 = 1;
    127: op1_07_inv28 = 1;
    128: op1_07_inv28 = 1;
    129: op1_07_inv28 = 1;
    130: op1_07_inv28 = 1;
    default: op1_07_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in29 = reg_1018;
    53: op1_07_in29 = reg_0779;
    55: op1_07_in29 = reg_0030;
    86: op1_07_in29 = imem04_in[3:0];
    69: op1_07_in29 = reg_0237;
    73: op1_07_in29 = reg_0373;
    50: op1_07_in29 = reg_0468;
    54: op1_07_in29 = reg_0898;
    71: op1_07_in29 = reg_0290;
    74: op1_07_in29 = reg_0162;
    68: op1_07_in29 = reg_0794;
    116: op1_07_in29 = reg_0794;
    75: op1_07_in29 = reg_1415;
    61: op1_07_in29 = reg_0588;
    56: op1_07_in29 = reg_0930;
    87: op1_07_in29 = reg_1514;
    76: op1_07_in29 = reg_1094;
    57: op1_07_in29 = reg_0878;
    77: op1_07_in29 = reg_0116;
    60: op1_07_in29 = reg_0021;
    78: op1_07_in29 = reg_0755;
    70: op1_07_in29 = reg_0109;
    46: op1_07_in29 = reg_0180;
    88: op1_07_in29 = reg_0088;
    91: op1_07_in29 = reg_0088;
    79: op1_07_in29 = reg_0637;
    48: op1_07_in29 = reg_0636;
    106: op1_07_in29 = reg_0636;
    80: op1_07_in29 = reg_0053;
    62: op1_07_in29 = reg_0309;
    52: op1_07_in29 = reg_0489;
    81: op1_07_in29 = reg_0892;
    63: op1_07_in29 = imem06_in[15:12];
    82: op1_07_in29 = reg_0113;
    89: op1_07_in29 = reg_0412;
    83: op1_07_in29 = reg_0400;
    64: op1_07_in29 = reg_0019;
    84: op1_07_in29 = reg_0065;
    85: op1_07_in29 = reg_0141;
    90: op1_07_in29 = reg_0932;
    66: op1_07_in29 = reg_0147;
    129: op1_07_in29 = reg_0147;
    92: op1_07_in29 = reg_0578;
    93: op1_07_in29 = reg_0484;
    94: op1_07_in29 = reg_0213;
    95: op1_07_in29 = imem03_in[3:0];
    44: op1_07_in29 = reg_0118;
    96: op1_07_in29 = reg_0270;
    97: op1_07_in29 = imem07_in[15:12];
    98: op1_07_in29 = reg_0125;
    99: op1_07_in29 = reg_0191;
    100: op1_07_in29 = imem05_in[15:12];
    101: op1_07_in29 = imem05_in[15:12];
    103: op1_07_in29 = reg_0901;
    104: op1_07_in29 = reg_0377;
    105: op1_07_in29 = reg_0456;
    107: op1_07_in29 = reg_1009;
    108: op1_07_in29 = reg_0819;
    109: op1_07_in29 = reg_0146;
    110: op1_07_in29 = reg_0316;
    127: op1_07_in29 = reg_0316;
    111: op1_07_in29 = reg_0595;
    112: op1_07_in29 = reg_1237;
    113: op1_07_in29 = reg_0572;
    114: op1_07_in29 = reg_0103;
    115: op1_07_in29 = reg_0999;
    117: op1_07_in29 = reg_0070;
    118: op1_07_in29 = reg_0604;
    119: op1_07_in29 = reg_1198;
    42: op1_07_in29 = reg_0495;
    120: op1_07_in29 = reg_0903;
    122: op1_07_in29 = reg_0620;
    123: op1_07_in29 = reg_1253;
    125: op1_07_in29 = reg_0176;
    126: op1_07_in29 = reg_0158;
    128: op1_07_in29 = reg_0040;
    130: op1_07_in29 = reg_0236;
    default: op1_07_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv29 = 1;
    53: op1_07_inv29 = 1;
    73: op1_07_inv29 = 1;
    75: op1_07_inv29 = 1;
    61: op1_07_inv29 = 1;
    76: op1_07_inv29 = 1;
    57: op1_07_inv29 = 1;
    77: op1_07_inv29 = 1;
    79: op1_07_inv29 = 1;
    62: op1_07_inv29 = 1;
    52: op1_07_inv29 = 1;
    63: op1_07_inv29 = 1;
    82: op1_07_inv29 = 1;
    89: op1_07_inv29 = 1;
    83: op1_07_inv29 = 1;
    66: op1_07_inv29 = 1;
    92: op1_07_inv29 = 1;
    94: op1_07_inv29 = 1;
    97: op1_07_inv29 = 1;
    98: op1_07_inv29 = 1;
    99: op1_07_inv29 = 1;
    100: op1_07_inv29 = 1;
    101: op1_07_inv29 = 1;
    107: op1_07_inv29 = 1;
    108: op1_07_inv29 = 1;
    109: op1_07_inv29 = 1;
    111: op1_07_inv29 = 1;
    114: op1_07_inv29 = 1;
    117: op1_07_inv29 = 1;
    118: op1_07_inv29 = 1;
    119: op1_07_inv29 = 1;
    42: op1_07_inv29 = 1;
    122: op1_07_inv29 = 1;
    125: op1_07_inv29 = 1;
    126: op1_07_inv29 = 1;
    128: op1_07_inv29 = 1;
    default: op1_07_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_07_in30 = imem02_in[15:12];
    53: op1_07_in30 = reg_0031;
    55: op1_07_in30 = reg_0661;
    86: op1_07_in30 = imem04_in[11:8];
    69: op1_07_in30 = reg_0117;
    73: op1_07_in30 = reg_0570;
    50: op1_07_in30 = reg_0967;
    54: op1_07_in30 = reg_0878;
    71: op1_07_in30 = reg_0222;
    74: op1_07_in30 = reg_0025;
    68: op1_07_in30 = reg_0579;
    64: op1_07_in30 = reg_0579;
    75: op1_07_in30 = reg_1315;
    61: op1_07_in30 = reg_0560;
    56: op1_07_in30 = reg_0291;
    107: op1_07_in30 = reg_0291;
    87: op1_07_in30 = reg_0303;
    76: op1_07_in30 = reg_0285;
    57: op1_07_in30 = reg_0877;
    77: op1_07_in30 = reg_0109;
    60: op1_07_in30 = reg_0020;
    78: op1_07_in30 = reg_1509;
    70: op1_07_in30 = reg_0717;
    46: op1_07_in30 = reg_0178;
    88: op1_07_in30 = reg_0264;
    91: op1_07_in30 = reg_0264;
    79: op1_07_in30 = reg_0398;
    48: op1_07_in30 = reg_0637;
    106: op1_07_in30 = reg_0637;
    80: op1_07_in30 = reg_0084;
    62: op1_07_in30 = reg_0674;
    52: op1_07_in30 = reg_0139;
    81: op1_07_in30 = reg_1351;
    63: op1_07_in30 = reg_0859;
    82: op1_07_in30 = reg_0885;
    89: op1_07_in30 = reg_0097;
    83: op1_07_in30 = reg_0403;
    84: op1_07_in30 = reg_0708;
    85: op1_07_in30 = reg_0617;
    90: op1_07_in30 = reg_0095;
    66: op1_07_in30 = reg_0149;
    92: op1_07_in30 = reg_1431;
    94: op1_07_in30 = reg_0018;
    95: op1_07_in30 = reg_0699;
    44: op1_07_in30 = reg_0240;
    96: op1_07_in30 = reg_0213;
    97: op1_07_in30 = reg_0867;
    98: op1_07_in30 = reg_0111;
    99: op1_07_in30 = reg_0234;
    100: op1_07_in30 = reg_0833;
    101: op1_07_in30 = reg_1059;
    103: op1_07_in30 = reg_0595;
    104: op1_07_in30 = reg_0328;
    130: op1_07_in30 = reg_0328;
    105: op1_07_in30 = reg_0626;
    108: op1_07_in30 = reg_0430;
    109: op1_07_in30 = reg_0290;
    110: op1_07_in30 = reg_1323;
    111: op1_07_in30 = reg_0079;
    112: op1_07_in30 = reg_0236;
    113: op1_07_in30 = reg_0966;
    114: op1_07_in30 = reg_0114;
    115: op1_07_in30 = reg_0750;
    116: op1_07_in30 = reg_0492;
    117: op1_07_in30 = reg_0349;
    118: op1_07_in30 = reg_0045;
    119: op1_07_in30 = reg_0421;
    42: op1_07_in30 = reg_0474;
    120: op1_07_in30 = reg_0824;
    122: op1_07_in30 = reg_0593;
    123: op1_07_in30 = reg_1034;
    125: op1_07_in30 = reg_0793;
    126: op1_07_in30 = reg_0923;
    127: op1_07_in30 = reg_1179;
    128: op1_07_in30 = reg_1164;
    129: op1_07_in30 = reg_1032;
    default: op1_07_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_07_inv30 = 1;
    55: op1_07_inv30 = 1;
    54: op1_07_inv30 = 1;
    75: op1_07_inv30 = 1;
    56: op1_07_inv30 = 1;
    87: op1_07_inv30 = 1;
    57: op1_07_inv30 = 1;
    77: op1_07_inv30 = 1;
    60: op1_07_inv30 = 1;
    78: op1_07_inv30 = 1;
    46: op1_07_inv30 = 1;
    48: op1_07_inv30 = 1;
    62: op1_07_inv30 = 1;
    52: op1_07_inv30 = 1;
    81: op1_07_inv30 = 1;
    84: op1_07_inv30 = 1;
    85: op1_07_inv30 = 1;
    90: op1_07_inv30 = 1;
    92: op1_07_inv30 = 1;
    44: op1_07_inv30 = 1;
    96: op1_07_inv30 = 1;
    97: op1_07_inv30 = 1;
    101: op1_07_inv30 = 1;
    103: op1_07_inv30 = 1;
    104: op1_07_inv30 = 1;
    106: op1_07_inv30 = 1;
    107: op1_07_inv30 = 1;
    109: op1_07_inv30 = 1;
    111: op1_07_inv30 = 1;
    112: op1_07_inv30 = 1;
    113: op1_07_inv30 = 1;
    114: op1_07_inv30 = 1;
    129: op1_07_inv30 = 1;
    default: op1_07_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_07_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#7の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_07_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in00 = imem05_in[7:4];
    53: op1_08_in00 = imem01_in[3:0];
    55: op1_08_in00 = reg_0527;
    86: op1_08_in00 = imem03_in[7:4];
    40: op1_08_in00 = imem03_in[7:4];
    73: op1_08_in00 = reg_0196;
    116: op1_08_in00 = reg_0196;
    69: op1_08_in00 = reg_0365;
    109: op1_08_in00 = reg_0365;
    49: op1_08_in00 = imem07_in[11:8];
    94: op1_08_in00 = imem07_in[11:8];
    50: op1_08_in00 = reg_0386;
    54: op1_08_in00 = reg_0166;
    74: op1_08_in00 = reg_0219;
    62: op1_08_in00 = reg_0219;
    68: op1_08_in00 = reg_0329;
    71: op1_08_in00 = reg_0554;
    75: op1_08_in00 = reg_0580;
    61: op1_08_in00 = reg_1277;
    56: op1_08_in00 = reg_0291;
    87: op1_08_in00 = reg_0711;
    76: op1_08_in00 = imem00_in[11:8];
    83: op1_08_in00 = imem00_in[11:8];
    57: op1_08_in00 = reg_0295;
    77: op1_08_in00 = reg_0983;
    58: op1_08_in00 = reg_0238;
    78: op1_08_in00 = reg_0397;
    70: op1_08_in00 = reg_0473;
    51: op1_08_in00 = reg_0271;
    88: op1_08_in00 = reg_0314;
    46: op1_08_in00 = reg_0532;
    59: op1_08_in00 = imem03_in[15:12];
    79: op1_08_in00 = reg_0418;
    60: op1_08_in00 = reg_0330;
    80: op1_08_in00 = reg_0616;
    33: op1_08_in00 = reg_0158;
    48: op1_08_in00 = reg_0369;
    52: op1_08_in00 = reg_0646;
    81: op1_08_in00 = imem00_in[3:0];
    63: op1_08_in00 = reg_1313;
    82: op1_08_in00 = imem05_in[3:0];
    89: op1_08_in00 = reg_0190;
    28: op1_08_in00 = reg_0028;
    64: op1_08_in00 = reg_0578;
    84: op1_08_in00 = reg_1299;
    65: op1_08_in00 = reg_0967;
    85: op1_08_in00 = reg_0350;
    90: op1_08_in00 = reg_1503;
    37: op1_08_in00 = imem07_in[3:0];
    66: op1_08_in00 = reg_0383;
    91: op1_08_in00 = reg_0034;
    67: op1_08_in00 = reg_1280;
    92: op1_08_in00 = reg_0562;
    93: op1_08_in00 = reg_1470;
    95: op1_08_in00 = reg_0710;
    96: op1_08_in00 = reg_0022;
    97: op1_08_in00 = reg_0498;
    98: op1_08_in00 = reg_0106;
    99: op1_08_in00 = reg_0965;
    44: op1_08_in00 = reg_0346;
    100: op1_08_in00 = reg_0791;
    114: op1_08_in00 = reg_0791;
    47: op1_08_in00 = reg_0735;
    101: op1_08_in00 = reg_1430;
    102: op1_08_in00 = reg_0866;
    103: op1_08_in00 = reg_0400;
    104: op1_08_in00 = reg_0732;
    105: op1_08_in00 = reg_0056;
    106: op1_08_in00 = reg_0569;
    107: op1_08_in00 = reg_0864;
    108: op1_08_in00 = reg_1457;
    110: op1_08_in00 = reg_1504;
    111: op1_08_in00 = reg_0634;
    112: op1_08_in00 = reg_0064;
    113: op1_08_in00 = reg_0819;
    115: op1_08_in00 = reg_0246;
    117: op1_08_in00 = reg_1314;
    118: op1_08_in00 = reg_0051;
    119: op1_08_in00 = reg_1104;
    34: op1_08_in00 = reg_0156;
    120: op1_08_in00 = reg_1078;
    121: op1_08_in00 = reg_0725;
    122: op1_08_in00 = reg_0248;
    123: op1_08_in00 = reg_0360;
    124: op1_08_in00 = reg_0581;
    125: op1_08_in00 = reg_0391;
    126: op1_08_in00 = reg_0843;
    38: op1_08_in00 = reg_0442;
    127: op1_08_in00 = reg_0714;
    42: op1_08_in00 = reg_0363;
    128: op1_08_in00 = reg_0604;
    129: op1_08_in00 = reg_0269;
    22: op1_08_in00 = reg_0102;
    130: op1_08_in00 = reg_0978;
    131: op1_08_in00 = imem00_in[7:4];
    default: op1_08_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv00 = 1;
    53: op1_08_inv00 = 1;
    86: op1_08_inv00 = 1;
    49: op1_08_inv00 = 1;
    54: op1_08_inv00 = 1;
    74: op1_08_inv00 = 1;
    71: op1_08_inv00 = 1;
    87: op1_08_inv00 = 1;
    57: op1_08_inv00 = 1;
    78: op1_08_inv00 = 1;
    88: op1_08_inv00 = 1;
    46: op1_08_inv00 = 1;
    60: op1_08_inv00 = 1;
    80: op1_08_inv00 = 1;
    33: op1_08_inv00 = 1;
    62: op1_08_inv00 = 1;
    82: op1_08_inv00 = 1;
    28: op1_08_inv00 = 1;
    64: op1_08_inv00 = 1;
    65: op1_08_inv00 = 1;
    85: op1_08_inv00 = 1;
    90: op1_08_inv00 = 1;
    37: op1_08_inv00 = 1;
    66: op1_08_inv00 = 1;
    92: op1_08_inv00 = 1;
    94: op1_08_inv00 = 1;
    95: op1_08_inv00 = 1;
    96: op1_08_inv00 = 1;
    97: op1_08_inv00 = 1;
    100: op1_08_inv00 = 1;
    47: op1_08_inv00 = 1;
    40: op1_08_inv00 = 1;
    102: op1_08_inv00 = 1;
    103: op1_08_inv00 = 1;
    105: op1_08_inv00 = 1;
    106: op1_08_inv00 = 1;
    108: op1_08_inv00 = 1;
    112: op1_08_inv00 = 1;
    116: op1_08_inv00 = 1;
    119: op1_08_inv00 = 1;
    125: op1_08_inv00 = 1;
    126: op1_08_inv00 = 1;
    129: op1_08_inv00 = 1;
    22: op1_08_inv00 = 1;
    130: op1_08_inv00 = 1;
    131: op1_08_inv00 = 1;
    default: op1_08_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in01 = reg_0864;
    53: op1_08_in01 = imem01_in[15:12];
    55: op1_08_in01 = reg_0171;
    86: op1_08_in01 = reg_0348;
    67: op1_08_in01 = reg_0348;
    73: op1_08_in01 = reg_0118;
    69: op1_08_in01 = reg_0901;
    49: op1_08_in01 = reg_0623;
    50: op1_08_in01 = reg_0362;
    66: op1_08_in01 = reg_0362;
    108: op1_08_in01 = reg_0362;
    54: op1_08_in01 = reg_0259;
    74: op1_08_in01 = reg_0616;
    62: op1_08_in01 = reg_0616;
    68: op1_08_in01 = reg_0178;
    71: op1_08_in01 = reg_0615;
    75: op1_08_in01 = imem00_in[7:4];
    61: op1_08_in01 = reg_1243;
    56: op1_08_in01 = reg_0282;
    87: op1_08_in01 = reg_0801;
    76: op1_08_in01 = reg_0613;
    57: op1_08_in01 = reg_0289;
    77: op1_08_in01 = imem00_in[11:8];
    58: op1_08_in01 = reg_0819;
    78: op1_08_in01 = reg_0863;
    70: op1_08_in01 = reg_0474;
    51: op1_08_in01 = reg_0152;
    106: op1_08_in01 = reg_0152;
    88: op1_08_in01 = reg_1313;
    46: op1_08_in01 = reg_0473;
    59: op1_08_in01 = reg_0425;
    79: op1_08_in01 = reg_0872;
    60: op1_08_in01 = reg_1280;
    80: op1_08_in01 = reg_1279;
    121: op1_08_in01 = reg_1279;
    33: op1_08_in01 = reg_0285;
    48: op1_08_in01 = reg_0262;
    52: op1_08_in01 = reg_0648;
    81: op1_08_in01 = reg_0552;
    63: op1_08_in01 = reg_0957;
    117: op1_08_in01 = reg_0957;
    82: op1_08_in01 = imem05_in[7:4];
    89: op1_08_in01 = reg_1300;
    28: op1_08_in01 = reg_0002;
    83: op1_08_in01 = reg_0983;
    102: op1_08_in01 = reg_0983;
    122: op1_08_in01 = reg_0983;
    64: op1_08_in01 = reg_1299;
    84: op1_08_in01 = reg_0251;
    65: op1_08_in01 = reg_0930;
    85: op1_08_in01 = imem00_in[15:12];
    90: op1_08_in01 = reg_0019;
    37: op1_08_in01 = reg_0100;
    91: op1_08_in01 = reg_1198;
    92: op1_08_in01 = reg_0701;
    93: op1_08_in01 = reg_1141;
    94: op1_08_in01 = reg_0868;
    95: op1_08_in01 = reg_0312;
    96: op1_08_in01 = reg_0498;
    97: op1_08_in01 = reg_1010;
    98: op1_08_in01 = reg_0684;
    99: op1_08_in01 = reg_1516;
    44: op1_08_in01 = reg_0174;
    100: op1_08_in01 = reg_1439;
    47: op1_08_in01 = reg_0832;
    101: op1_08_in01 = reg_0833;
    40: op1_08_in01 = reg_0537;
    103: op1_08_in01 = reg_0896;
    104: op1_08_in01 = reg_0261;
    105: op1_08_in01 = reg_0276;
    107: op1_08_in01 = reg_0038;
    109: op1_08_in01 = reg_0899;
    123: op1_08_in01 = reg_0899;
    110: op1_08_in01 = reg_0265;
    111: op1_08_in01 = reg_0043;
    112: op1_08_in01 = reg_1503;
    113: op1_08_in01 = reg_0438;
    114: op1_08_in01 = reg_1490;
    115: op1_08_in01 = reg_0049;
    116: op1_08_in01 = reg_0130;
    118: op1_08_in01 = reg_0394;
    119: op1_08_in01 = reg_0045;
    34: op1_08_in01 = reg_0157;
    120: op1_08_in01 = reg_0227;
    124: op1_08_in01 = imem00_in[3:0];
    125: op1_08_in01 = reg_1104;
    126: op1_08_in01 = reg_1491;
    38: op1_08_in01 = reg_0738;
    127: op1_08_in01 = reg_1302;
    42: op1_08_in01 = reg_0091;
    128: op1_08_in01 = reg_0697;
    129: op1_08_in01 = reg_0363;
    22: op1_08_in01 = reg_0103;
    130: op1_08_in01 = reg_0421;
    131: op1_08_in01 = reg_1242;
    default: op1_08_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv01 = 1;
    55: op1_08_inv01 = 1;
    73: op1_08_inv01 = 1;
    49: op1_08_inv01 = 1;
    54: op1_08_inv01 = 1;
    68: op1_08_inv01 = 1;
    75: op1_08_inv01 = 1;
    61: op1_08_inv01 = 1;
    56: op1_08_inv01 = 1;
    76: op1_08_inv01 = 1;
    58: op1_08_inv01 = 1;
    78: op1_08_inv01 = 1;
    51: op1_08_inv01 = 1;
    88: op1_08_inv01 = 1;
    59: op1_08_inv01 = 1;
    79: op1_08_inv01 = 1;
    48: op1_08_inv01 = 1;
    52: op1_08_inv01 = 1;
    81: op1_08_inv01 = 1;
    82: op1_08_inv01 = 1;
    28: op1_08_inv01 = 1;
    83: op1_08_inv01 = 1;
    90: op1_08_inv01 = 1;
    66: op1_08_inv01 = 1;
    92: op1_08_inv01 = 1;
    93: op1_08_inv01 = 1;
    95: op1_08_inv01 = 1;
    96: op1_08_inv01 = 1;
    97: op1_08_inv01 = 1;
    99: op1_08_inv01 = 1;
    100: op1_08_inv01 = 1;
    47: op1_08_inv01 = 1;
    40: op1_08_inv01 = 1;
    104: op1_08_inv01 = 1;
    106: op1_08_inv01 = 1;
    109: op1_08_inv01 = 1;
    111: op1_08_inv01 = 1;
    114: op1_08_inv01 = 1;
    116: op1_08_inv01 = 1;
    117: op1_08_inv01 = 1;
    119: op1_08_inv01 = 1;
    34: op1_08_inv01 = 1;
    120: op1_08_inv01 = 1;
    124: op1_08_inv01 = 1;
    125: op1_08_inv01 = 1;
    38: op1_08_inv01 = 1;
    127: op1_08_inv01 = 1;
    42: op1_08_inv01 = 1;
    129: op1_08_inv01 = 1;
    default: op1_08_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in02 = reg_0828;
    53: op1_08_in02 = reg_0439;
    55: op1_08_in02 = reg_0419;
    86: op1_08_in02 = reg_0425;
    73: op1_08_in02 = reg_1348;
    69: op1_08_in02 = reg_0078;
    66: op1_08_in02 = reg_0078;
    49: op1_08_in02 = reg_0593;
    50: op1_08_in02 = reg_0360;
    54: op1_08_in02 = reg_0982;
    74: op1_08_in02 = imem00_in[7:4];
    93: op1_08_in02 = imem00_in[7:4];
    68: op1_08_in02 = reg_1208;
    71: op1_08_in02 = reg_0614;
    75: op1_08_in02 = imem00_in[15:12];
    61: op1_08_in02 = reg_1052;
    56: op1_08_in02 = reg_1029;
    87: op1_08_in02 = reg_0217;
    76: op1_08_in02 = reg_0841;
    57: op1_08_in02 = reg_1179;
    77: op1_08_in02 = reg_1079;
    80: op1_08_in02 = reg_1079;
    58: op1_08_in02 = reg_0930;
    78: op1_08_in02 = reg_0669;
    70: op1_08_in02 = reg_0495;
    51: op1_08_in02 = reg_0018;
    88: op1_08_in02 = reg_0954;
    46: op1_08_in02 = reg_0475;
    59: op1_08_in02 = reg_0443;
    79: op1_08_in02 = reg_0601;
    60: op1_08_in02 = reg_0427;
    67: op1_08_in02 = reg_0427;
    33: op1_08_in02 = imem07_in[3:0];
    62: op1_08_in02 = reg_0748;
    48: op1_08_in02 = reg_0129;
    52: op1_08_in02 = reg_0992;
    81: op1_08_in02 = reg_0562;
    63: op1_08_in02 = reg_0220;
    82: op1_08_in02 = reg_0566;
    125: op1_08_in02 = reg_0566;
    89: op1_08_in02 = reg_1301;
    28: op1_08_in02 = imem07_in[7:4];
    83: op1_08_in02 = reg_0868;
    64: op1_08_in02 = reg_0737;
    84: op1_08_in02 = reg_1163;
    65: op1_08_in02 = reg_0384;
    85: op1_08_in02 = reg_0983;
    90: op1_08_in02 = reg_0016;
    37: op1_08_in02 = reg_0001;
    91: op1_08_in02 = reg_1200;
    92: op1_08_in02 = reg_0182;
    94: op1_08_in02 = reg_0135;
    95: op1_08_in02 = reg_0000;
    96: op1_08_in02 = reg_0465;
    97: op1_08_in02 = reg_1440;
    98: op1_08_in02 = reg_0628;
    99: op1_08_in02 = reg_1517;
    44: op1_08_in02 = reg_0602;
    100: op1_08_in02 = reg_0667;
    47: op1_08_in02 = reg_0176;
    101: op1_08_in02 = reg_0733;
    40: op1_08_in02 = reg_0488;
    102: op1_08_in02 = reg_0445;
    103: op1_08_in02 = reg_0634;
    104: op1_08_in02 = reg_1001;
    105: op1_08_in02 = reg_1260;
    106: op1_08_in02 = reg_1010;
    107: op1_08_in02 = reg_0039;
    108: op1_08_in02 = reg_0365;
    109: op1_08_in02 = reg_0901;
    129: op1_08_in02 = reg_0901;
    110: op1_08_in02 = reg_0115;
    111: op1_08_in02 = reg_0895;
    112: op1_08_in02 = reg_0470;
    113: op1_08_in02 = reg_0726;
    114: op1_08_in02 = reg_0803;
    115: op1_08_in02 = reg_0709;
    116: op1_08_in02 = reg_0243;
    117: op1_08_in02 = reg_0952;
    118: op1_08_in02 = reg_0993;
    119: op1_08_in02 = reg_0697;
    34: op1_08_in02 = reg_0286;
    120: op1_08_in02 = imem03_in[11:8];
    121: op1_08_in02 = reg_1489;
    122: op1_08_in02 = reg_1081;
    123: op1_08_in02 = reg_0175;
    124: op1_08_in02 = reg_1277;
    126: op1_08_in02 = imem00_in[11:8];
    38: op1_08_in02 = reg_0621;
    127: op1_08_in02 = reg_0636;
    42: op1_08_in02 = imem01_in[7:4];
    128: op1_08_in02 = reg_1404;
    22: op1_08_in02 = reg_0031;
    130: op1_08_in02 = reg_0199;
    131: op1_08_in02 = reg_0005;
    default: op1_08_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv02 = 1;
    53: op1_08_inv02 = 1;
    69: op1_08_inv02 = 1;
    68: op1_08_inv02 = 1;
    61: op1_08_inv02 = 1;
    76: op1_08_inv02 = 1;
    58: op1_08_inv02 = 1;
    78: op1_08_inv02 = 1;
    70: op1_08_inv02 = 1;
    51: op1_08_inv02 = 1;
    88: op1_08_inv02 = 1;
    59: op1_08_inv02 = 1;
    33: op1_08_inv02 = 1;
    62: op1_08_inv02 = 1;
    63: op1_08_inv02 = 1;
    83: op1_08_inv02 = 1;
    64: op1_08_inv02 = 1;
    84: op1_08_inv02 = 1;
    65: op1_08_inv02 = 1;
    85: op1_08_inv02 = 1;
    37: op1_08_inv02 = 1;
    66: op1_08_inv02 = 1;
    91: op1_08_inv02 = 1;
    67: op1_08_inv02 = 1;
    92: op1_08_inv02 = 1;
    93: op1_08_inv02 = 1;
    94: op1_08_inv02 = 1;
    98: op1_08_inv02 = 1;
    40: op1_08_inv02 = 1;
    102: op1_08_inv02 = 1;
    103: op1_08_inv02 = 1;
    104: op1_08_inv02 = 1;
    106: op1_08_inv02 = 1;
    107: op1_08_inv02 = 1;
    108: op1_08_inv02 = 1;
    110: op1_08_inv02 = 1;
    113: op1_08_inv02 = 1;
    115: op1_08_inv02 = 1;
    117: op1_08_inv02 = 1;
    118: op1_08_inv02 = 1;
    34: op1_08_inv02 = 1;
    121: op1_08_inv02 = 1;
    122: op1_08_inv02 = 1;
    124: op1_08_inv02 = 1;
    38: op1_08_inv02 = 1;
    127: op1_08_inv02 = 1;
    128: op1_08_inv02 = 1;
    131: op1_08_inv02 = 1;
    default: op1_08_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in03 = reg_0317;
    53: op1_08_in03 = reg_0386;
    65: op1_08_in03 = reg_0386;
    55: op1_08_in03 = reg_0119;
    86: op1_08_in03 = reg_0898;
    73: op1_08_in03 = reg_1346;
    69: op1_08_in03 = reg_0290;
    49: op1_08_in03 = reg_0004;
    50: op1_08_in03 = reg_0093;
    54: op1_08_in03 = reg_0439;
    74: op1_08_in03 = imem00_in[15:12];
    93: op1_08_in03 = imem00_in[15:12];
    68: op1_08_in03 = reg_0107;
    71: op1_08_in03 = reg_0791;
    75: op1_08_in03 = reg_1279;
    122: op1_08_in03 = reg_1279;
    61: op1_08_in03 = reg_0293;
    56: op1_08_in03 = reg_0563;
    87: op1_08_in03 = reg_0279;
    76: op1_08_in03 = reg_1078;
    57: op1_08_in03 = reg_0152;
    77: op1_08_in03 = reg_1490;
    80: op1_08_in03 = reg_1490;
    58: op1_08_in03 = reg_0727;
    109: op1_08_in03 = reg_0727;
    78: op1_08_in03 = reg_0109;
    70: op1_08_in03 = reg_0970;
    51: op1_08_in03 = reg_0230;
    88: op1_08_in03 = reg_0597;
    46: op1_08_in03 = reg_0429;
    59: op1_08_in03 = reg_0582;
    79: op1_08_in03 = reg_0240;
    60: op1_08_in03 = reg_0411;
    33: op1_08_in03 = reg_0028;
    62: op1_08_in03 = reg_0701;
    48: op1_08_in03 = reg_0065;
    52: op1_08_in03 = reg_0045;
    81: op1_08_in03 = reg_0868;
    85: op1_08_in03 = reg_0868;
    63: op1_08_in03 = reg_0884;
    82: op1_08_in03 = reg_0334;
    89: op1_08_in03 = reg_1199;
    83: op1_08_in03 = reg_0616;
    64: op1_08_in03 = reg_0735;
    84: op1_08_in03 = imem05_in[7:4];
    90: op1_08_in03 = reg_0470;
    40: op1_08_in03 = reg_0470;
    37: op1_08_in03 = reg_0086;
    66: op1_08_in03 = reg_0088;
    91: op1_08_in03 = reg_0488;
    67: op1_08_in03 = imem04_in[3:0];
    92: op1_08_in03 = reg_0564;
    94: op1_08_in03 = reg_0140;
    95: op1_08_in03 = reg_1494;
    96: op1_08_in03 = reg_0665;
    97: op1_08_in03 = reg_0158;
    98: op1_08_in03 = reg_0631;
    99: op1_08_in03 = reg_0246;
    44: op1_08_in03 = reg_0567;
    100: op1_08_in03 = reg_0457;
    47: op1_08_in03 = reg_0650;
    101: op1_08_in03 = reg_1164;
    102: op1_08_in03 = imem00_in[7:4];
    103: op1_08_in03 = reg_0044;
    104: op1_08_in03 = reg_0600;
    105: op1_08_in03 = reg_1207;
    106: op1_08_in03 = reg_0922;
    107: op1_08_in03 = imem06_in[7:4];
    108: op1_08_in03 = reg_0363;
    110: op1_08_in03 = reg_0714;
    111: op1_08_in03 = reg_0845;
    112: op1_08_in03 = reg_1059;
    113: op1_08_in03 = reg_1456;
    114: op1_08_in03 = reg_0613;
    115: op1_08_in03 = reg_0261;
    116: op1_08_in03 = reg_0602;
    117: op1_08_in03 = reg_0329;
    118: op1_08_in03 = reg_0667;
    119: op1_08_in03 = reg_0792;
    128: op1_08_in03 = reg_0792;
    34: op1_08_in03 = reg_0366;
    120: op1_08_in03 = reg_0234;
    121: op1_08_in03 = reg_0485;
    123: op1_08_in03 = reg_0724;
    124: op1_08_in03 = reg_1028;
    125: op1_08_in03 = reg_0266;
    126: op1_08_in03 = reg_0186;
    38: op1_08_in03 = reg_0620;
    127: op1_08_in03 = reg_0194;
    42: op1_08_in03 = imem01_in[15:12];
    129: op1_08_in03 = reg_0080;
    22: op1_08_in03 = reg_0030;
    130: op1_08_in03 = reg_0698;
    131: op1_08_in03 = reg_0026;
    default: op1_08_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv03 = 1;
    53: op1_08_inv03 = 1;
    55: op1_08_inv03 = 1;
    69: op1_08_inv03 = 1;
    49: op1_08_inv03 = 1;
    50: op1_08_inv03 = 1;
    54: op1_08_inv03 = 1;
    61: op1_08_inv03 = 1;
    56: op1_08_inv03 = 1;
    87: op1_08_inv03 = 1;
    77: op1_08_inv03 = 1;
    78: op1_08_inv03 = 1;
    88: op1_08_inv03 = 1;
    79: op1_08_inv03 = 1;
    60: op1_08_inv03 = 1;
    62: op1_08_inv03 = 1;
    48: op1_08_inv03 = 1;
    81: op1_08_inv03 = 1;
    63: op1_08_inv03 = 1;
    82: op1_08_inv03 = 1;
    89: op1_08_inv03 = 1;
    83: op1_08_inv03 = 1;
    64: op1_08_inv03 = 1;
    65: op1_08_inv03 = 1;
    90: op1_08_inv03 = 1;
    91: op1_08_inv03 = 1;
    95: op1_08_inv03 = 1;
    96: op1_08_inv03 = 1;
    97: op1_08_inv03 = 1;
    98: op1_08_inv03 = 1;
    100: op1_08_inv03 = 1;
    101: op1_08_inv03 = 1;
    40: op1_08_inv03 = 1;
    105: op1_08_inv03 = 1;
    107: op1_08_inv03 = 1;
    108: op1_08_inv03 = 1;
    110: op1_08_inv03 = 1;
    112: op1_08_inv03 = 1;
    113: op1_08_inv03 = 1;
    114: op1_08_inv03 = 1;
    115: op1_08_inv03 = 1;
    118: op1_08_inv03 = 1;
    119: op1_08_inv03 = 1;
    121: op1_08_inv03 = 1;
    122: op1_08_inv03 = 1;
    123: op1_08_inv03 = 1;
    124: op1_08_inv03 = 1;
    125: op1_08_inv03 = 1;
    127: op1_08_inv03 = 1;
    128: op1_08_inv03 = 1;
    129: op1_08_inv03 = 1;
    22: op1_08_inv03 = 1;
    130: op1_08_inv03 = 1;
    default: op1_08_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in04 = reg_0754;
    53: op1_08_in04 = reg_0385;
    55: op1_08_in04 = reg_0152;
    86: op1_08_in04 = reg_0696;
    73: op1_08_in04 = reg_0014;
    69: op1_08_in04 = reg_0679;
    49: op1_08_in04 = reg_0123;
    50: op1_08_in04 = reg_0899;
    108: op1_08_in04 = reg_0899;
    54: op1_08_in04 = reg_0384;
    74: op1_08_in04 = reg_1278;
    68: op1_08_in04 = reg_0113;
    71: op1_08_in04 = reg_0866;
    75: op1_08_in04 = reg_1081;
    61: op1_08_in04 = reg_0155;
    56: op1_08_in04 = reg_0530;
    87: op1_08_in04 = reg_1495;
    76: op1_08_in04 = reg_1491;
    131: op1_08_in04 = reg_1491;
    57: op1_08_in04 = reg_0215;
    77: op1_08_in04 = reg_1242;
    58: op1_08_in04 = reg_0402;
    123: op1_08_in04 = reg_0402;
    78: op1_08_in04 = reg_0718;
    70: op1_08_in04 = reg_0972;
    51: op1_08_in04 = reg_0135;
    88: op1_08_in04 = reg_1301;
    99: op1_08_in04 = reg_1301;
    117: op1_08_in04 = reg_1301;
    46: op1_08_in04 = imem02_in[3:0];
    59: op1_08_in04 = reg_1143;
    79: op1_08_in04 = reg_0799;
    60: op1_08_in04 = reg_0582;
    80: op1_08_in04 = reg_0580;
    114: op1_08_in04 = reg_0580;
    33: op1_08_in04 = reg_0228;
    62: op1_08_in04 = reg_0445;
    48: op1_08_in04 = reg_0210;
    52: op1_08_in04 = reg_0940;
    81: op1_08_in04 = reg_1489;
    102: op1_08_in04 = reg_1489;
    63: op1_08_in04 = reg_0232;
    82: op1_08_in04 = reg_1070;
    89: op1_08_in04 = reg_1208;
    83: op1_08_in04 = reg_1487;
    64: op1_08_in04 = reg_0702;
    84: op1_08_in04 = reg_0392;
    65: op1_08_in04 = reg_0365;
    85: op1_08_in04 = reg_1277;
    90: op1_08_in04 = imem05_in[15:12];
    66: op1_08_in04 = reg_0044;
    91: op1_08_in04 = reg_1215;
    67: op1_08_in04 = imem04_in[11:8];
    92: op1_08_in04 = reg_1181;
    93: op1_08_in04 = reg_0672;
    94: op1_08_in04 = reg_0157;
    95: op1_08_in04 = reg_0556;
    96: op1_08_in04 = reg_0284;
    97: op1_08_in04 = reg_0924;
    98: op1_08_in04 = reg_0473;
    44: op1_08_in04 = reg_0318;
    100: op1_08_in04 = reg_1347;
    47: op1_08_in04 = reg_0567;
    101: op1_08_in04 = reg_0251;
    40: op1_08_in04 = reg_0721;
    103: op1_08_in04 = reg_0010;
    104: op1_08_in04 = reg_0145;
    105: op1_08_in04 = reg_0433;
    106: op1_08_in04 = reg_0894;
    107: op1_08_in04 = reg_0755;
    109: op1_08_in04 = reg_0400;
    110: op1_08_in04 = reg_0374;
    111: op1_08_in04 = reg_0423;
    112: op1_08_in04 = reg_0338;
    113: op1_08_in04 = reg_0042;
    115: op1_08_in04 = reg_0177;
    116: op1_08_in04 = reg_1346;
    118: op1_08_in04 = reg_0922;
    119: op1_08_in04 = reg_0300;
    34: op1_08_in04 = reg_0442;
    120: op1_08_in04 = reg_0375;
    121: op1_08_in04 = reg_1459;
    122: op1_08_in04 = reg_0748;
    124: op1_08_in04 = reg_1027;
    125: op1_08_in04 = reg_1514;
    126: op1_08_in04 = reg_0523;
    38: op1_08_in04 = reg_0592;
    127: op1_08_in04 = reg_0624;
    42: op1_08_in04 = reg_0291;
    128: op1_08_in04 = reg_1163;
    129: op1_08_in04 = reg_0162;
    22: op1_08_in04 = imem07_in[15:12];
    130: op1_08_in04 = reg_0268;
    default: op1_08_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv04 = 1;
    53: op1_08_inv04 = 1;
    55: op1_08_inv04 = 1;
    73: op1_08_inv04 = 1;
    49: op1_08_inv04 = 1;
    50: op1_08_inv04 = 1;
    54: op1_08_inv04 = 1;
    74: op1_08_inv04 = 1;
    71: op1_08_inv04 = 1;
    61: op1_08_inv04 = 1;
    56: op1_08_inv04 = 1;
    77: op1_08_inv04 = 1;
    88: op1_08_inv04 = 1;
    46: op1_08_inv04 = 1;
    59: op1_08_inv04 = 1;
    79: op1_08_inv04 = 1;
    60: op1_08_inv04 = 1;
    80: op1_08_inv04 = 1;
    48: op1_08_inv04 = 1;
    81: op1_08_inv04 = 1;
    63: op1_08_inv04 = 1;
    82: op1_08_inv04 = 1;
    89: op1_08_inv04 = 1;
    83: op1_08_inv04 = 1;
    64: op1_08_inv04 = 1;
    90: op1_08_inv04 = 1;
    66: op1_08_inv04 = 1;
    91: op1_08_inv04 = 1;
    97: op1_08_inv04 = 1;
    98: op1_08_inv04 = 1;
    47: op1_08_inv04 = 1;
    40: op1_08_inv04 = 1;
    102: op1_08_inv04 = 1;
    103: op1_08_inv04 = 1;
    104: op1_08_inv04 = 1;
    107: op1_08_inv04 = 1;
    108: op1_08_inv04 = 1;
    109: op1_08_inv04 = 1;
    110: op1_08_inv04 = 1;
    111: op1_08_inv04 = 1;
    115: op1_08_inv04 = 1;
    118: op1_08_inv04 = 1;
    119: op1_08_inv04 = 1;
    34: op1_08_inv04 = 1;
    121: op1_08_inv04 = 1;
    124: op1_08_inv04 = 1;
    38: op1_08_inv04 = 1;
    130: op1_08_inv04 = 1;
    default: op1_08_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in05 = imem06_in[15:12];
    53: op1_08_in05 = reg_0362;
    54: op1_08_in05 = reg_0362;
    55: op1_08_in05 = reg_0212;
    86: op1_08_in05 = reg_0032;
    73: op1_08_in05 = reg_0458;
    69: op1_08_in05 = reg_0457;
    50: op1_08_in05 = reg_0871;
    74: op1_08_in05 = reg_1279;
    68: op1_08_in05 = reg_0885;
    89: op1_08_in05 = reg_0885;
    71: op1_08_in05 = reg_1081;
    75: op1_08_in05 = reg_0552;
    77: op1_08_in05 = reg_0552;
    61: op1_08_in05 = reg_0172;
    56: op1_08_in05 = reg_0981;
    87: op1_08_in05 = reg_0999;
    76: op1_08_in05 = reg_1243;
    57: op1_08_in05 = reg_0213;
    58: op1_08_in05 = reg_0047;
    78: op1_08_in05 = reg_0624;
    70: op1_08_in05 = imem02_in[7:4];
    51: op1_08_in05 = reg_0162;
    88: op1_08_in05 = reg_1093;
    117: op1_08_in05 = reg_1093;
    46: op1_08_in05 = reg_0106;
    59: op1_08_in05 = reg_0535;
    79: op1_08_in05 = imem06_in[11:8];
    60: op1_08_in05 = imem04_in[11:8];
    80: op1_08_in05 = reg_1470;
    33: op1_08_in05 = reg_0053;
    62: op1_08_in05 = reg_0791;
    48: op1_08_in05 = reg_0208;
    52: op1_08_in05 = reg_0184;
    81: op1_08_in05 = reg_0841;
    63: op1_08_in05 = reg_0268;
    82: op1_08_in05 = reg_0939;
    83: op1_08_in05 = reg_1242;
    64: op1_08_in05 = reg_1164;
    84: op1_08_in05 = reg_0173;
    65: op1_08_in05 = reg_0291;
    85: op1_08_in05 = reg_0613;
    90: op1_08_in05 = reg_0736;
    66: op1_08_in05 = reg_0012;
    91: op1_08_in05 = reg_0281;
    67: op1_08_in05 = reg_0694;
    92: op1_08_in05 = reg_1180;
    93: op1_08_in05 = reg_1487;
    94: op1_08_in05 = reg_0923;
    95: op1_08_in05 = reg_0965;
    120: op1_08_in05 = reg_0965;
    96: op1_08_in05 = reg_0404;
    34: op1_08_in05 = reg_0404;
    97: op1_08_in05 = reg_0441;
    98: op1_08_in05 = reg_1098;
    99: op1_08_in05 = reg_0178;
    44: op1_08_in05 = reg_0539;
    100: op1_08_in05 = reg_0157;
    47: op1_08_in05 = reg_0066;
    101: op1_08_in05 = reg_0176;
    40: op1_08_in05 = reg_0466;
    102: op1_08_in05 = reg_0907;
    103: op1_08_in05 = reg_0456;
    104: op1_08_in05 = reg_0000;
    105: op1_08_in05 = reg_0326;
    106: op1_08_in05 = reg_0225;
    107: op1_08_in05 = reg_0269;
    108: op1_08_in05 = reg_0092;
    109: op1_08_in05 = reg_0335;
    110: op1_08_in05 = reg_0373;
    111: op1_08_in05 = reg_0138;
    112: op1_08_in05 = reg_0367;
    113: op1_08_in05 = reg_0044;
    114: op1_08_in05 = reg_0486;
    115: op1_08_in05 = reg_1001;
    116: op1_08_in05 = reg_0317;
    118: op1_08_in05 = reg_0892;
    119: op1_08_in05 = reg_0151;
    121: op1_08_in05 = reg_1205;
    122: op1_08_in05 = reg_0615;
    123: op1_08_in05 = reg_0043;
    124: op1_08_in05 = reg_0221;
    125: op1_08_in05 = reg_0492;
    126: op1_08_in05 = reg_1027;
    38: op1_08_in05 = reg_0103;
    127: op1_08_in05 = reg_0529;
    42: op1_08_in05 = reg_0277;
    128: op1_08_in05 = reg_0302;
    129: op1_08_in05 = reg_0634;
    22: op1_08_in05 = reg_0002;
    130: op1_08_in05 = reg_0862;
    131: op1_08_in05 = reg_0250;
    default: op1_08_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv05 = 1;
    53: op1_08_inv05 = 1;
    73: op1_08_inv05 = 1;
    69: op1_08_inv05 = 1;
    50: op1_08_inv05 = 1;
    54: op1_08_inv05 = 1;
    74: op1_08_inv05 = 1;
    68: op1_08_inv05 = 1;
    71: op1_08_inv05 = 1;
    75: op1_08_inv05 = 1;
    78: op1_08_inv05 = 1;
    70: op1_08_inv05 = 1;
    46: op1_08_inv05 = 1;
    59: op1_08_inv05 = 1;
    60: op1_08_inv05 = 1;
    80: op1_08_inv05 = 1;
    33: op1_08_inv05 = 1;
    48: op1_08_inv05 = 1;
    52: op1_08_inv05 = 1;
    63: op1_08_inv05 = 1;
    89: op1_08_inv05 = 1;
    83: op1_08_inv05 = 1;
    64: op1_08_inv05 = 1;
    84: op1_08_inv05 = 1;
    90: op1_08_inv05 = 1;
    66: op1_08_inv05 = 1;
    93: op1_08_inv05 = 1;
    94: op1_08_inv05 = 1;
    95: op1_08_inv05 = 1;
    98: op1_08_inv05 = 1;
    99: op1_08_inv05 = 1;
    47: op1_08_inv05 = 1;
    40: op1_08_inv05 = 1;
    102: op1_08_inv05 = 1;
    103: op1_08_inv05 = 1;
    105: op1_08_inv05 = 1;
    106: op1_08_inv05 = 1;
    109: op1_08_inv05 = 1;
    110: op1_08_inv05 = 1;
    111: op1_08_inv05 = 1;
    112: op1_08_inv05 = 1;
    115: op1_08_inv05 = 1;
    116: op1_08_inv05 = 1;
    117: op1_08_inv05 = 1;
    123: op1_08_inv05 = 1;
    124: op1_08_inv05 = 1;
    125: op1_08_inv05 = 1;
    130: op1_08_inv05 = 1;
    131: op1_08_inv05 = 1;
    default: op1_08_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in06 = reg_0192;
    53: op1_08_in06 = reg_0047;
    55: op1_08_in06 = reg_0214;
    86: op1_08_in06 = imem04_in[7:4];
    73: op1_08_in06 = reg_0377;
    69: op1_08_in06 = reg_1029;
    50: op1_08_in06 = reg_0874;
    54: op1_08_in06 = reg_0091;
    74: op1_08_in06 = reg_1078;
    68: op1_08_in06 = reg_0504;
    71: op1_08_in06 = reg_1241;
    75: op1_08_in06 = reg_0562;
    61: op1_08_in06 = reg_0725;
    56: op1_08_in06 = reg_0495;
    87: op1_08_in06 = reg_0559;
    76: op1_08_in06 = reg_0121;
    57: op1_08_in06 = reg_1170;
    77: op1_08_in06 = reg_1028;
    58: op1_08_in06 = reg_0093;
    78: op1_08_in06 = reg_0132;
    70: op1_08_in06 = imem02_in[11:8];
    51: op1_08_in06 = reg_1057;
    88: op1_08_in06 = reg_1208;
    99: op1_08_in06 = reg_1208;
    46: op1_08_in06 = reg_0382;
    59: op1_08_in06 = reg_0534;
    79: op1_08_in06 = imem06_in[15:12];
    60: op1_08_in06 = reg_0463;
    80: op1_08_in06 = reg_0218;
    33: op1_08_in06 = reg_0124;
    62: op1_08_in06 = reg_1279;
    48: op1_08_in06 = reg_0792;
    52: op1_08_in06 = reg_0130;
    81: op1_08_in06 = reg_0580;
    122: op1_08_in06 = reg_0580;
    63: op1_08_in06 = reg_0537;
    82: op1_08_in06 = reg_0938;
    92: op1_08_in06 = reg_0938;
    89: op1_08_in06 = reg_0479;
    83: op1_08_in06 = reg_0806;
    85: op1_08_in06 = reg_0806;
    64: op1_08_in06 = reg_0176;
    84: op1_08_in06 = reg_0131;
    65: op1_08_in06 = reg_0042;
    42: op1_08_in06 = reg_0042;
    90: op1_08_in06 = reg_0735;
    66: op1_08_in06 = reg_0662;
    91: op1_08_in06 = reg_0796;
    67: op1_08_in06 = reg_0208;
    93: op1_08_in06 = reg_0613;
    94: op1_08_in06 = reg_0489;
    44: op1_08_in06 = reg_0489;
    95: op1_08_in06 = reg_0314;
    96: op1_08_in06 = reg_0408;
    97: op1_08_in06 = reg_0002;
    98: op1_08_in06 = reg_0711;
    100: op1_08_in06 = reg_0921;
    106: op1_08_in06 = reg_0921;
    47: op1_08_in06 = reg_0182;
    101: op1_08_in06 = reg_0649;
    40: op1_08_in06 = reg_0633;
    102: op1_08_in06 = reg_0803;
    103: op1_08_in06 = imem02_in[3:0];
    104: op1_08_in06 = reg_0180;
    105: op1_08_in06 = reg_0778;
    107: op1_08_in06 = reg_1209;
    108: op1_08_in06 = reg_0400;
    109: op1_08_in06 = reg_0044;
    123: op1_08_in06 = reg_0044;
    110: op1_08_in06 = reg_0622;
    111: op1_08_in06 = reg_0608;
    112: op1_08_in06 = reg_0833;
    113: op1_08_in06 = reg_0626;
    114: op1_08_in06 = reg_1027;
    115: op1_08_in06 = reg_0234;
    116: op1_08_in06 = imem06_in[3:0];
    117: op1_08_in06 = reg_1199;
    118: op1_08_in06 = reg_0310;
    119: op1_08_in06 = reg_0039;
    34: op1_08_in06 = reg_0415;
    120: op1_08_in06 = reg_0070;
    121: op1_08_in06 = reg_1418;
    124: op1_08_in06 = reg_0886;
    125: op1_08_in06 = reg_0118;
    126: op1_08_in06 = reg_1454;
    131: op1_08_in06 = reg_1454;
    38: op1_08_in06 = reg_0100;
    127: op1_08_in06 = reg_0345;
    128: op1_08_in06 = reg_0066;
    129: op1_08_in06 = reg_0041;
    130: op1_08_in06 = reg_0837;
    default: op1_08_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_08_inv06 = 1;
    73: op1_08_inv06 = 1;
    69: op1_08_inv06 = 1;
    54: op1_08_inv06 = 1;
    75: op1_08_inv06 = 1;
    61: op1_08_inv06 = 1;
    87: op1_08_inv06 = 1;
    58: op1_08_inv06 = 1;
    51: op1_08_inv06 = 1;
    88: op1_08_inv06 = 1;
    59: op1_08_inv06 = 1;
    33: op1_08_inv06 = 1;
    48: op1_08_inv06 = 1;
    52: op1_08_inv06 = 1;
    81: op1_08_inv06 = 1;
    82: op1_08_inv06 = 1;
    83: op1_08_inv06 = 1;
    84: op1_08_inv06 = 1;
    90: op1_08_inv06 = 1;
    67: op1_08_inv06 = 1;
    92: op1_08_inv06 = 1;
    93: op1_08_inv06 = 1;
    95: op1_08_inv06 = 1;
    96: op1_08_inv06 = 1;
    97: op1_08_inv06 = 1;
    98: op1_08_inv06 = 1;
    99: op1_08_inv06 = 1;
    100: op1_08_inv06 = 1;
    47: op1_08_inv06 = 1;
    40: op1_08_inv06 = 1;
    103: op1_08_inv06 = 1;
    104: op1_08_inv06 = 1;
    105: op1_08_inv06 = 1;
    106: op1_08_inv06 = 1;
    107: op1_08_inv06 = 1;
    109: op1_08_inv06 = 1;
    110: op1_08_inv06 = 1;
    111: op1_08_inv06 = 1;
    112: op1_08_inv06 = 1;
    113: op1_08_inv06 = 1;
    115: op1_08_inv06 = 1;
    117: op1_08_inv06 = 1;
    118: op1_08_inv06 = 1;
    119: op1_08_inv06 = 1;
    120: op1_08_inv06 = 1;
    121: op1_08_inv06 = 1;
    125: op1_08_inv06 = 1;
    126: op1_08_inv06 = 1;
    127: op1_08_inv06 = 1;
    42: op1_08_inv06 = 1;
    130: op1_08_inv06 = 1;
    131: op1_08_inv06 = 1;
    default: op1_08_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in07 = reg_0870;
    53: op1_08_in07 = reg_0093;
    55: op1_08_in07 = reg_0213;
    86: op1_08_in07 = reg_1214;
    73: op1_08_in07 = reg_0795;
    69: op1_08_in07 = reg_0455;
    50: op1_08_in07 = reg_0290;
    54: op1_08_in07 = reg_0047;
    74: op1_08_in07 = reg_1243;
    68: op1_08_in07 = reg_0506;
    71: op1_08_in07 = imem00_in[15:12];
    75: op1_08_in07 = reg_1470;
    61: op1_08_in07 = reg_0881;
    56: op1_08_in07 = reg_0776;
    87: op1_08_in07 = reg_0154;
    76: op1_08_in07 = reg_0806;
    57: op1_08_in07 = reg_1096;
    77: op1_08_in07 = reg_0485;
    122: op1_08_in07 = reg_0485;
    58: op1_08_in07 = reg_0899;
    78: op1_08_in07 = reg_0165;
    70: op1_08_in07 = reg_0128;
    51: op1_08_in07 = reg_0226;
    88: op1_08_in07 = reg_0350;
    46: op1_08_in07 = reg_0903;
    59: op1_08_in07 = imem04_in[11:8];
    79: op1_08_in07 = reg_1468;
    60: op1_08_in07 = reg_0978;
    80: op1_08_in07 = reg_0293;
    62: op1_08_in07 = reg_1080;
    48: op1_08_in07 = reg_0793;
    52: op1_08_in07 = reg_0272;
    81: op1_08_in07 = reg_1028;
    63: op1_08_in07 = reg_0263;
    82: op1_08_in07 = reg_0986;
    92: op1_08_in07 = reg_0986;
    89: op1_08_in07 = reg_0291;
    83: op1_08_in07 = reg_0805;
    85: op1_08_in07 = reg_0805;
    64: op1_08_in07 = reg_0333;
    84: op1_08_in07 = reg_0794;
    65: op1_08_in07 = reg_0662;
    90: op1_08_in07 = reg_0315;
    66: op1_08_in07 = reg_0742;
    91: op1_08_in07 = reg_0421;
    40: op1_08_in07 = reg_0421;
    67: op1_08_in07 = reg_0252;
    93: op1_08_in07 = reg_0580;
    94: op1_08_in07 = reg_0665;
    95: op1_08_in07 = reg_0349;
    96: op1_08_in07 = reg_0100;
    97: op1_08_in07 = reg_0053;
    98: op1_08_in07 = reg_0801;
    99: op1_08_in07 = reg_0107;
    117: op1_08_in07 = reg_0107;
    44: op1_08_in07 = reg_0492;
    100: op1_08_in07 = reg_0489;
    47: op1_08_in07 = reg_0167;
    101: op1_08_in07 = reg_0630;
    102: op1_08_in07 = reg_0153;
    103: op1_08_in07 = imem02_in[11:8];
    104: op1_08_in07 = reg_0789;
    105: op1_08_in07 = reg_0971;
    106: op1_08_in07 = reg_1094;
    107: op1_08_in07 = reg_1437;
    108: op1_08_in07 = reg_0078;
    109: op1_08_in07 = reg_0785;
    110: op1_08_in07 = reg_0619;
    111: op1_08_in07 = reg_0588;
    112: op1_08_in07 = reg_0832;
    113: op1_08_in07 = reg_0877;
    114: op1_08_in07 = reg_0221;
    115: op1_08_in07 = reg_0000;
    116: op1_08_in07 = imem06_in[7:4];
    118: op1_08_in07 = reg_1440;
    119: op1_08_in07 = reg_0929;
    34: op1_08_in07 = reg_0620;
    120: op1_08_in07 = reg_1516;
    121: op1_08_in07 = reg_0887;
    123: op1_08_in07 = reg_0845;
    124: op1_08_in07 = reg_0353;
    125: op1_08_in07 = reg_0602;
    126: op1_08_in07 = reg_1227;
    38: op1_08_in07 = reg_0114;
    127: op1_08_in07 = reg_1228;
    42: op1_08_in07 = reg_0044;
    128: op1_08_in07 = reg_1259;
    129: op1_08_in07 = reg_0012;
    130: op1_08_in07 = reg_1340;
    131: op1_08_in07 = reg_1229;
    default: op1_08_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv07 = 1;
    55: op1_08_inv07 = 1;
    86: op1_08_inv07 = 1;
    69: op1_08_inv07 = 1;
    54: op1_08_inv07 = 1;
    74: op1_08_inv07 = 1;
    71: op1_08_inv07 = 1;
    77: op1_08_inv07 = 1;
    58: op1_08_inv07 = 1;
    78: op1_08_inv07 = 1;
    59: op1_08_inv07 = 1;
    79: op1_08_inv07 = 1;
    80: op1_08_inv07 = 1;
    62: op1_08_inv07 = 1;
    52: op1_08_inv07 = 1;
    81: op1_08_inv07 = 1;
    89: op1_08_inv07 = 1;
    66: op1_08_inv07 = 1;
    91: op1_08_inv07 = 1;
    67: op1_08_inv07 = 1;
    99: op1_08_inv07 = 1;
    44: op1_08_inv07 = 1;
    100: op1_08_inv07 = 1;
    101: op1_08_inv07 = 1;
    102: op1_08_inv07 = 1;
    106: op1_08_inv07 = 1;
    108: op1_08_inv07 = 1;
    109: op1_08_inv07 = 1;
    111: op1_08_inv07 = 1;
    112: op1_08_inv07 = 1;
    117: op1_08_inv07 = 1;
    118: op1_08_inv07 = 1;
    119: op1_08_inv07 = 1;
    34: op1_08_inv07 = 1;
    122: op1_08_inv07 = 1;
    123: op1_08_inv07 = 1;
    126: op1_08_inv07 = 1;
    127: op1_08_inv07 = 1;
    129: op1_08_inv07 = 1;
    131: op1_08_inv07 = 1;
    default: op1_08_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in08 = reg_0397;
    53: op1_08_in08 = reg_0724;
    55: op1_08_in08 = reg_0230;
    86: op1_08_in08 = reg_0406;
    73: op1_08_in08 = reg_0905;
    69: op1_08_in08 = reg_1018;
    50: op1_08_in08 = reg_0041;
    42: op1_08_in08 = reg_0041;
    54: op1_08_in08 = reg_0093;
    74: op1_08_in08 = reg_1241;
    68: op1_08_in08 = reg_0480;
    71: op1_08_in08 = reg_0250;
    75: op1_08_in08 = reg_0485;
    61: op1_08_in08 = reg_0887;
    56: op1_08_in08 = reg_0778;
    87: op1_08_in08 = reg_0179;
    76: op1_08_in08 = reg_1470;
    85: op1_08_in08 = reg_1470;
    57: op1_08_in08 = reg_1183;
    77: op1_08_in08 = reg_1453;
    58: op1_08_in08 = reg_0078;
    78: op1_08_in08 = reg_0269;
    70: op1_08_in08 = reg_0105;
    51: op1_08_in08 = reg_0672;
    88: op1_08_in08 = reg_1149;
    46: op1_08_in08 = reg_0712;
    59: op1_08_in08 = reg_1216;
    79: op1_08_in08 = reg_0120;
    60: op1_08_in08 = reg_1203;
    80: op1_08_in08 = reg_0249;
    62: op1_08_in08 = reg_0844;
    48: op1_08_in08 = reg_0736;
    52: op1_08_in08 = reg_0864;
    81: op1_08_in08 = reg_0927;
    63: op1_08_in08 = reg_1198;
    82: op1_08_in08 = reg_0477;
    89: op1_08_in08 = reg_0673;
    83: op1_08_in08 = reg_0218;
    64: op1_08_in08 = reg_1181;
    84: op1_08_in08 = reg_0303;
    65: op1_08_in08 = reg_0606;
    90: op1_08_in08 = reg_0702;
    66: op1_08_in08 = reg_1140;
    91: op1_08_in08 = reg_0407;
    67: op1_08_in08 = reg_0978;
    92: op1_08_in08 = reg_0301;
    93: op1_08_in08 = reg_0186;
    94: op1_08_in08 = reg_0661;
    106: op1_08_in08 = reg_0661;
    95: op1_08_in08 = reg_1300;
    96: op1_08_in08 = reg_0087;
    97: op1_08_in08 = reg_0085;
    98: op1_08_in08 = reg_0294;
    99: op1_08_in08 = reg_0880;
    44: op1_08_in08 = reg_0491;
    100: op1_08_in08 = reg_1094;
    47: op1_08_in08 = reg_0183;
    101: op1_08_in08 = reg_1180;
    40: op1_08_in08 = reg_0796;
    102: op1_08_in08 = reg_1027;
    103: op1_08_in08 = reg_0254;
    123: op1_08_in08 = reg_0254;
    104: op1_08_in08 = reg_0375;
    105: op1_08_in08 = reg_0111;
    107: op1_08_in08 = reg_0860;
    108: op1_08_in08 = reg_0634;
    109: op1_08_in08 = reg_1071;
    110: op1_08_in08 = reg_0132;
    111: op1_08_in08 = reg_0975;
    112: op1_08_in08 = reg_0332;
    113: op1_08_in08 = reg_0845;
    114: op1_08_in08 = reg_0961;
    115: op1_08_in08 = reg_1494;
    116: op1_08_in08 = imem06_in[15:12];
    117: op1_08_in08 = imem04_in[3:0];
    118: op1_08_in08 = reg_0309;
    119: op1_08_in08 = reg_0161;
    34: op1_08_in08 = reg_0103;
    120: op1_08_in08 = reg_1517;
    121: op1_08_in08 = reg_0188;
    122: op1_08_in08 = reg_1227;
    124: op1_08_in08 = reg_0431;
    125: op1_08_in08 = reg_0151;
    126: op1_08_in08 = reg_0987;
    38: op1_08_in08 = reg_0001;
    127: op1_08_in08 = reg_0244;
    128: op1_08_in08 = reg_0601;
    129: op1_08_in08 = reg_0011;
    130: op1_08_in08 = reg_0256;
    131: op1_08_in08 = reg_0821;
    default: op1_08_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_08_inv08 = 1;
    86: op1_08_inv08 = 1;
    50: op1_08_inv08 = 1;
    74: op1_08_inv08 = 1;
    61: op1_08_inv08 = 1;
    87: op1_08_inv08 = 1;
    57: op1_08_inv08 = 1;
    70: op1_08_inv08 = 1;
    59: op1_08_inv08 = 1;
    48: op1_08_inv08 = 1;
    81: op1_08_inv08 = 1;
    63: op1_08_inv08 = 1;
    82: op1_08_inv08 = 1;
    84: op1_08_inv08 = 1;
    66: op1_08_inv08 = 1;
    91: op1_08_inv08 = 1;
    92: op1_08_inv08 = 1;
    93: op1_08_inv08 = 1;
    94: op1_08_inv08 = 1;
    95: op1_08_inv08 = 1;
    96: op1_08_inv08 = 1;
    97: op1_08_inv08 = 1;
    102: op1_08_inv08 = 1;
    103: op1_08_inv08 = 1;
    107: op1_08_inv08 = 1;
    108: op1_08_inv08 = 1;
    110: op1_08_inv08 = 1;
    115: op1_08_inv08 = 1;
    117: op1_08_inv08 = 1;
    118: op1_08_inv08 = 1;
    34: op1_08_inv08 = 1;
    120: op1_08_inv08 = 1;
    122: op1_08_inv08 = 1;
    123: op1_08_inv08 = 1;
    125: op1_08_inv08 = 1;
    126: op1_08_inv08 = 1;
    38: op1_08_inv08 = 1;
    42: op1_08_inv08 = 1;
    130: op1_08_inv08 = 1;
    131: op1_08_inv08 = 1;
    default: op1_08_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in09 = reg_1334;
    119: op1_08_in09 = reg_1334;
    53: op1_08_in09 = reg_0875;
    55: op1_08_in09 = reg_0191;
    86: op1_08_in09 = reg_0451;
    73: op1_08_in09 = reg_0160;
    69: op1_08_in09 = reg_0589;
    50: op1_08_in09 = reg_0011;
    54: op1_08_in09 = reg_0724;
    74: op1_08_in09 = reg_0121;
    68: op1_08_in09 = imem03_in[11:8];
    71: op1_08_in09 = reg_0293;
    75: op1_08_in09 = reg_1454;
    61: op1_08_in09 = reg_0883;
    56: op1_08_in09 = reg_0127;
    87: op1_08_in09 = reg_0706;
    76: op1_08_in09 = reg_0987;
    57: op1_08_in09 = reg_0245;
    77: op1_08_in09 = reg_1201;
    58: op1_08_in09 = reg_0291;
    78: op1_08_in09 = reg_0271;
    70: op1_08_in09 = reg_0382;
    51: op1_08_in09 = reg_0777;
    88: op1_08_in09 = reg_0025;
    46: op1_08_in09 = reg_0294;
    59: op1_08_in09 = reg_1203;
    79: op1_08_in09 = reg_1209;
    60: op1_08_in09 = reg_1077;
    80: op1_08_in09 = reg_1417;
    122: op1_08_in09 = reg_1417;
    62: op1_08_in09 = reg_0841;
    48: op1_08_in09 = reg_0175;
    52: op1_08_in09 = reg_0151;
    81: op1_08_in09 = reg_0886;
    63: op1_08_in09 = reg_1083;
    82: op1_08_in09 = reg_1514;
    89: op1_08_in09 = reg_0534;
    83: op1_08_in09 = reg_1052;
    64: op1_08_in09 = reg_0540;
    84: op1_08_in09 = reg_0130;
    65: op1_08_in09 = reg_1018;
    85: op1_08_in09 = reg_1230;
    90: op1_08_in09 = reg_0332;
    66: op1_08_in09 = reg_1029;
    91: op1_08_in09 = reg_1041;
    67: op1_08_in09 = reg_1198;
    92: op1_08_in09 = reg_1484;
    93: op1_08_in09 = reg_0640;
    94: op1_08_in09 = reg_0441;
    95: op1_08_in09 = reg_1301;
    96: op1_08_in09 = reg_0521;
    97: op1_08_in09 = reg_1182;
    98: op1_08_in09 = reg_0007;
    99: op1_08_in09 = reg_0288;
    44: op1_08_in09 = imem05_in[15:12];
    100: op1_08_in09 = reg_0774;
    47: op1_08_in09 = reg_0240;
    101: op1_08_in09 = reg_0697;
    40: op1_08_in09 = reg_0369;
    102: op1_08_in09 = reg_1459;
    103: op1_08_in09 = reg_0822;
    104: op1_08_in09 = reg_0314;
    105: op1_08_in09 = reg_0629;
    106: op1_08_in09 = reg_0286;
    107: op1_08_in09 = reg_0869;
    108: op1_08_in09 = reg_0042;
    109: op1_08_in09 = reg_0662;
    42: op1_08_in09 = reg_0662;
    110: op1_08_in09 = reg_0165;
    111: op1_08_in09 = reg_0776;
    112: op1_08_in09 = reg_0333;
    113: op1_08_in09 = reg_0055;
    114: op1_08_in09 = reg_0460;
    115: op1_08_in09 = reg_1313;
    116: op1_08_in09 = reg_1030;
    117: op1_08_in09 = reg_0208;
    118: op1_08_in09 = reg_0159;
    34: op1_08_in09 = reg_0050;
    120: op1_08_in09 = reg_1447;
    121: op1_08_in09 = reg_0722;
    123: op1_08_in09 = reg_1493;
    124: op1_08_in09 = reg_0416;
    125: op1_08_in09 = reg_0206;
    126: op1_08_in09 = reg_1418;
    38: op1_08_in09 = reg_0085;
    127: op1_08_in09 = reg_0195;
    128: op1_08_in09 = reg_0393;
    129: op1_08_in09 = reg_0447;
    130: op1_08_in09 = reg_0096;
    131: op1_08_in09 = reg_0887;
    default: op1_08_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv09 = 1;
    53: op1_08_inv09 = 1;
    55: op1_08_inv09 = 1;
    86: op1_08_inv09 = 1;
    73: op1_08_inv09 = 1;
    69: op1_08_inv09 = 1;
    50: op1_08_inv09 = 1;
    54: op1_08_inv09 = 1;
    74: op1_08_inv09 = 1;
    68: op1_08_inv09 = 1;
    71: op1_08_inv09 = 1;
    75: op1_08_inv09 = 1;
    61: op1_08_inv09 = 1;
    87: op1_08_inv09 = 1;
    76: op1_08_inv09 = 1;
    57: op1_08_inv09 = 1;
    77: op1_08_inv09 = 1;
    58: op1_08_inv09 = 1;
    59: op1_08_inv09 = 1;
    60: op1_08_inv09 = 1;
    63: op1_08_inv09 = 1;
    64: op1_08_inv09 = 1;
    84: op1_08_inv09 = 1;
    65: op1_08_inv09 = 1;
    85: op1_08_inv09 = 1;
    67: op1_08_inv09 = 1;
    92: op1_08_inv09 = 1;
    94: op1_08_inv09 = 1;
    95: op1_08_inv09 = 1;
    96: op1_08_inv09 = 1;
    97: op1_08_inv09 = 1;
    99: op1_08_inv09 = 1;
    44: op1_08_inv09 = 1;
    47: op1_08_inv09 = 1;
    101: op1_08_inv09 = 1;
    40: op1_08_inv09 = 1;
    102: op1_08_inv09 = 1;
    103: op1_08_inv09 = 1;
    104: op1_08_inv09 = 1;
    106: op1_08_inv09 = 1;
    110: op1_08_inv09 = 1;
    111: op1_08_inv09 = 1;
    113: op1_08_inv09 = 1;
    114: op1_08_inv09 = 1;
    118: op1_08_inv09 = 1;
    122: op1_08_inv09 = 1;
    125: op1_08_inv09 = 1;
    127: op1_08_inv09 = 1;
    42: op1_08_inv09 = 1;
    default: op1_08_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in10 = reg_0869;
    79: op1_08_in10 = reg_0869;
    53: op1_08_in10 = reg_0291;
    55: op1_08_in10 = reg_0998;
    86: op1_08_in10 = reg_0097;
    73: op1_08_in10 = reg_0860;
    69: op1_08_in10 = reg_0560;
    50: op1_08_in10 = reg_0662;
    54: op1_08_in10 = reg_0899;
    74: op1_08_in10 = reg_1471;
    68: op1_08_in10 = reg_0247;
    71: op1_08_in10 = reg_1453;
    75: op1_08_in10 = reg_1432;
    77: op1_08_in10 = reg_1432;
    61: op1_08_in10 = reg_0350;
    95: op1_08_in10 = reg_0350;
    56: op1_08_in10 = reg_0112;
    87: op1_08_in10 = reg_0378;
    76: op1_08_in10 = reg_1205;
    57: op1_08_in10 = reg_0324;
    58: op1_08_in10 = reg_0012;
    78: op1_08_in10 = reg_0046;
    70: op1_08_in10 = reg_0381;
    51: op1_08_in10 = reg_0029;
    88: op1_08_in10 = reg_0218;
    46: op1_08_in10 = reg_0877;
    59: op1_08_in10 = reg_0676;
    60: op1_08_in10 = reg_1083;
    80: op1_08_in10 = reg_0524;
    62: op1_08_in10 = reg_0804;
    48: op1_08_in10 = reg_0646;
    52: op1_08_in10 = reg_0204;
    81: op1_08_in10 = reg_0202;
    131: op1_08_in10 = reg_0202;
    63: op1_08_in10 = reg_0414;
    82: op1_08_in10 = reg_1346;
    89: op1_08_in10 = reg_0341;
    83: op1_08_in10 = reg_0250;
    64: op1_08_in10 = reg_0538;
    84: op1_08_in10 = reg_0631;
    65: op1_08_in10 = reg_0563;
    85: op1_08_in10 = reg_1229;
    90: op1_08_in10 = reg_0333;
    66: op1_08_in10 = reg_0497;
    91: op1_08_in10 = reg_1151;
    67: op1_08_in10 = reg_1077;
    92: op1_08_in10 = reg_0344;
    93: op1_08_in10 = reg_1206;
    94: op1_08_in10 = reg_0741;
    98: op1_08_in10 = reg_0255;
    99: op1_08_in10 = reg_0088;
    44: op1_08_in10 = reg_0090;
    100: op1_08_in10 = reg_0663;
    47: op1_08_in10 = reg_0151;
    101: op1_08_in10 = reg_0318;
    40: op1_08_in10 = reg_0304;
    102: op1_08_in10 = reg_0987;
    103: op1_08_in10 = reg_0256;
    104: op1_08_in10 = reg_0178;
    105: op1_08_in10 = reg_0007;
    106: op1_08_in10 = reg_0437;
    107: op1_08_in10 = reg_0115;
    108: op1_08_in10 = reg_0011;
    109: op1_08_in10 = reg_0327;
    110: op1_08_in10 = reg_0754;
    111: op1_08_in10 = reg_0778;
    123: op1_08_in10 = reg_0778;
    112: op1_08_in10 = reg_0347;
    113: op1_08_in10 = reg_0898;
    114: op1_08_in10 = reg_0881;
    115: op1_08_in10 = reg_0952;
    116: op1_08_in10 = reg_1058;
    117: op1_08_in10 = reg_0534;
    118: op1_08_in10 = reg_0921;
    119: op1_08_in10 = reg_1420;
    34: op1_08_in10 = reg_0051;
    120: op1_08_in10 = reg_1301;
    121: op1_08_in10 = reg_0134;
    122: op1_08_in10 = reg_1418;
    124: op1_08_in10 = reg_0388;
    125: op1_08_in10 = reg_0270;
    126: op1_08_in10 = reg_0459;
    38: op1_08_in10 = reg_0519;
    127: op1_08_in10 = reg_0084;
    42: op1_08_in10 = reg_0254;
    128: op1_08_in10 = reg_0206;
    129: op1_08_in10 = reg_0659;
    130: op1_08_in10 = reg_0536;
    default: op1_08_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv10 = 1;
    55: op1_08_inv10 = 1;
    73: op1_08_inv10 = 1;
    69: op1_08_inv10 = 1;
    50: op1_08_inv10 = 1;
    74: op1_08_inv10 = 1;
    75: op1_08_inv10 = 1;
    56: op1_08_inv10 = 1;
    87: op1_08_inv10 = 1;
    76: op1_08_inv10 = 1;
    57: op1_08_inv10 = 1;
    77: op1_08_inv10 = 1;
    88: op1_08_inv10 = 1;
    60: op1_08_inv10 = 1;
    83: op1_08_inv10 = 1;
    91: op1_08_inv10 = 1;
    94: op1_08_inv10 = 1;
    95: op1_08_inv10 = 1;
    47: op1_08_inv10 = 1;
    101: op1_08_inv10 = 1;
    104: op1_08_inv10 = 1;
    105: op1_08_inv10 = 1;
    107: op1_08_inv10 = 1;
    113: op1_08_inv10 = 1;
    119: op1_08_inv10 = 1;
    34: op1_08_inv10 = 1;
    120: op1_08_inv10 = 1;
    121: op1_08_inv10 = 1;
    124: op1_08_inv10 = 1;
    126: op1_08_inv10 = 1;
    128: op1_08_inv10 = 1;
    129: op1_08_inv10 = 1;
    130: op1_08_inv10 = 1;
    default: op1_08_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in11 = reg_0585;
    53: op1_08_in11 = reg_0282;
    55: op1_08_in11 = imem07_in[7:4];
    86: op1_08_in11 = reg_0582;
    73: op1_08_in11 = reg_1323;
    69: op1_08_in11 = reg_0494;
    50: op1_08_in11 = reg_0255;
    54: op1_08_in11 = reg_0080;
    74: op1_08_in11 = reg_1406;
    126: op1_08_in11 = reg_1406;
    68: op1_08_in11 = reg_0341;
    71: op1_08_in11 = reg_1205;
    75: op1_08_in11 = reg_1405;
    122: op1_08_in11 = reg_1405;
    61: op1_08_in11 = reg_0071;
    56: op1_08_in11 = reg_0382;
    87: op1_08_in11 = reg_0145;
    76: op1_08_in11 = reg_0821;
    57: op1_08_in11 = reg_0893;
    77: op1_08_in11 = reg_0229;
    58: op1_08_in11 = reg_0446;
    78: op1_08_in11 = reg_0152;
    70: op1_08_in11 = reg_0379;
    51: op1_08_in11 = reg_0286;
    88: op1_08_in11 = reg_0288;
    46: op1_08_in11 = reg_0024;
    59: op1_08_in11 = reg_0414;
    79: op1_08_in11 = reg_1504;
    60: op1_08_in11 = reg_0681;
    80: op1_08_in11 = reg_0883;
    62: op1_08_in11 = reg_0805;
    48: op1_08_in11 = reg_0066;
    52: op1_08_in11 = reg_0207;
    81: op1_08_in11 = reg_0722;
    63: op1_08_in11 = reg_0407;
    82: op1_08_in11 = reg_0589;
    92: op1_08_in11 = reg_0589;
    42: op1_08_in11 = reg_0589;
    89: op1_08_in11 = reg_0032;
    83: op1_08_in11 = reg_1459;
    64: op1_08_in11 = reg_0896;
    84: op1_08_in11 = reg_0864;
    65: op1_08_in11 = reg_0474;
    85: op1_08_in11 = reg_1206;
    90: op1_08_in11 = reg_0395;
    112: op1_08_in11 = reg_0395;
    66: op1_08_in11 = reg_0981;
    91: op1_08_in11 = reg_0236;
    67: op1_08_in11 = reg_1147;
    93: op1_08_in11 = reg_0155;
    94: op1_08_in11 = reg_0740;
    95: op1_08_in11 = reg_0378;
    98: op1_08_in11 = reg_0507;
    99: op1_08_in11 = reg_0500;
    44: op1_08_in11 = reg_0873;
    100: op1_08_in11 = reg_0285;
    47: op1_08_in11 = imem06_in[11:8];
    101: op1_08_in11 = reg_1486;
    40: op1_08_in11 = reg_0199;
    102: op1_08_in11 = reg_1432;
    103: op1_08_in11 = reg_0433;
    104: op1_08_in11 = reg_0882;
    105: op1_08_in11 = reg_0008;
    106: op1_08_in11 = reg_0739;
    107: op1_08_in11 = reg_0637;
    108: op1_08_in11 = reg_1068;
    109: op1_08_in11 = reg_1018;
    110: op1_08_in11 = reg_0212;
    111: op1_08_in11 = reg_1455;
    123: op1_08_in11 = reg_1455;
    113: op1_08_in11 = reg_0054;
    114: op1_08_in11 = reg_0435;
    115: op1_08_in11 = reg_1447;
    116: op1_08_in11 = reg_0929;
    117: op1_08_in11 = reg_0694;
    118: op1_08_in11 = reg_0489;
    119: op1_08_in11 = reg_0271;
    34: op1_08_in11 = reg_0085;
    120: op1_08_in11 = reg_1092;
    121: op1_08_in11 = reg_0005;
    124: op1_08_in11 = reg_0267;
    125: op1_08_in11 = reg_0333;
    38: op1_08_in11 = reg_0518;
    127: op1_08_in11 = reg_1055;
    128: op1_08_in11 = reg_1299;
    129: op1_08_in11 = reg_0495;
    130: op1_08_in11 = reg_1488;
    131: op1_08_in11 = reg_0352;
    default: op1_08_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv11 = 1;
    53: op1_08_inv11 = 1;
    73: op1_08_inv11 = 1;
    68: op1_08_inv11 = 1;
    71: op1_08_inv11 = 1;
    61: op1_08_inv11 = 1;
    87: op1_08_inv11 = 1;
    76: op1_08_inv11 = 1;
    77: op1_08_inv11 = 1;
    58: op1_08_inv11 = 1;
    51: op1_08_inv11 = 1;
    88: op1_08_inv11 = 1;
    59: op1_08_inv11 = 1;
    79: op1_08_inv11 = 1;
    48: op1_08_inv11 = 1;
    52: op1_08_inv11 = 1;
    81: op1_08_inv11 = 1;
    63: op1_08_inv11 = 1;
    64: op1_08_inv11 = 1;
    85: op1_08_inv11 = 1;
    91: op1_08_inv11 = 1;
    95: op1_08_inv11 = 1;
    98: op1_08_inv11 = 1;
    99: op1_08_inv11 = 1;
    100: op1_08_inv11 = 1;
    101: op1_08_inv11 = 1;
    104: op1_08_inv11 = 1;
    105: op1_08_inv11 = 1;
    106: op1_08_inv11 = 1;
    107: op1_08_inv11 = 1;
    108: op1_08_inv11 = 1;
    109: op1_08_inv11 = 1;
    111: op1_08_inv11 = 1;
    113: op1_08_inv11 = 1;
    115: op1_08_inv11 = 1;
    116: op1_08_inv11 = 1;
    117: op1_08_inv11 = 1;
    118: op1_08_inv11 = 1;
    34: op1_08_inv11 = 1;
    120: op1_08_inv11 = 1;
    123: op1_08_inv11 = 1;
    125: op1_08_inv11 = 1;
    42: op1_08_inv11 = 1;
    default: op1_08_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in12 = reg_0622;
    53: op1_08_in12 = reg_0012;
    55: op1_08_in12 = reg_0225;
    86: op1_08_in12 = reg_0340;
    73: op1_08_in12 = imem06_in[3:0];
    69: op1_08_in12 = reg_0971;
    50: op1_08_in12 = reg_0631;
    54: op1_08_in12 = reg_0077;
    74: op1_08_in12 = reg_1405;
    68: op1_08_in12 = reg_1383;
    71: op1_08_in12 = reg_0887;
    75: op1_08_in12 = reg_0476;
    93: op1_08_in12 = reg_0476;
    61: op1_08_in12 = reg_0059;
    56: op1_08_in12 = reg_0708;
    87: op1_08_in12 = reg_0314;
    76: op1_08_in12 = reg_0881;
    57: op1_08_in12 = reg_0867;
    77: op1_08_in12 = reg_0155;
    58: op1_08_in12 = reg_0486;
    78: op1_08_in12 = reg_0213;
    70: op1_08_in12 = reg_0897;
    51: op1_08_in12 = reg_0740;
    88: op1_08_in12 = reg_0427;
    46: op1_08_in12 = reg_0217;
    59: op1_08_in12 = reg_0797;
    79: op1_08_in12 = reg_0116;
    60: op1_08_in12 = reg_0552;
    80: op1_08_in12 = reg_0201;
    62: op1_08_in12 = reg_1027;
    48: op1_08_in12 = reg_0182;
    52: op1_08_in12 = reg_0014;
    81: op1_08_in12 = reg_0416;
    63: op1_08_in12 = reg_0598;
    82: op1_08_in12 = reg_0206;
    84: op1_08_in12 = reg_0206;
    89: op1_08_in12 = reg_0493;
    83: op1_08_in12 = reg_1417;
    64: op1_08_in12 = reg_0895;
    108: op1_08_in12 = reg_0895;
    65: op1_08_in12 = reg_0326;
    85: op1_08_in12 = reg_0927;
    90: op1_08_in12 = reg_0700;
    66: op1_08_in12 = reg_1260;
    91: op1_08_in12 = reg_0063;
    67: op1_08_in12 = reg_0412;
    92: op1_08_in12 = imem06_in[11:8];
    94: op1_08_in12 = reg_0137;
    95: op1_08_in12 = reg_1282;
    98: op1_08_in12 = reg_0999;
    99: op1_08_in12 = reg_1147;
    44: op1_08_in12 = reg_0251;
    100: op1_08_in12 = reg_0413;
    47: op1_08_in12 = reg_0120;
    101: op1_08_in12 = reg_0197;
    40: op1_08_in12 = imem04_in[11:8];
    102: op1_08_in12 = reg_1418;
    103: op1_08_in12 = reg_1450;
    104: op1_08_in12 = reg_1009;
    105: op1_08_in12 = reg_1448;
    106: op1_08_in12 = reg_0103;
    107: op1_08_in12 = reg_1228;
    109: op1_08_in12 = reg_0839;
    110: op1_08_in12 = reg_0215;
    111: op1_08_in12 = reg_0111;
    123: op1_08_in12 = reg_0111;
    112: op1_08_in12 = reg_0176;
    113: op1_08_in12 = reg_0776;
    114: op1_08_in12 = reg_0409;
    115: op1_08_in12 = reg_0756;
    116: op1_08_in12 = reg_0669;
    117: op1_08_in12 = reg_1083;
    118: op1_08_in12 = reg_0224;
    119: op1_08_in12 = reg_0827;
    34: op1_08_in12 = reg_0519;
    120: op1_08_in12 = reg_0790;
    121: op1_08_in12 = reg_0267;
    122: op1_08_in12 = reg_1393;
    124: op1_08_in12 = reg_1152;
    125: op1_08_in12 = reg_0372;
    126: op1_08_in12 = reg_0886;
    127: op1_08_in12 = reg_0050;
    42: op1_08_in12 = reg_0531;
    128: op1_08_in12 = reg_0261;
    129: op1_08_in12 = reg_0399;
    130: op1_08_in12 = reg_0038;
    131: op1_08_in12 = reg_0440;
    default: op1_08_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv12 = 1;
    53: op1_08_inv12 = 1;
    86: op1_08_inv12 = 1;
    68: op1_08_inv12 = 1;
    71: op1_08_inv12 = 1;
    75: op1_08_inv12 = 1;
    58: op1_08_inv12 = 1;
    88: op1_08_inv12 = 1;
    46: op1_08_inv12 = 1;
    79: op1_08_inv12 = 1;
    60: op1_08_inv12 = 1;
    80: op1_08_inv12 = 1;
    62: op1_08_inv12 = 1;
    48: op1_08_inv12 = 1;
    81: op1_08_inv12 = 1;
    63: op1_08_inv12 = 1;
    64: op1_08_inv12 = 1;
    84: op1_08_inv12 = 1;
    90: op1_08_inv12 = 1;
    66: op1_08_inv12 = 1;
    91: op1_08_inv12 = 1;
    92: op1_08_inv12 = 1;
    94: op1_08_inv12 = 1;
    98: op1_08_inv12 = 1;
    99: op1_08_inv12 = 1;
    100: op1_08_inv12 = 1;
    47: op1_08_inv12 = 1;
    101: op1_08_inv12 = 1;
    40: op1_08_inv12 = 1;
    103: op1_08_inv12 = 1;
    104: op1_08_inv12 = 1;
    105: op1_08_inv12 = 1;
    106: op1_08_inv12 = 1;
    109: op1_08_inv12 = 1;
    111: op1_08_inv12 = 1;
    113: op1_08_inv12 = 1;
    115: op1_08_inv12 = 1;
    116: op1_08_inv12 = 1;
    117: op1_08_inv12 = 1;
    118: op1_08_inv12 = 1;
    34: op1_08_inv12 = 1;
    122: op1_08_inv12 = 1;
    123: op1_08_inv12 = 1;
    124: op1_08_inv12 = 1;
    42: op1_08_inv12 = 1;
    128: op1_08_inv12 = 1;
    129: op1_08_inv12 = 1;
    130: op1_08_inv12 = 1;
    default: op1_08_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in13 = reg_0624;
    53: op1_08_in13 = reg_0662;
    58: op1_08_in13 = reg_0662;
    55: op1_08_in13 = reg_0310;
    86: op1_08_in13 = reg_0487;
    73: op1_08_in13 = reg_0714;
    69: op1_08_in13 = reg_0626;
    50: op1_08_in13 = imem02_in[3:0];
    109: op1_08_in13 = imem02_in[3:0];
    54: op1_08_in13 = reg_0290;
    74: op1_08_in13 = reg_0883;
    76: op1_08_in13 = reg_0883;
    68: op1_08_in13 = reg_1258;
    71: op1_08_in13 = reg_0202;
    75: op1_08_in13 = reg_0887;
    61: op1_08_in13 = reg_0058;
    56: op1_08_in13 = reg_0153;
    87: op1_08_in13 = reg_0349;
    57: op1_08_in13 = reg_0309;
    77: op1_08_in13 = reg_0927;
    78: op1_08_in13 = imem07_in[3:0];
    110: op1_08_in13 = imem07_in[3:0];
    70: op1_08_in13 = reg_0846;
    51: op1_08_in13 = reg_0415;
    88: op1_08_in13 = imem04_in[7:4];
    46: op1_08_in13 = reg_0069;
    59: op1_08_in13 = reg_0341;
    79: op1_08_in13 = reg_0110;
    60: op1_08_in13 = reg_0421;
    99: op1_08_in13 = reg_0421;
    80: op1_08_in13 = reg_0428;
    85: op1_08_in13 = reg_0428;
    62: op1_08_in13 = reg_0221;
    48: op1_08_in13 = reg_0331;
    124: op1_08_in13 = reg_0331;
    52: op1_08_in13 = reg_0931;
    81: op1_08_in13 = reg_0134;
    63: op1_08_in13 = reg_0796;
    82: op1_08_in13 = reg_1468;
    89: op1_08_in13 = reg_0535;
    83: op1_08_in13 = reg_0821;
    102: op1_08_in13 = reg_0821;
    64: op1_08_in13 = reg_0090;
    84: op1_08_in13 = reg_1064;
    65: op1_08_in13 = reg_0106;
    90: op1_08_in13 = reg_0604;
    66: op1_08_in13 = reg_0631;
    91: op1_08_in13 = reg_0370;
    67: op1_08_in13 = reg_0406;
    92: op1_08_in13 = reg_0195;
    93: op1_08_in13 = reg_0928;
    94: op1_08_in13 = reg_0100;
    95: op1_08_in13 = reg_1280;
    120: op1_08_in13 = reg_1280;
    98: op1_08_in13 = reg_0233;
    44: op1_08_in13 = reg_0197;
    100: op1_08_in13 = reg_0623;
    47: op1_08_in13 = reg_0141;
    101: op1_08_in13 = reg_0196;
    40: op1_08_in13 = imem04_in[15:12];
    103: op1_08_in13 = reg_0745;
    104: op1_08_in13 = reg_0218;
    105: op1_08_in13 = reg_0312;
    106: op1_08_in13 = reg_0050;
    107: op1_08_in13 = reg_0289;
    108: op1_08_in13 = reg_0530;
    111: op1_08_in13 = reg_0496;
    112: op1_08_in13 = reg_0066;
    113: op1_08_in13 = reg_0128;
    114: op1_08_in13 = reg_0075;
    115: op1_08_in13 = reg_0962;
    116: op1_08_in13 = reg_0782;
    117: op1_08_in13 = reg_1200;
    118: op1_08_in13 = reg_0777;
    119: op1_08_in13 = reg_0265;
    34: op1_08_in13 = reg_0520;
    121: op1_08_in13 = reg_1255;
    122: op1_08_in13 = reg_0188;
    123: op1_08_in13 = reg_0379;
    125: op1_08_in13 = reg_0669;
    126: op1_08_in13 = reg_0351;
    127: op1_08_in13 = reg_1056;
    42: op1_08_in13 = reg_0497;
    128: op1_08_in13 = reg_1467;
    129: op1_08_in13 = reg_0879;
    130: op1_08_in13 = imem05_in[15:12];
    131: op1_08_in13 = reg_0122;
    default: op1_08_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_08_inv13 = 1;
    73: op1_08_inv13 = 1;
    50: op1_08_inv13 = 1;
    54: op1_08_inv13 = 1;
    68: op1_08_inv13 = 1;
    71: op1_08_inv13 = 1;
    75: op1_08_inv13 = 1;
    61: op1_08_inv13 = 1;
    56: op1_08_inv13 = 1;
    58: op1_08_inv13 = 1;
    70: op1_08_inv13 = 1;
    60: op1_08_inv13 = 1;
    80: op1_08_inv13 = 1;
    62: op1_08_inv13 = 1;
    81: op1_08_inv13 = 1;
    63: op1_08_inv13 = 1;
    82: op1_08_inv13 = 1;
    89: op1_08_inv13 = 1;
    83: op1_08_inv13 = 1;
    64: op1_08_inv13 = 1;
    65: op1_08_inv13 = 1;
    85: op1_08_inv13 = 1;
    90: op1_08_inv13 = 1;
    67: op1_08_inv13 = 1;
    95: op1_08_inv13 = 1;
    98: op1_08_inv13 = 1;
    99: op1_08_inv13 = 1;
    100: op1_08_inv13 = 1;
    105: op1_08_inv13 = 1;
    109: op1_08_inv13 = 1;
    114: op1_08_inv13 = 1;
    116: op1_08_inv13 = 1;
    117: op1_08_inv13 = 1;
    118: op1_08_inv13 = 1;
    119: op1_08_inv13 = 1;
    120: op1_08_inv13 = 1;
    126: op1_08_inv13 = 1;
    127: op1_08_inv13 = 1;
    129: op1_08_inv13 = 1;
    131: op1_08_inv13 = 1;
    default: op1_08_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in14 = reg_0132;
    53: op1_08_in14 = reg_0133;
    55: op1_08_in14 = reg_0867;
    86: op1_08_in14 = reg_0336;
    73: op1_08_in14 = reg_0585;
    69: op1_08_in14 = reg_0935;
    50: op1_08_in14 = reg_0975;
    54: op1_08_in14 = reg_0291;
    74: op1_08_in14 = reg_0188;
    68: op1_08_in14 = reg_1065;
    71: op1_08_in14 = reg_0431;
    85: op1_08_in14 = reg_0431;
    75: op1_08_in14 = reg_0351;
    61: op1_08_in14 = reg_0005;
    56: op1_08_in14 = reg_0008;
    87: op1_08_in14 = reg_0246;
    76: op1_08_in14 = reg_0202;
    57: op1_08_in14 = reg_0673;
    77: op1_08_in14 = reg_0883;
    102: op1_08_in14 = reg_0883;
    58: op1_08_in14 = reg_0632;
    78: op1_08_in14 = reg_0706;
    70: op1_08_in14 = reg_0327;
    51: op1_08_in14 = reg_0620;
    88: op1_08_in14 = imem04_in[11:8];
    46: op1_08_in14 = reg_0325;
    59: op1_08_in14 = reg_0305;
    79: op1_08_in14 = reg_0398;
    60: op1_08_in14 = reg_0414;
    80: op1_08_in14 = reg_0440;
    62: op1_08_in14 = reg_1230;
    48: op1_08_in14 = reg_0332;
    52: op1_08_in14 = reg_0866;
    81: op1_08_in14 = reg_0389;
    63: op1_08_in14 = reg_0370;
    82: op1_08_in14 = reg_0120;
    89: op1_08_in14 = reg_0531;
    83: op1_08_in14 = reg_0881;
    64: op1_08_in14 = reg_0872;
    84: op1_08_in14 = reg_0905;
    65: op1_08_in14 = reg_0380;
    90: op1_08_in14 = reg_0392;
    66: op1_08_in14 = reg_1207;
    91: op1_08_in14 = reg_0750;
    67: op1_08_in14 = reg_0797;
    92: op1_08_in14 = reg_1064;
    93: op1_08_in14 = reg_0887;
    94: op1_08_in14 = reg_0004;
    95: op1_08_in14 = reg_1368;
    98: op1_08_in14 = reg_0699;
    99: op1_08_in14 = reg_0599;
    44: op1_08_in14 = reg_0243;
    100: op1_08_in14 = reg_0591;
    47: op1_08_in14 = reg_0397;
    125: op1_08_in14 = reg_0397;
    101: op1_08_in14 = reg_1348;
    40: op1_08_in14 = reg_0096;
    103: op1_08_in14 = reg_0560;
    104: op1_08_in14 = reg_0427;
    105: op1_08_in14 = reg_0144;
    106: op1_08_in14 = reg_0003;
    107: op1_08_in14 = reg_0165;
    108: op1_08_in14 = reg_0138;
    109: op1_08_in14 = imem02_in[15:12];
    110: op1_08_in14 = imem07_in[7:4];
    111: op1_08_in14 = reg_0878;
    112: op1_08_in14 = reg_0167;
    113: op1_08_in14 = reg_1140;
    114: op1_08_in14 = reg_0059;
    115: op1_08_in14 = reg_1301;
    116: op1_08_in14 = reg_0696;
    117: op1_08_in14 = reg_0681;
    118: op1_08_in14 = reg_0774;
    119: op1_08_in14 = reg_0780;
    34: op1_08_in14 = reg_0483;
    120: op1_08_in14 = reg_0425;
    121: op1_08_in14 = imem01_in[7:4];
    122: op1_08_in14 = reg_0416;
    123: op1_08_in14 = reg_1492;
    124: op1_08_in14 = reg_0746;
    126: op1_08_in14 = reg_0409;
    127: op1_08_in14 = reg_0140;
    42: op1_08_in14 = reg_0128;
    128: op1_08_in14 = reg_0265;
    129: op1_08_in14 = reg_0934;
    130: op1_08_in14 = reg_0648;
    131: op1_08_in14 = reg_0238;
    default: op1_08_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_08_inv14 = 1;
    55: op1_08_inv14 = 1;
    50: op1_08_inv14 = 1;
    74: op1_08_inv14 = 1;
    68: op1_08_inv14 = 1;
    71: op1_08_inv14 = 1;
    61: op1_08_inv14 = 1;
    76: op1_08_inv14 = 1;
    77: op1_08_inv14 = 1;
    58: op1_08_inv14 = 1;
    78: op1_08_inv14 = 1;
    79: op1_08_inv14 = 1;
    60: op1_08_inv14 = 1;
    80: op1_08_inv14 = 1;
    62: op1_08_inv14 = 1;
    81: op1_08_inv14 = 1;
    89: op1_08_inv14 = 1;
    83: op1_08_inv14 = 1;
    64: op1_08_inv14 = 1;
    84: op1_08_inv14 = 1;
    85: op1_08_inv14 = 1;
    90: op1_08_inv14 = 1;
    67: op1_08_inv14 = 1;
    93: op1_08_inv14 = 1;
    94: op1_08_inv14 = 1;
    98: op1_08_inv14 = 1;
    99: op1_08_inv14 = 1;
    100: op1_08_inv14 = 1;
    102: op1_08_inv14 = 1;
    103: op1_08_inv14 = 1;
    104: op1_08_inv14 = 1;
    105: op1_08_inv14 = 1;
    110: op1_08_inv14 = 1;
    112: op1_08_inv14 = 1;
    114: op1_08_inv14 = 1;
    115: op1_08_inv14 = 1;
    116: op1_08_inv14 = 1;
    118: op1_08_inv14 = 1;
    119: op1_08_inv14 = 1;
    34: op1_08_inv14 = 1;
    123: op1_08_inv14 = 1;
    125: op1_08_inv14 = 1;
    127: op1_08_inv14 = 1;
    42: op1_08_inv14 = 1;
    129: op1_08_inv14 = 1;
    130: op1_08_inv14 = 1;
    131: op1_08_inv14 = 1;
    default: op1_08_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in15 = reg_0171;
    53: op1_08_in15 = reg_0606;
    55: op1_08_in15 = reg_0297;
    86: op1_08_in15 = reg_0096;
    73: op1_08_in15 = reg_0617;
    69: op1_08_in15 = reg_0126;
    50: op1_08_in15 = reg_0922;
    54: op1_08_in15 = imem02_in[11:8];
    74: op1_08_in15 = reg_0435;
    68: op1_08_in15 = reg_1082;
    71: op1_08_in15 = reg_0203;
    81: op1_08_in15 = reg_0203;
    75: op1_08_in15 = reg_0431;
    61: op1_08_in15 = imem00_in[3:0];
    56: op1_08_in15 = reg_0006;
    87: op1_08_in15 = imem03_in[15:12];
    76: op1_08_in15 = reg_0351;
    102: op1_08_in15 = reg_0351;
    57: op1_08_in15 = reg_0169;
    77: op1_08_in15 = reg_0188;
    58: op1_08_in15 = reg_0133;
    78: op1_08_in15 = reg_1439;
    70: op1_08_in15 = reg_0008;
    51: op1_08_in15 = reg_0100;
    88: op1_08_in15 = reg_0535;
    46: op1_08_in15 = reg_0281;
    59: op1_08_in15 = reg_0319;
    79: op1_08_in15 = reg_0585;
    60: op1_08_in15 = reg_0412;
    80: op1_08_in15 = reg_0058;
    114: op1_08_in15 = reg_0058;
    62: op1_08_in15 = reg_0460;
    48: op1_08_in15 = reg_0540;
    52: op1_08_in15 = reg_0397;
    63: op1_08_in15 = reg_0342;
    99: op1_08_in15 = reg_0342;
    82: op1_08_in15 = reg_0974;
    89: op1_08_in15 = reg_0500;
    117: op1_08_in15 = reg_0500;
    83: op1_08_in15 = reg_0405;
    64: op1_08_in15 = reg_0602;
    101: op1_08_in15 = reg_0602;
    84: op1_08_in15 = reg_1426;
    65: op1_08_in15 = reg_0898;
    85: op1_08_in15 = reg_0389;
    90: op1_08_in15 = reg_0701;
    66: op1_08_in15 = reg_0432;
    91: op1_08_in15 = reg_0333;
    67: op1_08_in15 = reg_0932;
    92: op1_08_in15 = reg_0931;
    93: op1_08_in15 = reg_0189;
    94: op1_08_in15 = reg_0053;
    95: op1_08_in15 = reg_1258;
    98: op1_08_in15 = reg_0121;
    44: op1_08_in15 = reg_0449;
    100: op1_08_in15 = reg_0228;
    47: op1_08_in15 = reg_0825;
    40: op1_08_in15 = reg_0236;
    103: op1_08_in15 = reg_0800;
    104: op1_08_in15 = imem04_in[3:0];
    105: op1_08_in15 = reg_0964;
    106: op1_08_in15 = reg_0001;
    107: op1_08_in15 = reg_0015;
    108: op1_08_in15 = reg_0934;
    109: op1_08_in15 = reg_0495;
    110: op1_08_in15 = reg_0867;
    111: op1_08_in15 = reg_0380;
    112: op1_08_in15 = reg_0939;
    113: op1_08_in15 = reg_0631;
    115: op1_08_in15 = reg_1092;
    116: op1_08_in15 = reg_1326;
    118: op1_08_in15 = reg_0031;
    119: op1_08_in15 = reg_0115;
    120: op1_08_in15 = reg_0427;
    121: op1_08_in15 = reg_0576;
    122: op1_08_in15 = reg_0409;
    123: op1_08_in15 = reg_0903;
    124: op1_08_in15 = reg_1473;
    125: op1_08_in15 = reg_0192;
    126: op1_08_in15 = reg_0071;
    127: op1_08_in15 = reg_0309;
    42: op1_08_in15 = reg_0382;
    128: op1_08_in15 = reg_0109;
    129: op1_08_in15 = reg_0975;
    130: op1_08_in15 = reg_0650;
    131: op1_08_in15 = reg_0242;
    default: op1_08_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_08_inv15 = 1;
    86: op1_08_inv15 = 1;
    73: op1_08_inv15 = 1;
    69: op1_08_inv15 = 1;
    54: op1_08_inv15 = 1;
    75: op1_08_inv15 = 1;
    61: op1_08_inv15 = 1;
    56: op1_08_inv15 = 1;
    87: op1_08_inv15 = 1;
    57: op1_08_inv15 = 1;
    70: op1_08_inv15 = 1;
    88: op1_08_inv15 = 1;
    79: op1_08_inv15 = 1;
    80: op1_08_inv15 = 1;
    63: op1_08_inv15 = 1;
    83: op1_08_inv15 = 1;
    64: op1_08_inv15 = 1;
    65: op1_08_inv15 = 1;
    66: op1_08_inv15 = 1;
    67: op1_08_inv15 = 1;
    93: op1_08_inv15 = 1;
    47: op1_08_inv15 = 1;
    40: op1_08_inv15 = 1;
    104: op1_08_inv15 = 1;
    105: op1_08_inv15 = 1;
    108: op1_08_inv15 = 1;
    109: op1_08_inv15 = 1;
    111: op1_08_inv15 = 1;
    112: op1_08_inv15 = 1;
    114: op1_08_inv15 = 1;
    115: op1_08_inv15 = 1;
    117: op1_08_inv15 = 1;
    120: op1_08_inv15 = 1;
    121: op1_08_inv15 = 1;
    123: op1_08_inv15 = 1;
    125: op1_08_inv15 = 1;
    126: op1_08_inv15 = 1;
    127: op1_08_inv15 = 1;
    42: op1_08_inv15 = 1;
    129: op1_08_inv15 = 1;
    130: op1_08_inv15 = 1;
    131: op1_08_inv15 = 1;
    default: op1_08_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in16 = reg_0289;
    53: op1_08_in16 = reg_0455;
    55: op1_08_in16 = reg_0489;
    86: op1_08_in16 = reg_0211;
    73: op1_08_in16 = reg_1228;
    69: op1_08_in16 = reg_0105;
    50: op1_08_in16 = reg_0976;
    54: op1_08_in16 = reg_0629;
    74: op1_08_in16 = reg_0134;
    83: op1_08_in16 = reg_0134;
    68: op1_08_in16 = reg_0421;
    71: op1_08_in16 = reg_1321;
    75: op1_08_in16 = reg_1322;
    61: op1_08_in16 = imem01_in[3:0];
    56: op1_08_in16 = reg_0311;
    87: op1_08_in16 = reg_0425;
    76: op1_08_in16 = reg_0428;
    57: op1_08_in16 = reg_0777;
    77: op1_08_in16 = reg_0722;
    58: op1_08_in16 = reg_0606;
    78: op1_08_in16 = reg_1440;
    70: op1_08_in16 = reg_1392;
    51: op1_08_in16 = reg_0321;
    88: op1_08_in16 = reg_0088;
    46: op1_08_in16 = reg_0313;
    59: op1_08_in16 = reg_0835;
    79: op1_08_in16 = reg_0584;
    60: op1_08_in16 = reg_0320;
    80: op1_08_in16 = reg_0917;
    62: op1_08_in16 = reg_0492;
    48: op1_08_in16 = reg_0167;
    52: op1_08_in16 = reg_0109;
    81: op1_08_in16 = reg_1254;
    63: op1_08_in16 = reg_0904;
    82: op1_08_in16 = reg_0133;
    89: op1_08_in16 = reg_1147;
    64: op1_08_in16 = reg_0449;
    84: op1_08_in16 = reg_1209;
    125: op1_08_in16 = reg_1209;
    65: op1_08_in16 = reg_0306;
    85: op1_08_in16 = reg_0059;
    90: op1_08_in16 = reg_0182;
    66: op1_08_in16 = reg_0973;
    91: op1_08_in16 = reg_1168;
    67: op1_08_in16 = reg_0199;
    92: op1_08_in16 = reg_0977;
    93: op1_08_in16 = reg_0440;
    94: op1_08_in16 = reg_0085;
    95: op1_08_in16 = reg_0462;
    98: op1_08_in16 = reg_0185;
    99: op1_08_in16 = reg_0698;
    44: op1_08_in16 = reg_0780;
    100: op1_08_in16 = reg_0087;
    106: op1_08_in16 = reg_0087;
    47: op1_08_in16 = reg_0717;
    101: op1_08_in16 = reg_0317;
    40: op1_08_in16 = reg_0150;
    102: op1_08_in16 = reg_0189;
    103: op1_08_in16 = reg_0294;
    104: op1_08_in16 = imem04_in[11:8];
    105: op1_08_in16 = reg_0954;
    107: op1_08_in16 = reg_0018;
    108: op1_08_in16 = reg_0839;
    109: op1_08_in16 = reg_0494;
    110: op1_08_in16 = reg_0893;
    111: op1_08_in16 = reg_0801;
    112: op1_08_in16 = reg_0938;
    113: op1_08_in16 = reg_0878;
    114: op1_08_in16 = reg_0026;
    115: op1_08_in16 = reg_0107;
    116: op1_08_in16 = reg_0860;
    117: op1_08_in16 = reg_0407;
    118: op1_08_in16 = reg_0030;
    119: op1_08_in16 = reg_1225;
    120: op1_08_in16 = reg_0264;
    121: op1_08_in16 = reg_0902;
    122: op1_08_in16 = reg_0389;
    123: op1_08_in16 = reg_1006;
    124: op1_08_in16 = reg_0430;
    126: op1_08_in16 = reg_0075;
    127: op1_08_in16 = reg_1094;
    42: op1_08_in16 = reg_0712;
    129: op1_08_in16 = reg_0712;
    128: op1_08_in16 = reg_0718;
    130: op1_08_in16 = reg_0579;
    131: op1_08_in16 = reg_0239;
    default: op1_08_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_08_inv16 = 1;
    55: op1_08_inv16 = 1;
    73: op1_08_inv16 = 1;
    69: op1_08_inv16 = 1;
    50: op1_08_inv16 = 1;
    74: op1_08_inv16 = 1;
    68: op1_08_inv16 = 1;
    61: op1_08_inv16 = 1;
    87: op1_08_inv16 = 1;
    76: op1_08_inv16 = 1;
    57: op1_08_inv16 = 1;
    58: op1_08_inv16 = 1;
    51: op1_08_inv16 = 1;
    46: op1_08_inv16 = 1;
    79: op1_08_inv16 = 1;
    52: op1_08_inv16 = 1;
    84: op1_08_inv16 = 1;
    65: op1_08_inv16 = 1;
    94: op1_08_inv16 = 1;
    99: op1_08_inv16 = 1;
    44: op1_08_inv16 = 1;
    100: op1_08_inv16 = 1;
    101: op1_08_inv16 = 1;
    40: op1_08_inv16 = 1;
    102: op1_08_inv16 = 1;
    105: op1_08_inv16 = 1;
    106: op1_08_inv16 = 1;
    108: op1_08_inv16 = 1;
    113: op1_08_inv16 = 1;
    115: op1_08_inv16 = 1;
    119: op1_08_inv16 = 1;
    120: op1_08_inv16 = 1;
    121: op1_08_inv16 = 1;
    122: op1_08_inv16 = 1;
    124: op1_08_inv16 = 1;
    126: op1_08_inv16 = 1;
    127: op1_08_inv16 = 1;
    128: op1_08_inv16 = 1;
    131: op1_08_inv16 = 1;
    default: op1_08_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in17 = reg_0119;
    53: op1_08_in17 = reg_0531;
    95: op1_08_in17 = reg_0531;
    55: op1_08_in17 = reg_0791;
    86: op1_08_in17 = reg_0205;
    73: op1_08_in17 = reg_0171;
    69: op1_08_in17 = reg_0708;
    50: op1_08_in17 = reg_0455;
    54: op1_08_in17 = reg_0133;
    74: op1_08_in17 = reg_0387;
    68: op1_08_in17 = reg_0412;
    71: op1_08_in17 = reg_1322;
    75: op1_08_in17 = reg_0027;
    61: op1_08_in17 = imem01_in[11:8];
    56: op1_08_in17 = reg_0312;
    87: op1_08_in17 = reg_0411;
    76: op1_08_in17 = reg_0435;
    93: op1_08_in17 = reg_0435;
    57: op1_08_in17 = reg_0775;
    77: op1_08_in17 = reg_0410;
    58: op1_08_in17 = reg_0605;
    78: op1_08_in17 = reg_0491;
    70: op1_08_in17 = reg_0820;
    51: op1_08_in17 = reg_0086;
    88: op1_08_in17 = reg_0252;
    46: op1_08_in17 = reg_0755;
    59: op1_08_in17 = reg_0337;
    63: op1_08_in17 = reg_0337;
    79: op1_08_in17 = reg_0529;
    60: op1_08_in17 = reg_0341;
    80: op1_08_in17 = reg_1071;
    62: op1_08_in17 = reg_0928;
    48: op1_08_in17 = reg_0450;
    90: op1_08_in17 = reg_0450;
    52: op1_08_in17 = reg_0714;
    81: op1_08_in17 = reg_0222;
    82: op1_08_in17 = reg_1334;
    89: op1_08_in17 = reg_0199;
    83: op1_08_in17 = reg_1290;
    64: op1_08_in17 = reg_1035;
    84: op1_08_in17 = reg_0730;
    92: op1_08_in17 = reg_0730;
    125: op1_08_in17 = reg_0730;
    65: op1_08_in17 = reg_0878;
    85: op1_08_in17 = reg_0464;
    66: op1_08_in17 = reg_0972;
    91: op1_08_in17 = reg_1169;
    67: op1_08_in17 = reg_0262;
    94: op1_08_in17 = reg_0484;
    98: op1_08_in17 = reg_0573;
    99: op1_08_in17 = reg_1143;
    44: op1_08_in17 = reg_0373;
    100: op1_08_in17 = reg_0520;
    47: op1_08_in17 = reg_0524;
    101: op1_08_in17 = reg_0039;
    40: op1_08_in17 = reg_0035;
    102: op1_08_in17 = reg_0409;
    103: op1_08_in17 = reg_1078;
    104: op1_08_in17 = reg_1144;
    105: op1_08_in17 = reg_1149;
    107: op1_08_in17 = reg_1060;
    108: op1_08_in17 = reg_0744;
    109: op1_08_in17 = reg_0054;
    110: op1_08_in17 = reg_0324;
    111: op1_08_in17 = reg_0294;
    112: op1_08_in17 = reg_0794;
    113: op1_08_in17 = reg_1492;
    114: op1_08_in17 = reg_0282;
    115: op1_08_in17 = reg_0707;
    116: op1_08_in17 = reg_1323;
    117: op1_08_in17 = reg_0452;
    118: op1_08_in17 = reg_0286;
    119: op1_08_in17 = reg_0132;
    120: op1_08_in17 = reg_1203;
    121: op1_08_in17 = reg_0163;
    122: op1_08_in17 = reg_0075;
    123: op1_08_in17 = reg_0217;
    124: op1_08_in17 = reg_0726;
    126: op1_08_in17 = reg_0072;
    127: op1_08_in17 = reg_0661;
    42: op1_08_in17 = reg_0846;
    128: op1_08_in17 = reg_1303;
    129: op1_08_in17 = reg_0839;
    130: op1_08_in17 = reg_0832;
    131: op1_08_in17 = reg_0553;
    default: op1_08_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_08_inv17 = 1;
    86: op1_08_inv17 = 1;
    69: op1_08_inv17 = 1;
    50: op1_08_inv17 = 1;
    54: op1_08_inv17 = 1;
    74: op1_08_inv17 = 1;
    71: op1_08_inv17 = 1;
    75: op1_08_inv17 = 1;
    61: op1_08_inv17 = 1;
    56: op1_08_inv17 = 1;
    87: op1_08_inv17 = 1;
    57: op1_08_inv17 = 1;
    77: op1_08_inv17 = 1;
    78: op1_08_inv17 = 1;
    51: op1_08_inv17 = 1;
    88: op1_08_inv17 = 1;
    60: op1_08_inv17 = 1;
    80: op1_08_inv17 = 1;
    83: op1_08_inv17 = 1;
    64: op1_08_inv17 = 1;
    85: op1_08_inv17 = 1;
    90: op1_08_inv17 = 1;
    94: op1_08_inv17 = 1;
    44: op1_08_inv17 = 1;
    100: op1_08_inv17 = 1;
    102: op1_08_inv17 = 1;
    104: op1_08_inv17 = 1;
    109: op1_08_inv17 = 1;
    115: op1_08_inv17 = 1;
    116: op1_08_inv17 = 1;
    117: op1_08_inv17 = 1;
    119: op1_08_inv17 = 1;
    120: op1_08_inv17 = 1;
    121: op1_08_inv17 = 1;
    122: op1_08_inv17 = 1;
    124: op1_08_inv17 = 1;
    125: op1_08_inv17 = 1;
    126: op1_08_inv17 = 1;
    127: op1_08_inv17 = 1;
    131: op1_08_inv17 = 1;
    default: op1_08_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in18 = reg_0023;
    53: op1_08_in18 = imem02_in[11:8];
    55: op1_08_in18 = reg_0029;
    86: op1_08_in18 = reg_0578;
    73: op1_08_in18 = reg_0244;
    69: op1_08_in18 = reg_0705;
    50: op1_08_in18 = reg_0472;
    54: op1_08_in18 = reg_0606;
    74: op1_08_in18 = reg_0075;
    68: op1_08_in18 = reg_0936;
    71: op1_08_in18 = reg_0786;
    75: op1_08_in18 = reg_1068;
    61: op1_08_in18 = reg_0166;
    56: op1_08_in18 = reg_0755;
    87: op1_08_in18 = reg_1372;
    76: op1_08_in18 = reg_0405;
    77: op1_08_in18 = reg_0405;
    57: op1_08_in18 = reg_0465;
    58: op1_08_in18 = reg_0455;
    78: op1_08_in18 = reg_0461;
    70: op1_08_in18 = reg_1132;
    88: op1_08_in18 = reg_1338;
    46: op1_08_in18 = reg_0227;
    111: op1_08_in18 = reg_0227;
    59: op1_08_in18 = reg_0164;
    79: op1_08_in18 = reg_0672;
    60: op1_08_in18 = reg_0487;
    67: op1_08_in18 = reg_0487;
    80: op1_08_in18 = reg_1253;
    62: op1_08_in18 = reg_0883;
    48: op1_08_in18 = reg_0418;
    52: op1_08_in18 = reg_0671;
    81: op1_08_in18 = reg_1474;
    63: op1_08_in18 = reg_0097;
    82: op1_08_in18 = reg_0860;
    89: op1_08_in18 = reg_1077;
    83: op1_08_in18 = reg_0788;
    114: op1_08_in18 = reg_0788;
    64: op1_08_in18 = reg_0754;
    84: op1_08_in18 = reg_0752;
    116: op1_08_in18 = reg_0752;
    65: op1_08_in18 = reg_0839;
    85: op1_08_in18 = reg_1291;
    90: op1_08_in18 = reg_0118;
    66: op1_08_in18 = reg_0626;
    91: op1_08_in18 = reg_0831;
    92: op1_08_in18 = reg_0974;
    93: op1_08_in18 = reg_0134;
    95: op1_08_in18 = reg_0552;
    98: op1_08_in18 = reg_0823;
    99: op1_08_in18 = reg_0339;
    44: op1_08_in18 = reg_0115;
    47: op1_08_in18 = reg_0635;
    101: op1_08_in18 = reg_1058;
    40: op1_08_in18 = reg_0034;
    102: op1_08_in18 = reg_0410;
    103: op1_08_in18 = reg_0009;
    104: op1_08_in18 = reg_0467;
    105: op1_08_in18 = reg_0707;
    107: op1_08_in18 = reg_0667;
    108: op1_08_in18 = reg_0971;
    109: op1_08_in18 = reg_0127;
    110: op1_08_in18 = reg_1415;
    112: op1_08_in18 = reg_0197;
    113: op1_08_in18 = reg_0802;
    115: op1_08_in18 = reg_0541;
    117: op1_08_in18 = reg_1419;
    118: op1_08_in18 = reg_0321;
    119: op1_08_in18 = reg_0419;
    120: op1_08_in18 = reg_0796;
    121: op1_08_in18 = reg_0549;
    122: op1_08_in18 = reg_0723;
    123: op1_08_in18 = reg_0758;
    124: op1_08_in18 = reg_0147;
    125: op1_08_in18 = reg_1505;
    126: op1_08_in18 = reg_1324;
    127: op1_08_in18 = reg_0664;
    42: op1_08_in18 = reg_0217;
    128: op1_08_in18 = reg_0374;
    129: op1_08_in18 = reg_0744;
    130: op1_08_in18 = reg_0986;
    131: op1_08_in18 = reg_0013;
    default: op1_08_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv18 = 1;
    53: op1_08_inv18 = 1;
    86: op1_08_inv18 = 1;
    73: op1_08_inv18 = 1;
    69: op1_08_inv18 = 1;
    71: op1_08_inv18 = 1;
    75: op1_08_inv18 = 1;
    56: op1_08_inv18 = 1;
    70: op1_08_inv18 = 1;
    88: op1_08_inv18 = 1;
    46: op1_08_inv18 = 1;
    62: op1_08_inv18 = 1;
    52: op1_08_inv18 = 1;
    81: op1_08_inv18 = 1;
    63: op1_08_inv18 = 1;
    82: op1_08_inv18 = 1;
    64: op1_08_inv18 = 1;
    90: op1_08_inv18 = 1;
    66: op1_08_inv18 = 1;
    67: op1_08_inv18 = 1;
    92: op1_08_inv18 = 1;
    95: op1_08_inv18 = 1;
    99: op1_08_inv18 = 1;
    44: op1_08_inv18 = 1;
    47: op1_08_inv18 = 1;
    101: op1_08_inv18 = 1;
    40: op1_08_inv18 = 1;
    104: op1_08_inv18 = 1;
    105: op1_08_inv18 = 1;
    109: op1_08_inv18 = 1;
    114: op1_08_inv18 = 1;
    116: op1_08_inv18 = 1;
    117: op1_08_inv18 = 1;
    118: op1_08_inv18 = 1;
    119: op1_08_inv18 = 1;
    120: op1_08_inv18 = 1;
    125: op1_08_inv18 = 1;
    126: op1_08_inv18 = 1;
    129: op1_08_inv18 = 1;
    default: op1_08_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in19 = reg_0065;
    53: op1_08_in19 = imem02_in[15:12];
    55: op1_08_in19 = reg_0665;
    86: op1_08_in19 = reg_0733;
    73: op1_08_in19 = reg_0165;
    69: op1_08_in19 = reg_0306;
    50: op1_08_in19 = reg_0474;
    54: op1_08_in19 = reg_0532;
    129: op1_08_in19 = reg_0532;
    74: op1_08_in19 = reg_0122;
    68: op1_08_in19 = reg_0452;
    71: op1_08_in19 = reg_1069;
    75: op1_08_in19 = reg_1070;
    61: op1_08_in19 = reg_1291;
    56: op1_08_in19 = reg_0678;
    87: op1_08_in19 = reg_1368;
    76: op1_08_in19 = reg_0134;
    57: op1_08_in19 = reg_0030;
    77: op1_08_in19 = reg_0389;
    58: op1_08_in19 = reg_0589;
    78: op1_08_in19 = reg_0673;
    70: op1_08_in19 = reg_0677;
    88: op1_08_in19 = reg_0531;
    46: op1_08_in19 = reg_0710;
    111: op1_08_in19 = reg_0710;
    59: op1_08_in19 = reg_0021;
    79: op1_08_in19 = reg_0391;
    60: op1_08_in19 = reg_0337;
    80: op1_08_in19 = reg_0166;
    85: op1_08_in19 = reg_0166;
    62: op1_08_in19 = reg_0642;
    48: op1_08_in19 = reg_0890;
    130: op1_08_in19 = reg_0890;
    52: op1_08_in19 = reg_0247;
    81: op1_08_in19 = reg_0430;
    63: op1_08_in19 = reg_0181;
    82: op1_08_in19 = reg_0863;
    89: op1_08_in19 = reg_1065;
    83: op1_08_in19 = reg_0047;
    64: op1_08_in19 = reg_0195;
    84: op1_08_in19 = reg_1504;
    65: op1_08_in19 = imem02_in[3:0];
    90: op1_08_in19 = reg_0240;
    66: op1_08_in19 = reg_0106;
    91: op1_08_in19 = reg_0167;
    67: op1_08_in19 = reg_0251;
    92: op1_08_in19 = reg_0133;
    93: op1_08_in19 = reg_0071;
    95: op1_08_in19 = reg_1200;
    98: op1_08_in19 = reg_1494;
    99: op1_08_in19 = reg_0211;
    44: op1_08_in19 = reg_0634;
    47: op1_08_in19 = reg_0584;
    101: op1_08_in19 = reg_0795;
    40: op1_08_in19 = reg_0579;
    102: op1_08_in19 = reg_0073;
    103: op1_08_in19 = reg_0006;
    104: op1_08_in19 = reg_0208;
    105: op1_08_in19 = reg_0025;
    107: op1_08_in19 = reg_0922;
    108: op1_08_in19 = reg_0126;
    109: op1_08_in19 = reg_0897;
    110: op1_08_in19 = reg_0994;
    112: op1_08_in19 = reg_0275;
    113: op1_08_in19 = reg_0989;
    114: op1_08_in19 = reg_0463;
    115: op1_08_in19 = reg_0411;
    116: op1_08_in19 = reg_0116;
    117: op1_08_in19 = reg_1143;
    118: op1_08_in19 = reg_0361;
    119: op1_08_in19 = reg_0023;
    120: op1_08_in19 = reg_0471;
    121: op1_08_in19 = reg_0743;
    122: op1_08_in19 = reg_0966;
    123: op1_08_in19 = reg_0840;
    124: op1_08_in19 = reg_1034;
    125: op1_08_in19 = reg_0172;
    126: op1_08_in19 = reg_0917;
    127: op1_08_in19 = reg_0285;
    42: op1_08_in19 = reg_0325;
    128: op1_08_in19 = reg_0624;
    131: op1_08_in19 = reg_0747;
    default: op1_08_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv19 = 1;
    53: op1_08_inv19 = 1;
    55: op1_08_inv19 = 1;
    86: op1_08_inv19 = 1;
    73: op1_08_inv19 = 1;
    69: op1_08_inv19 = 1;
    50: op1_08_inv19 = 1;
    74: op1_08_inv19 = 1;
    68: op1_08_inv19 = 1;
    71: op1_08_inv19 = 1;
    61: op1_08_inv19 = 1;
    56: op1_08_inv19 = 1;
    76: op1_08_inv19 = 1;
    77: op1_08_inv19 = 1;
    70: op1_08_inv19 = 1;
    88: op1_08_inv19 = 1;
    46: op1_08_inv19 = 1;
    59: op1_08_inv19 = 1;
    60: op1_08_inv19 = 1;
    48: op1_08_inv19 = 1;
    63: op1_08_inv19 = 1;
    82: op1_08_inv19 = 1;
    83: op1_08_inv19 = 1;
    66: op1_08_inv19 = 1;
    67: op1_08_inv19 = 1;
    92: op1_08_inv19 = 1;
    93: op1_08_inv19 = 1;
    95: op1_08_inv19 = 1;
    98: op1_08_inv19 = 1;
    99: op1_08_inv19 = 1;
    40: op1_08_inv19 = 1;
    102: op1_08_inv19 = 1;
    103: op1_08_inv19 = 1;
    104: op1_08_inv19 = 1;
    108: op1_08_inv19 = 1;
    109: op1_08_inv19 = 1;
    110: op1_08_inv19 = 1;
    116: op1_08_inv19 = 1;
    118: op1_08_inv19 = 1;
    119: op1_08_inv19 = 1;
    120: op1_08_inv19 = 1;
    121: op1_08_inv19 = 1;
    123: op1_08_inv19 = 1;
    124: op1_08_inv19 = 1;
    126: op1_08_inv19 = 1;
    127: op1_08_inv19 = 1;
    128: op1_08_inv19 = 1;
    129: op1_08_inv19 = 1;
    131: op1_08_inv19 = 1;
    default: op1_08_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in20 = reg_0461;
    53: op1_08_in20 = reg_0496;
    55: op1_08_in20 = reg_0442;
    86: op1_08_in20 = reg_1169;
    73: op1_08_in20 = reg_1202;
    69: op1_08_in20 = reg_0009;
    50: op1_08_in20 = reg_0432;
    129: op1_08_in20 = reg_0432;
    54: op1_08_in20 = reg_1140;
    74: op1_08_in20 = reg_0027;
    68: op1_08_in20 = reg_0340;
    71: op1_08_in20 = reg_0259;
    75: op1_08_in20 = imem01_in[7:4];
    61: op1_08_in20 = reg_1068;
    56: op1_08_in20 = reg_0709;
    87: op1_08_in20 = reg_0535;
    76: op1_08_in20 = reg_0387;
    57: op1_08_in20 = reg_0663;
    77: op1_08_in20 = reg_0060;
    58: op1_08_in20 = reg_0532;
    78: op1_08_in20 = reg_0894;
    70: op1_08_in20 = reg_0710;
    88: op1_08_in20 = reg_1083;
    46: op1_08_in20 = reg_0375;
    59: op1_08_in20 = reg_0794;
    79: op1_08_in20 = reg_0162;
    60: op1_08_in20 = reg_0097;
    80: op1_08_in20 = reg_0553;
    83: op1_08_in20 = reg_0553;
    62: op1_08_in20 = reg_0640;
    48: op1_08_in20 = reg_0888;
    52: op1_08_in20 = reg_0568;
    81: op1_08_in20 = reg_0434;
    63: op1_08_in20 = reg_0065;
    82: op1_08_in20 = reg_0859;
    89: op1_08_in20 = reg_0582;
    64: op1_08_in20 = reg_0780;
    84: op1_08_in20 = reg_0372;
    65: op1_08_in20 = imem02_in[11:8];
    85: op1_08_in20 = reg_0746;
    90: op1_08_in20 = reg_0797;
    66: op1_08_in20 = reg_0105;
    91: op1_08_in20 = reg_1181;
    67: op1_08_in20 = reg_0833;
    92: op1_08_in20 = reg_0984;
    93: op1_08_in20 = reg_1324;
    95: op1_08_in20 = reg_0500;
    98: op1_08_in20 = reg_0952;
    99: op1_08_in20 = reg_0236;
    44: op1_08_in20 = reg_0637;
    47: op1_08_in20 = reg_0527;
    101: op1_08_in20 = reg_0974;
    40: op1_08_in20 = reg_0736;
    102: op1_08_in20 = reg_0058;
    103: op1_08_in20 = imem03_in[3:0];
    104: op1_08_in20 = reg_0493;
    105: op1_08_in20 = reg_1139;
    107: op1_08_in20 = reg_0139;
    108: op1_08_in20 = reg_0112;
    109: op1_08_in20 = reg_0695;
    110: op1_08_in20 = reg_1055;
    111: op1_08_in20 = reg_0185;
    112: op1_08_in20 = reg_0196;
    113: op1_08_in20 = reg_0732;
    114: op1_08_in20 = reg_0550;
    115: op1_08_in20 = reg_0032;
    116: op1_08_in20 = reg_0718;
    117: op1_08_in20 = reg_0117;
    118: op1_08_in20 = reg_0087;
    119: op1_08_in20 = reg_0015;
    120: op1_08_in20 = reg_0537;
    121: op1_08_in20 = reg_0820;
    122: op1_08_in20 = reg_0788;
    123: op1_08_in20 = reg_0479;
    124: op1_08_in20 = reg_0360;
    125: op1_08_in20 = reg_1179;
    126: op1_08_in20 = reg_0723;
    127: op1_08_in20 = reg_0228;
    42: op1_08_in20 = reg_0314;
    128: op1_08_in20 = reg_0152;
    130: op1_08_in20 = reg_1268;
    131: op1_08_in20 = reg_0610;
    default: op1_08_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_08_inv20 = 1;
    74: op1_08_inv20 = 1;
    61: op1_08_inv20 = 1;
    87: op1_08_inv20 = 1;
    76: op1_08_inv20 = 1;
    58: op1_08_inv20 = 1;
    88: op1_08_inv20 = 1;
    59: op1_08_inv20 = 1;
    79: op1_08_inv20 = 1;
    60: op1_08_inv20 = 1;
    80: op1_08_inv20 = 1;
    48: op1_08_inv20 = 1;
    63: op1_08_inv20 = 1;
    83: op1_08_inv20 = 1;
    85: op1_08_inv20 = 1;
    66: op1_08_inv20 = 1;
    67: op1_08_inv20 = 1;
    93: op1_08_inv20 = 1;
    95: op1_08_inv20 = 1;
    98: op1_08_inv20 = 1;
    99: op1_08_inv20 = 1;
    44: op1_08_inv20 = 1;
    102: op1_08_inv20 = 1;
    104: op1_08_inv20 = 1;
    108: op1_08_inv20 = 1;
    109: op1_08_inv20 = 1;
    110: op1_08_inv20 = 1;
    111: op1_08_inv20 = 1;
    112: op1_08_inv20 = 1;
    113: op1_08_inv20 = 1;
    115: op1_08_inv20 = 1;
    117: op1_08_inv20 = 1;
    120: op1_08_inv20 = 1;
    121: op1_08_inv20 = 1;
    124: op1_08_inv20 = 1;
    127: op1_08_inv20 = 1;
    128: op1_08_inv20 = 1;
    129: op1_08_inv20 = 1;
    130: op1_08_inv20 = 1;
    131: op1_08_inv20 = 1;
    default: op1_08_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in21 = reg_1416;
    53: op1_08_in21 = reg_0494;
    55: op1_08_in21 = reg_0739;
    86: op1_08_in21 = reg_0392;
    73: op1_08_in21 = reg_0152;
    69: op1_08_in21 = reg_0379;
    50: op1_08_in21 = reg_0054;
    54: op1_08_in21 = reg_1139;
    74: op1_08_in21 = reg_0785;
    68: op1_08_in21 = reg_0305;
    71: op1_08_in21 = reg_0547;
    80: op1_08_in21 = reg_0547;
    75: op1_08_in21 = imem01_in[15:12];
    61: op1_08_in21 = reg_1031;
    56: op1_08_in21 = reg_1064;
    87: op1_08_in21 = reg_0088;
    104: op1_08_in21 = reg_0088;
    76: op1_08_in21 = reg_1324;
    57: op1_08_in21 = reg_0442;
    77: op1_08_in21 = reg_1100;
    58: op1_08_in21 = imem02_in[15:12];
    78: op1_08_in21 = reg_0135;
    70: op1_08_in21 = reg_0375;
    88: op1_08_in21 = reg_1200;
    46: op1_08_in21 = reg_0234;
    59: op1_08_in21 = reg_0331;
    79: op1_08_in21 = reg_0667;
    60: op1_08_in21 = reg_0164;
    62: op1_08_in21 = reg_0189;
    48: op1_08_in21 = reg_0303;
    52: op1_08_in21 = reg_0569;
    81: op1_08_in21 = reg_0438;
    63: op1_08_in21 = reg_0062;
    82: op1_08_in21 = reg_1323;
    89: op1_08_in21 = reg_0337;
    83: op1_08_in21 = reg_0242;
    85: op1_08_in21 = reg_0242;
    64: op1_08_in21 = reg_1105;
    84: op1_08_in21 = reg_0116;
    65: op1_08_in21 = reg_0069;
    90: op1_08_in21 = reg_0864;
    66: op1_08_in21 = reg_0876;
    91: op1_08_in21 = reg_1401;
    67: op1_08_in21 = reg_1164;
    92: op1_08_in21 = reg_0860;
    93: op1_08_in21 = reg_0089;
    95: op1_08_in21 = reg_0412;
    98: op1_08_in21 = reg_0190;
    99: op1_08_in21 = reg_0420;
    44: op1_08_in21 = reg_0624;
    47: op1_08_in21 = reg_0295;
    101: op1_08_in21 = reg_1467;
    40: op1_08_in21 = imem05_in[15:12];
    102: op1_08_in21 = reg_0027;
    103: op1_08_in21 = imem03_in[7:4];
    105: op1_08_in21 = reg_1340;
    107: op1_08_in21 = reg_0030;
    108: op1_08_in21 = reg_1433;
    109: op1_08_in21 = reg_1078;
    110: op1_08_in21 = reg_1056;
    111: op1_08_in21 = reg_0706;
    112: op1_08_in21 = reg_0243;
    113: op1_08_in21 = reg_0597;
    114: op1_08_in21 = reg_1473;
    115: op1_08_in21 = reg_0534;
    116: op1_08_in21 = reg_0636;
    117: op1_08_in21 = reg_0019;
    118: op1_08_in21 = reg_0124;
    119: op1_08_in21 = reg_1097;
    120: op1_08_in21 = reg_1004;
    121: op1_08_in21 = reg_0967;
    122: op1_08_in21 = reg_0183;
    123: op1_08_in21 = reg_1063;
    124: op1_08_in21 = reg_0899;
    125: op1_08_in21 = reg_0265;
    126: op1_08_in21 = reg_0788;
    127: op1_08_in21 = reg_0085;
    42: op1_08_in21 = reg_0755;
    128: op1_08_in21 = reg_0215;
    129: op1_08_in21 = reg_0776;
    130: op1_08_in21 = reg_1059;
    131: op1_08_in21 = reg_0572;
    default: op1_08_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_08_inv21 = 1;
    50: op1_08_inv21 = 1;
    54: op1_08_inv21 = 1;
    74: op1_08_inv21 = 1;
    61: op1_08_inv21 = 1;
    56: op1_08_inv21 = 1;
    57: op1_08_inv21 = 1;
    77: op1_08_inv21 = 1;
    70: op1_08_inv21 = 1;
    88: op1_08_inv21 = 1;
    59: op1_08_inv21 = 1;
    60: op1_08_inv21 = 1;
    80: op1_08_inv21 = 1;
    62: op1_08_inv21 = 1;
    81: op1_08_inv21 = 1;
    63: op1_08_inv21 = 1;
    82: op1_08_inv21 = 1;
    89: op1_08_inv21 = 1;
    83: op1_08_inv21 = 1;
    65: op1_08_inv21 = 1;
    85: op1_08_inv21 = 1;
    66: op1_08_inv21 = 1;
    91: op1_08_inv21 = 1;
    92: op1_08_inv21 = 1;
    93: op1_08_inv21 = 1;
    95: op1_08_inv21 = 1;
    44: op1_08_inv21 = 1;
    47: op1_08_inv21 = 1;
    101: op1_08_inv21 = 1;
    102: op1_08_inv21 = 1;
    103: op1_08_inv21 = 1;
    104: op1_08_inv21 = 1;
    110: op1_08_inv21 = 1;
    111: op1_08_inv21 = 1;
    112: op1_08_inv21 = 1;
    113: op1_08_inv21 = 1;
    114: op1_08_inv21 = 1;
    115: op1_08_inv21 = 1;
    117: op1_08_inv21 = 1;
    118: op1_08_inv21 = 1;
    120: op1_08_inv21 = 1;
    121: op1_08_inv21 = 1;
    123: op1_08_inv21 = 1;
    124: op1_08_inv21 = 1;
    125: op1_08_inv21 = 1;
    42: op1_08_inv21 = 1;
    128: op1_08_inv21 = 1;
    129: op1_08_inv21 = 1;
    131: op1_08_inv21 = 1;
    default: op1_08_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in22 = reg_1415;
    53: op1_08_in22 = reg_0474;
    55: op1_08_in22 = reg_0137;
    86: op1_08_in22 = reg_0491;
    73: op1_08_in22 = reg_0213;
    69: op1_08_in22 = reg_0217;
    50: op1_08_in22 = reg_0379;
    54: op1_08_in22 = reg_0128;
    74: op1_08_in22 = reg_0175;
    68: op1_08_in22 = reg_0487;
    71: op1_08_in22 = reg_0868;
    75: op1_08_in22 = reg_0930;
    61: op1_08_in22 = reg_0819;
    121: op1_08_in22 = reg_0819;
    56: op1_08_in22 = reg_0377;
    87: op1_08_in22 = reg_1339;
    76: op1_08_in22 = reg_0122;
    57: op1_08_in22 = reg_0408;
    77: op1_08_in22 = reg_0372;
    58: op1_08_in22 = reg_0475;
    78: op1_08_in22 = reg_0674;
    70: op1_08_in22 = reg_0789;
    88: op1_08_in22 = reg_0488;
    46: op1_08_in22 = reg_0349;
    59: op1_08_in22 = reg_0750;
    79: op1_08_in22 = reg_0309;
    60: op1_08_in22 = reg_0117;
    80: op1_08_in22 = reg_0549;
    62: op1_08_in22 = reg_0440;
    48: op1_08_in22 = reg_0873;
    52: op1_08_in22 = reg_0528;
    81: op1_08_in22 = reg_1452;
    63: op1_08_in22 = reg_0021;
    99: op1_08_in22 = reg_0021;
    82: op1_08_in22 = reg_0780;
    89: op1_08_in22 = reg_1151;
    83: op1_08_in22 = reg_0239;
    64: op1_08_in22 = reg_0906;
    84: op1_08_in22 = reg_0714;
    65: op1_08_in22 = reg_0325;
    85: op1_08_in22 = reg_0742;
    90: op1_08_in22 = imem06_in[3:0];
    66: op1_08_in22 = reg_0878;
    91: op1_08_in22 = reg_0450;
    67: op1_08_in22 = reg_0538;
    92: op1_08_in22 = reg_0720;
    93: op1_08_in22 = reg_0723;
    95: op1_08_in22 = reg_1041;
    98: op1_08_in22 = reg_0597;
    44: op1_08_in22 = reg_0527;
    47: op1_08_in22 = reg_0419;
    101: op1_08_in22 = reg_0751;
    40: op1_08_in22 = reg_0173;
    102: op1_08_in22 = reg_0183;
    103: op1_08_in22 = imem03_in[11:8];
    104: op1_08_in22 = reg_0797;
    105: op1_08_in22 = reg_0264;
    107: op1_08_in22 = reg_0738;
    108: op1_08_in22 = reg_1492;
    109: op1_08_in22 = reg_1091;
    110: op1_08_in22 = reg_0157;
    111: op1_08_in22 = reg_0999;
    112: op1_08_in22 = reg_0206;
    113: op1_08_in22 = reg_0220;
    114: op1_08_in22 = reg_0612;
    115: op1_08_in22 = reg_0181;
    116: op1_08_in22 = reg_0622;
    117: op1_08_in22 = reg_0540;
    119: op1_08_in22 = reg_1096;
    120: op1_08_in22 = reg_0452;
    122: op1_08_in22 = reg_1152;
    123: op1_08_in22 = reg_0216;
    124: op1_08_in22 = reg_0875;
    125: op1_08_in22 = reg_0110;
    126: op1_08_in22 = reg_0577;
    127: op1_08_in22 = reg_0226;
    42: op1_08_in22 = reg_0734;
    128: op1_08_in22 = reg_0017;
    129: op1_08_in22 = reg_0127;
    130: op1_08_in22 = reg_0340;
    131: op1_08_in22 = reg_0439;
    default: op1_08_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv22 = 1;
    69: op1_08_inv22 = 1;
    50: op1_08_inv22 = 1;
    54: op1_08_inv22 = 1;
    74: op1_08_inv22 = 1;
    56: op1_08_inv22 = 1;
    76: op1_08_inv22 = 1;
    77: op1_08_inv22 = 1;
    58: op1_08_inv22 = 1;
    70: op1_08_inv22 = 1;
    88: op1_08_inv22 = 1;
    46: op1_08_inv22 = 1;
    59: op1_08_inv22 = 1;
    81: op1_08_inv22 = 1;
    82: op1_08_inv22 = 1;
    89: op1_08_inv22 = 1;
    83: op1_08_inv22 = 1;
    65: op1_08_inv22 = 1;
    90: op1_08_inv22 = 1;
    91: op1_08_inv22 = 1;
    92: op1_08_inv22 = 1;
    95: op1_08_inv22 = 1;
    98: op1_08_inv22 = 1;
    47: op1_08_inv22 = 1;
    40: op1_08_inv22 = 1;
    103: op1_08_inv22 = 1;
    104: op1_08_inv22 = 1;
    105: op1_08_inv22 = 1;
    108: op1_08_inv22 = 1;
    110: op1_08_inv22 = 1;
    112: op1_08_inv22 = 1;
    113: op1_08_inv22 = 1;
    114: op1_08_inv22 = 1;
    116: op1_08_inv22 = 1;
    117: op1_08_inv22 = 1;
    119: op1_08_inv22 = 1;
    120: op1_08_inv22 = 1;
    121: op1_08_inv22 = 1;
    126: op1_08_inv22 = 1;
    42: op1_08_inv22 = 1;
    128: op1_08_inv22 = 1;
    default: op1_08_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in23 = reg_0703;
    53: op1_08_in23 = reg_0990;
    55: op1_08_in23 = reg_0103;
    86: op1_08_in23 = reg_0182;
    73: op1_08_in23 = reg_0015;
    69: op1_08_in23 = reg_0325;
    50: op1_08_in23 = reg_0154;
    54: op1_08_in23 = reg_0105;
    74: op1_08_in23 = reg_1032;
    102: op1_08_in23 = reg_1032;
    68: op1_08_in23 = reg_0862;
    71: op1_08_in23 = reg_0966;
    114: op1_08_in23 = reg_0966;
    75: op1_08_in23 = reg_0093;
    61: op1_08_in23 = reg_0434;
    56: op1_08_in23 = reg_0314;
    87: op1_08_in23 = reg_0252;
    76: op1_08_in23 = reg_0785;
    57: op1_08_in23 = reg_0415;
    77: op1_08_in23 = reg_0611;
    58: op1_08_in23 = reg_1207;
    78: op1_08_in23 = reg_0187;
    70: op1_08_in23 = reg_0999;
    88: op1_08_in23 = reg_1233;
    46: op1_08_in23 = reg_0179;
    59: op1_08_in23 = reg_0733;
    79: op1_08_in23 = reg_0139;
    60: op1_08_in23 = imem05_in[11:8];
    80: op1_08_in23 = reg_0548;
    62: op1_08_in23 = reg_0409;
    48: op1_08_in23 = reg_0861;
    52: op1_08_in23 = reg_0522;
    81: op1_08_in23 = reg_0360;
    63: op1_08_in23 = reg_0273;
    82: op1_08_in23 = reg_0115;
    89: op1_08_in23 = reg_0420;
    83: op1_08_in23 = reg_0238;
    64: op1_08_in23 = reg_0696;
    84: op1_08_in23 = reg_0636;
    65: op1_08_in23 = reg_0525;
    85: op1_08_in23 = reg_0968;
    90: op1_08_in23 = imem06_in[15:12];
    112: op1_08_in23 = imem06_in[15:12];
    66: op1_08_in23 = reg_0845;
    91: op1_08_in23 = reg_1514;
    67: op1_08_in23 = reg_0167;
    92: op1_08_in23 = reg_0869;
    93: op1_08_in23 = imem01_in[3:0];
    95: op1_08_in23 = reg_1077;
    98: op1_08_in23 = reg_1226;
    99: op1_08_in23 = reg_0020;
    44: op1_08_in23 = reg_0459;
    47: op1_08_in23 = reg_0461;
    101: op1_08_in23 = reg_0718;
    125: op1_08_in23 = reg_0718;
    40: op1_08_in23 = reg_0648;
    103: op1_08_in23 = reg_0328;
    104: op1_08_in23 = reg_0462;
    105: op1_08_in23 = reg_0094;
    107: op1_08_in23 = reg_0413;
    108: op1_08_in23 = reg_0632;
    109: op1_08_in23 = reg_0068;
    110: op1_08_in23 = reg_0223;
    111: op1_08_in23 = reg_0823;
    113: op1_08_in23 = reg_0261;
    115: op1_08_in23 = reg_1369;
    116: op1_08_in23 = reg_0624;
    117: op1_08_in23 = reg_0038;
    119: op1_08_in23 = reg_1183;
    120: op1_08_in23 = reg_0487;
    121: op1_08_in23 = reg_0439;
    122: op1_08_in23 = reg_0401;
    123: op1_08_in23 = reg_0847;
    124: op1_08_in23 = reg_0335;
    126: op1_08_in23 = reg_0985;
    42: op1_08_in23 = reg_0216;
    128: op1_08_in23 = reg_1170;
    129: op1_08_in23 = reg_0106;
    130: op1_08_in23 = reg_0562;
    131: op1_08_in23 = reg_1457;
    default: op1_08_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    50: op1_08_inv23 = 1;
    54: op1_08_inv23 = 1;
    75: op1_08_inv23 = 1;
    56: op1_08_inv23 = 1;
    76: op1_08_inv23 = 1;
    58: op1_08_inv23 = 1;
    46: op1_08_inv23 = 1;
    59: op1_08_inv23 = 1;
    79: op1_08_inv23 = 1;
    60: op1_08_inv23 = 1;
    80: op1_08_inv23 = 1;
    62: op1_08_inv23 = 1;
    63: op1_08_inv23 = 1;
    64: op1_08_inv23 = 1;
    85: op1_08_inv23 = 1;
    90: op1_08_inv23 = 1;
    66: op1_08_inv23 = 1;
    91: op1_08_inv23 = 1;
    67: op1_08_inv23 = 1;
    92: op1_08_inv23 = 1;
    98: op1_08_inv23 = 1;
    44: op1_08_inv23 = 1;
    101: op1_08_inv23 = 1;
    40: op1_08_inv23 = 1;
    102: op1_08_inv23 = 1;
    103: op1_08_inv23 = 1;
    105: op1_08_inv23 = 1;
    108: op1_08_inv23 = 1;
    109: op1_08_inv23 = 1;
    110: op1_08_inv23 = 1;
    114: op1_08_inv23 = 1;
    116: op1_08_inv23 = 1;
    117: op1_08_inv23 = 1;
    122: op1_08_inv23 = 1;
    125: op1_08_inv23 = 1;
    129: op1_08_inv23 = 1;
    130: op1_08_inv23 = 1;
    131: op1_08_inv23 = 1;
    default: op1_08_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in24 = reg_0297;
    53: op1_08_in24 = reg_0436;
    55: op1_08_in24 = reg_0228;
    86: op1_08_in24 = reg_0630;
    73: op1_08_in24 = reg_0065;
    69: op1_08_in24 = reg_0280;
    50: op1_08_in24 = reg_0325;
    54: op1_08_in24 = reg_0138;
    74: op1_08_in24 = reg_0047;
    68: op1_08_in24 = reg_0837;
    71: op1_08_in24 = reg_0430;
    75: op1_08_in24 = reg_0609;
    61: op1_08_in24 = reg_0438;
    114: op1_08_in24 = reg_0438;
    56: op1_08_in24 = reg_0185;
    87: op1_08_in24 = reg_1257;
    76: op1_08_in24 = reg_1290;
    57: op1_08_in24 = reg_0623;
    77: op1_08_in24 = reg_0166;
    58: op1_08_in24 = reg_0970;
    78: op1_08_in24 = reg_0703;
    70: op1_08_in24 = reg_0963;
    88: op1_08_in24 = reg_1214;
    46: op1_08_in24 = reg_0293;
    59: op1_08_in24 = reg_0168;
    79: op1_08_in24 = reg_0029;
    60: op1_08_in24 = reg_0395;
    80: op1_08_in24 = reg_0222;
    62: op1_08_in24 = reg_0352;
    48: op1_08_in24 = reg_0204;
    52: op1_08_in24 = reg_0067;
    81: op1_08_in24 = reg_0724;
    63: op1_08_in24 = reg_1164;
    82: op1_08_in24 = reg_0636;
    89: op1_08_in24 = reg_1502;
    83: op1_08_in24 = reg_0241;
    64: op1_08_in24 = reg_0397;
    112: op1_08_in24 = reg_0397;
    84: op1_08_in24 = reg_0398;
    65: op1_08_in24 = reg_0573;
    85: op1_08_in24 = reg_0434;
    121: op1_08_in24 = reg_0434;
    90: op1_08_in24 = reg_0906;
    66: op1_08_in24 = reg_0695;
    91: op1_08_in24 = reg_0300;
    67: op1_08_in24 = reg_0873;
    92: op1_08_in24 = reg_0110;
    93: op1_08_in24 = reg_0871;
    95: op1_08_in24 = reg_1004;
    98: op1_08_in24 = reg_1199;
    99: op1_08_in24 = imem05_in[15:12];
    44: op1_08_in24 = reg_0269;
    47: op1_08_in24 = reg_0459;
    101: op1_08_in24 = reg_0714;
    125: op1_08_in24 = reg_0714;
    40: op1_08_in24 = reg_0604;
    102: op1_08_in24 = reg_1254;
    103: op1_08_in24 = reg_0732;
    104: op1_08_in24 = reg_1198;
    105: op1_08_in24 = reg_0414;
    107: op1_08_in24 = reg_0114;
    108: op1_08_in24 = reg_0505;
    109: op1_08_in24 = reg_0563;
    110: op1_08_in24 = reg_0224;
    111: op1_08_in24 = reg_0600;
    113: op1_08_in24 = reg_0557;
    115: op1_08_in24 = reg_0088;
    116: op1_08_in24 = reg_1228;
    117: op1_08_in24 = reg_1298;
    119: op1_08_in24 = reg_0084;
    120: op1_08_in24 = reg_1312;
    122: op1_08_in24 = reg_0553;
    123: op1_08_in24 = reg_0144;
    124: op1_08_in24 = reg_0896;
    126: op1_08_in24 = reg_0902;
    42: op1_08_in24 = reg_0288;
    128: op1_08_in24 = imem07_in[15:12];
    129: op1_08_in24 = reg_0382;
    130: op1_08_in24 = reg_0167;
    131: op1_08_in24 = reg_1456;
    default: op1_08_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_08_inv24 = 1;
    55: op1_08_inv24 = 1;
    73: op1_08_inv24 = 1;
    69: op1_08_inv24 = 1;
    54: op1_08_inv24 = 1;
    56: op1_08_inv24 = 1;
    87: op1_08_inv24 = 1;
    57: op1_08_inv24 = 1;
    77: op1_08_inv24 = 1;
    88: op1_08_inv24 = 1;
    46: op1_08_inv24 = 1;
    59: op1_08_inv24 = 1;
    79: op1_08_inv24 = 1;
    82: op1_08_inv24 = 1;
    89: op1_08_inv24 = 1;
    83: op1_08_inv24 = 1;
    64: op1_08_inv24 = 1;
    65: op1_08_inv24 = 1;
    85: op1_08_inv24 = 1;
    90: op1_08_inv24 = 1;
    91: op1_08_inv24 = 1;
    92: op1_08_inv24 = 1;
    98: op1_08_inv24 = 1;
    99: op1_08_inv24 = 1;
    44: op1_08_inv24 = 1;
    40: op1_08_inv24 = 1;
    104: op1_08_inv24 = 1;
    107: op1_08_inv24 = 1;
    108: op1_08_inv24 = 1;
    111: op1_08_inv24 = 1;
    112: op1_08_inv24 = 1;
    115: op1_08_inv24 = 1;
    117: op1_08_inv24 = 1;
    120: op1_08_inv24 = 1;
    122: op1_08_inv24 = 1;
    123: op1_08_inv24 = 1;
    125: op1_08_inv24 = 1;
    128: op1_08_inv24 = 1;
    131: op1_08_inv24 = 1;
    default: op1_08_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in25 = reg_1347;
    53: op1_08_in25 = reg_0326;
    55: op1_08_in25 = reg_0052;
    86: op1_08_in25 = reg_1402;
    73: op1_08_in25 = reg_0490;
    69: op1_08_in25 = reg_0732;
    50: op1_08_in25 = reg_0758;
    54: op1_08_in25 = reg_0712;
    74: op1_08_in25 = reg_0553;
    68: op1_08_in25 = reg_0338;
    71: op1_08_in25 = reg_0383;
    75: op1_08_in25 = reg_0241;
    61: op1_08_in25 = reg_0727;
    56: op1_08_in25 = reg_0179;
    87: op1_08_in25 = reg_0297;
    76: op1_08_in25 = reg_1291;
    57: op1_08_in25 = reg_0591;
    77: op1_08_in25 = reg_1512;
    58: op1_08_in25 = reg_0972;
    78: op1_08_in25 = reg_0851;
    70: op1_08_in25 = reg_0220;
    88: op1_08_in25 = reg_1147;
    46: op1_08_in25 = reg_0145;
    59: op1_08_in25 = reg_0565;
    79: op1_08_in25 = reg_0284;
    60: op1_08_in25 = reg_1169;
    80: op1_08_in25 = reg_0242;
    62: op1_08_in25 = reg_1100;
    48: op1_08_in25 = reg_0206;
    52: op1_08_in25 = reg_0215;
    81: op1_08_in25 = reg_0875;
    63: op1_08_in25 = reg_0996;
    82: op1_08_in25 = reg_0979;
    89: op1_08_in25 = reg_0633;
    83: op1_08_in25 = reg_0742;
    64: op1_08_in25 = reg_0720;
    84: op1_08_in25 = reg_0585;
    65: op1_08_in25 = reg_0121;
    85: op1_08_in25 = reg_0091;
    90: op1_08_in25 = reg_0960;
    66: op1_08_in25 = reg_0024;
    91: op1_08_in25 = reg_1484;
    67: op1_08_in25 = reg_0301;
    92: op1_08_in25 = reg_0716;
    93: op1_08_in25 = reg_1253;
    95: op1_08_in25 = reg_0452;
    98: op1_08_in25 = reg_0178;
    99: op1_08_in25 = reg_0890;
    44: op1_08_in25 = reg_0023;
    47: op1_08_in25 = reg_0046;
    101: op1_08_in25 = reg_0619;
    40: op1_08_in25 = reg_0602;
    102: op1_08_in25 = reg_0166;
    103: op1_08_in25 = reg_0049;
    104: op1_08_in25 = reg_1200;
    105: op1_08_in25 = reg_0969;
    107: op1_08_in25 = reg_0228;
    108: op1_08_in25 = imem03_in[3:0];
    109: op1_08_in25 = reg_0233;
    110: op1_08_in25 = reg_0774;
    111: op1_08_in25 = reg_1495;
    112: op1_08_in25 = reg_0925;
    113: op1_08_in25 = reg_0823;
    114: op1_08_in25 = reg_1457;
    115: op1_08_in25 = reg_1258;
    116: op1_08_in25 = reg_0522;
    117: op1_08_in25 = imem05_in[3:0];
    119: op1_08_in25 = reg_1060;
    120: op1_08_in25 = reg_0117;
    121: op1_08_in25 = reg_0438;
    122: op1_08_in25 = reg_0550;
    123: op1_08_in25 = reg_1517;
    124: op1_08_in25 = reg_0162;
    125: op1_08_in25 = reg_0398;
    126: op1_08_in25 = reg_0163;
    42: op1_08_in25 = reg_0627;
    128: op1_08_in25 = reg_1055;
    129: op1_08_in25 = reg_0381;
    130: op1_08_in25 = reg_1181;
    131: op1_08_in25 = reg_0147;
    default: op1_08_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_08_inv25 = 1;
    50: op1_08_inv25 = 1;
    54: op1_08_inv25 = 1;
    68: op1_08_inv25 = 1;
    61: op1_08_inv25 = 1;
    87: op1_08_inv25 = 1;
    76: op1_08_inv25 = 1;
    57: op1_08_inv25 = 1;
    77: op1_08_inv25 = 1;
    58: op1_08_inv25 = 1;
    88: op1_08_inv25 = 1;
    59: op1_08_inv25 = 1;
    79: op1_08_inv25 = 1;
    52: op1_08_inv25 = 1;
    81: op1_08_inv25 = 1;
    63: op1_08_inv25 = 1;
    89: op1_08_inv25 = 1;
    83: op1_08_inv25 = 1;
    84: op1_08_inv25 = 1;
    85: op1_08_inv25 = 1;
    66: op1_08_inv25 = 1;
    91: op1_08_inv25 = 1;
    92: op1_08_inv25 = 1;
    40: op1_08_inv25 = 1;
    102: op1_08_inv25 = 1;
    103: op1_08_inv25 = 1;
    104: op1_08_inv25 = 1;
    105: op1_08_inv25 = 1;
    107: op1_08_inv25 = 1;
    108: op1_08_inv25 = 1;
    110: op1_08_inv25 = 1;
    113: op1_08_inv25 = 1;
    120: op1_08_inv25 = 1;
    125: op1_08_inv25 = 1;
    126: op1_08_inv25 = 1;
    129: op1_08_inv25 = 1;
    130: op1_08_inv25 = 1;
    default: op1_08_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in26 = reg_1345;
    53: op1_08_in26 = reg_0778;
    55: op1_08_in26 = reg_0053;
    86: op1_08_in26 = reg_1070;
    73: op1_08_in26 = reg_0491;
    69: op1_08_in26 = reg_0121;
    50: op1_08_in26 = reg_0734;
    54: op1_08_in26 = reg_0217;
    74: op1_08_in26 = reg_0241;
    68: op1_08_in26 = reg_0236;
    71: op1_08_in26 = reg_0091;
    75: op1_08_in26 = reg_1474;
    61: op1_08_in26 = reg_0147;
    56: op1_08_in26 = reg_0144;
    87: op1_08_in26 = reg_0574;
    76: op1_08_in26 = reg_1513;
    57: op1_08_in26 = reg_0103;
    77: op1_08_in26 = reg_0047;
    58: op1_08_in26 = reg_0935;
    78: op1_08_in26 = reg_0297;
    70: op1_08_in26 = reg_1301;
    88: op1_08_in26 = reg_0342;
    46: op1_08_in26 = reg_0559;
    59: op1_08_in26 = reg_0045;
    79: op1_08_in26 = reg_0286;
    60: op1_08_in26 = reg_0174;
    80: op1_08_in26 = reg_0438;
    62: op1_08_in26 = reg_1253;
    48: op1_08_in26 = reg_0784;
    52: op1_08_in26 = reg_0022;
    81: op1_08_in26 = reg_0874;
    63: op1_08_in26 = reg_0131;
    82: op1_08_in26 = reg_0522;
    89: op1_08_in26 = reg_1488;
    83: op1_08_in26 = reg_0612;
    64: op1_08_in26 = reg_1323;
    84: op1_08_in26 = reg_0373;
    65: op1_08_in26 = reg_0216;
    85: op1_08_in26 = imem01_in[3:0];
    90: op1_08_in26 = reg_0133;
    66: op1_08_in26 = reg_0325;
    91: op1_08_in26 = reg_0492;
    67: op1_08_in26 = reg_0274;
    92: op1_08_in26 = reg_0636;
    93: op1_08_in26 = reg_0277;
    95: op1_08_in26 = reg_0033;
    98: op1_08_in26 = reg_1208;
    99: op1_08_in26 = reg_1059;
    44: op1_08_in26 = reg_0215;
    47: op1_08_in26 = imem07_in[3:0];
    101: op1_08_in26 = reg_0570;
    40: op1_08_in26 = reg_0603;
    102: op1_08_in26 = reg_0902;
    103: op1_08_in26 = reg_1449;
    104: op1_08_in26 = reg_0488;
    105: op1_08_in26 = reg_0599;
    107: op1_08_in26 = reg_0001;
    108: op1_08_in26 = imem03_in[7:4];
    109: op1_08_in26 = reg_0049;
    110: op1_08_in26 = reg_0287;
    111: op1_08_in26 = reg_0965;
    112: op1_08_in26 = reg_0870;
    113: op1_08_in26 = reg_0143;
    114: op1_08_in26 = reg_0868;
    115: op1_08_in26 = reg_0978;
    116: op1_08_in26 = reg_0323;
    117: op1_08_in26 = imem05_in[15:12];
    119: op1_08_in26 = reg_0703;
    120: op1_08_in26 = reg_0065;
    121: op1_08_in26 = reg_0360;
    122: op1_08_in26 = reg_0609;
    123: op1_08_in26 = reg_0505;
    124: op1_08_in26 = reg_0041;
    125: op1_08_in26 = reg_0619;
    126: op1_08_in26 = reg_0331;
    42: op1_08_in26 = reg_0377;
    128: op1_08_in26 = reg_1315;
    129: op1_08_in26 = reg_0829;
    130: op1_08_in26 = reg_1404;
    131: op1_08_in26 = reg_0963;
    default: op1_08_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_08_inv26 = 1;
    73: op1_08_inv26 = 1;
    69: op1_08_inv26 = 1;
    50: op1_08_inv26 = 1;
    68: op1_08_inv26 = 1;
    71: op1_08_inv26 = 1;
    75: op1_08_inv26 = 1;
    61: op1_08_inv26 = 1;
    87: op1_08_inv26 = 1;
    76: op1_08_inv26 = 1;
    57: op1_08_inv26 = 1;
    77: op1_08_inv26 = 1;
    58: op1_08_inv26 = 1;
    70: op1_08_inv26 = 1;
    46: op1_08_inv26 = 1;
    80: op1_08_inv26 = 1;
    48: op1_08_inv26 = 1;
    52: op1_08_inv26 = 1;
    63: op1_08_inv26 = 1;
    89: op1_08_inv26 = 1;
    64: op1_08_inv26 = 1;
    90: op1_08_inv26 = 1;
    66: op1_08_inv26 = 1;
    93: op1_08_inv26 = 1;
    44: op1_08_inv26 = 1;
    47: op1_08_inv26 = 1;
    101: op1_08_inv26 = 1;
    102: op1_08_inv26 = 1;
    103: op1_08_inv26 = 1;
    108: op1_08_inv26 = 1;
    109: op1_08_inv26 = 1;
    110: op1_08_inv26 = 1;
    112: op1_08_inv26 = 1;
    113: op1_08_inv26 = 1;
    116: op1_08_inv26 = 1;
    121: op1_08_inv26 = 1;
    122: op1_08_inv26 = 1;
    128: op1_08_inv26 = 1;
    131: op1_08_inv26 = 1;
    default: op1_08_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in27 = reg_0777;
    53: op1_08_in27 = reg_0973;
    86: op1_08_in27 = reg_0090;
    73: op1_08_in27 = reg_0025;
    69: op1_08_in27 = reg_0216;
    50: op1_08_in27 = reg_0677;
    54: op1_08_in27 = reg_0325;
    74: op1_08_in27 = reg_0798;
    68: op1_08_in27 = reg_0237;
    71: op1_08_in27 = reg_0291;
    75: op1_08_in27 = reg_0819;
    61: op1_08_in27 = reg_0149;
    56: op1_08_in27 = reg_0954;
    87: op1_08_in27 = reg_0412;
    76: op1_08_in27 = reg_0463;
    77: op1_08_in27 = reg_0463;
    57: op1_08_in27 = reg_0100;
    58: op1_08_in27 = reg_0933;
    78: op1_08_in27 = reg_1350;
    70: op1_08_in27 = reg_0178;
    88: op1_08_in27 = reg_0097;
    46: op1_08_in27 = reg_0104;
    59: op1_08_in27 = reg_1180;
    79: op1_08_in27 = reg_0366;
    60: op1_08_in27 = reg_0066;
    80: op1_08_in27 = reg_0146;
    62: op1_08_in27 = reg_1254;
    48: op1_08_in27 = reg_0192;
    52: op1_08_in27 = imem07_in[3:0];
    81: op1_08_in27 = reg_0080;
    63: op1_08_in27 = reg_0045;
    40: op1_08_in27 = reg_0045;
    82: op1_08_in27 = reg_0419;
    89: op1_08_in27 = imem05_in[11:8];
    83: op1_08_in27 = reg_0430;
    64: op1_08_in27 = reg_0827;
    84: op1_08_in27 = reg_0584;
    65: op1_08_in27 = reg_0630;
    85: op1_08_in27 = imem01_in[7:4];
    90: op1_08_in27 = reg_0860;
    66: op1_08_in27 = reg_1132;
    91: op1_08_in27 = imem05_in[7:4];
    67: op1_08_in27 = reg_0602;
    92: op1_08_in27 = reg_0194;
    93: op1_08_in27 = reg_0258;
    95: op1_08_in27 = reg_0369;
    98: op1_08_in27 = reg_0107;
    99: op1_08_in27 = reg_0793;
    120: op1_08_in27 = reg_0793;
    44: op1_08_in27 = reg_0022;
    47: op1_08_in27 = reg_0324;
    101: op1_08_in27 = reg_0979;
    102: op1_08_in27 = reg_0553;
    103: op1_08_in27 = reg_1063;
    104: op1_08_in27 = reg_1233;
    105: op1_08_in27 = reg_1237;
    108: op1_08_in27 = reg_0049;
    109: op1_08_in27 = reg_1003;
    110: op1_08_in27 = reg_0741;
    111: op1_08_in27 = reg_0627;
    112: op1_08_in27 = reg_0730;
    113: op1_08_in27 = reg_0000;
    114: op1_08_in27 = reg_1513;
    115: op1_08_in27 = reg_0462;
    116: op1_08_in27 = reg_0394;
    117: op1_08_in27 = reg_0136;
    119: op1_08_in27 = reg_0309;
    121: op1_08_in27 = reg_0899;
    122: op1_08_in27 = reg_0242;
    123: op1_08_in27 = reg_0329;
    124: op1_08_in27 = reg_1103;
    125: op1_08_in27 = reg_0528;
    126: op1_08_in27 = reg_0549;
    42: op1_08_in27 = reg_0235;
    128: op1_08_in27 = reg_0457;
    129: op1_08_in27 = reg_0745;
    130: op1_08_in27 = reg_0940;
    131: op1_08_in27 = reg_0464;
    default: op1_08_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv27 = 1;
    53: op1_08_inv27 = 1;
    86: op1_08_inv27 = 1;
    73: op1_08_inv27 = 1;
    69: op1_08_inv27 = 1;
    50: op1_08_inv27 = 1;
    54: op1_08_inv27 = 1;
    74: op1_08_inv27 = 1;
    68: op1_08_inv27 = 1;
    71: op1_08_inv27 = 1;
    61: op1_08_inv27 = 1;
    56: op1_08_inv27 = 1;
    87: op1_08_inv27 = 1;
    57: op1_08_inv27 = 1;
    46: op1_08_inv27 = 1;
    59: op1_08_inv27 = 1;
    79: op1_08_inv27 = 1;
    48: op1_08_inv27 = 1;
    63: op1_08_inv27 = 1;
    82: op1_08_inv27 = 1;
    64: op1_08_inv27 = 1;
    65: op1_08_inv27 = 1;
    85: op1_08_inv27 = 1;
    90: op1_08_inv27 = 1;
    66: op1_08_inv27 = 1;
    67: op1_08_inv27 = 1;
    92: op1_08_inv27 = 1;
    98: op1_08_inv27 = 1;
    44: op1_08_inv27 = 1;
    47: op1_08_inv27 = 1;
    103: op1_08_inv27 = 1;
    105: op1_08_inv27 = 1;
    110: op1_08_inv27 = 1;
    114: op1_08_inv27 = 1;
    120: op1_08_inv27 = 1;
    121: op1_08_inv27 = 1;
    123: op1_08_inv27 = 1;
    126: op1_08_inv27 = 1;
    42: op1_08_inv27 = 1;
    128: op1_08_inv27 = 1;
    129: op1_08_inv27 = 1;
    131: op1_08_inv27 = 1;
    default: op1_08_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in28 = reg_0664;
    53: op1_08_in28 = reg_0106;
    58: op1_08_in28 = reg_0106;
    86: op1_08_in28 = reg_0872;
    73: op1_08_in28 = reg_0667;
    69: op1_08_in28 = imem03_in[11:8];
    50: op1_08_in28 = reg_0216;
    54: op1_08_in28 = reg_0573;
    74: op1_08_in28 = reg_0820;
    68: op1_08_in28 = reg_0117;
    71: op1_08_in28 = reg_0277;
    75: op1_08_in28 = reg_0385;
    61: op1_08_in28 = reg_0148;
    56: op1_08_in28 = reg_0107;
    70: op1_08_in28 = reg_0107;
    87: op1_08_in28 = reg_0097;
    76: op1_08_in28 = reg_0260;
    57: op1_08_in28 = reg_0321;
    77: op1_08_in28 = reg_0331;
    78: op1_08_in28 = reg_1345;
    88: op1_08_in28 = reg_0305;
    46: op1_08_in28 = reg_0884;
    59: op1_08_in28 = reg_0316;
    79: op1_08_in28 = reg_0620;
    60: op1_08_in28 = reg_1212;
    80: op1_08_in28 = reg_0384;
    62: op1_08_in28 = reg_1070;
    48: op1_08_in28 = imem06_in[15:12];
    52: op1_08_in28 = imem07_in[15:12];
    81: op1_08_in28 = reg_0077;
    63: op1_08_in28 = reg_0938;
    82: op1_08_in28 = reg_1202;
    89: op1_08_in28 = reg_0737;
    83: op1_08_in28 = reg_0726;
    64: op1_08_in28 = reg_0110;
    84: op1_08_in28 = reg_1228;
    65: op1_08_in28 = reg_0707;
    85: op1_08_in28 = reg_0043;
    90: op1_08_in28 = reg_0827;
    66: op1_08_in28 = reg_0525;
    91: op1_08_in28 = reg_0449;
    67: op1_08_in28 = reg_1346;
    92: op1_08_in28 = reg_0584;
    93: op1_08_in28 = reg_0547;
    95: op1_08_in28 = reg_0262;
    98: op1_08_in28 = reg_0291;
    99: op1_08_in28 = reg_0136;
    44: op1_08_in28 = reg_0252;
    47: op1_08_in28 = reg_0894;
    101: op1_08_in28 = reg_0308;
    40: op1_08_in28 = reg_0490;
    102: op1_08_in28 = reg_0258;
    103: op1_08_in28 = reg_1425;
    104: op1_08_in28 = reg_0281;
    105: op1_08_in28 = reg_0096;
    108: op1_08_in28 = reg_1063;
    109: op1_08_in28 = reg_0840;
    110: op1_08_in28 = reg_0102;
    111: op1_08_in28 = reg_1093;
    123: op1_08_in28 = reg_1093;
    112: op1_08_in28 = reg_0265;
    113: op1_08_in28 = reg_1518;
    114: op1_08_in28 = reg_0362;
    115: op1_08_in28 = reg_0531;
    116: op1_08_in28 = reg_1095;
    117: op1_08_in28 = reg_0272;
    119: op1_08_in28 = reg_0457;
    120: op1_08_in28 = reg_0205;
    121: op1_08_in28 = reg_0464;
    122: op1_08_in28 = reg_0967;
    124: op1_08_in28 = imem02_in[11:8];
    125: op1_08_in28 = reg_0571;
    126: op1_08_in28 = reg_0550;
    42: op1_08_in28 = reg_0234;
    128: op1_08_in28 = reg_1349;
    129: op1_08_in28 = reg_0294;
    130: op1_08_in28 = reg_0792;
    131: op1_08_in28 = reg_0400;
    default: op1_08_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv28 = 1;
    53: op1_08_inv28 = 1;
    86: op1_08_inv28 = 1;
    54: op1_08_inv28 = 1;
    74: op1_08_inv28 = 1;
    87: op1_08_inv28 = 1;
    57: op1_08_inv28 = 1;
    88: op1_08_inv28 = 1;
    79: op1_08_inv28 = 1;
    80: op1_08_inv28 = 1;
    63: op1_08_inv28 = 1;
    83: op1_08_inv28 = 1;
    65: op1_08_inv28 = 1;
    93: op1_08_inv28 = 1;
    95: op1_08_inv28 = 1;
    44: op1_08_inv28 = 1;
    101: op1_08_inv28 = 1;
    40: op1_08_inv28 = 1;
    103: op1_08_inv28 = 1;
    104: op1_08_inv28 = 1;
    105: op1_08_inv28 = 1;
    111: op1_08_inv28 = 1;
    112: op1_08_inv28 = 1;
    114: op1_08_inv28 = 1;
    116: op1_08_inv28 = 1;
    120: op1_08_inv28 = 1;
    121: op1_08_inv28 = 1;
    122: op1_08_inv28 = 1;
    123: op1_08_inv28 = 1;
    125: op1_08_inv28 = 1;
    128: op1_08_inv28 = 1;
    129: op1_08_inv28 = 1;
    default: op1_08_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in29 = reg_0286;
    53: op1_08_in29 = reg_0380;
    86: op1_08_in29 = reg_1486;
    73: op1_08_in29 = reg_0703;
    69: op1_08_in29 = reg_1139;
    50: op1_08_in29 = reg_0227;
    54: op1_08_in29 = reg_0198;
    74: op1_08_in29 = reg_0257;
    68: op1_08_in29 = reg_0211;
    71: op1_08_in29 = reg_0011;
    75: op1_08_in29 = reg_0383;
    61: op1_08_in29 = reg_0146;
    56: op1_08_in29 = reg_0113;
    87: op1_08_in29 = reg_0061;
    76: op1_08_in29 = reg_1473;
    57: op1_08_in29 = reg_0050;
    77: op1_08_in29 = reg_0548;
    58: op1_08_in29 = reg_0055;
    78: op1_08_in29 = reg_1349;
    70: op1_08_in29 = reg_0481;
    88: op1_08_in29 = reg_0339;
    46: op1_08_in29 = reg_0507;
    59: op1_08_in29 = reg_0939;
    79: op1_08_in29 = reg_0103;
    60: op1_08_in29 = reg_0541;
    80: op1_08_in29 = reg_0385;
    62: op1_08_in29 = reg_1033;
    48: op1_08_in29 = reg_0977;
    52: op1_08_in29 = reg_1060;
    81: op1_08_in29 = reg_0042;
    63: op1_08_in29 = imem05_in[15:12];
    82: op1_08_in29 = reg_1179;
    89: op1_08_in29 = reg_0205;
    83: op1_08_in29 = reg_0148;
    64: op1_08_in29 = reg_0373;
    84: op1_08_in29 = reg_0119;
    65: op1_08_in29 = reg_0375;
    85: op1_08_in29 = reg_0332;
    90: op1_08_in29 = reg_1501;
    66: op1_08_in29 = reg_0734;
    91: op1_08_in29 = imem06_in[15:12];
    67: op1_08_in29 = reg_0864;
    92: op1_08_in29 = reg_0244;
    93: op1_08_in29 = reg_0747;
    102: op1_08_in29 = reg_0747;
    126: op1_08_in29 = reg_0747;
    95: op1_08_in29 = reg_0836;
    98: op1_08_in29 = reg_0348;
    42: op1_08_in29 = reg_0348;
    99: op1_08_in29 = reg_0702;
    44: op1_08_in29 = imem07_in[3:0];
    47: op1_08_in29 = reg_0893;
    101: op1_08_in29 = reg_1202;
    40: op1_08_in29 = reg_0418;
    103: op1_08_in29 = reg_1001;
    104: op1_08_in29 = reg_0500;
    105: op1_08_in29 = reg_1189;
    108: op1_08_in29 = reg_0216;
    109: op1_08_in29 = reg_0312;
    110: op1_08_in29 = reg_0361;
    111: op1_08_in29 = reg_0884;
    112: op1_08_in29 = reg_0585;
    113: op1_08_in29 = reg_0627;
    114: op1_08_in29 = reg_0360;
    115: op1_08_in29 = reg_0552;
    116: op1_08_in29 = reg_0298;
    117: op1_08_in29 = reg_0176;
    119: op1_08_in29 = reg_1350;
    120: op1_08_in29 = reg_0251;
    121: op1_08_in29 = reg_0292;
    122: op1_08_in29 = reg_0430;
    123: op1_08_in29 = reg_0882;
    124: op1_08_in29 = reg_0423;
    125: op1_08_in29 = reg_0979;
    128: op1_08_in29 = reg_0031;
    129: op1_08_in29 = reg_1091;
    130: op1_08_in29 = reg_0937;
    131: op1_08_in29 = reg_0043;
    default: op1_08_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv29 = 1;
    86: op1_08_inv29 = 1;
    69: op1_08_inv29 = 1;
    68: op1_08_inv29 = 1;
    71: op1_08_inv29 = 1;
    75: op1_08_inv29 = 1;
    61: op1_08_inv29 = 1;
    76: op1_08_inv29 = 1;
    58: op1_08_inv29 = 1;
    70: op1_08_inv29 = 1;
    46: op1_08_inv29 = 1;
    60: op1_08_inv29 = 1;
    80: op1_08_inv29 = 1;
    48: op1_08_inv29 = 1;
    81: op1_08_inv29 = 1;
    89: op1_08_inv29 = 1;
    83: op1_08_inv29 = 1;
    64: op1_08_inv29 = 1;
    84: op1_08_inv29 = 1;
    65: op1_08_inv29 = 1;
    90: op1_08_inv29 = 1;
    91: op1_08_inv29 = 1;
    67: op1_08_inv29 = 1;
    93: op1_08_inv29 = 1;
    95: op1_08_inv29 = 1;
    98: op1_08_inv29 = 1;
    99: op1_08_inv29 = 1;
    44: op1_08_inv29 = 1;
    102: op1_08_inv29 = 1;
    104: op1_08_inv29 = 1;
    105: op1_08_inv29 = 1;
    111: op1_08_inv29 = 1;
    112: op1_08_inv29 = 1;
    114: op1_08_inv29 = 1;
    115: op1_08_inv29 = 1;
    117: op1_08_inv29 = 1;
    121: op1_08_inv29 = 1;
    124: op1_08_inv29 = 1;
    125: op1_08_inv29 = 1;
    42: op1_08_inv29 = 1;
    131: op1_08_inv29 = 1;
    default: op1_08_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_08_in30 = reg_0366;
    53: op1_08_in30 = reg_0712;
    58: op1_08_in30 = reg_0712;
    86: op1_08_in30 = reg_1484;
    73: op1_08_in30 = reg_0140;
    69: op1_08_in30 = reg_0638;
    50: op1_08_in30 = reg_0288;
    54: op1_08_in30 = reg_1064;
    74: op1_08_in30 = reg_0875;
    80: op1_08_in30 = reg_0875;
    68: op1_08_in30 = reg_0064;
    71: op1_08_in30 = reg_0010;
    75: op1_08_in30 = reg_0362;
    61: op1_08_in30 = reg_0360;
    56: op1_08_in30 = reg_0507;
    87: op1_08_in30 = reg_0582;
    76: op1_08_in30 = reg_0468;
    57: op1_08_in30 = reg_0004;
    77: op1_08_in30 = reg_0746;
    78: op1_08_in30 = reg_0157;
    70: op1_08_in30 = reg_0831;
    88: op1_08_in30 = reg_0904;
    46: op1_08_in30 = reg_0481;
    59: op1_08_in30 = reg_0167;
    79: op1_08_in30 = reg_0028;
    60: op1_08_in30 = reg_0450;
    62: op1_08_in30 = reg_0547;
    48: op1_08_in30 = reg_0906;
    52: op1_08_in30 = reg_0998;
    81: op1_08_in30 = reg_0332;
    63: op1_08_in30 = reg_0861;
    82: op1_08_in30 = reg_0270;
    89: op1_08_in30 = reg_0315;
    83: op1_08_in30 = reg_0384;
    64: op1_08_in30 = reg_0529;
    84: op1_08_in30 = reg_1202;
    92: op1_08_in30 = reg_1202;
    65: op1_08_in30 = reg_1139;
    85: op1_08_in30 = reg_0744;
    90: op1_08_in30 = reg_0635;
    66: op1_08_in30 = reg_0675;
    91: op1_08_in30 = reg_0870;
    67: op1_08_in30 = reg_0828;
    93: op1_08_in30 = reg_0239;
    95: op1_08_in30 = reg_0835;
    98: op1_08_in30 = reg_0427;
    99: op1_08_in30 = reg_0395;
    44: op1_08_in30 = imem07_in[7:4];
    47: op1_08_in30 = reg_0187;
    101: op1_08_in30 = reg_0371;
    40: op1_08_in30 = reg_0090;
    102: op1_08_in30 = reg_0787;
    103: op1_08_in30 = reg_0600;
    104: op1_08_in30 = reg_0421;
    105: op1_08_in30 = reg_0470;
    108: op1_08_in30 = reg_0180;
    109: op1_08_in30 = reg_0180;
    110: op1_08_in30 = reg_0050;
    111: op1_08_in30 = reg_0458;
    112: op1_08_in30 = reg_0622;
    113: op1_08_in30 = reg_0756;
    114: op1_08_in30 = reg_0899;
    115: op1_08_in30 = reg_1203;
    116: op1_08_in30 = reg_1056;
    117: op1_08_in30 = reg_0391;
    119: op1_08_in30 = reg_0223;
    120: op1_08_in30 = reg_0174;
    121: op1_08_in30 = reg_0162;
    122: op1_08_in30 = reg_0434;
    123: op1_08_in30 = reg_0673;
    124: op1_08_in30 = reg_0588;
    125: op1_08_in30 = reg_0244;
    126: op1_08_in30 = reg_0609;
    42: op1_08_in30 = reg_0597;
    128: op1_08_in30 = reg_0665;
    129: op1_08_in30 = reg_0068;
    130: op1_08_in30 = reg_0300;
    131: op1_08_in30 = reg_0125;
    default: op1_08_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_08_inv30 = 1;
    53: op1_08_inv30 = 1;
    73: op1_08_inv30 = 1;
    74: op1_08_inv30 = 1;
    61: op1_08_inv30 = 1;
    56: op1_08_inv30 = 1;
    57: op1_08_inv30 = 1;
    78: op1_08_inv30 = 1;
    88: op1_08_inv30 = 1;
    46: op1_08_inv30 = 1;
    59: op1_08_inv30 = 1;
    60: op1_08_inv30 = 1;
    48: op1_08_inv30 = 1;
    52: op1_08_inv30 = 1;
    84: op1_08_inv30 = 1;
    65: op1_08_inv30 = 1;
    85: op1_08_inv30 = 1;
    90: op1_08_inv30 = 1;
    91: op1_08_inv30 = 1;
    67: op1_08_inv30 = 1;
    98: op1_08_inv30 = 1;
    47: op1_08_inv30 = 1;
    101: op1_08_inv30 = 1;
    103: op1_08_inv30 = 1;
    105: op1_08_inv30 = 1;
    110: op1_08_inv30 = 1;
    112: op1_08_inv30 = 1;
    113: op1_08_inv30 = 1;
    114: op1_08_inv30 = 1;
    115: op1_08_inv30 = 1;
    116: op1_08_inv30 = 1;
    117: op1_08_inv30 = 1;
    119: op1_08_inv30 = 1;
    121: op1_08_inv30 = 1;
    123: op1_08_inv30 = 1;
    125: op1_08_inv30 = 1;
    126: op1_08_inv30 = 1;
    128: op1_08_inv30 = 1;
    default: op1_08_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_08_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#8の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_08_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in00 = reg_0182;
    53: op1_09_in00 = reg_0574;
    86: op1_09_in00 = reg_0848;
    55: op1_09_in00 = reg_0527;
    73: op1_09_in00 = reg_0219;
    69: op1_09_in00 = reg_0839;
    49: op1_09_in00 = reg_0310;
    74: op1_09_in00 = reg_0735;
    54: op1_09_in00 = reg_0383;
    68: op1_09_in00 = reg_0048;
    75: op1_09_in00 = reg_1430;
    50: op1_09_in00 = reg_0585;
    56: op1_09_in00 = reg_0394;
    71: op1_09_in00 = reg_0554;
    87: op1_09_in00 = reg_0179;
    76: op1_09_in00 = imem05_in[7:4];
    61: op1_09_in00 = reg_0803;
    57: op1_09_in00 = reg_1151;
    77: op1_09_in00 = reg_0210;
    58: op1_09_in00 = reg_0419;
    78: op1_09_in00 = reg_1510;
    82: op1_09_in00 = reg_1510;
    70: op1_09_in00 = imem03_in[7:4];
    51: op1_09_in00 = reg_0297;
    79: op1_09_in00 = reg_0555;
    59: op1_09_in00 = reg_0403;
    88: op1_09_in00 = reg_0559;
    60: op1_09_in00 = reg_0301;
    46: op1_09_in00 = reg_0702;
    62: op1_09_in00 = reg_0550;
    80: op1_09_in00 = reg_0575;
    48: op1_09_in00 = reg_0726;
    81: op1_09_in00 = reg_0457;
    52: op1_09_in00 = reg_0305;
    33: op1_09_in00 = imem07_in[11:8];
    28: op1_09_in00 = imem07_in[11:8];
    63: op1_09_in00 = reg_0615;
    89: op1_09_in00 = reg_0326;
    83: op1_09_in00 = reg_0037;
    64: op1_09_in00 = reg_0568;
    84: op1_09_in00 = reg_1278;
    85: op1_09_in00 = reg_0530;
    65: op1_09_in00 = reg_1300;
    90: op1_09_in00 = reg_0780;
    66: op1_09_in00 = imem07_in[15:12];
    37: op1_09_in00 = reg_0673;
    111: op1_09_in00 = reg_0673;
    91: op1_09_in00 = reg_1079;
    67: op1_09_in00 = imem06_in[11:8];
    92: op1_09_in00 = imem00_in[11:8];
    93: op1_09_in00 = reg_0742;
    94: op1_09_in00 = imem00_in[3:0];
    118: op1_09_in00 = imem00_in[3:0];
    128: op1_09_in00 = imem00_in[3:0];
    95: op1_09_in00 = reg_0344;
    96: op1_09_in00 = imem00_in[15:12];
    110: op1_09_in00 = imem00_in[15:12];
    97: op1_09_in00 = reg_1241;
    98: op1_09_in00 = reg_1372;
    99: op1_09_in00 = reg_0992;
    100: op1_09_in00 = reg_1281;
    101: op1_09_in00 = reg_0023;
    102: op1_09_in00 = reg_0222;
    103: op1_09_in00 = reg_1495;
    44: op1_09_in00 = reg_0796;
    104: op1_09_in00 = imem06_in[15:12];
    47: op1_09_in00 = reg_0459;
    105: op1_09_in00 = reg_0370;
    106: op1_09_in00 = imem00_in[7:4];
    119: op1_09_in00 = imem00_in[7:4];
    107: op1_09_in00 = reg_1244;
    108: op1_09_in00 = reg_0891;
    109: op1_09_in00 = reg_0375;
    112: op1_09_in00 = reg_0619;
    113: op1_09_in00 = reg_0558;
    114: op1_09_in00 = reg_0078;
    115: op1_09_in00 = reg_1200;
    116: op1_09_in00 = reg_1101;
    117: op1_09_in00 = reg_0701;
    40: op1_09_in00 = reg_0412;
    120: op1_09_in00 = reg_0926;
    121: op1_09_in00 = reg_0728;
    122: op1_09_in00 = reg_1032;
    34: op1_09_in00 = reg_0139;
    123: op1_09_in00 = reg_1280;
    124: op1_09_in00 = reg_0055;
    125: op1_09_in00 = reg_1204;
    126: op1_09_in00 = reg_0241;
    127: op1_09_in00 = reg_1080;
    38: op1_09_in00 = reg_0029;
    42: op1_09_in00 = reg_0167;
    129: op1_09_in00 = reg_0279;
    130: op1_09_in00 = reg_0196;
    131: op1_09_in00 = reg_0561;
    default: op1_09_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_09_inv00 = 1;
    69: op1_09_inv00 = 1;
    49: op1_09_inv00 = 1;
    74: op1_09_inv00 = 1;
    68: op1_09_inv00 = 1;
    87: op1_09_inv00 = 1;
    76: op1_09_inv00 = 1;
    61: op1_09_inv00 = 1;
    57: op1_09_inv00 = 1;
    77: op1_09_inv00 = 1;
    58: op1_09_inv00 = 1;
    70: op1_09_inv00 = 1;
    51: op1_09_inv00 = 1;
    88: op1_09_inv00 = 1;
    46: op1_09_inv00 = 1;
    62: op1_09_inv00 = 1;
    48: op1_09_inv00 = 1;
    81: op1_09_inv00 = 1;
    63: op1_09_inv00 = 1;
    89: op1_09_inv00 = 1;
    64: op1_09_inv00 = 1;
    84: op1_09_inv00 = 1;
    85: op1_09_inv00 = 1;
    65: op1_09_inv00 = 1;
    28: op1_09_inv00 = 1;
    90: op1_09_inv00 = 1;
    37: op1_09_inv00 = 1;
    91: op1_09_inv00 = 1;
    67: op1_09_inv00 = 1;
    93: op1_09_inv00 = 1;
    95: op1_09_inv00 = 1;
    96: op1_09_inv00 = 1;
    98: op1_09_inv00 = 1;
    100: op1_09_inv00 = 1;
    44: op1_09_inv00 = 1;
    104: op1_09_inv00 = 1;
    47: op1_09_inv00 = 1;
    105: op1_09_inv00 = 1;
    108: op1_09_inv00 = 1;
    109: op1_09_inv00 = 1;
    111: op1_09_inv00 = 1;
    112: op1_09_inv00 = 1;
    113: op1_09_inv00 = 1;
    114: op1_09_inv00 = 1;
    116: op1_09_inv00 = 1;
    117: op1_09_inv00 = 1;
    118: op1_09_inv00 = 1;
    119: op1_09_inv00 = 1;
    121: op1_09_inv00 = 1;
    122: op1_09_inv00 = 1;
    34: op1_09_inv00 = 1;
    124: op1_09_inv00 = 1;
    126: op1_09_inv00 = 1;
    127: op1_09_inv00 = 1;
    38: op1_09_inv00 = 1;
    42: op1_09_inv00 = 1;
    130: op1_09_inv00 = 1;
    131: op1_09_inv00 = 1;
    default: op1_09_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in01 = reg_0045;
    53: op1_09_in01 = reg_0464;
    86: op1_09_in01 = reg_0009;
    55: op1_09_in01 = imem06_in[7:4];
    73: op1_09_in01 = reg_0701;
    69: op1_09_in01 = reg_0846;
    49: op1_09_in01 = reg_0297;
    56: op1_09_in01 = reg_0297;
    74: op1_09_in01 = reg_0251;
    54: op1_09_in01 = reg_0724;
    68: op1_09_in01 = reg_0329;
    75: op1_09_in01 = reg_1164;
    50: op1_09_in01 = reg_0586;
    71: op1_09_in01 = reg_0844;
    87: op1_09_in01 = reg_1033;
    76: op1_09_in01 = reg_0937;
    61: op1_09_in01 = reg_0523;
    57: op1_09_in01 = reg_0982;
    77: op1_09_in01 = reg_0736;
    58: op1_09_in01 = reg_0289;
    78: op1_09_in01 = reg_1081;
    94: op1_09_in01 = reg_1081;
    127: op1_09_in01 = reg_1081;
    70: op1_09_in01 = imem03_in[11:8];
    51: op1_09_in01 = reg_0673;
    79: op1_09_in01 = imem00_in[7:4];
    118: op1_09_in01 = imem00_in[7:4];
    59: op1_09_in01 = reg_0384;
    88: op1_09_in01 = reg_0233;
    60: op1_09_in01 = reg_0243;
    46: op1_09_in01 = reg_0176;
    62: op1_09_in01 = reg_0548;
    80: op1_09_in01 = reg_0799;
    48: op1_09_in01 = reg_0401;
    81: op1_09_in01 = reg_0626;
    52: op1_09_in01 = reg_0262;
    33: op1_09_in01 = reg_0137;
    63: op1_09_in01 = reg_0445;
    91: op1_09_in01 = reg_0445;
    82: op1_09_in01 = reg_0868;
    89: op1_09_in01 = reg_1458;
    83: op1_09_in01 = reg_0751;
    64: op1_09_in01 = reg_0522;
    84: op1_09_in01 = reg_0841;
    85: op1_09_in01 = reg_0607;
    65: op1_09_in01 = reg_0048;
    90: op1_09_in01 = reg_1035;
    66: op1_09_in01 = reg_0461;
    37: op1_09_in01 = reg_0156;
    67: op1_09_in01 = reg_0977;
    92: op1_09_in01 = reg_1241;
    96: op1_09_in01 = reg_1241;
    93: op1_09_in01 = reg_0439;
    95: op1_09_in01 = reg_0449;
    97: op1_09_in01 = reg_0672;
    98: op1_09_in01 = reg_1368;
    123: op1_09_in01 = reg_1368;
    99: op1_09_in01 = reg_0334;
    100: op1_09_in01 = imem00_in[3:0];
    101: op1_09_in01 = reg_0791;
    106: op1_09_in01 = reg_0791;
    102: op1_09_in01 = reg_0242;
    103: op1_09_in01 = reg_0142;
    44: op1_09_in01 = reg_0797;
    104: op1_09_in01 = reg_1105;
    47: op1_09_in01 = reg_0268;
    105: op1_09_in01 = reg_1298;
    107: op1_09_in01 = reg_1487;
    108: op1_09_in01 = reg_1495;
    109: op1_09_in01 = reg_0957;
    110: op1_09_in01 = reg_0983;
    111: op1_09_in01 = reg_1325;
    112: op1_09_in01 = reg_0570;
    113: op1_09_in01 = reg_0448;
    114: op1_09_in01 = reg_0079;
    115: op1_09_in01 = reg_0421;
    116: op1_09_in01 = reg_0555;
    117: op1_09_in01 = reg_0630;
    40: op1_09_in01 = reg_0796;
    119: op1_09_in01 = reg_1244;
    120: op1_09_in01 = reg_1101;
    121: op1_09_in01 = reg_1071;
    122: op1_09_in01 = reg_1253;
    34: op1_09_in01 = reg_0140;
    124: op1_09_in01 = reg_1074;
    125: op1_09_in01 = reg_0583;
    126: op1_09_in01 = reg_0830;
    38: op1_09_in01 = reg_0740;
    128: op1_09_in01 = imem00_in[11:8];
    42: op1_09_in01 = reg_0120;
    129: op1_09_in01 = reg_0255;
    130: op1_09_in01 = reg_0130;
    131: op1_09_in01 = reg_0975;
    default: op1_09_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv01 = 1;
    73: op1_09_inv01 = 1;
    74: op1_09_inv01 = 1;
    75: op1_09_inv01 = 1;
    50: op1_09_inv01 = 1;
    76: op1_09_inv01 = 1;
    61: op1_09_inv01 = 1;
    78: op1_09_inv01 = 1;
    51: op1_09_inv01 = 1;
    79: op1_09_inv01 = 1;
    59: op1_09_inv01 = 1;
    88: op1_09_inv01 = 1;
    60: op1_09_inv01 = 1;
    62: op1_09_inv01 = 1;
    80: op1_09_inv01 = 1;
    48: op1_09_inv01 = 1;
    81: op1_09_inv01 = 1;
    52: op1_09_inv01 = 1;
    82: op1_09_inv01 = 1;
    83: op1_09_inv01 = 1;
    64: op1_09_inv01 = 1;
    84: op1_09_inv01 = 1;
    65: op1_09_inv01 = 1;
    66: op1_09_inv01 = 1;
    37: op1_09_inv01 = 1;
    91: op1_09_inv01 = 1;
    92: op1_09_inv01 = 1;
    94: op1_09_inv01 = 1;
    96: op1_09_inv01 = 1;
    99: op1_09_inv01 = 1;
    100: op1_09_inv01 = 1;
    103: op1_09_inv01 = 1;
    44: op1_09_inv01 = 1;
    104: op1_09_inv01 = 1;
    47: op1_09_inv01 = 1;
    107: op1_09_inv01 = 1;
    111: op1_09_inv01 = 1;
    116: op1_09_inv01 = 1;
    117: op1_09_inv01 = 1;
    40: op1_09_inv01 = 1;
    119: op1_09_inv01 = 1;
    126: op1_09_inv01 = 1;
    38: op1_09_inv01 = 1;
    128: op1_09_inv01 = 1;
    42: op1_09_inv01 = 1;
    129: op1_09_inv01 = 1;
    130: op1_09_inv01 = 1;
    default: op1_09_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in02 = reg_0334;
    53: op1_09_in02 = reg_0462;
    86: op1_09_in02 = reg_0227;
    55: op1_09_in02 = imem06_in[15:12];
    73: op1_09_in02 = reg_0866;
    63: op1_09_in02 = reg_0866;
    69: op1_09_in02 = reg_0327;
    49: op1_09_in02 = reg_0672;
    74: op1_09_in02 = reg_0702;
    54: op1_09_in02 = reg_0901;
    68: op1_09_in02 = reg_1092;
    75: op1_09_in02 = reg_1163;
    50: op1_09_in02 = reg_0171;
    56: op1_09_in02 = reg_0673;
    71: op1_09_in02 = reg_0841;
    87: op1_09_in02 = reg_1001;
    76: op1_09_in02 = reg_0301;
    61: op1_09_in02 = reg_0293;
    57: op1_09_in02 = reg_0966;
    77: op1_09_in02 = reg_0735;
    58: op1_09_in02 = reg_0119;
    78: op1_09_in02 = reg_1241;
    70: op1_09_in02 = reg_0232;
    51: op1_09_in02 = reg_0923;
    79: op1_09_in02 = reg_0868;
    59: op1_09_in02 = reg_0362;
    88: op1_09_in02 = reg_1063;
    60: op1_09_in02 = reg_0449;
    46: op1_09_in02 = imem05_in[11:8];
    62: op1_09_in02 = reg_0747;
    80: op1_09_in02 = reg_0207;
    48: op1_09_in02 = reg_0291;
    81: op1_09_in02 = reg_0608;
    52: op1_09_in02 = reg_0117;
    33: op1_09_in02 = reg_0361;
    82: op1_09_in02 = reg_1278;
    89: op1_09_in02 = reg_0380;
    83: op1_09_in02 = reg_0195;
    125: op1_09_in02 = reg_0195;
    64: op1_09_in02 = reg_1204;
    84: op1_09_in02 = reg_0250;
    85: op1_09_in02 = reg_0456;
    65: op1_09_in02 = reg_1301;
    90: op1_09_in02 = reg_0116;
    66: op1_09_in02 = reg_0600;
    37: op1_09_in02 = reg_0157;
    91: op1_09_in02 = reg_0501;
    67: op1_09_in02 = reg_0268;
    92: op1_09_in02 = reg_1101;
    93: op1_09_in02 = reg_0726;
    94: op1_09_in02 = reg_0638;
    95: op1_09_in02 = reg_0040;
    96: op1_09_in02 = reg_0926;
    106: op1_09_in02 = reg_0926;
    119: op1_09_in02 = reg_0926;
    97: op1_09_in02 = reg_0153;
    98: op1_09_in02 = reg_1258;
    99: op1_09_in02 = reg_0697;
    100: op1_09_in02 = reg_0806;
    101: op1_09_in02 = reg_1097;
    102: op1_09_in02 = reg_0241;
    103: op1_09_in02 = reg_1300;
    44: op1_09_in02 = reg_0598;
    104: op1_09_in02 = reg_0270;
    47: op1_09_in02 = reg_0152;
    105: op1_09_in02 = imem05_in[7:4];
    107: op1_09_in02 = reg_1491;
    108: op1_09_in02 = reg_1518;
    109: op1_09_in02 = reg_0107;
    110: op1_09_in02 = reg_0958;
    111: op1_09_in02 = reg_1280;
    112: op1_09_in02 = reg_0132;
    113: op1_09_in02 = reg_1009;
    114: op1_09_in02 = reg_0724;
    115: op1_09_in02 = reg_0599;
    116: op1_09_in02 = reg_1028;
    117: op1_09_in02 = reg_1181;
    118: op1_09_in02 = imem00_in[15:12];
    40: op1_09_in02 = reg_0795;
    120: op1_09_in02 = reg_0748;
    121: op1_09_in02 = imem02_in[15:12];
    122: op1_09_in02 = reg_0384;
    34: op1_09_in02 = imem07_in[7:4];
    123: op1_09_in02 = imem04_in[11:8];
    124: op1_09_in02 = reg_0900;
    126: op1_09_in02 = reg_0968;
    127: op1_09_in02 = reg_1279;
    38: op1_09_in02 = reg_0738;
    128: op1_09_in02 = reg_0959;
    42: op1_09_in02 = reg_0239;
    129: op1_09_in02 = reg_0168;
    130: op1_09_in02 = reg_0575;
    131: op1_09_in02 = reg_1493;
    default: op1_09_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv02 = 1;
    86: op1_09_inv02 = 1;
    55: op1_09_inv02 = 1;
    73: op1_09_inv02 = 1;
    69: op1_09_inv02 = 1;
    49: op1_09_inv02 = 1;
    74: op1_09_inv02 = 1;
    50: op1_09_inv02 = 1;
    56: op1_09_inv02 = 1;
    71: op1_09_inv02 = 1;
    76: op1_09_inv02 = 1;
    61: op1_09_inv02 = 1;
    57: op1_09_inv02 = 1;
    58: op1_09_inv02 = 1;
    78: op1_09_inv02 = 1;
    51: op1_09_inv02 = 1;
    59: op1_09_inv02 = 1;
    88: op1_09_inv02 = 1;
    62: op1_09_inv02 = 1;
    33: op1_09_inv02 = 1;
    82: op1_09_inv02 = 1;
    64: op1_09_inv02 = 1;
    84: op1_09_inv02 = 1;
    65: op1_09_inv02 = 1;
    66: op1_09_inv02 = 1;
    91: op1_09_inv02 = 1;
    67: op1_09_inv02 = 1;
    92: op1_09_inv02 = 1;
    93: op1_09_inv02 = 1;
    94: op1_09_inv02 = 1;
    99: op1_09_inv02 = 1;
    100: op1_09_inv02 = 1;
    101: op1_09_inv02 = 1;
    103: op1_09_inv02 = 1;
    104: op1_09_inv02 = 1;
    47: op1_09_inv02 = 1;
    106: op1_09_inv02 = 1;
    111: op1_09_inv02 = 1;
    112: op1_09_inv02 = 1;
    113: op1_09_inv02 = 1;
    114: op1_09_inv02 = 1;
    115: op1_09_inv02 = 1;
    117: op1_09_inv02 = 1;
    40: op1_09_inv02 = 1;
    119: op1_09_inv02 = 1;
    122: op1_09_inv02 = 1;
    127: op1_09_inv02 = 1;
    38: op1_09_inv02 = 1;
    130: op1_09_inv02 = 1;
    default: op1_09_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in03 = reg_1181;
    53: op1_09_in03 = reg_0978;
    86: op1_09_in03 = reg_0006;
    129: op1_09_in03 = reg_0006;
    55: op1_09_in03 = reg_0152;
    73: op1_09_in03 = reg_1281;
    79: op1_09_in03 = reg_1281;
    96: op1_09_in03 = reg_1281;
    69: op1_09_in03 = reg_0632;
    49: op1_09_in03 = imem07_in[7:4];
    74: op1_09_in03 = reg_0395;
    54: op1_09_in03 = reg_0868;
    68: op1_09_in03 = reg_0178;
    103: op1_09_in03 = reg_0178;
    75: op1_09_in03 = reg_0066;
    50: op1_09_in03 = reg_0289;
    56: op1_09_in03 = reg_0674;
    71: op1_09_in03 = reg_1241;
    82: op1_09_in03 = reg_1241;
    87: op1_09_in03 = reg_0783;
    76: op1_09_in03 = reg_1484;
    61: op1_09_in03 = reg_0221;
    57: op1_09_in03 = reg_0146;
    77: op1_09_in03 = reg_0204;
    58: op1_09_in03 = reg_0165;
    78: op1_09_in03 = imem00_in[11:8];
    70: op1_09_in03 = reg_1149;
    51: op1_09_in03 = reg_0169;
    59: op1_09_in03 = reg_0360;
    88: op1_09_in03 = reg_0216;
    60: op1_09_in03 = reg_1030;
    46: op1_09_in03 = reg_0540;
    62: op1_09_in03 = imem01_in[11:8];
    80: op1_09_in03 = reg_0193;
    48: op1_09_in03 = reg_0283;
    81: op1_09_in03 = reg_0588;
    52: op1_09_in03 = reg_0209;
    33: op1_09_in03 = reg_0052;
    63: op1_09_in03 = reg_1080;
    89: op1_09_in03 = reg_0381;
    83: op1_09_in03 = reg_1064;
    64: op1_09_in03 = reg_0046;
    84: op1_09_in03 = reg_1028;
    85: op1_09_in03 = reg_0276;
    65: op1_09_in03 = reg_1093;
    90: op1_09_in03 = reg_0714;
    66: op1_09_in03 = reg_1183;
    37: op1_09_in03 = reg_0140;
    91: op1_09_in03 = reg_0803;
    67: op1_09_in03 = reg_0192;
    92: op1_09_in03 = reg_1079;
    93: op1_09_in03 = reg_0402;
    94: op1_09_in03 = reg_0445;
    95: op1_09_in03 = reg_0859;
    97: op1_09_in03 = reg_0186;
    98: op1_09_in03 = reg_1083;
    99: op1_09_in03 = reg_1402;
    100: op1_09_in03 = reg_0804;
    101: op1_09_in03 = reg_0498;
    102: op1_09_in03 = reg_0798;
    44: op1_09_in03 = imem04_in[15:12];
    123: op1_09_in03 = imem04_in[15:12];
    104: op1_09_in03 = reg_0795;
    47: op1_09_in03 = reg_0215;
    105: op1_09_in03 = reg_0315;
    106: op1_09_in03 = reg_1101;
    107: op1_09_in03 = reg_0293;
    108: op1_09_in03 = reg_0314;
    109: op1_09_in03 = reg_0104;
    110: op1_09_in03 = reg_1278;
    111: op1_09_in03 = reg_1338;
    112: op1_09_in03 = reg_0419;
    113: op1_09_in03 = reg_0025;
    114: op1_09_in03 = reg_0403;
    115: op1_09_in03 = reg_1040;
    116: op1_09_in03 = reg_1459;
    117: op1_09_in03 = reg_1070;
    118: op1_09_in03 = reg_1244;
    40: op1_09_in03 = reg_0596;
    119: op1_09_in03 = reg_0866;
    120: op1_09_in03 = reg_1491;
    121: op1_09_in03 = reg_0877;
    122: op1_09_in03 = reg_0385;
    34: op1_09_in03 = reg_0284;
    124: op1_09_in03 = reg_0495;
    125: op1_09_in03 = reg_0214;
    126: op1_09_in03 = reg_0434;
    127: op1_09_in03 = reg_1490;
    38: op1_09_in03 = reg_0408;
    128: op1_09_in03 = reg_0926;
    42: op1_09_in03 = reg_0241;
    130: op1_09_in03 = reg_0864;
    131: op1_09_in03 = reg_1074;
    default: op1_09_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv03 = 1;
    53: op1_09_inv03 = 1;
    55: op1_09_inv03 = 1;
    69: op1_09_inv03 = 1;
    74: op1_09_inv03 = 1;
    68: op1_09_inv03 = 1;
    75: op1_09_inv03 = 1;
    56: op1_09_inv03 = 1;
    87: op1_09_inv03 = 1;
    76: op1_09_inv03 = 1;
    61: op1_09_inv03 = 1;
    57: op1_09_inv03 = 1;
    58: op1_09_inv03 = 1;
    78: op1_09_inv03 = 1;
    70: op1_09_inv03 = 1;
    59: op1_09_inv03 = 1;
    48: op1_09_inv03 = 1;
    81: op1_09_inv03 = 1;
    52: op1_09_inv03 = 1;
    33: op1_09_inv03 = 1;
    63: op1_09_inv03 = 1;
    82: op1_09_inv03 = 1;
    65: op1_09_inv03 = 1;
    37: op1_09_inv03 = 1;
    91: op1_09_inv03 = 1;
    103: op1_09_inv03 = 1;
    44: op1_09_inv03 = 1;
    47: op1_09_inv03 = 1;
    107: op1_09_inv03 = 1;
    108: op1_09_inv03 = 1;
    109: op1_09_inv03 = 1;
    111: op1_09_inv03 = 1;
    115: op1_09_inv03 = 1;
    116: op1_09_inv03 = 1;
    40: op1_09_inv03 = 1;
    122: op1_09_inv03 = 1;
    34: op1_09_inv03 = 1;
    123: op1_09_inv03 = 1;
    125: op1_09_inv03 = 1;
    126: op1_09_inv03 = 1;
    38: op1_09_inv03 = 1;
    128: op1_09_inv03 = 1;
    42: op1_09_inv03 = 1;
    default: op1_09_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in04 = reg_1402;
    53: op1_09_in04 = reg_1077;
    86: op1_09_in04 = reg_0233;
    55: op1_09_in04 = reg_0214;
    73: op1_09_in04 = reg_1080;
    69: op1_09_in04 = reg_0325;
    49: op1_09_in04 = reg_0774;
    74: op1_09_in04 = reg_0168;
    77: op1_09_in04 = reg_0168;
    54: op1_09_in04 = reg_0010;
    68: op1_09_in04 = reg_1208;
    75: op1_09_in04 = reg_0564;
    50: op1_09_in04 = reg_0460;
    56: op1_09_in04 = reg_0159;
    71: op1_09_in04 = reg_0806;
    120: op1_09_in04 = reg_0806;
    127: op1_09_in04 = reg_0806;
    87: op1_09_in04 = reg_1313;
    76: op1_09_in04 = reg_0576;
    61: op1_09_in04 = reg_0249;
    57: op1_09_in04 = reg_0385;
    58: op1_09_in04 = reg_0046;
    78: op1_09_in04 = reg_0803;
    70: op1_09_in04 = reg_0199;
    115: op1_09_in04 = reg_0199;
    51: op1_09_in04 = reg_0791;
    79: op1_09_in04 = reg_1277;
    59: op1_09_in04 = reg_0092;
    88: op1_09_in04 = reg_0541;
    60: op1_09_in04 = reg_0783;
    46: op1_09_in04 = reg_0450;
    62: op1_09_in04 = imem01_in[15:12];
    80: op1_09_in04 = reg_0751;
    48: op1_09_in04 = reg_0043;
    81: op1_09_in04 = reg_0934;
    52: op1_09_in04 = reg_0793;
    33: op1_09_in04 = reg_0085;
    63: op1_09_in04 = reg_1244;
    82: op1_09_in04 = reg_0580;
    94: op1_09_in04 = reg_0580;
    89: op1_09_in04 = reg_0307;
    83: op1_09_in04 = reg_0906;
    64: op1_09_in04 = reg_0212;
    84: op1_09_in04 = reg_1230;
    85: op1_09_in04 = reg_1260;
    65: op1_09_in04 = reg_1092;
    90: op1_09_in04 = reg_1302;
    66: op1_09_in04 = reg_1350;
    37: op1_09_in04 = reg_0664;
    91: op1_09_in04 = reg_0841;
    67: op1_09_in04 = reg_0120;
    92: op1_09_in04 = reg_1490;
    96: op1_09_in04 = reg_1490;
    93: op1_09_in04 = reg_0464;
    95: op1_09_in04 = reg_0752;
    97: op1_09_in04 = reg_1205;
    98: op1_09_in04 = reg_0500;
    99: op1_09_in04 = reg_0303;
    100: op1_09_in04 = reg_0615;
    101: op1_09_in04 = reg_0667;
    102: op1_09_in04 = reg_0612;
    103: op1_09_in04 = reg_0104;
    44: op1_09_in04 = reg_0305;
    104: op1_09_in04 = reg_0397;
    47: op1_09_in04 = imem07_in[11:8];
    105: op1_09_in04 = reg_0367;
    106: op1_09_in04 = reg_0613;
    107: op1_09_in04 = reg_1453;
    108: op1_09_in04 = reg_0597;
    109: op1_09_in04 = reg_0880;
    110: op1_09_in04 = reg_1491;
    111: op1_09_in04 = reg_1144;
    112: op1_09_in04 = reg_0289;
    113: op1_09_in04 = reg_0291;
    114: op1_09_in04 = imem01_in[3:0];
    116: op1_09_in04 = reg_1206;
    117: op1_09_in04 = reg_1514;
    118: op1_09_in04 = reg_1470;
    40: op1_09_in04 = reg_0341;
    119: op1_09_in04 = reg_0843;
    121: op1_09_in04 = reg_0423;
    122: op1_09_in04 = reg_0899;
    34: op1_09_in04 = reg_0441;
    123: op1_09_in04 = reg_0297;
    124: op1_09_in04 = reg_0436;
    125: op1_09_in04 = reg_0017;
    126: op1_09_in04 = reg_0438;
    38: op1_09_in04 = reg_0621;
    128: op1_09_in04 = reg_0725;
    42: op1_09_in04 = reg_0149;
    129: op1_09_in04 = reg_0377;
    130: op1_09_in04 = reg_0617;
    131: op1_09_in04 = reg_0900;
    default: op1_09_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv04 = 1;
    73: op1_09_inv04 = 1;
    49: op1_09_inv04 = 1;
    74: op1_09_inv04 = 1;
    54: op1_09_inv04 = 1;
    75: op1_09_inv04 = 1;
    56: op1_09_inv04 = 1;
    71: op1_09_inv04 = 1;
    87: op1_09_inv04 = 1;
    61: op1_09_inv04 = 1;
    57: op1_09_inv04 = 1;
    77: op1_09_inv04 = 1;
    58: op1_09_inv04 = 1;
    78: op1_09_inv04 = 1;
    79: op1_09_inv04 = 1;
    59: op1_09_inv04 = 1;
    88: op1_09_inv04 = 1;
    48: op1_09_inv04 = 1;
    52: op1_09_inv04 = 1;
    33: op1_09_inv04 = 1;
    63: op1_09_inv04 = 1;
    82: op1_09_inv04 = 1;
    83: op1_09_inv04 = 1;
    64: op1_09_inv04 = 1;
    84: op1_09_inv04 = 1;
    85: op1_09_inv04 = 1;
    65: op1_09_inv04 = 1;
    90: op1_09_inv04 = 1;
    66: op1_09_inv04 = 1;
    91: op1_09_inv04 = 1;
    67: op1_09_inv04 = 1;
    92: op1_09_inv04 = 1;
    93: op1_09_inv04 = 1;
    94: op1_09_inv04 = 1;
    96: op1_09_inv04 = 1;
    97: op1_09_inv04 = 1;
    98: op1_09_inv04 = 1;
    100: op1_09_inv04 = 1;
    101: op1_09_inv04 = 1;
    102: op1_09_inv04 = 1;
    103: op1_09_inv04 = 1;
    47: op1_09_inv04 = 1;
    105: op1_09_inv04 = 1;
    107: op1_09_inv04 = 1;
    109: op1_09_inv04 = 1;
    112: op1_09_inv04 = 1;
    114: op1_09_inv04 = 1;
    115: op1_09_inv04 = 1;
    117: op1_09_inv04 = 1;
    118: op1_09_inv04 = 1;
    40: op1_09_inv04 = 1;
    120: op1_09_inv04 = 1;
    121: op1_09_inv04 = 1;
    122: op1_09_inv04 = 1;
    123: op1_09_inv04 = 1;
    124: op1_09_inv04 = 1;
    125: op1_09_inv04 = 1;
    126: op1_09_inv04 = 1;
    127: op1_09_inv04 = 1;
    38: op1_09_inv04 = 1;
    129: op1_09_inv04 = 1;
    130: op1_09_inv04 = 1;
    default: op1_09_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in05 = reg_0541;
    103: op1_09_in05 = reg_0541;
    53: op1_09_in05 = reg_0412;
    86: op1_09_in05 = reg_0699;
    55: op1_09_in05 = reg_0162;
    73: op1_09_in05 = reg_0562;
    69: op1_09_in05 = reg_0276;
    121: op1_09_in05 = reg_0276;
    49: op1_09_in05 = reg_0738;
    74: op1_09_in05 = reg_0347;
    54: op1_09_in05 = reg_0486;
    68: op1_09_in05 = reg_0104;
    75: op1_09_in05 = reg_1403;
    50: op1_09_in05 = reg_0046;
    56: op1_09_in05 = reg_0158;
    71: op1_09_in05 = imem00_in[7:4];
    87: op1_09_in05 = reg_0190;
    76: op1_09_in05 = reg_0197;
    99: op1_09_in05 = reg_0197;
    61: op1_09_in05 = reg_0987;
    84: op1_09_in05 = reg_0987;
    57: op1_09_in05 = reg_0362;
    77: op1_09_in05 = reg_1169;
    58: op1_09_in05 = reg_0152;
    78: op1_09_in05 = reg_1028;
    70: op1_09_in05 = reg_1139;
    51: op1_09_in05 = reg_0465;
    79: op1_09_in05 = reg_1078;
    59: op1_09_in05 = reg_0724;
    88: op1_09_in05 = reg_0962;
    60: op1_09_in05 = reg_0192;
    46: op1_09_in05 = reg_0070;
    62: op1_09_in05 = reg_0242;
    80: op1_09_in05 = reg_1105;
    48: op1_09_in05 = reg_0010;
    81: op1_09_in05 = reg_1343;
    52: op1_09_in05 = imem05_in[15:12];
    33: op1_09_in05 = reg_0084;
    63: op1_09_in05 = reg_1242;
    82: op1_09_in05 = reg_0806;
    89: op1_09_in05 = reg_0473;
    83: op1_09_in05 = reg_1426;
    64: op1_09_in05 = reg_0215;
    85: op1_09_in05 = reg_0666;
    65: op1_09_in05 = reg_0113;
    90: op1_09_in05 = reg_1303;
    66: op1_09_in05 = reg_0139;
    37: op1_09_in05 = reg_0286;
    91: op1_09_in05 = reg_0615;
    67: op1_09_in05 = reg_1326;
    92: op1_09_in05 = reg_0613;
    93: op1_09_in05 = reg_0257;
    94: op1_09_in05 = reg_0555;
    95: op1_09_in05 = reg_1501;
    96: op1_09_in05 = reg_1489;
    97: op1_09_in05 = reg_0476;
    98: op1_09_in05 = reg_0094;
    100: op1_09_in05 = reg_0805;
    101: op1_09_in05 = reg_0225;
    102: op1_09_in05 = reg_0572;
    44: op1_09_in05 = reg_0487;
    104: op1_09_in05 = reg_0161;
    47: op1_09_in05 = reg_0704;
    105: op1_09_in05 = reg_0136;
    106: op1_09_in05 = reg_0841;
    110: op1_09_in05 = reg_0841;
    107: op1_09_in05 = reg_1459;
    108: op1_09_in05 = reg_1300;
    109: op1_09_in05 = reg_0350;
    111: op1_09_in05 = reg_0336;
    112: op1_09_in05 = reg_0213;
    113: op1_09_in05 = reg_0411;
    114: op1_09_in05 = reg_0895;
    115: op1_09_in05 = reg_1143;
    116: op1_09_in05 = reg_0961;
    117: op1_09_in05 = reg_0736;
    118: op1_09_in05 = reg_0926;
    40: op1_09_in05 = imem04_in[15:12];
    119: op1_09_in05 = reg_1278;
    120: op1_09_in05 = reg_1418;
    122: op1_09_in05 = reg_0901;
    34: op1_09_in05 = reg_0442;
    123: op1_09_in05 = reg_1200;
    124: op1_09_in05 = reg_0326;
    125: op1_09_in05 = reg_1170;
    126: op1_09_in05 = reg_1452;
    127: op1_09_in05 = reg_0616;
    38: op1_09_in05 = reg_0103;
    128: op1_09_in05 = reg_1277;
    42: op1_09_in05 = reg_0400;
    129: op1_09_in05 = imem03_in[7:4];
    130: op1_09_in05 = reg_0133;
    131: op1_09_in05 = reg_0778;
    default: op1_09_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    49: op1_09_inv05 = 1;
    74: op1_09_inv05 = 1;
    54: op1_09_inv05 = 1;
    50: op1_09_inv05 = 1;
    87: op1_09_inv05 = 1;
    76: op1_09_inv05 = 1;
    61: op1_09_inv05 = 1;
    57: op1_09_inv05 = 1;
    78: op1_09_inv05 = 1;
    51: op1_09_inv05 = 1;
    79: op1_09_inv05 = 1;
    59: op1_09_inv05 = 1;
    60: op1_09_inv05 = 1;
    62: op1_09_inv05 = 1;
    80: op1_09_inv05 = 1;
    48: op1_09_inv05 = 1;
    81: op1_09_inv05 = 1;
    33: op1_09_inv05 = 1;
    82: op1_09_inv05 = 1;
    89: op1_09_inv05 = 1;
    83: op1_09_inv05 = 1;
    84: op1_09_inv05 = 1;
    85: op1_09_inv05 = 1;
    65: op1_09_inv05 = 1;
    90: op1_09_inv05 = 1;
    66: op1_09_inv05 = 1;
    37: op1_09_inv05 = 1;
    91: op1_09_inv05 = 1;
    93: op1_09_inv05 = 1;
    94: op1_09_inv05 = 1;
    97: op1_09_inv05 = 1;
    98: op1_09_inv05 = 1;
    99: op1_09_inv05 = 1;
    100: op1_09_inv05 = 1;
    44: op1_09_inv05 = 1;
    104: op1_09_inv05 = 1;
    47: op1_09_inv05 = 1;
    105: op1_09_inv05 = 1;
    106: op1_09_inv05 = 1;
    107: op1_09_inv05 = 1;
    108: op1_09_inv05 = 1;
    112: op1_09_inv05 = 1;
    113: op1_09_inv05 = 1;
    116: op1_09_inv05 = 1;
    117: op1_09_inv05 = 1;
    40: op1_09_inv05 = 1;
    120: op1_09_inv05 = 1;
    121: op1_09_inv05 = 1;
    34: op1_09_inv05 = 1;
    123: op1_09_inv05 = 1;
    130: op1_09_inv05 = 1;
    131: op1_09_inv05 = 1;
    default: op1_09_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in06 = reg_0539;
    53: op1_09_in06 = reg_0796;
    86: op1_09_in06 = reg_0710;
    55: op1_09_in06 = reg_0229;
    73: op1_09_in06 = reg_0155;
    69: op1_09_in06 = reg_0280;
    49: op1_09_in06 = reg_0228;
    74: op1_09_in06 = reg_0176;
    54: op1_09_in06 = imem02_in[11:8];
    68: op1_09_in06 = reg_0481;
    75: op1_09_in06 = reg_0540;
    50: op1_09_in06 = imem07_in[7:4];
    56: op1_09_in06 = reg_0661;
    71: op1_09_in06 = imem00_in[11:8];
    87: op1_09_in06 = reg_1231;
    76: op1_09_in06 = reg_0492;
    61: op1_09_in06 = reg_1206;
    57: op1_09_in06 = reg_0047;
    77: op1_09_in06 = reg_0346;
    52: op1_09_in06 = reg_0346;
    58: op1_09_in06 = reg_0215;
    78: op1_09_in06 = reg_0821;
    107: op1_09_in06 = reg_0821;
    70: op1_09_in06 = reg_0638;
    51: op1_09_in06 = reg_0664;
    79: op1_09_in06 = reg_1489;
    59: op1_09_in06 = reg_0088;
    88: op1_09_in06 = reg_0377;
    60: op1_09_in06 = reg_0869;
    46: op1_09_in06 = reg_0418;
    62: op1_09_in06 = reg_0241;
    80: op1_09_in06 = reg_1426;
    48: op1_09_in06 = reg_0446;
    81: op1_09_in06 = reg_0255;
    33: op1_09_in06 = reg_0483;
    63: op1_09_in06 = reg_0293;
    82: op1_09_in06 = reg_0805;
    89: op1_09_in06 = reg_1000;
    83: op1_09_in06 = reg_0316;
    64: op1_09_in06 = reg_0214;
    84: op1_09_in06 = reg_1201;
    85: op1_09_in06 = reg_0474;
    65: op1_09_in06 = reg_0885;
    90: op1_09_in06 = reg_0194;
    66: op1_09_in06 = reg_0224;
    37: op1_09_in06 = reg_0366;
    91: op1_09_in06 = reg_0555;
    100: op1_09_in06 = reg_0555;
    127: op1_09_in06 = reg_0555;
    67: op1_09_in06 = reg_0160;
    92: op1_09_in06 = reg_0153;
    93: op1_09_in06 = reg_0120;
    94: op1_09_in06 = reg_0250;
    95: op1_09_in06 = reg_0635;
    96: op1_09_in06 = reg_0615;
    97: op1_09_in06 = reg_0928;
    120: op1_09_in06 = reg_0928;
    98: op1_09_in06 = reg_1147;
    99: op1_09_in06 = reg_0118;
    101: op1_09_in06 = reg_0309;
    102: op1_09_in06 = reg_0868;
    103: op1_09_in06 = reg_0218;
    44: op1_09_in06 = reg_0368;
    104: op1_09_in06 = reg_0192;
    47: op1_09_in06 = reg_0140;
    105: op1_09_in06 = reg_0347;
    106: op1_09_in06 = reg_0580;
    108: op1_09_in06 = reg_1199;
    109: op1_09_in06 = reg_0291;
    110: op1_09_in06 = reg_0640;
    111: op1_09_in06 = reg_0467;
    112: op1_09_in06 = reg_0017;
    113: op1_09_in06 = reg_1339;
    114: op1_09_in06 = reg_0447;
    115: op1_09_in06 = reg_0062;
    116: op1_09_in06 = reg_1417;
    117: op1_09_in06 = reg_0888;
    118: op1_09_in06 = reg_0866;
    40: op1_09_in06 = reg_0097;
    119: op1_09_in06 = reg_0803;
    121: op1_09_in06 = reg_0898;
    122: op1_09_in06 = reg_0080;
    34: op1_09_in06 = reg_0103;
    123: op1_09_in06 = reg_0281;
    124: op1_09_in06 = reg_0778;
    125: op1_09_in06 = reg_0169;
    126: op1_09_in06 = reg_0148;
    38: op1_09_in06 = reg_0361;
    128: op1_09_in06 = reg_0748;
    42: op1_09_in06 = reg_0384;
    129: op1_09_in06 = reg_0444;
    130: op1_09_in06 = reg_0670;
    131: op1_09_in06 = reg_0971;
    default: op1_09_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv06 = 1;
    86: op1_09_inv06 = 1;
    55: op1_09_inv06 = 1;
    73: op1_09_inv06 = 1;
    74: op1_09_inv06 = 1;
    75: op1_09_inv06 = 1;
    50: op1_09_inv06 = 1;
    71: op1_09_inv06 = 1;
    87: op1_09_inv06 = 1;
    76: op1_09_inv06 = 1;
    61: op1_09_inv06 = 1;
    57: op1_09_inv06 = 1;
    77: op1_09_inv06 = 1;
    78: op1_09_inv06 = 1;
    60: op1_09_inv06 = 1;
    46: op1_09_inv06 = 1;
    48: op1_09_inv06 = 1;
    81: op1_09_inv06 = 1;
    52: op1_09_inv06 = 1;
    82: op1_09_inv06 = 1;
    65: op1_09_inv06 = 1;
    66: op1_09_inv06 = 1;
    67: op1_09_inv06 = 1;
    97: op1_09_inv06 = 1;
    98: op1_09_inv06 = 1;
    101: op1_09_inv06 = 1;
    102: op1_09_inv06 = 1;
    103: op1_09_inv06 = 1;
    47: op1_09_inv06 = 1;
    105: op1_09_inv06 = 1;
    107: op1_09_inv06 = 1;
    108: op1_09_inv06 = 1;
    109: op1_09_inv06 = 1;
    110: op1_09_inv06 = 1;
    111: op1_09_inv06 = 1;
    112: op1_09_inv06 = 1;
    113: op1_09_inv06 = 1;
    118: op1_09_inv06 = 1;
    121: op1_09_inv06 = 1;
    34: op1_09_inv06 = 1;
    123: op1_09_inv06 = 1;
    125: op1_09_inv06 = 1;
    126: op1_09_inv06 = 1;
    127: op1_09_inv06 = 1;
    38: op1_09_inv06 = 1;
    42: op1_09_inv06 = 1;
    129: op1_09_inv06 = 1;
    130: op1_09_inv06 = 1;
    131: op1_09_inv06 = 1;
    default: op1_09_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in07 = reg_0937;
    53: op1_09_in07 = reg_0797;
    86: op1_09_in07 = reg_0179;
    129: op1_09_in07 = reg_0179;
    55: op1_09_in07 = reg_0821;
    73: op1_09_in07 = reg_0881;
    69: op1_09_in07 = reg_0312;
    49: op1_09_in07 = reg_0050;
    74: op1_09_in07 = reg_0992;
    54: op1_09_in07 = reg_0255;
    68: op1_09_in07 = imem03_in[3:0];
    75: op1_09_in07 = reg_0541;
    50: op1_09_in07 = reg_0998;
    56: op1_09_in07 = reg_0053;
    38: op1_09_in07 = reg_0053;
    71: op1_09_in07 = reg_1053;
    87: op1_09_in07 = reg_1199;
    76: op1_09_in07 = reg_0275;
    61: op1_09_in07 = reg_0460;
    57: op1_09_in07 = reg_0092;
    77: op1_09_in07 = reg_0333;
    58: op1_09_in07 = reg_0018;
    64: op1_09_in07 = reg_0018;
    78: op1_09_in07 = reg_0928;
    70: op1_09_in07 = reg_0144;
    51: op1_09_in07 = reg_0287;
    79: op1_09_in07 = reg_1244;
    59: op1_09_in07 = reg_0291;
    103: op1_09_in07 = reg_0291;
    88: op1_09_in07 = reg_0964;
    60: op1_09_in07 = reg_0827;
    46: op1_09_in07 = reg_0873;
    62: op1_09_in07 = reg_0743;
    80: op1_09_in07 = reg_1508;
    48: op1_09_in07 = reg_0629;
    81: op1_09_in07 = reg_0475;
    52: op1_09_in07 = reg_0392;
    63: op1_09_in07 = reg_0249;
    82: op1_09_in07 = reg_1471;
    89: op1_09_in07 = reg_0759;
    83: op1_09_in07 = reg_1509;
    84: op1_09_in07 = reg_0524;
    85: op1_09_in07 = reg_0054;
    65: op1_09_in07 = reg_0507;
    90: op1_09_in07 = reg_0141;
    66: op1_09_in07 = reg_0779;
    37: op1_09_in07 = reg_0442;
    91: op1_09_in07 = reg_0523;
    110: op1_09_in07 = reg_0523;
    67: op1_09_in07 = reg_0860;
    92: op1_09_in07 = reg_0554;
    93: op1_09_in07 = reg_0041;
    94: op1_09_in07 = reg_1418;
    95: op1_09_in07 = reg_0585;
    96: op1_09_in07 = reg_0580;
    97: op1_09_in07 = reg_0353;
    98: op1_09_in07 = reg_0421;
    99: op1_09_in07 = reg_0240;
    100: op1_09_in07 = reg_0640;
    101: op1_09_in07 = reg_0159;
    102: op1_09_in07 = reg_0091;
    44: op1_09_in07 = reg_0837;
    104: op1_09_in07 = reg_0782;
    47: op1_09_in07 = reg_0774;
    105: op1_09_in07 = reg_0184;
    106: op1_09_in07 = reg_0153;
    107: op1_09_in07 = reg_0476;
    116: op1_09_in07 = reg_0476;
    108: op1_09_in07 = reg_0885;
    109: op1_09_in07 = reg_0288;
    111: op1_09_in07 = reg_1369;
    112: op1_09_in07 = reg_1096;
    113: op1_09_in07 = reg_0336;
    114: op1_09_in07 = reg_0662;
    115: op1_09_in07 = reg_0236;
    117: op1_09_in07 = reg_0393;
    118: op1_09_in07 = reg_1081;
    40: op1_09_in07 = reg_0094;
    119: op1_09_in07 = reg_0805;
    120: op1_09_in07 = reg_0927;
    121: op1_09_in07 = reg_0776;
    122: op1_09_in07 = reg_0079;
    34: op1_09_in07 = reg_0361;
    123: op1_09_in07 = reg_0500;
    124: op1_09_in07 = reg_0307;
    125: op1_09_in07 = reg_0087;
    126: op1_09_in07 = reg_1032;
    127: op1_09_in07 = reg_1454;
    128: op1_09_in07 = reg_1487;
    42: op1_09_in07 = reg_0047;
    130: op1_09_in07 = reg_0729;
    131: op1_09_in07 = reg_0973;
    default: op1_09_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_09_inv07 = 1;
    55: op1_09_inv07 = 1;
    73: op1_09_inv07 = 1;
    69: op1_09_inv07 = 1;
    49: op1_09_inv07 = 1;
    74: op1_09_inv07 = 1;
    50: op1_09_inv07 = 1;
    56: op1_09_inv07 = 1;
    76: op1_09_inv07 = 1;
    57: op1_09_inv07 = 1;
    58: op1_09_inv07 = 1;
    70: op1_09_inv07 = 1;
    51: op1_09_inv07 = 1;
    79: op1_09_inv07 = 1;
    88: op1_09_inv07 = 1;
    46: op1_09_inv07 = 1;
    62: op1_09_inv07 = 1;
    48: op1_09_inv07 = 1;
    81: op1_09_inv07 = 1;
    52: op1_09_inv07 = 1;
    63: op1_09_inv07 = 1;
    82: op1_09_inv07 = 1;
    83: op1_09_inv07 = 1;
    65: op1_09_inv07 = 1;
    66: op1_09_inv07 = 1;
    91: op1_09_inv07 = 1;
    67: op1_09_inv07 = 1;
    93: op1_09_inv07 = 1;
    94: op1_09_inv07 = 1;
    95: op1_09_inv07 = 1;
    96: op1_09_inv07 = 1;
    99: op1_09_inv07 = 1;
    100: op1_09_inv07 = 1;
    44: op1_09_inv07 = 1;
    105: op1_09_inv07 = 1;
    106: op1_09_inv07 = 1;
    110: op1_09_inv07 = 1;
    111: op1_09_inv07 = 1;
    116: op1_09_inv07 = 1;
    117: op1_09_inv07 = 1;
    40: op1_09_inv07 = 1;
    119: op1_09_inv07 = 1;
    120: op1_09_inv07 = 1;
    121: op1_09_inv07 = 1;
    122: op1_09_inv07 = 1;
    123: op1_09_inv07 = 1;
    124: op1_09_inv07 = 1;
    125: op1_09_inv07 = 1;
    126: op1_09_inv07 = 1;
    38: op1_09_inv07 = 1;
    42: op1_09_inv07 = 1;
    default: op1_09_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in08 = reg_0163;
    53: op1_09_in08 = reg_0454;
    86: op1_09_in08 = reg_1425;
    55: op1_09_in08 = reg_1095;
    73: op1_09_in08 = reg_0353;
    69: op1_09_in08 = reg_0758;
    49: op1_09_in08 = reg_0052;
    74: op1_09_in08 = reg_1180;
    54: op1_09_in08 = reg_0629;
    68: op1_09_in08 = reg_0790;
    75: op1_09_in08 = reg_0303;
    50: op1_09_in08 = reg_0223;
    56: op1_09_in08 = reg_0085;
    71: op1_09_in08 = reg_0523;
    87: op1_09_in08 = reg_1092;
    76: op1_09_in08 = reg_1373;
    61: op1_09_in08 = reg_0459;
    57: op1_09_in08 = reg_0724;
    122: op1_09_in08 = reg_0724;
    77: op1_09_in08 = reg_0272;
    58: op1_09_in08 = reg_0022;
    78: op1_09_in08 = reg_0881;
    70: op1_09_in08 = reg_1314;
    51: op1_09_in08 = reg_0591;
    79: op1_09_in08 = reg_0613;
    59: op1_09_in08 = reg_0277;
    88: op1_09_in08 = reg_0957;
    60: op1_09_in08 = reg_0115;
    46: op1_09_in08 = reg_0872;
    62: op1_09_in08 = reg_1152;
    80: op1_09_in08 = reg_1326;
    48: op1_09_in08 = reg_0631;
    81: op1_09_in08 = reg_0495;
    52: op1_09_in08 = reg_0174;
    63: op1_09_in08 = reg_1201;
    82: op1_09_in08 = reg_1230;
    89: op1_09_in08 = reg_0573;
    83: op1_09_in08 = reg_0720;
    64: op1_09_in08 = reg_0230;
    84: op1_09_in08 = reg_0387;
    85: op1_09_in08 = reg_0972;
    131: op1_09_in08 = reg_0972;
    65: op1_09_in08 = reg_0425;
    90: op1_09_in08 = reg_0583;
    66: op1_09_in08 = reg_0664;
    37: op1_09_in08 = imem07_in[11:8];
    91: op1_09_in08 = reg_0221;
    67: op1_09_in08 = reg_0264;
    92: op1_09_in08 = reg_0640;
    93: op1_09_in08 = reg_1068;
    94: op1_09_in08 = reg_0928;
    95: op1_09_in08 = reg_0617;
    96: op1_09_in08 = reg_0616;
    97: op1_09_in08 = reg_0409;
    98: op1_09_in08 = reg_0407;
    99: op1_09_in08 = reg_0039;
    100: op1_09_in08 = reg_1052;
    101: op1_09_in08 = reg_0489;
    102: op1_09_in08 = reg_0899;
    103: op1_09_in08 = reg_0411;
    44: op1_09_in08 = reg_0337;
    104: op1_09_in08 = reg_0696;
    47: op1_09_in08 = reg_0031;
    105: op1_09_in08 = reg_0395;
    106: op1_09_in08 = reg_0554;
    107: op1_09_in08 = reg_0927;
    108: op1_09_in08 = reg_0707;
    109: op1_09_in08 = reg_1280;
    110: op1_09_in08 = reg_1453;
    111: op1_09_in08 = imem04_in[7:4];
    112: op1_09_in08 = reg_1183;
    113: op1_09_in08 = reg_0208;
    114: op1_09_in08 = imem02_in[15:12];
    115: op1_09_in08 = reg_0020;
    116: op1_09_in08 = reg_1393;
    117: op1_09_in08 = reg_0243;
    118: op1_09_in08 = reg_0725;
    40: op1_09_in08 = reg_0095;
    119: op1_09_in08 = reg_1027;
    120: op1_09_in08 = reg_0351;
    121: op1_09_in08 = reg_0326;
    34: op1_09_in08 = reg_0051;
    123: op1_09_in08 = reg_0406;
    124: op1_09_in08 = reg_0734;
    125: op1_09_in08 = reg_0394;
    126: op1_09_in08 = reg_0679;
    127: op1_09_in08 = reg_0155;
    38: op1_09_in08 = reg_0086;
    128: op1_09_in08 = reg_0806;
    42: op1_09_in08 = imem01_in[15:12];
    129: op1_09_in08 = reg_0706;
    130: op1_09_in08 = reg_0751;
    default: op1_09_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv08 = 1;
    86: op1_09_inv08 = 1;
    55: op1_09_inv08 = 1;
    69: op1_09_inv08 = 1;
    74: op1_09_inv08 = 1;
    54: op1_09_inv08 = 1;
    68: op1_09_inv08 = 1;
    56: op1_09_inv08 = 1;
    71: op1_09_inv08 = 1;
    76: op1_09_inv08 = 1;
    61: op1_09_inv08 = 1;
    57: op1_09_inv08 = 1;
    77: op1_09_inv08 = 1;
    70: op1_09_inv08 = 1;
    88: op1_09_inv08 = 1;
    60: op1_09_inv08 = 1;
    46: op1_09_inv08 = 1;
    80: op1_09_inv08 = 1;
    48: op1_09_inv08 = 1;
    52: op1_09_inv08 = 1;
    63: op1_09_inv08 = 1;
    82: op1_09_inv08 = 1;
    84: op1_09_inv08 = 1;
    85: op1_09_inv08 = 1;
    90: op1_09_inv08 = 1;
    37: op1_09_inv08 = 1;
    91: op1_09_inv08 = 1;
    67: op1_09_inv08 = 1;
    92: op1_09_inv08 = 1;
    93: op1_09_inv08 = 1;
    94: op1_09_inv08 = 1;
    95: op1_09_inv08 = 1;
    96: op1_09_inv08 = 1;
    97: op1_09_inv08 = 1;
    98: op1_09_inv08 = 1;
    100: op1_09_inv08 = 1;
    101: op1_09_inv08 = 1;
    103: op1_09_inv08 = 1;
    104: op1_09_inv08 = 1;
    105: op1_09_inv08 = 1;
    108: op1_09_inv08 = 1;
    111: op1_09_inv08 = 1;
    116: op1_09_inv08 = 1;
    117: op1_09_inv08 = 1;
    122: op1_09_inv08 = 1;
    34: op1_09_inv08 = 1;
    125: op1_09_inv08 = 1;
    126: op1_09_inv08 = 1;
    38: op1_09_inv08 = 1;
    128: op1_09_inv08 = 1;
    42: op1_09_inv08 = 1;
    default: op1_09_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in09 = reg_0450;
    53: op1_09_in09 = reg_0932;
    86: op1_09_in09 = reg_0823;
    89: op1_09_in09 = reg_0823;
    55: op1_09_in09 = imem07_in[11:8];
    73: op1_09_in09 = reg_0201;
    94: op1_09_in09 = reg_0201;
    69: op1_09_in09 = reg_0191;
    74: op1_09_in09 = reg_1403;
    54: op1_09_in09 = reg_0607;
    68: op1_09_in09 = reg_0427;
    75: op1_09_in09 = reg_0197;
    50: op1_09_in09 = reg_0225;
    56: op1_09_in09 = reg_0084;
    71: op1_09_in09 = reg_1027;
    87: op1_09_in09 = reg_0880;
    76: op1_09_in09 = reg_0118;
    61: op1_09_in09 = reg_1148;
    57: op1_09_in09 = reg_0902;
    77: op1_09_in09 = imem05_in[15:12];
    58: op1_09_in09 = reg_0490;
    78: op1_09_in09 = reg_0409;
    70: op1_09_in09 = reg_0627;
    51: op1_09_in09 = reg_0051;
    79: op1_09_in09 = reg_0580;
    59: op1_09_in09 = reg_0278;
    88: op1_09_in09 = reg_0558;
    60: op1_09_in09 = reg_0109;
    46: op1_09_in09 = reg_0130;
    62: op1_09_in09 = reg_0553;
    80: op1_09_in09 = reg_0860;
    48: op1_09_in09 = imem02_in[7:4];
    81: op1_09_in09 = reg_1207;
    52: op1_09_in09 = reg_0986;
    63: op1_09_in09 = reg_0492;
    82: op1_09_in09 = reg_1405;
    83: op1_09_in09 = reg_0780;
    64: op1_09_in09 = reg_0185;
    84: op1_09_in09 = reg_0058;
    85: op1_09_in09 = reg_0125;
    65: op1_09_in09 = reg_0458;
    90: op1_09_in09 = reg_1179;
    66: op1_09_in09 = reg_0102;
    37: op1_09_in09 = reg_0415;
    91: op1_09_in09 = reg_0485;
    119: op1_09_in09 = reg_0485;
    67: op1_09_in09 = reg_0116;
    92: op1_09_in09 = reg_0523;
    93: op1_09_in09 = reg_0447;
    95: op1_09_in09 = reg_0529;
    96: op1_09_in09 = reg_1052;
    106: op1_09_in09 = reg_1052;
    97: op1_09_in09 = reg_0134;
    98: op1_09_in09 = reg_1041;
    99: op1_09_in09 = reg_0265;
    100: op1_09_in09 = reg_1454;
    101: op1_09_in09 = reg_0620;
    102: op1_09_in09 = reg_0257;
    103: op1_09_in09 = imem04_in[11:8];
    44: op1_09_in09 = reg_0097;
    104: op1_09_in09 = reg_0984;
    47: op1_09_in09 = reg_0465;
    105: op1_09_in09 = reg_0700;
    107: op1_09_in09 = reg_0887;
    108: op1_09_in09 = reg_0378;
    109: op1_09_in09 = imem04_in[3:0];
    110: op1_09_in09 = reg_1459;
    111: op1_09_in09 = reg_1198;
    112: op1_09_in09 = reg_0140;
    113: op1_09_in09 = imem04_in[7:4];
    114: op1_09_in09 = reg_0889;
    115: op1_09_in09 = reg_0708;
    116: op1_09_in09 = reg_0410;
    117: op1_09_in09 = reg_1346;
    118: op1_09_in09 = reg_0843;
    40: op1_09_in09 = reg_0237;
    120: op1_09_in09 = reg_0352;
    121: op1_09_in09 = reg_0106;
    122: op1_09_in09 = reg_0162;
    34: op1_09_in09 = reg_0052;
    123: op1_09_in09 = reg_0599;
    124: op1_09_in09 = reg_0989;
    125: op1_09_in09 = reg_1095;
    126: op1_09_in09 = reg_0362;
    127: op1_09_in09 = reg_0524;
    38: op1_09_in09 = reg_0520;
    128: op1_09_in09 = reg_0248;
    42: op1_09_in09 = reg_0080;
    129: op1_09_in09 = reg_0220;
    130: op1_09_in09 = reg_1323;
    131: op1_09_in09 = reg_1458;
    default: op1_09_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv09 = 1;
    73: op1_09_inv09 = 1;
    69: op1_09_inv09 = 1;
    54: op1_09_inv09 = 1;
    68: op1_09_inv09 = 1;
    75: op1_09_inv09 = 1;
    50: op1_09_inv09 = 1;
    71: op1_09_inv09 = 1;
    58: op1_09_inv09 = 1;
    78: op1_09_inv09 = 1;
    70: op1_09_inv09 = 1;
    46: op1_09_inv09 = 1;
    62: op1_09_inv09 = 1;
    80: op1_09_inv09 = 1;
    48: op1_09_inv09 = 1;
    81: op1_09_inv09 = 1;
    52: op1_09_inv09 = 1;
    89: op1_09_inv09 = 1;
    64: op1_09_inv09 = 1;
    84: op1_09_inv09 = 1;
    66: op1_09_inv09 = 1;
    37: op1_09_inv09 = 1;
    96: op1_09_inv09 = 1;
    97: op1_09_inv09 = 1;
    98: op1_09_inv09 = 1;
    99: op1_09_inv09 = 1;
    100: op1_09_inv09 = 1;
    101: op1_09_inv09 = 1;
    102: op1_09_inv09 = 1;
    103: op1_09_inv09 = 1;
    104: op1_09_inv09 = 1;
    47: op1_09_inv09 = 1;
    105: op1_09_inv09 = 1;
    107: op1_09_inv09 = 1;
    110: op1_09_inv09 = 1;
    114: op1_09_inv09 = 1;
    115: op1_09_inv09 = 1;
    116: op1_09_inv09 = 1;
    117: op1_09_inv09 = 1;
    118: op1_09_inv09 = 1;
    119: op1_09_inv09 = 1;
    121: op1_09_inv09 = 1;
    124: op1_09_inv09 = 1;
    126: op1_09_inv09 = 1;
    38: op1_09_inv09 = 1;
    130: op1_09_inv09 = 1;
    default: op1_09_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in10 = reg_0477;
    53: op1_09_in10 = reg_0452;
    86: op1_09_in10 = reg_0144;
    55: op1_09_in10 = imem07_in[15:12];
    73: op1_09_in10 = reg_0189;
    120: op1_09_in10 = reg_0189;
    69: op1_09_in10 = reg_0677;
    74: op1_09_in10 = reg_1401;
    54: op1_09_in10 = reg_0455;
    68: op1_09_in10 = reg_0411;
    75: op1_09_in10 = reg_0601;
    50: op1_09_in10 = reg_0226;
    56: op1_09_in10 = reg_0518;
    71: op1_09_in10 = reg_1453;
    100: op1_09_in10 = reg_1453;
    106: op1_09_in10 = reg_1453;
    87: op1_09_in10 = imem03_in[3:0];
    76: op1_09_in10 = reg_1348;
    61: op1_09_in10 = reg_0886;
    107: op1_09_in10 = reg_0886;
    57: op1_09_in10 = reg_0291;
    77: op1_09_in10 = reg_0183;
    58: op1_09_in10 = reg_0668;
    93: op1_09_in10 = reg_0668;
    78: op1_09_in10 = reg_0203;
    70: op1_09_in10 = reg_0597;
    51: op1_09_in10 = reg_0053;
    79: op1_09_in10 = reg_0293;
    59: op1_09_in10 = reg_0662;
    88: op1_09_in10 = reg_0882;
    60: op1_09_in10 = reg_0194;
    46: op1_09_in10 = reg_0780;
    62: op1_09_in10 = reg_0982;
    80: op1_09_in10 = reg_0863;
    48: op1_09_in10 = reg_0587;
    81: op1_09_in10 = reg_0429;
    52: op1_09_in10 = reg_0565;
    63: op1_09_in10 = reg_1148;
    82: op1_09_in10 = reg_1393;
    89: op1_09_in10 = reg_0954;
    83: op1_09_in10 = reg_1302;
    64: op1_09_in10 = reg_0496;
    121: op1_09_in10 = reg_0496;
    84: op1_09_in10 = reg_1324;
    85: op1_09_in10 = reg_0112;
    65: op1_09_in10 = reg_0582;
    90: op1_09_in10 = reg_0023;
    66: op1_09_in10 = reg_0103;
    37: op1_09_in10 = reg_0621;
    91: op1_09_in10 = reg_1201;
    110: op1_09_in10 = reg_1201;
    67: op1_09_in10 = reg_0714;
    92: op1_09_in10 = reg_1230;
    94: op1_09_in10 = reg_0440;
    95: op1_09_in10 = reg_0571;
    96: op1_09_in10 = reg_0221;
    97: op1_09_in10 = reg_0073;
    98: op1_09_in10 = reg_1040;
    99: op1_09_in10 = reg_0784;
    101: op1_09_in10 = reg_0321;
    102: op1_09_in10 = reg_0043;
    103: op1_09_in10 = reg_0493;
    113: op1_09_in10 = reg_0493;
    44: op1_09_in10 = reg_0164;
    104: op1_09_in10 = reg_1467;
    47: op1_09_in10 = reg_0663;
    105: op1_09_in10 = reg_0996;
    108: op1_09_in10 = reg_0336;
    109: op1_09_in10 = imem04_in[7:4];
    111: op1_09_in10 = reg_0421;
    112: op1_09_in10 = reg_0921;
    114: op1_09_in10 = reg_0327;
    115: op1_09_in10 = reg_0538;
    116: op1_09_in10 = reg_0058;
    117: op1_09_in10 = reg_0861;
    118: op1_09_in10 = reg_1281;
    40: op1_09_in10 = reg_0181;
    119: op1_09_in10 = reg_0961;
    122: op1_09_in10 = reg_0041;
    34: op1_09_in10 = reg_0087;
    123: op1_09_in10 = reg_0320;
    124: op1_09_in10 = reg_0220;
    125: op1_09_in10 = reg_0922;
    126: op1_09_in10 = reg_0365;
    127: op1_09_in10 = reg_0405;
    128: op1_09_in10 = reg_1102;
    42: op1_09_in10 = reg_0290;
    129: op1_09_in10 = reg_0177;
    130: op1_09_in10 = reg_1505;
    131: op1_09_in10 = reg_1455;
    default: op1_09_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv10 = 1;
    73: op1_09_inv10 = 1;
    69: op1_09_inv10 = 1;
    74: op1_09_inv10 = 1;
    54: op1_09_inv10 = 1;
    68: op1_09_inv10 = 1;
    75: op1_09_inv10 = 1;
    50: op1_09_inv10 = 1;
    56: op1_09_inv10 = 1;
    71: op1_09_inv10 = 1;
    87: op1_09_inv10 = 1;
    76: op1_09_inv10 = 1;
    78: op1_09_inv10 = 1;
    51: op1_09_inv10 = 1;
    79: op1_09_inv10 = 1;
    88: op1_09_inv10 = 1;
    60: op1_09_inv10 = 1;
    46: op1_09_inv10 = 1;
    62: op1_09_inv10 = 1;
    80: op1_09_inv10 = 1;
    52: op1_09_inv10 = 1;
    82: op1_09_inv10 = 1;
    83: op1_09_inv10 = 1;
    84: op1_09_inv10 = 1;
    90: op1_09_inv10 = 1;
    37: op1_09_inv10 = 1;
    67: op1_09_inv10 = 1;
    94: op1_09_inv10 = 1;
    98: op1_09_inv10 = 1;
    99: op1_09_inv10 = 1;
    101: op1_09_inv10 = 1;
    103: op1_09_inv10 = 1;
    104: op1_09_inv10 = 1;
    106: op1_09_inv10 = 1;
    108: op1_09_inv10 = 1;
    110: op1_09_inv10 = 1;
    113: op1_09_inv10 = 1;
    116: op1_09_inv10 = 1;
    40: op1_09_inv10 = 1;
    121: op1_09_inv10 = 1;
    34: op1_09_inv10 = 1;
    123: op1_09_inv10 = 1;
    125: op1_09_inv10 = 1;
    42: op1_09_inv10 = 1;
    130: op1_09_inv10 = 1;
    131: op1_09_inv10 = 1;
    default: op1_09_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in11 = reg_0367;
    53: op1_09_in11 = reg_0369;
    86: op1_09_in11 = reg_0180;
    55: op1_09_in11 = reg_0225;
    73: op1_09_in11 = reg_0416;
    69: op1_09_in11 = reg_0216;
    74: op1_09_in11 = reg_0541;
    54: op1_09_in11 = reg_0587;
    68: op1_09_in11 = reg_0341;
    75: op1_09_in11 = reg_0130;
    50: op1_09_in11 = reg_0245;
    56: op1_09_in11 = reg_0483;
    34: op1_09_in11 = reg_0483;
    71: op1_09_in11 = reg_1230;
    87: op1_09_in11 = reg_0481;
    76: op1_09_in11 = reg_0797;
    61: op1_09_in11 = reg_0641;
    57: op1_09_in11 = reg_0662;
    77: op1_09_in11 = reg_0418;
    58: op1_09_in11 = reg_0893;
    78: op1_09_in11 = reg_0073;
    70: op1_09_in11 = reg_1300;
    51: op1_09_in11 = reg_0085;
    79: op1_09_in11 = reg_0476;
    59: op1_09_in11 = reg_0699;
    88: op1_09_in11 = reg_0218;
    60: op1_09_in11 = reg_0585;
    46: op1_09_in11 = reg_0192;
    62: op1_09_in11 = reg_0966;
    80: op1_09_in11 = reg_0116;
    48: op1_09_in11 = reg_0563;
    81: op1_09_in11 = reg_0776;
    52: op1_09_in11 = reg_0566;
    63: op1_09_in11 = reg_0927;
    82: op1_09_in11 = reg_0202;
    89: op1_09_in11 = reg_0597;
    83: op1_09_in11 = reg_0622;
    64: op1_09_in11 = reg_0922;
    84: op1_09_in11 = reg_0027;
    85: op1_09_in11 = reg_0105;
    65: op1_09_in11 = reg_0975;
    90: op1_09_in11 = reg_0215;
    66: op1_09_in11 = reg_0100;
    37: op1_09_in11 = reg_0228;
    101: op1_09_in11 = reg_0228;
    91: op1_09_in11 = reg_1432;
    67: op1_09_in11 = reg_0636;
    92: op1_09_in11 = reg_0524;
    93: op1_09_in11 = reg_0456;
    94: op1_09_in11 = reg_0388;
    95: op1_09_in11 = reg_0569;
    96: op1_09_in11 = reg_0485;
    97: op1_09_in11 = reg_0060;
    98: op1_09_in11 = reg_0320;
    99: op1_09_in11 = imem06_in[7:4];
    100: op1_09_in11 = reg_0987;
    102: op1_09_in11 = reg_0041;
    103: op1_09_in11 = reg_0264;
    44: op1_09_in11 = reg_0181;
    104: op1_09_in11 = reg_0860;
    47: op1_09_in11 = reg_0664;
    105: op1_09_in11 = reg_0649;
    106: op1_09_in11 = reg_1205;
    107: op1_09_in11 = reg_0410;
    120: op1_09_in11 = reg_0410;
    108: op1_09_in11 = reg_0467;
    109: op1_09_in11 = reg_0507;
    124: op1_09_in11 = reg_0507;
    110: op1_09_in11 = reg_0351;
    111: op1_09_in11 = reg_0598;
    112: op1_09_in11 = reg_0465;
    113: op1_09_in11 = reg_1203;
    114: op1_09_in11 = reg_0008;
    115: op1_09_in11 = reg_0579;
    116: op1_09_in11 = reg_1322;
    117: op1_09_in11 = reg_0317;
    118: op1_09_in11 = reg_1278;
    40: op1_09_in11 = reg_0117;
    119: op1_09_in11 = reg_1417;
    121: op1_09_in11 = reg_0745;
    122: op1_09_in11 = reg_0010;
    123: op1_09_in11 = reg_0452;
    125: op1_09_in11 = reg_1350;
    126: op1_09_in11 = reg_0727;
    127: op1_09_in11 = reg_0058;
    128: op1_09_in11 = reg_0640;
    42: op1_09_in11 = reg_0042;
    129: op1_09_in11 = reg_0198;
    130: op1_09_in11 = reg_1504;
    131: op1_09_in11 = reg_0128;
    default: op1_09_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv11 = 1;
    86: op1_09_inv11 = 1;
    54: op1_09_inv11 = 1;
    76: op1_09_inv11 = 1;
    77: op1_09_inv11 = 1;
    78: op1_09_inv11 = 1;
    59: op1_09_inv11 = 1;
    62: op1_09_inv11 = 1;
    80: op1_09_inv11 = 1;
    52: op1_09_inv11 = 1;
    84: op1_09_inv11 = 1;
    85: op1_09_inv11 = 1;
    65: op1_09_inv11 = 1;
    90: op1_09_inv11 = 1;
    37: op1_09_inv11 = 1;
    91: op1_09_inv11 = 1;
    67: op1_09_inv11 = 1;
    92: op1_09_inv11 = 1;
    93: op1_09_inv11 = 1;
    95: op1_09_inv11 = 1;
    96: op1_09_inv11 = 1;
    97: op1_09_inv11 = 1;
    99: op1_09_inv11 = 1;
    100: op1_09_inv11 = 1;
    101: op1_09_inv11 = 1;
    102: op1_09_inv11 = 1;
    44: op1_09_inv11 = 1;
    104: op1_09_inv11 = 1;
    112: op1_09_inv11 = 1;
    116: op1_09_inv11 = 1;
    117: op1_09_inv11 = 1;
    118: op1_09_inv11 = 1;
    40: op1_09_inv11 = 1;
    120: op1_09_inv11 = 1;
    121: op1_09_inv11 = 1;
    34: op1_09_inv11 = 1;
    124: op1_09_inv11 = 1;
    125: op1_09_inv11 = 1;
    127: op1_09_inv11 = 1;
    131: op1_09_inv11 = 1;
    default: op1_09_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in12 = reg_0303;
    53: op1_09_in12 = reg_0262;
    86: op1_09_in12 = reg_0954;
    55: op1_09_in12 = reg_0704;
    73: op1_09_in12 = reg_0409;
    69: op1_09_in12 = reg_0830;
    74: op1_09_in12 = reg_0939;
    54: op1_09_in12 = reg_0532;
    68: op1_09_in12 = reg_1339;
    75: op1_09_in12 = reg_0631;
    50: op1_09_in12 = reg_0324;
    71: op1_09_in12 = reg_1205;
    87: op1_09_in12 = reg_1139;
    76: op1_09_in12 = reg_0754;
    61: op1_09_in12 = reg_0642;
    63: op1_09_in12 = reg_0642;
    57: op1_09_in12 = reg_0699;
    77: op1_09_in12 = reg_0302;
    58: op1_09_in12 = reg_0672;
    78: op1_09_in12 = reg_0059;
    70: op1_09_in12 = reg_0558;
    51: op1_09_in12 = reg_0518;
    79: op1_09_in12 = reg_0928;
    59: op1_09_in12 = reg_0744;
    88: op1_09_in12 = reg_1325;
    60: op1_09_in12 = reg_0345;
    83: op1_09_in12 = reg_0345;
    46: op1_09_in12 = reg_0929;
    62: op1_09_in12 = reg_0430;
    80: op1_09_in12 = reg_0110;
    48: op1_09_in12 = reg_0562;
    81: op1_09_in12 = reg_0778;
    52: op1_09_in12 = reg_0334;
    82: op1_09_in12 = reg_0351;
    89: op1_09_in12 = reg_1301;
    64: op1_09_in12 = reg_0924;
    84: op1_09_in12 = reg_1034;
    85: op1_09_in12 = reg_0629;
    65: op1_09_in12 = reg_1369;
    90: op1_09_in12 = imem07_in[11:8];
    66: op1_09_in12 = reg_0028;
    37: op1_09_in12 = reg_0050;
    101: op1_09_in12 = reg_0050;
    91: op1_09_in12 = reg_0887;
    119: op1_09_in12 = reg_0887;
    67: op1_09_in12 = reg_0398;
    92: op1_09_in12 = reg_0440;
    93: op1_09_in12 = reg_0455;
    94: op1_09_in12 = reg_0058;
    95: op1_09_in12 = reg_0419;
    96: op1_09_in12 = reg_0476;
    97: op1_09_in12 = reg_1322;
    107: op1_09_in12 = reg_1322;
    98: op1_09_in12 = reg_0452;
    99: op1_09_in12 = reg_0906;
    100: op1_09_in12 = reg_1201;
    102: op1_09_in12 = reg_0456;
    103: op1_09_in12 = reg_0694;
    44: op1_09_in12 = reg_0117;
    104: op1_09_in12 = reg_0752;
    47: op1_09_in12 = reg_0287;
    105: op1_09_in12 = reg_0174;
    106: op1_09_in12 = reg_0821;
    108: op1_09_in12 = reg_1372;
    109: op1_09_in12 = reg_0336;
    110: op1_09_in12 = reg_0387;
    111: op1_09_in12 = reg_1065;
    112: op1_09_in12 = reg_0029;
    113: op1_09_in12 = reg_1040;
    114: op1_09_in12 = reg_0845;
    115: op1_09_in12 = reg_0136;
    116: op1_09_in12 = reg_0089;
    117: op1_09_in12 = reg_0014;
    118: op1_09_in12 = reg_1489;
    40: op1_09_in12 = reg_0211;
    120: op1_09_in12 = reg_0075;
    121: op1_09_in12 = reg_0711;
    122: op1_09_in12 = reg_0662;
    123: op1_09_in12 = reg_1312;
    124: op1_09_in12 = reg_1495;
    125: op1_09_in12 = reg_0366;
    126: op1_09_in12 = reg_0400;
    127: op1_09_in12 = reg_0122;
    128: op1_09_in12 = reg_1027;
    42: op1_09_in12 = reg_0044;
    129: op1_09_in12 = reg_0847;
    130: op1_09_in12 = reg_0265;
    131: op1_09_in12 = reg_0111;
    default: op1_09_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv12 = 1;
    86: op1_09_inv12 = 1;
    55: op1_09_inv12 = 1;
    73: op1_09_inv12 = 1;
    74: op1_09_inv12 = 1;
    68: op1_09_inv12 = 1;
    75: op1_09_inv12 = 1;
    50: op1_09_inv12 = 1;
    71: op1_09_inv12 = 1;
    57: op1_09_inv12 = 1;
    77: op1_09_inv12 = 1;
    58: op1_09_inv12 = 1;
    78: op1_09_inv12 = 1;
    70: op1_09_inv12 = 1;
    51: op1_09_inv12 = 1;
    79: op1_09_inv12 = 1;
    46: op1_09_inv12 = 1;
    62: op1_09_inv12 = 1;
    52: op1_09_inv12 = 1;
    89: op1_09_inv12 = 1;
    64: op1_09_inv12 = 1;
    85: op1_09_inv12 = 1;
    66: op1_09_inv12 = 1;
    37: op1_09_inv12 = 1;
    91: op1_09_inv12 = 1;
    67: op1_09_inv12 = 1;
    92: op1_09_inv12 = 1;
    93: op1_09_inv12 = 1;
    95: op1_09_inv12 = 1;
    99: op1_09_inv12 = 1;
    101: op1_09_inv12 = 1;
    44: op1_09_inv12 = 1;
    104: op1_09_inv12 = 1;
    47: op1_09_inv12 = 1;
    109: op1_09_inv12 = 1;
    110: op1_09_inv12 = 1;
    112: op1_09_inv12 = 1;
    113: op1_09_inv12 = 1;
    117: op1_09_inv12 = 1;
    40: op1_09_inv12 = 1;
    120: op1_09_inv12 = 1;
    121: op1_09_inv12 = 1;
    125: op1_09_inv12 = 1;
    42: op1_09_inv12 = 1;
    129: op1_09_inv12 = 1;
    default: op1_09_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in13 = reg_0300;
    53: op1_09_in13 = reg_0837;
    86: op1_09_in13 = reg_0220;
    55: op1_09_in13 = reg_0324;
    73: op1_09_in13 = reg_0073;
    69: op1_09_in13 = reg_0707;
    74: op1_09_in13 = reg_0938;
    54: op1_09_in13 = reg_0531;
    68: op1_09_in13 = reg_1258;
    75: op1_09_in13 = reg_0449;
    50: op1_09_in13 = reg_0867;
    71: op1_09_in13 = reg_0524;
    87: op1_09_in13 = reg_1280;
    76: op1_09_in13 = reg_0780;
    61: op1_09_in13 = reg_0189;
    106: op1_09_in13 = reg_0189;
    57: op1_09_in13 = reg_0254;
    77: op1_09_in13 = reg_0301;
    58: op1_09_in13 = reg_0158;
    78: op1_09_in13 = reg_0005;
    107: op1_09_in13 = reg_0005;
    70: op1_09_in13 = reg_0525;
    79: op1_09_in13 = reg_0881;
    59: op1_09_in13 = reg_0255;
    88: op1_09_in13 = reg_0443;
    60: op1_09_in13 = reg_1225;
    46: op1_09_in13 = reg_0160;
    62: op1_09_in13 = reg_0727;
    80: op1_09_in13 = reg_0109;
    48: op1_09_in13 = reg_0532;
    81: op1_09_in13 = reg_1458;
    52: op1_09_in13 = reg_0540;
    63: op1_09_in13 = reg_0722;
    82: op1_09_in13 = reg_0075;
    89: op1_09_in13 = reg_0113;
    83: op1_09_in13 = reg_0132;
    64: op1_09_in13 = reg_0741;
    84: op1_09_in13 = reg_1290;
    85: op1_09_in13 = reg_0380;
    65: op1_09_in13 = reg_1203;
    90: op1_09_in13 = reg_0394;
    66: op1_09_in13 = reg_0050;
    37: op1_09_in13 = reg_0004;
    91: op1_09_in13 = reg_0351;
    67: op1_09_in13 = reg_0569;
    92: op1_09_in13 = reg_0410;
    93: op1_09_in13 = reg_0055;
    94: op1_09_in13 = reg_1100;
    95: op1_09_in13 = reg_0269;
    96: op1_09_in13 = reg_0886;
    97: op1_09_in13 = reg_0355;
    98: op1_09_in13 = reg_0342;
    111: op1_09_in13 = reg_0342;
    99: op1_09_in13 = reg_0905;
    100: op1_09_in13 = reg_1205;
    101: op1_09_in13 = reg_0003;
    102: op1_09_in13 = reg_0608;
    103: op1_09_in13 = reg_0281;
    44: op1_09_in13 = reg_0211;
    104: op1_09_in13 = reg_1501;
    47: op1_09_in13 = reg_0415;
    105: op1_09_in13 = reg_0066;
    108: op1_09_in13 = reg_1369;
    109: op1_09_in13 = reg_1383;
    110: op1_09_in13 = reg_0072;
    112: op1_09_in13 = reg_0442;
    113: op1_09_in13 = reg_0454;
    114: op1_09_in13 = reg_1018;
    115: op1_09_in13 = reg_0333;
    116: op1_09_in13 = reg_0723;
    117: op1_09_in13 = reg_0565;
    118: op1_09_in13 = reg_1487;
    40: op1_09_in13 = reg_0064;
    119: op1_09_in13 = reg_0431;
    120: op1_09_in13 = reg_1322;
    121: op1_09_in13 = reg_1078;
    122: op1_09_in13 = imem02_in[3:0];
    123: op1_09_in13 = reg_0256;
    124: op1_09_in13 = reg_0965;
    125: op1_09_in13 = reg_0437;
    126: op1_09_in13 = reg_0724;
    127: op1_09_in13 = reg_0089;
    128: op1_09_in13 = reg_0249;
    42: op1_09_in13 = reg_0486;
    129: op1_09_in13 = reg_0556;
    130: op1_09_in13 = reg_1302;
    131: op1_09_in13 = reg_0876;
    default: op1_09_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_09_inv13 = 1;
    54: op1_09_inv13 = 1;
    75: op1_09_inv13 = 1;
    50: op1_09_inv13 = 1;
    61: op1_09_inv13 = 1;
    57: op1_09_inv13 = 1;
    77: op1_09_inv13 = 1;
    58: op1_09_inv13 = 1;
    78: op1_09_inv13 = 1;
    70: op1_09_inv13 = 1;
    79: op1_09_inv13 = 1;
    88: op1_09_inv13 = 1;
    46: op1_09_inv13 = 1;
    80: op1_09_inv13 = 1;
    81: op1_09_inv13 = 1;
    64: op1_09_inv13 = 1;
    84: op1_09_inv13 = 1;
    65: op1_09_inv13 = 1;
    66: op1_09_inv13 = 1;
    37: op1_09_inv13 = 1;
    67: op1_09_inv13 = 1;
    92: op1_09_inv13 = 1;
    96: op1_09_inv13 = 1;
    97: op1_09_inv13 = 1;
    98: op1_09_inv13 = 1;
    99: op1_09_inv13 = 1;
    100: op1_09_inv13 = 1;
    102: op1_09_inv13 = 1;
    103: op1_09_inv13 = 1;
    44: op1_09_inv13 = 1;
    104: op1_09_inv13 = 1;
    47: op1_09_inv13 = 1;
    106: op1_09_inv13 = 1;
    108: op1_09_inv13 = 1;
    109: op1_09_inv13 = 1;
    110: op1_09_inv13 = 1;
    113: op1_09_inv13 = 1;
    114: op1_09_inv13 = 1;
    115: op1_09_inv13 = 1;
    116: op1_09_inv13 = 1;
    118: op1_09_inv13 = 1;
    40: op1_09_inv13 = 1;
    122: op1_09_inv13 = 1;
    123: op1_09_inv13 = 1;
    125: op1_09_inv13 = 1;
    126: op1_09_inv13 = 1;
    127: op1_09_inv13 = 1;
    129: op1_09_inv13 = 1;
    130: op1_09_inv13 = 1;
    131: op1_09_inv13 = 1;
    default: op1_09_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in14 = reg_0197;
    53: op1_09_in14 = reg_0835;
    86: op1_09_in14 = reg_0246;
    55: op1_09_in14 = reg_0170;
    73: op1_09_in14 = reg_0058;
    110: op1_09_in14 = reg_0058;
    69: op1_09_in14 = imem03_in[7:4];
    74: op1_09_in14 = reg_0167;
    54: op1_09_in14 = reg_0256;
    111: op1_09_in14 = reg_0256;
    68: op1_09_in14 = reg_1065;
    75: op1_09_in14 = reg_0206;
    50: op1_09_in14 = reg_0673;
    71: op1_09_in14 = reg_1406;
    87: op1_09_in14 = reg_0425;
    76: op1_09_in14 = reg_0755;
    61: op1_09_in14 = reg_0389;
    57: op1_09_in14 = reg_0607;
    77: op1_09_in14 = reg_0576;
    58: op1_09_in14 = reg_0779;
    78: op1_09_in14 = reg_0446;
    70: op1_09_in14 = reg_1282;
    79: op1_09_in14 = reg_0353;
    59: op1_09_in14 = reg_0133;
    88: op1_09_in14 = imem04_in[7:4];
    60: op1_09_in14 = reg_0323;
    67: op1_09_in14 = reg_0323;
    46: op1_09_in14 = imem06_in[11:8];
    62: op1_09_in14 = reg_0146;
    80: op1_09_in14 = reg_1302;
    48: op1_09_in14 = reg_0533;
    81: op1_09_in14 = reg_1451;
    52: op1_09_in14 = reg_0888;
    63: op1_09_in14 = reg_1324;
    82: op1_09_in14 = reg_1321;
    89: op1_09_in14 = reg_0478;
    83: op1_09_in14 = reg_0308;
    64: op1_09_in14 = reg_0618;
    84: op1_09_in14 = reg_0463;
    85: op1_09_in14 = reg_0712;
    65: op1_09_in14 = reg_0574;
    90: op1_09_in14 = reg_0668;
    66: op1_09_in14 = reg_0051;
    37: op1_09_in14 = reg_0087;
    91: op1_09_in14 = reg_0440;
    92: op1_09_in14 = reg_0071;
    93: op1_09_in14 = reg_1344;
    94: op1_09_in14 = reg_1090;
    95: op1_09_in14 = reg_0022;
    96: op1_09_in14 = reg_0416;
    106: op1_09_in14 = reg_0416;
    97: op1_09_in14 = reg_0277;
    98: op1_09_in14 = reg_0698;
    99: op1_09_in14 = reg_0397;
    100: op1_09_in14 = reg_0202;
    101: op1_09_in14 = reg_0519;
    102: op1_09_in14 = imem02_in[15:12];
    103: op1_09_in14 = reg_1214;
    44: op1_09_in14 = reg_0799;
    104: op1_09_in14 = reg_1504;
    47: op1_09_in14 = reg_0413;
    105: op1_09_in14 = reg_0792;
    107: op1_09_in14 = reg_0788;
    108: op1_09_in14 = reg_0531;
    109: op1_09_in14 = reg_0208;
    112: op1_09_in14 = reg_0620;
    113: op1_09_in14 = reg_1004;
    114: op1_09_in14 = reg_0276;
    115: op1_09_in14 = reg_0346;
    116: op1_09_in14 = reg_1100;
    117: op1_09_in14 = imem06_in[7:4];
    118: op1_09_in14 = reg_1491;
    40: op1_09_in14 = reg_0016;
    119: op1_09_in14 = reg_0409;
    120: op1_09_in14 = reg_0027;
    121: op1_09_in14 = reg_1091;
    122: op1_09_in14 = imem02_in[11:8];
    123: op1_09_in14 = reg_0117;
    124: op1_09_in14 = reg_0290;
    125: op1_09_in14 = reg_0739;
    126: op1_09_in14 = reg_0162;
    127: op1_09_in14 = reg_0917;
    128: op1_09_in14 = reg_0460;
    42: op1_09_in14 = reg_0631;
    129: op1_09_in14 = reg_1314;
    130: op1_09_in14 = reg_0586;
    131: op1_09_in14 = reg_0829;
    default: op1_09_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv14 = 1;
    53: op1_09_inv14 = 1;
    86: op1_09_inv14 = 1;
    55: op1_09_inv14 = 1;
    73: op1_09_inv14 = 1;
    74: op1_09_inv14 = 1;
    68: op1_09_inv14 = 1;
    78: op1_09_inv14 = 1;
    70: op1_09_inv14 = 1;
    59: op1_09_inv14 = 1;
    88: op1_09_inv14 = 1;
    60: op1_09_inv14 = 1;
    46: op1_09_inv14 = 1;
    52: op1_09_inv14 = 1;
    82: op1_09_inv14 = 1;
    89: op1_09_inv14 = 1;
    83: op1_09_inv14 = 1;
    91: op1_09_inv14 = 1;
    100: op1_09_inv14 = 1;
    102: op1_09_inv14 = 1;
    44: op1_09_inv14 = 1;
    47: op1_09_inv14 = 1;
    105: op1_09_inv14 = 1;
    108: op1_09_inv14 = 1;
    109: op1_09_inv14 = 1;
    111: op1_09_inv14 = 1;
    114: op1_09_inv14 = 1;
    115: op1_09_inv14 = 1;
    118: op1_09_inv14 = 1;
    40: op1_09_inv14 = 1;
    120: op1_09_inv14 = 1;
    122: op1_09_inv14 = 1;
    123: op1_09_inv14 = 1;
    124: op1_09_inv14 = 1;
    125: op1_09_inv14 = 1;
    127: op1_09_inv14 = 1;
    128: op1_09_inv14 = 1;
    42: op1_09_inv14 = 1;
    130: op1_09_inv14 = 1;
    131: op1_09_inv14 = 1;
    default: op1_09_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in15 = reg_0601;
    53: op1_09_in15 = reg_0094;
    103: op1_09_in15 = reg_0094;
    86: op1_09_in15 = reg_0108;
    55: op1_09_in15 = reg_0186;
    73: op1_09_in15 = reg_0267;
    69: op1_09_in15 = imem03_in[11:8];
    74: op1_09_in15 = reg_0090;
    54: op1_09_in15 = reg_0496;
    48: op1_09_in15 = reg_0496;
    68: op1_09_in15 = reg_0676;
    75: op1_09_in15 = reg_0751;
    50: op1_09_in15 = reg_0924;
    71: op1_09_in15 = reg_0883;
    87: op1_09_in15 = reg_0534;
    76: op1_09_in15 = reg_1467;
    61: op1_09_in15 = reg_0351;
    57: op1_09_in15 = reg_0975;
    77: op1_09_in15 = reg_0197;
    58: op1_09_in15 = reg_0442;
    78: op1_09_in15 = reg_0372;
    107: op1_09_in15 = reg_0372;
    70: op1_09_in15 = reg_0790;
    79: op1_09_in15 = reg_0405;
    59: op1_09_in15 = reg_0606;
    42: op1_09_in15 = reg_0606;
    88: op1_09_in15 = imem04_in[11:8];
    60: op1_09_in15 = reg_1202;
    46: op1_09_in15 = reg_0866;
    62: op1_09_in15 = reg_0401;
    80: op1_09_in15 = reg_0194;
    81: op1_09_in15 = reg_1455;
    52: op1_09_in15 = reg_0873;
    63: op1_09_in15 = reg_1322;
    82: op1_09_in15 = reg_1100;
    89: op1_09_in15 = reg_0427;
    83: op1_09_in15 = reg_0270;
    67: op1_09_in15 = reg_0270;
    64: op1_09_in15 = reg_0593;
    84: op1_09_in15 = reg_0258;
    85: op1_09_in15 = reg_1492;
    65: op1_09_in15 = reg_1147;
    90: op1_09_in15 = reg_0786;
    66: op1_09_in15 = reg_0052;
    37: op1_09_in15 = reg_0483;
    91: op1_09_in15 = reg_0416;
    92: op1_09_in15 = reg_0058;
    93: op1_09_in15 = reg_0712;
    102: op1_09_in15 = reg_0712;
    94: op1_09_in15 = reg_1031;
    95: op1_09_in15 = reg_1170;
    96: op1_09_in15 = reg_0410;
    106: op1_09_in15 = reg_0410;
    119: op1_09_in15 = reg_0410;
    97: op1_09_in15 = reg_0785;
    98: op1_09_in15 = reg_1107;
    99: op1_09_in15 = reg_0960;
    100: op1_09_in15 = reg_0353;
    101: op1_09_in15 = reg_0124;
    44: op1_09_in15 = reg_0395;
    104: op1_09_in15 = reg_0172;
    47: op1_09_in15 = reg_0620;
    105: op1_09_in15 = reg_0303;
    108: op1_09_in15 = reg_0574;
    109: op1_09_in15 = reg_1367;
    110: op1_09_in15 = reg_0089;
    111: op1_09_in15 = reg_0096;
    112: op1_09_in15 = reg_0137;
    113: op1_09_in15 = reg_0097;
    114: op1_09_in15 = reg_0608;
    115: op1_09_in15 = reg_0562;
    116: op1_09_in15 = reg_0788;
    117: op1_09_in15 = imem06_in[15:12];
    118: op1_09_in15 = reg_0613;
    40: op1_09_in15 = reg_0020;
    120: op1_09_in15 = reg_0980;
    121: op1_09_in15 = reg_0255;
    122: op1_09_in15 = reg_0659;
    123: op1_09_in15 = reg_0633;
    124: op1_09_in15 = reg_0558;
    125: op1_09_in15 = reg_0740;
    126: op1_09_in15 = reg_0012;
    127: op1_09_in15 = reg_0723;
    128: op1_09_in15 = reg_0155;
    129: op1_09_in15 = reg_1313;
    130: op1_09_in15 = reg_0296;
    131: op1_09_in15 = reg_0745;
    default: op1_09_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv15 = 1;
    86: op1_09_inv15 = 1;
    69: op1_09_inv15 = 1;
    74: op1_09_inv15 = 1;
    54: op1_09_inv15 = 1;
    50: op1_09_inv15 = 1;
    71: op1_09_inv15 = 1;
    87: op1_09_inv15 = 1;
    76: op1_09_inv15 = 1;
    61: op1_09_inv15 = 1;
    58: op1_09_inv15 = 1;
    78: op1_09_inv15 = 1;
    70: op1_09_inv15 = 1;
    60: op1_09_inv15 = 1;
    80: op1_09_inv15 = 1;
    48: op1_09_inv15 = 1;
    81: op1_09_inv15 = 1;
    85: op1_09_inv15 = 1;
    37: op1_09_inv15 = 1;
    67: op1_09_inv15 = 1;
    93: op1_09_inv15 = 1;
    94: op1_09_inv15 = 1;
    95: op1_09_inv15 = 1;
    96: op1_09_inv15 = 1;
    97: op1_09_inv15 = 1;
    99: op1_09_inv15 = 1;
    100: op1_09_inv15 = 1;
    101: op1_09_inv15 = 1;
    104: op1_09_inv15 = 1;
    105: op1_09_inv15 = 1;
    107: op1_09_inv15 = 1;
    108: op1_09_inv15 = 1;
    109: op1_09_inv15 = 1;
    113: op1_09_inv15 = 1;
    116: op1_09_inv15 = 1;
    117: op1_09_inv15 = 1;
    118: op1_09_inv15 = 1;
    40: op1_09_inv15 = 1;
    122: op1_09_inv15 = 1;
    123: op1_09_inv15 = 1;
    124: op1_09_inv15 = 1;
    125: op1_09_inv15 = 1;
    42: op1_09_inv15 = 1;
    129: op1_09_inv15 = 1;
    131: op1_09_inv15 = 1;
    default: op1_09_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in16 = reg_0274;
    53: op1_09_in16 = reg_0096;
    86: op1_09_in16 = reg_0882;
    55: op1_09_in16 = reg_0139;
    73: op1_09_in16 = reg_0788;
    69: op1_09_in16 = reg_0640;
    74: op1_09_in16 = reg_0275;
    54: op1_09_in16 = reg_0971;
    68: op1_09_in16 = reg_0681;
    75: op1_09_in16 = reg_0261;
    50: op1_09_in16 = reg_0489;
    71: op1_09_in16 = reg_0353;
    87: op1_09_in16 = reg_1384;
    76: op1_09_in16 = reg_0268;
    61: op1_09_in16 = reg_0071;
    57: op1_09_in16 = reg_1029;
    77: op1_09_in16 = reg_0393;
    105: op1_09_in16 = reg_0393;
    58: op1_09_in16 = reg_0413;
    78: op1_09_in16 = reg_1256;
    70: op1_09_in16 = reg_0975;
    79: op1_09_in16 = reg_0203;
    59: op1_09_in16 = reg_0256;
    88: op1_09_in16 = reg_0694;
    60: op1_09_in16 = reg_0215;
    46: op1_09_in16 = reg_0720;
    62: op1_09_in16 = reg_0093;
    80: op1_09_in16 = reg_0141;
    48: op1_09_in16 = reg_0473;
    81: op1_09_in16 = reg_1433;
    52: op1_09_in16 = reg_0130;
    63: op1_09_in16 = reg_0448;
    82: op1_09_in16 = reg_1291;
    89: op1_09_in16 = reg_0443;
    83: op1_09_in16 = reg_0498;
    64: op1_09_in16 = reg_0137;
    84: op1_09_in16 = reg_0547;
    85: op1_09_in16 = reg_0800;
    65: op1_09_in16 = reg_0599;
    90: op1_09_in16 = reg_0219;
    66: op1_09_in16 = reg_0519;
    91: op1_09_in16 = reg_0389;
    67: op1_09_in16 = reg_0018;
    92: op1_09_in16 = reg_1322;
    93: op1_09_in16 = reg_0532;
    94: op1_09_in16 = reg_1254;
    95: op1_09_in16 = reg_0509;
    96: op1_09_in16 = reg_0005;
    97: op1_09_in16 = reg_0222;
    98: op1_09_in16 = reg_0064;
    99: op1_09_in16 = reg_0782;
    100: op1_09_in16 = reg_0351;
    102: op1_09_in16 = reg_0436;
    103: op1_09_in16 = reg_0452;
    44: op1_09_in16 = reg_0748;
    104: op1_09_in16 = reg_0780;
    47: op1_09_in16 = reg_0591;
    106: op1_09_in16 = reg_0072;
    107: op1_09_in16 = reg_1032;
    108: op1_09_in16 = reg_0796;
    109: op1_09_in16 = reg_0797;
    110: op1_09_in16 = reg_0980;
    111: op1_09_in16 = reg_1107;
    112: op1_09_in16 = reg_0103;
    113: op1_09_in16 = reg_0033;
    114: op1_09_in16 = reg_0744;
    115: op1_09_in16 = reg_0391;
    116: op1_09_in16 = reg_0930;
    117: op1_09_in16 = reg_0929;
    118: op1_09_in16 = reg_0615;
    40: op1_09_in16 = reg_0032;
    119: op1_09_in16 = reg_0059;
    120: op1_09_in16 = reg_0785;
    121: op1_09_in16 = reg_1515;
    122: op1_09_in16 = reg_0008;
    123: op1_09_in16 = reg_1503;
    124: op1_09_in16 = reg_1093;
    125: op1_09_in16 = reg_0408;
    126: op1_09_in16 = reg_0010;
    127: op1_09_in16 = reg_0677;
    128: op1_09_in16 = reg_0476;
    42: op1_09_in16 = reg_0607;
    129: op1_09_in16 = reg_0962;
    130: op1_09_in16 = reg_0119;
    131: op1_09_in16 = reg_0560;
    default: op1_09_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv16 = 1;
    53: op1_09_inv16 = 1;
    54: op1_09_inv16 = 1;
    75: op1_09_inv16 = 1;
    50: op1_09_inv16 = 1;
    76: op1_09_inv16 = 1;
    61: op1_09_inv16 = 1;
    77: op1_09_inv16 = 1;
    58: op1_09_inv16 = 1;
    79: op1_09_inv16 = 1;
    59: op1_09_inv16 = 1;
    60: op1_09_inv16 = 1;
    46: op1_09_inv16 = 1;
    62: op1_09_inv16 = 1;
    80: op1_09_inv16 = 1;
    48: op1_09_inv16 = 1;
    81: op1_09_inv16 = 1;
    52: op1_09_inv16 = 1;
    82: op1_09_inv16 = 1;
    64: op1_09_inv16 = 1;
    84: op1_09_inv16 = 1;
    85: op1_09_inv16 = 1;
    90: op1_09_inv16 = 1;
    92: op1_09_inv16 = 1;
    94: op1_09_inv16 = 1;
    96: op1_09_inv16 = 1;
    98: op1_09_inv16 = 1;
    99: op1_09_inv16 = 1;
    100: op1_09_inv16 = 1;
    103: op1_09_inv16 = 1;
    104: op1_09_inv16 = 1;
    105: op1_09_inv16 = 1;
    107: op1_09_inv16 = 1;
    108: op1_09_inv16 = 1;
    110: op1_09_inv16 = 1;
    111: op1_09_inv16 = 1;
    113: op1_09_inv16 = 1;
    114: op1_09_inv16 = 1;
    115: op1_09_inv16 = 1;
    116: op1_09_inv16 = 1;
    117: op1_09_inv16 = 1;
    118: op1_09_inv16 = 1;
    120: op1_09_inv16 = 1;
    121: op1_09_inv16 = 1;
    126: op1_09_inv16 = 1;
    127: op1_09_inv16 = 1;
    42: op1_09_inv16 = 1;
    130: op1_09_inv16 = 1;
    default: op1_09_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in17 = reg_0196;
    53: op1_09_in17 = reg_0236;
    86: op1_09_in17 = reg_0481;
    55: op1_09_in17 = reg_0791;
    73: op1_09_in17 = reg_1254;
    82: op1_09_in17 = reg_1254;
    69: op1_09_in17 = reg_1325;
    74: op1_09_in17 = reg_1373;
    54: op1_09_in17 = reg_0935;
    68: op1_09_in17 = reg_0407;
    75: op1_09_in17 = reg_0466;
    50: op1_09_in17 = reg_0665;
    71: op1_09_in17 = reg_0188;
    87: op1_09_in17 = reg_1383;
    76: op1_09_in17 = reg_0192;
    61: op1_09_in17 = reg_0267;
    106: op1_09_in17 = reg_0267;
    57: op1_09_in17 = reg_1140;
    77: op1_09_in17 = reg_0575;
    58: op1_09_in17 = reg_0620;
    78: op1_09_in17 = reg_0166;
    70: op1_09_in17 = reg_0181;
    79: op1_09_in17 = reg_0059;
    59: op1_09_in17 = reg_0889;
    88: op1_09_in17 = reg_1368;
    60: op1_09_in17 = reg_0490;
    95: op1_09_in17 = reg_0490;
    46: op1_09_in17 = reg_0863;
    62: op1_09_in17 = reg_0088;
    80: op1_09_in17 = reg_0585;
    48: op1_09_in17 = reg_0054;
    81: op1_09_in17 = reg_0381;
    52: op1_09_in17 = reg_0205;
    63: op1_09_in17 = reg_0372;
    89: op1_09_in17 = reg_0208;
    83: op1_09_in17 = reg_0867;
    64: op1_09_in17 = reg_0028;
    84: op1_09_in17 = reg_0550;
    85: op1_09_in17 = reg_0312;
    65: op1_09_in17 = reg_0796;
    90: op1_09_in17 = reg_1440;
    66: op1_09_in17 = reg_0521;
    91: op1_09_in17 = reg_0060;
    67: op1_09_in17 = reg_0491;
    92: op1_09_in17 = reg_0122;
    93: op1_09_in17 = reg_0256;
    94: op1_09_in17 = reg_0785;
    96: op1_09_in17 = reg_0723;
    97: op1_09_in17 = reg_0242;
    98: op1_09_in17 = reg_0021;
    123: op1_09_in17 = reg_0021;
    99: op1_09_in17 = reg_0271;
    100: op1_09_in17 = reg_0201;
    102: op1_09_in17 = reg_0326;
    103: op1_09_in17 = reg_0061;
    44: op1_09_in17 = reg_0831;
    104: op1_09_in17 = reg_0115;
    47: op1_09_in17 = reg_0592;
    105: op1_09_in17 = reg_0344;
    107: op1_09_in17 = reg_1253;
    108: op1_09_in17 = reg_0414;
    109: op1_09_in17 = reg_0297;
    110: op1_09_in17 = imem01_in[7:4];
    111: op1_09_in17 = reg_0536;
    112: op1_09_in17 = reg_0051;
    113: op1_09_in17 = reg_0368;
    114: op1_09_in17 = reg_0532;
    115: op1_09_in17 = reg_0564;
    116: op1_09_in17 = reg_0047;
    117: op1_09_in17 = reg_0397;
    118: op1_09_in17 = reg_0616;
    40: op1_09_in17 = reg_0035;
    119: op1_09_in17 = reg_1321;
    120: op1_09_in17 = reg_1152;
    121: op1_09_in17 = reg_0999;
    122: op1_09_in17 = reg_0712;
    124: op1_09_in17 = reg_0107;
    125: op1_09_in17 = reg_0623;
    126: op1_09_in17 = reg_0184;
    127: op1_09_in17 = reg_0982;
    128: op1_09_in17 = reg_1393;
    42: op1_09_in17 = reg_0608;
    129: op1_09_in17 = reg_1231;
    130: op1_09_in17 = reg_1204;
    131: op1_09_in17 = reg_1078;
    default: op1_09_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv17 = 1;
    55: op1_09_inv17 = 1;
    54: op1_09_inv17 = 1;
    68: op1_09_inv17 = 1;
    75: op1_09_inv17 = 1;
    87: op1_09_inv17 = 1;
    61: op1_09_inv17 = 1;
    58: op1_09_inv17 = 1;
    78: op1_09_inv17 = 1;
    70: op1_09_inv17 = 1;
    46: op1_09_inv17 = 1;
    80: op1_09_inv17 = 1;
    48: op1_09_inv17 = 1;
    63: op1_09_inv17 = 1;
    83: op1_09_inv17 = 1;
    64: op1_09_inv17 = 1;
    84: op1_09_inv17 = 1;
    85: op1_09_inv17 = 1;
    65: op1_09_inv17 = 1;
    66: op1_09_inv17 = 1;
    91: op1_09_inv17 = 1;
    67: op1_09_inv17 = 1;
    92: op1_09_inv17 = 1;
    93: op1_09_inv17 = 1;
    95: op1_09_inv17 = 1;
    97: op1_09_inv17 = 1;
    44: op1_09_inv17 = 1;
    104: op1_09_inv17 = 1;
    47: op1_09_inv17 = 1;
    106: op1_09_inv17 = 1;
    109: op1_09_inv17 = 1;
    110: op1_09_inv17 = 1;
    111: op1_09_inv17 = 1;
    114: op1_09_inv17 = 1;
    115: op1_09_inv17 = 1;
    116: op1_09_inv17 = 1;
    118: op1_09_inv17 = 1;
    123: op1_09_inv17 = 1;
    124: op1_09_inv17 = 1;
    125: op1_09_inv17 = 1;
    127: op1_09_inv17 = 1;
    default: op1_09_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in18 = reg_0130;
    53: op1_09_in18 = reg_0237;
    86: op1_09_in18 = reg_0478;
    55: op1_09_in18 = reg_0779;
    73: op1_09_in18 = reg_1069;
    69: op1_09_in18 = reg_0144;
    74: op1_09_in18 = reg_0039;
    54: op1_09_in18 = reg_0848;
    68: op1_09_in18 = reg_0969;
    75: op1_09_in18 = reg_0907;
    50: op1_09_in18 = reg_0663;
    71: op1_09_in18 = reg_0440;
    87: op1_09_in18 = reg_0208;
    76: op1_09_in18 = imem06_in[7:4];
    61: op1_09_in18 = reg_0723;
    57: op1_09_in18 = reg_0973;
    77: op1_09_in18 = reg_0797;
    58: op1_09_in18 = reg_0592;
    78: op1_09_in18 = reg_0463;
    70: op1_09_in18 = reg_0252;
    79: op1_09_in18 = reg_1322;
    119: op1_09_in18 = reg_1322;
    59: op1_09_in18 = reg_0778;
    48: op1_09_in18 = reg_0778;
    88: op1_09_in18 = reg_0034;
    60: op1_09_in18 = reg_1055;
    46: op1_09_in18 = reg_0374;
    62: op1_09_in18 = reg_0291;
    80: op1_09_in18 = reg_0586;
    81: op1_09_in18 = reg_0379;
    52: op1_09_in18 = reg_0206;
    63: op1_09_in18 = imem01_in[7:4];
    82: op1_09_in18 = reg_0747;
    89: op1_09_in18 = reg_0493;
    83: op1_09_in18 = reg_0560;
    64: op1_09_in18 = reg_0228;
    84: op1_09_in18 = reg_0746;
    85: op1_09_in18 = reg_0444;
    65: op1_09_in18 = reg_0342;
    90: op1_09_in18 = reg_0457;
    66: op1_09_in18 = reg_0520;
    91: op1_09_in18 = reg_0072;
    67: op1_09_in18 = reg_1056;
    92: op1_09_in18 = reg_1100;
    93: op1_09_in18 = reg_0436;
    94: op1_09_in18 = reg_1512;
    95: op1_09_in18 = reg_1439;
    96: op1_09_in18 = reg_0871;
    97: op1_09_in18 = reg_0966;
    98: op1_09_in18 = reg_0370;
    99: op1_09_in18 = reg_0115;
    100: op1_09_in18 = reg_0277;
    102: op1_09_in18 = reg_1458;
    103: op1_09_in18 = reg_0698;
    44: op1_09_in18 = reg_0701;
    104: op1_09_in18 = reg_0717;
    47: op1_09_in18 = reg_0102;
    105: op1_09_in18 = reg_0589;
    106: op1_09_in18 = reg_0917;
    107: op1_09_in18 = reg_0401;
    108: op1_09_in18 = reg_0599;
    109: op1_09_in18 = reg_1233;
    110: op1_09_in18 = reg_0635;
    111: op1_09_in18 = reg_1503;
    112: op1_09_in18 = reg_0053;
    113: op1_09_in18 = reg_0904;
    114: op1_09_in18 = reg_0898;
    115: op1_09_in18 = reg_0131;
    116: op1_09_in18 = reg_0553;
    117: op1_09_in18 = reg_0161;
    118: op1_09_in18 = reg_0554;
    40: op1_09_in18 = reg_0792;
    120: op1_09_in18 = reg_0874;
    121: op1_09_in18 = reg_0840;
    122: op1_09_in18 = reg_0839;
    126: op1_09_in18 = reg_0839;
    123: op1_09_in18 = reg_0210;
    124: op1_09_in18 = reg_0880;
    125: op1_09_in18 = reg_0593;
    127: op1_09_in18 = reg_0902;
    128: op1_09_in18 = reg_0887;
    42: op1_09_in18 = reg_0587;
    129: op1_09_in18 = reg_0448;
    130: op1_09_in18 = reg_0754;
    131: op1_09_in18 = reg_0068;
    default: op1_09_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv18 = 1;
    86: op1_09_inv18 = 1;
    55: op1_09_inv18 = 1;
    54: op1_09_inv18 = 1;
    75: op1_09_inv18 = 1;
    87: op1_09_inv18 = 1;
    61: op1_09_inv18 = 1;
    57: op1_09_inv18 = 1;
    77: op1_09_inv18 = 1;
    78: op1_09_inv18 = 1;
    70: op1_09_inv18 = 1;
    59: op1_09_inv18 = 1;
    88: op1_09_inv18 = 1;
    62: op1_09_inv18 = 1;
    80: op1_09_inv18 = 1;
    81: op1_09_inv18 = 1;
    52: op1_09_inv18 = 1;
    82: op1_09_inv18 = 1;
    89: op1_09_inv18 = 1;
    83: op1_09_inv18 = 1;
    64: op1_09_inv18 = 1;
    85: op1_09_inv18 = 1;
    65: op1_09_inv18 = 1;
    90: op1_09_inv18 = 1;
    66: op1_09_inv18 = 1;
    92: op1_09_inv18 = 1;
    96: op1_09_inv18 = 1;
    97: op1_09_inv18 = 1;
    98: op1_09_inv18 = 1;
    99: op1_09_inv18 = 1;
    100: op1_09_inv18 = 1;
    103: op1_09_inv18 = 1;
    44: op1_09_inv18 = 1;
    47: op1_09_inv18 = 1;
    110: op1_09_inv18 = 1;
    112: op1_09_inv18 = 1;
    113: op1_09_inv18 = 1;
    114: op1_09_inv18 = 1;
    115: op1_09_inv18 = 1;
    117: op1_09_inv18 = 1;
    40: op1_09_inv18 = 1;
    119: op1_09_inv18 = 1;
    120: op1_09_inv18 = 1;
    121: op1_09_inv18 = 1;
    122: op1_09_inv18 = 1;
    124: op1_09_inv18 = 1;
    125: op1_09_inv18 = 1;
    129: op1_09_inv18 = 1;
    131: op1_09_inv18 = 1;
    default: op1_09_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in19 = reg_0118;
    53: op1_09_in19 = reg_0117;
    86: op1_09_in19 = imem03_in[15:12];
    55: op1_09_in19 = reg_0665;
    73: op1_09_in19 = reg_0239;
    69: op1_09_in19 = reg_1003;
    74: op1_09_in19 = reg_0751;
    54: op1_09_in19 = reg_0839;
    68: op1_09_in19 = reg_0796;
    75: op1_09_in19 = reg_0172;
    50: op1_09_in19 = reg_0286;
    71: op1_09_in19 = reg_0416;
    87: op1_09_in19 = reg_0263;
    76: op1_09_in19 = reg_0160;
    61: op1_09_in19 = imem00_in[3:0];
    57: op1_09_in19 = reg_0626;
    77: op1_09_in19 = reg_0449;
    58: op1_09_in19 = reg_0114;
    47: op1_09_in19 = reg_0114;
    78: op1_09_in19 = reg_0547;
    70: op1_09_in19 = reg_0462;
    79: op1_09_in19 = reg_0089;
    59: op1_09_in19 = reg_0972;
    48: op1_09_in19 = reg_0972;
    88: op1_09_in19 = reg_0252;
    60: op1_09_in19 = reg_0600;
    46: op1_09_in19 = reg_0827;
    62: op1_09_in19 = reg_0283;
    80: op1_09_in19 = reg_0526;
    81: op1_09_in19 = reg_0531;
    52: op1_09_in19 = reg_0037;
    63: op1_09_in19 = imem01_in[15:12];
    82: op1_09_in19 = reg_0787;
    89: op1_09_in19 = reg_0088;
    83: op1_09_in19 = reg_0162;
    64: op1_09_in19 = reg_0004;
    84: op1_09_in19 = reg_0747;
    85: op1_09_in19 = reg_1448;
    121: op1_09_in19 = reg_1448;
    65: op1_09_in19 = reg_0368;
    103: op1_09_in19 = reg_0368;
    90: op1_09_in19 = reg_0924;
    66: op1_09_in19 = reg_0484;
    91: op1_09_in19 = reg_0723;
    106: op1_09_in19 = reg_0723;
    67: op1_09_in19 = reg_0185;
    92: op1_09_in19 = reg_1152;
    93: op1_09_in19 = reg_0971;
    94: op1_09_in19 = reg_1513;
    95: op1_09_in19 = imem07_in[11:8];
    96: op1_09_in19 = reg_1090;
    100: op1_09_in19 = reg_1090;
    97: op1_09_in19 = reg_0968;
    98: op1_09_in19 = imem05_in[11:8];
    99: op1_09_in19 = reg_0637;
    104: op1_09_in19 = reg_0637;
    102: op1_09_in19 = reg_0382;
    44: op1_09_in19 = reg_0175;
    105: op1_09_in19 = reg_0861;
    107: op1_09_in19 = reg_0743;
    108: op1_09_in19 = reg_1041;
    109: op1_09_in19 = reg_0281;
    110: op1_09_in19 = reg_0047;
    111: op1_09_in19 = reg_0016;
    113: op1_09_in19 = reg_1488;
    114: op1_09_in19 = reg_0533;
    115: op1_09_in19 = reg_1404;
    116: op1_09_in19 = reg_0260;
    117: op1_09_in19 = reg_1209;
    118: op1_09_in19 = reg_0486;
    40: op1_09_in19 = reg_0748;
    119: op1_09_in19 = reg_0005;
    120: op1_09_in19 = reg_0463;
    122: op1_09_in19 = reg_0822;
    123: op1_09_in19 = reg_0347;
    124: op1_09_in19 = reg_0458;
    125: op1_09_in19 = reg_0361;
    126: op1_09_in19 = reg_1493;
    127: op1_09_in19 = reg_0163;
    128: op1_09_in19 = reg_0353;
    42: op1_09_in19 = reg_0562;
    129: op1_09_in19 = reg_0350;
    130: op1_09_in19 = reg_0046;
    131: op1_09_in19 = reg_0217;
    default: op1_09_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv19 = 1;
    69: op1_09_inv19 = 1;
    74: op1_09_inv19 = 1;
    54: op1_09_inv19 = 1;
    75: op1_09_inv19 = 1;
    50: op1_09_inv19 = 1;
    87: op1_09_inv19 = 1;
    76: op1_09_inv19 = 1;
    79: op1_09_inv19 = 1;
    88: op1_09_inv19 = 1;
    60: op1_09_inv19 = 1;
    62: op1_09_inv19 = 1;
    80: op1_09_inv19 = 1;
    82: op1_09_inv19 = 1;
    83: op1_09_inv19 = 1;
    65: op1_09_inv19 = 1;
    91: op1_09_inv19 = 1;
    93: op1_09_inv19 = 1;
    94: op1_09_inv19 = 1;
    95: op1_09_inv19 = 1;
    97: op1_09_inv19 = 1;
    98: op1_09_inv19 = 1;
    99: op1_09_inv19 = 1;
    103: op1_09_inv19 = 1;
    104: op1_09_inv19 = 1;
    47: op1_09_inv19 = 1;
    105: op1_09_inv19 = 1;
    108: op1_09_inv19 = 1;
    115: op1_09_inv19 = 1;
    117: op1_09_inv19 = 1;
    118: op1_09_inv19 = 1;
    119: op1_09_inv19 = 1;
    120: op1_09_inv19 = 1;
    121: op1_09_inv19 = 1;
    122: op1_09_inv19 = 1;
    126: op1_09_inv19 = 1;
    128: op1_09_inv19 = 1;
    42: op1_09_inv19 = 1;
    130: op1_09_inv19 = 1;
    default: op1_09_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in20 = reg_0602;
    53: op1_09_in20 = reg_0129;
    86: op1_09_in20 = reg_0411;
    55: op1_09_in20 = reg_0366;
    73: op1_09_in20 = reg_0238;
    107: op1_09_in20 = reg_0238;
    69: op1_09_in20 = reg_0964;
    74: op1_09_in20 = reg_0261;
    54: op1_09_in20 = reg_0009;
    68: op1_09_in20 = reg_0798;
    75: op1_09_in20 = reg_0669;
    50: op1_09_in20 = reg_0415;
    71: op1_09_in20 = reg_0405;
    87: op1_09_in20 = reg_1372;
    76: op1_09_in20 = reg_0869;
    61: op1_09_in20 = reg_1253;
    57: op1_09_in20 = reg_0933;
    77: op1_09_in20 = reg_0151;
    58: op1_09_in20 = reg_0003;
    78: op1_09_in20 = reg_0747;
    70: op1_09_in20 = reg_0466;
    79: op1_09_in20 = reg_0026;
    59: op1_09_in20 = reg_0127;
    93: op1_09_in20 = reg_0127;
    88: op1_09_in20 = reg_1258;
    60: op1_09_in20 = reg_1183;
    67: op1_09_in20 = reg_1183;
    46: op1_09_in20 = reg_0110;
    62: op1_09_in20 = reg_0013;
    80: op1_09_in20 = reg_0345;
    48: op1_09_in20 = reg_0112;
    81: op1_09_in20 = reg_0294;
    52: op1_09_in20 = reg_0827;
    63: op1_09_in20 = reg_0547;
    82: op1_09_in20 = reg_0609;
    89: op1_09_in20 = reg_1200;
    83: op1_09_in20 = reg_0461;
    64: op1_09_in20 = reg_0001;
    84: op1_09_in20 = reg_0743;
    85: op1_09_in20 = reg_1425;
    65: op1_09_in20 = reg_0835;
    90: op1_09_in20 = reg_0287;
    91: op1_09_in20 = reg_1291;
    92: op1_09_in20 = imem01_in[11:8];
    94: op1_09_in20 = reg_0930;
    95: op1_09_in20 = reg_0667;
    96: op1_09_in20 = reg_1032;
    100: op1_09_in20 = reg_1032;
    97: op1_09_in20 = reg_0819;
    98: op1_09_in20 = reg_0266;
    115: op1_09_in20 = reg_0266;
    99: op1_09_in20 = reg_1228;
    102: op1_09_in20 = reg_0629;
    103: op1_09_in20 = reg_0862;
    44: op1_09_in20 = reg_0565;
    104: op1_09_in20 = reg_0194;
    47: op1_09_in20 = reg_0361;
    105: op1_09_in20 = reg_0207;
    106: op1_09_in20 = reg_1100;
    108: op1_09_in20 = reg_1004;
    109: op1_09_in20 = reg_0599;
    110: op1_09_in20 = reg_0093;
    111: op1_09_in20 = reg_0021;
    113: op1_09_in20 = reg_0370;
    114: op1_09_in20 = reg_0494;
    116: op1_09_in20 = reg_0830;
    117: op1_09_in20 = reg_0730;
    118: op1_09_in20 = reg_0555;
    40: op1_09_in20 = reg_0737;
    119: op1_09_in20 = reg_1512;
    120: op1_09_in20 = reg_0331;
    121: op1_09_in20 = reg_1145;
    122: op1_09_in20 = reg_0390;
    123: op1_09_in20 = reg_1259;
    124: op1_09_in20 = reg_0750;
    125: op1_09_in20 = reg_0052;
    126: op1_09_in20 = reg_0744;
    127: op1_09_in20 = reg_0610;
    128: op1_09_in20 = reg_0351;
    42: op1_09_in20 = reg_0531;
    129: op1_09_in20 = reg_1149;
    130: op1_09_in20 = reg_0152;
    131: op1_09_in20 = reg_0479;
    default: op1_09_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_09_inv20 = 1;
    86: op1_09_inv20 = 1;
    74: op1_09_inv20 = 1;
    68: op1_09_inv20 = 1;
    75: op1_09_inv20 = 1;
    50: op1_09_inv20 = 1;
    71: op1_09_inv20 = 1;
    57: op1_09_inv20 = 1;
    58: op1_09_inv20 = 1;
    78: op1_09_inv20 = 1;
    79: op1_09_inv20 = 1;
    88: op1_09_inv20 = 1;
    62: op1_09_inv20 = 1;
    80: op1_09_inv20 = 1;
    48: op1_09_inv20 = 1;
    81: op1_09_inv20 = 1;
    89: op1_09_inv20 = 1;
    83: op1_09_inv20 = 1;
    84: op1_09_inv20 = 1;
    65: op1_09_inv20 = 1;
    90: op1_09_inv20 = 1;
    91: op1_09_inv20 = 1;
    92: op1_09_inv20 = 1;
    94: op1_09_inv20 = 1;
    95: op1_09_inv20 = 1;
    97: op1_09_inv20 = 1;
    98: op1_09_inv20 = 1;
    103: op1_09_inv20 = 1;
    107: op1_09_inv20 = 1;
    108: op1_09_inv20 = 1;
    110: op1_09_inv20 = 1;
    111: op1_09_inv20 = 1;
    114: op1_09_inv20 = 1;
    115: op1_09_inv20 = 1;
    116: op1_09_inv20 = 1;
    120: op1_09_inv20 = 1;
    124: op1_09_inv20 = 1;
    125: op1_09_inv20 = 1;
    126: op1_09_inv20 = 1;
    127: op1_09_inv20 = 1;
    128: op1_09_inv20 = 1;
    130: op1_09_inv20 = 1;
    default: op1_09_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in21 = imem05_in[3:0];
    111: op1_09_in21 = imem05_in[3:0];
    53: op1_09_in21 = reg_0032;
    86: op1_09_in21 = reg_0247;
    55: op1_09_in21 = reg_0618;
    73: op1_09_in21 = reg_0820;
    69: op1_09_in21 = reg_0962;
    74: op1_09_in21 = reg_0755;
    54: op1_09_in21 = reg_0007;
    81: op1_09_in21 = reg_0007;
    68: op1_09_in21 = reg_0452;
    75: op1_09_in21 = reg_0115;
    50: op1_09_in21 = reg_0137;
    71: op1_09_in21 = reg_0388;
    87: op1_09_in21 = reg_0088;
    76: op1_09_in21 = reg_1504;
    61: op1_09_in21 = reg_1069;
    57: op1_09_in21 = reg_0128;
    77: op1_09_in21 = reg_0195;
    58: op1_09_in21 = reg_0085;
    78: op1_09_in21 = reg_0260;
    70: op1_09_in21 = reg_0414;
    79: op1_09_in21 = reg_1100;
    59: op1_09_in21 = reg_0106;
    88: op1_09_in21 = reg_1200;
    60: op1_09_in21 = reg_0226;
    46: op1_09_in21 = reg_0718;
    52: op1_09_in21 = reg_0718;
    62: op1_09_in21 = reg_0486;
    80: op1_09_in21 = reg_0067;
    48: op1_09_in21 = reg_0900;
    63: op1_09_in21 = reg_0550;
    82: op1_09_in21 = reg_0239;
    89: op1_09_in21 = reg_0281;
    83: op1_09_in21 = reg_0894;
    67: op1_09_in21 = reg_0894;
    95: op1_09_in21 = reg_0894;
    64: op1_09_in21 = reg_0084;
    84: op1_09_in21 = reg_0238;
    85: op1_09_in21 = reg_0177;
    65: op1_09_in21 = reg_0097;
    90: op1_09_in21 = reg_0286;
    91: op1_09_in21 = reg_0930;
    92: op1_09_in21 = reg_1511;
    93: op1_09_in21 = reg_0629;
    94: op1_09_in21 = reg_0047;
    96: op1_09_in21 = reg_0282;
    100: op1_09_in21 = reg_0282;
    97: op1_09_in21 = reg_0439;
    98: op1_09_in21 = reg_0367;
    99: op1_09_in21 = reg_0295;
    102: op1_09_in21 = reg_0897;
    103: op1_09_in21 = reg_0835;
    44: op1_09_in21 = reg_0315;
    104: op1_09_in21 = reg_0374;
    47: op1_09_in21 = reg_0002;
    105: op1_09_in21 = reg_0040;
    106: op1_09_in21 = reg_0277;
    107: op1_09_in21 = reg_0241;
    108: op1_09_in21 = reg_0342;
    109: op1_09_in21 = reg_0454;
    110: op1_09_in21 = reg_0547;
    113: op1_09_in21 = reg_0332;
    114: op1_09_in21 = reg_0054;
    115: op1_09_in21 = reg_0937;
    116: op1_09_in21 = reg_0742;
    117: op1_09_in21 = reg_0696;
    118: op1_09_in21 = reg_0640;
    40: op1_09_in21 = reg_0735;
    119: op1_09_in21 = reg_0269;
    120: op1_09_in21 = reg_0549;
    121: op1_09_in21 = reg_0706;
    122: op1_09_in21 = reg_1207;
    123: op1_09_in21 = reg_0708;
    124: op1_09_in21 = reg_0443;
    125: op1_09_in21 = reg_1182;
    126: op1_09_in21 = reg_0532;
    127: op1_09_in21 = reg_0222;
    128: op1_09_in21 = reg_0201;
    42: op1_09_in21 = reg_0495;
    129: op1_09_in21 = reg_0559;
    130: op1_09_in21 = reg_0215;
    131: op1_09_in21 = reg_0185;
    default: op1_09_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv21 = 1;
    86: op1_09_inv21 = 1;
    73: op1_09_inv21 = 1;
    50: op1_09_inv21 = 1;
    71: op1_09_inv21 = 1;
    87: op1_09_inv21 = 1;
    76: op1_09_inv21 = 1;
    61: op1_09_inv21 = 1;
    59: op1_09_inv21 = 1;
    88: op1_09_inv21 = 1;
    60: op1_09_inv21 = 1;
    62: op1_09_inv21 = 1;
    80: op1_09_inv21 = 1;
    48: op1_09_inv21 = 1;
    81: op1_09_inv21 = 1;
    63: op1_09_inv21 = 1;
    82: op1_09_inv21 = 1;
    89: op1_09_inv21 = 1;
    83: op1_09_inv21 = 1;
    84: op1_09_inv21 = 1;
    85: op1_09_inv21 = 1;
    65: op1_09_inv21 = 1;
    91: op1_09_inv21 = 1;
    98: op1_09_inv21 = 1;
    99: op1_09_inv21 = 1;
    102: op1_09_inv21 = 1;
    44: op1_09_inv21 = 1;
    106: op1_09_inv21 = 1;
    109: op1_09_inv21 = 1;
    111: op1_09_inv21 = 1;
    117: op1_09_inv21 = 1;
    118: op1_09_inv21 = 1;
    119: op1_09_inv21 = 1;
    121: op1_09_inv21 = 1;
    127: op1_09_inv21 = 1;
    42: op1_09_inv21 = 1;
    130: op1_09_inv21 = 1;
    default: op1_09_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in22 = imem05_in[7:4];
    44: op1_09_in22 = imem05_in[7:4];
    53: op1_09_in22 = reg_0034;
    86: op1_09_in22 = reg_0534;
    55: op1_09_in22 = reg_0484;
    73: op1_09_in22 = reg_0742;
    84: op1_09_in22 = reg_0742;
    69: op1_09_in22 = reg_0349;
    74: op1_09_in22 = reg_1435;
    54: op1_09_in22 = reg_0327;
    68: op1_09_in22 = reg_0721;
    75: op1_09_in22 = reg_0716;
    50: op1_09_in22 = reg_0100;
    71: op1_09_in22 = reg_0072;
    87: op1_09_in22 = reg_0264;
    76: op1_09_in22 = reg_0172;
    61: op1_09_in22 = reg_1031;
    57: op1_09_in22 = reg_0112;
    77: op1_09_in22 = reg_1467;
    78: op1_09_in22 = reg_0241;
    70: op1_09_in22 = reg_0412;
    79: op1_09_in22 = reg_0930;
    59: op1_09_in22 = reg_0381;
    88: op1_09_in22 = reg_1215;
    60: op1_09_in22 = reg_0245;
    46: op1_09_in22 = reg_0714;
    52: op1_09_in22 = reg_0714;
    62: op1_09_in22 = reg_0457;
    80: op1_09_in22 = reg_0023;
    48: op1_09_in22 = reg_0712;
    81: op1_09_in22 = reg_0325;
    63: op1_09_in22 = reg_0548;
    120: op1_09_in22 = reg_0548;
    82: op1_09_in22 = reg_1474;
    89: op1_09_in22 = reg_0796;
    83: op1_09_in22 = reg_0310;
    64: op1_09_in22 = reg_0521;
    85: op1_09_in22 = reg_0198;
    65: op1_09_in22 = reg_0237;
    90: op1_09_in22 = reg_0740;
    91: op1_09_in22 = reg_0258;
    67: op1_09_in22 = reg_0139;
    92: op1_09_in22 = reg_0047;
    93: op1_09_in22 = reg_0684;
    94: op1_09_in22 = reg_0093;
    95: op1_09_in22 = reg_0135;
    96: op1_09_in22 = reg_1254;
    97: op1_09_in22 = reg_0290;
    98: op1_09_in22 = reg_0735;
    99: op1_09_in22 = reg_0289;
    100: op1_09_in22 = reg_1253;
    106: op1_09_in22 = reg_1253;
    102: op1_09_in22 = reg_0711;
    103: op1_09_in22 = reg_0904;
    104: op1_09_in22 = reg_0619;
    47: op1_09_in22 = reg_0086;
    105: op1_09_in22 = reg_0270;
    107: op1_09_in22 = reg_0430;
    108: op1_09_in22 = reg_0487;
    109: op1_09_in22 = reg_0835;
    110: op1_09_in22 = reg_0610;
    111: op1_09_in22 = reg_0708;
    113: op1_09_in22 = reg_0184;
    114: op1_09_in22 = reg_0778;
    115: op1_09_in22 = reg_0318;
    116: op1_09_in22 = reg_0469;
    117: op1_09_in22 = reg_0720;
    118: op1_09_in22 = reg_1027;
    40: op1_09_in22 = reg_0345;
    119: op1_09_in22 = reg_0980;
    121: op1_09_in22 = reg_0216;
    122: op1_09_in22 = reg_0494;
    123: op1_09_in22 = reg_0367;
    124: op1_09_in22 = reg_1144;
    126: op1_09_in22 = reg_1074;
    127: op1_09_in22 = reg_0820;
    128: op1_09_in22 = reg_0189;
    42: op1_09_in22 = reg_0456;
    129: op1_09_in22 = reg_0218;
    130: op1_09_in22 = reg_0022;
    131: op1_09_in22 = reg_0311;
    default: op1_09_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv22 = 1;
    53: op1_09_inv22 = 1;
    86: op1_09_inv22 = 1;
    73: op1_09_inv22 = 1;
    74: op1_09_inv22 = 1;
    54: op1_09_inv22 = 1;
    76: op1_09_inv22 = 1;
    61: op1_09_inv22 = 1;
    57: op1_09_inv22 = 1;
    70: op1_09_inv22 = 1;
    79: op1_09_inv22 = 1;
    59: op1_09_inv22 = 1;
    80: op1_09_inv22 = 1;
    48: op1_09_inv22 = 1;
    63: op1_09_inv22 = 1;
    82: op1_09_inv22 = 1;
    83: op1_09_inv22 = 1;
    85: op1_09_inv22 = 1;
    65: op1_09_inv22 = 1;
    67: op1_09_inv22 = 1;
    94: op1_09_inv22 = 1;
    95: op1_09_inv22 = 1;
    96: op1_09_inv22 = 1;
    98: op1_09_inv22 = 1;
    99: op1_09_inv22 = 1;
    102: op1_09_inv22 = 1;
    103: op1_09_inv22 = 1;
    105: op1_09_inv22 = 1;
    106: op1_09_inv22 = 1;
    107: op1_09_inv22 = 1;
    108: op1_09_inv22 = 1;
    109: op1_09_inv22 = 1;
    110: op1_09_inv22 = 1;
    118: op1_09_inv22 = 1;
    122: op1_09_inv22 = 1;
    124: op1_09_inv22 = 1;
    127: op1_09_inv22 = 1;
    42: op1_09_inv22 = 1;
    129: op1_09_inv22 = 1;
    130: op1_09_inv22 = 1;
    131: op1_09_inv22 = 1;
    default: op1_09_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in23 = reg_0449;
    53: op1_09_in23 = reg_0794;
    86: op1_09_in23 = reg_1367;
    73: op1_09_in23 = reg_0612;
    69: op1_09_in23 = reg_1314;
    74: op1_09_in23 = reg_0925;
    105: op1_09_in23 = reg_0925;
    54: op1_09_in23 = reg_0154;
    68: op1_09_in23 = imem04_in[7:4];
    75: op1_09_in23 = reg_0717;
    50: op1_09_in23 = reg_0114;
    71: op1_09_in23 = reg_1322;
    87: op1_09_in23 = reg_0531;
    76: op1_09_in23 = reg_0109;
    61: op1_09_in23 = reg_1034;
    57: op1_09_in23 = reg_0390;
    59: op1_09_in23 = reg_0390;
    77: op1_09_in23 = reg_0316;
    78: op1_09_in23 = reg_0742;
    62: op1_09_in23 = reg_0742;
    127: op1_09_in23 = reg_0742;
    70: op1_09_in23 = reg_0599;
    79: op1_09_in23 = reg_0547;
    94: op1_09_in23 = reg_0547;
    88: op1_09_in23 = reg_0281;
    81: op1_09_in23 = reg_0281;
    60: op1_09_in23 = reg_0704;
    46: op1_09_in23 = reg_0261;
    80: op1_09_in23 = reg_0212;
    48: op1_09_in23 = reg_0708;
    52: op1_09_in23 = reg_0671;
    63: op1_09_in23 = reg_0610;
    82: op1_09_in23 = reg_0385;
    89: op1_09_in23 = reg_1147;
    83: op1_09_in23 = reg_1349;
    64: op1_09_in23 = reg_0520;
    47: op1_09_in23 = reg_0520;
    84: op1_09_in23 = reg_1473;
    85: op1_09_in23 = reg_0847;
    65: op1_09_in23 = reg_0019;
    90: op1_09_in23 = reg_0484;
    91: op1_09_in23 = reg_0550;
    67: op1_09_in23 = reg_0224;
    92: op1_09_in23 = reg_0163;
    93: op1_09_in23 = reg_0876;
    95: op1_09_in23 = reg_0786;
    96: op1_09_in23 = reg_0576;
    97: op1_09_in23 = reg_1513;
    98: op1_09_in23 = reg_0702;
    123: op1_09_in23 = reg_0702;
    99: op1_09_in23 = reg_0371;
    100: op1_09_in23 = reg_0239;
    102: op1_09_in23 = reg_0008;
    103: op1_09_in23 = reg_0016;
    44: op1_09_in23 = imem05_in[11:8];
    40: op1_09_in23 = imem05_in[11:8];
    104: op1_09_in23 = reg_0570;
    106: op1_09_in23 = reg_0874;
    107: op1_09_in23 = reg_1452;
    108: op1_09_in23 = reg_0837;
    109: op1_09_in23 = reg_0096;
    110: op1_09_in23 = reg_0222;
    120: op1_09_in23 = reg_0222;
    111: op1_09_in23 = reg_0347;
    113: op1_09_in23 = reg_0566;
    114: op1_09_in23 = reg_0973;
    115: op1_09_in23 = reg_0736;
    116: op1_09_in23 = reg_0966;
    117: op1_09_in23 = reg_1501;
    118: op1_09_in23 = reg_1454;
    119: op1_09_in23 = reg_0785;
    121: op1_09_in23 = reg_1033;
    122: op1_09_in23 = reg_0970;
    124: op1_09_in23 = reg_0574;
    126: op1_09_in23 = reg_0429;
    128: op1_09_in23 = reg_0060;
    42: op1_09_in23 = reg_0455;
    129: op1_09_in23 = reg_0291;
    130: op1_09_in23 = reg_0156;
    131: op1_09_in23 = reg_0144;
    default: op1_09_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv23 = 1;
    86: op1_09_inv23 = 1;
    73: op1_09_inv23 = 1;
    69: op1_09_inv23 = 1;
    74: op1_09_inv23 = 1;
    54: op1_09_inv23 = 1;
    75: op1_09_inv23 = 1;
    87: op1_09_inv23 = 1;
    57: op1_09_inv23 = 1;
    78: op1_09_inv23 = 1;
    79: op1_09_inv23 = 1;
    59: op1_09_inv23 = 1;
    88: op1_09_inv23 = 1;
    60: op1_09_inv23 = 1;
    46: op1_09_inv23 = 1;
    80: op1_09_inv23 = 1;
    81: op1_09_inv23 = 1;
    52: op1_09_inv23 = 1;
    63: op1_09_inv23 = 1;
    89: op1_09_inv23 = 1;
    64: op1_09_inv23 = 1;
    65: op1_09_inv23 = 1;
    91: op1_09_inv23 = 1;
    93: op1_09_inv23 = 1;
    96: op1_09_inv23 = 1;
    97: op1_09_inv23 = 1;
    98: op1_09_inv23 = 1;
    99: op1_09_inv23 = 1;
    102: op1_09_inv23 = 1;
    104: op1_09_inv23 = 1;
    47: op1_09_inv23 = 1;
    106: op1_09_inv23 = 1;
    108: op1_09_inv23 = 1;
    109: op1_09_inv23 = 1;
    113: op1_09_inv23 = 1;
    114: op1_09_inv23 = 1;
    119: op1_09_inv23 = 1;
    120: op1_09_inv23 = 1;
    122: op1_09_inv23 = 1;
    124: op1_09_inv23 = 1;
    126: op1_09_inv23 = 1;
    127: op1_09_inv23 = 1;
    129: op1_09_inv23 = 1;
    130: op1_09_inv23 = 1;
    131: op1_09_inv23 = 1;
    default: op1_09_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in24 = reg_0038;
    53: op1_09_in24 = reg_0733;
    86: op1_09_in24 = imem04_in[7:4];
    73: op1_09_in24 = reg_0439;
    69: op1_09_in24 = reg_1300;
    74: op1_09_in24 = reg_0860;
    54: op1_09_in24 = reg_0829;
    68: op1_09_in24 = reg_0368;
    75: op1_09_in24 = reg_0374;
    50: op1_09_in24 = reg_0518;
    71: op1_09_in24 = reg_0917;
    87: op1_09_in24 = reg_1203;
    76: op1_09_in24 = reg_1302;
    61: op1_09_in24 = reg_0634;
    57: op1_09_in24 = reg_0306;
    77: op1_09_in24 = reg_1420;
    78: op1_09_in24 = reg_0612;
    127: op1_09_in24 = reg_0612;
    70: op1_09_in24 = reg_0342;
    79: op1_09_in24 = reg_0222;
    59: op1_09_in24 = reg_0708;
    88: op1_09_in24 = reg_0500;
    60: op1_09_in24 = reg_0324;
    46: op1_09_in24 = reg_0619;
    62: op1_09_in24 = reg_0820;
    80: op1_09_in24 = reg_0213;
    48: op1_09_in24 = reg_0153;
    81: op1_09_in24 = reg_0279;
    52: op1_09_in24 = reg_0586;
    63: op1_09_in24 = reg_1152;
    82: op1_09_in24 = reg_0362;
    89: op1_09_in24 = reg_0421;
    83: op1_09_in24 = reg_0157;
    84: op1_09_in24 = reg_1475;
    85: op1_09_in24 = reg_0143;
    65: op1_09_in24 = reg_0020;
    90: op1_09_in24 = reg_0123;
    91: op1_09_in24 = reg_0548;
    67: op1_09_in24 = reg_0775;
    92: op1_09_in24 = reg_0258;
    93: op1_09_in24 = reg_0801;
    94: op1_09_in24 = reg_0787;
    95: op1_09_in24 = reg_0703;
    96: op1_09_in24 = reg_0401;
    97: op1_09_in24 = reg_0595;
    98: op1_09_in24 = reg_0205;
    99: op1_09_in24 = reg_0214;
    100: op1_09_in24 = reg_0241;
    102: op1_09_in24 = reg_1006;
    103: op1_09_in24 = reg_0750;
    44: op1_09_in24 = reg_0418;
    104: op1_09_in24 = reg_0345;
    105: op1_09_in24 = reg_1209;
    106: op1_09_in24 = reg_0902;
    107: op1_09_in24 = reg_1457;
    108: op1_09_in24 = reg_0211;
    109: op1_09_in24 = reg_0904;
    110: op1_09_in24 = reg_0242;
    111: op1_09_in24 = reg_0992;
    113: op1_09_in24 = reg_1181;
    114: op1_09_in24 = reg_0106;
    115: op1_09_in24 = reg_0130;
    116: op1_09_in24 = reg_0434;
    117: op1_09_in24 = reg_0172;
    118: op1_09_in24 = reg_1201;
    40: op1_09_in24 = reg_0702;
    119: op1_09_in24 = reg_0183;
    120: op1_09_in24 = reg_1473;
    121: op1_09_in24 = reg_0198;
    122: op1_09_in24 = reg_0973;
    123: op1_09_in24 = reg_1268;
    124: op1_09_in24 = reg_1200;
    126: op1_09_in24 = reg_0970;
    128: op1_09_in24 = reg_0058;
    42: op1_09_in24 = reg_0054;
    129: op1_09_in24 = reg_1282;
    130: op1_09_in24 = reg_0025;
    131: op1_09_in24 = reg_0180;
    default: op1_09_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv24 = 1;
    53: op1_09_inv24 = 1;
    86: op1_09_inv24 = 1;
    69: op1_09_inv24 = 1;
    75: op1_09_inv24 = 1;
    61: op1_09_inv24 = 1;
    57: op1_09_inv24 = 1;
    77: op1_09_inv24 = 1;
    78: op1_09_inv24 = 1;
    88: op1_09_inv24 = 1;
    60: op1_09_inv24 = 1;
    46: op1_09_inv24 = 1;
    52: op1_09_inv24 = 1;
    89: op1_09_inv24 = 1;
    85: op1_09_inv24 = 1;
    90: op1_09_inv24 = 1;
    91: op1_09_inv24 = 1;
    67: op1_09_inv24 = 1;
    92: op1_09_inv24 = 1;
    93: op1_09_inv24 = 1;
    96: op1_09_inv24 = 1;
    97: op1_09_inv24 = 1;
    98: op1_09_inv24 = 1;
    100: op1_09_inv24 = 1;
    102: op1_09_inv24 = 1;
    44: op1_09_inv24 = 1;
    104: op1_09_inv24 = 1;
    106: op1_09_inv24 = 1;
    107: op1_09_inv24 = 1;
    108: op1_09_inv24 = 1;
    109: op1_09_inv24 = 1;
    110: op1_09_inv24 = 1;
    111: op1_09_inv24 = 1;
    113: op1_09_inv24 = 1;
    114: op1_09_inv24 = 1;
    115: op1_09_inv24 = 1;
    40: op1_09_inv24 = 1;
    119: op1_09_inv24 = 1;
    120: op1_09_inv24 = 1;
    121: op1_09_inv24 = 1;
    122: op1_09_inv24 = 1;
    123: op1_09_inv24 = 1;
    124: op1_09_inv24 = 1;
    126: op1_09_inv24 = 1;
    128: op1_09_inv24 = 1;
    129: op1_09_inv24 = 1;
    130: op1_09_inv24 = 1;
    default: op1_09_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in25 = reg_0751;
    53: op1_09_in25 = reg_0735;
    86: op1_09_in25 = reg_0462;
    73: op1_09_in25 = reg_1452;
    69: op1_09_in25 = reg_0558;
    74: op1_09_in25 = reg_1323;
    54: op1_09_in25 = reg_0069;
    68: op1_09_in25 = reg_0150;
    75: op1_09_in25 = reg_0373;
    71: op1_09_in25 = reg_0786;
    87: op1_09_in25 = reg_1200;
    76: op1_09_in25 = reg_0637;
    61: op1_09_in25 = reg_0601;
    57: op1_09_in25 = reg_0878;
    77: op1_09_in25 = reg_0264;
    78: op1_09_in25 = reg_0715;
    110: op1_09_in25 = reg_0715;
    120: op1_09_in25 = reg_0715;
    70: op1_09_in25 = reg_0487;
    79: op1_09_in25 = reg_0820;
    59: op1_09_in25 = reg_0153;
    88: op1_09_in25 = reg_0406;
    60: op1_09_in25 = reg_0892;
    46: op1_09_in25 = reg_0585;
    62: op1_09_in25 = reg_0632;
    80: op1_09_in25 = reg_0018;
    48: op1_09_in25 = reg_0845;
    81: op1_09_in25 = reg_0999;
    52: op1_09_in25 = reg_0569;
    63: op1_09_in25 = reg_0982;
    82: op1_09_in25 = reg_0365;
    89: op1_09_in25 = reg_0598;
    83: op1_09_in25 = reg_0921;
    84: op1_09_in25 = reg_0572;
    85: op1_09_in25 = reg_0891;
    65: op1_09_in25 = reg_0035;
    109: op1_09_in25 = reg_0035;
    91: op1_09_in25 = reg_0260;
    67: op1_09_in25 = reg_0029;
    92: op1_09_in25 = reg_0547;
    93: op1_09_in25 = reg_0800;
    94: op1_09_in25 = reg_0830;
    95: op1_09_in25 = reg_0157;
    96: op1_09_in25 = reg_0550;
    97: op1_09_in25 = reg_0464;
    98: op1_09_in25 = reg_1268;
    99: op1_09_in25 = reg_0213;
    100: op1_09_in25 = reg_1475;
    102: op1_09_in25 = reg_0235;
    103: op1_09_in25 = reg_0538;
    44: op1_09_in25 = reg_0300;
    104: op1_09_in25 = reg_0979;
    105: op1_09_in25 = reg_0960;
    106: op1_09_in25 = reg_0163;
    107: op1_09_in25 = reg_1456;
    127: op1_09_in25 = reg_1456;
    108: op1_09_in25 = reg_0021;
    111: op1_09_in25 = reg_0392;
    113: op1_09_in25 = reg_1070;
    114: op1_09_in25 = reg_0381;
    115: op1_09_in25 = reg_0344;
    116: op1_09_in25 = reg_0078;
    117: op1_09_in25 = reg_0586;
    118: op1_09_in25 = reg_1206;
    40: op1_09_in25 = reg_0697;
    119: op1_09_in25 = reg_0576;
    121: op1_09_in25 = reg_0180;
    122: op1_09_in25 = reg_0126;
    123: op1_09_in25 = reg_0700;
    124: op1_09_in25 = reg_0412;
    126: op1_09_in25 = reg_0972;
    128: op1_09_in25 = reg_0057;
    42: op1_09_in25 = reg_0390;
    129: op1_09_in25 = reg_0790;
    130: op1_09_in25 = reg_0050;
    131: op1_09_in25 = reg_0789;
    default: op1_09_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv25 = 1;
    53: op1_09_inv25 = 1;
    86: op1_09_inv25 = 1;
    69: op1_09_inv25 = 1;
    75: op1_09_inv25 = 1;
    77: op1_09_inv25 = 1;
    78: op1_09_inv25 = 1;
    79: op1_09_inv25 = 1;
    60: op1_09_inv25 = 1;
    62: op1_09_inv25 = 1;
    48: op1_09_inv25 = 1;
    81: op1_09_inv25 = 1;
    63: op1_09_inv25 = 1;
    82: op1_09_inv25 = 1;
    83: op1_09_inv25 = 1;
    65: op1_09_inv25 = 1;
    67: op1_09_inv25 = 1;
    94: op1_09_inv25 = 1;
    95: op1_09_inv25 = 1;
    97: op1_09_inv25 = 1;
    98: op1_09_inv25 = 1;
    99: op1_09_inv25 = 1;
    100: op1_09_inv25 = 1;
    104: op1_09_inv25 = 1;
    106: op1_09_inv25 = 1;
    107: op1_09_inv25 = 1;
    109: op1_09_inv25 = 1;
    111: op1_09_inv25 = 1;
    114: op1_09_inv25 = 1;
    115: op1_09_inv25 = 1;
    116: op1_09_inv25 = 1;
    117: op1_09_inv25 = 1;
    120: op1_09_inv25 = 1;
    121: op1_09_inv25 = 1;
    122: op1_09_inv25 = 1;
    123: op1_09_inv25 = 1;
    124: op1_09_inv25 = 1;
    128: op1_09_inv25 = 1;
    129: op1_09_inv25 = 1;
    default: op1_09_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in26 = imem06_in[7:4];
    74: op1_09_in26 = imem06_in[7:4];
    53: op1_09_in26 = imem05_in[3:0];
    86: op1_09_in26 = reg_0406;
    73: op1_09_in26 = reg_1456;
    69: op1_09_in26 = reg_1092;
    54: op1_09_in26 = reg_0279;
    68: op1_09_in26 = reg_0064;
    75: op1_09_in26 = reg_0619;
    71: op1_09_in26 = reg_0611;
    87: op1_09_in26 = reg_0488;
    76: op1_09_in26 = reg_0141;
    61: op1_09_in26 = reg_0548;
    92: op1_09_in26 = reg_0548;
    96: op1_09_in26 = reg_0548;
    57: op1_09_in26 = reg_0839;
    77: op1_09_in26 = reg_1334;
    78: op1_09_in26 = reg_0966;
    70: op1_09_in26 = reg_0337;
    79: op1_09_in26 = reg_0572;
    110: op1_09_in26 = reg_0572;
    59: op1_09_in26 = reg_0294;
    88: op1_09_in26 = reg_1041;
    60: op1_09_in26 = imem07_in[15:12];
    46: op1_09_in26 = reg_0526;
    62: op1_09_in26 = reg_1029;
    80: op1_09_in26 = reg_0560;
    48: op1_09_in26 = reg_0024;
    81: op1_09_in26 = reg_0227;
    93: op1_09_in26 = reg_0227;
    52: op1_09_in26 = reg_0460;
    118: op1_09_in26 = reg_0460;
    63: op1_09_in26 = reg_0715;
    82: op1_09_in26 = reg_0363;
    89: op1_09_in26 = reg_0471;
    83: op1_09_in26 = reg_0924;
    84: op1_09_in26 = reg_0147;
    85: op1_09_in26 = reg_1003;
    65: op1_09_in26 = reg_0792;
    91: op1_09_in26 = reg_0609;
    67: op1_09_in26 = reg_0665;
    94: op1_09_in26 = reg_1474;
    95: op1_09_in26 = reg_0223;
    97: op1_09_in26 = reg_0078;
    98: op1_09_in26 = reg_0251;
    99: op1_09_in26 = reg_0394;
    100: op1_09_in26 = reg_0968;
    102: op1_09_in26 = reg_0179;
    103: op1_09_in26 = reg_0136;
    44: op1_09_in26 = reg_0197;
    104: op1_09_in26 = reg_1228;
    105: op1_09_in26 = reg_0316;
    106: op1_09_in26 = reg_0610;
    107: op1_09_in26 = reg_0362;
    108: op1_09_in26 = reg_0020;
    109: op1_09_in26 = reg_0370;
    111: op1_09_in26 = reg_0173;
    113: op1_09_in26 = reg_0938;
    114: op1_09_in26 = reg_0307;
    115: op1_09_in26 = reg_0449;
    116: op1_09_in26 = reg_0724;
    117: op1_09_in26 = reg_0979;
    40: op1_09_in26 = reg_0648;
    119: op1_09_in26 = reg_0902;
    120: op1_09_in26 = reg_0438;
    121: op1_09_in26 = reg_0891;
    122: op1_09_in26 = reg_0106;
    123: op1_09_in26 = reg_1404;
    124: op1_09_in26 = reg_0454;
    126: op1_09_in26 = reg_0125;
    127: op1_09_in26 = reg_1511;
    128: op1_09_in26 = reg_0547;
    42: op1_09_in26 = reg_0105;
    129: op1_09_in26 = reg_0032;
    130: op1_09_in26 = reg_0786;
    131: op1_09_in26 = reg_0142;
    default: op1_09_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv26 = 1;
    86: op1_09_inv26 = 1;
    73: op1_09_inv26 = 1;
    69: op1_09_inv26 = 1;
    54: op1_09_inv26 = 1;
    68: op1_09_inv26 = 1;
    71: op1_09_inv26 = 1;
    87: op1_09_inv26 = 1;
    61: op1_09_inv26 = 1;
    59: op1_09_inv26 = 1;
    88: op1_09_inv26 = 1;
    46: op1_09_inv26 = 1;
    62: op1_09_inv26 = 1;
    80: op1_09_inv26 = 1;
    48: op1_09_inv26 = 1;
    81: op1_09_inv26 = 1;
    52: op1_09_inv26 = 1;
    82: op1_09_inv26 = 1;
    89: op1_09_inv26 = 1;
    67: op1_09_inv26 = 1;
    93: op1_09_inv26 = 1;
    99: op1_09_inv26 = 1;
    100: op1_09_inv26 = 1;
    44: op1_09_inv26 = 1;
    104: op1_09_inv26 = 1;
    105: op1_09_inv26 = 1;
    109: op1_09_inv26 = 1;
    111: op1_09_inv26 = 1;
    114: op1_09_inv26 = 1;
    115: op1_09_inv26 = 1;
    116: op1_09_inv26 = 1;
    40: op1_09_inv26 = 1;
    120: op1_09_inv26 = 1;
    121: op1_09_inv26 = 1;
    122: op1_09_inv26 = 1;
    124: op1_09_inv26 = 1;
    128: op1_09_inv26 = 1;
    42: op1_09_inv26 = 1;
    130: op1_09_inv26 = 1;
    default: op1_09_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in27 = reg_0795;
    53: op1_09_in27 = imem05_in[7:4];
    86: op1_09_in27 = reg_0454;
    73: op1_09_in27 = reg_0400;
    78: op1_09_in27 = reg_0400;
    69: op1_09_in27 = reg_1208;
    74: op1_09_in27 = reg_0984;
    54: op1_09_in27 = reg_0311;
    68: op1_09_in27 = reg_0061;
    75: op1_09_in27 = reg_0528;
    71: op1_09_in27 = reg_0372;
    87: op1_09_in27 = reg_0421;
    76: op1_09_in27 = reg_0584;
    61: op1_09_in27 = reg_0241;
    57: op1_09_in27 = reg_0845;
    77: op1_09_in27 = reg_0160;
    70: op1_09_in27 = reg_0338;
    79: op1_09_in27 = reg_0967;
    63: op1_09_in27 = reg_0967;
    59: op1_09_in27 = reg_0878;
    88: op1_09_in27 = reg_0537;
    60: op1_09_in27 = reg_0673;
    46: op1_09_in27 = reg_0527;
    62: op1_09_in27 = reg_0606;
    80: op1_09_in27 = reg_0162;
    116: op1_09_in27 = reg_0162;
    48: op1_09_in27 = reg_0800;
    81: op1_09_in27 = reg_0198;
    52: op1_09_in27 = reg_0023;
    82: op1_09_in27 = reg_0899;
    89: op1_09_in27 = reg_0451;
    124: op1_09_in27 = reg_0451;
    83: op1_09_in27 = reg_0139;
    84: op1_09_in27 = reg_0362;
    85: op1_09_in27 = reg_0965;
    65: op1_09_in27 = reg_0737;
    91: op1_09_in27 = reg_0239;
    67: op1_09_in27 = reg_0285;
    92: op1_09_in27 = reg_0746;
    96: op1_09_in27 = reg_0746;
    93: op1_09_in27 = reg_0559;
    94: op1_09_in27 = reg_0572;
    95: op1_09_in27 = reg_0030;
    97: op1_09_in27 = reg_0077;
    98: op1_09_in27 = reg_0831;
    99: op1_09_in27 = reg_1010;
    100: op1_09_in27 = reg_0439;
    102: op1_09_in27 = reg_1448;
    103: op1_09_in27 = reg_0347;
    44: op1_09_in27 = reg_0864;
    104: op1_09_in27 = reg_0296;
    105: op1_09_in27 = reg_0974;
    106: op1_09_in27 = reg_0798;
    107: op1_09_in27 = reg_0092;
    108: op1_09_in27 = reg_0210;
    109: op1_09_in27 = reg_0890;
    110: op1_09_in27 = reg_0147;
    120: op1_09_in27 = reg_0147;
    111: op1_09_in27 = reg_0491;
    113: op1_09_in27 = reg_1514;
    114: op1_09_in27 = reg_0829;
    115: op1_09_in27 = reg_0461;
    117: op1_09_in27 = reg_0522;
    118: op1_09_in27 = reg_0524;
    40: op1_09_in27 = reg_0650;
    119: op1_09_in27 = reg_0401;
    121: op1_09_in27 = reg_0789;
    122: op1_09_in27 = reg_0629;
    123: op1_09_in27 = reg_0302;
    126: op1_09_in27 = reg_0111;
    127: op1_09_in27 = reg_0091;
    128: op1_09_in27 = reg_0120;
    42: op1_09_in27 = reg_0342;
    129: op1_09_in27 = reg_0236;
    130: op1_09_in27 = reg_0225;
    131: op1_09_in27 = reg_0962;
    default: op1_09_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_09_inv27 = 1;
    73: op1_09_inv27 = 1;
    75: op1_09_inv27 = 1;
    87: op1_09_inv27 = 1;
    76: op1_09_inv27 = 1;
    79: op1_09_inv27 = 1;
    60: op1_09_inv27 = 1;
    46: op1_09_inv27 = 1;
    62: op1_09_inv27 = 1;
    80: op1_09_inv27 = 1;
    48: op1_09_inv27 = 1;
    52: op1_09_inv27 = 1;
    89: op1_09_inv27 = 1;
    83: op1_09_inv27 = 1;
    85: op1_09_inv27 = 1;
    65: op1_09_inv27 = 1;
    91: op1_09_inv27 = 1;
    67: op1_09_inv27 = 1;
    94: op1_09_inv27 = 1;
    95: op1_09_inv27 = 1;
    98: op1_09_inv27 = 1;
    99: op1_09_inv27 = 1;
    100: op1_09_inv27 = 1;
    102: op1_09_inv27 = 1;
    103: op1_09_inv27 = 1;
    107: op1_09_inv27 = 1;
    110: op1_09_inv27 = 1;
    113: op1_09_inv27 = 1;
    115: op1_09_inv27 = 1;
    40: op1_09_inv27 = 1;
    119: op1_09_inv27 = 1;
    120: op1_09_inv27 = 1;
    121: op1_09_inv27 = 1;
    122: op1_09_inv27 = 1;
    124: op1_09_inv27 = 1;
    129: op1_09_inv27 = 1;
    default: op1_09_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in28 = reg_1436;
    53: op1_09_in28 = reg_0646;
    86: op1_09_in28 = reg_0342;
    73: op1_09_in28 = reg_0362;
    69: op1_09_in28 = reg_0108;
    74: op1_09_in28 = reg_0718;
    54: op1_09_in28 = reg_0757;
    68: op1_09_in28 = reg_0021;
    75: op1_09_in28 = reg_0570;
    71: op1_09_in28 = reg_1253;
    87: op1_09_in28 = reg_0414;
    76: op1_09_in28 = reg_0571;
    61: op1_09_in28 = reg_0984;
    57: op1_09_in28 = reg_0006;
    77: op1_09_in28 = reg_0161;
    78: op1_09_in28 = reg_0077;
    70: op1_09_in28 = reg_0336;
    79: op1_09_in28 = reg_0438;
    59: op1_09_in28 = reg_0877;
    88: op1_09_in28 = reg_1040;
    60: op1_09_in28 = reg_0921;
    46: op1_09_in28 = reg_0522;
    62: op1_09_in28 = reg_0608;
    80: op1_09_in28 = reg_0922;
    48: op1_09_in28 = reg_0198;
    81: op1_09_in28 = reg_0378;
    52: op1_09_in28 = reg_0152;
    63: op1_09_in28 = reg_0146;
    110: op1_09_in28 = reg_0146;
    82: op1_09_in28 = reg_0901;
    89: op1_09_in28 = reg_0452;
    83: op1_09_in28 = reg_0779;
    84: op1_09_in28 = reg_0091;
    120: op1_09_in28 = reg_0091;
    85: op1_09_in28 = reg_0964;
    65: op1_09_in28 = reg_0833;
    91: op1_09_in28 = reg_0241;
    67: op1_09_in28 = reg_0103;
    92: op1_09_in28 = reg_0260;
    93: op1_09_in28 = reg_0709;
    94: op1_09_in28 = reg_0966;
    95: op1_09_in28 = reg_0441;
    96: op1_09_in28 = reg_0787;
    97: op1_09_in28 = reg_0011;
    98: op1_09_in28 = reg_0562;
    99: op1_09_in28 = reg_1060;
    100: op1_09_in28 = reg_1452;
    102: op1_09_in28 = reg_1425;
    103: op1_09_in28 = reg_0066;
    44: op1_09_in28 = reg_0204;
    104: op1_09_in28 = reg_0171;
    105: op1_09_in28 = reg_0115;
    106: op1_09_in28 = reg_0469;
    107: op1_09_in28 = reg_0078;
    108: op1_09_in28 = reg_0035;
    109: op1_09_in28 = reg_1298;
    111: op1_09_in28 = reg_1104;
    113: op1_09_in28 = reg_0302;
    114: op1_09_in28 = reg_0802;
    115: op1_09_in28 = reg_0270;
    116: op1_09_in28 = reg_0010;
    117: op1_09_in28 = reg_0132;
    118: op1_09_in28 = reg_1405;
    40: op1_09_in28 = reg_0601;
    119: op1_09_in28 = reg_0930;
    121: op1_09_in28 = imem03_in[3:0];
    122: op1_09_in28 = reg_1433;
    123: op1_09_in28 = reg_0492;
    124: op1_09_in28 = reg_0320;
    126: op1_09_in28 = reg_0106;
    127: op1_09_in28 = reg_0080;
    128: op1_09_in28 = imem01_in[7:4];
    42: op1_09_in28 = reg_0705;
    129: op1_09_in28 = reg_0337;
    130: op1_09_in28 = reg_0159;
    131: op1_09_in28 = reg_0376;
    default: op1_09_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv28 = 1;
    73: op1_09_inv28 = 1;
    74: op1_09_inv28 = 1;
    54: op1_09_inv28 = 1;
    68: op1_09_inv28 = 1;
    75: op1_09_inv28 = 1;
    71: op1_09_inv28 = 1;
    87: op1_09_inv28 = 1;
    78: op1_09_inv28 = 1;
    70: op1_09_inv28 = 1;
    59: op1_09_inv28 = 1;
    88: op1_09_inv28 = 1;
    46: op1_09_inv28 = 1;
    62: op1_09_inv28 = 1;
    80: op1_09_inv28 = 1;
    82: op1_09_inv28 = 1;
    89: op1_09_inv28 = 1;
    83: op1_09_inv28 = 1;
    84: op1_09_inv28 = 1;
    85: op1_09_inv28 = 1;
    65: op1_09_inv28 = 1;
    67: op1_09_inv28 = 1;
    93: op1_09_inv28 = 1;
    95: op1_09_inv28 = 1;
    96: op1_09_inv28 = 1;
    98: op1_09_inv28 = 1;
    99: op1_09_inv28 = 1;
    100: op1_09_inv28 = 1;
    102: op1_09_inv28 = 1;
    103: op1_09_inv28 = 1;
    105: op1_09_inv28 = 1;
    107: op1_09_inv28 = 1;
    108: op1_09_inv28 = 1;
    111: op1_09_inv28 = 1;
    115: op1_09_inv28 = 1;
    40: op1_09_inv28 = 1;
    120: op1_09_inv28 = 1;
    122: op1_09_inv28 = 1;
    124: op1_09_inv28 = 1;
    126: op1_09_inv28 = 1;
    42: op1_09_inv28 = 1;
    default: op1_09_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in29 = reg_1426;
    53: op1_09_in29 = reg_0996;
    86: op1_09_in29 = reg_0698;
    73: op1_09_in29 = reg_0727;
    69: op1_09_in29 = reg_0107;
    74: op1_09_in29 = reg_0617;
    54: op1_09_in29 = reg_0756;
    68: op1_09_in29 = reg_0033;
    75: op1_09_in29 = reg_1228;
    71: op1_09_in29 = reg_1254;
    87: op1_09_in29 = reg_1040;
    76: op1_09_in29 = reg_0979;
    61: op1_09_in29 = reg_0743;
    57: op1_09_in29 = reg_0154;
    77: op1_09_in29 = reg_0115;
    78: op1_09_in29 = reg_0291;
    70: op1_09_in29 = reg_0096;
    79: op1_09_in29 = reg_1456;
    59: op1_09_in29 = reg_0008;
    88: op1_09_in29 = reg_0199;
    60: op1_09_in29 = reg_0489;
    46: op1_09_in29 = reg_0295;
    62: op1_09_in29 = reg_0561;
    80: op1_09_in29 = reg_0309;
    48: op1_09_in29 = reg_0707;
    81: op1_09_in29 = reg_0541;
    52: op1_09_in29 = reg_0457;
    63: op1_09_in29 = reg_0400;
    82: op1_09_in29 = reg_0257;
    89: op1_09_in29 = reg_0342;
    83: op1_09_in29 = reg_0740;
    84: op1_09_in29 = reg_0901;
    85: op1_09_in29 = reg_0314;
    65: op1_09_in29 = reg_1168;
    91: op1_09_in29 = reg_0830;
    92: op1_09_in29 = reg_0830;
    67: op1_09_in29 = reg_0100;
    93: op1_09_in29 = reg_1449;
    94: op1_09_in29 = reg_0149;
    95: op1_09_in29 = reg_0593;
    96: op1_09_in29 = reg_0222;
    97: op1_09_in29 = reg_1068;
    98: op1_09_in29 = reg_0173;
    99: op1_09_in29 = reg_0892;
    100: op1_09_in29 = reg_0726;
    102: op1_09_in29 = reg_0177;
    103: op1_09_in29 = reg_0167;
    44: op1_09_in29 = reg_0207;
    104: op1_09_in29 = reg_0244;
    105: op1_09_in29 = reg_0109;
    106: op1_09_in29 = reg_0147;
    107: op1_09_in29 = reg_0042;
    108: op1_09_in29 = imem05_in[3:0];
    109: op1_09_in29 = reg_1485;
    110: op1_09_in29 = reg_0290;
    111: op1_09_in29 = reg_0697;
    113: op1_09_in29 = reg_0090;
    114: op1_09_in29 = reg_0800;
    115: op1_09_in29 = imem06_in[7:4];
    116: op1_09_in29 = reg_0845;
    117: op1_09_in29 = reg_1202;
    118: op1_09_in29 = reg_0887;
    40: op1_09_in29 = reg_0602;
    119: op1_09_in29 = reg_0548;
    120: op1_09_in29 = reg_0899;
    121: op1_09_in29 = reg_0458;
    122: op1_09_in29 = reg_1140;
    123: op1_09_in29 = reg_1346;
    124: op1_09_in29 = reg_1340;
    126: op1_09_in29 = reg_0105;
    127: op1_09_in29 = reg_0896;
    128: op1_09_in29 = reg_0183;
    42: op1_09_in29 = reg_0848;
    129: op1_09_in29 = reg_1258;
    130: op1_09_in29 = reg_0139;
    131: op1_09_in29 = reg_1231;
    default: op1_09_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv29 = 1;
    86: op1_09_inv29 = 1;
    73: op1_09_inv29 = 1;
    69: op1_09_inv29 = 1;
    68: op1_09_inv29 = 1;
    75: op1_09_inv29 = 1;
    76: op1_09_inv29 = 1;
    77: op1_09_inv29 = 1;
    78: op1_09_inv29 = 1;
    79: op1_09_inv29 = 1;
    59: op1_09_inv29 = 1;
    88: op1_09_inv29 = 1;
    60: op1_09_inv29 = 1;
    46: op1_09_inv29 = 1;
    81: op1_09_inv29 = 1;
    63: op1_09_inv29 = 1;
    82: op1_09_inv29 = 1;
    89: op1_09_inv29 = 1;
    84: op1_09_inv29 = 1;
    65: op1_09_inv29 = 1;
    67: op1_09_inv29 = 1;
    92: op1_09_inv29 = 1;
    93: op1_09_inv29 = 1;
    94: op1_09_inv29 = 1;
    96: op1_09_inv29 = 1;
    105: op1_09_inv29 = 1;
    108: op1_09_inv29 = 1;
    109: op1_09_inv29 = 1;
    111: op1_09_inv29 = 1;
    115: op1_09_inv29 = 1;
    116: op1_09_inv29 = 1;
    117: op1_09_inv29 = 1;
    118: op1_09_inv29 = 1;
    40: op1_09_inv29 = 1;
    120: op1_09_inv29 = 1;
    122: op1_09_inv29 = 1;
    123: op1_09_inv29 = 1;
    124: op1_09_inv29 = 1;
    126: op1_09_inv29 = 1;
    128: op1_09_inv29 = 1;
    129: op1_09_inv29 = 1;
    default: op1_09_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_09_in30 = reg_0907;
    53: op1_09_in30 = reg_0997;
    86: op1_09_in30 = reg_0319;
    73: op1_09_in30 = reg_0078;
    84: op1_09_in30 = reg_0078;
    69: op1_09_in30 = reg_0504;
    74: op1_09_in30 = reg_0624;
    54: op1_09_in30 = reg_0525;
    68: op1_09_in30 = reg_0035;
    75: op1_09_in30 = reg_0171;
    46: op1_09_in30 = reg_0171;
    71: op1_09_in30 = reg_1032;
    87: op1_09_in30 = reg_0199;
    76: op1_09_in30 = reg_0522;
    61: op1_09_in30 = reg_0982;
    57: op1_09_in30 = reg_0069;
    77: op1_09_in30 = reg_0716;
    78: op1_09_in30 = reg_0278;
    70: op1_09_in30 = reg_0209;
    79: op1_09_in30 = reg_0400;
    59: op1_09_in30 = reg_0830;
    88: op1_09_in30 = reg_1077;
    60: op1_09_in30 = reg_0777;
    62: op1_09_in30 = reg_0497;
    80: op1_09_in30 = reg_0159;
    48: op1_09_in30 = reg_0706;
    81: op1_09_in30 = reg_0962;
    52: op1_09_in30 = reg_1057;
    63: op1_09_in30 = reg_0093;
    82: op1_09_in30 = reg_0595;
    89: op1_09_in30 = reg_0369;
    83: op1_09_in30 = reg_0408;
    85: op1_09_in30 = reg_0957;
    65: op1_09_in30 = reg_0174;
    91: op1_09_in30 = reg_0798;
    92: op1_09_in30 = reg_0798;
    67: op1_09_in30 = reg_0003;
    93: op1_09_in30 = reg_1033;
    94: op1_09_in30 = reg_0148;
    95: op1_09_in30 = reg_0592;
    96: op1_09_in30 = reg_0241;
    97: op1_09_in30 = reg_0662;
    98: op1_09_in30 = reg_0391;
    99: op1_09_in30 = reg_0786;
    100: op1_09_in30 = reg_1511;
    102: op1_09_in30 = reg_0600;
    103: op1_09_in30 = reg_1401;
    44: op1_09_in30 = reg_0040;
    104: op1_09_in30 = reg_0165;
    105: op1_09_in30 = reg_1303;
    106: op1_09_in30 = reg_0175;
    107: op1_09_in30 = reg_0533;
    108: op1_09_in30 = reg_0702;
    109: op1_09_in30 = reg_1259;
    110: op1_09_in30 = reg_0335;
    111: op1_09_in30 = reg_1404;
    113: op1_09_in30 = reg_0872;
    114: op1_09_in30 = reg_1006;
    115: op1_09_in30 = reg_0161;
    116: op1_09_in30 = reg_0879;
    117: op1_09_in30 = reg_0195;
    118: op1_09_in30 = reg_0352;
    40: op1_09_in30 = reg_0603;
    119: op1_09_in30 = reg_0222;
    120: op1_09_in30 = reg_0464;
    121: op1_09_in30 = reg_0313;
    122: op1_09_in30 = reg_0628;
    123: op1_09_in30 = reg_0864;
    124: op1_09_in30 = reg_1502;
    126: op1_09_in30 = reg_0496;
    127: op1_09_in30 = reg_0042;
    128: op1_09_in30 = reg_0746;
    42: op1_09_in30 = reg_0845;
    129: op1_09_in30 = reg_0978;
    130: op1_09_in30 = reg_0665;
    131: op1_09_in30 = reg_1092;
    default: op1_09_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_09_inv30 = 1;
    53: op1_09_inv30 = 1;
    86: op1_09_inv30 = 1;
    69: op1_09_inv30 = 1;
    54: op1_09_inv30 = 1;
    71: op1_09_inv30 = 1;
    76: op1_09_inv30 = 1;
    61: op1_09_inv30 = 1;
    77: op1_09_inv30 = 1;
    79: op1_09_inv30 = 1;
    62: op1_09_inv30 = 1;
    80: op1_09_inv30 = 1;
    48: op1_09_inv30 = 1;
    81: op1_09_inv30 = 1;
    52: op1_09_inv30 = 1;
    63: op1_09_inv30 = 1;
    82: op1_09_inv30 = 1;
    83: op1_09_inv30 = 1;
    85: op1_09_inv30 = 1;
    65: op1_09_inv30 = 1;
    91: op1_09_inv30 = 1;
    67: op1_09_inv30 = 1;
    92: op1_09_inv30 = 1;
    93: op1_09_inv30 = 1;
    96: op1_09_inv30 = 1;
    98: op1_09_inv30 = 1;
    100: op1_09_inv30 = 1;
    104: op1_09_inv30 = 1;
    105: op1_09_inv30 = 1;
    106: op1_09_inv30 = 1;
    108: op1_09_inv30 = 1;
    110: op1_09_inv30 = 1;
    113: op1_09_inv30 = 1;
    117: op1_09_inv30 = 1;
    40: op1_09_inv30 = 1;
    119: op1_09_inv30 = 1;
    122: op1_09_inv30 = 1;
    124: op1_09_inv30 = 1;
    42: op1_09_inv30 = 1;
    130: op1_09_inv30 = 1;
    default: op1_09_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_09_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#9の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_09_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in00 = reg_0368;
    53: op1_10_in00 = reg_0798;
    86: op1_10_in00 = reg_1098;
    55: op1_10_in00 = reg_0464;
    73: op1_10_in00 = reg_0750;
    69: op1_10_in00 = reg_0557;
    49: op1_10_in00 = reg_0583;
    74: op1_10_in00 = reg_0906;
    54: op1_10_in00 = reg_0020;
    68: op1_10_in00 = reg_0964;
    75: op1_10_in00 = reg_0554;
    77: op1_10_in00 = reg_0554;
    67: op1_10_in00 = reg_0554;
    50: op1_10_in00 = reg_0786;
    56: op1_10_in00 = reg_0305;
    71: op1_10_in00 = reg_0866;
    61: op1_10_in00 = reg_0866;
    87: op1_10_in00 = reg_0032;
    76: op1_10_in00 = reg_0346;
    57: op1_10_in00 = reg_0195;
    58: op1_10_in00 = reg_0434;
    78: op1_10_in00 = reg_1346;
    70: op1_10_in00 = reg_0261;
    89: op1_10_in00 = reg_0261;
    79: op1_10_in00 = reg_0579;
    51: op1_10_in00 = reg_0308;
    59: op1_10_in00 = reg_0598;
    60: op1_10_in00 = reg_0277;
    88: op1_10_in00 = reg_1226;
    46: op1_10_in00 = reg_0574;
    129: op1_10_in00 = reg_0574;
    80: op1_10_in00 = imem00_in[7:4];
    62: op1_10_in00 = reg_1182;
    81: op1_10_in00 = reg_1151;
    52: op1_10_in00 = reg_0998;
    63: op1_10_in00 = reg_0023;
    82: op1_10_in00 = reg_0133;
    33: op1_10_in00 = imem07_in[11:8];
    37: op1_10_in00 = imem07_in[11:8];
    83: op1_10_in00 = reg_0907;
    64: op1_10_in00 = imem02_in[11:8];
    84: op1_10_in00 = reg_0088;
    48: op1_10_in00 = reg_0754;
    85: op1_10_in00 = reg_0566;
    65: op1_10_in00 = reg_0270;
    90: op1_10_in00 = reg_0983;
    101: op1_10_in00 = reg_0983;
    66: op1_10_in00 = reg_1256;
    91: op1_10_in00 = reg_1448;
    28: op1_10_in00 = reg_0003;
    92: op1_10_in00 = reg_0350;
    93: op1_10_in00 = imem03_in[3:0];
    94: op1_10_in00 = reg_0383;
    95: op1_10_in00 = reg_0319;
    96: op1_10_in00 = reg_0631;
    97: op1_10_in00 = reg_0666;
    98: op1_10_in00 = reg_0491;
    99: op1_10_in00 = reg_1440;
    100: op1_10_in00 = reg_0365;
    102: op1_10_in00 = reg_0145;
    103: op1_10_in00 = reg_0940;
    104: op1_10_in00 = reg_1202;
    47: op1_10_in00 = reg_0445;
    105: op1_10_in00 = reg_0398;
    106: op1_10_in00 = reg_0080;
    44: op1_10_in00 = reg_0745;
    107: op1_10_in00 = reg_0626;
    108: op1_10_in00 = reg_0395;
    109: op1_10_in00 = reg_0315;
    110: op1_10_in00 = reg_0162;
    111: op1_10_in00 = reg_0792;
    112: op1_10_in00 = reg_1277;
    113: op1_10_in00 = reg_0450;
    114: op1_10_in00 = reg_0068;
    115: op1_10_in00 = reg_1334;
    116: op1_10_in00 = reg_0138;
    117: op1_10_in00 = reg_0067;
    118: op1_10_in00 = reg_0189;
    119: op1_10_in00 = reg_1207;
    120: op1_10_in00 = reg_0043;
    121: op1_10_in00 = reg_0208;
    122: op1_10_in00 = reg_0306;
    123: op1_10_in00 = reg_0207;
    34: op1_10_in00 = reg_0404;
    124: op1_10_in00 = reg_0019;
    125: op1_10_in00 = reg_0843;
    126: op1_10_in00 = reg_1433;
    127: op1_10_in00 = reg_0447;
    38: op1_10_in00 = reg_0284;
    128: op1_10_in00 = reg_0253;
    130: op1_10_in00 = reg_1489;
    42: op1_10_in00 = reg_0550;
    131: op1_10_in00 = reg_0113;
    default: op1_10_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv00 = 1;
    74: op1_10_inv00 = 1;
    56: op1_10_inv00 = 1;
    87: op1_10_inv00 = 1;
    59: op1_10_inv00 = 1;
    88: op1_10_inv00 = 1;
    46: op1_10_inv00 = 1;
    52: op1_10_inv00 = 1;
    63: op1_10_inv00 = 1;
    89: op1_10_inv00 = 1;
    33: op1_10_inv00 = 1;
    83: op1_10_inv00 = 1;
    64: op1_10_inv00 = 1;
    84: op1_10_inv00 = 1;
    85: op1_10_inv00 = 1;
    91: op1_10_inv00 = 1;
    28: op1_10_inv00 = 1;
    98: op1_10_inv00 = 1;
    100: op1_10_inv00 = 1;
    101: op1_10_inv00 = 1;
    105: op1_10_inv00 = 1;
    44: op1_10_inv00 = 1;
    107: op1_10_inv00 = 1;
    109: op1_10_inv00 = 1;
    110: op1_10_inv00 = 1;
    113: op1_10_inv00 = 1;
    114: op1_10_inv00 = 1;
    118: op1_10_inv00 = 1;
    121: op1_10_inv00 = 1;
    123: op1_10_inv00 = 1;
    38: op1_10_inv00 = 1;
    131: op1_10_inv00 = 1;
    default: op1_10_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in01 = reg_0835;
    53: op1_10_in01 = reg_0795;
    86: op1_10_in01 = reg_0695;
    55: op1_10_in01 = reg_0978;
    73: op1_10_in01 = reg_0833;
    69: op1_10_in01 = reg_0177;
    49: op1_10_in01 = reg_0568;
    74: op1_10_in01 = reg_0863;
    54: op1_10_in01 = reg_0579;
    68: op1_10_in01 = reg_0627;
    75: op1_10_in01 = reg_0616;
    50: op1_10_in01 = reg_0601;
    56: op1_10_in01 = reg_0338;
    71: op1_10_in01 = reg_1244;
    87: op1_10_in01 = reg_1368;
    76: op1_10_in01 = reg_0646;
    61: op1_10_in01 = reg_0841;
    57: op1_10_in01 = reg_0141;
    77: op1_10_in01 = reg_0748;
    44: op1_10_in01 = reg_0748;
    58: op1_10_in01 = reg_0383;
    78: op1_10_in01 = reg_0589;
    70: op1_10_in01 = reg_1000;
    79: op1_10_in01 = reg_1430;
    51: op1_10_in01 = reg_0212;
    59: op1_10_in01 = reg_0969;
    60: op1_10_in01 = reg_0283;
    88: op1_10_in01 = reg_0025;
    46: op1_10_in01 = reg_0582;
    80: op1_10_in01 = reg_0552;
    81: op1_10_in01 = reg_0063;
    52: op1_10_in01 = reg_0298;
    63: op1_10_in01 = reg_0214;
    82: op1_10_in01 = reg_0869;
    89: op1_10_in01 = reg_0143;
    33: op1_10_in01 = reg_0591;
    83: op1_10_in01 = reg_1079;
    64: op1_10_in01 = reg_0184;
    84: op1_10_in01 = reg_0291;
    48: op1_10_in01 = reg_0195;
    104: op1_10_in01 = reg_0195;
    85: op1_10_in01 = reg_0334;
    65: op1_10_in01 = reg_0995;
    90: op1_10_in01 = reg_1243;
    66: op1_10_in01 = reg_1069;
    37: op1_10_in01 = reg_0623;
    91: op1_10_in01 = reg_1063;
    28: op1_10_in01 = reg_0086;
    67: op1_10_in01 = reg_0613;
    92: op1_10_in01 = reg_0541;
    93: op1_10_in01 = reg_0965;
    94: op1_10_in01 = reg_0595;
    95: op1_10_in01 = reg_0501;
    96: op1_10_in01 = reg_0802;
    97: op1_10_in01 = reg_0474;
    98: op1_10_in01 = reg_0630;
    99: op1_10_in01 = reg_0156;
    100: op1_10_in01 = reg_0175;
    101: op1_10_in01 = reg_0926;
    102: op1_10_in01 = reg_0180;
    103: op1_10_in01 = imem05_in[11:8];
    47: op1_10_in01 = reg_0648;
    105: op1_10_in01 = reg_0586;
    106: op1_10_in01 = reg_0402;
    107: op1_10_in01 = reg_0138;
    108: op1_10_in01 = reg_0391;
    109: op1_10_in01 = imem05_in[7:4];
    110: op1_10_in01 = reg_0043;
    111: op1_10_in01 = reg_0303;
    112: op1_10_in01 = reg_1491;
    113: op1_10_in01 = reg_0118;
    114: op1_10_in01 = reg_0217;
    115: op1_10_in01 = reg_0192;
    116: op1_10_in01 = reg_0934;
    117: op1_10_in01 = reg_0152;
    118: op1_10_in01 = reg_0428;
    119: op1_10_in01 = reg_0054;
    120: op1_10_in01 = reg_0042;
    121: op1_10_in01 = reg_0032;
    122: op1_10_in01 = reg_0897;
    123: op1_10_in01 = reg_0206;
    34: op1_10_in01 = reg_0408;
    124: op1_10_in01 = reg_0210;
    125: op1_10_in01 = reg_1277;
    126: op1_10_in01 = reg_0381;
    127: op1_10_in01 = imem02_in[3:0];
    38: op1_10_in01 = reg_0740;
    128: op1_10_in01 = reg_0227;
    129: op1_10_in01 = reg_0488;
    130: op1_10_in01 = reg_0805;
    42: op1_10_in01 = reg_0167;
    131: op1_10_in01 = reg_0885;
    default: op1_10_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv01 = 1;
    86: op1_10_inv01 = 1;
    73: op1_10_inv01 = 1;
    69: op1_10_inv01 = 1;
    49: op1_10_inv01 = 1;
    74: op1_10_inv01 = 1;
    68: op1_10_inv01 = 1;
    75: op1_10_inv01 = 1;
    50: op1_10_inv01 = 1;
    71: op1_10_inv01 = 1;
    57: op1_10_inv01 = 1;
    77: op1_10_inv01 = 1;
    58: op1_10_inv01 = 1;
    78: op1_10_inv01 = 1;
    70: op1_10_inv01 = 1;
    51: op1_10_inv01 = 1;
    88: op1_10_inv01 = 1;
    46: op1_10_inv01 = 1;
    63: op1_10_inv01 = 1;
    89: op1_10_inv01 = 1;
    84: op1_10_inv01 = 1;
    48: op1_10_inv01 = 1;
    85: op1_10_inv01 = 1;
    65: op1_10_inv01 = 1;
    90: op1_10_inv01 = 1;
    67: op1_10_inv01 = 1;
    97: op1_10_inv01 = 1;
    100: op1_10_inv01 = 1;
    101: op1_10_inv01 = 1;
    102: op1_10_inv01 = 1;
    105: op1_10_inv01 = 1;
    108: op1_10_inv01 = 1;
    109: op1_10_inv01 = 1;
    112: op1_10_inv01 = 1;
    114: op1_10_inv01 = 1;
    117: op1_10_inv01 = 1;
    118: op1_10_inv01 = 1;
    120: op1_10_inv01 = 1;
    122: op1_10_inv01 = 1;
    123: op1_10_inv01 = 1;
    34: op1_10_inv01 = 1;
    126: op1_10_inv01 = 1;
    127: op1_10_inv01 = 1;
    128: op1_10_inv01 = 1;
    129: op1_10_inv01 = 1;
    131: op1_10_inv01 = 1;
    default: op1_10_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in02 = reg_0117;
    53: op1_10_in02 = reg_0488;
    86: op1_10_in02 = reg_0006;
    55: op1_10_in02 = imem04_in[3:0];
    73: op1_10_in02 = reg_0182;
    108: op1_10_in02 = reg_0182;
    69: op1_10_in02 = imem03_in[7:4];
    49: op1_10_in02 = reg_0323;
    74: op1_10_in02 = reg_1323;
    82: op1_10_in02 = reg_1323;
    54: op1_10_in02 = reg_0578;
    68: op1_10_in02 = reg_0957;
    75: op1_10_in02 = imem00_in[3:0];
    71: op1_10_in02 = imem00_in[3:0];
    50: op1_10_in02 = reg_0548;
    56: op1_10_in02 = reg_0336;
    87: op1_10_in02 = reg_0088;
    76: op1_10_in02 = reg_0648;
    61: op1_10_in02 = reg_0293;
    57: op1_10_in02 = reg_0720;
    77: op1_10_in02 = reg_0791;
    58: op1_10_in02 = reg_0363;
    78: op1_10_in02 = reg_0799;
    70: op1_10_in02 = reg_0329;
    79: op1_10_in02 = reg_0702;
    51: op1_10_in02 = reg_0394;
    59: op1_10_in02 = reg_0342;
    60: op1_10_in02 = reg_0742;
    88: op1_10_in02 = reg_0313;
    46: op1_10_in02 = reg_0625;
    80: op1_10_in02 = reg_0562;
    81: op1_10_in02 = reg_0095;
    52: op1_10_in02 = reg_0299;
    63: op1_10_in02 = reg_0230;
    89: op1_10_in02 = reg_0989;
    33: op1_10_in02 = reg_0361;
    83: op1_10_in02 = reg_0841;
    64: op1_10_in02 = reg_0608;
    84: op1_10_in02 = reg_0042;
    48: op1_10_in02 = reg_0193;
    85: op1_10_in02 = reg_0938;
    65: op1_10_in02 = reg_0667;
    90: op1_10_in02 = reg_1277;
    66: op1_10_in02 = reg_1032;
    37: op1_10_in02 = reg_0618;
    91: op1_10_in02 = reg_0198;
    28: op1_10_in02 = reg_0050;
    67: op1_10_in02 = reg_0672;
    92: op1_10_in02 = reg_1009;
    93: op1_10_in02 = reg_1184;
    94: op1_10_in02 = reg_0896;
    95: op1_10_in02 = reg_0804;
    96: op1_10_in02 = reg_1098;
    97: op1_10_in02 = reg_0845;
    98: op1_10_in02 = reg_1181;
    99: op1_10_in02 = reg_0924;
    100: op1_10_in02 = reg_0162;
    101: op1_10_in02 = reg_1278;
    102: op1_10_in02 = reg_1494;
    103: op1_10_in02 = reg_0090;
    104: op1_10_in02 = reg_0213;
    47: op1_10_in02 = reg_0565;
    105: op1_10_in02 = reg_0624;
    106: op1_10_in02 = reg_0634;
    44: op1_10_in02 = reg_0735;
    107: op1_10_in02 = reg_0712;
    109: op1_10_in02 = reg_0833;
    110: op1_10_in02 = reg_0895;
    111: op1_10_in02 = reg_0872;
    112: op1_10_in02 = reg_0153;
    113: op1_10_in02 = reg_0575;
    114: op1_10_in02 = reg_0479;
    115: op1_10_in02 = reg_0870;
    116: op1_10_in02 = reg_0055;
    117: op1_10_in02 = reg_0214;
    118: op1_10_in02 = reg_0410;
    119: op1_10_in02 = reg_0778;
    120: op1_10_in02 = reg_0010;
    121: op1_10_in02 = reg_0337;
    122: op1_10_in02 = reg_0560;
    123: op1_10_in02 = imem06_in[15:12];
    34: op1_10_in02 = reg_0413;
    124: op1_10_in02 = reg_0567;
    125: op1_10_in02 = reg_0501;
    126: op1_10_in02 = reg_0306;
    127: op1_10_in02 = reg_0138;
    38: op1_10_in02 = reg_0620;
    128: op1_10_in02 = reg_0168;
    129: op1_10_in02 = reg_1215;
    130: op1_10_in02 = reg_0523;
    42: op1_10_in02 = reg_0120;
    131: op1_10_in02 = reg_0448;
    default: op1_10_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv02 = 1;
    55: op1_10_inv02 = 1;
    54: op1_10_inv02 = 1;
    68: op1_10_inv02 = 1;
    50: op1_10_inv02 = 1;
    56: op1_10_inv02 = 1;
    87: op1_10_inv02 = 1;
    76: op1_10_inv02 = 1;
    61: op1_10_inv02 = 1;
    57: op1_10_inv02 = 1;
    58: op1_10_inv02 = 1;
    78: op1_10_inv02 = 1;
    51: op1_10_inv02 = 1;
    82: op1_10_inv02 = 1;
    84: op1_10_inv02 = 1;
    65: op1_10_inv02 = 1;
    66: op1_10_inv02 = 1;
    28: op1_10_inv02 = 1;
    94: op1_10_inv02 = 1;
    95: op1_10_inv02 = 1;
    96: op1_10_inv02 = 1;
    98: op1_10_inv02 = 1;
    100: op1_10_inv02 = 1;
    102: op1_10_inv02 = 1;
    47: op1_10_inv02 = 1;
    105: op1_10_inv02 = 1;
    107: op1_10_inv02 = 1;
    108: op1_10_inv02 = 1;
    109: op1_10_inv02 = 1;
    110: op1_10_inv02 = 1;
    111: op1_10_inv02 = 1;
    113: op1_10_inv02 = 1;
    129: op1_10_inv02 = 1;
    42: op1_10_inv02 = 1;
    default: op1_10_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in03 = reg_0129;
    53: op1_10_in03 = reg_0596;
    86: op1_10_in03 = reg_1132;
    55: op1_10_in03 = reg_1065;
    73: op1_10_in03 = reg_1401;
    69: op1_10_in03 = reg_1033;
    49: op1_10_in03 = reg_0296;
    74: op1_10_in03 = reg_0984;
    54: op1_10_in03 = reg_0749;
    68: op1_10_in03 = reg_0952;
    75: op1_10_in03 = imem00_in[7:4];
    50: op1_10_in03 = reg_0260;
    56: op1_10_in03 = reg_0065;
    71: op1_10_in03 = reg_1052;
    87: op1_10_in03 = reg_0978;
    76: op1_10_in03 = reg_0650;
    61: op1_10_in03 = reg_1028;
    130: op1_10_in03 = reg_1028;
    57: op1_10_in03 = reg_0825;
    77: op1_10_in03 = reg_0983;
    58: op1_10_in03 = reg_0901;
    78: op1_10_in03 = reg_1035;
    82: op1_10_in03 = reg_1035;
    70: op1_10_in03 = reg_0558;
    79: op1_10_in03 = reg_0136;
    51: op1_10_in03 = reg_0191;
    59: op1_10_in03 = reg_0262;
    60: op1_10_in03 = reg_0744;
    88: op1_10_in03 = reg_1139;
    46: op1_10_in03 = reg_0536;
    80: op1_10_in03 = reg_1510;
    81: op1_10_in03 = reg_0019;
    52: op1_10_in03 = reg_0186;
    112: op1_10_in03 = reg_0186;
    63: op1_10_in03 = reg_0490;
    89: op1_10_in03 = reg_0314;
    33: op1_10_in03 = reg_0003;
    83: op1_10_in03 = reg_1471;
    64: op1_10_in03 = reg_0169;
    84: op1_10_in03 = reg_0895;
    48: op1_10_in03 = imem06_in[11:8];
    85: op1_10_in03 = reg_0418;
    65: op1_10_in03 = imem07_in[11:8];
    28: op1_10_in03 = imem07_in[11:8];
    90: op1_10_in03 = reg_0672;
    66: op1_10_in03 = reg_0161;
    37: op1_10_in03 = reg_0102;
    91: op1_10_in03 = reg_1001;
    67: op1_10_in03 = reg_0669;
    92: op1_10_in03 = reg_0025;
    93: op1_10_in03 = reg_1516;
    94: op1_10_in03 = reg_0120;
    95: op1_10_in03 = reg_0805;
    96: op1_10_in03 = reg_0007;
    97: op1_10_in03 = reg_0608;
    98: op1_10_in03 = reg_1402;
    99: op1_10_in03 = reg_0139;
    100: op1_10_in03 = reg_0402;
    101: op1_10_in03 = reg_1279;
    102: op1_10_in03 = reg_1495;
    103: op1_10_in03 = reg_0492;
    104: op1_10_in03 = reg_0394;
    47: op1_10_in03 = reg_0566;
    105: op1_10_in03 = reg_0570;
    106: op1_10_in03 = reg_1068;
    120: op1_10_in03 = reg_1068;
    44: op1_10_in03 = reg_0702;
    107: op1_10_in03 = reg_0472;
    108: op1_10_in03 = reg_0334;
    109: op1_10_in03 = reg_0333;
    110: op1_10_in03 = reg_0447;
    111: op1_10_in03 = reg_0318;
    113: op1_10_in03 = reg_1346;
    114: op1_10_in03 = reg_0507;
    115: op1_10_in03 = reg_0730;
    116: op1_10_in03 = reg_0975;
    117: op1_10_in03 = reg_1170;
    118: op1_10_in03 = reg_0071;
    119: op1_10_in03 = reg_1455;
    121: op1_10_in03 = reg_0731;
    122: op1_10_in03 = reg_0802;
    126: op1_10_in03 = reg_0802;
    123: op1_10_in03 = reg_0729;
    34: op1_10_in03 = reg_0621;
    124: op1_10_in03 = reg_1259;
    125: op1_10_in03 = reg_0554;
    127: op1_10_in03 = reg_0934;
    38: op1_10_in03 = reg_0002;
    128: op1_10_in03 = reg_0759;
    129: op1_10_in03 = reg_0407;
    42: op1_10_in03 = reg_0259;
    131: op1_10_in03 = reg_0350;
    default: op1_10_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv03 = 1;
    73: op1_10_inv03 = 1;
    69: op1_10_inv03 = 1;
    75: op1_10_inv03 = 1;
    50: op1_10_inv03 = 1;
    87: op1_10_inv03 = 1;
    76: op1_10_inv03 = 1;
    58: op1_10_inv03 = 1;
    78: op1_10_inv03 = 1;
    79: op1_10_inv03 = 1;
    88: op1_10_inv03 = 1;
    46: op1_10_inv03 = 1;
    80: op1_10_inv03 = 1;
    52: op1_10_inv03 = 1;
    63: op1_10_inv03 = 1;
    82: op1_10_inv03 = 1;
    33: op1_10_inv03 = 1;
    64: op1_10_inv03 = 1;
    48: op1_10_inv03 = 1;
    66: op1_10_inv03 = 1;
    37: op1_10_inv03 = 1;
    91: op1_10_inv03 = 1;
    93: op1_10_inv03 = 1;
    94: op1_10_inv03 = 1;
    96: op1_10_inv03 = 1;
    98: op1_10_inv03 = 1;
    101: op1_10_inv03 = 1;
    102: op1_10_inv03 = 1;
    106: op1_10_inv03 = 1;
    107: op1_10_inv03 = 1;
    108: op1_10_inv03 = 1;
    110: op1_10_inv03 = 1;
    111: op1_10_inv03 = 1;
    112: op1_10_inv03 = 1;
    113: op1_10_inv03 = 1;
    116: op1_10_inv03 = 1;
    117: op1_10_inv03 = 1;
    118: op1_10_inv03 = 1;
    119: op1_10_inv03 = 1;
    121: op1_10_inv03 = 1;
    34: op1_10_inv03 = 1;
    125: op1_10_inv03 = 1;
    42: op1_10_inv03 = 1;
    default: op1_10_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in04 = reg_0064;
    53: op1_10_in04 = reg_0304;
    86: op1_10_in04 = reg_1000;
    55: op1_10_in04 = reg_1082;
    73: op1_10_in04 = reg_0938;
    69: op1_10_in04 = reg_0638;
    49: op1_10_in04 = reg_0295;
    74: op1_10_in04 = reg_0115;
    57: op1_10_in04 = reg_0115;
    54: op1_10_in04 = reg_0750;
    68: op1_10_in04 = reg_0190;
    75: op1_10_in04 = imem00_in[11:8];
    50: op1_10_in04 = reg_0258;
    56: op1_10_in04 = reg_0033;
    71: op1_10_in04 = reg_0887;
    87: op1_10_in04 = reg_0531;
    76: op1_10_in04 = reg_0131;
    61: op1_10_in04 = reg_1027;
    77: op1_10_in04 = reg_1510;
    58: op1_10_in04 = reg_0277;
    78: op1_10_in04 = reg_1467;
    70: op1_10_in04 = reg_1226;
    79: op1_10_in04 = reg_0992;
    51: op1_10_in04 = imem07_in[7:4];
    117: op1_10_in04 = imem07_in[7:4];
    59: op1_10_in04 = reg_0837;
    60: op1_10_in04 = reg_0608;
    88: op1_10_in04 = reg_1282;
    46: op1_10_in04 = reg_0493;
    80: op1_10_in04 = reg_1490;
    81: op1_10_in04 = reg_0470;
    52: op1_10_in04 = reg_0921;
    63: op1_10_in04 = reg_0667;
    82: op1_10_in04 = reg_0141;
    89: op1_10_in04 = reg_0627;
    33: op1_10_in04 = reg_0087;
    83: op1_10_in04 = reg_0293;
    64: op1_10_in04 = reg_0253;
    84: op1_10_in04 = reg_1493;
    48: op1_10_in04 = reg_0133;
    85: op1_10_in04 = reg_0303;
    65: op1_10_in04 = reg_0187;
    90: op1_10_in04 = reg_0501;
    66: op1_10_in04 = reg_0982;
    37: op1_10_in04 = reg_0103;
    91: op1_10_in04 = reg_0375;
    67: op1_10_in04 = reg_0842;
    92: op1_10_in04 = reg_0313;
    131: op1_10_in04 = reg_0313;
    93: op1_10_in04 = reg_0558;
    94: op1_10_in04 = reg_0044;
    95: op1_10_in04 = reg_0250;
    125: op1_10_in04 = reg_0250;
    96: op1_10_in04 = reg_1006;
    97: op1_10_in04 = reg_0588;
    98: op1_10_in04 = reg_1070;
    99: op1_10_in04 = reg_0465;
    100: op1_10_in04 = reg_0895;
    101: op1_10_in04 = reg_0580;
    102: op1_10_in04 = reg_0142;
    103: op1_10_in04 = reg_1373;
    104: op1_10_in04 = reg_0498;
    47: op1_10_in04 = reg_0045;
    105: op1_10_in04 = reg_1228;
    106: op1_10_in04 = reg_0447;
    44: op1_10_in04 = reg_0649;
    107: op1_10_in04 = reg_0432;
    108: op1_10_in04 = reg_1401;
    109: op1_10_in04 = reg_0346;
    110: op1_10_in04 = reg_1071;
    111: op1_10_in04 = reg_0589;
    112: op1_10_in04 = reg_1028;
    113: op1_10_in04 = reg_0039;
    114: op1_10_in04 = reg_0600;
    115: op1_10_in04 = reg_0271;
    116: op1_10_in04 = reg_0494;
    118: op1_10_in04 = reg_0203;
    119: op1_10_in04 = reg_0126;
    120: op1_10_in04 = imem02_in[3:0];
    121: op1_10_in04 = reg_0297;
    122: op1_10_in04 = reg_0695;
    123: op1_10_in04 = reg_0669;
    34: op1_10_in04 = reg_0137;
    124: op1_10_in04 = reg_1164;
    126: op1_10_in04 = reg_1098;
    127: op1_10_in04 = reg_0561;
    38: op1_10_in04 = reg_0085;
    128: op1_10_in04 = reg_0233;
    129: op1_10_in04 = reg_0598;
    130: op1_10_in04 = reg_1206;
    42: op1_10_in04 = reg_0241;
    default: op1_10_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_10_inv04 = 1;
    55: op1_10_inv04 = 1;
    69: op1_10_inv04 = 1;
    50: op1_10_inv04 = 1;
    76: op1_10_inv04 = 1;
    61: op1_10_inv04 = 1;
    57: op1_10_inv04 = 1;
    77: op1_10_inv04 = 1;
    78: op1_10_inv04 = 1;
    70: op1_10_inv04 = 1;
    79: op1_10_inv04 = 1;
    51: op1_10_inv04 = 1;
    88: op1_10_inv04 = 1;
    82: op1_10_inv04 = 1;
    33: op1_10_inv04 = 1;
    83: op1_10_inv04 = 1;
    90: op1_10_inv04 = 1;
    92: op1_10_inv04 = 1;
    93: op1_10_inv04 = 1;
    94: op1_10_inv04 = 1;
    95: op1_10_inv04 = 1;
    98: op1_10_inv04 = 1;
    100: op1_10_inv04 = 1;
    104: op1_10_inv04 = 1;
    47: op1_10_inv04 = 1;
    105: op1_10_inv04 = 1;
    44: op1_10_inv04 = 1;
    108: op1_10_inv04 = 1;
    110: op1_10_inv04 = 1;
    111: op1_10_inv04 = 1;
    112: op1_10_inv04 = 1;
    113: op1_10_inv04 = 1;
    114: op1_10_inv04 = 1;
    117: op1_10_inv04 = 1;
    121: op1_10_inv04 = 1;
    123: op1_10_inv04 = 1;
    126: op1_10_inv04 = 1;
    127: op1_10_inv04 = 1;
    38: op1_10_inv04 = 1;
    129: op1_10_inv04 = 1;
    130: op1_10_inv04 = 1;
    42: op1_10_inv04 = 1;
    default: op1_10_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in05 = reg_0063;
    53: op1_10_in05 = reg_0837;
    86: op1_10_in05 = reg_0233;
    55: op1_10_in05 = reg_0420;
    73: op1_10_in05 = reg_0477;
    69: op1_10_in05 = reg_0891;
    49: op1_10_in05 = reg_0289;
    74: op1_10_in05 = reg_0717;
    54: op1_10_in05 = reg_1059;
    68: op1_10_in05 = reg_1300;
    75: op1_10_in05 = reg_1278;
    50: op1_10_in05 = reg_0239;
    56: op1_10_in05 = reg_0034;
    71: op1_10_in05 = reg_0351;
    87: op1_10_in05 = reg_1233;
    76: op1_10_in05 = reg_0334;
    47: op1_10_in05 = reg_0334;
    61: op1_10_in05 = reg_1227;
    57: op1_10_in05 = reg_0671;
    77: op1_10_in05 = reg_1277;
    58: op1_10_in05 = reg_0278;
    78: op1_10_in05 = reg_0906;
    70: op1_10_in05 = reg_1199;
    79: op1_10_in05 = reg_0173;
    51: op1_10_in05 = imem07_in[11:8];
    59: op1_10_in05 = reg_0094;
    60: op1_10_in05 = reg_1018;
    88: op1_10_in05 = reg_0975;
    127: op1_10_in05 = reg_0975;
    46: op1_10_in05 = reg_0731;
    80: op1_10_in05 = reg_1241;
    81: op1_10_in05 = reg_0175;
    52: op1_10_in05 = reg_0924;
    63: op1_10_in05 = reg_0892;
    82: op1_10_in05 = reg_0619;
    89: op1_10_in05 = reg_0957;
    33: op1_10_in05 = reg_0123;
    83: op1_10_in05 = reg_0221;
    125: op1_10_in05 = reg_0221;
    64: op1_10_in05 = reg_0456;
    84: op1_10_in05 = reg_1343;
    48: op1_10_in05 = reg_0979;
    85: op1_10_in05 = reg_0302;
    65: op1_10_in05 = reg_0299;
    90: op1_10_in05 = reg_0153;
    66: op1_10_in05 = reg_0469;
    37: op1_10_in05 = reg_0321;
    91: op1_10_in05 = reg_0070;
    67: op1_10_in05 = reg_1053;
    92: op1_10_in05 = reg_0467;
    93: op1_10_in05 = reg_1093;
    94: op1_10_in05 = reg_0041;
    95: op1_10_in05 = reg_1028;
    101: op1_10_in05 = reg_1028;
    96: op1_10_in05 = reg_0069;
    97: op1_10_in05 = reg_0497;
    98: op1_10_in05 = reg_0938;
    99: op1_10_in05 = reg_0030;
    100: op1_10_in05 = imem02_in[7:4];
    102: op1_10_in05 = reg_1518;
    103: op1_10_in05 = reg_0274;
    104: op1_10_in05 = reg_1315;
    105: op1_10_in05 = reg_1225;
    106: op1_10_in05 = reg_0845;
    44: op1_10_in05 = reg_0317;
    107: op1_10_in05 = reg_0429;
    108: op1_10_in05 = reg_0939;
    109: op1_10_in05 = reg_0272;
    110: op1_10_in05 = reg_1344;
    111: op1_10_in05 = reg_0828;
    112: op1_10_in05 = reg_1205;
    113: op1_10_in05 = imem06_in[11:8];
    114: op1_10_in05 = reg_0143;
    115: op1_10_in05 = reg_0863;
    116: op1_10_in05 = reg_0971;
    117: op1_10_in05 = reg_0893;
    118: op1_10_in05 = reg_0075;
    119: op1_10_in05 = reg_0105;
    120: op1_10_in05 = reg_0099;
    121: op1_10_in05 = reg_1200;
    122: op1_10_in05 = reg_1006;
    123: op1_10_in05 = reg_0397;
    34: op1_10_in05 = reg_0102;
    124: op1_10_in05 = reg_0340;
    126: op1_10_in05 = reg_0800;
    38: op1_10_in05 = reg_0084;
    128: op1_10_in05 = reg_1009;
    129: op1_10_in05 = reg_1041;
    130: op1_10_in05 = reg_1432;
    42: op1_10_in05 = reg_0746;
    131: op1_10_in05 = reg_0035;
    default: op1_10_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv05 = 1;
    53: op1_10_inv05 = 1;
    86: op1_10_inv05 = 1;
    55: op1_10_inv05 = 1;
    73: op1_10_inv05 = 1;
    74: op1_10_inv05 = 1;
    68: op1_10_inv05 = 1;
    50: op1_10_inv05 = 1;
    56: op1_10_inv05 = 1;
    71: op1_10_inv05 = 1;
    87: op1_10_inv05 = 1;
    76: op1_10_inv05 = 1;
    61: op1_10_inv05 = 1;
    57: op1_10_inv05 = 1;
    58: op1_10_inv05 = 1;
    79: op1_10_inv05 = 1;
    51: op1_10_inv05 = 1;
    60: op1_10_inv05 = 1;
    88: op1_10_inv05 = 1;
    46: op1_10_inv05 = 1;
    80: op1_10_inv05 = 1;
    81: op1_10_inv05 = 1;
    33: op1_10_inv05 = 1;
    83: op1_10_inv05 = 1;
    48: op1_10_inv05 = 1;
    85: op1_10_inv05 = 1;
    66: op1_10_inv05 = 1;
    37: op1_10_inv05 = 1;
    91: op1_10_inv05 = 1;
    67: op1_10_inv05 = 1;
    93: op1_10_inv05 = 1;
    97: op1_10_inv05 = 1;
    98: op1_10_inv05 = 1;
    100: op1_10_inv05 = 1;
    104: op1_10_inv05 = 1;
    47: op1_10_inv05 = 1;
    44: op1_10_inv05 = 1;
    109: op1_10_inv05 = 1;
    111: op1_10_inv05 = 1;
    112: op1_10_inv05 = 1;
    113: op1_10_inv05 = 1;
    115: op1_10_inv05 = 1;
    116: op1_10_inv05 = 1;
    119: op1_10_inv05 = 1;
    120: op1_10_inv05 = 1;
    121: op1_10_inv05 = 1;
    123: op1_10_inv05 = 1;
    125: op1_10_inv05 = 1;
    42: op1_10_inv05 = 1;
    default: op1_10_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in06 = reg_0204;
    53: op1_10_in06 = reg_0719;
    86: op1_10_in06 = reg_0709;
    55: op1_10_in06 = reg_0421;
    73: op1_10_in06 = reg_0196;
    69: op1_10_in06 = reg_0261;
    49: op1_10_in06 = reg_0271;
    74: op1_10_in06 = reg_1302;
    54: op1_10_in06 = reg_0345;
    68: op1_10_in06 = reg_1208;
    75: op1_10_in06 = reg_1079;
    50: op1_10_in06 = reg_0238;
    56: op1_10_in06 = reg_0794;
    71: op1_10_in06 = reg_0352;
    87: op1_10_in06 = reg_1214;
    76: op1_10_in06 = reg_1181;
    61: op1_10_in06 = reg_0203;
    57: op1_10_in06 = reg_0635;
    77: op1_10_in06 = reg_1241;
    58: op1_10_in06 = reg_0041;
    78: op1_10_in06 = reg_0120;
    70: op1_10_in06 = reg_0479;
    79: op1_10_in06 = reg_0346;
    51: op1_10_in06 = reg_1057;
    59: op1_10_in06 = reg_0181;
    60: op1_10_in06 = reg_0590;
    88: op1_10_in06 = reg_0208;
    46: op1_10_in06 = reg_0698;
    80: op1_10_in06 = reg_0841;
    81: op1_10_in06 = reg_0736;
    108: op1_10_in06 = reg_0736;
    52: op1_10_in06 = reg_0923;
    63: op1_10_in06 = reg_0309;
    82: op1_10_in06 = reg_0617;
    89: op1_10_in06 = reg_0190;
    83: op1_10_in06 = reg_1230;
    64: op1_10_in06 = reg_0562;
    84: op1_10_in06 = reg_0532;
    127: op1_10_in06 = reg_0532;
    48: op1_10_in06 = reg_0730;
    85: op1_10_in06 = reg_1484;
    65: op1_10_in06 = reg_0170;
    90: op1_10_in06 = reg_0616;
    66: op1_10_in06 = reg_0146;
    37: op1_10_in06 = reg_0050;
    91: op1_10_in06 = reg_1314;
    67: op1_10_in06 = reg_1052;
    92: op1_10_in06 = reg_0237;
    93: op1_10_in06 = reg_1092;
    94: op1_10_in06 = reg_0895;
    95: op1_10_in06 = reg_1027;
    96: op1_10_in06 = reg_0255;
    97: op1_10_in06 = reg_1002;
    98: op1_10_in06 = reg_0183;
    99: op1_10_in06 = reg_0665;
    100: op1_10_in06 = reg_0530;
    101: op1_10_in06 = reg_1229;
    102: op1_10_in06 = reg_0220;
    103: op1_10_in06 = reg_0118;
    104: op1_10_in06 = reg_0298;
    47: op1_10_in06 = reg_0316;
    105: op1_10_in06 = reg_0419;
    106: op1_10_in06 = reg_0276;
    44: op1_10_in06 = reg_0367;
    107: op1_10_in06 = reg_0970;
    109: op1_10_in06 = reg_0251;
    110: op1_10_in06 = reg_0721;
    111: op1_10_in06 = reg_0317;
    112: op1_10_in06 = reg_1432;
    113: op1_10_in06 = reg_0795;
    114: op1_10_in06 = reg_1495;
    115: op1_10_in06 = reg_0859;
    116: op1_10_in06 = reg_0112;
    117: op1_10_in06 = reg_0051;
    118: op1_10_in06 = reg_0060;
    119: op1_10_in06 = reg_0631;
    120: op1_10_in06 = reg_0138;
    121: op1_10_in06 = reg_0488;
    122: op1_10_in06 = reg_0168;
    123: op1_10_in06 = reg_0925;
    34: op1_10_in06 = reg_0114;
    124: op1_10_in06 = reg_0167;
    125: op1_10_in06 = reg_0155;
    126: op1_10_in06 = reg_1078;
    38: op1_10_in06 = reg_0087;
    128: op1_10_in06 = reg_0732;
    129: op1_10_in06 = reg_0537;
    130: op1_10_in06 = reg_1405;
    42: op1_10_in06 = reg_0726;
    131: op1_10_in06 = reg_0319;
    default: op1_10_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv06 = 1;
    53: op1_10_inv06 = 1;
    86: op1_10_inv06 = 1;
    73: op1_10_inv06 = 1;
    49: op1_10_inv06 = 1;
    74: op1_10_inv06 = 1;
    50: op1_10_inv06 = 1;
    76: op1_10_inv06 = 1;
    70: op1_10_inv06 = 1;
    59: op1_10_inv06 = 1;
    80: op1_10_inv06 = 1;
    81: op1_10_inv06 = 1;
    52: op1_10_inv06 = 1;
    82: op1_10_inv06 = 1;
    89: op1_10_inv06 = 1;
    84: op1_10_inv06 = 1;
    90: op1_10_inv06 = 1;
    66: op1_10_inv06 = 1;
    37: op1_10_inv06 = 1;
    91: op1_10_inv06 = 1;
    94: op1_10_inv06 = 1;
    96: op1_10_inv06 = 1;
    98: op1_10_inv06 = 1;
    99: op1_10_inv06 = 1;
    100: op1_10_inv06 = 1;
    101: op1_10_inv06 = 1;
    102: op1_10_inv06 = 1;
    103: op1_10_inv06 = 1;
    106: op1_10_inv06 = 1;
    108: op1_10_inv06 = 1;
    109: op1_10_inv06 = 1;
    112: op1_10_inv06 = 1;
    113: op1_10_inv06 = 1;
    118: op1_10_inv06 = 1;
    120: op1_10_inv06 = 1;
    121: op1_10_inv06 = 1;
    34: op1_10_inv06 = 1;
    125: op1_10_inv06 = 1;
    38: op1_10_inv06 = 1;
    128: op1_10_inv06 = 1;
    130: op1_10_inv06 = 1;
    default: op1_10_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in07 = reg_1431;
    53: op1_10_in07 = reg_0094;
    86: op1_10_in07 = reg_1001;
    55: op1_10_in07 = reg_0412;
    73: op1_10_in07 = reg_0799;
    69: op1_10_in07 = reg_0999;
    49: op1_10_in07 = reg_0213;
    74: op1_10_in07 = reg_0141;
    54: op1_10_in07 = reg_1169;
    68: op1_10_in07 = reg_0107;
    75: op1_10_in07 = reg_1080;
    50: op1_10_in07 = reg_0980;
    56: op1_10_in07 = reg_0631;
    71: op1_10_in07 = reg_0405;
    87: op1_10_in07 = reg_0796;
    76: op1_10_in07 = reg_0697;
    61: op1_10_in07 = reg_0460;
    83: op1_10_in07 = reg_0460;
    57: op1_10_in07 = reg_0636;
    77: op1_10_in07 = reg_0562;
    58: op1_10_in07 = reg_0446;
    78: op1_10_in07 = reg_0870;
    70: op1_10_in07 = reg_0573;
    79: op1_10_in07 = reg_0174;
    51: op1_10_in07 = reg_0993;
    59: op1_10_in07 = reg_0117;
    60: op1_10_in07 = reg_0561;
    64: op1_10_in07 = reg_0561;
    88: op1_10_in07 = reg_0032;
    46: op1_10_in07 = reg_0633;
    80: op1_10_in07 = reg_0293;
    81: op1_10_in07 = reg_0579;
    52: op1_10_in07 = reg_0777;
    63: op1_10_in07 = imem07_in[7:4];
    82: op1_10_in07 = reg_0569;
    89: op1_10_in07 = reg_1226;
    91: op1_10_in07 = reg_1226;
    84: op1_10_in07 = reg_0474;
    48: op1_10_in07 = reg_0860;
    85: op1_10_in07 = reg_0492;
    65: op1_10_in07 = reg_1347;
    90: op1_10_in07 = reg_0486;
    66: op1_10_in07 = reg_0091;
    37: op1_10_in07 = reg_0051;
    67: op1_10_in07 = reg_0987;
    92: op1_10_in07 = reg_0577;
    93: op1_10_in07 = reg_0104;
    94: op1_10_in07 = reg_0666;
    95: op1_10_in07 = reg_0249;
    96: op1_10_in07 = reg_0632;
    97: op1_10_in07 = reg_0973;
    98: op1_10_in07 = reg_0477;
    99: op1_10_in07 = reg_0739;
    100: op1_10_in07 = reg_0254;
    101: op1_10_in07 = reg_1201;
    102: op1_10_in07 = reg_1231;
    103: op1_10_in07 = reg_1346;
    104: op1_10_in07 = reg_0892;
    47: op1_10_in07 = reg_0318;
    105: op1_10_in07 = reg_0583;
    106: op1_10_in07 = reg_1493;
    44: op1_10_in07 = reg_0896;
    107: op1_10_in07 = reg_0125;
    108: op1_10_in07 = reg_0450;
    109: op1_10_in07 = reg_0996;
    110: op1_10_in07 = reg_0530;
    111: op1_10_in07 = reg_0038;
    112: op1_10_in07 = reg_0524;
    113: op1_10_in07 = reg_0925;
    114: op1_10_in07 = reg_1516;
    115: op1_10_in07 = reg_0827;
    116: op1_10_in07 = reg_1140;
    117: op1_10_in07 = reg_0084;
    118: op1_10_in07 = reg_0269;
    119: op1_10_in07 = reg_0306;
    120: op1_10_in07 = reg_0975;
    121: op1_10_in07 = reg_0281;
    122: op1_10_in07 = reg_1515;
    123: op1_10_in07 = reg_0869;
    34: op1_10_in07 = reg_0050;
    124: op1_10_in07 = reg_0630;
    125: op1_10_in07 = reg_0351;
    126: op1_10_in07 = reg_0006;
    127: op1_10_in07 = reg_0898;
    38: op1_10_in07 = reg_0484;
    128: op1_10_in07 = reg_0049;
    129: op1_10_in07 = reg_1040;
    130: op1_10_in07 = reg_0928;
    42: op1_10_in07 = reg_0727;
    131: op1_10_in07 = reg_0164;
    default: op1_10_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv07 = 1;
    86: op1_10_inv07 = 1;
    55: op1_10_inv07 = 1;
    69: op1_10_inv07 = 1;
    74: op1_10_inv07 = 1;
    54: op1_10_inv07 = 1;
    68: op1_10_inv07 = 1;
    50: op1_10_inv07 = 1;
    71: op1_10_inv07 = 1;
    87: op1_10_inv07 = 1;
    70: op1_10_inv07 = 1;
    79: op1_10_inv07 = 1;
    51: op1_10_inv07 = 1;
    60: op1_10_inv07 = 1;
    46: op1_10_inv07 = 1;
    52: op1_10_inv07 = 1;
    63: op1_10_inv07 = 1;
    82: op1_10_inv07 = 1;
    83: op1_10_inv07 = 1;
    84: op1_10_inv07 = 1;
    48: op1_10_inv07 = 1;
    85: op1_10_inv07 = 1;
    65: op1_10_inv07 = 1;
    90: op1_10_inv07 = 1;
    91: op1_10_inv07 = 1;
    92: op1_10_inv07 = 1;
    93: op1_10_inv07 = 1;
    97: op1_10_inv07 = 1;
    99: op1_10_inv07 = 1;
    101: op1_10_inv07 = 1;
    104: op1_10_inv07 = 1;
    47: op1_10_inv07 = 1;
    105: op1_10_inv07 = 1;
    107: op1_10_inv07 = 1;
    109: op1_10_inv07 = 1;
    110: op1_10_inv07 = 1;
    112: op1_10_inv07 = 1;
    113: op1_10_inv07 = 1;
    114: op1_10_inv07 = 1;
    116: op1_10_inv07 = 1;
    119: op1_10_inv07 = 1;
    121: op1_10_inv07 = 1;
    122: op1_10_inv07 = 1;
    123: op1_10_inv07 = 1;
    126: op1_10_inv07 = 1;
    38: op1_10_inv07 = 1;
    128: op1_10_inv07 = 1;
    131: op1_10_inv07 = 1;
    default: op1_10_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in08 = reg_0136;
    53: op1_10_in08 = reg_0096;
    86: op1_10_in08 = reg_0541;
    55: op1_10_in08 = reg_0406;
    73: op1_10_in08 = reg_0797;
    69: op1_10_in08 = reg_1003;
    49: op1_10_in08 = reg_0162;
    74: op1_10_in08 = reg_0296;
    54: op1_10_in08 = reg_0333;
    68: op1_10_in08 = imem03_in[3:0];
    96: op1_10_in08 = imem03_in[3:0];
    75: op1_10_in08 = reg_0552;
    50: op1_10_in08 = reg_0967;
    56: op1_10_in08 = reg_0393;
    71: op1_10_in08 = reg_0073;
    87: op1_10_in08 = reg_0094;
    76: op1_10_in08 = imem05_in[15:12];
    61: op1_10_in08 = reg_0958;
    57: op1_10_in08 = reg_0264;
    77: op1_10_in08 = reg_0803;
    58: op1_10_in08 = reg_0606;
    78: op1_10_in08 = reg_0730;
    70: op1_10_in08 = reg_0328;
    79: op1_10_in08 = reg_0567;
    51: op1_10_in08 = reg_0995;
    59: op1_10_in08 = reg_0129;
    60: op1_10_in08 = reg_0612;
    88: op1_10_in08 = reg_0088;
    46: op1_10_in08 = imem04_in[7:4];
    80: op1_10_in08 = reg_0485;
    81: op1_10_in08 = reg_0833;
    52: op1_10_in08 = reg_0779;
    63: op1_10_in08 = reg_0158;
    82: op1_10_in08 = reg_0570;
    89: op1_10_in08 = reg_1208;
    83: op1_10_in08 = reg_0229;
    64: op1_10_in08 = reg_0254;
    84: op1_10_in08 = reg_1455;
    48: op1_10_in08 = reg_0859;
    85: op1_10_in08 = reg_0274;
    65: op1_10_in08 = reg_0923;
    90: op1_10_in08 = reg_0555;
    66: op1_10_in08 = reg_0092;
    37: op1_10_in08 = reg_0002;
    91: op1_10_in08 = reg_0178;
    67: op1_10_in08 = reg_0460;
    92: op1_10_in08 = reg_0263;
    93: op1_10_in08 = reg_1149;
    94: op1_10_in08 = reg_0975;
    95: op1_10_in08 = reg_0961;
    101: op1_10_in08 = reg_0961;
    97: op1_10_in08 = reg_0111;
    98: op1_10_in08 = reg_0090;
    99: op1_10_in08 = reg_0618;
    100: op1_10_in08 = reg_0822;
    102: op1_10_in08 = reg_1092;
    103: op1_10_in08 = reg_0344;
    104: op1_10_in08 = reg_0786;
    47: op1_10_in08 = reg_0163;
    105: op1_10_in08 = reg_0023;
    106: op1_10_in08 = reg_0497;
    44: op1_10_in08 = reg_0301;
    107: op1_10_in08 = reg_0105;
    108: op1_10_in08 = reg_0118;
    109: op1_10_in08 = reg_0649;
    110: op1_10_in08 = reg_0608;
    111: op1_10_in08 = reg_0161;
    112: op1_10_in08 = reg_0928;
    113: op1_10_in08 = reg_0780;
    114: op1_10_in08 = reg_1517;
    115: op1_10_in08 = reg_1505;
    116: op1_10_in08 = reg_0380;
    117: op1_10_in08 = reg_0922;
    118: op1_10_in08 = reg_1032;
    119: op1_10_in08 = reg_0897;
    120: op1_10_in08 = reg_0455;
    121: op1_10_in08 = reg_0421;
    122: op1_10_in08 = imem03_in[15:12];
    123: op1_10_in08 = reg_0109;
    34: op1_10_in08 = reg_0001;
    124: op1_10_in08 = reg_1180;
    125: op1_10_in08 = reg_0388;
    126: op1_10_in08 = imem03_in[7:4];
    127: op1_10_in08 = reg_0533;
    128: op1_10_in08 = reg_0185;
    129: op1_10_in08 = reg_0452;
    130: op1_10_in08 = reg_0202;
    42: op1_10_in08 = reg_0572;
    131: op1_10_in08 = reg_0694;
    default: op1_10_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_10_inv08 = 1;
    55: op1_10_inv08 = 1;
    73: op1_10_inv08 = 1;
    69: op1_10_inv08 = 1;
    49: op1_10_inv08 = 1;
    68: op1_10_inv08 = 1;
    50: op1_10_inv08 = 1;
    71: op1_10_inv08 = 1;
    87: op1_10_inv08 = 1;
    76: op1_10_inv08 = 1;
    57: op1_10_inv08 = 1;
    77: op1_10_inv08 = 1;
    70: op1_10_inv08 = 1;
    79: op1_10_inv08 = 1;
    46: op1_10_inv08 = 1;
    52: op1_10_inv08 = 1;
    63: op1_10_inv08 = 1;
    82: op1_10_inv08 = 1;
    89: op1_10_inv08 = 1;
    84: op1_10_inv08 = 1;
    48: op1_10_inv08 = 1;
    85: op1_10_inv08 = 1;
    90: op1_10_inv08 = 1;
    66: op1_10_inv08 = 1;
    67: op1_10_inv08 = 1;
    92: op1_10_inv08 = 1;
    93: op1_10_inv08 = 1;
    94: op1_10_inv08 = 1;
    95: op1_10_inv08 = 1;
    96: op1_10_inv08 = 1;
    98: op1_10_inv08 = 1;
    99: op1_10_inv08 = 1;
    103: op1_10_inv08 = 1;
    47: op1_10_inv08 = 1;
    105: op1_10_inv08 = 1;
    109: op1_10_inv08 = 1;
    111: op1_10_inv08 = 1;
    113: op1_10_inv08 = 1;
    115: op1_10_inv08 = 1;
    116: op1_10_inv08 = 1;
    118: op1_10_inv08 = 1;
    119: op1_10_inv08 = 1;
    120: op1_10_inv08 = 1;
    122: op1_10_inv08 = 1;
    123: op1_10_inv08 = 1;
    34: op1_10_inv08 = 1;
    128: op1_10_inv08 = 1;
    129: op1_10_inv08 = 1;
    131: op1_10_inv08 = 1;
    default: op1_10_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in09 = reg_0879;
    53: op1_10_in09 = reg_0117;
    86: op1_10_in09 = reg_0891;
    55: op1_10_in09 = reg_0407;
    73: op1_10_in09 = reg_0317;
    69: op1_10_in09 = reg_1314;
    49: op1_10_in09 = reg_0892;
    74: op1_10_in09 = reg_0165;
    54: op1_10_in09 = reg_0650;
    68: op1_10_in09 = imem03_in[7:4];
    75: op1_10_in09 = reg_1470;
    77: op1_10_in09 = reg_1470;
    50: op1_10_in09 = reg_0728;
    56: op1_10_in09 = reg_0750;
    71: op1_10_in09 = reg_0059;
    87: op1_10_in09 = reg_0421;
    76: op1_10_in09 = reg_0090;
    61: op1_10_in09 = reg_0725;
    57: op1_10_in09 = reg_0622;
    58: op1_10_in09 = reg_0605;
    78: op1_10_in09 = reg_0714;
    70: op1_10_in09 = reg_0790;
    79: op1_10_in09 = reg_1404;
    51: op1_10_in09 = reg_0703;
    104: op1_10_in09 = reg_0703;
    59: op1_10_in09 = reg_0020;
    60: op1_10_in09 = reg_0981;
    88: op1_10_in09 = reg_1339;
    46: op1_10_in09 = reg_0470;
    80: op1_10_in09 = reg_1417;
    95: op1_10_in09 = reg_1417;
    101: op1_10_in09 = reg_1417;
    81: op1_10_in09 = reg_0136;
    52: op1_10_in09 = reg_0774;
    63: op1_10_in09 = reg_0921;
    82: op1_10_in09 = reg_0419;
    89: op1_10_in09 = reg_0880;
    83: op1_10_in09 = reg_0155;
    64: op1_10_in09 = reg_1260;
    100: op1_10_in09 = reg_1260;
    84: op1_10_in09 = reg_0127;
    48: op1_10_in09 = reg_0827;
    85: op1_10_in09 = reg_0589;
    65: op1_10_in09 = reg_0779;
    90: op1_10_in09 = reg_1052;
    66: op1_10_in09 = reg_0093;
    37: op1_10_in09 = reg_0052;
    91: op1_10_in09 = reg_1208;
    67: op1_10_in09 = reg_0959;
    92: op1_10_in09 = reg_0462;
    93: op1_10_in09 = reg_0025;
    94: op1_10_in09 = reg_0845;
    96: op1_10_in09 = reg_0328;
    97: op1_10_in09 = reg_0112;
    98: op1_10_in09 = reg_0197;
    99: op1_10_in09 = reg_0592;
    102: op1_10_in09 = reg_0104;
    103: op1_10_in09 = reg_0799;
    108: op1_10_in09 = reg_0799;
    47: op1_10_in09 = reg_0367;
    105: op1_10_in09 = reg_0215;
    106: op1_10_in09 = reg_0433;
    44: op1_10_in09 = reg_0130;
    107: op1_10_in09 = reg_0684;
    109: op1_10_in09 = reg_1104;
    110: op1_10_in09 = reg_0839;
    111: op1_10_in09 = reg_0730;
    112: op1_10_in09 = reg_0927;
    113: op1_10_in09 = reg_1228;
    114: op1_10_in09 = reg_0627;
    115: op1_10_in09 = reg_1508;
    116: op1_10_in09 = reg_0897;
    117: op1_10_in09 = reg_0894;
    118: op1_10_in09 = reg_0734;
    119: op1_10_in09 = reg_0802;
    120: op1_10_in09 = reg_0472;
    121: op1_10_in09 = reg_0471;
    122: op1_10_in09 = reg_0233;
    123: op1_10_in09 = reg_0717;
    34: op1_10_in09 = reg_0484;
    124: op1_10_in09 = reg_0939;
    125: op1_10_in09 = reg_0071;
    126: op1_10_in09 = reg_0732;
    127: op1_10_in09 = reg_0973;
    128: op1_10_in09 = reg_1063;
    129: op1_10_in09 = reg_0262;
    130: op1_10_in09 = reg_0353;
    42: op1_10_in09 = reg_0451;
    131: op1_10_in09 = reg_0531;
    default: op1_10_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv09 = 1;
    86: op1_10_inv09 = 1;
    69: op1_10_inv09 = 1;
    75: op1_10_inv09 = 1;
    50: op1_10_inv09 = 1;
    71: op1_10_inv09 = 1;
    76: op1_10_inv09 = 1;
    57: op1_10_inv09 = 1;
    78: op1_10_inv09 = 1;
    59: op1_10_inv09 = 1;
    60: op1_10_inv09 = 1;
    81: op1_10_inv09 = 1;
    63: op1_10_inv09 = 1;
    82: op1_10_inv09 = 1;
    83: op1_10_inv09 = 1;
    84: op1_10_inv09 = 1;
    90: op1_10_inv09 = 1;
    92: op1_10_inv09 = 1;
    93: op1_10_inv09 = 1;
    94: op1_10_inv09 = 1;
    98: op1_10_inv09 = 1;
    103: op1_10_inv09 = 1;
    105: op1_10_inv09 = 1;
    44: op1_10_inv09 = 1;
    112: op1_10_inv09 = 1;
    113: op1_10_inv09 = 1;
    115: op1_10_inv09 = 1;
    117: op1_10_inv09 = 1;
    120: op1_10_inv09 = 1;
    121: op1_10_inv09 = 1;
    123: op1_10_inv09 = 1;
    125: op1_10_inv09 = 1;
    42: op1_10_inv09 = 1;
    131: op1_10_inv09 = 1;
    default: op1_10_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in10 = reg_0538;
    53: op1_10_in10 = reg_0129;
    86: op1_10_in10 = reg_0375;
    55: op1_10_in10 = reg_0598;
    73: op1_10_in10 = reg_0207;
    69: op1_10_in10 = reg_0190;
    49: op1_10_in10 = reg_0299;
    74: op1_10_in10 = reg_0371;
    54: op1_10_in10 = reg_0567;
    68: op1_10_in10 = imem03_in[15:12];
    75: op1_10_in10 = reg_1053;
    50: op1_10_in10 = reg_0386;
    56: op1_10_in10 = reg_0736;
    71: op1_10_in10 = reg_1254;
    87: op1_10_in10 = reg_0412;
    76: op1_10_in10 = reg_0873;
    61: op1_10_in10 = reg_0928;
    77: op1_10_in10 = reg_0928;
    57: op1_10_in10 = imem06_in[11:8];
    58: op1_10_in10 = reg_0607;
    78: op1_10_in10 = reg_0637;
    70: op1_10_in10 = reg_1280;
    79: op1_10_in10 = reg_0492;
    98: op1_10_in10 = reg_0492;
    51: op1_10_in10 = reg_0324;
    59: op1_10_in10 = imem05_in[15:12];
    60: op1_10_in10 = reg_0889;
    88: op1_10_in10 = reg_1338;
    46: op1_10_in10 = reg_0337;
    80: op1_10_in10 = reg_0155;
    81: op1_10_in10 = reg_1169;
    52: op1_10_in10 = reg_0663;
    63: op1_10_in10 = reg_0031;
    82: op1_10_in10 = reg_1202;
    89: op1_10_in10 = reg_0884;
    83: op1_10_in10 = reg_0524;
    64: op1_10_in10 = reg_0631;
    84: op1_10_in10 = reg_0382;
    48: op1_10_in10 = reg_0716;
    115: op1_10_in10 = reg_0716;
    85: op1_10_in10 = reg_0449;
    65: op1_10_in10 = reg_0661;
    90: op1_10_in10 = reg_0250;
    66: op1_10_in10 = reg_0899;
    37: op1_10_in10 = reg_0053;
    91: op1_10_in10 = reg_0108;
    67: op1_10_in10 = reg_1393;
    92: op1_10_in10 = reg_0574;
    93: op1_10_in10 = reg_0218;
    94: op1_10_in10 = reg_0608;
    95: op1_10_in10 = reg_0352;
    130: op1_10_in10 = reg_0352;
    96: op1_10_in10 = reg_0233;
    97: op1_10_in10 = reg_0106;
    99: op1_10_in10 = reg_0004;
    100: op1_10_in10 = reg_0054;
    101: op1_10_in10 = reg_1418;
    102: op1_10_in10 = reg_0291;
    103: op1_10_in10 = reg_0014;
    104: op1_10_in10 = reg_1350;
    47: op1_10_in10 = reg_0895;
    105: op1_10_in10 = reg_1170;
    106: op1_10_in10 = reg_0436;
    44: op1_10_in10 = reg_0243;
    107: op1_10_in10 = reg_0829;
    108: op1_10_in10 = reg_0151;
    109: op1_10_in10 = reg_0182;
    110: op1_10_in10 = reg_0390;
    111: op1_10_in10 = reg_0974;
    112: op1_10_in10 = reg_0189;
    113: op1_10_in10 = reg_0067;
    114: op1_10_in10 = reg_1447;
    116: op1_10_in10 = reg_0800;
    117: op1_10_in10 = reg_0219;
    118: op1_10_in10 = imem01_in[15:12];
    119: op1_10_in10 = reg_0903;
    120: op1_10_in10 = reg_0494;
    121: op1_10_in10 = reg_0454;
    122: op1_10_in10 = reg_0049;
    123: op1_10_in10 = reg_0374;
    124: op1_10_in10 = reg_0477;
    125: op1_10_in10 = reg_1321;
    126: op1_10_in10 = reg_0154;
    127: op1_10_in10 = reg_0628;
    128: op1_10_in10 = reg_0216;
    129: op1_10_in10 = reg_1340;
    42: op1_10_in10 = reg_0430;
    131: op1_10_in10 = reg_1083;
    default: op1_10_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv10 = 1;
    53: op1_10_inv10 = 1;
    55: op1_10_inv10 = 1;
    73: op1_10_inv10 = 1;
    69: op1_10_inv10 = 1;
    74: op1_10_inv10 = 1;
    68: op1_10_inv10 = 1;
    50: op1_10_inv10 = 1;
    71: op1_10_inv10 = 1;
    87: op1_10_inv10 = 1;
    57: op1_10_inv10 = 1;
    58: op1_10_inv10 = 1;
    60: op1_10_inv10 = 1;
    88: op1_10_inv10 = 1;
    46: op1_10_inv10 = 1;
    81: op1_10_inv10 = 1;
    52: op1_10_inv10 = 1;
    89: op1_10_inv10 = 1;
    83: op1_10_inv10 = 1;
    64: op1_10_inv10 = 1;
    48: op1_10_inv10 = 1;
    85: op1_10_inv10 = 1;
    65: op1_10_inv10 = 1;
    37: op1_10_inv10 = 1;
    67: op1_10_inv10 = 1;
    93: op1_10_inv10 = 1;
    95: op1_10_inv10 = 1;
    98: op1_10_inv10 = 1;
    99: op1_10_inv10 = 1;
    47: op1_10_inv10 = 1;
    105: op1_10_inv10 = 1;
    106: op1_10_inv10 = 1;
    107: op1_10_inv10 = 1;
    109: op1_10_inv10 = 1;
    112: op1_10_inv10 = 1;
    116: op1_10_inv10 = 1;
    117: op1_10_inv10 = 1;
    121: op1_10_inv10 = 1;
    122: op1_10_inv10 = 1;
    125: op1_10_inv10 = 1;
    127: op1_10_inv10 = 1;
    128: op1_10_inv10 = 1;
    130: op1_10_inv10 = 1;
    131: op1_10_inv10 = 1;
    default: op1_10_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in11 = reg_0541;
    53: op1_10_in11 = reg_0150;
    86: op1_10_in11 = reg_0377;
    55: op1_10_in11 = reg_0471;
    73: op1_10_in11 = reg_0038;
    69: op1_10_in11 = reg_0597;
    49: op1_10_in11 = imem07_in[11:8];
    74: op1_10_in11 = reg_0271;
    54: op1_10_in11 = reg_0418;
    68: op1_10_in11 = reg_1282;
    75: op1_10_in11 = reg_1052;
    50: op1_10_in11 = reg_0362;
    56: op1_10_in11 = reg_1059;
    71: op1_10_in11 = reg_1068;
    87: op1_10_in11 = reg_0537;
    76: op1_10_in11 = reg_1484;
    61: op1_10_in11 = reg_0387;
    57: op1_10_in11 = reg_0979;
    77: op1_10_in11 = reg_0927;
    58: op1_10_in11 = reg_0455;
    78: op1_10_in11 = reg_0373;
    70: op1_10_in11 = reg_0411;
    79: op1_10_in11 = reg_0118;
    51: op1_10_in11 = reg_0157;
    59: op1_10_in11 = reg_0832;
    60: op1_10_in11 = reg_0128;
    88: op1_10_in11 = reg_0531;
    46: op1_10_in11 = reg_0094;
    80: op1_10_in11 = reg_0476;
    81: op1_10_in11 = reg_0176;
    52: op1_10_in11 = reg_0739;
    63: op1_10_in11 = reg_0029;
    82: op1_10_in11 = reg_0270;
    89: op1_10_in11 = reg_0350;
    83: op1_10_in11 = reg_0353;
    64: op1_10_in11 = reg_0666;
    84: op1_10_in11 = reg_1032;
    48: op1_10_in11 = reg_0714;
    85: op1_10_in11 = reg_0861;
    65: op1_10_in11 = reg_0664;
    90: op1_10_in11 = reg_1229;
    66: op1_10_in11 = reg_0078;
    37: op1_10_in11 = reg_0084;
    91: op1_10_in11 = reg_0113;
    67: op1_10_in11 = reg_0431;
    92: op1_10_in11 = reg_1215;
    93: op1_10_in11 = reg_0288;
    94: op1_10_in11 = reg_0561;
    95: op1_10_in11 = reg_0201;
    96: op1_10_in11 = reg_0709;
    97: op1_10_in11 = reg_1140;
    98: op1_10_in11 = reg_1373;
    100: op1_10_in11 = reg_1451;
    106: op1_10_in11 = reg_1451;
    101: op1_10_in11 = reg_1405;
    102: op1_10_in11 = reg_0425;
    103: op1_10_in11 = imem06_in[3:0];
    104: op1_10_in11 = reg_1349;
    47: op1_10_in11 = reg_0243;
    105: op1_10_in11 = imem07_in[15:12];
    44: op1_10_in11 = reg_0240;
    107: op1_10_in11 = reg_0711;
    108: op1_10_in11 = reg_0729;
    109: op1_10_in11 = reg_1180;
    110: op1_10_in11 = reg_0973;
    111: op1_10_in11 = reg_0984;
    112: op1_10_in11 = reg_0389;
    113: op1_10_in11 = reg_0046;
    114: op1_10_in11 = reg_1301;
    115: op1_10_in11 = reg_0717;
    116: op1_10_in11 = reg_1006;
    117: op1_10_in11 = reg_1347;
    118: op1_10_in11 = reg_1152;
    119: op1_10_in11 = reg_1091;
    120: op1_10_in11 = reg_0054;
    121: op1_10_in11 = reg_0451;
    122: op1_10_in11 = reg_0185;
    123: op1_10_in11 = reg_0584;
    124: op1_10_in11 = reg_0303;
    125: op1_10_in11 = reg_0026;
    126: op1_10_in11 = reg_1001;
    127: op1_10_in11 = reg_0380;
    128: op1_10_in11 = reg_0312;
    129: op1_10_in11 = reg_1146;
    130: op1_10_in11 = reg_0722;
    42: op1_10_in11 = reg_0163;
    131: op1_10_in11 = reg_0421;
    default: op1_10_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv11 = 1;
    53: op1_10_inv11 = 1;
    86: op1_10_inv11 = 1;
    55: op1_10_inv11 = 1;
    69: op1_10_inv11 = 1;
    49: op1_10_inv11 = 1;
    54: op1_10_inv11 = 1;
    68: op1_10_inv11 = 1;
    87: op1_10_inv11 = 1;
    77: op1_10_inv11 = 1;
    80: op1_10_inv11 = 1;
    64: op1_10_inv11 = 1;
    84: op1_10_inv11 = 1;
    48: op1_10_inv11 = 1;
    66: op1_10_inv11 = 1;
    37: op1_10_inv11 = 1;
    91: op1_10_inv11 = 1;
    92: op1_10_inv11 = 1;
    93: op1_10_inv11 = 1;
    97: op1_10_inv11 = 1;
    101: op1_10_inv11 = 1;
    102: op1_10_inv11 = 1;
    103: op1_10_inv11 = 1;
    104: op1_10_inv11 = 1;
    106: op1_10_inv11 = 1;
    44: op1_10_inv11 = 1;
    107: op1_10_inv11 = 1;
    111: op1_10_inv11 = 1;
    112: op1_10_inv11 = 1;
    116: op1_10_inv11 = 1;
    117: op1_10_inv11 = 1;
    119: op1_10_inv11 = 1;
    122: op1_10_inv11 = 1;
    125: op1_10_inv11 = 1;
    127: op1_10_inv11 = 1;
    131: op1_10_inv11 = 1;
    default: op1_10_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in12 = reg_0167;
    53: op1_10_in12 = reg_0209;
    86: op1_10_in12 = reg_1314;
    55: op1_10_in12 = reg_0797;
    73: op1_10_in12 = reg_0466;
    69: op1_10_in12 = reg_1208;
    49: op1_10_in12 = reg_0777;
    74: op1_10_in12 = reg_0152;
    54: op1_10_in12 = reg_0302;
    68: op1_10_in12 = reg_0443;
    75: op1_10_in12 = reg_0523;
    50: op1_10_in12 = reg_0724;
    56: op1_10_in12 = reg_1164;
    59: op1_10_in12 = reg_1164;
    71: op1_10_in12 = reg_1069;
    87: op1_10_in12 = reg_0454;
    76: op1_10_in12 = reg_0275;
    61: op1_10_in12 = reg_0075;
    112: op1_10_in12 = reg_0075;
    57: op1_10_in12 = reg_0419;
    77: op1_10_in12 = reg_0883;
    58: op1_10_in12 = reg_0590;
    78: op1_10_in12 = reg_0979;
    70: op1_10_in12 = reg_0488;
    79: op1_10_in12 = reg_0240;
    51: op1_10_in12 = reg_0661;
    60: op1_10_in12 = reg_0126;
    88: op1_10_in12 = reg_0552;
    46: op1_10_in12 = reg_0211;
    80: op1_10_in12 = reg_0928;
    81: op1_10_in12 = reg_0392;
    52: op1_10_in12 = reg_0051;
    63: op1_10_in12 = reg_0437;
    82: op1_10_in12 = reg_0023;
    89: op1_10_in12 = reg_1149;
    83: op1_10_in12 = reg_0416;
    64: op1_10_in12 = reg_0934;
    84: op1_10_in12 = reg_0306;
    48: op1_10_in12 = reg_0669;
    85: op1_10_in12 = reg_0317;
    65: op1_10_in12 = reg_0286;
    90: op1_10_in12 = reg_1432;
    66: op1_10_in12 = reg_0278;
    37: op1_10_in12 = reg_0519;
    91: op1_10_in12 = reg_1009;
    67: op1_10_in12 = reg_0059;
    92: op1_10_in12 = reg_0414;
    131: op1_10_in12 = reg_0414;
    93: op1_10_in12 = reg_1282;
    94: op1_10_in12 = reg_1344;
    95: op1_10_in12 = reg_0189;
    96: op1_10_in12 = reg_0261;
    97: op1_10_in12 = reg_0381;
    127: op1_10_in12 = reg_0381;
    98: op1_10_in12 = reg_0274;
    100: op1_10_in12 = reg_0128;
    101: op1_10_in12 = reg_0352;
    102: op1_10_in12 = reg_0426;
    103: op1_10_in12 = reg_0784;
    104: op1_10_in12 = reg_0156;
    47: op1_10_in12 = reg_0118;
    105: op1_10_in12 = reg_0963;
    106: op1_10_in12 = reg_0629;
    44: op1_10_in12 = reg_0272;
    107: op1_10_in12 = imem02_in[3:0];
    108: op1_10_in12 = imem06_in[7:4];
    109: op1_10_in12 = reg_1402;
    110: op1_10_in12 = reg_0125;
    111: op1_10_in12 = reg_0751;
    113: op1_10_in12 = reg_0018;
    114: op1_10_in12 = reg_1231;
    115: op1_10_in12 = reg_0637;
    116: op1_10_in12 = reg_0009;
    117: op1_10_in12 = reg_0157;
    118: op1_10_in12 = reg_0930;
    119: op1_10_in12 = imem03_in[7:4];
    120: op1_10_in12 = reg_0972;
    121: op1_10_in12 = reg_1419;
    122: op1_10_in12 = reg_0706;
    123: op1_10_in12 = reg_0624;
    124: op1_10_in12 = reg_0318;
    125: op1_10_in12 = reg_0027;
    126: op1_10_in12 = reg_0783;
    128: op1_10_in12 = reg_0180;
    129: op1_10_in12 = imem04_in[3:0];
    130: op1_10_in12 = reg_0073;
    42: op1_10_in12 = reg_0402;
    default: op1_10_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_10_inv12 = 1;
    55: op1_10_inv12 = 1;
    73: op1_10_inv12 = 1;
    49: op1_10_inv12 = 1;
    74: op1_10_inv12 = 1;
    54: op1_10_inv12 = 1;
    68: op1_10_inv12 = 1;
    50: op1_10_inv12 = 1;
    56: op1_10_inv12 = 1;
    87: op1_10_inv12 = 1;
    76: op1_10_inv12 = 1;
    61: op1_10_inv12 = 1;
    78: op1_10_inv12 = 1;
    70: op1_10_inv12 = 1;
    51: op1_10_inv12 = 1;
    60: op1_10_inv12 = 1;
    46: op1_10_inv12 = 1;
    82: op1_10_inv12 = 1;
    89: op1_10_inv12 = 1;
    83: op1_10_inv12 = 1;
    84: op1_10_inv12 = 1;
    65: op1_10_inv12 = 1;
    91: op1_10_inv12 = 1;
    92: op1_10_inv12 = 1;
    93: op1_10_inv12 = 1;
    94: op1_10_inv12 = 1;
    95: op1_10_inv12 = 1;
    97: op1_10_inv12 = 1;
    98: op1_10_inv12 = 1;
    101: op1_10_inv12 = 1;
    47: op1_10_inv12 = 1;
    105: op1_10_inv12 = 1;
    106: op1_10_inv12 = 1;
    44: op1_10_inv12 = 1;
    110: op1_10_inv12 = 1;
    111: op1_10_inv12 = 1;
    112: op1_10_inv12 = 1;
    113: op1_10_inv12 = 1;
    116: op1_10_inv12 = 1;
    117: op1_10_inv12 = 1;
    118: op1_10_inv12 = 1;
    120: op1_10_inv12 = 1;
    121: op1_10_inv12 = 1;
    124: op1_10_inv12 = 1;
    126: op1_10_inv12 = 1;
    127: op1_10_inv12 = 1;
    129: op1_10_inv12 = 1;
    130: op1_10_inv12 = 1;
    42: op1_10_inv12 = 1;
    default: op1_10_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in13 = reg_0418;
    53: op1_10_in13 = reg_0035;
    86: op1_10_in13 = reg_0627;
    55: op1_10_in13 = reg_0369;
    73: op1_10_in13 = reg_1435;
    69: op1_10_in13 = reg_0885;
    49: op1_10_in13 = reg_0775;
    74: op1_10_in13 = imem07_in[3:0];
    54: op1_10_in13 = reg_0197;
    68: op1_10_in13 = reg_1384;
    75: op1_10_in13 = reg_0221;
    50: op1_10_in13 = reg_0871;
    56: op1_10_in13 = reg_0173;
    71: op1_10_in13 = reg_1071;
    87: op1_10_in13 = reg_0320;
    76: op1_10_in13 = reg_0601;
    61: op1_10_in13 = imem01_in[15:12];
    57: op1_10_in13 = reg_0289;
    77: op1_10_in13 = reg_1324;
    58: op1_10_in13 = reg_0530;
    78: op1_10_in13 = reg_1228;
    70: op1_10_in13 = reg_0181;
    79: op1_10_in13 = reg_0575;
    51: op1_10_in13 = reg_0664;
    59: op1_10_in13 = reg_1163;
    60: op1_10_in13 = reg_0111;
    88: op1_10_in13 = reg_0406;
    46: op1_10_in13 = reg_0064;
    80: op1_10_in13 = reg_0881;
    81: op1_10_in13 = reg_0066;
    63: op1_10_in13 = reg_0740;
    82: op1_10_in13 = reg_0215;
    89: op1_10_in13 = reg_0673;
    83: op1_10_in13 = reg_0410;
    64: op1_10_in13 = reg_0056;
    84: op1_10_in13 = reg_0294;
    48: op1_10_in13 = reg_0622;
    85: op1_10_in13 = reg_1468;
    65: op1_10_in13 = reg_0441;
    90: op1_10_in13 = reg_1417;
    66: op1_10_in13 = reg_0044;
    37: op1_10_in13 = reg_0521;
    91: op1_10_in13 = reg_0218;
    67: op1_10_in13 = reg_0917;
    92: op1_10_in13 = reg_0407;
    93: op1_10_in13 = reg_0237;
    94: op1_10_in13 = reg_0254;
    95: op1_10_in13 = reg_0416;
    101: op1_10_in13 = reg_0416;
    96: op1_10_in13 = reg_0557;
    97: op1_10_in13 = reg_0473;
    127: op1_10_in13 = reg_0473;
    98: op1_10_in13 = reg_0602;
    100: op1_10_in13 = reg_0127;
    102: op1_10_in13 = reg_0427;
    103: op1_10_in13 = reg_0795;
    108: op1_10_in13 = reg_0795;
    104: op1_10_in13 = reg_0924;
    47: op1_10_in13 = reg_0204;
    105: op1_10_in13 = reg_0394;
    106: op1_10_in13 = reg_0496;
    44: op1_10_in13 = reg_0205;
    107: op1_10_in13 = imem02_in[15:12];
    109: op1_10_in13 = reg_0090;
    110: op1_10_in13 = reg_0105;
    111: op1_10_in13 = reg_1323;
    112: op1_10_in13 = reg_0059;
    113: op1_10_in13 = reg_0017;
    114: op1_10_in13 = reg_1093;
    115: op1_10_in13 = reg_0585;
    116: op1_10_in13 = reg_0227;
    117: op1_10_in13 = reg_0139;
    118: op1_10_in13 = reg_0553;
    119: op1_10_in13 = reg_0190;
    120: op1_10_in13 = reg_0628;
    121: op1_10_in13 = reg_0582;
    122: op1_10_in13 = reg_0597;
    123: op1_10_in13 = reg_0529;
    124: op1_10_in13 = reg_0196;
    125: op1_10_in13 = reg_0267;
    126: op1_10_in13 = reg_0311;
    128: op1_10_in13 = reg_0789;
    129: op1_10_in13 = imem04_in[15:12];
    130: op1_10_in13 = reg_0072;
    42: op1_10_in13 = reg_0384;
    131: op1_10_in13 = reg_0412;
    default: op1_10_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv13 = 1;
    86: op1_10_inv13 = 1;
    74: op1_10_inv13 = 1;
    54: op1_10_inv13 = 1;
    68: op1_10_inv13 = 1;
    50: op1_10_inv13 = 1;
    56: op1_10_inv13 = 1;
    61: op1_10_inv13 = 1;
    57: op1_10_inv13 = 1;
    77: op1_10_inv13 = 1;
    58: op1_10_inv13 = 1;
    51: op1_10_inv13 = 1;
    59: op1_10_inv13 = 1;
    89: op1_10_inv13 = 1;
    83: op1_10_inv13 = 1;
    64: op1_10_inv13 = 1;
    84: op1_10_inv13 = 1;
    90: op1_10_inv13 = 1;
    92: op1_10_inv13 = 1;
    93: op1_10_inv13 = 1;
    98: op1_10_inv13 = 1;
    100: op1_10_inv13 = 1;
    102: op1_10_inv13 = 1;
    104: op1_10_inv13 = 1;
    106: op1_10_inv13 = 1;
    108: op1_10_inv13 = 1;
    110: op1_10_inv13 = 1;
    111: op1_10_inv13 = 1;
    113: op1_10_inv13 = 1;
    114: op1_10_inv13 = 1;
    117: op1_10_inv13 = 1;
    120: op1_10_inv13 = 1;
    121: op1_10_inv13 = 1;
    122: op1_10_inv13 = 1;
    123: op1_10_inv13 = 1;
    124: op1_10_inv13 = 1;
    125: op1_10_inv13 = 1;
    126: op1_10_inv13 = 1;
    127: op1_10_inv13 = 1;
    128: op1_10_inv13 = 1;
    42: op1_10_inv13 = 1;
    default: op1_10_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in14 = reg_0872;
    53: op1_10_in14 = reg_0331;
    86: op1_10_in14 = reg_0048;
    55: op1_10_in14 = reg_0488;
    73: op1_10_in14 = reg_0905;
    69: op1_10_in14 = reg_0880;
    49: op1_10_in14 = reg_0029;
    74: op1_10_in14 = reg_0391;
    54: op1_10_in14 = reg_0196;
    76: op1_10_in14 = reg_0196;
    68: op1_10_in14 = reg_1372;
    75: op1_10_in14 = reg_1201;
    50: op1_10_in14 = reg_0013;
    56: op1_10_in14 = reg_0648;
    71: op1_10_in14 = reg_0553;
    87: op1_10_in14 = reg_0369;
    61: op1_10_in14 = reg_1254;
    125: op1_10_in14 = reg_1254;
    57: op1_10_in14 = reg_0023;
    77: op1_10_in14 = reg_1322;
    58: op1_10_in14 = reg_0533;
    78: op1_10_in14 = reg_1225;
    70: op1_10_in14 = reg_1369;
    79: op1_10_in14 = reg_1348;
    51: op1_10_in14 = reg_0366;
    59: op1_10_in14 = reg_0173;
    60: op1_10_in14 = reg_0112;
    88: op1_10_in14 = reg_0599;
    46: op1_10_in14 = reg_0021;
    80: op1_10_in14 = reg_0353;
    81: op1_10_in14 = imem05_in[3:0];
    63: op1_10_in14 = reg_0623;
    82: op1_10_in14 = reg_0213;
    89: op1_10_in14 = reg_0348;
    83: op1_10_in14 = reg_0075;
    64: op1_10_in14 = reg_0390;
    84: op1_10_in14 = reg_0311;
    48: op1_10_in14 = reg_0624;
    85: op1_10_in14 = reg_0396;
    65: op1_10_in14 = reg_0408;
    90: op1_10_in14 = reg_0524;
    66: op1_10_in14 = reg_0012;
    91: op1_10_in14 = reg_0291;
    67: op1_10_in14 = reg_0822;
    92: op1_10_in14 = reg_0969;
    93: op1_10_in14 = reg_0696;
    94: op1_10_in14 = reg_0712;
    95: op1_10_in14 = reg_0388;
    96: op1_10_in14 = reg_0198;
    97: op1_10_in14 = reg_0327;
    98: op1_10_in14 = reg_0344;
    100: op1_10_in14 = reg_0111;
    101: op1_10_in14 = reg_0409;
    102: op1_10_in14 = imem04_in[7:4];
    103: op1_10_in14 = reg_0397;
    104: op1_10_in14 = reg_0923;
    47: op1_10_in14 = reg_0014;
    105: op1_10_in14 = reg_1060;
    106: op1_10_in14 = reg_0878;
    44: op1_10_in14 = reg_0038;
    107: op1_10_in14 = reg_0024;
    108: op1_10_in14 = reg_0316;
    109: op1_10_in14 = reg_0828;
    124: op1_10_in14 = reg_0828;
    110: op1_10_in14 = reg_0496;
    111: op1_10_in14 = reg_1501;
    112: op1_10_in14 = reg_1321;
    113: op1_10_in14 = reg_1170;
    114: op1_10_in14 = reg_1092;
    115: op1_10_in14 = reg_0571;
    116: op1_10_in14 = reg_0190;
    117: op1_10_in14 = reg_0030;
    118: op1_10_in14 = reg_0550;
    119: op1_10_in14 = reg_0989;
    120: op1_10_in14 = reg_0381;
    121: op1_10_in14 = reg_0062;
    122: op1_10_in14 = reg_0220;
    123: op1_10_in14 = reg_0527;
    126: op1_10_in14 = reg_0312;
    127: op1_10_in14 = reg_0253;
    128: op1_10_in14 = reg_0964;
    129: op1_10_in14 = reg_0064;
    130: op1_10_in14 = reg_0057;
    42: op1_10_in14 = reg_0385;
    131: op1_10_in14 = reg_1065;
    default: op1_10_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_10_inv14 = 1;
    73: op1_10_inv14 = 1;
    49: op1_10_inv14 = 1;
    74: op1_10_inv14 = 1;
    68: op1_10_inv14 = 1;
    56: op1_10_inv14 = 1;
    71: op1_10_inv14 = 1;
    79: op1_10_inv14 = 1;
    60: op1_10_inv14 = 1;
    46: op1_10_inv14 = 1;
    80: op1_10_inv14 = 1;
    81: op1_10_inv14 = 1;
    89: op1_10_inv14 = 1;
    64: op1_10_inv14 = 1;
    85: op1_10_inv14 = 1;
    90: op1_10_inv14 = 1;
    66: op1_10_inv14 = 1;
    92: op1_10_inv14 = 1;
    93: op1_10_inv14 = 1;
    95: op1_10_inv14 = 1;
    97: op1_10_inv14 = 1;
    98: op1_10_inv14 = 1;
    100: op1_10_inv14 = 1;
    102: op1_10_inv14 = 1;
    104: op1_10_inv14 = 1;
    47: op1_10_inv14 = 1;
    106: op1_10_inv14 = 1;
    110: op1_10_inv14 = 1;
    114: op1_10_inv14 = 1;
    115: op1_10_inv14 = 1;
    116: op1_10_inv14 = 1;
    118: op1_10_inv14 = 1;
    119: op1_10_inv14 = 1;
    121: op1_10_inv14 = 1;
    123: op1_10_inv14 = 1;
    128: op1_10_inv14 = 1;
    130: op1_10_inv14 = 1;
    default: op1_10_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in15 = reg_0303;
    53: op1_10_in15 = reg_0748;
    86: op1_10_in15 = reg_1226;
    55: op1_10_in15 = reg_0487;
    73: op1_10_in15 = reg_0133;
    69: op1_10_in15 = reg_0507;
    49: op1_10_in15 = reg_0740;
    74: op1_10_in15 = reg_1440;
    54: op1_10_in15 = reg_0243;
    68: op1_10_in15 = reg_1369;
    75: op1_10_in15 = reg_0459;
    50: op1_10_in15 = reg_0486;
    56: op1_10_in15 = reg_0650;
    71: op1_10_in15 = reg_0547;
    87: op1_10_in15 = reg_0582;
    76: op1_10_in15 = reg_0631;
    100: op1_10_in15 = reg_0631;
    61: op1_10_in15 = reg_1071;
    57: op1_10_in15 = reg_0152;
    77: op1_10_in15 = reg_1034;
    58: op1_10_in15 = imem02_in[7:4];
    78: op1_10_in15 = reg_0419;
    70: op1_10_in15 = reg_0577;
    79: op1_10_in15 = reg_0014;
    109: op1_10_in15 = reg_0014;
    124: op1_10_in15 = reg_0014;
    51: op1_10_in15 = reg_0592;
    59: op1_10_in15 = reg_0646;
    60: op1_10_in15 = reg_0138;
    88: op1_10_in15 = reg_1040;
    92: op1_10_in15 = reg_1040;
    46: op1_10_in15 = reg_0020;
    80: op1_10_in15 = reg_0189;
    81: op1_10_in15 = reg_0167;
    63: op1_10_in15 = reg_0618;
    65: op1_10_in15 = reg_0618;
    82: op1_10_in15 = reg_0017;
    89: op1_10_in15 = reg_0425;
    83: op1_10_in15 = reg_0060;
    64: op1_10_in15 = reg_0306;
    84: op1_10_in15 = reg_0313;
    48: op1_10_in15 = reg_0526;
    85: op1_10_in15 = reg_0466;
    90: op1_10_in15 = reg_0881;
    66: op1_10_in15 = reg_0010;
    91: op1_10_in15 = reg_0443;
    67: op1_10_in15 = reg_0335;
    93: op1_10_in15 = reg_1372;
    94: op1_10_in15 = reg_0532;
    95: op1_10_in15 = reg_0026;
    96: op1_10_in15 = reg_0312;
    97: op1_10_in15 = reg_1078;
    98: op1_10_in15 = reg_0589;
    101: op1_10_in15 = reg_0134;
    102: op1_10_in15 = imem04_in[11:8];
    103: op1_10_in15 = reg_1334;
    104: op1_10_in15 = reg_0663;
    47: op1_10_in15 = reg_0754;
    44: op1_10_in15 = reg_0754;
    105: op1_10_in15 = reg_0892;
    106: op1_10_in15 = reg_0307;
    107: op1_10_in15 = reg_0759;
    108: op1_10_in15 = reg_0751;
    110: op1_10_in15 = reg_1140;
    111: op1_10_in15 = reg_0717;
    112: op1_10_in15 = reg_1322;
    113: op1_10_in15 = reg_1096;
    114: op1_10_in15 = reg_1208;
    115: op1_10_in15 = reg_0522;
    116: op1_10_in15 = reg_0179;
    117: op1_10_in15 = reg_0664;
    118: op1_10_in15 = reg_0548;
    119: op1_10_in15 = reg_1448;
    120: op1_10_in15 = reg_0253;
    121: op1_10_in15 = reg_1340;
    122: op1_10_in15 = reg_0177;
    123: op1_10_in15 = reg_0308;
    125: op1_10_in15 = reg_0902;
    126: op1_10_in15 = reg_1300;
    127: op1_10_in15 = reg_0007;
    128: op1_10_in15 = reg_1314;
    129: op1_10_in15 = reg_1502;
    130: op1_10_in15 = reg_0267;
    42: op1_10_in15 = reg_0362;
    131: op1_10_in15 = reg_1419;
    default: op1_10_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_10_inv15 = 1;
    55: op1_10_inv15 = 1;
    73: op1_10_inv15 = 1;
    69: op1_10_inv15 = 1;
    49: op1_10_inv15 = 1;
    74: op1_10_inv15 = 1;
    54: op1_10_inv15 = 1;
    71: op1_10_inv15 = 1;
    76: op1_10_inv15 = 1;
    57: op1_10_inv15 = 1;
    58: op1_10_inv15 = 1;
    78: op1_10_inv15 = 1;
    70: op1_10_inv15 = 1;
    79: op1_10_inv15 = 1;
    59: op1_10_inv15 = 1;
    46: op1_10_inv15 = 1;
    80: op1_10_inv15 = 1;
    81: op1_10_inv15 = 1;
    83: op1_10_inv15 = 1;
    64: op1_10_inv15 = 1;
    48: op1_10_inv15 = 1;
    85: op1_10_inv15 = 1;
    91: op1_10_inv15 = 1;
    67: op1_10_inv15 = 1;
    93: op1_10_inv15 = 1;
    94: op1_10_inv15 = 1;
    95: op1_10_inv15 = 1;
    97: op1_10_inv15 = 1;
    98: op1_10_inv15 = 1;
    100: op1_10_inv15 = 1;
    101: op1_10_inv15 = 1;
    102: op1_10_inv15 = 1;
    103: op1_10_inv15 = 1;
    104: op1_10_inv15 = 1;
    47: op1_10_inv15 = 1;
    106: op1_10_inv15 = 1;
    107: op1_10_inv15 = 1;
    110: op1_10_inv15 = 1;
    111: op1_10_inv15 = 1;
    113: op1_10_inv15 = 1;
    114: op1_10_inv15 = 1;
    115: op1_10_inv15 = 1;
    116: op1_10_inv15 = 1;
    117: op1_10_inv15 = 1;
    118: op1_10_inv15 = 1;
    119: op1_10_inv15 = 1;
    120: op1_10_inv15 = 1;
    123: op1_10_inv15 = 1;
    124: op1_10_inv15 = 1;
    125: op1_10_inv15 = 1;
    129: op1_10_inv15 = 1;
    130: op1_10_inv15 = 1;
    42: op1_10_inv15 = 1;
    default: op1_10_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in16 = reg_0302;
    53: op1_10_in16 = reg_0750;
    86: op1_10_in16 = reg_1199;
    55: op1_10_in16 = reg_0836;
    73: op1_10_in16 = imem06_in[3:0];
    69: op1_10_in16 = reg_0479;
    49: op1_10_in16 = reg_0408;
    74: op1_10_in16 = reg_1416;
    54: op1_10_in16 = reg_0864;
    68: op1_10_in16 = reg_1200;
    75: op1_10_in16 = reg_1405;
    50: op1_10_in16 = imem02_in[7:4];
    56: op1_10_in16 = reg_0334;
    71: op1_10_in16 = reg_0549;
    87: op1_10_in16 = reg_0862;
    76: op1_10_in16 = reg_0449;
    61: op1_10_in16 = reg_0547;
    125: op1_10_in16 = reg_0547;
    57: op1_10_in16 = reg_0215;
    77: op1_10_in16 = reg_1256;
    58: op1_10_in16 = reg_0473;
    106: op1_10_in16 = reg_0473;
    78: op1_10_in16 = reg_1179;
    70: op1_10_in16 = reg_1083;
    79: op1_10_in16 = imem06_in[15:12];
    109: op1_10_in16 = imem06_in[15:12];
    51: op1_10_in16 = reg_0004;
    59: op1_10_in16 = reg_0650;
    60: op1_10_in16 = reg_0007;
    88: op1_10_in16 = reg_1077;
    46: op1_10_in16 = reg_0793;
    80: op1_10_in16 = reg_0428;
    81: op1_10_in16 = reg_0630;
    63: op1_10_in16 = reg_0321;
    82: op1_10_in16 = reg_0034;
    89: op1_10_in16 = reg_1312;
    83: op1_10_in16 = reg_0072;
    64: op1_10_in16 = reg_0008;
    84: op1_10_in16 = reg_1495;
    48: op1_10_in16 = reg_0529;
    85: op1_10_in16 = reg_1437;
    65: op1_10_in16 = reg_0591;
    90: op1_10_in16 = reg_0887;
    66: op1_10_in16 = reg_0486;
    91: op1_10_in16 = reg_0411;
    67: op1_10_in16 = reg_1254;
    92: op1_10_in16 = reg_0199;
    93: op1_10_in16 = reg_0181;
    94: op1_10_in16 = reg_0432;
    95: op1_10_in16 = reg_0005;
    96: op1_10_in16 = reg_1313;
    97: op1_10_in16 = imem03_in[7:4];
    98: op1_10_in16 = reg_0828;
    100: op1_10_in16 = reg_1392;
    101: op1_10_in16 = reg_0387;
    102: op1_10_in16 = reg_0577;
    103: op1_10_in16 = reg_1209;
    104: op1_10_in16 = reg_0664;
    47: op1_10_in16 = reg_0751;
    105: op1_10_in16 = reg_1347;
    44: op1_10_in16 = reg_0753;
    107: op1_10_in16 = reg_0377;
    108: op1_10_in16 = reg_1505;
    110: op1_10_in16 = reg_0876;
    111: op1_10_in16 = reg_0398;
    112: op1_10_in16 = reg_0027;
    113: op1_10_in16 = reg_1060;
    114: op1_10_in16 = reg_0882;
    115: op1_10_in16 = reg_0132;
    116: op1_10_in16 = reg_0311;
    117: op1_10_in16 = reg_0284;
    118: op1_10_in16 = reg_0787;
    119: op1_10_in16 = reg_0049;
    120: op1_10_in16 = reg_0848;
    121: op1_10_in16 = reg_1107;
    122: op1_10_in16 = reg_1001;
    123: op1_10_in16 = reg_0119;
    124: op1_10_in16 = reg_0908;
    126: op1_10_in16 = reg_0558;
    127: op1_10_in16 = reg_0903;
    128: op1_10_in16 = reg_0756;
    129: op1_10_in16 = reg_0633;
    130: op1_10_in16 = reg_0635;
    42: op1_10_in16 = reg_0365;
    131: op1_10_in16 = reg_1144;
    default: op1_10_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv16 = 1;
    69: op1_10_inv16 = 1;
    74: op1_10_inv16 = 1;
    68: op1_10_inv16 = 1;
    75: op1_10_inv16 = 1;
    76: op1_10_inv16 = 1;
    61: op1_10_inv16 = 1;
    57: op1_10_inv16 = 1;
    58: op1_10_inv16 = 1;
    78: op1_10_inv16 = 1;
    70: op1_10_inv16 = 1;
    79: op1_10_inv16 = 1;
    51: op1_10_inv16 = 1;
    60: op1_10_inv16 = 1;
    88: op1_10_inv16 = 1;
    46: op1_10_inv16 = 1;
    80: op1_10_inv16 = 1;
    83: op1_10_inv16 = 1;
    48: op1_10_inv16 = 1;
    65: op1_10_inv16 = 1;
    93: op1_10_inv16 = 1;
    94: op1_10_inv16 = 1;
    96: op1_10_inv16 = 1;
    98: op1_10_inv16 = 1;
    102: op1_10_inv16 = 1;
    103: op1_10_inv16 = 1;
    104: op1_10_inv16 = 1;
    108: op1_10_inv16 = 1;
    112: op1_10_inv16 = 1;
    113: op1_10_inv16 = 1;
    114: op1_10_inv16 = 1;
    115: op1_10_inv16 = 1;
    116: op1_10_inv16 = 1;
    119: op1_10_inv16 = 1;
    121: op1_10_inv16 = 1;
    124: op1_10_inv16 = 1;
    126: op1_10_inv16 = 1;
    127: op1_10_inv16 = 1;
    129: op1_10_inv16 = 1;
    130: op1_10_inv16 = 1;
    default: op1_10_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in17 = reg_0301;
    53: op1_10_in17 = reg_0733;
    86: op1_10_in17 = reg_0178;
    55: op1_10_in17 = reg_0794;
    73: op1_10_in17 = reg_0718;
    69: op1_10_in17 = reg_0478;
    49: op1_10_in17 = reg_0621;
    74: op1_10_in17 = reg_0667;
    54: op1_10_in17 = reg_0207;
    68: op1_10_in17 = reg_1082;
    70: op1_10_in17 = reg_1082;
    93: op1_10_in17 = reg_1082;
    75: op1_10_in17 = reg_0881;
    50: op1_10_in17 = reg_1029;
    56: op1_10_in17 = reg_0540;
    71: op1_10_in17 = reg_0463;
    87: op1_10_in17 = reg_1237;
    76: op1_10_in17 = reg_0861;
    61: op1_10_in17 = reg_0242;
    57: op1_10_in17 = reg_0213;
    77: op1_10_in17 = reg_1513;
    58: op1_10_in17 = reg_0475;
    78: op1_10_in17 = reg_0269;
    109: op1_10_in17 = reg_0269;
    79: op1_10_in17 = reg_0195;
    44: op1_10_in17 = reg_0195;
    51: op1_10_in17 = reg_0123;
    59: op1_10_in17 = reg_0333;
    60: op1_10_in17 = reg_0327;
    88: op1_10_in17 = reg_1065;
    46: op1_10_in17 = reg_0748;
    80: op1_10_in17 = reg_0134;
    81: op1_10_in17 = reg_1181;
    63: op1_10_in17 = reg_0086;
    82: op1_10_in17 = reg_1183;
    89: op1_10_in17 = reg_0493;
    83: op1_10_in17 = reg_1324;
    64: op1_10_in17 = reg_0830;
    84: op1_10_in17 = imem03_in[3:0];
    48: op1_10_in17 = reg_0527;
    85: op1_10_in17 = reg_0825;
    65: op1_10_in17 = reg_0103;
    90: op1_10_in17 = reg_1321;
    66: op1_10_in17 = reg_0606;
    91: op1_10_in17 = reg_1144;
    67: op1_10_in17 = reg_1071;
    92: op1_10_in17 = reg_1077;
    94: op1_10_in17 = reg_0433;
    95: op1_10_in17 = reg_0734;
    96: op1_10_in17 = reg_1301;
    97: op1_10_in17 = reg_0840;
    98: op1_10_in17 = reg_0039;
    100: op1_10_in17 = reg_1078;
    101: op1_10_in17 = reg_0071;
    102: op1_10_in17 = reg_1383;
    103: op1_10_in17 = reg_0316;
    104: op1_10_in17 = reg_0618;
    47: op1_10_in17 = reg_0193;
    105: op1_10_in17 = reg_0157;
    106: op1_10_in17 = reg_0306;
    107: op1_10_in17 = reg_0750;
    108: op1_10_in17 = reg_0780;
    110: op1_10_in17 = reg_0381;
    111: op1_10_in17 = reg_0374;
    112: op1_10_in17 = reg_0917;
    113: op1_10_in17 = reg_0135;
    114: op1_10_in17 = reg_0458;
    115: op1_10_in17 = reg_0296;
    116: op1_10_in17 = reg_1184;
    117: op1_10_in17 = reg_0415;
    118: op1_10_in17 = reg_0222;
    119: op1_10_in17 = reg_0444;
    120: op1_10_in17 = reg_0217;
    121: op1_10_in17 = reg_0063;
    122: op1_10_in17 = reg_0823;
    123: op1_10_in17 = reg_0371;
    124: op1_10_in17 = reg_1064;
    125: op1_10_in17 = reg_0550;
    126: op1_10_in17 = reg_1199;
    127: op1_10_in17 = reg_0848;
    128: op1_10_in17 = reg_1300;
    129: op1_10_in17 = reg_0019;
    130: op1_10_in17 = imem01_in[3:0];
    42: op1_10_in17 = reg_0320;
    131: op1_10_in17 = reg_0065;
    default: op1_10_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv17 = 1;
    86: op1_10_inv17 = 1;
    55: op1_10_inv17 = 1;
    73: op1_10_inv17 = 1;
    69: op1_10_inv17 = 1;
    74: op1_10_inv17 = 1;
    54: op1_10_inv17 = 1;
    68: op1_10_inv17 = 1;
    56: op1_10_inv17 = 1;
    87: op1_10_inv17 = 1;
    57: op1_10_inv17 = 1;
    77: op1_10_inv17 = 1;
    58: op1_10_inv17 = 1;
    70: op1_10_inv17 = 1;
    79: op1_10_inv17 = 1;
    51: op1_10_inv17 = 1;
    60: op1_10_inv17 = 1;
    88: op1_10_inv17 = 1;
    81: op1_10_inv17 = 1;
    82: op1_10_inv17 = 1;
    48: op1_10_inv17 = 1;
    90: op1_10_inv17 = 1;
    91: op1_10_inv17 = 1;
    94: op1_10_inv17 = 1;
    97: op1_10_inv17 = 1;
    98: op1_10_inv17 = 1;
    100: op1_10_inv17 = 1;
    101: op1_10_inv17 = 1;
    104: op1_10_inv17 = 1;
    105: op1_10_inv17 = 1;
    106: op1_10_inv17 = 1;
    107: op1_10_inv17 = 1;
    108: op1_10_inv17 = 1;
    112: op1_10_inv17 = 1;
    113: op1_10_inv17 = 1;
    114: op1_10_inv17 = 1;
    115: op1_10_inv17 = 1;
    116: op1_10_inv17 = 1;
    119: op1_10_inv17 = 1;
    120: op1_10_inv17 = 1;
    123: op1_10_inv17 = 1;
    125: op1_10_inv17 = 1;
    127: op1_10_inv17 = 1;
    129: op1_10_inv17 = 1;
    default: op1_10_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in18 = imem05_in[3:0];
    53: op1_10_in18 = reg_0832;
    86: op1_10_in18 = reg_0108;
    55: op1_10_in18 = reg_0578;
    73: op1_10_in18 = reg_0637;
    69: op1_10_in18 = reg_1282;
    49: op1_10_in18 = reg_0137;
    74: op1_10_in18 = reg_0170;
    54: op1_10_in18 = reg_0037;
    68: op1_10_in18 = reg_0406;
    75: op1_10_in18 = reg_0883;
    50: op1_10_in18 = reg_0563;
    56: op1_10_in18 = reg_0937;
    71: op1_10_in18 = imem01_in[7:4];
    87: op1_10_in18 = reg_0117;
    76: op1_10_in18 = reg_0039;
    61: op1_10_in18 = reg_1152;
    57: op1_10_in18 = reg_0490;
    77: op1_10_in18 = reg_0047;
    58: op1_10_in18 = reg_0472;
    78: op1_10_in18 = reg_0706;
    70: op1_10_in18 = reg_0421;
    79: op1_10_in18 = reg_1064;
    59: op1_10_in18 = reg_0539;
    60: op1_10_in18 = reg_0068;
    88: op1_10_in18 = reg_0319;
    46: op1_10_in18 = reg_0733;
    80: op1_10_in18 = reg_0072;
    81: op1_10_in18 = reg_0697;
    63: op1_10_in18 = reg_1182;
    82: op1_10_in18 = reg_0922;
    89: op1_10_in18 = reg_0264;
    83: op1_10_in18 = reg_0917;
    64: op1_10_in18 = reg_0069;
    84: op1_10_in18 = imem03_in[15:12];
    48: op1_10_in18 = reg_0458;
    85: op1_10_in18 = reg_0908;
    65: op1_10_in18 = reg_0100;
    90: op1_10_in18 = reg_0026;
    66: op1_10_in18 = reg_0532;
    91: op1_10_in18 = reg_0062;
    67: op1_10_in18 = reg_1032;
    92: op1_10_in18 = reg_0304;
    93: op1_10_in18 = reg_1147;
    94: op1_10_in18 = reg_0970;
    95: op1_10_in18 = reg_1031;
    96: op1_10_in18 = reg_1093;
    97: op1_10_in18 = reg_0559;
    98: op1_10_in18 = reg_0014;
    100: op1_10_in18 = reg_0227;
    101: op1_10_in18 = reg_0059;
    102: op1_10_in18 = reg_0263;
    103: op1_10_in18 = reg_1420;
    104: op1_10_in18 = reg_0591;
    47: op1_10_in18 = reg_0192;
    124: op1_10_in18 = reg_0192;
    105: op1_10_in18 = reg_0489;
    106: op1_10_in18 = reg_0897;
    44: op1_10_in18 = imem06_in[15:12];
    107: op1_10_in18 = reg_0261;
    108: op1_10_in18 = reg_0586;
    109: op1_10_in18 = reg_0795;
    110: op1_10_in18 = reg_0307;
    111: op1_10_in18 = reg_0529;
    112: op1_10_in18 = reg_1253;
    113: op1_10_in18 = reg_0310;
    114: op1_10_in18 = reg_0707;
    115: op1_10_in18 = reg_0295;
    116: op1_10_in18 = reg_0964;
    117: op1_10_in18 = reg_0085;
    118: op1_10_in18 = reg_0609;
    119: op1_10_in18 = reg_0709;
    120: op1_10_in18 = reg_0006;
    121: op1_10_in18 = reg_0065;
    122: op1_10_in18 = reg_0312;
    123: op1_10_in18 = reg_0977;
    125: op1_10_in18 = reg_0787;
    126: op1_10_in18 = reg_0178;
    127: op1_10_in18 = reg_0024;
    128: op1_10_in18 = reg_0290;
    129: op1_10_in18 = imem05_in[15:12];
    130: op1_10_in18 = reg_0078;
    42: op1_10_in18 = reg_0091;
    131: op1_10_in18 = reg_0095;
    default: op1_10_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    49: op1_10_inv18 = 1;
    68: op1_10_inv18 = 1;
    75: op1_10_inv18 = 1;
    50: op1_10_inv18 = 1;
    71: op1_10_inv18 = 1;
    87: op1_10_inv18 = 1;
    76: op1_10_inv18 = 1;
    61: op1_10_inv18 = 1;
    70: op1_10_inv18 = 1;
    60: op1_10_inv18 = 1;
    46: op1_10_inv18 = 1;
    80: op1_10_inv18 = 1;
    82: op1_10_inv18 = 1;
    83: op1_10_inv18 = 1;
    64: op1_10_inv18 = 1;
    84: op1_10_inv18 = 1;
    65: op1_10_inv18 = 1;
    90: op1_10_inv18 = 1;
    92: op1_10_inv18 = 1;
    93: op1_10_inv18 = 1;
    94: op1_10_inv18 = 1;
    96: op1_10_inv18 = 1;
    98: op1_10_inv18 = 1;
    104: op1_10_inv18 = 1;
    47: op1_10_inv18 = 1;
    105: op1_10_inv18 = 1;
    106: op1_10_inv18 = 1;
    44: op1_10_inv18 = 1;
    109: op1_10_inv18 = 1;
    110: op1_10_inv18 = 1;
    112: op1_10_inv18 = 1;
    120: op1_10_inv18 = 1;
    123: op1_10_inv18 = 1;
    124: op1_10_inv18 = 1;
    126: op1_10_inv18 = 1;
    129: op1_10_inv18 = 1;
    130: op1_10_inv18 = 1;
    42: op1_10_inv18 = 1;
    default: op1_10_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in19 = reg_0864;
    53: op1_10_in19 = reg_0700;
    86: op1_10_in19 = reg_0107;
    55: op1_10_in19 = reg_0176;
    73: op1_10_in19 = reg_0979;
    69: op1_10_in19 = reg_0443;
    49: op1_10_in19 = reg_0004;
    74: op1_10_in19 = reg_1345;
    54: op1_10_in19 = reg_0751;
    68: op1_10_in19 = reg_0598;
    75: op1_10_in19 = reg_0416;
    50: op1_10_in19 = reg_0533;
    56: op1_10_in19 = reg_0070;
    116: op1_10_in19 = reg_0070;
    71: op1_10_in19 = imem01_in[15:12];
    87: op1_10_in19 = reg_0536;
    76: op1_10_in19 = reg_0466;
    61: op1_10_in19 = reg_0468;
    57: op1_10_in19 = reg_0821;
    77: op1_10_in19 = reg_0572;
    58: op1_10_in19 = reg_0433;
    78: op1_10_in19 = reg_0461;
    70: op1_10_in19 = reg_0414;
    79: op1_10_in19 = reg_0264;
    59: op1_10_in19 = reg_0938;
    60: op1_10_in19 = reg_0325;
    88: op1_10_in19 = reg_0487;
    46: op1_10_in19 = reg_0828;
    80: op1_10_in19 = reg_0057;
    81: op1_10_in19 = reg_1402;
    82: op1_10_in19 = reg_0894;
    89: op1_10_in19 = reg_1339;
    83: op1_10_in19 = reg_1100;
    64: op1_10_in19 = reg_0198;
    84: op1_10_in19 = reg_0444;
    48: op1_10_in19 = reg_0023;
    85: op1_10_in19 = reg_1209;
    124: op1_10_in19 = reg_1209;
    65: op1_10_in19 = reg_0086;
    117: op1_10_in19 = reg_0086;
    90: op1_10_in19 = reg_0747;
    66: op1_10_in19 = reg_0562;
    91: op1_10_in19 = reg_1372;
    67: op1_10_in19 = reg_0634;
    92: op1_10_in19 = reg_0319;
    93: op1_10_in19 = reg_0407;
    94: op1_10_in19 = reg_1451;
    95: op1_10_in19 = reg_1256;
    96: op1_10_in19 = reg_1092;
    97: op1_10_in19 = reg_0710;
    98: op1_10_in19 = reg_0265;
    100: op1_10_in19 = reg_0233;
    101: op1_10_in19 = reg_0058;
    102: op1_10_in19 = reg_0535;
    103: op1_10_in19 = reg_0984;
    104: op1_10_in19 = reg_0137;
    47: op1_10_in19 = imem06_in[11:8];
    105: op1_10_in19 = reg_0465;
    106: op1_10_in19 = reg_1098;
    44: op1_10_in19 = reg_0826;
    107: op1_10_in19 = reg_1425;
    108: op1_10_in19 = reg_0584;
    109: op1_10_in19 = reg_0906;
    110: op1_10_in19 = reg_0829;
    111: op1_10_in19 = reg_0527;
    112: op1_10_in19 = imem01_in[3:0];
    42: op1_10_in19 = imem01_in[3:0];
    113: op1_10_in19 = reg_0786;
    114: op1_10_in19 = reg_0378;
    115: op1_10_in19 = reg_0583;
    118: op1_10_in19 = reg_0239;
    119: op1_10_in19 = reg_0261;
    120: op1_10_in19 = reg_0963;
    121: op1_10_in19 = reg_0420;
    122: op1_10_in19 = reg_0964;
    123: op1_10_in19 = reg_0067;
    125: op1_10_in19 = reg_0609;
    126: op1_10_in19 = reg_0291;
    127: op1_10_in19 = reg_0279;
    128: op1_10_in19 = reg_0376;
    129: op1_10_in19 = reg_0648;
    130: op1_10_in19 = reg_0013;
    131: op1_10_in19 = reg_0278;
    default: op1_10_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv19 = 1;
    53: op1_10_inv19 = 1;
    86: op1_10_inv19 = 1;
    55: op1_10_inv19 = 1;
    69: op1_10_inv19 = 1;
    74: op1_10_inv19 = 1;
    68: op1_10_inv19 = 1;
    71: op1_10_inv19 = 1;
    87: op1_10_inv19 = 1;
    76: op1_10_inv19 = 1;
    77: op1_10_inv19 = 1;
    60: op1_10_inv19 = 1;
    46: op1_10_inv19 = 1;
    64: op1_10_inv19 = 1;
    84: op1_10_inv19 = 1;
    48: op1_10_inv19 = 1;
    65: op1_10_inv19 = 1;
    91: op1_10_inv19 = 1;
    92: op1_10_inv19 = 1;
    95: op1_10_inv19 = 1;
    97: op1_10_inv19 = 1;
    98: op1_10_inv19 = 1;
    100: op1_10_inv19 = 1;
    102: op1_10_inv19 = 1;
    104: op1_10_inv19 = 1;
    106: op1_10_inv19 = 1;
    44: op1_10_inv19 = 1;
    107: op1_10_inv19 = 1;
    110: op1_10_inv19 = 1;
    111: op1_10_inv19 = 1;
    115: op1_10_inv19 = 1;
    120: op1_10_inv19 = 1;
    123: op1_10_inv19 = 1;
    127: op1_10_inv19 = 1;
    129: op1_10_inv19 = 1;
    default: op1_10_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in20 = reg_0039;
    53: op1_10_in20 = imem05_in[15:12];
    86: op1_10_in20 = reg_0113;
    96: op1_10_in20 = reg_0113;
    55: op1_10_in20 = reg_1169;
    73: op1_10_in20 = reg_1202;
    69: op1_10_in20 = reg_1384;
    49: op1_10_in20 = reg_0001;
    74: op1_10_in20 = reg_0158;
    54: op1_10_in20 = reg_0784;
    98: op1_10_in20 = reg_0784;
    68: op1_10_in20 = reg_0797;
    75: op1_10_in20 = reg_0134;
    50: op1_10_in20 = reg_0531;
    56: op1_10_in20 = reg_0418;
    71: op1_10_in20 = reg_0715;
    87: op1_10_in20 = reg_0020;
    76: op1_10_in20 = reg_1467;
    61: op1_10_in20 = reg_0434;
    57: op1_10_in20 = reg_1096;
    77: op1_10_in20 = reg_0146;
    58: op1_10_in20 = reg_0111;
    78: op1_10_in20 = reg_0922;
    70: op1_10_in20 = reg_0599;
    79: op1_10_in20 = reg_0863;
    59: op1_10_in20 = reg_0450;
    60: op1_10_in20 = reg_0313;
    126: op1_10_in20 = reg_0313;
    88: op1_10_in20 = reg_0337;
    92: op1_10_in20 = reg_0337;
    46: op1_10_in20 = reg_0702;
    80: op1_10_in20 = reg_1324;
    101: op1_10_in20 = reg_1324;
    81: op1_10_in20 = reg_0939;
    82: op1_10_in20 = reg_0310;
    89: op1_10_in20 = reg_1258;
    83: op1_10_in20 = reg_0335;
    64: op1_10_in20 = imem03_in[7:4];
    84: op1_10_in20 = reg_0049;
    100: op1_10_in20 = reg_0049;
    48: op1_10_in20 = reg_0017;
    85: op1_10_in20 = imem06_in[3:0];
    65: op1_10_in20 = reg_0087;
    90: op1_10_in20 = reg_0609;
    66: op1_10_in20 = reg_0254;
    91: op1_10_in20 = reg_1368;
    67: op1_10_in20 = reg_0258;
    93: op1_10_in20 = reg_0471;
    94: op1_10_in20 = reg_1140;
    95: op1_10_in20 = reg_0553;
    97: op1_10_in20 = reg_0444;
    102: op1_10_in20 = reg_1257;
    103: op1_10_in20 = reg_1504;
    104: op1_10_in20 = reg_0592;
    47: op1_10_in20 = reg_0960;
    105: op1_10_in20 = reg_0738;
    106: op1_10_in20 = reg_1078;
    44: op1_10_in20 = reg_0115;
    107: op1_10_in20 = reg_0600;
    108: op1_10_in20 = reg_0571;
    109: op1_10_in20 = reg_0908;
    110: op1_10_in20 = reg_1492;
    111: op1_10_in20 = reg_0569;
    112: op1_10_in20 = reg_1034;
    113: op1_10_in20 = reg_0170;
    114: op1_10_in20 = reg_1367;
    115: op1_10_in20 = reg_0754;
    116: op1_10_in20 = reg_1518;
    117: op1_10_in20 = reg_0518;
    118: op1_10_in20 = reg_0241;
    119: op1_10_in20 = reg_0216;
    120: op1_10_in20 = reg_0480;
    121: op1_10_in20 = reg_0633;
    122: op1_10_in20 = reg_0952;
    123: op1_10_in20 = reg_0213;
    124: op1_10_in20 = reg_1420;
    125: op1_10_in20 = reg_0242;
    127: op1_10_in20 = reg_0378;
    128: op1_10_in20 = reg_0108;
    129: op1_10_in20 = reg_0579;
    130: op1_10_in20 = reg_0331;
    42: op1_10_in20 = reg_0078;
    131: op1_10_in20 = reg_0648;
    default: op1_10_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv20 = 1;
    55: op1_10_inv20 = 1;
    73: op1_10_inv20 = 1;
    69: op1_10_inv20 = 1;
    68: op1_10_inv20 = 1;
    75: op1_10_inv20 = 1;
    50: op1_10_inv20 = 1;
    56: op1_10_inv20 = 1;
    71: op1_10_inv20 = 1;
    76: op1_10_inv20 = 1;
    61: op1_10_inv20 = 1;
    57: op1_10_inv20 = 1;
    77: op1_10_inv20 = 1;
    79: op1_10_inv20 = 1;
    59: op1_10_inv20 = 1;
    60: op1_10_inv20 = 1;
    89: op1_10_inv20 = 1;
    83: op1_10_inv20 = 1;
    85: op1_10_inv20 = 1;
    65: op1_10_inv20 = 1;
    67: op1_10_inv20 = 1;
    92: op1_10_inv20 = 1;
    94: op1_10_inv20 = 1;
    95: op1_10_inv20 = 1;
    96: op1_10_inv20 = 1;
    97: op1_10_inv20 = 1;
    100: op1_10_inv20 = 1;
    101: op1_10_inv20 = 1;
    102: op1_10_inv20 = 1;
    47: op1_10_inv20 = 1;
    44: op1_10_inv20 = 1;
    111: op1_10_inv20 = 1;
    114: op1_10_inv20 = 1;
    116: op1_10_inv20 = 1;
    117: op1_10_inv20 = 1;
    119: op1_10_inv20 = 1;
    120: op1_10_inv20 = 1;
    122: op1_10_inv20 = 1;
    125: op1_10_inv20 = 1;
    128: op1_10_inv20 = 1;
    129: op1_10_inv20 = 1;
    42: op1_10_inv20 = 1;
    131: op1_10_inv20 = 1;
    default: op1_10_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in21 = reg_0458;
    53: op1_10_in21 = reg_0347;
    86: op1_10_in21 = reg_0885;
    96: op1_10_in21 = reg_0885;
    55: op1_10_in21 = reg_0346;
    73: op1_10_in21 = reg_1179;
    69: op1_10_in21 = reg_0263;
    49: op1_10_in21 = reg_0086;
    74: op1_10_in21 = reg_0921;
    54: op1_10_in21 = reg_0782;
    68: op1_10_in21 = reg_0936;
    75: op1_10_in21 = reg_0389;
    50: op1_10_in21 = reg_0497;
    56: op1_10_in21 = reg_0303;
    71: op1_10_in21 = reg_0469;
    87: op1_10_in21 = reg_0470;
    76: op1_10_in21 = imem06_in[7:4];
    85: op1_10_in21 = imem06_in[7:4];
    61: op1_10_in21 = reg_0147;
    57: op1_10_in21 = reg_1183;
    77: op1_10_in21 = reg_0091;
    58: op1_10_in21 = reg_0381;
    78: op1_10_in21 = reg_0894;
    70: op1_10_in21 = reg_0320;
    79: op1_10_in21 = reg_1504;
    59: op1_10_in21 = reg_0301;
    60: op1_10_in21 = reg_0218;
    88: op1_10_in21 = reg_0336;
    46: op1_10_in21 = reg_0603;
    80: op1_10_in21 = reg_0122;
    81: op1_10_in21 = reg_0418;
    82: op1_10_in21 = reg_0245;
    89: op1_10_in21 = reg_1203;
    83: op1_10_in21 = reg_0982;
    64: op1_10_in21 = imem03_in[11:8];
    84: op1_10_in21 = reg_0198;
    48: op1_10_in21 = imem07_in[3:0];
    65: op1_10_in21 = reg_0483;
    117: op1_10_in21 = reg_0483;
    90: op1_10_in21 = reg_0572;
    66: op1_10_in21 = reg_1260;
    91: op1_10_in21 = reg_1367;
    67: op1_10_in21 = reg_0548;
    92: op1_10_in21 = reg_0338;
    93: op1_10_in21 = reg_0452;
    94: op1_10_in21 = reg_0306;
    95: op1_10_in21 = reg_0463;
    97: op1_10_in21 = reg_0573;
    98: op1_10_in21 = reg_0193;
    100: op1_10_in21 = reg_0847;
    101: op1_10_in21 = imem01_in[15:12];
    102: op1_10_in21 = reg_0552;
    103: op1_10_in21 = reg_0172;
    104: op1_10_in21 = reg_0100;
    47: op1_10_in21 = reg_0866;
    105: op1_10_in21 = reg_0415;
    106: op1_10_in21 = reg_1006;
    44: op1_10_in21 = reg_0264;
    107: op1_10_in21 = reg_0789;
    108: op1_10_in21 = reg_0289;
    109: op1_10_in21 = reg_0905;
    110: op1_10_in21 = reg_0802;
    111: op1_10_in21 = reg_0119;
    112: op1_10_in21 = reg_0930;
    113: op1_10_in21 = reg_0156;
    114: op1_10_in21 = reg_0535;
    115: op1_10_in21 = reg_0977;
    116: op1_10_in21 = reg_0957;
    118: op1_10_in21 = reg_0830;
    119: op1_10_in21 = reg_0600;
    120: op1_10_in21 = imem03_in[7:4];
    121: op1_10_in21 = reg_0020;
    122: op1_10_in21 = reg_1231;
    123: op1_10_in21 = reg_0518;
    124: op1_10_in21 = reg_0271;
    125: op1_10_in21 = reg_0241;
    126: op1_10_in21 = reg_0443;
    127: op1_10_in21 = reg_0234;
    128: op1_10_in21 = reg_0831;
    129: op1_10_in21 = reg_0702;
    130: op1_10_in21 = reg_0222;
    42: op1_10_in21 = reg_0079;
    131: op1_10_in21 = reg_0986;
    default: op1_10_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_10_inv21 = 1;
    49: op1_10_inv21 = 1;
    68: op1_10_inv21 = 1;
    75: op1_10_inv21 = 1;
    56: op1_10_inv21 = 1;
    71: op1_10_inv21 = 1;
    61: op1_10_inv21 = 1;
    77: op1_10_inv21 = 1;
    58: op1_10_inv21 = 1;
    88: op1_10_inv21 = 1;
    80: op1_10_inv21 = 1;
    81: op1_10_inv21 = 1;
    64: op1_10_inv21 = 1;
    84: op1_10_inv21 = 1;
    90: op1_10_inv21 = 1;
    66: op1_10_inv21 = 1;
    93: op1_10_inv21 = 1;
    94: op1_10_inv21 = 1;
    96: op1_10_inv21 = 1;
    98: op1_10_inv21 = 1;
    100: op1_10_inv21 = 1;
    103: op1_10_inv21 = 1;
    104: op1_10_inv21 = 1;
    47: op1_10_inv21 = 1;
    106: op1_10_inv21 = 1;
    108: op1_10_inv21 = 1;
    109: op1_10_inv21 = 1;
    112: op1_10_inv21 = 1;
    116: op1_10_inv21 = 1;
    117: op1_10_inv21 = 1;
    119: op1_10_inv21 = 1;
    126: op1_10_inv21 = 1;
    129: op1_10_inv21 = 1;
    42: op1_10_inv21 = 1;
    default: op1_10_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in22 = reg_0195;
    53: op1_10_in22 = reg_0648;
    55: op1_10_in22 = reg_0648;
    86: op1_10_in22 = reg_0884;
    73: op1_10_in22 = reg_0215;
    69: op1_10_in22 = reg_1372;
    49: op1_10_in22 = reg_0084;
    104: op1_10_in22 = reg_0084;
    74: op1_10_in22 = reg_1094;
    54: op1_10_in22 = reg_1058;
    68: op1_10_in22 = reg_0451;
    75: op1_10_in22 = reg_0059;
    50: op1_10_in22 = reg_0495;
    56: op1_10_in22 = reg_0300;
    71: op1_10_in22 = reg_0968;
    87: op1_10_in22 = reg_0205;
    76: op1_10_in22 = reg_0974;
    61: op1_10_in22 = reg_0902;
    57: op1_10_in22 = reg_0224;
    77: op1_10_in22 = reg_0901;
    58: op1_10_in22 = reg_0138;
    78: op1_10_in22 = reg_0703;
    82: op1_10_in22 = reg_0703;
    70: op1_10_in22 = reg_1419;
    79: op1_10_in22 = reg_0161;
    59: op1_10_in22 = reg_0090;
    60: op1_10_in22 = reg_0444;
    88: op1_10_in22 = reg_1151;
    46: op1_10_in22 = reg_0066;
    80: op1_10_in22 = reg_0917;
    81: op1_10_in22 = reg_1486;
    89: op1_10_in22 = reg_1198;
    83: op1_10_in22 = reg_1255;
    64: op1_10_in22 = imem03_in[15:12];
    84: op1_10_in22 = reg_1001;
    48: op1_10_in22 = reg_0225;
    85: op1_10_in22 = reg_0827;
    65: op1_10_in22 = reg_1182;
    90: op1_10_in22 = reg_0402;
    66: op1_10_in22 = reg_0475;
    91: op1_10_in22 = reg_0034;
    67: op1_10_in22 = reg_0819;
    92: op1_10_in22 = reg_0236;
    93: op1_10_in22 = reg_1107;
    94: op1_10_in22 = reg_0560;
    95: op1_10_in22 = reg_0547;
    96: op1_10_in22 = reg_0880;
    97: op1_10_in22 = reg_0261;
    98: op1_10_in22 = reg_0906;
    100: op1_10_in22 = reg_0600;
    101: op1_10_in22 = reg_1032;
    102: op1_10_in22 = reg_1200;
    103: op1_10_in22 = reg_1179;
    47: op1_10_in22 = reg_0635;
    105: op1_10_in22 = reg_0593;
    106: op1_10_in22 = reg_0217;
    44: op1_10_in22 = reg_0624;
    107: op1_10_in22 = reg_0142;
    108: op1_10_in22 = reg_0244;
    109: op1_10_in22 = reg_0696;
    110: op1_10_in22 = reg_0711;
    111: op1_10_in22 = reg_0165;
    112: op1_10_in22 = reg_0463;
    113: op1_10_in22 = reg_0157;
    114: op1_10_in22 = reg_0088;
    115: op1_10_in22 = reg_0067;
    116: op1_10_in22 = reg_1447;
    117: op1_10_in22 = reg_0123;
    118: op1_10_in22 = reg_0715;
    119: op1_10_in22 = reg_0312;
    120: op1_10_in22 = reg_0989;
    121: op1_10_in22 = reg_0210;
    122: op1_10_in22 = reg_1208;
    123: op1_10_in22 = reg_0169;
    124: op1_10_in22 = reg_1467;
    125: op1_10_in22 = reg_0830;
    130: op1_10_in22 = reg_0830;
    126: op1_10_in22 = imem04_in[3:0];
    127: op1_10_in22 = reg_1495;
    128: op1_10_in22 = reg_0291;
    129: op1_10_in22 = reg_1168;
    42: op1_10_in22 = reg_0290;
    131: op1_10_in22 = reg_0735;
    default: op1_10_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv22 = 1;
    73: op1_10_inv22 = 1;
    69: op1_10_inv22 = 1;
    74: op1_10_inv22 = 1;
    54: op1_10_inv22 = 1;
    75: op1_10_inv22 = 1;
    50: op1_10_inv22 = 1;
    56: op1_10_inv22 = 1;
    57: op1_10_inv22 = 1;
    77: op1_10_inv22 = 1;
    78: op1_10_inv22 = 1;
    81: op1_10_inv22 = 1;
    64: op1_10_inv22 = 1;
    84: op1_10_inv22 = 1;
    85: op1_10_inv22 = 1;
    65: op1_10_inv22 = 1;
    67: op1_10_inv22 = 1;
    92: op1_10_inv22 = 1;
    93: op1_10_inv22 = 1;
    95: op1_10_inv22 = 1;
    96: op1_10_inv22 = 1;
    97: op1_10_inv22 = 1;
    98: op1_10_inv22 = 1;
    102: op1_10_inv22 = 1;
    104: op1_10_inv22 = 1;
    105: op1_10_inv22 = 1;
    112: op1_10_inv22 = 1;
    116: op1_10_inv22 = 1;
    117: op1_10_inv22 = 1;
    122: op1_10_inv22 = 1;
    123: op1_10_inv22 = 1;
    124: op1_10_inv22 = 1;
    128: op1_10_inv22 = 1;
    129: op1_10_inv22 = 1;
    42: op1_10_inv22 = 1;
    default: op1_10_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in23 = reg_0755;
    53: op1_10_in23 = reg_0566;
    86: op1_10_in23 = reg_0411;
    55: op1_10_in23 = reg_0996;
    73: op1_10_in23 = reg_0213;
    69: op1_10_in23 = reg_1215;
    49: op1_10_in23 = reg_0087;
    104: op1_10_in23 = reg_0087;
    123: op1_10_in23 = reg_0087;
    74: op1_10_in23 = reg_0775;
    54: op1_10_in23 = reg_0720;
    68: op1_10_in23 = reg_0452;
    75: op1_10_in23 = reg_0005;
    50: op1_10_in23 = reg_0472;
    56: op1_10_in23 = reg_0873;
    59: op1_10_in23 = reg_0873;
    71: op1_10_in23 = reg_0430;
    87: op1_10_in23 = reg_0578;
    76: op1_10_in23 = reg_0133;
    61: op1_10_in23 = reg_0088;
    57: op1_10_in23 = reg_0703;
    77: op1_10_in23 = reg_0724;
    58: op1_10_in23 = reg_0307;
    78: op1_10_in23 = reg_0170;
    70: op1_10_in23 = reg_0369;
    79: op1_10_in23 = reg_0115;
    60: op1_10_in23 = reg_1064;
    88: op1_10_in23 = reg_1189;
    46: op1_10_in23 = reg_0182;
    80: op1_10_in23 = imem01_in[7:4];
    81: op1_10_in23 = reg_0492;
    82: op1_10_in23 = reg_1347;
    89: op1_10_in23 = reg_0488;
    83: op1_10_in23 = reg_0754;
    64: op1_10_in23 = reg_0234;
    84: op1_10_in23 = reg_0541;
    48: op1_10_in23 = reg_0226;
    85: op1_10_in23 = reg_0635;
    65: op1_10_in23 = reg_0618;
    90: op1_10_in23 = reg_0464;
    66: op1_10_in23 = reg_1207;
    91: op1_10_in23 = reg_0252;
    67: op1_10_in23 = reg_0149;
    92: op1_10_in23 = reg_0016;
    93: op1_10_in23 = reg_0536;
    94: op1_10_in23 = reg_1098;
    95: op1_10_in23 = reg_0747;
    96: op1_10_in23 = reg_0291;
    97: op1_10_in23 = reg_1001;
    98: op1_10_in23 = reg_0397;
    100: op1_10_in23 = reg_0142;
    101: op1_10_in23 = reg_0282;
    102: op1_10_in23 = reg_0062;
    103: op1_10_in23 = reg_0116;
    47: op1_10_in23 = reg_0636;
    105: op1_10_in23 = reg_0001;
    106: op1_10_in23 = reg_0632;
    44: op1_10_in23 = reg_0526;
    107: op1_10_in23 = reg_1208;
    108: op1_10_in23 = reg_0165;
    109: op1_10_in23 = reg_1467;
    110: op1_10_in23 = reg_0479;
    111: op1_10_in23 = reg_0046;
    112: op1_10_in23 = reg_0746;
    113: op1_10_in23 = reg_0661;
    114: op1_10_in23 = reg_0694;
    115: op1_10_in23 = imem07_in[11:8];
    116: op1_10_in23 = reg_0048;
    117: op1_10_in23 = reg_1182;
    118: op1_10_in23 = reg_0967;
    119: op1_10_in23 = reg_0000;
    120: op1_10_in23 = reg_0233;
    121: op1_10_in23 = reg_0315;
    122: op1_10_in23 = reg_0108;
    124: op1_10_in23 = reg_1505;
    125: op1_10_in23 = reg_1474;
    126: op1_10_in23 = reg_0129;
    127: op1_10_in23 = reg_1518;
    128: op1_10_in23 = imem04_in[7:4];
    129: op1_10_in23 = reg_0890;
    130: op1_10_in23 = reg_0820;
    42: op1_10_in23 = reg_0042;
    131: op1_10_in23 = reg_0702;
    default: op1_10_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_10_inv23 = 1;
    55: op1_10_inv23 = 1;
    49: op1_10_inv23 = 1;
    54: op1_10_inv23 = 1;
    61: op1_10_inv23 = 1;
    77: op1_10_inv23 = 1;
    58: op1_10_inv23 = 1;
    79: op1_10_inv23 = 1;
    60: op1_10_inv23 = 1;
    80: op1_10_inv23 = 1;
    81: op1_10_inv23 = 1;
    82: op1_10_inv23 = 1;
    89: op1_10_inv23 = 1;
    84: op1_10_inv23 = 1;
    85: op1_10_inv23 = 1;
    91: op1_10_inv23 = 1;
    92: op1_10_inv23 = 1;
    96: op1_10_inv23 = 1;
    97: op1_10_inv23 = 1;
    102: op1_10_inv23 = 1;
    47: op1_10_inv23 = 1;
    105: op1_10_inv23 = 1;
    44: op1_10_inv23 = 1;
    111: op1_10_inv23 = 1;
    112: op1_10_inv23 = 1;
    113: op1_10_inv23 = 1;
    114: op1_10_inv23 = 1;
    115: op1_10_inv23 = 1;
    116: op1_10_inv23 = 1;
    119: op1_10_inv23 = 1;
    120: op1_10_inv23 = 1;
    124: op1_10_inv23 = 1;
    125: op1_10_inv23 = 1;
    126: op1_10_inv23 = 1;
    129: op1_10_inv23 = 1;
    default: op1_10_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in24 = reg_1437;
    53: op1_10_in24 = reg_0045;
    86: op1_10_in24 = reg_0263;
    55: op1_10_in24 = reg_1181;
    73: op1_10_in24 = reg_0018;
    69: op1_10_in24 = reg_1198;
    49: op1_10_in24 = reg_0484;
    74: op1_10_in24 = reg_0442;
    54: op1_10_in24 = reg_0372;
    68: op1_10_in24 = imem04_in[11:8];
    75: op1_10_in24 = reg_0917;
    50: op1_10_in24 = reg_0473;
    56: op1_10_in24 = reg_0251;
    71: op1_10_in24 = reg_0149;
    87: op1_10_in24 = reg_0204;
    76: op1_10_in24 = reg_0397;
    61: op1_10_in24 = reg_0277;
    57: op1_10_in24 = reg_0299;
    77: op1_10_in24 = reg_0896;
    58: op1_10_in24 = reg_0294;
    78: op1_10_in24 = reg_0158;
    70: op1_10_in24 = reg_0304;
    79: op1_10_in24 = reg_0373;
    59: op1_10_in24 = reg_0243;
    60: op1_10_in24 = reg_1149;
    88: op1_10_in24 = reg_1107;
    46: op1_10_in24 = imem05_in[15:12];
    80: op1_10_in24 = reg_0788;
    81: op1_10_in24 = reg_0196;
    82: op1_10_in24 = reg_0779;
    89: op1_10_in24 = reg_1147;
    83: op1_10_in24 = reg_1512;
    64: op1_10_in24 = reg_0954;
    84: op1_10_in24 = reg_0375;
    48: op1_10_in24 = reg_0893;
    85: op1_10_in24 = reg_0116;
    90: op1_10_in24 = reg_0080;
    66: op1_10_in24 = reg_0433;
    91: op1_10_in24 = reg_1257;
    114: op1_10_in24 = reg_1257;
    67: op1_10_in24 = imem01_in[11:8];
    92: op1_10_in24 = reg_1488;
    93: op1_10_in24 = reg_1503;
    94: op1_10_in24 = reg_0711;
    95: op1_10_in24 = reg_0222;
    96: op1_10_in24 = reg_0313;
    97: op1_10_in24 = reg_1495;
    98: op1_10_in24 = reg_0925;
    100: op1_10_in24 = reg_1314;
    101: op1_10_in24 = reg_0553;
    102: op1_10_in24 = reg_0862;
    103: op1_10_in24 = reg_0398;
    104: op1_10_in24 = reg_0483;
    47: op1_10_in24 = reg_0569;
    105: op1_10_in24 = reg_0520;
    106: op1_10_in24 = reg_0049;
    44: op1_10_in24 = reg_0522;
    107: op1_10_in24 = reg_0108;
    108: op1_10_in24 = reg_1202;
    109: op1_10_in24 = reg_0869;
    110: op1_10_in24 = reg_0246;
    111: op1_10_in24 = reg_0084;
    112: op1_10_in24 = reg_0743;
    113: op1_10_in24 = reg_0663;
    115: op1_10_in24 = reg_0298;
    116: op1_10_in24 = reg_0329;
    118: op1_10_in24 = reg_0439;
    119: op1_10_in24 = reg_0180;
    120: op1_10_in24 = reg_1001;
    121: op1_10_in24 = imem05_in[11:8];
    122: op1_10_in24 = reg_0113;
    123: op1_10_in24 = imem07_in[3:0];
    124: op1_10_in24 = reg_0265;
    125: op1_10_in24 = reg_0819;
    126: op1_10_in24 = reg_0534;
    127: op1_10_in24 = reg_0627;
    128: op1_10_in24 = reg_1384;
    129: op1_10_in24 = reg_0346;
    130: op1_10_in24 = reg_0438;
    42: op1_10_in24 = reg_0011;
    131: op1_10_in24 = reg_0040;
    default: op1_10_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv24 = 1;
    55: op1_10_inv24 = 1;
    69: op1_10_inv24 = 1;
    49: op1_10_inv24 = 1;
    74: op1_10_inv24 = 1;
    54: op1_10_inv24 = 1;
    68: op1_10_inv24 = 1;
    75: op1_10_inv24 = 1;
    50: op1_10_inv24 = 1;
    56: op1_10_inv24 = 1;
    76: op1_10_inv24 = 1;
    61: op1_10_inv24 = 1;
    57: op1_10_inv24 = 1;
    58: op1_10_inv24 = 1;
    78: op1_10_inv24 = 1;
    70: op1_10_inv24 = 1;
    79: op1_10_inv24 = 1;
    88: op1_10_inv24 = 1;
    46: op1_10_inv24 = 1;
    89: op1_10_inv24 = 1;
    64: op1_10_inv24 = 1;
    48: op1_10_inv24 = 1;
    92: op1_10_inv24 = 1;
    93: op1_10_inv24 = 1;
    97: op1_10_inv24 = 1;
    98: op1_10_inv24 = 1;
    100: op1_10_inv24 = 1;
    101: op1_10_inv24 = 1;
    103: op1_10_inv24 = 1;
    104: op1_10_inv24 = 1;
    47: op1_10_inv24 = 1;
    106: op1_10_inv24 = 1;
    107: op1_10_inv24 = 1;
    114: op1_10_inv24 = 1;
    115: op1_10_inv24 = 1;
    123: op1_10_inv24 = 1;
    124: op1_10_inv24 = 1;
    127: op1_10_inv24 = 1;
    129: op1_10_inv24 = 1;
    default: op1_10_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in25 = reg_0192;
    53: op1_10_in25 = reg_0316;
    86: op1_10_in25 = reg_1372;
    55: op1_10_in25 = reg_0318;
    73: op1_10_in25 = reg_0017;
    69: op1_10_in25 = reg_1200;
    74: op1_10_in25 = reg_0739;
    54: op1_10_in25 = reg_0827;
    68: op1_10_in25 = imem04_in[15:12];
    75: op1_10_in25 = reg_1068;
    50: op1_10_in25 = reg_0433;
    56: op1_10_in25 = reg_0168;
    71: op1_10_in25 = reg_0148;
    87: op1_10_in25 = reg_0832;
    76: op1_10_in25 = reg_0160;
    61: op1_10_in25 = reg_0486;
    57: op1_10_in25 = reg_0924;
    77: op1_10_in25 = reg_0679;
    42: op1_10_in25 = reg_0679;
    58: op1_10_in25 = reg_0879;
    78: op1_10_in25 = reg_0223;
    70: op1_10_in25 = reg_0836;
    79: op1_10_in25 = reg_0584;
    59: op1_10_in25 = reg_0864;
    60: op1_10_in25 = reg_0049;
    88: op1_10_in25 = reg_1502;
    46: op1_10_in25 = reg_0163;
    80: op1_10_in25 = reg_0277;
    81: op1_10_in25 = reg_0589;
    82: op1_10_in25 = reg_0663;
    89: op1_10_in25 = reg_0421;
    83: op1_10_in25 = reg_0047;
    64: op1_10_in25 = reg_0246;
    84: op1_10_in25 = reg_0965;
    48: op1_10_in25 = reg_0867;
    85: op1_10_in25 = reg_0714;
    90: op1_10_in25 = reg_0257;
    66: op1_10_in25 = reg_0054;
    91: op1_10_in25 = reg_1233;
    67: op1_10_in25 = reg_0874;
    92: op1_10_in25 = reg_0737;
    93: op1_10_in25 = reg_0016;
    94: op1_10_in25 = reg_0007;
    95: op1_10_in25 = reg_0830;
    96: op1_10_in25 = reg_1139;
    97: op1_10_in25 = reg_0349;
    98: op1_10_in25 = reg_0870;
    100: op1_10_in25 = reg_1313;
    101: op1_10_in25 = reg_0463;
    102: op1_10_in25 = reg_0096;
    103: op1_10_in25 = reg_0585;
    104: op1_10_in25 = reg_1182;
    47: op1_10_in25 = imem07_in[3:0];
    106: op1_10_in25 = reg_0154;
    44: op1_10_in25 = reg_0295;
    107: op1_10_in25 = reg_0448;
    108: op1_10_in25 = reg_0754;
    109: op1_10_in25 = reg_1501;
    110: op1_10_in25 = reg_1003;
    111: op1_10_in25 = reg_0226;
    112: op1_10_in25 = reg_0798;
    113: op1_10_in25 = reg_0437;
    114: op1_10_in25 = reg_0412;
    115: op1_10_in25 = reg_0310;
    116: op1_10_in25 = reg_1231;
    118: op1_10_in25 = reg_0868;
    119: op1_10_in25 = reg_0070;
    120: op1_10_in25 = reg_0312;
    121: op1_10_in25 = reg_0890;
    122: op1_10_in25 = reg_0885;
    123: op1_10_in25 = reg_0170;
    124: op1_10_in25 = reg_0115;
    125: op1_10_in25 = reg_0430;
    126: op1_10_in25 = reg_0535;
    127: op1_10_in25 = reg_0290;
    128: op1_10_in25 = reg_0252;
    129: op1_10_in25 = reg_0733;
    131: op1_10_in25 = reg_0733;
    130: op1_10_in25 = reg_1457;
    default: op1_10_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv25 = 1;
    53: op1_10_inv25 = 1;
    86: op1_10_inv25 = 1;
    55: op1_10_inv25 = 1;
    68: op1_10_inv25 = 1;
    56: op1_10_inv25 = 1;
    71: op1_10_inv25 = 1;
    76: op1_10_inv25 = 1;
    61: op1_10_inv25 = 1;
    58: op1_10_inv25 = 1;
    78: op1_10_inv25 = 1;
    81: op1_10_inv25 = 1;
    82: op1_10_inv25 = 1;
    89: op1_10_inv25 = 1;
    85: op1_10_inv25 = 1;
    91: op1_10_inv25 = 1;
    67: op1_10_inv25 = 1;
    93: op1_10_inv25 = 1;
    97: op1_10_inv25 = 1;
    103: op1_10_inv25 = 1;
    47: op1_10_inv25 = 1;
    106: op1_10_inv25 = 1;
    44: op1_10_inv25 = 1;
    112: op1_10_inv25 = 1;
    113: op1_10_inv25 = 1;
    115: op1_10_inv25 = 1;
    116: op1_10_inv25 = 1;
    118: op1_10_inv25 = 1;
    120: op1_10_inv25 = 1;
    122: op1_10_inv25 = 1;
    124: op1_10_inv25 = 1;
    126: op1_10_inv25 = 1;
    127: op1_10_inv25 = 1;
    128: op1_10_inv25 = 1;
    131: op1_10_inv25 = 1;
    default: op1_10_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in26 = reg_0907;
    53: op1_10_in26 = reg_0540;
    86: op1_10_in26 = reg_0181;
    55: op1_10_in26 = reg_0539;
    73: op1_10_in26 = reg_0226;
    47: op1_10_in26 = reg_0226;
    69: op1_10_in26 = reg_0676;
    74: op1_10_in26 = reg_0621;
    54: op1_10_in26 = reg_0718;
    124: op1_10_in26 = reg_0718;
    68: op1_10_in26 = reg_0338;
    75: op1_10_in26 = reg_1071;
    50: op1_10_in26 = reg_0972;
    56: op1_10_in26 = reg_0240;
    71: op1_10_in26 = reg_0400;
    87: op1_10_in26 = imem05_in[3:0];
    76: op1_10_in26 = reg_0172;
    61: op1_10_in26 = reg_0632;
    57: op1_10_in26 = reg_0139;
    77: op1_10_in26 = reg_0457;
    58: op1_10_in26 = reg_0839;
    78: op1_10_in26 = reg_0777;
    70: op1_10_in26 = reg_0096;
    79: op1_10_in26 = reg_0619;
    59: op1_10_in26 = reg_0449;
    60: op1_10_in26 = reg_0234;
    88: op1_10_in26 = reg_0019;
    46: op1_10_in26 = reg_0450;
    80: op1_10_in26 = reg_1511;
    81: op1_10_in26 = reg_0207;
    82: op1_10_in26 = reg_0740;
    89: op1_10_in26 = reg_1040;
    83: op1_10_in26 = reg_1474;
    64: op1_10_in26 = reg_1300;
    84: op1_10_in26 = reg_1314;
    119: op1_10_in26 = reg_1314;
    48: op1_10_in26 = reg_0299;
    85: op1_10_in26 = reg_0528;
    90: op1_10_in26 = reg_1068;
    66: op1_10_in26 = reg_0326;
    91: op1_10_in26 = reg_0281;
    67: op1_10_in26 = reg_0077;
    92: op1_10_in26 = reg_0204;
    93: op1_10_in26 = reg_0370;
    94: op1_10_in26 = reg_0279;
    95: op1_10_in26 = reg_0820;
    96: op1_10_in26 = reg_1280;
    97: op1_10_in26 = reg_0558;
    98: op1_10_in26 = reg_1209;
    100: op1_10_in26 = reg_0220;
    101: op1_10_in26 = reg_0163;
    102: op1_10_in26 = reg_1189;
    103: op1_10_in26 = reg_0165;
    106: op1_10_in26 = reg_0706;
    44: op1_10_in26 = reg_0458;
    107: op1_10_in26 = reg_0378;
    108: op1_10_in26 = reg_0213;
    109: op1_10_in26 = reg_0780;
    110: op1_10_in26 = reg_1063;
    111: op1_10_in26 = imem07_in[7:4];
    112: op1_10_in26 = reg_0434;
    113: op1_10_in26 = reg_0404;
    114: op1_10_in26 = reg_1041;
    115: op1_10_in26 = reg_0786;
    116: op1_10_in26 = reg_1325;
    118: op1_10_in26 = reg_0385;
    120: op1_10_in26 = reg_0789;
    121: op1_10_in26 = reg_0205;
    131: op1_10_in26 = reg_0205;
    122: op1_10_in26 = reg_0448;
    123: op1_10_in26 = reg_1349;
    125: op1_10_in26 = reg_0146;
    126: op1_10_in26 = reg_0797;
    127: op1_10_in26 = reg_1199;
    128: op1_10_in26 = reg_1216;
    129: op1_10_in26 = reg_0272;
    130: op1_10_in26 = reg_1034;
    42: op1_10_in26 = reg_0446;
    default: op1_10_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_10_inv26 = 1;
    69: op1_10_inv26 = 1;
    74: op1_10_inv26 = 1;
    54: op1_10_inv26 = 1;
    68: op1_10_inv26 = 1;
    50: op1_10_inv26 = 1;
    71: op1_10_inv26 = 1;
    61: op1_10_inv26 = 1;
    57: op1_10_inv26 = 1;
    78: op1_10_inv26 = 1;
    70: op1_10_inv26 = 1;
    79: op1_10_inv26 = 1;
    59: op1_10_inv26 = 1;
    88: op1_10_inv26 = 1;
    46: op1_10_inv26 = 1;
    80: op1_10_inv26 = 1;
    83: op1_10_inv26 = 1;
    64: op1_10_inv26 = 1;
    84: op1_10_inv26 = 1;
    90: op1_10_inv26 = 1;
    67: op1_10_inv26 = 1;
    92: op1_10_inv26 = 1;
    94: op1_10_inv26 = 1;
    95: op1_10_inv26 = 1;
    98: op1_10_inv26 = 1;
    102: op1_10_inv26 = 1;
    103: op1_10_inv26 = 1;
    47: op1_10_inv26 = 1;
    106: op1_10_inv26 = 1;
    107: op1_10_inv26 = 1;
    108: op1_10_inv26 = 1;
    110: op1_10_inv26 = 1;
    112: op1_10_inv26 = 1;
    121: op1_10_inv26 = 1;
    123: op1_10_inv26 = 1;
    127: op1_10_inv26 = 1;
    128: op1_10_inv26 = 1;
    129: op1_10_inv26 = 1;
    130: op1_10_inv26 = 1;
    131: op1_10_inv26 = 1;
    default: op1_10_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in27 = reg_0172;
    53: op1_10_in27 = reg_0939;
    86: op1_10_in27 = imem04_in[3:0];
    55: op1_10_in27 = reg_0938;
    73: op1_10_in27 = reg_1416;
    69: op1_10_in27 = reg_0464;
    118: op1_10_in27 = reg_0464;
    74: op1_10_in27 = reg_0620;
    54: op1_10_in27 = reg_0634;
    68: op1_10_in27 = reg_0210;
    75: op1_10_in27 = reg_0093;
    50: op1_10_in27 = reg_0125;
    56: op1_10_in27 = reg_0037;
    71: op1_10_in27 = reg_0091;
    87: op1_10_in27 = reg_0333;
    76: op1_10_in27 = reg_0109;
    61: op1_10_in27 = reg_0455;
    57: op1_10_in27 = reg_0779;
    77: op1_10_in27 = reg_1029;
    58: op1_10_in27 = reg_0845;
    78: op1_10_in27 = reg_0665;
    70: op1_10_in27 = reg_0095;
    79: op1_10_in27 = reg_0624;
    59: op1_10_in27 = reg_0205;
    60: op1_10_in27 = reg_1001;
    88: op1_10_in27 = reg_0470;
    46: op1_10_in27 = reg_0183;
    80: op1_10_in27 = reg_0548;
    81: op1_10_in27 = reg_0014;
    82: op1_10_in27 = reg_0593;
    89: op1_10_in27 = reg_0033;
    83: op1_10_in27 = reg_0469;
    95: op1_10_in27 = reg_0469;
    64: op1_10_in27 = reg_1301;
    84: op1_10_in27 = reg_0957;
    48: op1_10_in27 = reg_0309;
    85: op1_10_in27 = reg_0569;
    90: op1_10_in27 = reg_0626;
    66: op1_10_in27 = reg_0626;
    91: op1_10_in27 = reg_1082;
    67: op1_10_in27 = reg_0290;
    92: op1_10_in27 = reg_1430;
    93: op1_10_in27 = reg_0136;
    94: op1_10_in27 = reg_0255;
    96: op1_10_in27 = reg_0348;
    97: op1_10_in27 = reg_0108;
    98: op1_10_in27 = reg_0960;
    100: op1_10_in27 = reg_1300;
    101: op1_10_in27 = reg_0239;
    102: op1_10_in27 = reg_0064;
    103: op1_10_in27 = reg_1204;
    47: op1_10_in27 = reg_0894;
    106: op1_10_in27 = reg_0600;
    44: op1_10_in27 = reg_0459;
    107: op1_10_in27 = reg_0025;
    108: op1_10_in27 = reg_0015;
    109: op1_10_in27 = reg_0398;
    110: op1_10_in27 = reg_1425;
    111: op1_10_in27 = reg_0786;
    112: op1_10_in27 = reg_1457;
    113: op1_10_in27 = reg_0408;
    114: op1_10_in27 = reg_0537;
    115: op1_10_in27 = reg_1056;
    116: op1_10_in27 = reg_1282;
    119: op1_10_in27 = reg_1313;
    120: op1_10_in27 = reg_1495;
    121: op1_10_in27 = reg_0182;
    122: op1_10_in27 = reg_0291;
    123: op1_10_in27 = reg_0156;
    124: op1_10_in27 = reg_0194;
    125: op1_10_in27 = reg_1032;
    126: op1_10_in27 = reg_1083;
    127: op1_10_in27 = reg_0350;
    128: op1_10_in27 = reg_0978;
    129: op1_10_in27 = reg_0996;
    130: op1_10_in27 = reg_0963;
    42: op1_10_in27 = reg_0662;
    131: op1_10_in27 = reg_0176;
    default: op1_10_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv27 = 1;
    53: op1_10_inv27 = 1;
    55: op1_10_inv27 = 1;
    69: op1_10_inv27 = 1;
    54: op1_10_inv27 = 1;
    68: op1_10_inv27 = 1;
    50: op1_10_inv27 = 1;
    87: op1_10_inv27 = 1;
    76: op1_10_inv27 = 1;
    61: op1_10_inv27 = 1;
    57: op1_10_inv27 = 1;
    70: op1_10_inv27 = 1;
    88: op1_10_inv27 = 1;
    46: op1_10_inv27 = 1;
    80: op1_10_inv27 = 1;
    81: op1_10_inv27 = 1;
    64: op1_10_inv27 = 1;
    84: op1_10_inv27 = 1;
    48: op1_10_inv27 = 1;
    85: op1_10_inv27 = 1;
    91: op1_10_inv27 = 1;
    67: op1_10_inv27 = 1;
    92: op1_10_inv27 = 1;
    94: op1_10_inv27 = 1;
    95: op1_10_inv27 = 1;
    97: op1_10_inv27 = 1;
    101: op1_10_inv27 = 1;
    102: op1_10_inv27 = 1;
    103: op1_10_inv27 = 1;
    47: op1_10_inv27 = 1;
    44: op1_10_inv27 = 1;
    107: op1_10_inv27 = 1;
    109: op1_10_inv27 = 1;
    110: op1_10_inv27 = 1;
    112: op1_10_inv27 = 1;
    113: op1_10_inv27 = 1;
    118: op1_10_inv27 = 1;
    119: op1_10_inv27 = 1;
    120: op1_10_inv27 = 1;
    122: op1_10_inv27 = 1;
    124: op1_10_inv27 = 1;
    126: op1_10_inv27 = 1;
    131: op1_10_inv27 = 1;
    default: op1_10_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in28 = reg_1334;
    53: op1_10_in28 = reg_0163;
    86: op1_10_in28 = imem04_in[7:4];
    55: op1_10_in28 = reg_0450;
    73: op1_10_in28 = reg_0673;
    69: op1_10_in28 = reg_0421;
    91: op1_10_in28 = reg_0421;
    74: op1_10_in28 = reg_0003;
    54: op1_10_in28 = reg_0529;
    68: op1_10_in28 = reg_0064;
    75: op1_10_in28 = reg_0550;
    50: op1_10_in28 = reg_0126;
    56: op1_10_in28 = reg_0039;
    71: op1_10_in28 = reg_0899;
    87: op1_10_in28 = reg_0184;
    76: op1_10_in28 = reg_0584;
    61: op1_10_in28 = reg_1140;
    57: op1_10_in28 = reg_0031;
    77: op1_10_in28 = reg_0607;
    58: op1_10_in28 = reg_0154;
    78: op1_10_in28 = reg_0102;
    70: op1_10_in28 = reg_0150;
    79: op1_10_in28 = reg_0569;
    59: op1_10_in28 = reg_1036;
    60: op1_10_in28 = reg_0963;
    88: op1_10_in28 = reg_0735;
    46: op1_10_in28 = reg_0302;
    80: op1_10_in28 = reg_0238;
    81: op1_10_in28 = imem06_in[7:4];
    82: op1_10_in28 = reg_0591;
    89: op1_10_in28 = reg_0369;
    83: op1_10_in28 = reg_0968;
    64: op1_10_in28 = reg_0884;
    84: op1_10_in28 = reg_0220;
    48: op1_10_in28 = reg_0851;
    85: op1_10_in28 = reg_0979;
    90: op1_10_in28 = reg_0399;
    66: op1_10_in28 = reg_0934;
    67: op1_10_in28 = reg_0043;
    92: op1_10_in28 = reg_0332;
    93: op1_10_in28 = reg_0347;
    94: op1_10_in28 = imem03_in[11:8];
    95: op1_10_in28 = reg_0438;
    96: op1_10_in28 = reg_0443;
    97: op1_10_in28 = reg_0350;
    98: op1_10_in28 = reg_0316;
    100: op1_10_in28 = reg_0558;
    101: op1_10_in28 = reg_0742;
    102: op1_10_in28 = reg_0065;
    103: op1_10_in28 = reg_0195;
    47: op1_10_in28 = reg_0867;
    106: op1_10_in28 = reg_0965;
    44: op1_10_in28 = reg_0460;
    107: op1_10_in28 = reg_1139;
    108: op1_10_in28 = imem07_in[15:12];
    109: op1_10_in28 = reg_0374;
    124: op1_10_in28 = reg_0374;
    110: op1_10_in28 = reg_1033;
    111: op1_10_in28 = reg_0225;
    112: op1_10_in28 = reg_0149;
    113: op1_10_in28 = reg_0620;
    114: op1_10_in28 = reg_1040;
    115: op1_10_in28 = reg_0457;
    116: op1_10_in28 = reg_0319;
    118: op1_10_in28 = reg_0080;
    119: op1_10_in28 = reg_1300;
    120: op1_10_in28 = reg_1518;
    121: op1_10_in28 = reg_1402;
    122: op1_10_in28 = reg_1383;
    123: op1_10_in28 = reg_1094;
    125: op1_10_in28 = reg_0362;
    130: op1_10_in28 = reg_0362;
    126: op1_10_in28 = reg_0094;
    127: op1_10_in28 = reg_0559;
    128: op1_10_in28 = reg_0531;
    129: op1_10_in28 = reg_0391;
    42: op1_10_in28 = reg_0666;
    131: op1_10_in28 = reg_0793;
    default: op1_10_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_10_inv28 = 1;
    73: op1_10_inv28 = 1;
    54: op1_10_inv28 = 1;
    68: op1_10_inv28 = 1;
    50: op1_10_inv28 = 1;
    56: op1_10_inv28 = 1;
    87: op1_10_inv28 = 1;
    76: op1_10_inv28 = 1;
    77: op1_10_inv28 = 1;
    78: op1_10_inv28 = 1;
    88: op1_10_inv28 = 1;
    80: op1_10_inv28 = 1;
    82: op1_10_inv28 = 1;
    83: op1_10_inv28 = 1;
    64: op1_10_inv28 = 1;
    84: op1_10_inv28 = 1;
    48: op1_10_inv28 = 1;
    85: op1_10_inv28 = 1;
    66: op1_10_inv28 = 1;
    67: op1_10_inv28 = 1;
    93: op1_10_inv28 = 1;
    103: op1_10_inv28 = 1;
    47: op1_10_inv28 = 1;
    44: op1_10_inv28 = 1;
    107: op1_10_inv28 = 1;
    109: op1_10_inv28 = 1;
    110: op1_10_inv28 = 1;
    112: op1_10_inv28 = 1;
    113: op1_10_inv28 = 1;
    118: op1_10_inv28 = 1;
    121: op1_10_inv28 = 1;
    122: op1_10_inv28 = 1;
    123: op1_10_inv28 = 1;
    128: op1_10_inv28 = 1;
    42: op1_10_inv28 = 1;
    131: op1_10_inv28 = 1;
    default: op1_10_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in29 = reg_0827;
    53: op1_10_in29 = reg_0450;
    86: op1_10_in29 = reg_1339;
    55: op1_10_in29 = reg_0300;
    46: op1_10_in29 = reg_0300;
    73: op1_10_in29 = reg_0667;
    42: op1_10_in29 = reg_0667;
    69: op1_10_in29 = reg_0598;
    74: op1_10_in29 = reg_0052;
    54: op1_10_in29 = reg_0527;
    68: op1_10_in29 = reg_0020;
    75: op1_10_in29 = reg_0742;
    80: op1_10_in29 = reg_0742;
    50: op1_10_in29 = reg_0106;
    56: op1_10_in29 = reg_0014;
    71: op1_10_in29 = reg_0257;
    87: op1_10_in29 = reg_0395;
    92: op1_10_in29 = reg_0395;
    76: op1_10_in29 = reg_0624;
    61: op1_10_in29 = reg_0399;
    57: op1_10_in29 = reg_0663;
    77: op1_10_in29 = reg_0530;
    58: op1_10_in29 = reg_0829;
    78: op1_10_in29 = reg_0321;
    70: op1_10_in29 = reg_0034;
    79: op1_10_in29 = reg_0979;
    59: op1_10_in29 = reg_0751;
    60: op1_10_in29 = imem03_in[3:0];
    88: op1_10_in29 = reg_1431;
    81: op1_10_in29 = reg_0120;
    82: op1_10_in29 = reg_0592;
    89: op1_10_in29 = reg_1237;
    83: op1_10_in29 = reg_0438;
    64: op1_10_in29 = reg_0481;
    84: op1_10_in29 = reg_0246;
    48: op1_10_in29 = reg_0674;
    85: op1_10_in29 = reg_0244;
    90: op1_10_in29 = reg_0456;
    66: op1_10_in29 = reg_0128;
    91: op1_10_in29 = reg_0412;
    67: op1_10_in29 = reg_0044;
    93: op1_10_in29 = reg_0205;
    94: op1_10_in29 = reg_0999;
    95: op1_10_in29 = reg_0149;
    96: op1_10_in29 = reg_0252;
    97: op1_10_in29 = reg_0313;
    98: op1_10_in29 = reg_0696;
    100: op1_10_in29 = reg_0885;
    101: op1_10_in29 = reg_0968;
    102: op1_10_in29 = reg_0490;
    103: op1_10_in29 = reg_0396;
    47: op1_10_in29 = reg_0791;
    106: op1_10_in29 = reg_1518;
    44: op1_10_in29 = reg_0268;
    107: op1_10_in29 = reg_1325;
    108: op1_10_in29 = reg_0226;
    109: op1_10_in29 = reg_0141;
    110: op1_10_in29 = reg_0557;
    111: op1_10_in29 = reg_0170;
    112: op1_10_in29 = reg_0595;
    113: op1_10_in29 = reg_0137;
    114: op1_10_in29 = reg_0698;
    115: op1_10_in29 = reg_1349;
    116: op1_10_in29 = reg_0577;
    118: op1_10_in29 = reg_0079;
    119: op1_10_in29 = reg_0882;
    120: op1_10_in29 = reg_0957;
    121: op1_10_in29 = reg_0792;
    122: op1_10_in29 = imem04_in[7:4];
    123: op1_10_in29 = reg_0774;
    124: op1_10_in29 = reg_0617;
    125: op1_10_in29 = reg_0092;
    126: op1_10_in29 = reg_0421;
    127: op1_10_in29 = reg_0025;
    128: op1_10_in29 = reg_0500;
    129: op1_10_in29 = reg_0182;
    130: op1_10_in29 = reg_0091;
    131: op1_10_in29 = reg_0392;
    default: op1_10_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv29 = 1;
    86: op1_10_inv29 = 1;
    69: op1_10_inv29 = 1;
    54: op1_10_inv29 = 1;
    75: op1_10_inv29 = 1;
    61: op1_10_inv29 = 1;
    78: op1_10_inv29 = 1;
    79: op1_10_inv29 = 1;
    88: op1_10_inv29 = 1;
    81: op1_10_inv29 = 1;
    48: op1_10_inv29 = 1;
    85: op1_10_inv29 = 1;
    66: op1_10_inv29 = 1;
    91: op1_10_inv29 = 1;
    92: op1_10_inv29 = 1;
    93: op1_10_inv29 = 1;
    100: op1_10_inv29 = 1;
    102: op1_10_inv29 = 1;
    103: op1_10_inv29 = 1;
    106: op1_10_inv29 = 1;
    108: op1_10_inv29 = 1;
    110: op1_10_inv29 = 1;
    114: op1_10_inv29 = 1;
    115: op1_10_inv29 = 1;
    116: op1_10_inv29 = 1;
    121: op1_10_inv29 = 1;
    123: op1_10_inv29 = 1;
    124: op1_10_inv29 = 1;
    126: op1_10_inv29 = 1;
    129: op1_10_inv29 = 1;
    131: op1_10_inv29 = 1;
    default: op1_10_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_10_in30 = reg_0264;
    53: op1_10_in30 = reg_0890;
    86: op1_10_in30 = reg_1338;
    55: op1_10_in30 = reg_0197;
    73: op1_10_in30 = reg_1351;
    69: op1_10_in30 = reg_1419;
    74: op1_10_in30 = reg_0053;
    54: op1_10_in30 = reg_0244;
    68: op1_10_in30 = reg_0799;
    75: op1_10_in30 = reg_0469;
    50: op1_10_in30 = reg_0379;
    56: op1_10_in30 = reg_0120;
    71: op1_10_in30 = reg_0595;
    87: op1_10_in30 = reg_0346;
    76: op1_10_in30 = reg_0569;
    61: op1_10_in30 = reg_0497;
    57: op1_10_in30 = reg_0442;
    77: op1_10_in30 = reg_0138;
    58: op1_10_in30 = reg_0800;
    78: op1_10_in30 = reg_0050;
    70: op1_10_in30 = reg_0136;
    88: op1_10_in30 = reg_0136;
    79: op1_10_in30 = reg_0296;
    59: op1_10_in30 = reg_0906;
    60: op1_10_in30 = reg_0558;
    46: op1_10_in30 = reg_0243;
    80: op1_10_in30 = reg_0966;
    81: op1_10_in30 = reg_1509;
    82: op1_10_in30 = reg_0102;
    89: op1_10_in30 = reg_0932;
    83: op1_10_in30 = reg_0901;
    125: op1_10_in30 = reg_0901;
    64: op1_10_in30 = reg_0443;
    84: op1_10_in30 = reg_1301;
    48: op1_10_in30 = reg_0159;
    85: op1_10_in30 = reg_1204;
    90: op1_10_in30 = reg_0276;
    66: op1_10_in30 = reg_0380;
    91: op1_10_in30 = reg_0969;
    126: op1_10_in30 = reg_0969;
    67: op1_10_in30 = reg_0011;
    92: op1_10_in30 = reg_0996;
    93: op1_10_in30 = reg_1164;
    94: op1_10_in30 = reg_0233;
    95: op1_10_in30 = reg_0403;
    96: op1_10_in30 = imem04_in[3:0];
    97: op1_10_in30 = reg_1144;
    98: op1_10_in30 = reg_0271;
    100: op1_10_in30 = reg_0880;
    101: op1_10_in30 = reg_0148;
    102: op1_10_in30 = reg_0538;
    103: op1_10_in30 = reg_0023;
    47: op1_10_in30 = reg_0030;
    106: op1_10_in30 = reg_0954;
    44: op1_10_in30 = reg_0215;
    107: op1_10_in30 = reg_0493;
    108: op1_10_in30 = reg_0498;
    109: op1_10_in30 = reg_0584;
    110: op1_10_in30 = reg_0783;
    111: op1_10_in30 = reg_0309;
    112: op1_10_in30 = reg_0875;
    113: op1_10_in30 = reg_0592;
    114: op1_10_in30 = reg_0340;
    115: op1_10_in30 = reg_0489;
    116: op1_10_in30 = reg_1369;
    118: op1_10_in30 = reg_0402;
    119: op1_10_in30 = reg_0378;
    120: op1_10_in30 = reg_1231;
    121: op1_10_in30 = reg_0477;
    122: op1_10_in30 = reg_0252;
    123: op1_10_in30 = reg_0664;
    124: op1_10_in30 = reg_0526;
    127: op1_10_in30 = reg_0218;
    128: op1_10_in30 = reg_1214;
    129: op1_10_in30 = reg_0334;
    130: op1_10_in30 = reg_0727;
    42: op1_10_in30 = reg_0608;
    131: op1_10_in30 = reg_0701;
    default: op1_10_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_10_inv30 = 1;
    53: op1_10_inv30 = 1;
    86: op1_10_inv30 = 1;
    55: op1_10_inv30 = 1;
    73: op1_10_inv30 = 1;
    69: op1_10_inv30 = 1;
    68: op1_10_inv30 = 1;
    75: op1_10_inv30 = 1;
    71: op1_10_inv30 = 1;
    87: op1_10_inv30 = 1;
    76: op1_10_inv30 = 1;
    77: op1_10_inv30 = 1;
    58: op1_10_inv30 = 1;
    78: op1_10_inv30 = 1;
    79: op1_10_inv30 = 1;
    59: op1_10_inv30 = 1;
    60: op1_10_inv30 = 1;
    46: op1_10_inv30 = 1;
    81: op1_10_inv30 = 1;
    82: op1_10_inv30 = 1;
    89: op1_10_inv30 = 1;
    83: op1_10_inv30 = 1;
    85: op1_10_inv30 = 1;
    91: op1_10_inv30 = 1;
    67: op1_10_inv30 = 1;
    92: op1_10_inv30 = 1;
    93: op1_10_inv30 = 1;
    94: op1_10_inv30 = 1;
    95: op1_10_inv30 = 1;
    96: op1_10_inv30 = 1;
    100: op1_10_inv30 = 1;
    101: op1_10_inv30 = 1;
    47: op1_10_inv30 = 1;
    106: op1_10_inv30 = 1;
    44: op1_10_inv30 = 1;
    107: op1_10_inv30 = 1;
    109: op1_10_inv30 = 1;
    110: op1_10_inv30 = 1;
    111: op1_10_inv30 = 1;
    112: op1_10_inv30 = 1;
    118: op1_10_inv30 = 1;
    120: op1_10_inv30 = 1;
    122: op1_10_inv30 = 1;
    125: op1_10_inv30 = 1;
    127: op1_10_inv30 = 1;
    131: op1_10_inv30 = 1;
    default: op1_10_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_10_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#10の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_10_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in00 = reg_0554;
    53: op1_11_in00 = reg_0468;
    55: op1_11_in00 = reg_0962;
    73: op1_11_in00 = reg_0320;
    86: op1_11_in00 = reg_0143;
    74: op1_11_in00 = reg_0615;
    69: op1_11_in00 = reg_0377;
    49: op1_11_in00 = reg_0157;
    54: op1_11_in00 = reg_0091;
    75: op1_11_in00 = reg_1419;
    50: op1_11_in00 = reg_0890;
    56: op1_11_in00 = reg_1183;
    68: op1_11_in00 = reg_0708;
    76: op1_11_in00 = reg_0088;
    71: op1_11_in00 = reg_0219;
    59: op1_11_in00 = reg_0219;
    85: op1_11_in00 = reg_0219;
    87: op1_11_in00 = reg_1367;
    57: op1_11_in00 = reg_0137;
    77: op1_11_in00 = imem05_in[15:12];
    61: op1_11_in00 = reg_0445;
    62: op1_11_in00 = reg_0445;
    58: op1_11_in00 = reg_0797;
    44: op1_11_in00 = reg_0797;
    78: op1_11_in00 = reg_1281;
    70: op1_11_in00 = reg_0360;
    79: op1_11_in00 = imem00_in[11:8];
    81: op1_11_in00 = imem00_in[11:8];
    51: op1_11_in00 = reg_0869;
    60: op1_11_in00 = reg_0119;
    88: op1_11_in00 = reg_0734;
    80: op1_11_in00 = reg_0710;
    46: op1_11_in00 = reg_0932;
    52: op1_11_in00 = reg_0899;
    63: op1_11_in00 = reg_0078;
    82: op1_11_in00 = reg_0121;
    89: op1_11_in00 = reg_0000;
    47: op1_11_in00 = reg_0000;
    83: op1_11_in00 = reg_0350;
    84: op1_11_in00 = reg_0350;
    64: op1_11_in00 = reg_0698;
    33: op1_11_in00 = reg_0286;
    38: op1_11_in00 = reg_0286;
    48: op1_11_in00 = reg_0743;
    65: op1_11_in00 = reg_0743;
    90: op1_11_in00 = imem04_in[3:0];
    66: op1_11_in00 = reg_0462;
    91: op1_11_in00 = imem00_in[3:0];
    111: op1_11_in00 = imem00_in[3:0];
    28: op1_11_in00 = reg_0002;
    67: op1_11_in00 = reg_0013;
    92: op1_11_in00 = reg_0176;
    93: op1_11_in00 = reg_0700;
    94: op1_11_in00 = reg_0759;
    95: op1_11_in00 = reg_0363;
    96: op1_11_in00 = reg_0577;
    97: op1_11_in00 = imem04_in[7:4];
    98: op1_11_in00 = reg_0984;
    37: op1_11_in00 = imem07_in[11:8];
    99: op1_11_in00 = imem00_in[7:4];
    105: op1_11_in00 = imem00_in[7:4];
    117: op1_11_in00 = imem00_in[7:4];
    100: op1_11_in00 = reg_0025;
    101: op1_11_in00 = reg_0290;
    102: op1_11_in00 = reg_1104;
    103: op1_11_in00 = reg_0994;
    104: op1_11_in00 = reg_1277;
    106: op1_11_in00 = reg_0178;
    120: op1_11_in00 = reg_0178;
    107: op1_11_in00 = reg_0275;
    108: op1_11_in00 = reg_0725;
    109: op1_11_in00 = reg_0617;
    110: op1_11_in00 = reg_0191;
    112: op1_11_in00 = reg_0077;
    113: op1_11_in00 = reg_0638;
    114: op1_11_in00 = reg_0236;
    115: op1_11_in00 = reg_0926;
    116: op1_11_in00 = reg_1203;
    118: op1_11_in00 = reg_0728;
    119: op1_11_in00 = reg_1009;
    121: op1_11_in00 = reg_0937;
    122: op1_11_in00 = reg_1216;
    123: op1_11_in00 = reg_1244;
    124: op1_11_in00 = reg_0295;
    125: op1_11_in00 = reg_0595;
    34: op1_11_in00 = reg_0156;
    126: op1_11_in00 = reg_0931;
    127: op1_11_in00 = reg_1280;
    128: op1_11_in00 = reg_0414;
    129: op1_11_in00 = reg_1180;
    130: op1_11_in00 = reg_0292;
    131: op1_11_in00 = reg_0045;
    default: op1_11_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv00 = 1;
    86: op1_11_inv00 = 1;
    74: op1_11_inv00 = 1;
    69: op1_11_inv00 = 1;
    54: op1_11_inv00 = 1;
    50: op1_11_inv00 = 1;
    56: op1_11_inv00 = 1;
    68: op1_11_inv00 = 1;
    76: op1_11_inv00 = 1;
    87: op1_11_inv00 = 1;
    77: op1_11_inv00 = 1;
    61: op1_11_inv00 = 1;
    58: op1_11_inv00 = 1;
    78: op1_11_inv00 = 1;
    70: op1_11_inv00 = 1;
    51: op1_11_inv00 = 1;
    88: op1_11_inv00 = 1;
    81: op1_11_inv00 = 1;
    46: op1_11_inv00 = 1;
    52: op1_11_inv00 = 1;
    64: op1_11_inv00 = 1;
    33: op1_11_inv00 = 1;
    84: op1_11_inv00 = 1;
    85: op1_11_inv00 = 1;
    90: op1_11_inv00 = 1;
    66: op1_11_inv00 = 1;
    91: op1_11_inv00 = 1;
    67: op1_11_inv00 = 1;
    92: op1_11_inv00 = 1;
    94: op1_11_inv00 = 1;
    97: op1_11_inv00 = 1;
    98: op1_11_inv00 = 1;
    99: op1_11_inv00 = 1;
    101: op1_11_inv00 = 1;
    102: op1_11_inv00 = 1;
    104: op1_11_inv00 = 1;
    105: op1_11_inv00 = 1;
    106: op1_11_inv00 = 1;
    47: op1_11_inv00 = 1;
    107: op1_11_inv00 = 1;
    109: op1_11_inv00 = 1;
    111: op1_11_inv00 = 1;
    113: op1_11_inv00 = 1;
    114: op1_11_inv00 = 1;
    115: op1_11_inv00 = 1;
    116: op1_11_inv00 = 1;
    117: op1_11_inv00 = 1;
    120: op1_11_inv00 = 1;
    122: op1_11_inv00 = 1;
    44: op1_11_inv00 = 1;
    34: op1_11_inv00 = 1;
    128: op1_11_inv00 = 1;
    38: op1_11_inv00 = 1;
    130: op1_11_inv00 = 1;
    131: op1_11_inv00 = 1;
    default: op1_11_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in01 = reg_0616;
    53: op1_11_in01 = reg_0966;
    55: op1_11_in01 = reg_0145;
    110: op1_11_in01 = reg_0145;
    73: op1_11_in01 = reg_1151;
    86: op1_11_in01 = reg_0789;
    74: op1_11_in01 = reg_0614;
    59: op1_11_in01 = reg_0614;
    105: op1_11_in01 = reg_0614;
    69: op1_11_in01 = reg_0709;
    49: op1_11_in01 = imem07_in[11:8];
    54: op1_11_in01 = reg_0899;
    75: op1_11_in01 = reg_0698;
    50: op1_11_in01 = reg_0888;
    56: op1_11_in01 = reg_0223;
    68: op1_11_in01 = reg_0306;
    76: op1_11_in01 = reg_0590;
    71: op1_11_in01 = reg_0748;
    87: op1_11_in01 = reg_0493;
    57: op1_11_in01 = reg_0102;
    77: op1_11_in01 = reg_0450;
    61: op1_11_in01 = reg_1081;
    58: op1_11_in01 = reg_0795;
    126: op1_11_in01 = reg_0795;
    78: op1_11_in01 = reg_1277;
    70: op1_11_in01 = reg_0896;
    79: op1_11_in01 = reg_0983;
    83: op1_11_in01 = reg_0983;
    51: op1_11_in01 = reg_0870;
    60: op1_11_in01 = reg_0271;
    88: op1_11_in01 = imem02_in[7:4];
    80: op1_11_in01 = reg_0049;
    62: op1_11_in01 = reg_0669;
    81: op1_11_in01 = reg_0907;
    46: op1_11_in01 = reg_0452;
    52: op1_11_in01 = reg_0283;
    63: op1_11_in01 = reg_0290;
    82: op1_11_in01 = reg_1281;
    89: op1_11_in01 = reg_0375;
    64: op1_11_in01 = reg_0595;
    33: op1_11_in01 = reg_0441;
    84: op1_11_in01 = reg_0554;
    48: op1_11_in01 = reg_0468;
    85: op1_11_in01 = imem00_in[7:4];
    65: op1_11_in01 = reg_0161;
    90: op1_11_in01 = reg_0032;
    66: op1_11_in01 = reg_1203;
    91: op1_11_in01 = imem00_in[11:8];
    111: op1_11_in01 = imem00_in[11:8];
    117: op1_11_in01 = imem00_in[11:8];
    28: op1_11_in01 = reg_0085;
    67: op1_11_in01 = reg_1103;
    92: op1_11_in01 = reg_0174;
    93: op1_11_in01 = reg_0176;
    94: op1_11_in01 = reg_1447;
    95: op1_11_in01 = reg_0464;
    96: op1_11_in01 = reg_1383;
    97: op1_11_in01 = reg_0577;
    98: op1_11_in01 = reg_0827;
    37: op1_11_in01 = reg_0404;
    99: op1_11_in01 = reg_0866;
    100: op1_11_in01 = reg_1325;
    101: op1_11_in01 = reg_0362;
    102: op1_11_in01 = reg_0167;
    103: op1_11_in01 = reg_1055;
    104: op1_11_in01 = reg_1099;
    106: op1_11_in01 = reg_1208;
    120: op1_11_in01 = reg_1208;
    47: op1_11_in01 = reg_0329;
    107: op1_11_in01 = reg_0118;
    108: op1_11_in01 = reg_1101;
    113: op1_11_in01 = reg_1101;
    123: op1_11_in01 = reg_1101;
    109: op1_11_in01 = reg_0529;
    112: op1_11_in01 = reg_0257;
    114: op1_11_in01 = reg_0117;
    115: op1_11_in01 = imem00_in[15:12];
    116: op1_11_in01 = reg_0574;
    118: op1_11_in01 = reg_0010;
    119: op1_11_in01 = reg_0313;
    121: op1_11_in01 = reg_0418;
    122: op1_11_in01 = reg_1367;
    124: op1_11_in01 = reg_0119;
    125: op1_11_in01 = reg_0727;
    44: op1_11_in01 = imem04_in[3:0];
    34: op1_11_in01 = reg_0157;
    127: op1_11_in01 = reg_0699;
    128: op1_11_in01 = reg_0412;
    38: op1_11_in01 = reg_0741;
    129: op1_11_in01 = reg_1163;
    130: op1_11_in01 = reg_0077;
    131: op1_11_in01 = reg_0564;
    default: op1_11_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv01 = 1;
    55: op1_11_inv01 = 1;
    74: op1_11_inv01 = 1;
    49: op1_11_inv01 = 1;
    54: op1_11_inv01 = 1;
    75: op1_11_inv01 = 1;
    87: op1_11_inv01 = 1;
    57: op1_11_inv01 = 1;
    58: op1_11_inv01 = 1;
    78: op1_11_inv01 = 1;
    70: op1_11_inv01 = 1;
    79: op1_11_inv01 = 1;
    51: op1_11_inv01 = 1;
    59: op1_11_inv01 = 1;
    60: op1_11_inv01 = 1;
    80: op1_11_inv01 = 1;
    62: op1_11_inv01 = 1;
    81: op1_11_inv01 = 1;
    46: op1_11_inv01 = 1;
    52: op1_11_inv01 = 1;
    82: op1_11_inv01 = 1;
    64: op1_11_inv01 = 1;
    48: op1_11_inv01 = 1;
    85: op1_11_inv01 = 1;
    90: op1_11_inv01 = 1;
    28: op1_11_inv01 = 1;
    95: op1_11_inv01 = 1;
    96: op1_11_inv01 = 1;
    97: op1_11_inv01 = 1;
    99: op1_11_inv01 = 1;
    102: op1_11_inv01 = 1;
    109: op1_11_inv01 = 1;
    110: op1_11_inv01 = 1;
    111: op1_11_inv01 = 1;
    112: op1_11_inv01 = 1;
    113: op1_11_inv01 = 1;
    115: op1_11_inv01 = 1;
    117: op1_11_inv01 = 1;
    119: op1_11_inv01 = 1;
    120: op1_11_inv01 = 1;
    121: op1_11_inv01 = 1;
    124: op1_11_inv01 = 1;
    34: op1_11_inv01 = 1;
    126: op1_11_inv01 = 1;
    131: op1_11_inv01 = 1;
    default: op1_11_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in02 = reg_0748;
    53: op1_11_in02 = reg_0147;
    55: op1_11_in02 = reg_0142;
    73: op1_11_in02 = reg_0537;
    64: op1_11_in02 = reg_0537;
    86: op1_11_in02 = reg_0965;
    74: op1_11_in02 = reg_0445;
    69: op1_11_in02 = reg_1063;
    49: op1_11_in02 = reg_0169;
    54: op1_11_in02 = reg_0283;
    75: op1_11_in02 = reg_0582;
    50: op1_11_in02 = reg_0300;
    56: op1_11_in02 = reg_0245;
    68: op1_11_in02 = reg_0379;
    76: op1_11_in02 = reg_1103;
    71: op1_11_in02 = reg_0701;
    87: op1_11_in02 = reg_0034;
    97: op1_11_in02 = reg_0034;
    57: op1_11_in02 = reg_0228;
    77: op1_11_in02 = reg_0872;
    61: op1_11_in02 = reg_1241;
    58: op1_11_in02 = reg_0454;
    78: op1_11_in02 = reg_1081;
    70: op1_11_in02 = reg_0079;
    79: op1_11_in02 = reg_1489;
    51: op1_11_in02 = reg_0860;
    59: op1_11_in02 = reg_1099;
    60: op1_11_in02 = reg_0214;
    88: op1_11_in02 = reg_0607;
    80: op1_11_in02 = reg_1001;
    62: op1_11_in02 = reg_0842;
    81: op1_11_in02 = reg_0640;
    46: op1_11_in02 = reg_0904;
    52: op1_11_in02 = reg_0043;
    63: op1_11_in02 = reg_0278;
    82: op1_11_in02 = reg_1278;
    89: op1_11_in02 = reg_1518;
    83: op1_11_in02 = reg_1490;
    33: op1_11_in02 = reg_0408;
    38: op1_11_in02 = reg_0408;
    84: op1_11_in02 = reg_1471;
    48: op1_11_in02 = reg_0728;
    112: op1_11_in02 = reg_0728;
    85: op1_11_in02 = reg_1277;
    65: op1_11_in02 = reg_0982;
    90: op1_11_in02 = reg_1338;
    66: op1_11_in02 = reg_1200;
    91: op1_11_in02 = reg_0725;
    28: op1_11_in02 = reg_0086;
    67: op1_11_in02 = reg_0455;
    92: op1_11_in02 = reg_0392;
    93: op1_11_in02 = reg_0831;
    94: op1_11_in02 = reg_0049;
    95: op1_11_in02 = reg_0335;
    96: op1_11_in02 = reg_1372;
    98: op1_11_in02 = reg_1504;
    37: op1_11_in02 = reg_0618;
    99: op1_11_in02 = reg_1491;
    100: op1_11_in02 = reg_0181;
    101: op1_11_in02 = reg_0175;
    102: op1_11_in02 = reg_0131;
    131: op1_11_in02 = reg_0131;
    103: op1_11_in02 = reg_0478;
    104: op1_11_in02 = reg_1487;
    105: op1_11_in02 = reg_0638;
    106: op1_11_in02 = reg_0104;
    120: op1_11_in02 = reg_0104;
    47: op1_11_in02 = reg_0577;
    107: op1_11_in02 = reg_0603;
    108: op1_11_in02 = reg_0803;
    109: op1_11_in02 = reg_1225;
    110: op1_11_in02 = reg_0143;
    111: op1_11_in02 = imem00_in[15:12];
    113: op1_11_in02 = reg_0805;
    114: op1_11_in02 = reg_1503;
    115: op1_11_in02 = reg_0843;
    116: op1_11_in02 = reg_1233;
    117: op1_11_in02 = reg_0248;
    118: op1_11_in02 = reg_0662;
    119: op1_11_in02 = reg_0348;
    121: op1_11_in02 = reg_0736;
    122: op1_11_in02 = reg_1258;
    123: op1_11_in02 = reg_0958;
    124: op1_11_in02 = reg_0583;
    125: op1_11_in02 = reg_0077;
    44: op1_11_in02 = reg_0369;
    34: op1_11_in02 = reg_0031;
    126: op1_11_in02 = reg_0908;
    127: op1_11_in02 = reg_0164;
    128: op1_11_in02 = reg_0406;
    129: op1_11_in02 = reg_0937;
    130: op1_11_in02 = reg_0042;
    default: op1_11_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv02 = 1;
    74: op1_11_inv02 = 1;
    69: op1_11_inv02 = 1;
    49: op1_11_inv02 = 1;
    54: op1_11_inv02 = 1;
    75: op1_11_inv02 = 1;
    50: op1_11_inv02 = 1;
    56: op1_11_inv02 = 1;
    68: op1_11_inv02 = 1;
    71: op1_11_inv02 = 1;
    57: op1_11_inv02 = 1;
    77: op1_11_inv02 = 1;
    58: op1_11_inv02 = 1;
    78: op1_11_inv02 = 1;
    70: op1_11_inv02 = 1;
    79: op1_11_inv02 = 1;
    88: op1_11_inv02 = 1;
    81: op1_11_inv02 = 1;
    46: op1_11_inv02 = 1;
    63: op1_11_inv02 = 1;
    82: op1_11_inv02 = 1;
    83: op1_11_inv02 = 1;
    33: op1_11_inv02 = 1;
    84: op1_11_inv02 = 1;
    48: op1_11_inv02 = 1;
    66: op1_11_inv02 = 1;
    91: op1_11_inv02 = 1;
    28: op1_11_inv02 = 1;
    67: op1_11_inv02 = 1;
    94: op1_11_inv02 = 1;
    97: op1_11_inv02 = 1;
    98: op1_11_inv02 = 1;
    99: op1_11_inv02 = 1;
    100: op1_11_inv02 = 1;
    101: op1_11_inv02 = 1;
    106: op1_11_inv02 = 1;
    47: op1_11_inv02 = 1;
    107: op1_11_inv02 = 1;
    110: op1_11_inv02 = 1;
    111: op1_11_inv02 = 1;
    113: op1_11_inv02 = 1;
    114: op1_11_inv02 = 1;
    115: op1_11_inv02 = 1;
    116: op1_11_inv02 = 1;
    117: op1_11_inv02 = 1;
    118: op1_11_inv02 = 1;
    119: op1_11_inv02 = 1;
    121: op1_11_inv02 = 1;
    122: op1_11_inv02 = 1;
    123: op1_11_inv02 = 1;
    125: op1_11_inv02 = 1;
    34: op1_11_inv02 = 1;
    127: op1_11_inv02 = 1;
    128: op1_11_inv02 = 1;
    38: op1_11_inv02 = 1;
    default: op1_11_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in03 = reg_0824;
    53: op1_11_in03 = reg_0402;
    55: op1_11_in03 = reg_0952;
    73: op1_11_in03 = reg_0582;
    86: op1_11_in03 = reg_0964;
    74: op1_11_in03 = imem00_in[7:4];
    69: op1_11_in03 = imem03_in[7:4];
    49: op1_11_in03 = reg_0777;
    54: op1_11_in03 = reg_0629;
    75: op1_11_in03 = reg_0862;
    50: op1_11_in03 = reg_0872;
    56: op1_11_in03 = reg_0298;
    68: op1_11_in03 = reg_0897;
    76: op1_11_in03 = reg_0055;
    71: op1_11_in03 = reg_0445;
    87: op1_11_in03 = reg_0462;
    90: op1_11_in03 = reg_0462;
    57: op1_11_in03 = reg_0050;
    28: op1_11_in03 = reg_0050;
    77: op1_11_in03 = reg_1484;
    61: op1_11_in03 = reg_0293;
    58: op1_11_in03 = reg_0368;
    46: op1_11_in03 = reg_0368;
    78: op1_11_in03 = reg_1489;
    70: op1_11_in03 = reg_0282;
    79: op1_11_in03 = reg_1491;
    51: op1_11_in03 = reg_0720;
    59: op1_11_in03 = imem00_in[15:12];
    60: op1_11_in03 = reg_1056;
    88: op1_11_in03 = reg_0588;
    80: op1_11_in03 = reg_0823;
    62: op1_11_in03 = reg_1243;
    81: op1_11_in03 = reg_1281;
    52: op1_11_in03 = reg_0010;
    63: op1_11_in03 = reg_0042;
    82: op1_11_in03 = imem00_in[3:0];
    89: op1_11_in03 = reg_0954;
    83: op1_11_in03 = reg_1242;
    64: op1_11_in03 = reg_0978;
    122: op1_11_in03 = reg_0978;
    33: op1_11_in03 = imem07_in[11:8];
    84: op1_11_in03 = reg_1027;
    48: op1_11_in03 = reg_0726;
    85: op1_11_in03 = reg_1279;
    65: op1_11_in03 = reg_0468;
    66: op1_11_in03 = reg_1065;
    91: op1_11_in03 = reg_0791;
    67: op1_11_in03 = reg_0590;
    92: op1_11_in03 = reg_0562;
    93: op1_11_in03 = reg_0649;
    94: op1_11_in03 = reg_0198;
    95: op1_11_in03 = reg_0077;
    96: op1_11_in03 = reg_0493;
    97: op1_11_in03 = reg_1082;
    116: op1_11_in03 = reg_1082;
    98: op1_11_in03 = reg_0716;
    37: op1_11_in03 = reg_0620;
    99: op1_11_in03 = reg_0804;
    100: op1_11_in03 = reg_0731;
    101: op1_11_in03 = reg_0875;
    102: op1_11_in03 = reg_1404;
    103: op1_11_in03 = reg_1060;
    104: op1_11_in03 = reg_0803;
    105: op1_11_in03 = reg_0186;
    106: op1_11_in03 = reg_0025;
    47: op1_11_in03 = reg_0694;
    107: op1_11_in03 = reg_0931;
    108: op1_11_in03 = reg_0580;
    109: op1_11_in03 = reg_0132;
    110: op1_11_in03 = reg_1516;
    111: op1_11_in03 = reg_0248;
    112: op1_11_in03 = imem02_in[3:0];
    113: op1_11_in03 = reg_0523;
    114: op1_11_in03 = reg_0470;
    44: op1_11_in03 = reg_0470;
    115: op1_11_in03 = reg_1141;
    117: op1_11_in03 = reg_1081;
    118: op1_11_in03 = reg_0456;
    119: op1_11_in03 = reg_0426;
    120: op1_11_in03 = reg_0882;
    121: op1_11_in03 = reg_0794;
    123: op1_11_in03 = reg_0907;
    124: op1_11_in03 = reg_0754;
    125: op1_11_in03 = reg_0724;
    34: op1_11_in03 = reg_0029;
    126: op1_11_in03 = reg_0826;
    127: op1_11_in03 = reg_0236;
    128: op1_11_in03 = reg_1041;
    38: op1_11_in03 = reg_0415;
    129: op1_11_in03 = reg_0066;
    130: op1_11_in03 = reg_0166;
    131: op1_11_in03 = reg_0697;
    default: op1_11_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv03 = 1;
    55: op1_11_inv03 = 1;
    73: op1_11_inv03 = 1;
    50: op1_11_inv03 = 1;
    68: op1_11_inv03 = 1;
    76: op1_11_inv03 = 1;
    71: op1_11_inv03 = 1;
    57: op1_11_inv03 = 1;
    77: op1_11_inv03 = 1;
    61: op1_11_inv03 = 1;
    60: op1_11_inv03 = 1;
    88: op1_11_inv03 = 1;
    62: op1_11_inv03 = 1;
    52: op1_11_inv03 = 1;
    63: op1_11_inv03 = 1;
    82: op1_11_inv03 = 1;
    84: op1_11_inv03 = 1;
    90: op1_11_inv03 = 1;
    91: op1_11_inv03 = 1;
    28: op1_11_inv03 = 1;
    67: op1_11_inv03 = 1;
    96: op1_11_inv03 = 1;
    97: op1_11_inv03 = 1;
    37: op1_11_inv03 = 1;
    102: op1_11_inv03 = 1;
    106: op1_11_inv03 = 1;
    47: op1_11_inv03 = 1;
    111: op1_11_inv03 = 1;
    112: op1_11_inv03 = 1;
    114: op1_11_inv03 = 1;
    120: op1_11_inv03 = 1;
    124: op1_11_inv03 = 1;
    44: op1_11_inv03 = 1;
    127: op1_11_inv03 = 1;
    38: op1_11_inv03 = 1;
    131: op1_11_inv03 = 1;
    default: op1_11_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in04 = reg_1277;
    53: op1_11_in04 = reg_0384;
    55: op1_11_in04 = reg_0190;
    73: op1_11_in04 = reg_0719;
    46: op1_11_in04 = reg_0719;
    86: op1_11_in04 = reg_0314;
    74: op1_11_in04 = imem00_in[11:8];
    69: op1_11_in04 = imem03_in[11:8];
    49: op1_11_in04 = reg_0664;
    54: op1_11_in04 = reg_1098;
    75: op1_11_in04 = reg_0338;
    50: op1_11_in04 = reg_0184;
    56: op1_11_in04 = reg_0777;
    68: op1_11_in04 = reg_0007;
    76: op1_11_in04 = reg_1260;
    71: op1_11_in04 = reg_0824;
    87: op1_11_in04 = reg_0531;
    57: op1_11_in04 = reg_1182;
    77: op1_11_in04 = reg_0274;
    129: op1_11_in04 = reg_0274;
    61: op1_11_in04 = reg_0136;
    58: op1_11_in04 = reg_0862;
    78: op1_11_in04 = imem00_in[3:0];
    70: op1_11_in04 = reg_0446;
    79: op1_11_in04 = reg_1243;
    81: op1_11_in04 = reg_1243;
    51: op1_11_in04 = reg_0859;
    59: op1_11_in04 = reg_0843;
    60: op1_11_in04 = reg_0994;
    88: op1_11_in04 = reg_0934;
    80: op1_11_in04 = reg_0962;
    62: op1_11_in04 = reg_1244;
    82: op1_11_in04 = reg_1244;
    52: op1_11_in04 = reg_0133;
    63: op1_11_in04 = reg_0044;
    89: op1_11_in04 = reg_0952;
    83: op1_11_in04 = reg_0615;
    64: op1_11_in04 = reg_0462;
    33: op1_11_in04 = imem07_in[15:12];
    84: op1_11_in04 = reg_0221;
    48: op1_11_in04 = reg_0146;
    85: op1_11_in04 = reg_1079;
    65: op1_11_in04 = reg_0438;
    90: op1_11_in04 = reg_0574;
    66: op1_11_in04 = reg_1147;
    91: op1_11_in04 = reg_0866;
    28: op1_11_in04 = imem07_in[7:4];
    67: op1_11_in04 = reg_0981;
    92: op1_11_in04 = reg_0701;
    93: op1_11_in04 = reg_0562;
    94: op1_11_in04 = reg_0311;
    95: op1_11_in04 = reg_0724;
    96: op1_11_in04 = reg_0264;
    97: op1_11_in04 = reg_0412;
    98: op1_11_in04 = reg_0714;
    37: op1_11_in04 = reg_0591;
    99: op1_11_in04 = reg_0613;
    104: op1_11_in04 = reg_0613;
    100: op1_11_in04 = reg_0797;
    101: op1_11_in04 = reg_0464;
    102: op1_11_in04 = reg_0940;
    103: op1_11_in04 = reg_0667;
    105: op1_11_in04 = reg_0523;
    106: op1_11_in04 = imem04_in[7:4];
    47: op1_11_in04 = reg_0537;
    107: op1_11_in04 = reg_0192;
    108: op1_11_in04 = reg_1028;
    109: op1_11_in04 = reg_0295;
    110: op1_11_in04 = reg_0954;
    111: op1_11_in04 = reg_0672;
    112: op1_11_in04 = reg_0456;
    113: op1_11_in04 = reg_0293;
    114: op1_11_in04 = reg_0466;
    115: op1_11_in04 = reg_0486;
    116: op1_11_in04 = reg_0320;
    117: op1_11_in04 = reg_0725;
    118: op1_11_in04 = reg_0721;
    119: op1_11_in04 = imem04_in[3:0];
    120: op1_11_in04 = reg_0884;
    121: op1_11_in04 = reg_0492;
    122: op1_11_in04 = reg_1203;
    123: op1_11_in04 = reg_0153;
    124: op1_11_in04 = reg_1170;
    125: op1_11_in04 = reg_0041;
    44: op1_11_in04 = reg_0341;
    34: op1_11_in04 = reg_0030;
    126: op1_11_in04 = reg_0161;
    127: op1_11_in04 = reg_0337;
    128: op1_11_in04 = reg_1004;
    38: op1_11_in04 = reg_0321;
    130: op1_11_in04 = reg_0447;
    131: op1_11_in04 = reg_0938;
    default: op1_11_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv04 = 1;
    55: op1_11_inv04 = 1;
    69: op1_11_inv04 = 1;
    54: op1_11_inv04 = 1;
    75: op1_11_inv04 = 1;
    50: op1_11_inv04 = 1;
    56: op1_11_inv04 = 1;
    68: op1_11_inv04 = 1;
    76: op1_11_inv04 = 1;
    87: op1_11_inv04 = 1;
    57: op1_11_inv04 = 1;
    77: op1_11_inv04 = 1;
    70: op1_11_inv04 = 1;
    51: op1_11_inv04 = 1;
    59: op1_11_inv04 = 1;
    81: op1_11_inv04 = 1;
    46: op1_11_inv04 = 1;
    52: op1_11_inv04 = 1;
    89: op1_11_inv04 = 1;
    83: op1_11_inv04 = 1;
    64: op1_11_inv04 = 1;
    84: op1_11_inv04 = 1;
    91: op1_11_inv04 = 1;
    28: op1_11_inv04 = 1;
    67: op1_11_inv04 = 1;
    93: op1_11_inv04 = 1;
    95: op1_11_inv04 = 1;
    98: op1_11_inv04 = 1;
    37: op1_11_inv04 = 1;
    99: op1_11_inv04 = 1;
    100: op1_11_inv04 = 1;
    101: op1_11_inv04 = 1;
    103: op1_11_inv04 = 1;
    106: op1_11_inv04 = 1;
    47: op1_11_inv04 = 1;
    111: op1_11_inv04 = 1;
    112: op1_11_inv04 = 1;
    118: op1_11_inv04 = 1;
    121: op1_11_inv04 = 1;
    123: op1_11_inv04 = 1;
    124: op1_11_inv04 = 1;
    125: op1_11_inv04 = 1;
    44: op1_11_inv04 = 1;
    126: op1_11_inv04 = 1;
    128: op1_11_inv04 = 1;
    default: op1_11_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in05 = reg_1243;
    53: op1_11_in05 = reg_0091;
    55: op1_11_in05 = reg_0246;
    73: op1_11_in05 = reg_0336;
    86: op1_11_in05 = reg_1314;
    74: op1_11_in05 = reg_1078;
    69: op1_11_in05 = reg_1033;
    49: op1_11_in05 = reg_0442;
    56: op1_11_in05 = reg_0442;
    54: op1_11_in05 = reg_1029;
    75: op1_11_in05 = reg_0236;
    50: op1_11_in05 = reg_0130;
    68: op1_11_in05 = reg_0008;
    76: op1_11_in05 = reg_1207;
    71: op1_11_in05 = reg_0672;
    87: op1_11_in05 = reg_0297;
    127: op1_11_in05 = reg_0297;
    77: op1_11_in05 = reg_0243;
    61: op1_11_in05 = reg_1206;
    108: op1_11_in05 = reg_1206;
    58: op1_11_in05 = reg_0164;
    119: op1_11_in05 = reg_0164;
    78: op1_11_in05 = imem00_in[7:4];
    70: op1_11_in05 = reg_0699;
    79: op1_11_in05 = reg_0615;
    51: op1_11_in05 = reg_0374;
    59: op1_11_in05 = reg_0523;
    60: op1_11_in05 = reg_0668;
    88: op1_11_in05 = reg_0561;
    80: op1_11_in05 = reg_0234;
    62: op1_11_in05 = reg_1053;
    81: op1_11_in05 = reg_1244;
    46: op1_11_in05 = reg_0129;
    52: op1_11_in05 = reg_0606;
    63: op1_11_in05 = reg_0012;
    82: op1_11_in05 = reg_1241;
    89: op1_11_in05 = reg_0190;
    83: op1_11_in05 = reg_1470;
    64: op1_11_in05 = reg_1077;
    33: op1_11_in05 = reg_0103;
    84: op1_11_in05 = reg_1230;
    48: op1_11_in05 = reg_0386;
    85: op1_11_in05 = reg_1487;
    65: op1_11_in05 = reg_0148;
    90: op1_11_in05 = reg_0414;
    66: op1_11_in05 = reg_0421;
    91: op1_11_in05 = reg_1490;
    67: op1_11_in05 = reg_0473;
    92: op1_11_in05 = reg_1104;
    93: op1_11_in05 = reg_1180;
    94: op1_11_in05 = reg_0891;
    95: op1_11_in05 = reg_0011;
    96: op1_11_in05 = reg_0462;
    97: op1_11_in05 = reg_0471;
    98: op1_11_in05 = reg_0619;
    37: op1_11_in05 = reg_0137;
    99: op1_11_in05 = reg_0153;
    100: op1_11_in05 = reg_1257;
    101: op1_11_in05 = reg_0634;
    102: op1_11_in05 = reg_0938;
    103: op1_11_in05 = reg_0310;
    104: op1_11_in05 = reg_0616;
    105: op1_11_in05 = reg_0293;
    106: op1_11_in05 = reg_1383;
    47: op1_11_in05 = reg_0464;
    107: op1_11_in05 = reg_0863;
    109: op1_11_in05 = reg_0215;
    110: op1_11_in05 = reg_0952;
    111: op1_11_in05 = reg_1278;
    112: op1_11_in05 = reg_0056;
    113: op1_11_in05 = reg_1227;
    114: op1_11_in05 = reg_0278;
    115: op1_11_in05 = reg_0250;
    123: op1_11_in05 = reg_0250;
    116: op1_11_in05 = reg_1312;
    117: op1_11_in05 = reg_0638;
    118: op1_11_in05 = imem02_in[3:0];
    120: op1_11_in05 = reg_0350;
    121: op1_11_in05 = reg_0393;
    122: op1_11_in05 = reg_1198;
    124: op1_11_in05 = reg_0223;
    125: op1_11_in05 = reg_0895;
    44: op1_11_in05 = reg_0340;
    34: op1_11_in05 = imem07_in[7:4];
    126: op1_11_in05 = reg_0316;
    128: op1_11_in05 = reg_1419;
    38: op1_11_in05 = reg_0051;
    129: op1_11_in05 = reg_1431;
    130: op1_11_in05 = reg_1071;
    131: op1_11_in05 = reg_0589;
    default: op1_11_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    69: op1_11_inv05 = 1;
    54: op1_11_inv05 = 1;
    50: op1_11_inv05 = 1;
    87: op1_11_inv05 = 1;
    58: op1_11_inv05 = 1;
    59: op1_11_inv05 = 1;
    60: op1_11_inv05 = 1;
    88: op1_11_inv05 = 1;
    80: op1_11_inv05 = 1;
    62: op1_11_inv05 = 1;
    81: op1_11_inv05 = 1;
    46: op1_11_inv05 = 1;
    64: op1_11_inv05 = 1;
    84: op1_11_inv05 = 1;
    65: op1_11_inv05 = 1;
    66: op1_11_inv05 = 1;
    67: op1_11_inv05 = 1;
    96: op1_11_inv05 = 1;
    97: op1_11_inv05 = 1;
    102: op1_11_inv05 = 1;
    106: op1_11_inv05 = 1;
    47: op1_11_inv05 = 1;
    107: op1_11_inv05 = 1;
    108: op1_11_inv05 = 1;
    109: op1_11_inv05 = 1;
    111: op1_11_inv05 = 1;
    112: op1_11_inv05 = 1;
    117: op1_11_inv05 = 1;
    120: op1_11_inv05 = 1;
    121: op1_11_inv05 = 1;
    123: op1_11_inv05 = 1;
    44: op1_11_inv05 = 1;
    129: op1_11_inv05 = 1;
    131: op1_11_inv05 = 1;
    default: op1_11_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in06 = reg_1244;
    53: op1_11_in06 = reg_0724;
    55: op1_11_in06 = reg_0889;
    73: op1_11_in06 = reg_0237;
    86: op1_11_in06 = reg_0627;
    74: op1_11_in06 = reg_1489;
    69: op1_11_in06 = reg_0376;
    49: op1_11_in06 = reg_0437;
    54: op1_11_in06 = reg_0456;
    75: op1_11_in06 = imem04_in[3:0];
    50: op1_11_in06 = reg_0274;
    56: op1_11_in06 = reg_0741;
    68: op1_11_in06 = reg_0695;
    76: op1_11_in06 = reg_0429;
    71: op1_11_in06 = reg_0669;
    87: op1_11_in06 = reg_1083;
    100: op1_11_in06 = reg_1083;
    77: op1_11_in06 = reg_0864;
    61: op1_11_in06 = reg_0959;
    58: op1_11_in06 = reg_0211;
    78: op1_11_in06 = reg_0218;
    70: op1_11_in06 = reg_0184;
    79: op1_11_in06 = reg_0580;
    81: op1_11_in06 = reg_0580;
    51: op1_11_in06 = reg_0371;
    59: op1_11_in06 = reg_0250;
    60: op1_11_in06 = reg_0186;
    104: op1_11_in06 = reg_0186;
    88: op1_11_in06 = reg_0532;
    80: op1_11_in06 = reg_0891;
    62: op1_11_in06 = reg_1052;
    46: op1_11_in06 = reg_0019;
    52: op1_11_in06 = reg_1018;
    63: op1_11_in06 = reg_0010;
    82: op1_11_in06 = reg_0613;
    89: op1_11_in06 = reg_0113;
    83: op1_11_in06 = reg_0293;
    123: op1_11_in06 = reg_0293;
    64: op1_11_in06 = reg_0406;
    33: op1_11_in06 = reg_0100;
    84: op1_11_in06 = reg_1417;
    48: op1_11_in06 = reg_0902;
    85: op1_11_in06 = reg_1243;
    65: op1_11_in06 = reg_0402;
    90: op1_11_in06 = reg_0305;
    66: op1_11_in06 = reg_0797;
    91: op1_11_in06 = reg_0803;
    67: op1_11_in06 = reg_0495;
    130: op1_11_in06 = reg_0495;
    92: op1_11_in06 = reg_0939;
    93: op1_11_in06 = reg_0938;
    94: op1_11_in06 = reg_0789;
    95: op1_11_in06 = reg_0895;
    96: op1_11_in06 = reg_0488;
    122: op1_11_in06 = reg_0488;
    97: op1_11_in06 = reg_0199;
    98: op1_11_in06 = reg_0528;
    37: op1_11_in06 = reg_0102;
    99: op1_11_in06 = reg_0805;
    101: op1_11_in06 = reg_0253;
    102: op1_11_in06 = reg_1514;
    103: op1_11_in06 = reg_0299;
    105: op1_11_in06 = reg_1027;
    106: op1_11_in06 = reg_0263;
    47: op1_11_in06 = imem04_in[7:4];
    107: op1_11_in06 = reg_1179;
    108: op1_11_in06 = reg_0229;
    109: op1_11_in06 = reg_0015;
    110: op1_11_in06 = reg_0220;
    111: op1_11_in06 = reg_0615;
    112: op1_11_in06 = reg_0276;
    113: op1_11_in06 = reg_0987;
    114: op1_11_in06 = reg_0205;
    115: op1_11_in06 = reg_1028;
    116: op1_11_in06 = reg_1340;
    117: op1_11_in06 = reg_1278;
    118: op1_11_in06 = reg_1235;
    119: op1_11_in06 = reg_1372;
    120: op1_11_in06 = reg_0707;
    121: op1_11_in06 = reg_0240;
    124: op1_11_in06 = reg_0779;
    125: op1_11_in06 = reg_0662;
    44: op1_11_in06 = reg_0304;
    34: op1_11_in06 = reg_0404;
    126: op1_11_in06 = reg_0984;
    127: op1_11_in06 = reg_1203;
    128: op1_11_in06 = reg_0582;
    38: op1_11_in06 = reg_0087;
    129: op1_11_in06 = reg_0475;
    131: op1_11_in06 = reg_0799;
    default: op1_11_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv06 = 1;
    73: op1_11_inv06 = 1;
    86: op1_11_inv06 = 1;
    49: op1_11_inv06 = 1;
    54: op1_11_inv06 = 1;
    68: op1_11_inv06 = 1;
    76: op1_11_inv06 = 1;
    87: op1_11_inv06 = 1;
    77: op1_11_inv06 = 1;
    79: op1_11_inv06 = 1;
    51: op1_11_inv06 = 1;
    60: op1_11_inv06 = 1;
    62: op1_11_inv06 = 1;
    81: op1_11_inv06 = 1;
    46: op1_11_inv06 = 1;
    82: op1_11_inv06 = 1;
    48: op1_11_inv06 = 1;
    65: op1_11_inv06 = 1;
    90: op1_11_inv06 = 1;
    93: op1_11_inv06 = 1;
    94: op1_11_inv06 = 1;
    96: op1_11_inv06 = 1;
    98: op1_11_inv06 = 1;
    100: op1_11_inv06 = 1;
    103: op1_11_inv06 = 1;
    105: op1_11_inv06 = 1;
    106: op1_11_inv06 = 1;
    111: op1_11_inv06 = 1;
    113: op1_11_inv06 = 1;
    115: op1_11_inv06 = 1;
    116: op1_11_inv06 = 1;
    117: op1_11_inv06 = 1;
    118: op1_11_inv06 = 1;
    119: op1_11_inv06 = 1;
    122: op1_11_inv06 = 1;
    124: op1_11_inv06 = 1;
    125: op1_11_inv06 = 1;
    34: op1_11_inv06 = 1;
    38: op1_11_inv06 = 1;
    129: op1_11_inv06 = 1;
    130: op1_11_inv06 = 1;
    default: op1_11_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in07 = imem00_in[3:0];
    53: op1_11_in07 = reg_0077;
    55: op1_11_in07 = imem03_in[3:0];
    73: op1_11_in07 = reg_0117;
    86: op1_11_in07 = reg_0178;
    74: op1_11_in07 = reg_1243;
    69: op1_11_in07 = reg_0180;
    49: op1_11_in07 = reg_0740;
    56: op1_11_in07 = reg_0740;
    54: op1_11_in07 = reg_0530;
    75: op1_11_in07 = imem04_in[7:4];
    50: op1_11_in07 = reg_0861;
    68: op1_11_in07 = reg_1132;
    76: op1_11_in07 = reg_0126;
    71: op1_11_in07 = reg_1281;
    87: op1_11_in07 = reg_1198;
    77: op1_11_in07 = reg_0458;
    61: op1_11_in07 = reg_0883;
    58: op1_11_in07 = reg_0062;
    78: op1_11_in07 = reg_0293;
    59: op1_11_in07 = reg_0293;
    62: op1_11_in07 = reg_0293;
    70: op1_11_in07 = reg_1029;
    79: op1_11_in07 = reg_0485;
    83: op1_11_in07 = reg_0485;
    51: op1_11_in07 = reg_0636;
    60: op1_11_in07 = reg_0159;
    88: op1_11_in07 = reg_1074;
    80: op1_11_in07 = reg_1184;
    81: op1_11_in07 = reg_0803;
    46: op1_11_in07 = reg_0794;
    52: op1_11_in07 = reg_0560;
    63: op1_11_in07 = reg_0820;
    82: op1_11_in07 = reg_0580;
    89: op1_11_in07 = reg_0882;
    64: op1_11_in07 = reg_0797;
    33: op1_11_in07 = reg_0053;
    84: op1_11_in07 = reg_1418;
    48: op1_11_in07 = reg_0868;
    85: op1_11_in07 = reg_0615;
    91: op1_11_in07 = reg_0615;
    65: op1_11_in07 = reg_0363;
    90: op1_11_in07 = reg_0837;
    66: op1_11_in07 = reg_0454;
    67: op1_11_in07 = reg_0778;
    92: op1_11_in07 = reg_0937;
    93: op1_11_in07 = reg_0090;
    94: op1_11_in07 = reg_0349;
    95: op1_11_in07 = reg_0447;
    96: op1_11_in07 = reg_1214;
    97: op1_11_in07 = reg_0452;
    98: op1_11_in07 = reg_0569;
    37: op1_11_in07 = reg_0103;
    99: op1_11_in07 = reg_1053;
    100: op1_11_in07 = reg_1041;
    101: op1_11_in07 = reg_0456;
    102: op1_11_in07 = reg_0130;
    103: op1_11_in07 = reg_0851;
    104: op1_11_in07 = reg_0523;
    105: op1_11_in07 = reg_0961;
    106: op1_11_in07 = reg_0181;
    47: op1_11_in07 = reg_0699;
    107: op1_11_in07 = reg_0116;
    108: op1_11_in07 = reg_0428;
    109: op1_11_in07 = reg_1414;
    110: op1_11_in07 = reg_1300;
    111: op1_11_in07 = reg_0555;
    112: op1_11_in07 = reg_0133;
    113: op1_11_in07 = reg_1201;
    114: op1_11_in07 = reg_0392;
    115: op1_11_in07 = reg_0221;
    123: op1_11_in07 = reg_0221;
    116: op1_11_in07 = reg_0236;
    117: op1_11_in07 = reg_0186;
    118: op1_11_in07 = reg_1018;
    119: op1_11_in07 = reg_0032;
    120: op1_11_in07 = reg_1009;
    121: op1_11_in07 = reg_0575;
    122: op1_11_in07 = reg_0421;
    124: op1_11_in07 = reg_0661;
    125: op1_11_in07 = reg_1103;
    44: op1_11_in07 = reg_0487;
    34: op1_11_in07 = reg_0620;
    126: op1_11_in07 = reg_1467;
    127: op1_11_in07 = reg_0681;
    128: op1_11_in07 = reg_0719;
    38: op1_11_in07 = reg_0520;
    129: op1_11_in07 = reg_0397;
    130: op1_11_in07 = reg_0056;
    131: op1_11_in07 = reg_0864;
    default: op1_11_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv07 = 1;
    55: op1_11_inv07 = 1;
    86: op1_11_inv07 = 1;
    69: op1_11_inv07 = 1;
    75: op1_11_inv07 = 1;
    50: op1_11_inv07 = 1;
    77: op1_11_inv07 = 1;
    61: op1_11_inv07 = 1;
    78: op1_11_inv07 = 1;
    79: op1_11_inv07 = 1;
    51: op1_11_inv07 = 1;
    59: op1_11_inv07 = 1;
    80: op1_11_inv07 = 1;
    81: op1_11_inv07 = 1;
    63: op1_11_inv07 = 1;
    83: op1_11_inv07 = 1;
    33: op1_11_inv07 = 1;
    84: op1_11_inv07 = 1;
    65: op1_11_inv07 = 1;
    91: op1_11_inv07 = 1;
    92: op1_11_inv07 = 1;
    93: op1_11_inv07 = 1;
    94: op1_11_inv07 = 1;
    97: op1_11_inv07 = 1;
    98: op1_11_inv07 = 1;
    102: op1_11_inv07 = 1;
    103: op1_11_inv07 = 1;
    110: op1_11_inv07 = 1;
    112: op1_11_inv07 = 1;
    116: op1_11_inv07 = 1;
    118: op1_11_inv07 = 1;
    122: op1_11_inv07 = 1;
    44: op1_11_inv07 = 1;
    34: op1_11_inv07 = 1;
    127: op1_11_inv07 = 1;
    128: op1_11_inv07 = 1;
    38: op1_11_inv07 = 1;
    129: op1_11_inv07 = 1;
    default: op1_11_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in08 = reg_0806;
    53: op1_11_in08 = reg_0041;
    55: op1_11_in08 = imem03_in[7:4];
    73: op1_11_in08 = reg_0211;
    86: op1_11_in08 = reg_1208;
    74: op1_11_in08 = reg_0121;
    69: op1_11_in08 = reg_0349;
    49: op1_11_in08 = reg_0621;
    54: op1_11_in08 = reg_0533;
    75: op1_11_in08 = imem04_in[11:8];
    50: op1_11_in08 = reg_0207;
    56: op1_11_in08 = reg_0415;
    68: op1_11_in08 = reg_0757;
    76: op1_11_in08 = reg_0111;
    71: op1_11_in08 = reg_1080;
    87: op1_11_in08 = reg_0681;
    77: op1_11_in08 = imem06_in[7:4];
    61: op1_11_in08 = reg_0638;
    58: op1_11_in08 = reg_0061;
    78: op1_11_in08 = reg_0221;
    70: op1_11_in08 = reg_0607;
    79: op1_11_in08 = reg_1453;
    51: op1_11_in08 = reg_0568;
    59: op1_11_in08 = reg_0476;
    60: op1_11_in08 = reg_0924;
    88: op1_11_in08 = reg_0495;
    80: op1_11_in08 = reg_1518;
    62: op1_11_in08 = reg_0202;
    81: op1_11_in08 = reg_1470;
    46: op1_11_in08 = reg_0346;
    52: op1_11_in08 = reg_0530;
    63: op1_11_in08 = reg_0606;
    82: op1_11_in08 = reg_0804;
    85: op1_11_in08 = reg_0804;
    89: op1_11_in08 = reg_1282;
    83: op1_11_in08 = reg_1393;
    64: op1_11_in08 = reg_0454;
    33: op1_11_in08 = reg_0484;
    84: op1_11_in08 = reg_0524;
    48: op1_11_in08 = reg_0290;
    65: op1_11_in08 = reg_0047;
    90: op1_11_in08 = reg_0719;
    66: op1_11_in08 = reg_0451;
    91: op1_11_in08 = reg_0555;
    67: op1_11_in08 = reg_0626;
    92: op1_11_in08 = reg_0303;
    93: op1_11_in08 = reg_0872;
    94: op1_11_in08 = reg_0954;
    95: op1_11_in08 = reg_0133;
    121: op1_11_in08 = reg_0133;
    96: op1_11_in08 = reg_0796;
    127: op1_11_in08 = reg_0796;
    97: op1_11_in08 = reg_0033;
    98: op1_11_in08 = reg_0522;
    37: op1_11_in08 = reg_0321;
    99: op1_11_in08 = reg_0821;
    100: op1_11_in08 = reg_0232;
    101: op1_11_in08 = reg_0499;
    102: op1_11_in08 = reg_0243;
    103: op1_11_in08 = reg_0156;
    104: op1_11_in08 = reg_1027;
    105: op1_11_in08 = reg_1418;
    106: op1_11_in08 = reg_1369;
    119: op1_11_in08 = reg_1369;
    47: op1_11_in08 = reg_0414;
    107: op1_11_in08 = reg_0718;
    108: op1_11_in08 = reg_0440;
    109: op1_11_in08 = reg_1315;
    110: op1_11_in08 = reg_0558;
    111: op1_11_in08 = reg_0293;
    112: op1_11_in08 = reg_0971;
    113: op1_11_in08 = reg_0460;
    114: op1_11_in08 = reg_0938;
    115: op1_11_in08 = reg_0485;
    117: op1_11_in08 = reg_0485;
    116: op1_11_in08 = reg_0064;
    118: op1_11_in08 = reg_0588;
    120: op1_11_in08 = reg_0288;
    122: op1_11_in08 = reg_0598;
    123: op1_11_in08 = reg_1417;
    124: op1_11_in08 = reg_0664;
    125: op1_11_in08 = reg_0705;
    44: op1_11_in08 = reg_0338;
    34: op1_11_in08 = reg_0028;
    126: op1_11_in08 = reg_0265;
    128: op1_11_in08 = reg_1312;
    129: op1_11_in08 = reg_1334;
    130: op1_11_in08 = reg_0455;
    131: op1_11_in08 = imem06_in[3:0];
    default: op1_11_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv08 = 1;
    86: op1_11_inv08 = 1;
    54: op1_11_inv08 = 1;
    50: op1_11_inv08 = 1;
    56: op1_11_inv08 = 1;
    68: op1_11_inv08 = 1;
    71: op1_11_inv08 = 1;
    58: op1_11_inv08 = 1;
    78: op1_11_inv08 = 1;
    70: op1_11_inv08 = 1;
    79: op1_11_inv08 = 1;
    59: op1_11_inv08 = 1;
    62: op1_11_inv08 = 1;
    81: op1_11_inv08 = 1;
    63: op1_11_inv08 = 1;
    83: op1_11_inv08 = 1;
    33: op1_11_inv08 = 1;
    84: op1_11_inv08 = 1;
    85: op1_11_inv08 = 1;
    65: op1_11_inv08 = 1;
    66: op1_11_inv08 = 1;
    91: op1_11_inv08 = 1;
    92: op1_11_inv08 = 1;
    98: op1_11_inv08 = 1;
    99: op1_11_inv08 = 1;
    100: op1_11_inv08 = 1;
    101: op1_11_inv08 = 1;
    102: op1_11_inv08 = 1;
    103: op1_11_inv08 = 1;
    106: op1_11_inv08 = 1;
    107: op1_11_inv08 = 1;
    111: op1_11_inv08 = 1;
    113: op1_11_inv08 = 1;
    116: op1_11_inv08 = 1;
    118: op1_11_inv08 = 1;
    120: op1_11_inv08 = 1;
    121: op1_11_inv08 = 1;
    122: op1_11_inv08 = 1;
    44: op1_11_inv08 = 1;
    34: op1_11_inv08 = 1;
    128: op1_11_inv08 = 1;
    129: op1_11_inv08 = 1;
    131: op1_11_inv08 = 1;
    default: op1_11_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in09 = reg_1028;
    74: op1_11_in09 = reg_1028;
    53: op1_11_in09 = reg_0666;
    55: op1_11_in09 = reg_0113;
    73: op1_11_in09 = reg_0064;
    86: op1_11_in09 = reg_0885;
    69: op1_11_in09 = reg_0954;
    49: op1_11_in09 = reg_0137;
    54: op1_11_in09 = reg_0981;
    75: op1_11_in09 = reg_0420;
    50: op1_11_in09 = reg_0206;
    56: op1_11_in09 = reg_0593;
    68: op1_11_in09 = reg_0154;
    76: op1_11_in09 = reg_0105;
    71: op1_11_in09 = reg_1078;
    87: op1_11_in09 = reg_0500;
    77: op1_11_in09 = imem06_in[11:8];
    61: op1_11_in09 = reg_0201;
    58: op1_11_in09 = reg_0792;
    78: op1_11_in09 = reg_0485;
    81: op1_11_in09 = reg_0485;
    70: op1_11_in09 = reg_0456;
    79: op1_11_in09 = reg_1230;
    51: op1_11_in09 = reg_0569;
    59: op1_11_in09 = reg_0172;
    60: op1_11_in09 = reg_0224;
    88: op1_11_in09 = reg_0778;
    80: op1_11_in09 = reg_0314;
    62: op1_11_in09 = reg_0524;
    46: op1_11_in09 = reg_0700;
    52: op1_11_in09 = reg_0533;
    63: op1_11_in09 = reg_0608;
    82: op1_11_in09 = reg_0293;
    89: op1_11_in09 = reg_0790;
    83: op1_11_in09 = reg_0134;
    64: op1_11_in09 = reg_0470;
    84: op1_11_in09 = reg_1393;
    48: op1_11_in09 = reg_0291;
    85: op1_11_in09 = reg_1471;
    65: op1_11_in09 = reg_0724;
    90: op1_11_in09 = reg_0339;
    66: op1_11_in09 = reg_0721;
    91: op1_11_in09 = reg_1027;
    111: op1_11_in09 = reg_1027;
    67: op1_11_in09 = reg_0106;
    92: op1_11_in09 = reg_0576;
    93: op1_11_in09 = reg_1484;
    94: op1_11_in09 = reg_1300;
    95: op1_11_in09 = reg_0668;
    96: op1_11_in09 = reg_0412;
    97: op1_11_in09 = reg_0369;
    98: op1_11_in09 = reg_0244;
    37: op1_11_in09 = reg_0228;
    99: op1_11_in09 = reg_1405;
    113: op1_11_in09 = reg_1405;
    100: op1_11_in09 = reg_0836;
    101: op1_11_in09 = reg_0846;
    102: op1_11_in09 = reg_0602;
    103: op1_11_in09 = reg_1094;
    104: op1_11_in09 = reg_1453;
    105: op1_11_in09 = reg_0352;
    106: op1_11_in09 = reg_1083;
    47: op1_11_in09 = reg_0471;
    107: op1_11_in09 = reg_0585;
    108: op1_11_in09 = reg_0410;
    109: op1_11_in09 = reg_0135;
    110: op1_11_in09 = reg_0178;
    112: op1_11_in09 = reg_1458;
    114: op1_11_in09 = reg_0477;
    115: op1_11_in09 = reg_1459;
    116: op1_11_in09 = imem05_in[3:0];
    117: op1_11_in09 = reg_0249;
    118: op1_11_in09 = reg_0055;
    119: op1_11_in09 = reg_0493;
    120: op1_11_in09 = reg_1325;
    121: op1_11_in09 = reg_0729;
    122: op1_11_in09 = reg_0969;
    123: op1_11_in09 = reg_1406;
    124: op1_11_in09 = reg_0366;
    125: op1_11_in09 = reg_0889;
    44: op1_11_in09 = reg_0211;
    34: op1_11_in09 = reg_0052;
    126: op1_11_in09 = reg_1508;
    127: op1_11_in09 = reg_1147;
    128: op1_11_in09 = reg_0096;
    129: op1_11_in09 = reg_1209;
    130: op1_11_in09 = reg_1207;
    131: op1_11_in09 = imem06_in[7:4];
    default: op1_11_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_11_inv09 = 1;
    69: op1_11_inv09 = 1;
    49: op1_11_inv09 = 1;
    54: op1_11_inv09 = 1;
    50: op1_11_inv09 = 1;
    56: op1_11_inv09 = 1;
    68: op1_11_inv09 = 1;
    76: op1_11_inv09 = 1;
    71: op1_11_inv09 = 1;
    87: op1_11_inv09 = 1;
    61: op1_11_inv09 = 1;
    58: op1_11_inv09 = 1;
    70: op1_11_inv09 = 1;
    59: op1_11_inv09 = 1;
    80: op1_11_inv09 = 1;
    62: op1_11_inv09 = 1;
    52: op1_11_inv09 = 1;
    63: op1_11_inv09 = 1;
    64: op1_11_inv09 = 1;
    48: op1_11_inv09 = 1;
    85: op1_11_inv09 = 1;
    65: op1_11_inv09 = 1;
    91: op1_11_inv09 = 1;
    67: op1_11_inv09 = 1;
    95: op1_11_inv09 = 1;
    98: op1_11_inv09 = 1;
    37: op1_11_inv09 = 1;
    99: op1_11_inv09 = 1;
    100: op1_11_inv09 = 1;
    103: op1_11_inv09 = 1;
    106: op1_11_inv09 = 1;
    47: op1_11_inv09 = 1;
    107: op1_11_inv09 = 1;
    111: op1_11_inv09 = 1;
    112: op1_11_inv09 = 1;
    114: op1_11_inv09 = 1;
    116: op1_11_inv09 = 1;
    117: op1_11_inv09 = 1;
    119: op1_11_inv09 = 1;
    121: op1_11_inv09 = 1;
    123: op1_11_inv09 = 1;
    125: op1_11_inv09 = 1;
    44: op1_11_inv09 = 1;
    127: op1_11_inv09 = 1;
    128: op1_11_inv09 = 1;
    129: op1_11_inv09 = 1;
    131: op1_11_inv09 = 1;
    default: op1_11_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in10 = reg_1453;
    78: op1_11_in10 = reg_1453;
    53: op1_11_in10 = reg_0629;
    76: op1_11_in10 = reg_0629;
    55: op1_11_in10 = reg_0505;
    73: op1_11_in10 = reg_0063;
    86: op1_11_in10 = reg_0507;
    74: op1_11_in10 = reg_1454;
    81: op1_11_in10 = reg_1454;
    69: op1_11_in10 = reg_1300;
    49: op1_11_in10 = reg_0053;
    37: op1_11_in10 = reg_0053;
    54: op1_11_in10 = reg_0473;
    75: op1_11_in10 = reg_0587;
    50: op1_11_in10 = reg_1030;
    56: op1_11_in10 = reg_0591;
    68: op1_11_in10 = reg_1064;
    71: op1_11_in10 = imem00_in[3:0];
    87: op1_11_in10 = reg_0094;
    77: op1_11_in10 = reg_0133;
    118: op1_11_in10 = reg_0133;
    61: op1_11_in10 = reg_0440;
    58: op1_11_in10 = reg_0793;
    70: op1_11_in10 = reg_0455;
    79: op1_11_in10 = reg_0524;
    51: op1_11_in10 = reg_0570;
    59: op1_11_in10 = reg_1230;
    60: op1_11_in10 = reg_0661;
    88: op1_11_in10 = reg_0496;
    80: op1_11_in10 = reg_1314;
    62: op1_11_in10 = reg_0928;
    46: op1_11_in10 = reg_0250;
    52: op1_11_in10 = reg_0495;
    63: op1_11_in10 = reg_0169;
    95: op1_11_in10 = reg_0169;
    82: op1_11_in10 = reg_1027;
    89: op1_11_in10 = reg_0426;
    83: op1_11_in10 = reg_0387;
    108: op1_11_in10 = reg_0387;
    64: op1_11_in10 = reg_0304;
    84: op1_11_in10 = reg_0886;
    48: op1_11_in10 = reg_0042;
    85: op1_11_in10 = reg_0249;
    115: op1_11_in10 = reg_0249;
    65: op1_11_in10 = reg_0291;
    90: op1_11_in10 = reg_0236;
    66: op1_11_in10 = reg_0837;
    91: op1_11_in10 = reg_0485;
    67: op1_11_in10 = reg_0382;
    92: op1_11_in10 = reg_0130;
    93: op1_11_in10 = reg_0197;
    94: op1_11_in10 = reg_1093;
    96: op1_11_in10 = reg_0406;
    97: op1_11_in10 = reg_0062;
    98: op1_11_in10 = imem06_in[11:8];
    99: op1_11_in10 = reg_0431;
    100: op1_11_in10 = reg_0336;
    101: op1_11_in10 = imem02_in[7:4];
    102: op1_11_in10 = reg_1346;
    103: op1_11_in10 = reg_0779;
    104: op1_11_in10 = reg_0961;
    105: op1_11_in10 = reg_0188;
    106: op1_11_in10 = reg_0552;
    47: op1_11_in10 = reg_0721;
    125: op1_11_in10 = reg_0721;
    107: op1_11_in10 = reg_0584;
    109: op1_11_in10 = reg_0309;
    110: op1_11_in10 = reg_0108;
    111: op1_11_in10 = reg_0221;
    112: op1_11_in10 = reg_0126;
    113: op1_11_in10 = reg_0428;
    114: op1_11_in10 = reg_0243;
    116: op1_11_in10 = reg_0315;
    117: op1_11_in10 = reg_0460;
    119: op1_11_in10 = reg_0694;
    120: op1_11_in10 = reg_1280;
    121: op1_11_in10 = reg_0372;
    122: op1_11_in10 = reg_0471;
    123: op1_11_in10 = reg_1405;
    124: op1_11_in10 = reg_0739;
    44: op1_11_in10 = reg_0209;
    34: op1_11_in10 = reg_0085;
    126: op1_11_in10 = reg_0716;
    127: op1_11_in10 = reg_0421;
    128: op1_11_in10 = reg_0117;
    129: op1_11_in10 = reg_0782;
    130: op1_11_in10 = reg_0494;
    131: op1_11_in10 = reg_0192;
    default: op1_11_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_11_inv10 = 1;
    86: op1_11_inv10 = 1;
    69: op1_11_inv10 = 1;
    49: op1_11_inv10 = 1;
    75: op1_11_inv10 = 1;
    50: op1_11_inv10 = 1;
    71: op1_11_inv10 = 1;
    58: op1_11_inv10 = 1;
    70: op1_11_inv10 = 1;
    79: op1_11_inv10 = 1;
    59: op1_11_inv10 = 1;
    60: op1_11_inv10 = 1;
    88: op1_11_inv10 = 1;
    80: op1_11_inv10 = 1;
    81: op1_11_inv10 = 1;
    89: op1_11_inv10 = 1;
    64: op1_11_inv10 = 1;
    48: op1_11_inv10 = 1;
    85: op1_11_inv10 = 1;
    96: op1_11_inv10 = 1;
    37: op1_11_inv10 = 1;
    100: op1_11_inv10 = 1;
    101: op1_11_inv10 = 1;
    103: op1_11_inv10 = 1;
    104: op1_11_inv10 = 1;
    106: op1_11_inv10 = 1;
    47: op1_11_inv10 = 1;
    107: op1_11_inv10 = 1;
    108: op1_11_inv10 = 1;
    110: op1_11_inv10 = 1;
    111: op1_11_inv10 = 1;
    113: op1_11_inv10 = 1;
    114: op1_11_inv10 = 1;
    116: op1_11_inv10 = 1;
    118: op1_11_inv10 = 1;
    119: op1_11_inv10 = 1;
    125: op1_11_inv10 = 1;
    44: op1_11_inv10 = 1;
    34: op1_11_inv10 = 1;
    129: op1_11_inv10 = 1;
    130: op1_11_inv10 = 1;
    default: op1_11_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in11 = reg_0249;
    74: op1_11_in11 = reg_0249;
    53: op1_11_in11 = reg_0922;
    55: op1_11_in11 = reg_0840;
    73: op1_11_in11 = reg_0370;
    86: op1_11_in11 = reg_0479;
    69: op1_11_in11 = reg_1093;
    49: op1_11_in11 = reg_0519;
    37: op1_11_in11 = reg_0519;
    54: op1_11_in11 = reg_0474;
    75: op1_11_in11 = reg_0750;
    50: op1_11_in11 = reg_1035;
    56: op1_11_in11 = reg_0085;
    68: op1_11_in11 = reg_0704;
    76: op1_11_in11 = imem02_in[3:0];
    71: op1_11_in11 = reg_1206;
    87: op1_11_in11 = reg_0452;
    77: op1_11_in11 = reg_0720;
    61: op1_11_in11 = reg_0350;
    58: op1_11_in11 = reg_0393;
    78: op1_11_in11 = reg_1229;
    85: op1_11_in11 = reg_1229;
    70: op1_11_in11 = reg_1018;
    79: op1_11_in11 = reg_1406;
    51: op1_11_in11 = reg_0529;
    59: op1_11_in11 = reg_0987;
    60: op1_11_in11 = reg_0621;
    88: op1_11_in11 = reg_0839;
    125: op1_11_in11 = reg_0839;
    80: op1_11_in11 = reg_1313;
    62: op1_11_in11 = reg_0886;
    81: op1_11_in11 = reg_1459;
    46: op1_11_in11 = reg_0565;
    52: op1_11_in11 = reg_0432;
    63: op1_11_in11 = reg_0587;
    82: op1_11_in11 = reg_1453;
    91: op1_11_in11 = reg_1453;
    89: op1_11_in11 = reg_0208;
    83: op1_11_in11 = reg_0072;
    64: op1_11_in11 = reg_0368;
    84: op1_11_in11 = reg_0189;
    48: op1_11_in11 = reg_0041;
    65: op1_11_in11 = reg_0278;
    90: op1_11_in11 = reg_0536;
    66: op1_11_in11 = reg_0719;
    67: op1_11_in11 = reg_0705;
    92: op1_11_in11 = reg_0151;
    93: op1_11_in11 = reg_0601;
    94: op1_11_in11 = reg_0104;
    95: op1_11_in11 = reg_1235;
    96: op1_11_in11 = reg_0342;
    97: op1_11_in11 = reg_0268;
    98: op1_11_in11 = reg_0023;
    99: op1_11_in11 = reg_0405;
    100: op1_11_in11 = reg_0236;
    101: op1_11_in11 = reg_0138;
    102: op1_11_in11 = reg_0344;
    114: op1_11_in11 = reg_0344;
    103: op1_11_in11 = reg_0437;
    104: op1_11_in11 = reg_0821;
    105: op1_11_in11 = reg_0134;
    106: op1_11_in11 = reg_0681;
    47: op1_11_in11 = reg_0338;
    107: op1_11_in11 = reg_0571;
    108: op1_11_in11 = reg_0073;
    109: op1_11_in11 = reg_1345;
    110: op1_11_in11 = reg_0113;
    111: op1_11_in11 = reg_1230;
    112: op1_11_in11 = reg_0112;
    113: op1_11_in11 = reg_0409;
    115: op1_11_in11 = reg_1201;
    116: op1_11_in11 = reg_0793;
    117: op1_11_in11 = reg_0229;
    118: op1_11_in11 = reg_0532;
    119: op1_11_in11 = reg_1198;
    120: op1_11_in11 = reg_0425;
    121: op1_11_in11 = reg_0870;
    122: op1_11_in11 = reg_1041;
    123: op1_11_in11 = reg_0927;
    124: op1_11_in11 = reg_0028;
    44: op1_11_in11 = reg_0063;
    34: op1_11_in11 = reg_0086;
    126: op1_11_in11 = reg_0636;
    127: op1_11_in11 = reg_0598;
    128: op1_11_in11 = reg_0095;
    129: op1_11_in11 = reg_1467;
    130: op1_11_in11 = reg_0382;
    131: op1_11_in11 = reg_0714;
    default: op1_11_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv11 = 1;
    55: op1_11_inv11 = 1;
    86: op1_11_inv11 = 1;
    69: op1_11_inv11 = 1;
    54: op1_11_inv11 = 1;
    75: op1_11_inv11 = 1;
    68: op1_11_inv11 = 1;
    76: op1_11_inv11 = 1;
    87: op1_11_inv11 = 1;
    77: op1_11_inv11 = 1;
    61: op1_11_inv11 = 1;
    79: op1_11_inv11 = 1;
    60: op1_11_inv11 = 1;
    88: op1_11_inv11 = 1;
    80: op1_11_inv11 = 1;
    62: op1_11_inv11 = 1;
    82: op1_11_inv11 = 1;
    89: op1_11_inv11 = 1;
    84: op1_11_inv11 = 1;
    48: op1_11_inv11 = 1;
    91: op1_11_inv11 = 1;
    67: op1_11_inv11 = 1;
    92: op1_11_inv11 = 1;
    93: op1_11_inv11 = 1;
    98: op1_11_inv11 = 1;
    37: op1_11_inv11 = 1;
    102: op1_11_inv11 = 1;
    104: op1_11_inv11 = 1;
    105: op1_11_inv11 = 1;
    108: op1_11_inv11 = 1;
    109: op1_11_inv11 = 1;
    110: op1_11_inv11 = 1;
    111: op1_11_inv11 = 1;
    115: op1_11_inv11 = 1;
    116: op1_11_inv11 = 1;
    117: op1_11_inv11 = 1;
    118: op1_11_inv11 = 1;
    120: op1_11_inv11 = 1;
    121: op1_11_inv11 = 1;
    125: op1_11_inv11 = 1;
    128: op1_11_inv11 = 1;
    130: op1_11_inv11 = 1;
    default: op1_11_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in12 = reg_1205;
    81: op1_11_in12 = reg_1205;
    85: op1_11_in12 = reg_1205;
    53: op1_11_in12 = imem02_in[11:8];
    55: op1_11_in12 = reg_0849;
    73: op1_11_in12 = reg_1164;
    86: op1_11_in12 = imem03_in[3:0];
    74: op1_11_in12 = reg_1206;
    69: op1_11_in12 = reg_0478;
    54: op1_11_in12 = reg_0989;
    75: op1_11_in12 = reg_1298;
    50: op1_11_in12 = reg_0194;
    56: op1_11_in12 = reg_0124;
    37: op1_11_in12 = reg_0124;
    68: op1_11_in12 = reg_0376;
    76: op1_11_in12 = reg_0712;
    71: op1_11_in12 = reg_1406;
    87: op1_11_in12 = reg_0305;
    77: op1_11_in12 = reg_0869;
    61: op1_11_in12 = reg_0058;
    105: op1_11_in12 = reg_0058;
    108: op1_11_in12 = reg_0058;
    58: op1_11_in12 = reg_0578;
    78: op1_11_in12 = reg_0961;
    70: op1_11_in12 = reg_0590;
    79: op1_11_in12 = reg_0928;
    51: op1_11_in12 = reg_0527;
    59: op1_11_in12 = reg_0459;
    60: op1_11_in12 = reg_0592;
    88: op1_11_in12 = reg_1031;
    80: op1_11_in12 = reg_0558;
    62: op1_11_in12 = reg_0410;
    46: op1_11_in12 = reg_0316;
    52: op1_11_in12 = reg_0326;
    63: op1_11_in12 = reg_0562;
    82: op1_11_in12 = reg_0722;
    89: op1_11_in12 = reg_0263;
    83: op1_11_in12 = reg_0059;
    64: op1_11_in12 = reg_0065;
    84: op1_11_in12 = reg_0073;
    113: op1_11_in12 = reg_0073;
    48: op1_11_in12 = reg_0011;
    65: op1_11_in12 = reg_0043;
    90: op1_11_in12 = reg_0095;
    66: op1_11_in12 = reg_0211;
    91: op1_11_in12 = reg_1227;
    67: op1_11_in12 = reg_0711;
    92: op1_11_in12 = reg_0207;
    93: op1_11_in12 = reg_0393;
    94: op1_11_in12 = reg_0882;
    110: op1_11_in12 = reg_0882;
    95: op1_11_in12 = reg_0456;
    96: op1_11_in12 = reg_1143;
    97: op1_11_in12 = reg_0932;
    98: op1_11_in12 = reg_0213;
    99: op1_11_in12 = reg_0134;
    100: op1_11_in12 = reg_0035;
    101: op1_11_in12 = reg_0934;
    102: op1_11_in12 = reg_0799;
    103: op1_11_in12 = reg_0408;
    104: op1_11_in12 = reg_0476;
    106: op1_11_in12 = reg_0796;
    47: op1_11_in12 = reg_0096;
    107: op1_11_in12 = reg_0570;
    109: op1_11_in12 = reg_0157;
    111: op1_11_in12 = reg_0987;
    112: op1_11_in12 = reg_0897;
    114: op1_11_in12 = reg_0206;
    115: op1_11_in12 = reg_0460;
    116: op1_11_in12 = reg_0338;
    117: op1_11_in12 = reg_1417;
    118: op1_11_in12 = reg_0497;
    119: op1_11_in12 = reg_0574;
    120: op1_11_in12 = reg_0208;
    121: op1_11_in12 = reg_0730;
    122: op1_11_in12 = reg_1040;
    123: op1_11_in12 = reg_0060;
    124: op1_11_in12 = reg_1439;
    125: op1_11_in12 = reg_0054;
    44: op1_11_in12 = reg_0016;
    34: op1_11_in12 = reg_0519;
    126: op1_11_in12 = reg_0374;
    127: op1_11_in12 = reg_0969;
    128: op1_11_in12 = reg_0420;
    129: op1_11_in12 = reg_0827;
    130: op1_11_in12 = reg_0496;
    131: op1_11_in12 = reg_0751;
    default: op1_11_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv12 = 1;
    55: op1_11_inv12 = 1;
    73: op1_11_inv12 = 1;
    86: op1_11_inv12 = 1;
    74: op1_11_inv12 = 1;
    69: op1_11_inv12 = 1;
    54: op1_11_inv12 = 1;
    75: op1_11_inv12 = 1;
    56: op1_11_inv12 = 1;
    68: op1_11_inv12 = 1;
    76: op1_11_inv12 = 1;
    58: op1_11_inv12 = 1;
    70: op1_11_inv12 = 1;
    62: op1_11_inv12 = 1;
    81: op1_11_inv12 = 1;
    46: op1_11_inv12 = 1;
    52: op1_11_inv12 = 1;
    83: op1_11_inv12 = 1;
    48: op1_11_inv12 = 1;
    91: op1_11_inv12 = 1;
    67: op1_11_inv12 = 1;
    93: op1_11_inv12 = 1;
    94: op1_11_inv12 = 1;
    95: op1_11_inv12 = 1;
    97: op1_11_inv12 = 1;
    37: op1_11_inv12 = 1;
    103: op1_11_inv12 = 1;
    105: op1_11_inv12 = 1;
    108: op1_11_inv12 = 1;
    111: op1_11_inv12 = 1;
    114: op1_11_inv12 = 1;
    115: op1_11_inv12 = 1;
    124: op1_11_inv12 = 1;
    125: op1_11_inv12 = 1;
    44: op1_11_inv12 = 1;
    129: op1_11_inv12 = 1;
    default: op1_11_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in13 = reg_0459;
    53: op1_11_in13 = reg_0472;
    55: op1_11_in13 = reg_0426;
    73: op1_11_in13 = reg_1163;
    86: op1_11_in13 = reg_0427;
    74: op1_11_in13 = reg_0155;
    69: op1_11_in13 = reg_0849;
    54: op1_11_in13 = reg_0990;
    75: op1_11_in13 = reg_0833;
    116: op1_11_in13 = reg_0833;
    50: op1_11_in13 = reg_0195;
    68: op1_11_in13 = reg_1139;
    76: op1_11_in13 = reg_0708;
    71: op1_11_in13 = reg_0476;
    87: op1_11_in13 = reg_0338;
    77: op1_11_in13 = reg_0752;
    61: op1_11_in13 = reg_0089;
    58: op1_11_in13 = reg_0750;
    78: op1_11_in13 = reg_0229;
    70: op1_11_in13 = reg_0497;
    79: op1_11_in13 = reg_0886;
    91: op1_11_in13 = reg_0886;
    51: op1_11_in13 = reg_0522;
    59: op1_11_in13 = reg_1148;
    60: op1_11_in13 = reg_0361;
    88: op1_11_in13 = reg_0381;
    80: op1_11_in13 = reg_0178;
    62: op1_11_in13 = reg_0134;
    81: op1_11_in13 = reg_1432;
    85: op1_11_in13 = reg_1432;
    46: op1_11_in13 = reg_0163;
    52: op1_11_in13 = reg_0111;
    63: op1_11_in13 = reg_0561;
    101: op1_11_in13 = reg_0561;
    82: op1_11_in13 = reg_0428;
    89: op1_11_in13 = reg_1372;
    83: op1_11_in13 = reg_0057;
    113: op1_11_in13 = reg_0057;
    64: op1_11_in13 = reg_0208;
    84: op1_11_in13 = reg_0072;
    123: op1_11_in13 = reg_0072;
    48: op1_11_in13 = reg_0256;
    65: op1_11_in13 = reg_0679;
    90: op1_11_in13 = reg_0633;
    66: op1_11_in13 = reg_0064;
    67: op1_11_in13 = imem02_in[15:12];
    92: op1_11_in13 = reg_0040;
    114: op1_11_in13 = reg_0040;
    93: op1_11_in13 = reg_0344;
    94: op1_11_in13 = reg_1009;
    95: op1_11_in13 = reg_0934;
    96: op1_11_in13 = reg_0932;
    97: op1_11_in13 = reg_0536;
    98: op1_11_in13 = reg_0018;
    99: op1_11_in13 = reg_0387;
    100: op1_11_in13 = reg_0470;
    102: op1_11_in13 = reg_0864;
    103: op1_11_in13 = reg_0618;
    104: op1_11_in13 = reg_0887;
    105: op1_11_in13 = reg_0355;
    106: op1_11_in13 = reg_1040;
    47: op1_11_in13 = reg_0129;
    107: op1_11_in13 = reg_0396;
    108: op1_11_in13 = reg_0027;
    109: op1_11_in13 = reg_0921;
    110: op1_11_in13 = reg_1149;
    111: op1_11_in13 = reg_1201;
    112: op1_11_in13 = reg_0801;
    115: op1_11_in13 = reg_0821;
    117: op1_11_in13 = reg_1418;
    118: op1_11_in13 = reg_0533;
    119: op1_11_in13 = reg_0488;
    120: op1_11_in13 = reg_0164;
    121: op1_11_in13 = reg_1326;
    122: op1_11_in13 = reg_0199;
    124: op1_11_in13 = reg_0998;
    125: op1_11_in13 = reg_0105;
    44: op1_11_in13 = reg_0032;
    126: op1_11_in13 = reg_0585;
    127: op1_11_in13 = reg_0320;
    128: op1_11_in13 = imem05_in[11:8];
    129: op1_11_in13 = reg_0109;
    130: op1_11_in13 = reg_0876;
    131: op1_11_in13 = reg_0869;
    default: op1_11_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv13 = 1;
    55: op1_11_inv13 = 1;
    69: op1_11_inv13 = 1;
    54: op1_11_inv13 = 1;
    75: op1_11_inv13 = 1;
    50: op1_11_inv13 = 1;
    76: op1_11_inv13 = 1;
    71: op1_11_inv13 = 1;
    87: op1_11_inv13 = 1;
    70: op1_11_inv13 = 1;
    79: op1_11_inv13 = 1;
    60: op1_11_inv13 = 1;
    88: op1_11_inv13 = 1;
    62: op1_11_inv13 = 1;
    81: op1_11_inv13 = 1;
    82: op1_11_inv13 = 1;
    89: op1_11_inv13 = 1;
    48: op1_11_inv13 = 1;
    85: op1_11_inv13 = 1;
    65: op1_11_inv13 = 1;
    67: op1_11_inv13 = 1;
    92: op1_11_inv13 = 1;
    96: op1_11_inv13 = 1;
    98: op1_11_inv13 = 1;
    101: op1_11_inv13 = 1;
    103: op1_11_inv13 = 1;
    106: op1_11_inv13 = 1;
    108: op1_11_inv13 = 1;
    110: op1_11_inv13 = 1;
    112: op1_11_inv13 = 1;
    114: op1_11_inv13 = 1;
    115: op1_11_inv13 = 1;
    116: op1_11_inv13 = 1;
    117: op1_11_inv13 = 1;
    118: op1_11_inv13 = 1;
    119: op1_11_inv13 = 1;
    120: op1_11_inv13 = 1;
    121: op1_11_inv13 = 1;
    123: op1_11_inv13 = 1;
    124: op1_11_inv13 = 1;
    127: op1_11_inv13 = 1;
    131: op1_11_inv13 = 1;
    default: op1_11_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in14 = reg_0189;
    53: op1_11_in14 = reg_0473;
    55: op1_11_in14 = reg_0443;
    73: op1_11_in14 = reg_0173;
    86: op1_11_in14 = reg_0898;
    74: op1_11_in14 = reg_0524;
    69: op1_11_in14 = reg_0208;
    54: op1_11_in14 = reg_0972;
    75: op1_11_in14 = reg_0168;
    50: op1_11_in14 = reg_0870;
    68: op1_11_in14 = reg_0143;
    76: op1_11_in14 = reg_0294;
    71: op1_11_in14 = reg_0927;
    117: op1_11_in14 = reg_0927;
    87: op1_11_in14 = reg_0096;
    77: op1_11_in14 = reg_0984;
    61: op1_11_in14 = imem01_in[15:12];
    58: op1_11_in14 = imem05_in[3:0];
    78: op1_11_in14 = reg_0887;
    70: op1_11_in14 = reg_0631;
    79: op1_11_in14 = reg_0351;
    104: op1_11_in14 = reg_0351;
    111: op1_11_in14 = reg_0351;
    51: op1_11_in14 = reg_0323;
    59: op1_11_in14 = reg_0883;
    60: op1_11_in14 = reg_0051;
    88: op1_11_in14 = reg_0379;
    130: op1_11_in14 = reg_0379;
    80: op1_11_in14 = reg_0107;
    62: op1_11_in14 = reg_0075;
    81: op1_11_in14 = reg_1417;
    46: op1_11_in14 = reg_0418;
    52: op1_11_in14 = reg_0138;
    63: op1_11_in14 = reg_0560;
    82: op1_11_in14 = reg_0409;
    89: op1_11_in14 = reg_0181;
    83: op1_11_in14 = reg_0122;
    64: op1_11_in14 = reg_0064;
    84: op1_11_in14 = reg_0059;
    48: op1_11_in14 = reg_0629;
    125: op1_11_in14 = reg_0629;
    85: op1_11_in14 = reg_1406;
    65: op1_11_in14 = reg_0457;
    90: op1_11_in14 = reg_0370;
    66: op1_11_in14 = reg_0021;
    91: op1_11_in14 = reg_0202;
    115: op1_11_in14 = reg_0202;
    67: op1_11_in14 = reg_0632;
    92: op1_11_in14 = imem06_in[3:0];
    93: op1_11_in14 = reg_0753;
    94: op1_11_in14 = reg_0291;
    95: op1_11_in14 = reg_0055;
    96: op1_11_in14 = reg_0117;
    97: op1_11_in14 = reg_0095;
    98: op1_11_in14 = reg_1439;
    99: op1_11_in14 = reg_0389;
    100: op1_11_in14 = reg_0793;
    101: op1_11_in14 = reg_1344;
    102: op1_11_in14 = reg_1030;
    103: op1_11_in14 = reg_0103;
    105: op1_11_in14 = reg_0549;
    106: op1_11_in14 = reg_0452;
    47: op1_11_in14 = reg_0020;
    107: op1_11_in14 = reg_0215;
    108: op1_11_in14 = reg_0183;
    109: op1_11_in14 = reg_1094;
    110: op1_11_in14 = reg_0378;
    112: op1_11_in14 = reg_0253;
    113: op1_11_in14 = reg_1255;
    114: op1_11_in14 = reg_1058;
    116: op1_11_in14 = reg_0136;
    118: op1_11_in14 = reg_0900;
    119: op1_11_in14 = reg_1215;
    120: op1_11_in14 = reg_0263;
    121: op1_11_in14 = reg_1501;
    122: op1_11_in14 = reg_0320;
    123: op1_11_in14 = reg_0089;
    124: op1_11_in14 = reg_0519;
    44: op1_11_in14 = reg_0579;
    126: op1_11_in14 = reg_0622;
    127: op1_11_in14 = reg_0062;
    128: op1_11_in14 = reg_0567;
    129: op1_11_in14 = reg_0584;
    131: op1_11_in14 = reg_0752;
    default: op1_11_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv14 = 1;
    55: op1_11_inv14 = 1;
    86: op1_11_inv14 = 1;
    74: op1_11_inv14 = 1;
    54: op1_11_inv14 = 1;
    76: op1_11_inv14 = 1;
    77: op1_11_inv14 = 1;
    61: op1_11_inv14 = 1;
    78: op1_11_inv14 = 1;
    79: op1_11_inv14 = 1;
    51: op1_11_inv14 = 1;
    59: op1_11_inv14 = 1;
    60: op1_11_inv14 = 1;
    46: op1_11_inv14 = 1;
    52: op1_11_inv14 = 1;
    63: op1_11_inv14 = 1;
    82: op1_11_inv14 = 1;
    83: op1_11_inv14 = 1;
    64: op1_11_inv14 = 1;
    48: op1_11_inv14 = 1;
    90: op1_11_inv14 = 1;
    94: op1_11_inv14 = 1;
    99: op1_11_inv14 = 1;
    104: op1_11_inv14 = 1;
    47: op1_11_inv14 = 1;
    108: op1_11_inv14 = 1;
    109: op1_11_inv14 = 1;
    117: op1_11_inv14 = 1;
    118: op1_11_inv14 = 1;
    119: op1_11_inv14 = 1;
    120: op1_11_inv14 = 1;
    121: op1_11_inv14 = 1;
    122: op1_11_inv14 = 1;
    126: op1_11_inv14 = 1;
    127: op1_11_inv14 = 1;
    128: op1_11_inv14 = 1;
    130: op1_11_inv14 = 1;
    131: op1_11_inv14 = 1;
    default: op1_11_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in15 = reg_0059;
    53: op1_11_in15 = reg_0776;
    55: op1_11_in15 = reg_0594;
    73: op1_11_in15 = reg_0272;
    86: op1_11_in15 = reg_1372;
    74: op1_11_in15 = reg_0352;
    71: op1_11_in15 = reg_0352;
    69: op1_11_in15 = reg_1339;
    54: op1_11_in15 = reg_0934;
    75: op1_11_in15 = reg_0347;
    100: op1_11_in15 = reg_0347;
    50: op1_11_in15 = reg_0116;
    68: op1_11_in15 = reg_0234;
    76: op1_11_in15 = reg_0009;
    87: op1_11_in15 = reg_0065;
    77: op1_11_in15 = reg_0717;
    61: op1_11_in15 = reg_0160;
    58: op1_11_in15 = reg_1169;
    78: op1_11_in15 = reg_0188;
    70: op1_11_in15 = reg_0475;
    79: op1_11_in15 = reg_0431;
    115: op1_11_in15 = reg_0431;
    51: op1_11_in15 = reg_0419;
    59: op1_11_in15 = reg_0388;
    60: op1_11_in15 = reg_0086;
    88: op1_11_in15 = reg_0560;
    80: op1_11_in15 = reg_0113;
    62: op1_11_in15 = imem00_in[11:8];
    81: op1_11_in15 = reg_0410;
    46: op1_11_in15 = reg_0207;
    52: op1_11_in15 = reg_0712;
    101: op1_11_in15 = reg_0712;
    63: op1_11_in15 = reg_0497;
    82: op1_11_in15 = reg_0134;
    89: op1_11_in15 = reg_0034;
    83: op1_11_in15 = reg_0026;
    64: op1_11_in15 = reg_0020;
    84: op1_11_in15 = reg_1321;
    48: op1_11_in15 = reg_0608;
    85: op1_11_in15 = reg_0887;
    65: op1_11_in15 = reg_0744;
    90: op1_11_in15 = imem05_in[15:12];
    66: op1_11_in15 = reg_0391;
    91: op1_11_in15 = reg_0351;
    67: op1_11_in15 = reg_0006;
    92: op1_11_in15 = reg_1058;
    93: op1_11_in15 = reg_1508;
    94: op1_11_in15 = reg_1139;
    95: op1_11_in15 = reg_0839;
    96: op1_11_in15 = reg_0021;
    97: op1_11_in15 = reg_0633;
    98: op1_11_in15 = reg_1414;
    99: op1_11_in15 = reg_0058;
    102: op1_11_in15 = reg_0931;
    103: op1_11_in15 = reg_0028;
    104: op1_11_in15 = reg_0428;
    105: op1_11_in15 = reg_0747;
    106: op1_11_in15 = reg_0342;
    122: op1_11_in15 = reg_0342;
    47: op1_11_in15 = reg_0395;
    107: op1_11_in15 = reg_0214;
    108: op1_11_in15 = reg_0166;
    109: op1_11_in15 = reg_0774;
    110: op1_11_in15 = reg_0673;
    111: op1_11_in15 = reg_0389;
    112: op1_11_in15 = reg_1006;
    113: op1_11_in15 = reg_1253;
    114: op1_11_in15 = imem06_in[7:4];
    116: op1_11_in15 = reg_0332;
    117: op1_11_in15 = reg_0881;
    118: op1_11_in15 = reg_1207;
    119: op1_11_in15 = reg_0681;
    120: op1_11_in15 = imem04_in[3:0];
    121: op1_11_in15 = reg_0172;
    123: op1_11_in15 = reg_0723;
    124: op1_11_in15 = reg_0520;
    125: op1_11_in15 = reg_0684;
    44: op1_11_in15 = reg_0175;
    126: op1_11_in15 = reg_0529;
    127: op1_11_in15 = reg_0209;
    128: op1_11_in15 = reg_0278;
    129: op1_11_in15 = reg_0571;
    130: op1_11_in15 = reg_0897;
    131: op1_11_in15 = reg_1505;
    default: op1_11_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv15 = 1;
    53: op1_11_inv15 = 1;
    55: op1_11_inv15 = 1;
    73: op1_11_inv15 = 1;
    74: op1_11_inv15 = 1;
    50: op1_11_inv15 = 1;
    68: op1_11_inv15 = 1;
    76: op1_11_inv15 = 1;
    71: op1_11_inv15 = 1;
    77: op1_11_inv15 = 1;
    61: op1_11_inv15 = 1;
    58: op1_11_inv15 = 1;
    78: op1_11_inv15 = 1;
    70: op1_11_inv15 = 1;
    59: op1_11_inv15 = 1;
    60: op1_11_inv15 = 1;
    88: op1_11_inv15 = 1;
    80: op1_11_inv15 = 1;
    81: op1_11_inv15 = 1;
    63: op1_11_inv15 = 1;
    82: op1_11_inv15 = 1;
    89: op1_11_inv15 = 1;
    83: op1_11_inv15 = 1;
    84: op1_11_inv15 = 1;
    48: op1_11_inv15 = 1;
    65: op1_11_inv15 = 1;
    90: op1_11_inv15 = 1;
    67: op1_11_inv15 = 1;
    93: op1_11_inv15 = 1;
    97: op1_11_inv15 = 1;
    98: op1_11_inv15 = 1;
    102: op1_11_inv15 = 1;
    47: op1_11_inv15 = 1;
    108: op1_11_inv15 = 1;
    110: op1_11_inv15 = 1;
    112: op1_11_inv15 = 1;
    116: op1_11_inv15 = 1;
    118: op1_11_inv15 = 1;
    119: op1_11_inv15 = 1;
    120: op1_11_inv15 = 1;
    123: op1_11_inv15 = 1;
    124: op1_11_inv15 = 1;
    125: op1_11_inv15 = 1;
    128: op1_11_inv15 = 1;
    131: op1_11_inv15 = 1;
    default: op1_11_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in16 = reg_1322;
    53: op1_11_in16 = reg_0326;
    55: op1_11_in16 = reg_0463;
    73: op1_11_in16 = reg_1404;
    86: op1_11_in16 = imem04_in[7:4];
    74: op1_11_in16 = reg_0388;
    69: op1_11_in16 = reg_1215;
    54: op1_11_in16 = reg_0126;
    75: op1_11_in16 = reg_1169;
    50: op1_11_in16 = reg_0671;
    68: op1_11_in16 = reg_1000;
    76: op1_11_in16 = reg_0531;
    71: op1_11_in16 = reg_0188;
    87: op1_11_in16 = reg_0420;
    77: op1_11_in16 = reg_0637;
    61: op1_11_in16 = reg_0166;
    58: op1_11_in16 = reg_0334;
    78: op1_11_in16 = reg_0201;
    70: op1_11_in16 = reg_0432;
    118: op1_11_in16 = reg_0432;
    79: op1_11_in16 = reg_0387;
    82: op1_11_in16 = reg_0387;
    51: op1_11_in16 = reg_0119;
    59: op1_11_in16 = reg_0352;
    88: op1_11_in16 = reg_0711;
    80: op1_11_in16 = reg_0505;
    62: op1_11_in16 = reg_0788;
    81: op1_11_in16 = reg_0073;
    46: op1_11_in16 = reg_0782;
    52: op1_11_in16 = reg_0876;
    63: op1_11_in16 = reg_0889;
    89: op1_11_in16 = reg_0552;
    83: op1_11_in16 = reg_0027;
    99: op1_11_in16 = reg_0027;
    64: op1_11_in16 = reg_0792;
    96: op1_11_in16 = reg_0792;
    84: op1_11_in16 = reg_0026;
    48: op1_11_in16 = imem02_in[7:4];
    85: op1_11_in16 = reg_0431;
    91: op1_11_in16 = reg_0431;
    65: op1_11_in16 = reg_1029;
    90: op1_11_in16 = reg_0737;
    66: op1_11_in16 = reg_1299;
    67: op1_11_in16 = reg_0677;
    92: op1_11_in16 = reg_0193;
    93: op1_11_in16 = reg_1030;
    94: op1_11_in16 = reg_1280;
    95: op1_11_in16 = reg_1002;
    97: op1_11_in16 = reg_0367;
    98: op1_11_in16 = reg_1055;
    100: op1_11_in16 = reg_0648;
    101: op1_11_in16 = reg_0744;
    102: op1_11_in16 = reg_0161;
    103: op1_11_in16 = reg_0084;
    104: op1_11_in16 = reg_0409;
    105: op1_11_in16 = reg_1473;
    106: op1_11_in16 = reg_0061;
    47: op1_11_in16 = reg_0745;
    107: op1_11_in16 = reg_0018;
    108: op1_11_in16 = reg_1255;
    109: op1_11_in16 = reg_0031;
    110: op1_11_in16 = reg_0288;
    111: op1_11_in16 = reg_0075;
    112: op1_11_in16 = reg_0750;
    113: op1_11_in16 = reg_1031;
    114: op1_11_in16 = imem06_in[15:12];
    115: op1_11_in16 = reg_0440;
    116: op1_11_in16 = reg_0395;
    117: op1_11_in16 = reg_0883;
    119: op1_11_in16 = reg_1233;
    120: op1_11_in16 = imem04_in[11:8];
    121: op1_11_in16 = reg_0116;
    122: op1_11_in16 = reg_0837;
    123: op1_11_in16 = reg_0785;
    124: op1_11_in16 = reg_1182;
    125: op1_11_in16 = reg_0631;
    44: op1_11_in16 = reg_0066;
    126: op1_11_in16 = reg_1225;
    127: op1_11_in16 = reg_0633;
    128: op1_11_in16 = reg_0538;
    129: op1_11_in16 = reg_0522;
    130: op1_11_in16 = reg_0800;
    131: op1_11_in16 = reg_0571;
    default: op1_11_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv16 = 1;
    55: op1_11_inv16 = 1;
    74: op1_11_inv16 = 1;
    69: op1_11_inv16 = 1;
    68: op1_11_inv16 = 1;
    76: op1_11_inv16 = 1;
    70: op1_11_inv16 = 1;
    88: op1_11_inv16 = 1;
    80: op1_11_inv16 = 1;
    62: op1_11_inv16 = 1;
    81: op1_11_inv16 = 1;
    63: op1_11_inv16 = 1;
    82: op1_11_inv16 = 1;
    89: op1_11_inv16 = 1;
    83: op1_11_inv16 = 1;
    64: op1_11_inv16 = 1;
    84: op1_11_inv16 = 1;
    66: op1_11_inv16 = 1;
    92: op1_11_inv16 = 1;
    95: op1_11_inv16 = 1;
    96: op1_11_inv16 = 1;
    98: op1_11_inv16 = 1;
    99: op1_11_inv16 = 1;
    100: op1_11_inv16 = 1;
    102: op1_11_inv16 = 1;
    103: op1_11_inv16 = 1;
    109: op1_11_inv16 = 1;
    113: op1_11_inv16 = 1;
    114: op1_11_inv16 = 1;
    115: op1_11_inv16 = 1;
    116: op1_11_inv16 = 1;
    121: op1_11_inv16 = 1;
    123: op1_11_inv16 = 1;
    124: op1_11_inv16 = 1;
    125: op1_11_inv16 = 1;
    44: op1_11_inv16 = 1;
    default: op1_11_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in17 = reg_1100;
    53: op1_11_in17 = reg_0778;
    55: op1_11_in17 = reg_0462;
    73: op1_11_in17 = reg_0940;
    86: op1_11_in17 = reg_0421;
    74: op1_11_in17 = reg_0071;
    104: op1_11_in17 = reg_0071;
    69: op1_11_in17 = reg_1200;
    54: op1_11_in17 = reg_0381;
    75: op1_11_in17 = reg_0346;
    50: op1_11_in17 = reg_0670;
    68: op1_11_in17 = reg_1003;
    76: op1_11_in17 = reg_0846;
    71: op1_11_in17 = reg_0059;
    87: op1_11_in17 = reg_0021;
    77: op1_11_in17 = reg_0374;
    61: op1_11_in17 = reg_1291;
    58: op1_11_in17 = reg_0317;
    78: op1_11_in17 = reg_0440;
    70: op1_11_in17 = reg_0972;
    79: op1_11_in17 = reg_0389;
    91: op1_11_in17 = reg_0389;
    51: op1_11_in17 = reg_0067;
    59: op1_11_in17 = reg_0075;
    81: op1_11_in17 = reg_0075;
    88: op1_11_in17 = reg_1091;
    80: op1_11_in17 = reg_0525;
    62: op1_11_in17 = reg_1071;
    46: op1_11_in17 = reg_0780;
    52: op1_11_in17 = reg_0879;
    63: op1_11_in17 = reg_1207;
    82: op1_11_in17 = reg_1321;
    89: op1_11_in17 = reg_0574;
    83: op1_11_in17 = reg_0005;
    84: op1_11_in17 = reg_0005;
    64: op1_11_in17 = reg_1299;
    48: op1_11_in17 = reg_0588;
    85: op1_11_in17 = reg_0435;
    115: op1_11_in17 = reg_0435;
    65: op1_11_in17 = reg_0606;
    90: op1_11_in17 = reg_0579;
    128: op1_11_in17 = reg_0579;
    66: op1_11_in17 = reg_0733;
    67: op1_11_in17 = reg_0121;
    92: op1_11_in17 = reg_0397;
    93: op1_11_in17 = reg_0193;
    94: op1_11_in17 = reg_0341;
    95: op1_11_in17 = reg_0432;
    96: op1_11_in17 = reg_1169;
    97: op1_11_in17 = reg_0466;
    98: op1_11_in17 = reg_0478;
    99: op1_11_in17 = imem01_in[7:4];
    100: op1_11_in17 = reg_0701;
    101: op1_11_in17 = reg_1451;
    102: op1_11_in17 = reg_0870;
    103: op1_11_in17 = reg_0519;
    105: op1_11_in17 = reg_0726;
    106: op1_11_in17 = reg_0262;
    47: op1_11_in17 = reg_0347;
    107: op1_11_in17 = reg_0893;
    108: op1_11_in17 = reg_0549;
    109: op1_11_in17 = reg_0465;
    110: op1_11_in17 = reg_1282;
    111: op1_11_in17 = reg_0026;
    112: op1_11_in17 = reg_0709;
    113: op1_11_in17 = reg_0788;
    114: op1_11_in17 = reg_1209;
    116: op1_11_in17 = reg_1268;
    117: op1_11_in17 = reg_0189;
    118: op1_11_in17 = reg_0382;
    119: op1_11_in17 = reg_0281;
    120: op1_11_in17 = reg_0264;
    121: op1_11_in17 = reg_0637;
    122: op1_11_in17 = reg_1146;
    123: op1_11_in17 = reg_0576;
    125: op1_11_in17 = reg_0306;
    44: op1_11_in17 = reg_0334;
    126: op1_11_in17 = reg_0022;
    127: op1_11_in17 = reg_0338;
    129: op1_11_in17 = reg_0323;
    130: op1_11_in17 = reg_1006;
    131: op1_11_in17 = reg_0165;
    default: op1_11_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_11_inv17 = 1;
    74: op1_11_inv17 = 1;
    69: op1_11_inv17 = 1;
    54: op1_11_inv17 = 1;
    75: op1_11_inv17 = 1;
    76: op1_11_inv17 = 1;
    77: op1_11_inv17 = 1;
    61: op1_11_inv17 = 1;
    78: op1_11_inv17 = 1;
    79: op1_11_inv17 = 1;
    62: op1_11_inv17 = 1;
    81: op1_11_inv17 = 1;
    46: op1_11_inv17 = 1;
    52: op1_11_inv17 = 1;
    63: op1_11_inv17 = 1;
    82: op1_11_inv17 = 1;
    83: op1_11_inv17 = 1;
    84: op1_11_inv17 = 1;
    90: op1_11_inv17 = 1;
    66: op1_11_inv17 = 1;
    92: op1_11_inv17 = 1;
    94: op1_11_inv17 = 1;
    95: op1_11_inv17 = 1;
    96: op1_11_inv17 = 1;
    98: op1_11_inv17 = 1;
    99: op1_11_inv17 = 1;
    101: op1_11_inv17 = 1;
    103: op1_11_inv17 = 1;
    104: op1_11_inv17 = 1;
    105: op1_11_inv17 = 1;
    106: op1_11_inv17 = 1;
    47: op1_11_inv17 = 1;
    109: op1_11_inv17 = 1;
    112: op1_11_inv17 = 1;
    113: op1_11_inv17 = 1;
    117: op1_11_inv17 = 1;
    118: op1_11_inv17 = 1;
    121: op1_11_inv17 = 1;
    123: op1_11_inv17 = 1;
    44: op1_11_inv17 = 1;
    126: op1_11_inv17 = 1;
    128: op1_11_inv17 = 1;
    129: op1_11_inv17 = 1;
    131: op1_11_inv17 = 1;
    default: op1_11_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in18 = reg_0822;
    53: op1_11_in18 = reg_0935;
    55: op1_11_in18 = reg_0978;
    73: op1_11_in18 = reg_0070;
    86: op1_11_in18 = reg_0471;
    74: op1_11_in18 = reg_0089;
    69: op1_11_in18 = reg_1065;
    54: op1_11_in18 = reg_0839;
    75: op1_11_in18 = reg_0174;
    50: op1_11_in18 = reg_0634;
    68: op1_11_in18 = reg_1314;
    76: op1_11_in18 = reg_0695;
    71: op1_11_in18 = reg_0917;
    87: op1_11_in18 = reg_0035;
    77: op1_11_in18 = reg_0586;
    61: op1_11_in18 = reg_1031;
    58: op1_11_in18 = reg_0540;
    78: op1_11_in18 = reg_0409;
    70: op1_11_in18 = reg_0128;
    101: op1_11_in18 = reg_0128;
    79: op1_11_in18 = reg_0075;
    51: op1_11_in18 = reg_0023;
    59: op1_11_in18 = reg_0060;
    88: op1_11_in18 = reg_0328;
    80: op1_11_in18 = reg_0425;
    62: op1_11_in18 = reg_1032;
    81: op1_11_in18 = reg_0058;
    46: op1_11_in18 = reg_0751;
    52: op1_11_in18 = reg_0845;
    63: op1_11_in18 = reg_0432;
    82: op1_11_in18 = reg_0026;
    89: op1_11_in18 = reg_1214;
    83: op1_11_in18 = reg_0278;
    127: op1_11_in18 = reg_0278;
    64: op1_11_in18 = reg_0251;
    84: op1_11_in18 = reg_1100;
    48: op1_11_in18 = reg_0475;
    85: op1_11_in18 = reg_0203;
    91: op1_11_in18 = reg_0203;
    104: op1_11_in18 = reg_0203;
    65: op1_11_in18 = reg_0532;
    90: op1_11_in18 = reg_0315;
    66: op1_11_in18 = reg_0702;
    67: op1_11_in18 = reg_0707;
    92: op1_11_in18 = reg_0372;
    93: op1_11_in18 = reg_0795;
    94: op1_11_in18 = imem04_in[3:0];
    95: op1_11_in18 = reg_0127;
    96: op1_11_in18 = imem05_in[15:12];
    97: op1_11_in18 = reg_0184;
    98: op1_11_in18 = reg_0894;
    99: op1_11_in18 = reg_0785;
    100: op1_11_in18 = reg_0491;
    44: op1_11_in18 = reg_0491;
    102: op1_11_in18 = reg_1420;
    103: op1_11_in18 = reg_0520;
    105: op1_11_in18 = reg_0149;
    106: op1_11_in18 = reg_0338;
    47: op1_11_in18 = reg_0700;
    116: op1_11_in18 = reg_0700;
    107: op1_11_in18 = reg_1414;
    108: op1_11_in18 = reg_0747;
    109: op1_11_in18 = reg_0739;
    110: op1_11_in18 = reg_0426;
    111: op1_11_in18 = imem01_in[15:12];
    112: op1_11_in18 = reg_0330;
    113: op1_11_in18 = reg_0871;
    114: op1_11_in18 = reg_0960;
    115: op1_11_in18 = reg_0388;
    117: op1_11_in18 = reg_0440;
    118: op1_11_in18 = reg_0306;
    119: op1_11_in18 = reg_0500;
    120: op1_11_in18 = reg_0034;
    121: op1_11_in18 = reg_0398;
    122: op1_11_in18 = reg_0096;
    123: op1_11_in18 = reg_0746;
    125: op1_11_in18 = reg_0802;
    126: op1_11_in18 = reg_0017;
    128: op1_11_in18 = reg_0040;
    129: op1_11_in18 = reg_1204;
    130: op1_11_in18 = reg_0069;
    131: op1_11_in18 = reg_0067;
    default: op1_11_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv18 = 1;
    55: op1_11_inv18 = 1;
    74: op1_11_inv18 = 1;
    54: op1_11_inv18 = 1;
    50: op1_11_inv18 = 1;
    68: op1_11_inv18 = 1;
    76: op1_11_inv18 = 1;
    87: op1_11_inv18 = 1;
    77: op1_11_inv18 = 1;
    78: op1_11_inv18 = 1;
    70: op1_11_inv18 = 1;
    79: op1_11_inv18 = 1;
    46: op1_11_inv18 = 1;
    52: op1_11_inv18 = 1;
    89: op1_11_inv18 = 1;
    83: op1_11_inv18 = 1;
    64: op1_11_inv18 = 1;
    48: op1_11_inv18 = 1;
    85: op1_11_inv18 = 1;
    90: op1_11_inv18 = 1;
    66: op1_11_inv18 = 1;
    92: op1_11_inv18 = 1;
    96: op1_11_inv18 = 1;
    97: op1_11_inv18 = 1;
    98: op1_11_inv18 = 1;
    99: op1_11_inv18 = 1;
    100: op1_11_inv18 = 1;
    101: op1_11_inv18 = 1;
    104: op1_11_inv18 = 1;
    106: op1_11_inv18 = 1;
    108: op1_11_inv18 = 1;
    109: op1_11_inv18 = 1;
    110: op1_11_inv18 = 1;
    112: op1_11_inv18 = 1;
    113: op1_11_inv18 = 1;
    114: op1_11_inv18 = 1;
    115: op1_11_inv18 = 1;
    117: op1_11_inv18 = 1;
    125: op1_11_inv18 = 1;
    44: op1_11_inv18 = 1;
    126: op1_11_inv18 = 1;
    130: op1_11_inv18 = 1;
    131: op1_11_inv18 = 1;
    default: op1_11_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in19 = reg_0166;
    59: op1_11_in19 = reg_0166;
    53: op1_11_in19 = reg_0105;
    101: op1_11_in19 = reg_0105;
    55: op1_11_in19 = reg_0407;
    73: op1_11_in19 = reg_0090;
    86: op1_11_in19 = reg_1041;
    74: op1_11_in19 = reg_0027;
    69: op1_11_in19 = reg_0406;
    119: op1_11_in19 = reg_0406;
    54: op1_11_in19 = reg_0007;
    75: op1_11_in19 = reg_1212;
    50: op1_11_in19 = reg_0584;
    68: op1_11_in19 = reg_0957;
    76: op1_11_in19 = reg_0069;
    71: op1_11_in19 = reg_0786;
    87: op1_11_in19 = reg_0833;
    77: op1_11_in19 = reg_0568;
    61: op1_11_in19 = reg_1034;
    62: op1_11_in19 = reg_1034;
    58: op1_11_in19 = reg_0938;
    78: op1_11_in19 = reg_0388;
    70: op1_11_in19 = reg_0126;
    79: op1_11_in19 = reg_1321;
    51: op1_11_in19 = reg_0046;
    88: op1_11_in19 = reg_0707;
    80: op1_11_in19 = reg_0411;
    81: op1_11_in19 = reg_0057;
    46: op1_11_in19 = reg_0192;
    52: op1_11_in19 = reg_0068;
    63: op1_11_in19 = reg_0054;
    82: op1_11_in19 = imem01_in[3:0];
    89: op1_11_in19 = reg_1147;
    83: op1_11_in19 = reg_0982;
    64: op1_11_in19 = reg_0395;
    84: op1_11_in19 = reg_0679;
    48: op1_11_in19 = reg_0127;
    85: op1_11_in19 = reg_0060;
    104: op1_11_in19 = reg_0060;
    65: op1_11_in19 = reg_0253;
    90: op1_11_in19 = reg_1299;
    66: op1_11_in19 = reg_0831;
    91: op1_11_in19 = reg_0075;
    67: op1_11_in19 = reg_1064;
    92: op1_11_in19 = reg_0635;
    93: op1_11_in19 = reg_0397;
    94: op1_11_in19 = reg_0264;
    95: op1_11_in19 = reg_0631;
    96: op1_11_in19 = reg_1430;
    97: op1_11_in19 = reg_0992;
    98: op1_11_in19 = reg_0851;
    99: op1_11_in19 = reg_0963;
    100: op1_11_in19 = reg_1484;
    102: op1_11_in19 = reg_0782;
    103: op1_11_in19 = reg_0123;
    105: op1_11_in19 = reg_0895;
    106: op1_11_in19 = reg_0096;
    47: op1_11_in19 = reg_0697;
    107: op1_11_in19 = reg_1056;
    108: op1_11_in19 = reg_0820;
    109: op1_11_in19 = reg_0413;
    110: op1_11_in19 = reg_0443;
    111: op1_11_in19 = reg_0120;
    112: op1_11_in19 = imem03_in[7:4];
    113: op1_11_in19 = reg_0902;
    114: op1_11_in19 = reg_1467;
    115: op1_11_in19 = reg_0203;
    116: op1_11_in19 = reg_0996;
    117: op1_11_in19 = reg_0073;
    118: op1_11_in19 = reg_0800;
    125: op1_11_in19 = reg_0800;
    120: op1_11_in19 = reg_1258;
    121: op1_11_in19 = reg_0624;
    122: op1_11_in19 = reg_0064;
    123: op1_11_in19 = reg_0609;
    44: op1_11_in19 = imem05_in[7:4];
    126: op1_11_in19 = reg_0169;
    127: op1_11_in19 = reg_0648;
    128: op1_11_in19 = reg_0251;
    129: op1_11_in19 = reg_1202;
    130: op1_11_in19 = reg_1515;
    131: op1_11_in19 = reg_0213;
    default: op1_11_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_11_inv19 = 1;
    74: op1_11_inv19 = 1;
    54: op1_11_inv19 = 1;
    75: op1_11_inv19 = 1;
    50: op1_11_inv19 = 1;
    68: op1_11_inv19 = 1;
    77: op1_11_inv19 = 1;
    61: op1_11_inv19 = 1;
    70: op1_11_inv19 = 1;
    51: op1_11_inv19 = 1;
    88: op1_11_inv19 = 1;
    62: op1_11_inv19 = 1;
    46: op1_11_inv19 = 1;
    63: op1_11_inv19 = 1;
    82: op1_11_inv19 = 1;
    64: op1_11_inv19 = 1;
    84: op1_11_inv19 = 1;
    48: op1_11_inv19 = 1;
    90: op1_11_inv19 = 1;
    67: op1_11_inv19 = 1;
    97: op1_11_inv19 = 1;
    107: op1_11_inv19 = 1;
    108: op1_11_inv19 = 1;
    109: op1_11_inv19 = 1;
    113: op1_11_inv19 = 1;
    115: op1_11_inv19 = 1;
    116: op1_11_inv19 = 1;
    117: op1_11_inv19 = 1;
    119: op1_11_inv19 = 1;
    120: op1_11_inv19 = 1;
    123: op1_11_inv19 = 1;
    125: op1_11_inv19 = 1;
    44: op1_11_inv19 = 1;
    129: op1_11_inv19 = 1;
    130: op1_11_inv19 = 1;
    default: op1_11_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in20 = reg_0549;
    53: op1_11_in20 = reg_0138;
    55: op1_11_in20 = reg_0451;
    73: op1_11_in20 = imem05_in[11:8];
    86: op1_11_in20 = reg_1077;
    74: op1_11_in20 = reg_0917;
    69: op1_11_in20 = reg_0407;
    89: op1_11_in20 = reg_0407;
    54: op1_11_in20 = reg_0281;
    76: op1_11_in20 = reg_0281;
    75: op1_11_in20 = reg_0131;
    50: op1_11_in20 = reg_0526;
    68: op1_11_in20 = reg_0246;
    71: op1_11_in20 = reg_0788;
    87: op1_11_in20 = reg_0347;
    77: op1_11_in20 = reg_0570;
    61: op1_11_in20 = reg_0548;
    58: op1_11_in20 = reg_0163;
    78: op1_11_in20 = reg_0072;
    70: op1_11_in20 = reg_0382;
    79: op1_11_in20 = reg_1068;
    51: op1_11_in20 = reg_0213;
    59: op1_11_in20 = reg_0786;
    88: op1_11_in20 = reg_0143;
    80: op1_11_in20 = reg_0898;
    62: op1_11_in20 = reg_0611;
    81: op1_11_in20 = reg_0026;
    46: op1_11_in20 = imem06_in[3:0];
    52: op1_11_in20 = reg_0800;
    63: op1_11_in20 = reg_0973;
    82: op1_11_in20 = imem01_in[11:8];
    83: op1_11_in20 = reg_0448;
    64: op1_11_in20 = reg_1168;
    84: op1_11_in20 = reg_0278;
    48: op1_11_in20 = reg_0111;
    85: op1_11_in20 = reg_1321;
    65: op1_11_in20 = reg_0590;
    90: op1_11_in20 = reg_0332;
    66: op1_11_in20 = reg_0832;
    91: op1_11_in20 = reg_0060;
    67: op1_11_in20 = reg_0145;
    92: op1_11_in20 = reg_0717;
    93: op1_11_in20 = reg_0870;
    94: op1_11_in20 = reg_0797;
    95: op1_11_in20 = reg_0380;
    96: op1_11_in20 = reg_0136;
    97: op1_11_in20 = reg_0831;
    98: op1_11_in20 = reg_0457;
    107: op1_11_in20 = reg_0457;
    99: op1_11_in20 = reg_0553;
    100: op1_11_in20 = reg_0130;
    101: op1_11_in20 = reg_0381;
    102: op1_11_in20 = reg_1467;
    104: op1_11_in20 = reg_0122;
    117: op1_11_in20 = reg_0122;
    105: op1_11_in20 = reg_0447;
    106: op1_11_in20 = reg_0063;
    47: op1_11_in20 = reg_0175;
    108: op1_11_in20 = reg_0572;
    109: op1_11_in20 = reg_0100;
    110: op1_11_in20 = imem04_in[15:12];
    111: op1_11_in20 = reg_0282;
    112: op1_11_in20 = reg_0177;
    113: op1_11_in20 = reg_0047;
    114: op1_11_in20 = reg_0860;
    115: op1_11_in20 = reg_0013;
    116: op1_11_in20 = reg_1104;
    118: op1_11_in20 = reg_0903;
    119: op1_11_in20 = reg_0599;
    120: op1_11_in20 = reg_0552;
    121: op1_11_in20 = reg_1225;
    122: op1_11_in20 = reg_1503;
    123: op1_11_in20 = reg_0742;
    125: op1_11_in20 = reg_1078;
    44: op1_11_in20 = reg_0895;
    126: op1_11_in20 = reg_0084;
    127: op1_11_in20 = reg_0315;
    128: op1_11_in20 = reg_0996;
    129: op1_11_in20 = reg_0023;
    130: op1_11_in20 = reg_0330;
    131: op1_11_in20 = reg_0025;
    default: op1_11_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv20 = 1;
    73: op1_11_inv20 = 1;
    50: op1_11_inv20 = 1;
    76: op1_11_inv20 = 1;
    78: op1_11_inv20 = 1;
    79: op1_11_inv20 = 1;
    51: op1_11_inv20 = 1;
    59: op1_11_inv20 = 1;
    88: op1_11_inv20 = 1;
    80: op1_11_inv20 = 1;
    62: op1_11_inv20 = 1;
    81: op1_11_inv20 = 1;
    46: op1_11_inv20 = 1;
    82: op1_11_inv20 = 1;
    89: op1_11_inv20 = 1;
    84: op1_11_inv20 = 1;
    48: op1_11_inv20 = 1;
    65: op1_11_inv20 = 1;
    90: op1_11_inv20 = 1;
    91: op1_11_inv20 = 1;
    93: op1_11_inv20 = 1;
    95: op1_11_inv20 = 1;
    96: op1_11_inv20 = 1;
    101: op1_11_inv20 = 1;
    102: op1_11_inv20 = 1;
    111: op1_11_inv20 = 1;
    112: op1_11_inv20 = 1;
    117: op1_11_inv20 = 1;
    118: op1_11_inv20 = 1;
    119: op1_11_inv20 = 1;
    122: op1_11_inv20 = 1;
    125: op1_11_inv20 = 1;
    44: op1_11_inv20 = 1;
    126: op1_11_inv20 = 1;
    128: op1_11_inv20 = 1;
    default: op1_11_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in21 = reg_0550;
    53: op1_11_in21 = reg_0897;
    55: op1_11_in21 = reg_0320;
    73: op1_11_in21 = reg_1373;
    86: op1_11_in21 = reg_1004;
    74: op1_11_in21 = reg_0335;
    69: op1_11_in21 = reg_0599;
    54: op1_11_in21 = reg_0755;
    75: op1_11_in21 = reg_0567;
    50: op1_11_in21 = reg_0165;
    68: op1_11_in21 = reg_1300;
    76: op1_11_in21 = reg_1515;
    71: op1_11_in21 = reg_1032;
    87: op1_11_in21 = reg_0184;
    77: op1_11_in21 = reg_0296;
    61: op1_11_in21 = reg_0746;
    58: op1_11_in21 = reg_0896;
    78: op1_11_in21 = reg_0026;
    70: op1_11_in21 = reg_0695;
    79: op1_11_in21 = imem01_in[11:8];
    51: op1_11_in21 = reg_0191;
    59: op1_11_in21 = reg_0785;
    88: op1_11_in21 = reg_0220;
    80: op1_11_in21 = reg_1312;
    62: op1_11_in21 = reg_0372;
    81: op1_11_in21 = reg_0446;
    46: op1_11_in21 = reg_0397;
    52: op1_11_in21 = imem03_in[7:4];
    63: op1_11_in21 = reg_0106;
    48: op1_11_in21 = reg_0106;
    82: op1_11_in21 = reg_1512;
    89: op1_11_in21 = reg_0199;
    83: op1_11_in21 = reg_1291;
    64: op1_11_in21 = reg_1163;
    84: op1_11_in21 = reg_1290;
    115: op1_11_in21 = reg_1290;
    85: op1_11_in21 = reg_0089;
    65: op1_11_in21 = reg_0589;
    90: op1_11_in21 = reg_0278;
    66: op1_11_in21 = reg_1164;
    91: op1_11_in21 = reg_1322;
    67: op1_11_in21 = reg_0559;
    92: op1_11_in21 = reg_0714;
    93: op1_11_in21 = reg_1209;
    94: op1_11_in21 = reg_1258;
    95: op1_11_in21 = reg_0381;
    96: op1_11_in21 = reg_0333;
    97: op1_11_in21 = reg_0648;
    98: op1_11_in21 = reg_1345;
    99: op1_11_in21 = reg_0093;
    100: op1_11_in21 = reg_0118;
    101: op1_11_in21 = reg_0745;
    102: op1_11_in21 = reg_0860;
    104: op1_11_in21 = reg_1254;
    105: op1_11_in21 = reg_0662;
    106: op1_11_in21 = reg_0019;
    47: op1_11_in21 = reg_0250;
    107: op1_11_in21 = reg_1347;
    108: op1_11_in21 = reg_0967;
    109: op1_11_in21 = reg_0114;
    110: op1_11_in21 = reg_0252;
    111: op1_11_in21 = reg_1034;
    112: op1_11_in21 = reg_0145;
    113: op1_11_in21 = reg_0547;
    114: op1_11_in21 = reg_1501;
    116: op1_11_in21 = reg_0630;
    117: op1_11_in21 = reg_0027;
    118: op1_11_in21 = reg_1078;
    119: op1_11_in21 = reg_1041;
    120: op1_11_in21 = reg_0421;
    121: op1_11_in21 = reg_0132;
    122: op1_11_in21 = reg_0038;
    123: op1_11_in21 = reg_0726;
    125: op1_11_in21 = reg_0255;
    44: op1_11_in21 = reg_0873;
    126: op1_11_in21 = reg_0298;
    127: op1_11_in21 = reg_1168;
    128: op1_11_in21 = reg_0491;
    129: op1_11_in21 = reg_0152;
    130: op1_11_in21 = reg_0246;
    131: op1_11_in21 = reg_1055;
    default: op1_11_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv21 = 1;
    55: op1_11_inv21 = 1;
    73: op1_11_inv21 = 1;
    86: op1_11_inv21 = 1;
    74: op1_11_inv21 = 1;
    69: op1_11_inv21 = 1;
    68: op1_11_inv21 = 1;
    76: op1_11_inv21 = 1;
    61: op1_11_inv21 = 1;
    58: op1_11_inv21 = 1;
    78: op1_11_inv21 = 1;
    70: op1_11_inv21 = 1;
    88: op1_11_inv21 = 1;
    80: op1_11_inv21 = 1;
    62: op1_11_inv21 = 1;
    81: op1_11_inv21 = 1;
    52: op1_11_inv21 = 1;
    89: op1_11_inv21 = 1;
    83: op1_11_inv21 = 1;
    84: op1_11_inv21 = 1;
    85: op1_11_inv21 = 1;
    65: op1_11_inv21 = 1;
    66: op1_11_inv21 = 1;
    93: op1_11_inv21 = 1;
    94: op1_11_inv21 = 1;
    95: op1_11_inv21 = 1;
    96: op1_11_inv21 = 1;
    97: op1_11_inv21 = 1;
    99: op1_11_inv21 = 1;
    100: op1_11_inv21 = 1;
    101: op1_11_inv21 = 1;
    102: op1_11_inv21 = 1;
    105: op1_11_inv21 = 1;
    106: op1_11_inv21 = 1;
    107: op1_11_inv21 = 1;
    109: op1_11_inv21 = 1;
    114: op1_11_inv21 = 1;
    116: op1_11_inv21 = 1;
    118: op1_11_inv21 = 1;
    120: op1_11_inv21 = 1;
    123: op1_11_inv21 = 1;
    44: op1_11_inv21 = 1;
    127: op1_11_inv21 = 1;
    129: op1_11_inv21 = 1;
    130: op1_11_inv21 = 1;
    131: op1_11_inv21 = 1;
    default: op1_11_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in22 = reg_0610;
    113: op1_11_in22 = reg_0610;
    53: op1_11_in22 = reg_0708;
    63: op1_11_in22 = reg_0708;
    55: op1_11_in22 = reg_0904;
    73: op1_11_in22 = reg_0601;
    86: op1_11_in22 = reg_0452;
    89: op1_11_in22 = reg_0452;
    74: op1_11_in22 = reg_1254;
    83: op1_11_in22 = reg_1254;
    69: op1_11_in22 = reg_0797;
    54: op1_11_in22 = imem03_in[7:4];
    75: op1_11_in22 = reg_0272;
    50: op1_11_in22 = reg_0270;
    68: op1_11_in22 = reg_1231;
    76: op1_11_in22 = reg_1494;
    71: op1_11_in22 = reg_0166;
    87: op1_11_in22 = reg_0992;
    90: op1_11_in22 = reg_0992;
    77: op1_11_in22 = reg_0295;
    61: op1_11_in22 = reg_0259;
    58: op1_11_in22 = reg_0895;
    78: op1_11_in22 = reg_0027;
    70: op1_11_in22 = reg_0632;
    79: op1_11_in22 = reg_0553;
    51: op1_11_in22 = imem07_in[7:4];
    59: op1_11_in22 = imem01_in[15:12];
    88: op1_11_in22 = reg_0350;
    80: op1_11_in22 = reg_1339;
    62: op1_11_in22 = reg_0634;
    81: op1_11_in22 = reg_1071;
    46: op1_11_in22 = reg_0860;
    52: op1_11_in22 = imem03_in[15:12];
    82: op1_11_in22 = reg_0258;
    64: op1_11_in22 = reg_0346;
    84: op1_11_in22 = reg_0788;
    48: op1_11_in22 = reg_0105;
    85: op1_11_in22 = reg_0723;
    65: op1_11_in22 = reg_1343;
    66: op1_11_in22 = reg_0646;
    91: op1_11_in22 = reg_0985;
    67: op1_11_in22 = reg_1001;
    92: op1_11_in22 = reg_0584;
    93: op1_11_in22 = reg_0974;
    94: op1_11_in22 = reg_0462;
    95: op1_11_in22 = reg_0307;
    96: op1_11_in22 = reg_0347;
    97: op1_11_in22 = reg_1070;
    98: op1_11_in22 = reg_0159;
    99: op1_11_in22 = reg_0242;
    100: op1_11_in22 = reg_0861;
    101: op1_11_in22 = reg_0802;
    102: op1_11_in22 = reg_0752;
    104: op1_11_in22 = reg_0902;
    105: op1_11_in22 = imem02_in[3:0];
    106: op1_11_in22 = reg_0021;
    47: op1_11_in22 = reg_0523;
    107: op1_11_in22 = reg_1349;
    108: op1_11_in22 = reg_1456;
    109: op1_11_in22 = reg_0321;
    110: op1_11_in22 = reg_1372;
    111: op1_11_in22 = reg_1152;
    112: op1_11_in22 = reg_0891;
    114: op1_11_in22 = reg_0780;
    115: op1_11_in22 = reg_0047;
    116: op1_11_in22 = reg_1180;
    117: op1_11_in22 = reg_1100;
    118: op1_11_in22 = reg_1006;
    119: op1_11_in22 = reg_1040;
    120: op1_11_in22 = reg_0414;
    121: op1_11_in22 = reg_0296;
    122: op1_11_in22 = reg_0735;
    123: op1_11_in22 = reg_0400;
    125: op1_11_in22 = reg_0006;
    44: op1_11_in22 = reg_0184;
    126: op1_11_in22 = reg_0667;
    127: op1_11_in22 = reg_0395;
    128: op1_11_in22 = reg_0564;
    129: op1_11_in22 = reg_0029;
    130: op1_11_in22 = reg_1063;
    131: op1_11_in22 = reg_1315;
    default: op1_11_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv22 = 1;
    53: op1_11_inv22 = 1;
    55: op1_11_inv22 = 1;
    86: op1_11_inv22 = 1;
    69: op1_11_inv22 = 1;
    54: op1_11_inv22 = 1;
    50: op1_11_inv22 = 1;
    68: op1_11_inv22 = 1;
    76: op1_11_inv22 = 1;
    77: op1_11_inv22 = 1;
    79: op1_11_inv22 = 1;
    51: op1_11_inv22 = 1;
    59: op1_11_inv22 = 1;
    80: op1_11_inv22 = 1;
    62: op1_11_inv22 = 1;
    52: op1_11_inv22 = 1;
    63: op1_11_inv22 = 1;
    89: op1_11_inv22 = 1;
    83: op1_11_inv22 = 1;
    64: op1_11_inv22 = 1;
    84: op1_11_inv22 = 1;
    66: op1_11_inv22 = 1;
    92: op1_11_inv22 = 1;
    94: op1_11_inv22 = 1;
    97: op1_11_inv22 = 1;
    98: op1_11_inv22 = 1;
    99: op1_11_inv22 = 1;
    101: op1_11_inv22 = 1;
    102: op1_11_inv22 = 1;
    105: op1_11_inv22 = 1;
    107: op1_11_inv22 = 1;
    108: op1_11_inv22 = 1;
    111: op1_11_inv22 = 1;
    113: op1_11_inv22 = 1;
    114: op1_11_inv22 = 1;
    118: op1_11_inv22 = 1;
    120: op1_11_inv22 = 1;
    122: op1_11_inv22 = 1;
    123: op1_11_inv22 = 1;
    125: op1_11_inv22 = 1;
    44: op1_11_inv22 = 1;
    126: op1_11_inv22 = 1;
    129: op1_11_inv22 = 1;
    130: op1_11_inv22 = 1;
    131: op1_11_inv22 = 1;
    default: op1_11_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in23 = reg_0966;
    53: op1_11_in23 = reg_0307;
    55: op1_11_in23 = reg_0340;
    73: op1_11_in23 = reg_0196;
    86: op1_11_in23 = reg_0061;
    74: op1_11_in23 = reg_1256;
    78: op1_11_in23 = reg_1256;
    69: op1_11_in23 = imem04_in[11:8];
    54: op1_11_in23 = reg_0707;
    125: op1_11_in23 = reg_0707;
    75: op1_11_in23 = reg_1181;
    128: op1_11_in23 = reg_1181;
    50: op1_11_in23 = reg_0212;
    68: op1_11_in23 = reg_1208;
    76: op1_11_in23 = reg_0999;
    71: op1_11_in23 = reg_0547;
    62: op1_11_in23 = reg_0547;
    82: op1_11_in23 = reg_0547;
    87: op1_11_in23 = reg_0648;
    77: op1_11_in23 = reg_0371;
    46: op1_11_in23 = reg_0371;
    61: op1_11_in23 = reg_0553;
    104: op1_11_in23 = reg_0553;
    58: op1_11_in23 = reg_0300;
    70: op1_11_in23 = reg_0217;
    79: op1_11_in23 = reg_0163;
    51: op1_11_in23 = imem07_in[11:8];
    59: op1_11_in23 = reg_0576;
    111: op1_11_in23 = reg_0576;
    88: op1_11_in23 = reg_0288;
    80: op1_11_in23 = reg_1216;
    81: op1_11_in23 = imem01_in[3:0];
    52: op1_11_in23 = reg_0573;
    63: op1_11_in23 = reg_0306;
    89: op1_11_in23 = reg_0232;
    83: op1_11_in23 = reg_0047;
    64: op1_11_in23 = reg_0646;
    84: op1_11_in23 = reg_1291;
    48: op1_11_in23 = reg_0711;
    101: op1_11_in23 = reg_0711;
    85: op1_11_in23 = reg_0611;
    65: op1_11_in23 = reg_1207;
    90: op1_11_in23 = reg_0562;
    66: op1_11_in23 = reg_0066;
    91: op1_11_in23 = reg_0963;
    67: op1_11_in23 = reg_0965;
    92: op1_11_in23 = reg_0527;
    93: op1_11_in23 = reg_0859;
    94: op1_11_in23 = reg_0297;
    95: op1_11_in23 = reg_0829;
    96: op1_11_in23 = reg_1268;
    97: op1_11_in23 = reg_0873;
    98: op1_11_in23 = reg_0158;
    99: op1_11_in23 = reg_0238;
    100: op1_11_in23 = reg_0784;
    102: op1_11_in23 = reg_1501;
    105: op1_11_in23 = reg_0253;
    106: op1_11_in23 = reg_1488;
    47: op1_11_in23 = imem05_in[3:0];
    107: op1_11_in23 = reg_0159;
    108: op1_11_in23 = reg_0385;
    109: op1_11_in23 = reg_0003;
    110: op1_11_in23 = reg_1369;
    112: op1_11_in23 = reg_0556;
    113: op1_11_in23 = reg_0787;
    114: op1_11_in23 = reg_0115;
    115: op1_11_in23 = reg_0463;
    116: op1_11_in23 = reg_1402;
    117: op1_11_in23 = imem01_in[7:4];
    118: op1_11_in23 = reg_0068;
    119: op1_11_in23 = reg_1004;
    120: op1_11_in23 = reg_0487;
    121: op1_11_in23 = reg_1204;
    122: op1_11_in23 = reg_1168;
    123: op1_11_in23 = reg_0724;
    44: op1_11_in23 = reg_0130;
    126: op1_11_in23 = reg_0050;
    127: op1_11_in23 = reg_0272;
    129: op1_11_in23 = reg_0087;
    130: op1_11_in23 = reg_0783;
    131: op1_11_in23 = reg_0298;
    default: op1_11_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv23 = 1;
    55: op1_11_inv23 = 1;
    86: op1_11_inv23 = 1;
    74: op1_11_inv23 = 1;
    69: op1_11_inv23 = 1;
    54: op1_11_inv23 = 1;
    76: op1_11_inv23 = 1;
    61: op1_11_inv23 = 1;
    58: op1_11_inv23 = 1;
    70: op1_11_inv23 = 1;
    51: op1_11_inv23 = 1;
    59: op1_11_inv23 = 1;
    81: op1_11_inv23 = 1;
    82: op1_11_inv23 = 1;
    84: op1_11_inv23 = 1;
    48: op1_11_inv23 = 1;
    67: op1_11_inv23 = 1;
    93: op1_11_inv23 = 1;
    97: op1_11_inv23 = 1;
    98: op1_11_inv23 = 1;
    99: op1_11_inv23 = 1;
    100: op1_11_inv23 = 1;
    101: op1_11_inv23 = 1;
    102: op1_11_inv23 = 1;
    104: op1_11_inv23 = 1;
    105: op1_11_inv23 = 1;
    107: op1_11_inv23 = 1;
    108: op1_11_inv23 = 1;
    113: op1_11_inv23 = 1;
    115: op1_11_inv23 = 1;
    116: op1_11_inv23 = 1;
    117: op1_11_inv23 = 1;
    119: op1_11_inv23 = 1;
    120: op1_11_inv23 = 1;
    121: op1_11_inv23 = 1;
    122: op1_11_inv23 = 1;
    123: op1_11_inv23 = 1;
    44: op1_11_inv23 = 1;
    127: op1_11_inv23 = 1;
    130: op1_11_inv23 = 1;
    default: op1_11_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in24 = reg_0967;
    53: op1_11_in24 = reg_0839;
    55: op1_11_in24 = reg_0262;
    73: op1_11_in24 = reg_0797;
    86: op1_11_in24 = reg_0304;
    74: op1_11_in24 = reg_1031;
    69: op1_11_in24 = reg_0368;
    54: op1_11_in24 = reg_0314;
    75: op1_11_in24 = reg_0090;
    50: op1_11_in24 = reg_0017;
    68: op1_11_in24 = reg_0113;
    76: op1_11_in24 = reg_0235;
    71: op1_11_in24 = reg_0550;
    115: op1_11_in24 = reg_0550;
    87: op1_11_in24 = reg_0491;
    90: op1_11_in24 = reg_0491;
    77: op1_11_in24 = reg_0270;
    61: op1_11_in24 = reg_0715;
    58: op1_11_in24 = reg_0251;
    96: op1_11_in24 = reg_0251;
    78: op1_11_in24 = imem01_in[15:12];
    70: op1_11_in24 = reg_0311;
    79: op1_11_in24 = reg_0260;
    51: op1_11_in24 = reg_1060;
    59: op1_11_in24 = reg_0575;
    88: op1_11_in24 = reg_1282;
    80: op1_11_in24 = reg_1082;
    62: op1_11_in24 = imem01_in[7:4];
    81: op1_11_in24 = reg_0448;
    46: op1_11_in24 = reg_0826;
    52: op1_11_in24 = reg_1064;
    100: op1_11_in24 = reg_1064;
    63: op1_11_in24 = reg_0878;
    82: op1_11_in24 = reg_0548;
    89: op1_11_in24 = reg_0340;
    83: op1_11_in24 = reg_0258;
    64: op1_11_in24 = reg_0649;
    84: op1_11_in24 = reg_1253;
    48: op1_11_in24 = reg_0068;
    85: op1_11_in24 = reg_0982;
    65: op1_11_in24 = reg_0432;
    66: op1_11_in24 = reg_0333;
    91: op1_11_in24 = reg_1511;
    67: op1_11_in24 = reg_0963;
    92: op1_11_in24 = reg_1225;
    93: op1_11_in24 = reg_0869;
    94: op1_11_in24 = reg_1200;
    95: op1_11_in24 = reg_0560;
    97: op1_11_in24 = reg_1373;
    98: op1_11_in24 = reg_0921;
    99: op1_11_in24 = reg_0830;
    101: op1_11_in24 = reg_0695;
    102: op1_11_in24 = reg_0110;
    104: op1_11_in24 = reg_0798;
    105: op1_11_in24 = reg_0846;
    106: op1_11_in24 = reg_0370;
    47: op1_11_in24 = reg_0331;
    107: op1_11_in24 = reg_0158;
    108: op1_11_in24 = reg_0360;
    110: op1_11_in24 = reg_0535;
    111: op1_11_in24 = reg_0163;
    112: op1_11_in24 = reg_0964;
    113: op1_11_in24 = reg_0743;
    114: op1_11_in24 = reg_0619;
    116: op1_11_in24 = reg_0938;
    117: op1_11_in24 = reg_0747;
    118: op1_11_in24 = reg_0217;
    119: op1_11_in24 = reg_0451;
    120: op1_11_in24 = reg_0862;
    121: op1_11_in24 = reg_0371;
    122: op1_11_in24 = reg_0604;
    123: op1_11_in24 = reg_0162;
    125: op1_11_in24 = reg_0479;
    44: op1_11_in24 = reg_0272;
    126: op1_11_in24 = reg_0786;
    127: op1_11_in24 = reg_1268;
    128: op1_11_in24 = reg_1070;
    129: op1_11_in24 = reg_0003;
    130: op1_11_in24 = reg_0145;
    131: op1_11_in24 = reg_0170;
    default: op1_11_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_11_inv24 = 1;
    73: op1_11_inv24 = 1;
    74: op1_11_inv24 = 1;
    50: op1_11_inv24 = 1;
    71: op1_11_inv24 = 1;
    77: op1_11_inv24 = 1;
    58: op1_11_inv24 = 1;
    78: op1_11_inv24 = 1;
    51: op1_11_inv24 = 1;
    59: op1_11_inv24 = 1;
    88: op1_11_inv24 = 1;
    80: op1_11_inv24 = 1;
    46: op1_11_inv24 = 1;
    52: op1_11_inv24 = 1;
    63: op1_11_inv24 = 1;
    89: op1_11_inv24 = 1;
    65: op1_11_inv24 = 1;
    90: op1_11_inv24 = 1;
    91: op1_11_inv24 = 1;
    93: op1_11_inv24 = 1;
    95: op1_11_inv24 = 1;
    96: op1_11_inv24 = 1;
    98: op1_11_inv24 = 1;
    100: op1_11_inv24 = 1;
    110: op1_11_inv24 = 1;
    113: op1_11_inv24 = 1;
    116: op1_11_inv24 = 1;
    117: op1_11_inv24 = 1;
    119: op1_11_inv24 = 1;
    120: op1_11_inv24 = 1;
    121: op1_11_inv24 = 1;
    122: op1_11_inv24 = 1;
    123: op1_11_inv24 = 1;
    127: op1_11_inv24 = 1;
    130: op1_11_inv24 = 1;
    default: op1_11_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in25 = reg_0439;
    53: op1_11_in25 = reg_0069;
    55: op1_11_in25 = reg_0836;
    73: op1_11_in25 = reg_0828;
    86: op1_11_in25 = reg_0319;
    74: op1_11_in25 = reg_0047;
    69: op1_11_in25 = reg_0837;
    54: op1_11_in25 = reg_1145;
    75: op1_11_in25 = reg_0393;
    50: op1_11_in25 = reg_0391;
    68: op1_11_in25 = reg_0885;
    76: op1_11_in25 = reg_0707;
    71: op1_11_in25 = reg_0548;
    111: op1_11_in25 = reg_0548;
    87: op1_11_in25 = reg_0566;
    77: op1_11_in25 = reg_0461;
    61: op1_11_in25 = reg_0966;
    58: op1_11_in25 = reg_0197;
    78: op1_11_in25 = reg_0553;
    70: op1_11_in25 = reg_0756;
    79: op1_11_in25 = reg_0609;
    117: op1_11_in25 = reg_0609;
    51: op1_11_in25 = reg_0867;
    59: op1_11_in25 = reg_0747;
    88: op1_11_in25 = reg_1280;
    80: op1_11_in25 = reg_0396;
    62: op1_11_in25 = reg_0727;
    81: op1_11_in25 = reg_1256;
    46: op1_11_in25 = reg_0827;
    93: op1_11_in25 = reg_0827;
    52: op1_11_in25 = reg_0376;
    63: op1_11_in25 = reg_0327;
    82: op1_11_in25 = reg_0820;
    89: op1_11_in25 = reg_0096;
    83: op1_11_in25 = reg_1473;
    64: op1_11_in25 = reg_0131;
    84: op1_11_in25 = reg_0463;
    48: op1_11_in25 = reg_0325;
    85: op1_11_in25 = reg_0277;
    65: op1_11_in25 = reg_0436;
    90: op1_11_in25 = reg_0564;
    66: op1_11_in25 = reg_0334;
    91: op1_11_in25 = reg_1513;
    67: op1_11_in25 = reg_0190;
    92: op1_11_in25 = reg_0289;
    94: op1_11_in25 = reg_0414;
    95: op1_11_in25 = reg_1098;
    96: op1_11_in25 = reg_0996;
    97: op1_11_in25 = reg_0601;
    98: op1_11_in25 = reg_0139;
    99: op1_11_in25 = reg_0469;
    100: op1_11_in25 = reg_0925;
    101: op1_11_in25 = reg_1078;
    102: op1_11_in25 = reg_0373;
    104: op1_11_in25 = reg_0967;
    105: op1_11_in25 = reg_1018;
    106: op1_11_in25 = reg_0538;
    47: op1_11_in25 = reg_0541;
    107: op1_11_in25 = reg_0921;
    108: op1_11_in25 = reg_0595;
    110: op1_11_in25 = reg_0264;
    112: op1_11_in25 = reg_1517;
    113: op1_11_in25 = reg_0260;
    114: op1_11_in25 = reg_0571;
    115: op1_11_in25 = reg_0222;
    116: op1_11_in25 = reg_0792;
    118: op1_11_in25 = reg_0963;
    119: op1_11_in25 = reg_0452;
    120: op1_11_in25 = reg_0719;
    121: op1_11_in25 = reg_0246;
    122: op1_11_in25 = reg_1401;
    123: op1_11_in25 = reg_0043;
    125: op1_11_in25 = imem03_in[7:4];
    44: op1_11_in25 = reg_0151;
    126: op1_11_in25 = reg_1056;
    129: op1_11_in25 = reg_1056;
    127: op1_11_in25 = reg_0392;
    128: op1_11_in25 = reg_0939;
    130: op1_11_in25 = reg_1518;
    131: op1_11_in25 = reg_0457;
    default: op1_11_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv25 = 1;
    53: op1_11_inv25 = 1;
    86: op1_11_inv25 = 1;
    69: op1_11_inv25 = 1;
    75: op1_11_inv25 = 1;
    71: op1_11_inv25 = 1;
    61: op1_11_inv25 = 1;
    79: op1_11_inv25 = 1;
    51: op1_11_inv25 = 1;
    59: op1_11_inv25 = 1;
    63: op1_11_inv25 = 1;
    89: op1_11_inv25 = 1;
    83: op1_11_inv25 = 1;
    84: op1_11_inv25 = 1;
    65: op1_11_inv25 = 1;
    66: op1_11_inv25 = 1;
    67: op1_11_inv25 = 1;
    92: op1_11_inv25 = 1;
    94: op1_11_inv25 = 1;
    95: op1_11_inv25 = 1;
    97: op1_11_inv25 = 1;
    100: op1_11_inv25 = 1;
    102: op1_11_inv25 = 1;
    104: op1_11_inv25 = 1;
    107: op1_11_inv25 = 1;
    111: op1_11_inv25 = 1;
    112: op1_11_inv25 = 1;
    115: op1_11_inv25 = 1;
    119: op1_11_inv25 = 1;
    125: op1_11_inv25 = 1;
    44: op1_11_inv25 = 1;
    126: op1_11_inv25 = 1;
    127: op1_11_inv25 = 1;
    128: op1_11_inv25 = 1;
    129: op1_11_inv25 = 1;
    131: op1_11_inv25 = 1;
    default: op1_11_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in26 = reg_0146;
    53: op1_11_in26 = reg_0325;
    55: op1_11_in26 = reg_0338;
    73: op1_11_in26 = reg_0040;
    86: op1_11_in26 = reg_0368;
    74: op1_11_in26 = reg_0093;
    78: op1_11_in26 = reg_0093;
    69: op1_11_in26 = reg_0719;
    54: op1_11_in26 = reg_0600;
    75: op1_11_in26 = reg_0797;
    50: op1_11_in26 = reg_0457;
    68: op1_11_in26 = reg_0505;
    76: op1_11_in26 = reg_0049;
    71: op1_11_in26 = reg_0868;
    87: op1_11_in26 = reg_0303;
    128: op1_11_in26 = reg_0303;
    77: op1_11_in26 = reg_1315;
    61: op1_11_in26 = reg_0968;
    58: op1_11_in26 = reg_0184;
    70: op1_11_in26 = reg_0732;
    79: op1_11_in26 = reg_0742;
    82: op1_11_in26 = reg_0742;
    51: op1_11_in26 = reg_0297;
    59: op1_11_in26 = reg_0259;
    88: op1_11_in26 = reg_0426;
    80: op1_11_in26 = reg_1147;
    62: op1_11_in26 = reg_0360;
    81: op1_11_in26 = reg_0277;
    46: op1_11_in26 = reg_0718;
    52: op1_11_in26 = reg_0697;
    63: op1_11_in26 = reg_0830;
    89: op1_11_in26 = reg_1503;
    83: op1_11_in26 = reg_1474;
    64: op1_11_in26 = reg_0745;
    84: op1_11_in26 = reg_0548;
    48: op1_11_in26 = reg_0216;
    85: op1_11_in26 = reg_0785;
    65: op1_11_in26 = reg_0934;
    90: op1_11_in26 = reg_1180;
    66: op1_11_in26 = reg_1181;
    91: op1_11_in26 = reg_0553;
    67: op1_11_in26 = reg_0558;
    130: op1_11_in26 = reg_0558;
    92: op1_11_in26 = reg_0244;
    93: op1_11_in26 = reg_0109;
    94: op1_11_in26 = reg_0407;
    95: op1_11_in26 = reg_0007;
    96: op1_11_in26 = reg_0831;
    97: op1_11_in26 = reg_0243;
    98: op1_11_in26 = reg_0779;
    99: op1_11_in26 = reg_0572;
    100: op1_11_in26 = reg_0316;
    101: op1_11_in26 = reg_0069;
    102: op1_11_in26 = reg_0622;
    104: op1_11_in26 = reg_0434;
    105: op1_11_in26 = reg_1260;
    106: op1_11_in26 = imem05_in[3:0];
    47: op1_11_in26 = reg_0450;
    107: op1_11_in26 = reg_0441;
    108: op1_11_in26 = reg_0403;
    110: op1_11_in26 = reg_0034;
    111: op1_11_in26 = reg_0747;
    112: op1_11_in26 = reg_1199;
    113: op1_11_in26 = reg_0238;
    114: op1_11_in26 = reg_1228;
    115: op1_11_in26 = reg_0260;
    116: op1_11_in26 = reg_0266;
    117: op1_11_in26 = reg_1473;
    118: op1_11_in26 = imem03_in[3:0];
    119: op1_11_in26 = reg_0232;
    120: op1_11_in26 = reg_0256;
    121: op1_11_in26 = reg_0051;
    122: op1_11_in26 = reg_1404;
    123: op1_11_in26 = reg_0166;
    125: op1_11_in26 = reg_0190;
    44: op1_11_in26 = reg_0861;
    126: op1_11_in26 = reg_1440;
    127: op1_11_in26 = reg_0491;
    129: op1_11_in26 = reg_1350;
    131: op1_11_in26 = reg_0923;
    default: op1_11_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv26 = 1;
    86: op1_11_inv26 = 1;
    69: op1_11_inv26 = 1;
    54: op1_11_inv26 = 1;
    71: op1_11_inv26 = 1;
    58: op1_11_inv26 = 1;
    78: op1_11_inv26 = 1;
    70: op1_11_inv26 = 1;
    79: op1_11_inv26 = 1;
    51: op1_11_inv26 = 1;
    88: op1_11_inv26 = 1;
    52: op1_11_inv26 = 1;
    63: op1_11_inv26 = 1;
    82: op1_11_inv26 = 1;
    64: op1_11_inv26 = 1;
    84: op1_11_inv26 = 1;
    90: op1_11_inv26 = 1;
    67: op1_11_inv26 = 1;
    92: op1_11_inv26 = 1;
    93: op1_11_inv26 = 1;
    94: op1_11_inv26 = 1;
    99: op1_11_inv26 = 1;
    100: op1_11_inv26 = 1;
    104: op1_11_inv26 = 1;
    105: op1_11_inv26 = 1;
    106: op1_11_inv26 = 1;
    107: op1_11_inv26 = 1;
    110: op1_11_inv26 = 1;
    115: op1_11_inv26 = 1;
    116: op1_11_inv26 = 1;
    118: op1_11_inv26 = 1;
    120: op1_11_inv26 = 1;
    121: op1_11_inv26 = 1;
    123: op1_11_inv26 = 1;
    125: op1_11_inv26 = 1;
    126: op1_11_inv26 = 1;
    127: op1_11_inv26 = 1;
    128: op1_11_inv26 = 1;
    129: op1_11_inv26 = 1;
    130: op1_11_inv26 = 1;
    131: op1_11_inv26 = 1;
    default: op1_11_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in27 = reg_0091;
    53: op1_11_in27 = reg_0311;
    55: op1_11_in27 = reg_0061;
    73: op1_11_in27 = reg_0399;
    86: op1_11_in27 = reg_0719;
    74: op1_11_in27 = imem01_in[7:4];
    69: op1_11_in27 = reg_0337;
    54: op1_11_in27 = reg_0185;
    75: op1_11_in27 = reg_0151;
    50: op1_11_in27 = reg_0230;
    68: op1_11_in27 = reg_0480;
    76: op1_11_in27 = reg_0704;
    71: op1_11_in27 = reg_0331;
    87: op1_11_in27 = reg_0090;
    77: op1_11_in27 = reg_0667;
    61: op1_11_in27 = reg_0819;
    58: op1_11_in27 = reg_0130;
    78: op1_11_in27 = reg_0550;
    70: op1_11_in27 = reg_0678;
    79: op1_11_in27 = reg_1474;
    82: op1_11_in27 = reg_1474;
    117: op1_11_in27 = reg_1474;
    51: op1_11_in27 = reg_0169;
    59: op1_11_in27 = reg_0728;
    88: op1_11_in27 = reg_0443;
    80: op1_11_in27 = reg_0421;
    62: op1_11_in27 = reg_0047;
    81: op1_11_in27 = reg_1512;
    85: op1_11_in27 = reg_1512;
    46: op1_11_in27 = reg_0670;
    52: op1_11_in27 = reg_0698;
    63: op1_11_in27 = reg_0279;
    89: op1_11_in27 = reg_0016;
    83: op1_11_in27 = reg_0402;
    64: op1_11_in27 = reg_0541;
    84: op1_11_in27 = reg_0747;
    48: op1_11_in27 = reg_0709;
    65: op1_11_in27 = reg_0128;
    90: op1_11_in27 = reg_0301;
    66: op1_11_in27 = reg_0938;
    91: op1_11_in27 = reg_0547;
    67: op1_11_in27 = reg_1093;
    92: op1_11_in27 = reg_1202;
    93: op1_11_in27 = reg_0716;
    94: op1_11_in27 = reg_0599;
    95: op1_11_in27 = reg_1078;
    96: op1_11_in27 = reg_0391;
    97: op1_11_in27 = reg_0240;
    98: op1_11_in27 = reg_0775;
    99: op1_11_in27 = reg_0966;
    100: op1_11_in27 = reg_0974;
    101: op1_11_in27 = reg_0009;
    102: op1_11_in27 = reg_0619;
    104: op1_11_in27 = reg_0290;
    105: op1_11_in27 = reg_0495;
    106: op1_11_in27 = reg_0833;
    47: op1_11_in27 = reg_0895;
    107: op1_11_in27 = reg_0739;
    108: op1_11_in27 = reg_1493;
    110: op1_11_in27 = reg_0164;
    111: op1_11_in27 = reg_0610;
    112: op1_11_in27 = reg_0108;
    113: op1_11_in27 = reg_0798;
    114: op1_11_in27 = reg_0171;
    115: op1_11_in27 = reg_0830;
    116: op1_11_in27 = reg_1163;
    118: op1_11_in27 = imem03_in[7:4];
    119: op1_11_in27 = reg_0862;
    120: op1_11_in27 = reg_0236;
    121: op1_11_in27 = reg_0668;
    122: op1_11_in27 = reg_0939;
    123: op1_11_in27 = reg_1071;
    125: op1_11_in27 = reg_0732;
    44: op1_11_in27 = reg_0038;
    126: op1_11_in27 = reg_0140;
    127: op1_11_in27 = reg_0182;
    128: op1_11_in27 = reg_0302;
    129: op1_11_in27 = reg_0159;
    130: op1_11_in27 = reg_0884;
    131: op1_11_in27 = reg_0223;
    default: op1_11_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv27 = 1;
    53: op1_11_inv27 = 1;
    55: op1_11_inv27 = 1;
    73: op1_11_inv27 = 1;
    74: op1_11_inv27 = 1;
    69: op1_11_inv27 = 1;
    54: op1_11_inv27 = 1;
    68: op1_11_inv27 = 1;
    71: op1_11_inv27 = 1;
    77: op1_11_inv27 = 1;
    61: op1_11_inv27 = 1;
    78: op1_11_inv27 = 1;
    70: op1_11_inv27 = 1;
    59: op1_11_inv27 = 1;
    88: op1_11_inv27 = 1;
    62: op1_11_inv27 = 1;
    63: op1_11_inv27 = 1;
    82: op1_11_inv27 = 1;
    89: op1_11_inv27 = 1;
    64: op1_11_inv27 = 1;
    84: op1_11_inv27 = 1;
    48: op1_11_inv27 = 1;
    85: op1_11_inv27 = 1;
    65: op1_11_inv27 = 1;
    91: op1_11_inv27 = 1;
    67: op1_11_inv27 = 1;
    92: op1_11_inv27 = 1;
    93: op1_11_inv27 = 1;
    94: op1_11_inv27 = 1;
    98: op1_11_inv27 = 1;
    99: op1_11_inv27 = 1;
    104: op1_11_inv27 = 1;
    106: op1_11_inv27 = 1;
    108: op1_11_inv27 = 1;
    110: op1_11_inv27 = 1;
    113: op1_11_inv27 = 1;
    114: op1_11_inv27 = 1;
    115: op1_11_inv27 = 1;
    116: op1_11_inv27 = 1;
    117: op1_11_inv27 = 1;
    118: op1_11_inv27 = 1;
    119: op1_11_inv27 = 1;
    121: op1_11_inv27 = 1;
    122: op1_11_inv27 = 1;
    123: op1_11_inv27 = 1;
    44: op1_11_inv27 = 1;
    128: op1_11_inv27 = 1;
    130: op1_11_inv27 = 1;
    default: op1_11_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in28 = reg_0724;
    53: op1_11_in28 = reg_1092;
    55: op1_11_in28 = reg_0020;
    73: op1_11_in28 = reg_1436;
    86: op1_11_in28 = reg_0337;
    74: op1_11_in28 = reg_0968;
    69: op1_11_in28 = reg_0094;
    54: op1_11_in28 = reg_0179;
    75: op1_11_in28 = reg_0861;
    50: op1_11_in28 = imem07_in[3:0];
    68: op1_11_in28 = imem03_in[7:4];
    76: op1_11_in28 = reg_0378;
    71: op1_11_in28 = reg_0420;
    87: op1_11_in28 = reg_1373;
    77: op1_11_in28 = reg_0892;
    61: op1_11_in28 = reg_0434;
    82: op1_11_in28 = reg_0434;
    99: op1_11_in28 = reg_0434;
    58: op1_11_in28 = reg_0118;
    78: op1_11_in28 = reg_0787;
    70: op1_11_in28 = reg_0709;
    79: op1_11_in28 = reg_0572;
    51: op1_11_in28 = reg_0140;
    59: op1_11_in28 = reg_0402;
    88: op1_11_in28 = reg_0341;
    80: op1_11_in28 = reg_0969;
    62: op1_11_in28 = reg_0899;
    81: op1_11_in28 = reg_0093;
    46: op1_11_in28 = reg_0634;
    52: op1_11_in28 = reg_0699;
    63: op1_11_in28 = reg_1132;
    89: op1_11_in28 = reg_0021;
    83: op1_11_in28 = reg_0595;
    64: op1_11_in28 = reg_0070;
    84: op1_11_in28 = reg_0222;
    111: op1_11_in28 = reg_0222;
    48: op1_11_in28 = reg_0376;
    85: op1_11_in28 = reg_0331;
    65: op1_11_in28 = reg_0705;
    90: op1_11_in28 = reg_1484;
    66: op1_11_in28 = reg_0477;
    91: op1_11_in28 = reg_0549;
    67: op1_11_in28 = reg_0885;
    92: op1_11_in28 = reg_0022;
    93: op1_11_in28 = reg_0717;
    94: op1_11_in28 = reg_0454;
    95: op1_11_in28 = reg_0069;
    96: op1_11_in28 = reg_0045;
    97: op1_11_in28 = reg_1348;
    98: op1_11_in28 = reg_0465;
    126: op1_11_in28 = reg_0465;
    100: op1_11_in28 = reg_0751;
    101: op1_11_in28 = reg_0255;
    102: op1_11_in28 = reg_0571;
    104: op1_11_in28 = reg_0365;
    105: op1_11_in28 = reg_0436;
    106: op1_11_in28 = reg_0332;
    47: op1_11_in28 = reg_0168;
    107: op1_11_in28 = reg_0738;
    108: op1_11_in28 = reg_0822;
    110: op1_11_in28 = reg_1258;
    112: op1_11_in28 = reg_0104;
    113: op1_11_in28 = reg_0742;
    114: op1_11_in28 = reg_0419;
    115: op1_11_in28 = reg_0798;
    116: op1_11_in28 = reg_0736;
    117: op1_11_in28 = reg_1452;
    118: op1_11_in28 = imem03_in[11:8];
    119: op1_11_in28 = reg_0836;
    120: op1_11_in28 = reg_0904;
    121: op1_11_in28 = reg_1183;
    122: op1_11_in28 = reg_0302;
    123: op1_11_in28 = reg_0626;
    125: op1_11_in28 = reg_0049;
    44: op1_11_in28 = reg_0195;
    127: op1_11_in28 = reg_0266;
    128: op1_11_in28 = reg_0794;
    129: op1_11_in28 = reg_0779;
    130: op1_11_in28 = reg_0218;
    131: op1_11_in28 = reg_0441;
    default: op1_11_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_11_inv28 = 1;
    86: op1_11_inv28 = 1;
    69: op1_11_inv28 = 1;
    54: op1_11_inv28 = 1;
    75: op1_11_inv28 = 1;
    71: op1_11_inv28 = 1;
    77: op1_11_inv28 = 1;
    58: op1_11_inv28 = 1;
    70: op1_11_inv28 = 1;
    79: op1_11_inv28 = 1;
    88: op1_11_inv28 = 1;
    80: op1_11_inv28 = 1;
    81: op1_11_inv28 = 1;
    52: op1_11_inv28 = 1;
    83: op1_11_inv28 = 1;
    48: op1_11_inv28 = 1;
    85: op1_11_inv28 = 1;
    65: op1_11_inv28 = 1;
    90: op1_11_inv28 = 1;
    66: op1_11_inv28 = 1;
    93: op1_11_inv28 = 1;
    97: op1_11_inv28 = 1;
    99: op1_11_inv28 = 1;
    100: op1_11_inv28 = 1;
    102: op1_11_inv28 = 1;
    105: op1_11_inv28 = 1;
    106: op1_11_inv28 = 1;
    47: op1_11_inv28 = 1;
    107: op1_11_inv28 = 1;
    108: op1_11_inv28 = 1;
    112: op1_11_inv28 = 1;
    115: op1_11_inv28 = 1;
    117: op1_11_inv28 = 1;
    118: op1_11_inv28 = 1;
    119: op1_11_inv28 = 1;
    123: op1_11_inv28 = 1;
    125: op1_11_inv28 = 1;
    126: op1_11_inv28 = 1;
    127: op1_11_inv28 = 1;
    129: op1_11_inv28 = 1;
    default: op1_11_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in29 = reg_0282;
    53: op1_11_in29 = reg_1093;
    55: op1_11_in29 = reg_0793;
    73: op1_11_in29 = reg_0730;
    86: op1_11_in29 = reg_1151;
    74: op1_11_in29 = reg_0384;
    69: op1_11_in29 = reg_0236;
    54: op1_11_in29 = reg_1003;
    75: op1_11_in29 = reg_0039;
    50: op1_11_in29 = imem07_in[15:12];
    68: op1_11_in29 = reg_0849;
    76: op1_11_in29 = reg_1325;
    71: op1_11_in29 = reg_0468;
    87: op1_11_in29 = reg_0196;
    47: op1_11_in29 = reg_0196;
    77: op1_11_in29 = reg_0674;
    61: op1_11_in29 = reg_0401;
    58: op1_11_in29 = reg_0240;
    78: op1_11_in29 = reg_0439;
    70: op1_11_in29 = reg_0185;
    79: op1_11_in29 = reg_0434;
    51: op1_11_in29 = reg_0740;
    59: op1_11_in29 = reg_0386;
    88: op1_11_in29 = reg_0208;
    80: op1_11_in29 = reg_1233;
    62: op1_11_in29 = reg_0077;
    81: op1_11_in29 = reg_0463;
    46: op1_11_in29 = reg_0419;
    52: op1_11_in29 = reg_0600;
    63: op1_11_in29 = reg_0732;
    82: op1_11_in29 = reg_0148;
    99: op1_11_in29 = reg_0148;
    113: op1_11_in29 = reg_0148;
    117: op1_11_in29 = reg_0148;
    89: op1_11_in29 = imem05_in[11:8];
    83: op1_11_in29 = reg_0874;
    64: op1_11_in29 = imem05_in[15:12];
    84: op1_11_in29 = reg_0609;
    48: op1_11_in29 = reg_0348;
    85: op1_11_in29 = reg_0787;
    65: op1_11_in29 = reg_0845;
    90: op1_11_in29 = reg_0576;
    66: op1_11_in29 = reg_0274;
    91: op1_11_in29 = reg_0746;
    67: op1_11_in29 = reg_0880;
    92: op1_11_in29 = imem07_in[11:8];
    93: op1_11_in29 = reg_0373;
    94: op1_11_in29 = reg_0061;
    95: op1_11_in29 = reg_0168;
    96: op1_11_in29 = reg_0938;
    97: op1_11_in29 = reg_1346;
    98: op1_11_in29 = reg_0739;
    100: op1_11_in29 = reg_0827;
    101: op1_11_in29 = reg_0563;
    102: op1_11_in29 = reg_0345;
    104: op1_11_in29 = reg_0175;
    105: op1_11_in29 = reg_0054;
    106: op1_11_in29 = reg_0278;
    107: op1_11_in29 = reg_0593;
    108: op1_11_in29 = reg_1260;
    110: op1_11_in29 = reg_0531;
    111: op1_11_in29 = reg_0241;
    112: op1_11_in29 = reg_0707;
    114: op1_11_in29 = reg_0067;
    115: op1_11_in29 = reg_0966;
    116: op1_11_in29 = reg_0450;
    128: op1_11_in29 = reg_0450;
    118: op1_11_in29 = reg_0049;
    119: op1_11_in29 = reg_1312;
    120: op1_11_in29 = reg_0117;
    121: op1_11_in29 = reg_0922;
    122: op1_11_in29 = reg_0873;
    123: op1_11_in29 = reg_0606;
    125: op1_11_in29 = reg_0444;
    44: op1_11_in29 = reg_0192;
    126: op1_11_in29 = reg_0665;
    127: op1_11_in29 = reg_0302;
    129: op1_11_in29 = reg_0415;
    130: op1_11_in29 = reg_0313;
    131: op1_11_in29 = reg_0413;
    default: op1_11_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_11_inv29 = 1;
    53: op1_11_inv29 = 1;
    55: op1_11_inv29 = 1;
    73: op1_11_inv29 = 1;
    86: op1_11_inv29 = 1;
    69: op1_11_inv29 = 1;
    54: op1_11_inv29 = 1;
    50: op1_11_inv29 = 1;
    68: op1_11_inv29 = 1;
    76: op1_11_inv29 = 1;
    71: op1_11_inv29 = 1;
    61: op1_11_inv29 = 1;
    70: op1_11_inv29 = 1;
    88: op1_11_inv29 = 1;
    62: op1_11_inv29 = 1;
    81: op1_11_inv29 = 1;
    52: op1_11_inv29 = 1;
    85: op1_11_inv29 = 1;
    65: op1_11_inv29 = 1;
    90: op1_11_inv29 = 1;
    66: op1_11_inv29 = 1;
    91: op1_11_inv29 = 1;
    92: op1_11_inv29 = 1;
    93: op1_11_inv29 = 1;
    94: op1_11_inv29 = 1;
    95: op1_11_inv29 = 1;
    98: op1_11_inv29 = 1;
    99: op1_11_inv29 = 1;
    100: op1_11_inv29 = 1;
    102: op1_11_inv29 = 1;
    106: op1_11_inv29 = 1;
    47: op1_11_inv29 = 1;
    108: op1_11_inv29 = 1;
    110: op1_11_inv29 = 1;
    111: op1_11_inv29 = 1;
    117: op1_11_inv29 = 1;
    119: op1_11_inv29 = 1;
    120: op1_11_inv29 = 1;
    122: op1_11_inv29 = 1;
    44: op1_11_inv29 = 1;
    126: op1_11_inv29 = 1;
    128: op1_11_inv29 = 1;
    129: op1_11_inv29 = 1;
    default: op1_11_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_11_in30 = reg_0012;
    53: op1_11_in30 = reg_0706;
    55: op1_11_in30 = reg_0578;
    73: op1_11_in30 = reg_1323;
    86: op1_11_in30 = reg_0096;
    74: op1_11_in30 = reg_0386;
    69: op1_11_in30 = reg_0065;
    54: op1_11_in30 = reg_0220;
    75: op1_11_in30 = reg_0751;
    50: op1_11_in30 = reg_0998;
    68: op1_11_in30 = reg_1282;
    76: op1_11_in30 = reg_0145;
    71: op1_11_in30 = reg_0966;
    87: op1_11_in30 = reg_0240;
    77: op1_11_in30 = reg_0187;
    61: op1_11_in30 = reg_0093;
    58: op1_11_in30 = reg_0040;
    78: op1_11_in30 = reg_0438;
    70: op1_11_in30 = reg_0378;
    79: op1_11_in30 = reg_1457;
    51: op1_11_in30 = reg_0137;
    59: op1_11_in30 = reg_0385;
    88: op1_11_in30 = reg_0264;
    80: op1_11_in30 = reg_0342;
    62: op1_11_in30 = reg_0277;
    81: op1_11_in30 = reg_0239;
    46: op1_11_in30 = reg_0046;
    52: op1_11_in30 = reg_0178;
    63: op1_11_in30 = reg_0678;
    82: op1_11_in30 = reg_0384;
    89: op1_11_in30 = reg_0737;
    83: op1_11_in30 = reg_0291;
    64: op1_11_in30 = reg_0130;
    66: op1_11_in30 = reg_0130;
    47: op1_11_in30 = reg_0130;
    116: op1_11_in30 = reg_0130;
    84: op1_11_in30 = reg_0830;
    48: op1_11_in30 = reg_0790;
    85: op1_11_in30 = reg_0743;
    65: op1_11_in30 = imem02_in[7:4];
    90: op1_11_in30 = reg_0492;
    91: op1_11_in30 = reg_0222;
    67: op1_11_in30 = reg_0506;
    92: op1_11_in30 = reg_0675;
    93: op1_11_in30 = reg_0624;
    94: op1_11_in30 = reg_0369;
    95: op1_11_in30 = reg_0632;
    96: op1_11_in30 = reg_0450;
    97: op1_11_in30 = reg_0603;
    98: op1_11_in30 = reg_0103;
    99: op1_11_in30 = reg_0146;
    117: op1_11_in30 = reg_0146;
    100: op1_11_in30 = reg_1504;
    101: op1_11_in30 = reg_1515;
    102: op1_11_in30 = reg_0296;
    104: op1_11_in30 = reg_0335;
    105: op1_11_in30 = reg_0326;
    106: op1_11_in30 = reg_1164;
    107: op1_11_in30 = reg_0114;
    108: op1_11_in30 = reg_0495;
    110: op1_11_in30 = reg_0281;
    111: op1_11_in30 = reg_0820;
    112: op1_11_in30 = reg_0673;
    130: op1_11_in30 = reg_0673;
    113: op1_11_in30 = reg_0290;
    114: op1_11_in30 = reg_1170;
    115: op1_11_in30 = reg_0149;
    118: op1_11_in30 = reg_1003;
    119: op1_11_in30 = reg_0932;
    120: op1_11_in30 = reg_0536;
    121: op1_11_in30 = reg_1056;
    122: op1_11_in30 = reg_0197;
    123: op1_11_in30 = reg_0846;
    125: op1_11_in30 = reg_0330;
    44: op1_11_in30 = imem06_in[11:8];
    126: op1_11_in30 = reg_0663;
    127: op1_11_in30 = reg_0301;
    128: op1_11_in30 = reg_0274;
    129: op1_11_in30 = reg_0621;
    131: op1_11_in30 = reg_0593;
    default: op1_11_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_11_inv30 = 1;
    86: op1_11_inv30 = 1;
    74: op1_11_inv30 = 1;
    50: op1_11_inv30 = 1;
    71: op1_11_inv30 = 1;
    61: op1_11_inv30 = 1;
    78: op1_11_inv30 = 1;
    59: op1_11_inv30 = 1;
    62: op1_11_inv30 = 1;
    46: op1_11_inv30 = 1;
    52: op1_11_inv30 = 1;
    89: op1_11_inv30 = 1;
    64: op1_11_inv30 = 1;
    84: op1_11_inv30 = 1;
    48: op1_11_inv30 = 1;
    85: op1_11_inv30 = 1;
    67: op1_11_inv30 = 1;
    92: op1_11_inv30 = 1;
    98: op1_11_inv30 = 1;
    99: op1_11_inv30 = 1;
    100: op1_11_inv30 = 1;
    101: op1_11_inv30 = 1;
    104: op1_11_inv30 = 1;
    105: op1_11_inv30 = 1;
    106: op1_11_inv30 = 1;
    47: op1_11_inv30 = 1;
    113: op1_11_inv30 = 1;
    115: op1_11_inv30 = 1;
    116: op1_11_inv30 = 1;
    118: op1_11_inv30 = 1;
    121: op1_11_inv30 = 1;
    123: op1_11_inv30 = 1;
    125: op1_11_inv30 = 1;
    127: op1_11_inv30 = 1;
    129: op1_11_inv30 = 1;
    130: op1_11_inv30 = 1;
    131: op1_11_inv30 = 1;
    default: op1_11_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_11_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#11の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_11_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in00 = reg_0303;
    53: op1_12_in00 = imem01_in[7:4];
    55: op1_12_in00 = reg_0973;
    73: op1_12_in00 = reg_0129;
    86: op1_12_in00 = reg_0007;
    74: op1_12_in00 = reg_0615;
    69: op1_12_in00 = reg_0291;
    49: op1_12_in00 = reg_0752;
    54: op1_12_in00 = reg_0466;
    75: op1_12_in00 = reg_1105;
    56: op1_12_in00 = reg_0093;
    50: op1_12_in00 = reg_0116;
    76: op1_12_in00 = reg_0735;
    68: op1_12_in00 = reg_0789;
    71: op1_12_in00 = reg_0843;
    124: op1_12_in00 = reg_0843;
    87: op1_12_in00 = reg_0495;
    88: op1_12_in00 = reg_0495;
    57: op1_12_in00 = reg_0120;
    77: op1_12_in00 = reg_0799;
    61: op1_12_in00 = reg_0555;
    58: op1_12_in00 = reg_0044;
    78: op1_12_in00 = reg_0048;
    70: op1_12_in00 = reg_0145;
    59: op1_12_in00 = reg_0365;
    79: op1_12_in00 = reg_0905;
    51: op1_12_in00 = reg_0438;
    60: op1_12_in00 = reg_0445;
    80: op1_12_in00 = reg_1080;
    62: op1_12_in00 = reg_0391;
    81: op1_12_in00 = reg_0390;
    52: op1_12_in00 = reg_0207;
    63: op1_12_in00 = reg_0337;
    82: op1_12_in00 = reg_0368;
    46: op1_12_in00 = reg_0469;
    83: op1_12_in00 = reg_0983;
    64: op1_12_in00 = reg_0613;
    89: op1_12_in00 = reg_1199;
    84: op1_12_in00 = reg_0236;
    85: op1_12_in00 = reg_1091;
    65: op1_12_in00 = reg_0783;
    90: op1_12_in00 = reg_1448;
    48: op1_12_in00 = reg_0147;
    66: op1_12_in00 = reg_0929;
    91: op1_12_in00 = reg_0715;
    67: op1_12_in00 = reg_0371;
    92: op1_12_in00 = imem00_in[11:8];
    33: op1_12_in00 = imem07_in[3:0];
    93: op1_12_in00 = reg_0323;
    94: op1_12_in00 = reg_0698;
    47: op1_12_in00 = reg_0698;
    28: op1_12_in00 = reg_0228;
    95: op1_12_in00 = imem03_in[11:8];
    96: op1_12_in00 = reg_1514;
    97: op1_12_in00 = reg_0861;
    98: op1_12_in00 = reg_0100;
    99: op1_12_in00 = reg_0363;
    117: op1_12_in00 = reg_0363;
    100: op1_12_in00 = reg_0172;
    130: op1_12_in00 = reg_0172;
    101: op1_12_in00 = imem03_in[3:0];
    102: op1_12_in00 = reg_0308;
    37: op1_12_in00 = reg_0442;
    103: op1_12_in00 = reg_0121;
    104: op1_12_in00 = reg_0080;
    105: op1_12_in00 = reg_0778;
    106: op1_12_in00 = reg_0992;
    107: op1_12_in00 = reg_0028;
    108: op1_12_in00 = reg_0970;
    109: op1_12_in00 = reg_1243;
    110: op1_12_in00 = reg_0407;
    111: op1_12_in00 = reg_0383;
    112: op1_12_in00 = reg_0348;
    113: op1_12_in00 = reg_0875;
    114: op1_12_in00 = reg_1057;
    115: op1_12_in00 = reg_0290;
    116: op1_12_in00 = reg_0243;
    118: op1_12_in00 = reg_0185;
    119: op1_12_in00 = reg_0420;
    120: op1_12_in00 = reg_0065;
    121: op1_12_in00 = reg_1345;
    122: op1_12_in00 = reg_0602;
    123: op1_12_in00 = reg_0423;
    125: op1_12_in00 = reg_1000;
    44: op1_12_in00 = reg_0797;
    126: op1_12_in00 = reg_0959;
    127: op1_12_in00 = reg_0873;
    128: op1_12_in00 = reg_0118;
    129: op1_12_in00 = reg_0958;
    38: op1_12_in00 = reg_0661;
    34: op1_12_in00 = reg_0620;
    default: op1_12_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_12_inv00 = 1;
    86: op1_12_inv00 = 1;
    74: op1_12_inv00 = 1;
    49: op1_12_inv00 = 1;
    50: op1_12_inv00 = 1;
    71: op1_12_inv00 = 1;
    59: op1_12_inv00 = 1;
    62: op1_12_inv00 = 1;
    52: op1_12_inv00 = 1;
    82: op1_12_inv00 = 1;
    46: op1_12_inv00 = 1;
    64: op1_12_inv00 = 1;
    65: op1_12_inv00 = 1;
    48: op1_12_inv00 = 1;
    92: op1_12_inv00 = 1;
    33: op1_12_inv00 = 1;
    93: op1_12_inv00 = 1;
    95: op1_12_inv00 = 1;
    96: op1_12_inv00 = 1;
    98: op1_12_inv00 = 1;
    100: op1_12_inv00 = 1;
    101: op1_12_inv00 = 1;
    109: op1_12_inv00 = 1;
    110: op1_12_inv00 = 1;
    113: op1_12_inv00 = 1;
    115: op1_12_inv00 = 1;
    117: op1_12_inv00 = 1;
    120: op1_12_inv00 = 1;
    121: op1_12_inv00 = 1;
    126: op1_12_inv00 = 1;
    127: op1_12_inv00 = 1;
    128: op1_12_inv00 = 1;
    38: op1_12_inv00 = 1;
    130: op1_12_inv00 = 1;
    default: op1_12_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in01 = reg_0492;
    53: op1_12_in01 = imem01_in[15:12];
    46: op1_12_in01 = imem01_in[15:12];
    55: op1_12_in01 = reg_0056;
    73: op1_12_in01 = reg_0630;
    86: op1_12_in01 = reg_0008;
    74: op1_12_in01 = reg_1243;
    69: op1_12_in01 = reg_0278;
    49: op1_12_in01 = reg_0194;
    54: op1_12_in01 = reg_0681;
    75: op1_12_in01 = reg_0377;
    56: op1_12_in01 = reg_0043;
    50: op1_12_in01 = reg_0717;
    100: op1_12_in01 = reg_0717;
    76: op1_12_in01 = reg_0205;
    68: op1_12_in01 = reg_0964;
    71: op1_12_in01 = reg_1244;
    92: op1_12_in01 = reg_1244;
    87: op1_12_in01 = reg_1451;
    57: op1_12_in01 = reg_0866;
    77: op1_12_in01 = reg_0797;
    61: op1_12_in01 = reg_0445;
    58: op1_12_in01 = reg_0662;
    78: op1_12_in01 = reg_0882;
    70: op1_12_in01 = reg_0180;
    59: op1_12_in01 = reg_0092;
    79: op1_12_in01 = reg_0925;
    51: op1_12_in01 = reg_0147;
    60: op1_12_in01 = reg_1277;
    88: op1_12_in01 = reg_0111;
    80: op1_12_in01 = reg_1490;
    62: op1_12_in01 = reg_0315;
    81: op1_12_in01 = reg_0666;
    52: op1_12_in01 = reg_0206;
    63: op1_12_in01 = reg_0097;
    82: op1_12_in01 = reg_0211;
    83: op1_12_in01 = reg_1278;
    64: op1_12_in01 = reg_0669;
    89: op1_12_in01 = reg_0884;
    84: op1_12_in01 = reg_1107;
    85: op1_12_in01 = reg_0069;
    65: op1_12_in01 = reg_0730;
    90: op1_12_in01 = reg_0965;
    48: op1_12_in01 = reg_0149;
    66: op1_12_in01 = reg_0268;
    91: op1_12_in01 = reg_0383;
    67: op1_12_in01 = reg_0152;
    33: op1_12_in01 = imem07_in[15:12];
    93: op1_12_in01 = reg_1202;
    94: op1_12_in01 = reg_0305;
    28: op1_12_in01 = reg_0219;
    95: op1_12_in01 = reg_0504;
    96: op1_12_in01 = reg_0300;
    97: op1_12_in01 = reg_1030;
    98: op1_12_in01 = reg_0003;
    99: op1_12_in01 = reg_0400;
    101: op1_12_in01 = imem03_in[11:8];
    102: op1_12_in01 = reg_0289;
    37: op1_12_in01 = imem07_in[11:8];
    103: op1_12_in01 = imem00_in[11:8];
    104: op1_12_in01 = reg_0078;
    105: op1_12_in01 = reg_0973;
    106: op1_12_in01 = reg_0491;
    47: op1_12_in01 = reg_0466;
    107: op1_12_in01 = reg_0050;
    108: op1_12_in01 = reg_1433;
    109: op1_12_in01 = reg_0248;
    110: op1_12_in01 = reg_0969;
    111: op1_12_in01 = reg_0335;
    112: op1_12_in01 = reg_0425;
    113: op1_12_in01 = reg_0403;
    114: op1_12_in01 = reg_0478;
    115: op1_12_in01 = reg_0385;
    116: op1_12_in01 = reg_0589;
    117: op1_12_in01 = reg_0901;
    118: op1_12_in01 = reg_0706;
    119: op1_12_in01 = reg_0210;
    120: op1_12_in01 = reg_1502;
    121: op1_12_in01 = reg_0159;
    122: op1_12_in01 = reg_0603;
    123: op1_12_in01 = reg_0561;
    124: op1_12_in01 = reg_1080;
    125: op1_12_in01 = reg_0597;
    44: op1_12_in01 = reg_0795;
    126: op1_12_in01 = reg_0841;
    127: op1_12_in01 = reg_0794;
    128: op1_12_in01 = reg_0799;
    129: op1_12_in01 = reg_0387;
    38: op1_12_in01 = reg_0663;
    130: op1_12_in01 = reg_0316;
    34: op1_12_in01 = reg_0593;
    default: op1_12_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv01 = 1;
    55: op1_12_inv01 = 1;
    74: op1_12_inv01 = 1;
    49: op1_12_inv01 = 1;
    54: op1_12_inv01 = 1;
    75: op1_12_inv01 = 1;
    50: op1_12_inv01 = 1;
    76: op1_12_inv01 = 1;
    68: op1_12_inv01 = 1;
    87: op1_12_inv01 = 1;
    57: op1_12_inv01 = 1;
    77: op1_12_inv01 = 1;
    61: op1_12_inv01 = 1;
    58: op1_12_inv01 = 1;
    60: op1_12_inv01 = 1;
    80: op1_12_inv01 = 1;
    81: op1_12_inv01 = 1;
    64: op1_12_inv01 = 1;
    89: op1_12_inv01 = 1;
    84: op1_12_inv01 = 1;
    85: op1_12_inv01 = 1;
    90: op1_12_inv01 = 1;
    48: op1_12_inv01 = 1;
    67: op1_12_inv01 = 1;
    92: op1_12_inv01 = 1;
    33: op1_12_inv01 = 1;
    28: op1_12_inv01 = 1;
    95: op1_12_inv01 = 1;
    96: op1_12_inv01 = 1;
    97: op1_12_inv01 = 1;
    98: op1_12_inv01 = 1;
    101: op1_12_inv01 = 1;
    103: op1_12_inv01 = 1;
    104: op1_12_inv01 = 1;
    105: op1_12_inv01 = 1;
    47: op1_12_inv01 = 1;
    110: op1_12_inv01 = 1;
    112: op1_12_inv01 = 1;
    117: op1_12_inv01 = 1;
    118: op1_12_inv01 = 1;
    119: op1_12_inv01 = 1;
    121: op1_12_inv01 = 1;
    122: op1_12_inv01 = 1;
    123: op1_12_inv01 = 1;
    126: op1_12_inv01 = 1;
    129: op1_12_inv01 = 1;
    130: op1_12_inv01 = 1;
    34: op1_12_inv01 = 1;
    default: op1_12_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in02 = reg_0601;
    53: op1_12_in02 = reg_0572;
    55: op1_12_in02 = reg_0055;
    73: op1_12_in02 = reg_0587;
    86: op1_12_in02 = reg_1392;
    74: op1_12_in02 = reg_0552;
    54: op1_12_in02 = reg_0552;
    69: op1_12_in02 = reg_0457;
    49: op1_12_in02 = reg_0866;
    75: op1_12_in02 = reg_0795;
    56: op1_12_in02 = reg_0011;
    50: op1_12_in02 = reg_0263;
    76: op1_12_in02 = reg_1299;
    68: op1_12_in02 = reg_0314;
    71: op1_12_in02 = imem00_in[15:12];
    87: op1_12_in02 = reg_1450;
    57: op1_12_in02 = reg_0397;
    77: op1_12_in02 = reg_0730;
    61: op1_12_in02 = reg_1241;
    58: op1_12_in02 = reg_0820;
    78: op1_12_in02 = reg_0884;
    70: op1_12_in02 = reg_0559;
    59: op1_12_in02 = reg_0868;
    79: op1_12_in02 = reg_0133;
    51: op1_12_in02 = reg_0400;
    60: op1_12_in02 = reg_1279;
    126: op1_12_in02 = reg_1279;
    88: op1_12_in02 = reg_0496;
    105: op1_12_in02 = reg_0496;
    80: op1_12_in02 = reg_1489;
    62: op1_12_in02 = reg_0737;
    81: op1_12_in02 = reg_1207;
    52: op1_12_in02 = reg_0014;
    63: op1_12_in02 = reg_0094;
    82: op1_12_in02 = reg_0536;
    66: op1_12_in02 = reg_0536;
    46: op1_12_in02 = reg_0434;
    83: op1_12_in02 = reg_1242;
    64: op1_12_in02 = reg_1281;
    109: op1_12_in02 = reg_1281;
    129: op1_12_in02 = reg_1281;
    89: op1_12_in02 = reg_1149;
    84: op1_12_in02 = reg_0420;
    85: op1_12_in02 = reg_0006;
    65: op1_12_in02 = reg_0160;
    90: op1_12_in02 = reg_0142;
    48: op1_12_in02 = reg_0402;
    91: op1_12_in02 = reg_0899;
    67: op1_12_in02 = reg_0185;
    92: op1_12_in02 = reg_0791;
    33: op1_12_in02 = reg_0050;
    93: op1_12_in02 = reg_1179;
    94: op1_12_in02 = reg_0835;
    28: op1_12_in02 = reg_0003;
    95: op1_12_in02 = reg_0328;
    96: op1_12_in02 = reg_0301;
    97: op1_12_in02 = reg_0960;
    98: op1_12_in02 = reg_0519;
    99: op1_12_in02 = reg_0403;
    100: op1_12_in02 = reg_0619;
    101: op1_12_in02 = imem03_in[15:12];
    102: op1_12_in02 = reg_0023;
    37: op1_12_in02 = reg_0408;
    103: op1_12_in02 = reg_0983;
    104: op1_12_in02 = reg_0728;
    106: op1_12_in02 = reg_0566;
    47: op1_12_in02 = reg_0676;
    107: op1_12_in02 = reg_0004;
    108: op1_12_in02 = reg_1140;
    110: op1_12_in02 = reg_0537;
    111: op1_12_in02 = reg_0724;
    115: op1_12_in02 = reg_0724;
    112: op1_12_in02 = reg_0336;
    113: op1_12_in02 = reg_0895;
    114: op1_12_in02 = reg_1060;
    116: op1_12_in02 = imem06_in[3:0];
    117: op1_12_in02 = reg_0595;
    118: op1_12_in02 = reg_1033;
    119: op1_12_in02 = reg_0038;
    120: op1_12_in02 = reg_0540;
    121: op1_12_in02 = reg_0489;
    122: op1_12_in02 = reg_0449;
    123: op1_12_in02 = reg_0497;
    124: op1_12_in02 = reg_0804;
    125: op1_12_in02 = reg_1425;
    44: op1_12_in02 = reg_0599;
    127: op1_12_in02 = imem05_in[11:8];
    128: op1_12_in02 = reg_0317;
    38: op1_12_in02 = reg_0442;
    130: op1_12_in02 = reg_0212;
    34: op1_12_in02 = reg_0592;
    default: op1_12_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv02 = 1;
    53: op1_12_inv02 = 1;
    55: op1_12_inv02 = 1;
    69: op1_12_inv02 = 1;
    49: op1_12_inv02 = 1;
    54: op1_12_inv02 = 1;
    75: op1_12_inv02 = 1;
    68: op1_12_inv02 = 1;
    87: op1_12_inv02 = 1;
    57: op1_12_inv02 = 1;
    58: op1_12_inv02 = 1;
    70: op1_12_inv02 = 1;
    51: op1_12_inv02 = 1;
    80: op1_12_inv02 = 1;
    62: op1_12_inv02 = 1;
    81: op1_12_inv02 = 1;
    52: op1_12_inv02 = 1;
    63: op1_12_inv02 = 1;
    83: op1_12_inv02 = 1;
    84: op1_12_inv02 = 1;
    66: op1_12_inv02 = 1;
    93: op1_12_inv02 = 1;
    94: op1_12_inv02 = 1;
    95: op1_12_inv02 = 1;
    96: op1_12_inv02 = 1;
    98: op1_12_inv02 = 1;
    100: op1_12_inv02 = 1;
    102: op1_12_inv02 = 1;
    37: op1_12_inv02 = 1;
    104: op1_12_inv02 = 1;
    106: op1_12_inv02 = 1;
    107: op1_12_inv02 = 1;
    110: op1_12_inv02 = 1;
    112: op1_12_inv02 = 1;
    113: op1_12_inv02 = 1;
    114: op1_12_inv02 = 1;
    116: op1_12_inv02 = 1;
    121: op1_12_inv02 = 1;
    123: op1_12_inv02 = 1;
    44: op1_12_inv02 = 1;
    127: op1_12_inv02 = 1;
    128: op1_12_inv02 = 1;
    129: op1_12_inv02 = 1;
    34: op1_12_inv02 = 1;
    default: op1_12_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in03 = imem05_in[7:4];
    53: op1_12_in03 = reg_0966;
    55: op1_12_in03 = reg_0876;
    73: op1_12_in03 = reg_0205;
    86: op1_12_in03 = reg_0255;
    74: op1_12_in03 = reg_0806;
    69: op1_12_in03 = reg_0976;
    49: op1_12_in03 = reg_0822;
    54: op1_12_in03 = reg_0412;
    75: op1_12_in03 = reg_0907;
    126: op1_12_in03 = reg_0907;
    56: op1_12_in03 = reg_0589;
    50: op1_12_in03 = reg_0571;
    100: op1_12_in03 = reg_0571;
    76: op1_12_in03 = reg_0204;
    63: op1_12_in03 = reg_0204;
    68: op1_12_in03 = reg_0957;
    71: op1_12_in03 = reg_1230;
    87: op1_12_in03 = reg_0382;
    57: op1_12_in03 = reg_0399;
    77: op1_12_in03 = reg_0133;
    58: op1_12_in03 = reg_0133;
    61: op1_12_in03 = reg_1028;
    78: op1_12_in03 = reg_0504;
    70: op1_12_in03 = reg_1003;
    59: op1_12_in03 = reg_0043;
    79: op1_12_in03 = reg_1334;
    51: op1_12_in03 = reg_0383;
    60: op1_12_in03 = reg_1079;
    88: op1_12_in03 = reg_0745;
    80: op1_12_in03 = reg_0804;
    83: op1_12_in03 = reg_0804;
    62: op1_12_in03 = reg_1169;
    81: op1_12_in03 = reg_0494;
    52: op1_12_in03 = reg_0931;
    82: op1_12_in03 = reg_0633;
    46: op1_12_in03 = reg_0728;
    64: op1_12_in03 = reg_1244;
    89: op1_12_in03 = reg_0673;
    84: op1_12_in03 = reg_0708;
    85: op1_12_in03 = reg_0233;
    65: op1_12_in03 = reg_0859;
    90: op1_12_in03 = reg_0597;
    48: op1_12_in03 = reg_0400;
    66: op1_12_in03 = reg_0860;
    91: op1_12_in03 = reg_0175;
    67: op1_12_in03 = reg_0667;
    92: op1_12_in03 = reg_1510;
    33: op1_12_in03 = reg_0051;
    93: op1_12_in03 = reg_0067;
    94: op1_12_in03 = reg_0338;
    28: op1_12_in03 = reg_0084;
    95: op1_12_in03 = reg_0759;
    96: op1_12_in03 = reg_0090;
    97: op1_12_in03 = reg_0782;
    98: op1_12_in03 = reg_0520;
    99: op1_12_in03 = reg_0895;
    101: op1_12_in03 = reg_0377;
    102: op1_12_in03 = reg_1096;
    37: op1_12_in03 = reg_0415;
    103: op1_12_in03 = reg_0824;
    104: op1_12_in03 = reg_0403;
    105: op1_12_in03 = reg_0306;
    106: op1_12_in03 = reg_1181;
    47: op1_12_in03 = reg_0598;
    107: op1_12_in03 = reg_0003;
    108: op1_12_in03 = reg_0829;
    109: op1_12_in03 = reg_1278;
    110: op1_12_in03 = reg_1065;
    111: op1_12_in03 = reg_0041;
    112: op1_12_in03 = reg_1200;
    113: op1_12_in03 = imem02_in[7:4];
    114: op1_12_in03 = reg_0219;
    115: op1_12_in03 = reg_0162;
    116: op1_12_in03 = reg_0825;
    117: op1_12_in03 = reg_0402;
    118: op1_12_in03 = reg_0198;
    119: op1_12_in03 = reg_0833;
    120: op1_12_in03 = reg_1298;
    121: op1_12_in03 = reg_0031;
    122: op1_12_in03 = reg_0039;
    123: op1_12_in03 = reg_0495;
    124: op1_12_in03 = reg_0580;
    125: op1_12_in03 = reg_1001;
    44: op1_12_in03 = reg_0340;
    127: op1_12_in03 = reg_0393;
    128: op1_12_in03 = reg_0206;
    129: op1_12_in03 = reg_1279;
    38: op1_12_in03 = reg_0739;
    130: op1_12_in03 = imem06_in[3:0];
    34: op1_12_in03 = reg_0102;
    default: op1_12_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv03 = 1;
    53: op1_12_inv03 = 1;
    86: op1_12_inv03 = 1;
    74: op1_12_inv03 = 1;
    69: op1_12_inv03 = 1;
    54: op1_12_inv03 = 1;
    50: op1_12_inv03 = 1;
    76: op1_12_inv03 = 1;
    68: op1_12_inv03 = 1;
    57: op1_12_inv03 = 1;
    77: op1_12_inv03 = 1;
    79: op1_12_inv03 = 1;
    51: op1_12_inv03 = 1;
    60: op1_12_inv03 = 1;
    80: op1_12_inv03 = 1;
    62: op1_12_inv03 = 1;
    81: op1_12_inv03 = 1;
    52: op1_12_inv03 = 1;
    83: op1_12_inv03 = 1;
    84: op1_12_inv03 = 1;
    65: op1_12_inv03 = 1;
    90: op1_12_inv03 = 1;
    48: op1_12_inv03 = 1;
    66: op1_12_inv03 = 1;
    91: op1_12_inv03 = 1;
    67: op1_12_inv03 = 1;
    92: op1_12_inv03 = 1;
    33: op1_12_inv03 = 1;
    93: op1_12_inv03 = 1;
    28: op1_12_inv03 = 1;
    99: op1_12_inv03 = 1;
    100: op1_12_inv03 = 1;
    102: op1_12_inv03 = 1;
    37: op1_12_inv03 = 1;
    103: op1_12_inv03 = 1;
    104: op1_12_inv03 = 1;
    106: op1_12_inv03 = 1;
    107: op1_12_inv03 = 1;
    110: op1_12_inv03 = 1;
    111: op1_12_inv03 = 1;
    112: op1_12_inv03 = 1;
    114: op1_12_inv03 = 1;
    115: op1_12_inv03 = 1;
    116: op1_12_inv03 = 1;
    118: op1_12_inv03 = 1;
    119: op1_12_inv03 = 1;
    121: op1_12_inv03 = 1;
    123: op1_12_inv03 = 1;
    125: op1_12_inv03 = 1;
    127: op1_12_inv03 = 1;
    128: op1_12_inv03 = 1;
    38: op1_12_inv03 = 1;
    130: op1_12_inv03 = 1;
    34: op1_12_inv03 = 1;
    default: op1_12_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in04 = reg_0037;
    53: op1_12_in04 = reg_0967;
    55: op1_12_in04 = reg_0008;
    113: op1_12_in04 = reg_0008;
    73: op1_12_in04 = reg_1430;
    76: op1_12_in04 = reg_1430;
    86: op1_12_in04 = reg_0168;
    74: op1_12_in04 = reg_1471;
    69: op1_12_in04 = reg_1018;
    49: op1_12_in04 = reg_0116;
    54: op1_12_in04 = reg_0407;
    75: op1_12_in04 = reg_0906;
    56: op1_12_in04 = reg_0561;
    50: op1_12_in04 = reg_0529;
    68: op1_12_in04 = reg_0190;
    71: op1_12_in04 = reg_0961;
    87: op1_12_in04 = reg_0473;
    57: op1_12_in04 = reg_0115;
    77: op1_12_in04 = reg_1508;
    61: op1_12_in04 = reg_0172;
    58: op1_12_in04 = reg_0606;
    78: op1_12_in04 = reg_0734;
    70: op1_12_in04 = reg_1231;
    59: op1_12_in04 = reg_0044;
    104: op1_12_in04 = reg_0044;
    79: op1_12_in04 = reg_0863;
    51: op1_12_in04 = reg_0365;
    60: op1_12_in04 = reg_1241;
    88: op1_12_in04 = reg_0897;
    80: op1_12_in04 = reg_1470;
    62: op1_12_in04 = reg_1163;
    81: op1_12_in04 = reg_0432;
    52: op1_12_in04 = reg_0979;
    63: op1_12_in04 = reg_0347;
    82: op1_12_in04 = reg_0020;
    46: op1_12_in04 = reg_0400;
    83: op1_12_in04 = reg_0805;
    124: op1_12_in04 = reg_0805;
    64: op1_12_in04 = reg_0804;
    89: op1_12_in04 = reg_1282;
    84: op1_12_in04 = reg_0748;
    129: op1_12_in04 = reg_0748;
    85: op1_12_in04 = reg_0235;
    65: op1_12_in04 = reg_0752;
    90: op1_12_in04 = reg_0558;
    48: op1_12_in04 = reg_0386;
    66: op1_12_in04 = reg_1323;
    91: op1_12_in04 = reg_0895;
    67: op1_12_in04 = reg_0674;
    92: op1_12_in04 = reg_1490;
    33: op1_12_in04 = reg_0085;
    93: op1_12_in04 = reg_0046;
    94: op1_12_in04 = reg_1189;
    28: op1_12_in04 = reg_0050;
    95: op1_12_in04 = reg_0573;
    96: op1_12_in04 = reg_1486;
    97: op1_12_in04 = reg_0271;
    98: op1_12_in04 = reg_1182;
    99: op1_12_in04 = reg_0530;
    100: op1_12_in04 = reg_0569;
    101: op1_12_in04 = reg_0889;
    102: op1_12_in04 = reg_0894;
    37: op1_12_in04 = reg_0618;
    103: op1_12_in04 = reg_1278;
    105: op1_12_in04 = reg_0711;
    108: op1_12_in04 = reg_0711;
    106: op1_12_in04 = reg_1403;
    47: op1_12_in04 = reg_0797;
    107: op1_12_in04 = reg_0001;
    109: op1_12_in04 = reg_1277;
    110: op1_12_in04 = reg_0342;
    111: op1_12_in04 = reg_0447;
    112: op1_12_in04 = reg_0414;
    114: op1_12_in04 = reg_0170;
    115: op1_12_in04 = reg_0402;
    116: op1_12_in04 = reg_0795;
    117: op1_12_in04 = reg_0403;
    118: op1_12_in04 = reg_1001;
    119: op1_12_in04 = reg_0367;
    120: op1_12_in04 = imem05_in[11:8];
    121: op1_12_in04 = reg_0029;
    122: op1_12_in04 = reg_0670;
    123: op1_12_in04 = reg_1451;
    125: op1_12_in04 = reg_0823;
    44: op1_12_in04 = reg_0262;
    126: op1_12_in04 = reg_0486;
    127: op1_12_in04 = reg_0317;
    128: op1_12_in04 = reg_0014;
    38: op1_12_in04 = reg_0002;
    130: op1_12_in04 = reg_0870;
    34: op1_12_in04 = reg_0103;
    default: op1_12_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_12_inv04 = 1;
    54: op1_12_inv04 = 1;
    50: op1_12_inv04 = 1;
    68: op1_12_inv04 = 1;
    58: op1_12_inv04 = 1;
    78: op1_12_inv04 = 1;
    60: op1_12_inv04 = 1;
    62: op1_12_inv04 = 1;
    52: op1_12_inv04 = 1;
    63: op1_12_inv04 = 1;
    64: op1_12_inv04 = 1;
    84: op1_12_inv04 = 1;
    85: op1_12_inv04 = 1;
    66: op1_12_inv04 = 1;
    67: op1_12_inv04 = 1;
    93: op1_12_inv04 = 1;
    28: op1_12_inv04 = 1;
    95: op1_12_inv04 = 1;
    97: op1_12_inv04 = 1;
    99: op1_12_inv04 = 1;
    100: op1_12_inv04 = 1;
    102: op1_12_inv04 = 1;
    37: op1_12_inv04 = 1;
    104: op1_12_inv04 = 1;
    105: op1_12_inv04 = 1;
    47: op1_12_inv04 = 1;
    108: op1_12_inv04 = 1;
    109: op1_12_inv04 = 1;
    111: op1_12_inv04 = 1;
    113: op1_12_inv04 = 1;
    115: op1_12_inv04 = 1;
    116: op1_12_inv04 = 1;
    117: op1_12_inv04 = 1;
    118: op1_12_inv04 = 1;
    120: op1_12_inv04 = 1;
    122: op1_12_inv04 = 1;
    123: op1_12_inv04 = 1;
    44: op1_12_inv04 = 1;
    126: op1_12_inv04 = 1;
    129: op1_12_inv04 = 1;
    default: op1_12_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in05 = reg_0754;
    53: op1_12_in05 = reg_0434;
    55: op1_12_in05 = reg_0830;
    73: op1_12_in05 = reg_1431;
    127: op1_12_in05 = reg_1431;
    86: op1_12_in05 = reg_0311;
    74: op1_12_in05 = reg_1470;
    83: op1_12_in05 = reg_1470;
    69: op1_12_in05 = reg_0587;
    49: op1_12_in05 = reg_0109;
    54: op1_12_in05 = reg_0471;
    75: op1_12_in05 = reg_0905;
    56: op1_12_in05 = reg_1140;
    50: op1_12_in05 = reg_0323;
    76: op1_12_in05 = reg_1269;
    68: op1_12_in05 = reg_1300;
    71: op1_12_in05 = reg_0460;
    87: op1_12_in05 = reg_0829;
    57: op1_12_in05 = reg_0714;
    77: op1_12_in05 = reg_0720;
    61: op1_12_in05 = reg_1230;
    58: op1_12_in05 = reg_0605;
    78: op1_12_in05 = reg_0849;
    70: op1_12_in05 = reg_0178;
    59: op1_12_in05 = reg_0486;
    79: op1_12_in05 = reg_0669;
    116: op1_12_in05 = reg_0669;
    51: op1_12_in05 = reg_0047;
    60: op1_12_in05 = reg_0803;
    64: op1_12_in05 = reg_0803;
    88: op1_12_in05 = reg_0848;
    80: op1_12_in05 = reg_0218;
    62: op1_12_in05 = reg_0650;
    81: op1_12_in05 = reg_0970;
    52: op1_12_in05 = reg_0784;
    63: op1_12_in05 = reg_1169;
    82: op1_12_in05 = reg_0470;
    46: op1_12_in05 = reg_0385;
    89: op1_12_in05 = reg_1384;
    84: op1_12_in05 = reg_0579;
    85: op1_12_in05 = reg_0444;
    65: op1_12_in05 = reg_0751;
    90: op1_12_in05 = reg_0884;
    48: op1_12_in05 = reg_0365;
    66: op1_12_in05 = reg_0752;
    91: op1_12_in05 = reg_1071;
    67: op1_12_in05 = reg_0187;
    92: op1_12_in05 = reg_1491;
    93: op1_12_in05 = reg_1170;
    94: op1_12_in05 = reg_0016;
    28: op1_12_in05 = reg_0052;
    95: op1_12_in05 = reg_0330;
    96: op1_12_in05 = reg_1484;
    97: op1_12_in05 = reg_1501;
    99: op1_12_in05 = reg_0399;
    100: op1_12_in05 = reg_0345;
    101: op1_12_in05 = reg_0328;
    102: op1_12_in05 = reg_0135;
    37: op1_12_in05 = reg_0591;
    103: op1_12_in05 = reg_0804;
    104: op1_12_in05 = reg_0012;
    105: op1_12_in05 = reg_0235;
    106: op1_12_in05 = reg_1402;
    47: op1_12_in05 = reg_0932;
    107: op1_12_in05 = reg_0053;
    108: op1_12_in05 = reg_1091;
    109: op1_12_in05 = reg_0748;
    110: op1_12_in05 = reg_0097;
    111: op1_12_in05 = reg_0662;
    112: op1_12_in05 = reg_1040;
    113: op1_12_in05 = reg_0879;
    114: op1_12_in05 = reg_0741;
    115: op1_12_in05 = reg_0011;
    117: op1_12_in05 = reg_0634;
    118: op1_12_in05 = reg_0600;
    119: op1_12_in05 = reg_0136;
    120: op1_12_in05 = reg_1059;
    121: op1_12_in05 = reg_0284;
    122: op1_12_in05 = reg_0925;
    123: op1_12_in05 = reg_0105;
    124: op1_12_in05 = reg_1052;
    125: op1_12_in05 = reg_0312;
    44: op1_12_in05 = reg_0487;
    126: op1_12_in05 = reg_1053;
    128: op1_12_in05 = reg_0039;
    129: op1_12_in05 = reg_0806;
    38: op1_12_in05 = reg_0518;
    130: op1_12_in05 = reg_0782;
    34: op1_12_in05 = reg_0114;
    default: op1_12_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv05 = 1;
    53: op1_12_inv05 = 1;
    55: op1_12_inv05 = 1;
    73: op1_12_inv05 = 1;
    86: op1_12_inv05 = 1;
    69: op1_12_inv05 = 1;
    49: op1_12_inv05 = 1;
    54: op1_12_inv05 = 1;
    56: op1_12_inv05 = 1;
    68: op1_12_inv05 = 1;
    57: op1_12_inv05 = 1;
    77: op1_12_inv05 = 1;
    70: op1_12_inv05 = 1;
    59: op1_12_inv05 = 1;
    79: op1_12_inv05 = 1;
    51: op1_12_inv05 = 1;
    88: op1_12_inv05 = 1;
    81: op1_12_inv05 = 1;
    52: op1_12_inv05 = 1;
    63: op1_12_inv05 = 1;
    46: op1_12_inv05 = 1;
    85: op1_12_inv05 = 1;
    48: op1_12_inv05 = 1;
    66: op1_12_inv05 = 1;
    91: op1_12_inv05 = 1;
    67: op1_12_inv05 = 1;
    92: op1_12_inv05 = 1;
    93: op1_12_inv05 = 1;
    94: op1_12_inv05 = 1;
    96: op1_12_inv05 = 1;
    100: op1_12_inv05 = 1;
    101: op1_12_inv05 = 1;
    37: op1_12_inv05 = 1;
    104: op1_12_inv05 = 1;
    47: op1_12_inv05 = 1;
    111: op1_12_inv05 = 1;
    112: op1_12_inv05 = 1;
    115: op1_12_inv05 = 1;
    117: op1_12_inv05 = 1;
    119: op1_12_inv05 = 1;
    124: op1_12_inv05 = 1;
    125: op1_12_inv05 = 1;
    129: op1_12_inv05 = 1;
    38: op1_12_inv05 = 1;
    130: op1_12_inv05 = 1;
    34: op1_12_inv05 = 1;
    default: op1_12_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in06 = reg_0730;
    53: op1_12_in06 = reg_0384;
    55: op1_12_in06 = reg_0829;
    73: op1_12_in06 = reg_0395;
    76: op1_12_in06 = reg_0395;
    86: op1_12_in06 = reg_0312;
    118: op1_12_in06 = reg_0312;
    74: op1_12_in06 = reg_1454;
    69: op1_12_in06 = reg_0563;
    49: op1_12_in06 = reg_0670;
    54: op1_12_in06 = reg_0796;
    75: op1_12_in06 = reg_1420;
    56: op1_12_in06 = imem02_in[15:12];
    50: op1_12_in06 = reg_0244;
    68: op1_12_in06 = reg_1301;
    71: op1_12_in06 = reg_0459;
    87: op1_12_in06 = reg_0801;
    57: op1_12_in06 = reg_0634;
    77: op1_12_in06 = reg_1505;
    61: op1_12_in06 = reg_1206;
    58: op1_12_in06 = reg_0607;
    78: op1_12_in06 = reg_0790;
    70: op1_12_in06 = reg_0113;
    59: op1_12_in06 = reg_1029;
    79: op1_12_in06 = reg_0109;
    51: op1_12_in06 = reg_0901;
    60: op1_12_in06 = reg_0476;
    88: op1_12_in06 = reg_0069;
    80: op1_12_in06 = reg_1028;
    62: op1_12_in06 = reg_0300;
    81: op1_12_in06 = reg_0126;
    52: op1_12_in06 = reg_1058;
    63: op1_12_in06 = reg_0176;
    82: op1_12_in06 = reg_0370;
    46: op1_12_in06 = reg_0362;
    83: op1_12_in06 = reg_1053;
    64: op1_12_in06 = reg_1052;
    89: op1_12_in06 = reg_0535;
    84: op1_12_in06 = reg_0702;
    85: op1_12_in06 = reg_1448;
    65: op1_12_in06 = reg_0141;
    90: op1_12_in06 = imem03_in[15:12];
    48: op1_12_in06 = reg_0091;
    66: op1_12_in06 = reg_0827;
    91: op1_12_in06 = reg_0590;
    67: op1_12_in06 = reg_0703;
    92: op1_12_in06 = reg_0615;
    103: op1_12_in06 = reg_0615;
    93: op1_12_in06 = reg_0478;
    94: op1_12_in06 = reg_0315;
    28: op1_12_in06 = imem07_in[15:12];
    95: op1_12_in06 = reg_0216;
    96: op1_12_in06 = reg_0492;
    97: op1_12_in06 = reg_0115;
    99: op1_12_in06 = reg_0846;
    100: op1_12_in06 = reg_1228;
    101: op1_12_in06 = reg_0185;
    102: op1_12_in06 = reg_1440;
    37: op1_12_in06 = reg_0103;
    104: op1_12_in06 = reg_0447;
    105: op1_12_in06 = reg_0479;
    106: op1_12_in06 = reg_0940;
    47: op1_12_in06 = reg_0452;
    107: op1_12_in06 = reg_0123;
    108: op1_12_in06 = reg_0024;
    109: op1_12_in06 = reg_0501;
    110: op1_12_in06 = reg_0368;
    111: op1_12_in06 = imem02_in[11:8];
    112: op1_12_in06 = reg_0342;
    113: op1_12_in06 = reg_0276;
    114: op1_12_in06 = reg_0740;
    115: op1_12_in06 = reg_0166;
    116: op1_12_in06 = reg_0696;
    117: op1_12_in06 = reg_0043;
    119: op1_12_in06 = imem05_in[11:8];
    120: op1_12_in06 = reg_0735;
    121: op1_12_in06 = reg_0741;
    122: op1_12_in06 = reg_0870;
    123: op1_12_in06 = reg_0631;
    124: op1_12_in06 = reg_0293;
    125: op1_12_in06 = reg_0143;
    44: op1_12_in06 = reg_0835;
    126: op1_12_in06 = reg_0250;
    127: op1_12_in06 = imem06_in[3:0];
    128: op1_12_in06 = imem06_in[7:4];
    129: op1_12_in06 = reg_0803;
    130: op1_12_in06 = reg_1323;
    34: op1_12_in06 = reg_0050;
    default: op1_12_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_12_inv06 = 1;
    69: op1_12_inv06 = 1;
    56: op1_12_inv06 = 1;
    50: op1_12_inv06 = 1;
    87: op1_12_inv06 = 1;
    57: op1_12_inv06 = 1;
    77: op1_12_inv06 = 1;
    61: op1_12_inv06 = 1;
    58: op1_12_inv06 = 1;
    70: op1_12_inv06 = 1;
    59: op1_12_inv06 = 1;
    79: op1_12_inv06 = 1;
    60: op1_12_inv06 = 1;
    80: op1_12_inv06 = 1;
    62: op1_12_inv06 = 1;
    63: op1_12_inv06 = 1;
    46: op1_12_inv06 = 1;
    48: op1_12_inv06 = 1;
    94: op1_12_inv06 = 1;
    100: op1_12_inv06 = 1;
    101: op1_12_inv06 = 1;
    102: op1_12_inv06 = 1;
    103: op1_12_inv06 = 1;
    105: op1_12_inv06 = 1;
    108: op1_12_inv06 = 1;
    111: op1_12_inv06 = 1;
    114: op1_12_inv06 = 1;
    115: op1_12_inv06 = 1;
    116: op1_12_inv06 = 1;
    117: op1_12_inv06 = 1;
    118: op1_12_inv06 = 1;
    119: op1_12_inv06 = 1;
    122: op1_12_inv06 = 1;
    123: op1_12_inv06 = 1;
    124: op1_12_inv06 = 1;
    44: op1_12_inv06 = 1;
    128: op1_12_inv06 = 1;
    129: op1_12_inv06 = 1;
    130: op1_12_inv06 = 1;
    34: op1_12_inv06 = 1;
    default: op1_12_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in07 = reg_0316;
    66: op1_12_in07 = reg_0316;
    53: op1_12_in07 = reg_0385;
    55: op1_12_in07 = reg_0279;
    73: op1_12_in07 = reg_0996;
    86: op1_12_in07 = reg_0840;
    74: op1_12_in07 = reg_1230;
    69: op1_12_in07 = reg_0561;
    113: op1_12_in07 = reg_0561;
    49: op1_12_in07 = reg_0637;
    54: op1_12_in07 = reg_0797;
    75: op1_12_in07 = imem06_in[3:0];
    56: op1_12_in07 = reg_0776;
    50: op1_12_in07 = reg_0271;
    76: op1_12_in07 = reg_1259;
    68: op1_12_in07 = reg_0558;
    71: op1_12_in07 = reg_0388;
    87: op1_12_in07 = reg_0327;
    57: op1_12_in07 = reg_0619;
    77: op1_12_in07 = reg_1501;
    61: op1_12_in07 = reg_0202;
    60: op1_12_in07 = reg_0202;
    58: op1_12_in07 = reg_0531;
    78: op1_12_in07 = reg_0411;
    70: op1_12_in07 = reg_0481;
    59: op1_12_in07 = reg_0976;
    79: op1_12_in07 = reg_0586;
    51: op1_12_in07 = reg_0079;
    88: op1_12_in07 = reg_0168;
    80: op1_12_in07 = reg_1206;
    62: op1_12_in07 = reg_0197;
    81: op1_12_in07 = reg_1433;
    52: op1_12_in07 = reg_0908;
    63: op1_12_in07 = reg_0649;
    82: op1_12_in07 = reg_0347;
    84: op1_12_in07 = reg_0347;
    46: op1_12_in07 = reg_0047;
    83: op1_12_in07 = reg_1052;
    64: op1_12_in07 = reg_0476;
    89: op1_12_in07 = reg_1198;
    85: op1_12_in07 = reg_1063;
    65: op1_12_in07 = reg_0585;
    90: op1_12_in07 = reg_0313;
    48: op1_12_in07 = reg_0724;
    91: op1_12_in07 = reg_0138;
    67: op1_12_in07 = reg_0225;
    92: op1_12_in07 = reg_1053;
    93: op1_12_in07 = imem07_in[15:12];
    94: op1_12_in07 = reg_0204;
    95: op1_12_in07 = reg_1033;
    96: op1_12_in07 = reg_0275;
    97: op1_12_in07 = reg_0979;
    99: op1_12_in07 = reg_0455;
    100: op1_12_in07 = reg_0132;
    101: op1_12_in07 = reg_0216;
    102: op1_12_in07 = reg_0703;
    37: op1_12_in07 = reg_0228;
    103: op1_12_in07 = reg_0293;
    126: op1_12_in07 = reg_0293;
    104: op1_12_in07 = reg_1071;
    105: op1_12_in07 = reg_0732;
    106: op1_12_in07 = reg_0937;
    47: op1_12_in07 = reg_0721;
    107: op1_12_in07 = reg_1182;
    108: op1_12_in07 = reg_0068;
    109: op1_12_in07 = reg_1490;
    110: op1_12_in07 = reg_1312;
    111: op1_12_in07 = reg_1235;
    112: op1_12_in07 = reg_0698;
    114: op1_12_in07 = reg_0738;
    115: op1_12_in07 = reg_0662;
    117: op1_12_in07 = reg_0662;
    116: op1_12_in07 = reg_0827;
    118: op1_12_in07 = reg_0191;
    119: op1_12_in07 = reg_0272;
    120: op1_12_in07 = reg_0466;
    121: op1_12_in07 = reg_0404;
    122: op1_12_in07 = reg_0696;
    123: op1_12_in07 = reg_0379;
    124: op1_12_in07 = reg_0221;
    125: op1_12_in07 = reg_1494;
    44: op1_12_in07 = reg_0237;
    127: op1_12_in07 = reg_0729;
    128: op1_12_in07 = reg_0270;
    129: op1_12_in07 = reg_0248;
    130: op1_12_in07 = reg_1505;
    34: op1_12_in07 = reg_0051;
    default: op1_12_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv07 = 1;
    75: op1_12_inv07 = 1;
    76: op1_12_inv07 = 1;
    68: op1_12_inv07 = 1;
    71: op1_12_inv07 = 1;
    77: op1_12_inv07 = 1;
    58: op1_12_inv07 = 1;
    70: op1_12_inv07 = 1;
    59: op1_12_inv07 = 1;
    79: op1_12_inv07 = 1;
    51: op1_12_inv07 = 1;
    88: op1_12_inv07 = 1;
    81: op1_12_inv07 = 1;
    82: op1_12_inv07 = 1;
    46: op1_12_inv07 = 1;
    64: op1_12_inv07 = 1;
    84: op1_12_inv07 = 1;
    65: op1_12_inv07 = 1;
    66: op1_12_inv07 = 1;
    91: op1_12_inv07 = 1;
    67: op1_12_inv07 = 1;
    94: op1_12_inv07 = 1;
    97: op1_12_inv07 = 1;
    100: op1_12_inv07 = 1;
    37: op1_12_inv07 = 1;
    105: op1_12_inv07 = 1;
    108: op1_12_inv07 = 1;
    110: op1_12_inv07 = 1;
    111: op1_12_inv07 = 1;
    116: op1_12_inv07 = 1;
    117: op1_12_inv07 = 1;
    119: op1_12_inv07 = 1;
    120: op1_12_inv07 = 1;
    123: op1_12_inv07 = 1;
    124: op1_12_inv07 = 1;
    125: op1_12_inv07 = 1;
    44: op1_12_inv07 = 1;
    128: op1_12_inv07 = 1;
    129: op1_12_inv07 = 1;
    130: op1_12_inv07 = 1;
    default: op1_12_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in08 = reg_0172;
    77: op1_12_in08 = reg_0172;
    53: op1_12_in08 = reg_0077;
    55: op1_12_in08 = reg_0756;
    73: op1_12_in08 = reg_0992;
    86: op1_12_in08 = reg_0699;
    74: op1_12_in08 = reg_0460;
    61: op1_12_in08 = reg_0460;
    69: op1_12_in08 = reg_1260;
    49: op1_12_in08 = reg_0264;
    66: op1_12_in08 = reg_0264;
    54: op1_12_in08 = reg_0370;
    75: op1_12_in08 = reg_1334;
    56: op1_12_in08 = reg_0307;
    50: op1_12_in08 = reg_0215;
    76: op1_12_in08 = reg_1164;
    68: op1_12_in08 = reg_0880;
    71: op1_12_in08 = reg_0203;
    87: op1_12_in08 = reg_0227;
    57: op1_12_in08 = reg_0568;
    58: op1_12_in08 = imem02_in[11:8];
    104: op1_12_in08 = imem02_in[11:8];
    78: op1_12_in08 = reg_0898;
    70: op1_12_in08 = reg_0525;
    59: op1_12_in08 = reg_0455;
    79: op1_12_in08 = reg_0979;
    51: op1_12_in08 = reg_0043;
    60: op1_12_in08 = reg_0961;
    80: op1_12_in08 = reg_0961;
    92: op1_12_in08 = reg_0961;
    88: op1_12_in08 = reg_0559;
    62: op1_12_in08 = reg_0240;
    81: op1_12_in08 = reg_0711;
    52: op1_12_in08 = reg_0869;
    63: op1_12_in08 = reg_0567;
    82: op1_12_in08 = reg_1169;
    46: op1_12_in08 = reg_0899;
    83: op1_12_in08 = reg_1028;
    126: op1_12_in08 = reg_1028;
    64: op1_12_in08 = reg_1227;
    89: op1_12_in08 = reg_0488;
    84: op1_12_in08 = reg_1168;
    85: op1_12_in08 = reg_0783;
    65: op1_12_in08 = reg_0622;
    90: op1_12_in08 = reg_0673;
    48: op1_12_in08 = reg_0868;
    91: op1_12_in08 = reg_1344;
    67: op1_12_in08 = reg_0297;
    93: op1_12_in08 = reg_0461;
    94: op1_12_in08 = reg_0136;
    95: op1_12_in08 = reg_0145;
    96: op1_12_in08 = reg_1373;
    97: op1_12_in08 = reg_1225;
    99: op1_12_in08 = reg_1018;
    100: op1_12_in08 = reg_0396;
    101: op1_12_in08 = reg_0198;
    102: op1_12_in08 = reg_0299;
    37: op1_12_in08 = reg_0050;
    103: op1_12_in08 = reg_1459;
    105: op1_12_in08 = reg_0444;
    106: op1_12_in08 = reg_0197;
    47: op1_12_in08 = reg_0470;
    108: op1_12_in08 = reg_0962;
    109: op1_12_in08 = reg_0580;
    110: op1_12_in08 = reg_0536;
    111: op1_12_in08 = reg_0423;
    112: op1_12_in08 = reg_0582;
    113: op1_12_in08 = reg_0495;
    114: op1_12_in08 = reg_0103;
    115: op1_12_in08 = imem02_in[3:0];
    116: op1_12_in08 = reg_1501;
    117: op1_12_in08 = reg_0475;
    118: op1_12_in08 = reg_0234;
    119: op1_12_in08 = reg_1268;
    120: op1_12_in08 = reg_1268;
    121: op1_12_in08 = reg_0593;
    122: op1_12_in08 = reg_1467;
    123: op1_12_in08 = reg_1078;
    124: op1_12_in08 = reg_0485;
    125: op1_12_in08 = reg_0070;
    44: op1_12_in08 = reg_0117;
    127: op1_12_in08 = reg_0397;
    128: op1_12_in08 = reg_0859;
    129: op1_12_in08 = reg_0250;
    130: op1_12_in08 = reg_1179;
    34: op1_12_in08 = reg_0003;
    default: op1_12_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv08 = 1;
    55: op1_12_inv08 = 1;
    73: op1_12_inv08 = 1;
    74: op1_12_inv08 = 1;
    69: op1_12_inv08 = 1;
    49: op1_12_inv08 = 1;
    54: op1_12_inv08 = 1;
    87: op1_12_inv08 = 1;
    61: op1_12_inv08 = 1;
    79: op1_12_inv08 = 1;
    51: op1_12_inv08 = 1;
    80: op1_12_inv08 = 1;
    81: op1_12_inv08 = 1;
    52: op1_12_inv08 = 1;
    63: op1_12_inv08 = 1;
    82: op1_12_inv08 = 1;
    83: op1_12_inv08 = 1;
    89: op1_12_inv08 = 1;
    84: op1_12_inv08 = 1;
    85: op1_12_inv08 = 1;
    65: op1_12_inv08 = 1;
    66: op1_12_inv08 = 1;
    67: op1_12_inv08 = 1;
    93: op1_12_inv08 = 1;
    94: op1_12_inv08 = 1;
    97: op1_12_inv08 = 1;
    99: op1_12_inv08 = 1;
    100: op1_12_inv08 = 1;
    37: op1_12_inv08 = 1;
    104: op1_12_inv08 = 1;
    47: op1_12_inv08 = 1;
    108: op1_12_inv08 = 1;
    113: op1_12_inv08 = 1;
    116: op1_12_inv08 = 1;
    118: op1_12_inv08 = 1;
    120: op1_12_inv08 = 1;
    121: op1_12_inv08 = 1;
    125: op1_12_inv08 = 1;
    126: op1_12_inv08 = 1;
    default: op1_12_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in09 = reg_0714;
    53: op1_12_in09 = reg_0291;
    55: op1_12_in09 = reg_0677;
    73: op1_12_in09 = reg_0346;
    86: op1_12_in09 = reg_0573;
    105: op1_12_in09 = reg_0573;
    74: op1_12_in09 = reg_0476;
    69: op1_12_in09 = reg_0935;
    49: op1_12_in09 = reg_0247;
    54: op1_12_in09 = reg_0452;
    75: op1_12_in09 = reg_0869;
    56: op1_12_in09 = reg_0878;
    50: op1_12_in09 = reg_0391;
    76: op1_12_in09 = reg_0131;
    68: op1_12_in09 = reg_0479;
    71: op1_12_in09 = reg_0060;
    87: op1_12_in09 = reg_0168;
    57: op1_12_in09 = reg_0570;
    77: op1_12_in09 = reg_1065;
    61: op1_12_in09 = reg_0492;
    58: op1_12_in09 = reg_0669;
    78: op1_12_in09 = reg_0208;
    70: op1_12_in09 = reg_0411;
    59: op1_12_in09 = reg_0560;
    79: op1_12_in09 = reg_0244;
    51: op1_12_in09 = reg_0011;
    60: op1_12_in09 = reg_0725;
    88: op1_12_in09 = reg_0706;
    80: op1_12_in09 = reg_0459;
    62: op1_12_in09 = reg_0449;
    81: op1_12_in09 = reg_0009;
    52: op1_12_in09 = reg_0373;
    63: op1_12_in09 = reg_0566;
    82: op1_12_in09 = reg_0992;
    46: op1_12_in09 = reg_0277;
    83: op1_12_in09 = reg_1432;
    64: op1_12_in09 = reg_0987;
    89: op1_12_in09 = reg_0681;
    84: op1_12_in09 = imem05_in[7:4];
    85: op1_12_in09 = reg_0891;
    65: op1_12_in09 = reg_0571;
    90: op1_12_in09 = reg_0443;
    48: op1_12_in09 = reg_0078;
    66: op1_12_in09 = reg_0718;
    91: op1_12_in09 = reg_0776;
    67: op1_12_in09 = reg_1345;
    92: op1_12_in09 = reg_0722;
    93: op1_12_in09 = reg_1415;
    94: op1_12_in09 = reg_0466;
    95: op1_12_in09 = reg_0144;
    96: op1_12_in09 = reg_0196;
    97: op1_12_in09 = reg_0165;
    99: op1_12_in09 = reg_0608;
    100: op1_12_in09 = reg_0067;
    101: op1_12_in09 = reg_0312;
    102: op1_12_in09 = reg_0140;
    37: op1_12_in09 = reg_0051;
    114: op1_12_in09 = reg_0051;
    103: op1_12_in09 = reg_0249;
    104: op1_12_in09 = reg_0889;
    106: op1_12_in09 = reg_0601;
    47: op1_12_in09 = reg_0340;
    108: op1_12_in09 = reg_1003;
    109: op1_12_in09 = reg_0486;
    110: op1_12_in09 = reg_0016;
    111: op1_12_in09 = reg_0975;
    112: op1_12_in09 = reg_1143;
    113: op1_12_in09 = reg_1207;
    115: op1_12_in09 = reg_1002;
    116: op1_12_in09 = reg_0780;
    117: op1_12_in09 = reg_0322;
    118: op1_12_in09 = reg_0000;
    119: op1_12_in09 = reg_0176;
    120: op1_12_in09 = reg_0066;
    121: op1_12_in09 = reg_0086;
    122: op1_12_in09 = reg_0860;
    127: op1_12_in09 = reg_0860;
    123: op1_12_in09 = reg_1091;
    124: op1_12_in09 = reg_0460;
    125: op1_12_in09 = reg_1516;
    44: op1_12_in09 = reg_0211;
    126: op1_12_in09 = reg_1229;
    128: op1_12_in09 = reg_1467;
    129: op1_12_in09 = reg_1459;
    130: op1_12_in09 = reg_0265;
    34: op1_12_in09 = reg_0001;
    default: op1_12_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv09 = 1;
    73: op1_12_inv09 = 1;
    86: op1_12_inv09 = 1;
    54: op1_12_inv09 = 1;
    75: op1_12_inv09 = 1;
    56: op1_12_inv09 = 1;
    50: op1_12_inv09 = 1;
    76: op1_12_inv09 = 1;
    68: op1_12_inv09 = 1;
    71: op1_12_inv09 = 1;
    87: op1_12_inv09 = 1;
    57: op1_12_inv09 = 1;
    70: op1_12_inv09 = 1;
    59: op1_12_inv09 = 1;
    80: op1_12_inv09 = 1;
    63: op1_12_inv09 = 1;
    82: op1_12_inv09 = 1;
    46: op1_12_inv09 = 1;
    83: op1_12_inv09 = 1;
    89: op1_12_inv09 = 1;
    90: op1_12_inv09 = 1;
    67: op1_12_inv09 = 1;
    92: op1_12_inv09 = 1;
    94: op1_12_inv09 = 1;
    95: op1_12_inv09 = 1;
    96: op1_12_inv09 = 1;
    97: op1_12_inv09 = 1;
    100: op1_12_inv09 = 1;
    104: op1_12_inv09 = 1;
    106: op1_12_inv09 = 1;
    47: op1_12_inv09 = 1;
    108: op1_12_inv09 = 1;
    110: op1_12_inv09 = 1;
    111: op1_12_inv09 = 1;
    112: op1_12_inv09 = 1;
    113: op1_12_inv09 = 1;
    115: op1_12_inv09 = 1;
    120: op1_12_inv09 = 1;
    121: op1_12_inv09 = 1;
    125: op1_12_inv09 = 1;
    127: op1_12_inv09 = 1;
    default: op1_12_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in10 = reg_1302;
    53: op1_12_in10 = reg_0278;
    55: op1_12_in10 = reg_0675;
    73: op1_12_in10 = reg_0648;
    119: op1_12_in10 = reg_0648;
    86: op1_12_in10 = reg_0198;
    74: op1_12_in10 = reg_0351;
    69: op1_12_in10 = reg_0128;
    49: op1_12_in10 = reg_0528;
    54: op1_12_in10 = reg_0181;
    75: op1_12_in10 = reg_1323;
    56: op1_12_in10 = reg_0846;
    50: op1_12_in10 = reg_0230;
    76: op1_12_in10 = reg_0182;
    68: op1_12_in10 = imem03_in[3:0];
    71: op1_12_in10 = reg_0057;
    87: op1_12_in10 = reg_0006;
    57: op1_12_in10 = reg_0119;
    77: op1_12_in10 = reg_0115;
    61: op1_12_in10 = reg_0959;
    58: op1_12_in10 = reg_0475;
    78: op1_12_in10 = reg_1340;
    70: op1_12_in10 = reg_0898;
    59: op1_12_in10 = imem02_in[15:12];
    79: op1_12_in10 = reg_1204;
    51: op1_12_in10 = reg_0222;
    46: op1_12_in10 = reg_0222;
    60: op1_12_in10 = reg_0189;
    88: op1_12_in10 = reg_1447;
    80: op1_12_in10 = reg_0887;
    62: op1_12_in10 = imem05_in[15:12];
    81: op1_12_in10 = reg_0294;
    52: op1_12_in10 = reg_0826;
    63: op1_12_in10 = reg_0745;
    82: op1_12_in10 = reg_0650;
    83: op1_12_in10 = reg_0459;
    64: op1_12_in10 = reg_0459;
    89: op1_12_in10 = reg_0471;
    84: op1_12_in10 = reg_0391;
    120: op1_12_in10 = reg_0391;
    85: op1_12_in10 = reg_0989;
    65: op1_12_in10 = reg_0569;
    90: op1_12_in10 = reg_0034;
    48: op1_12_in10 = reg_0088;
    66: op1_12_in10 = reg_0717;
    91: op1_12_in10 = reg_0970;
    67: op1_12_in10 = reg_0921;
    92: op1_12_in10 = reg_0389;
    93: op1_12_in10 = reg_1056;
    94: op1_12_in10 = reg_0346;
    95: op1_12_in10 = reg_0965;
    96: op1_12_in10 = reg_0393;
    97: op1_12_in10 = reg_1202;
    99: op1_12_in10 = reg_0588;
    100: op1_12_in10 = reg_0212;
    101: op1_12_in10 = reg_0180;
    102: op1_12_in10 = reg_0159;
    37: op1_12_in10 = reg_0519;
    103: op1_12_in10 = reg_1432;
    104: op1_12_in10 = reg_0455;
    111: op1_12_in10 = reg_0455;
    105: op1_12_in10 = reg_0709;
    106: op1_12_in10 = reg_0118;
    47: op1_12_in10 = reg_0305;
    108: op1_12_in10 = reg_1033;
    109: op1_12_in10 = reg_0640;
    110: op1_12_in10 = reg_0021;
    112: op1_12_in10 = reg_0487;
    113: op1_12_in10 = reg_0494;
    114: op1_12_in10 = reg_0053;
    115: op1_12_in10 = reg_0169;
    116: op1_12_in10 = reg_1508;
    117: op1_12_in10 = imem02_in[7:4];
    118: op1_12_in10 = reg_0375;
    122: op1_12_in10 = reg_0859;
    123: op1_12_in10 = reg_0217;
    124: op1_12_in10 = reg_0060;
    125: op1_12_in10 = reg_1314;
    44: op1_12_in10 = reg_0063;
    126: op1_12_in10 = reg_0961;
    129: op1_12_in10 = reg_0961;
    127: op1_12_in10 = reg_0619;
    128: op1_12_in10 = reg_1505;
    130: op1_12_in10 = reg_0716;
    34: op1_12_in10 = reg_0002;
    default: op1_12_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv10 = 1;
    53: op1_12_inv10 = 1;
    74: op1_12_inv10 = 1;
    69: op1_12_inv10 = 1;
    49: op1_12_inv10 = 1;
    54: op1_12_inv10 = 1;
    56: op1_12_inv10 = 1;
    76: op1_12_inv10 = 1;
    68: op1_12_inv10 = 1;
    71: op1_12_inv10 = 1;
    57: op1_12_inv10 = 1;
    77: op1_12_inv10 = 1;
    58: op1_12_inv10 = 1;
    70: op1_12_inv10 = 1;
    59: op1_12_inv10 = 1;
    79: op1_12_inv10 = 1;
    51: op1_12_inv10 = 1;
    60: op1_12_inv10 = 1;
    80: op1_12_inv10 = 1;
    62: op1_12_inv10 = 1;
    82: op1_12_inv10 = 1;
    83: op1_12_inv10 = 1;
    84: op1_12_inv10 = 1;
    90: op1_12_inv10 = 1;
    48: op1_12_inv10 = 1;
    66: op1_12_inv10 = 1;
    91: op1_12_inv10 = 1;
    67: op1_12_inv10 = 1;
    92: op1_12_inv10 = 1;
    93: op1_12_inv10 = 1;
    96: op1_12_inv10 = 1;
    97: op1_12_inv10 = 1;
    101: op1_12_inv10 = 1;
    102: op1_12_inv10 = 1;
    106: op1_12_inv10 = 1;
    47: op1_12_inv10 = 1;
    112: op1_12_inv10 = 1;
    114: op1_12_inv10 = 1;
    115: op1_12_inv10 = 1;
    116: op1_12_inv10 = 1;
    119: op1_12_inv10 = 1;
    122: op1_12_inv10 = 1;
    124: op1_12_inv10 = 1;
    125: op1_12_inv10 = 1;
    126: op1_12_inv10 = 1;
    129: op1_12_inv10 = 1;
    130: op1_12_inv10 = 1;
    default: op1_12_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in11 = reg_0619;
    53: op1_12_in11 = reg_0283;
    55: op1_12_in11 = reg_0556;
    118: op1_12_in11 = reg_0556;
    73: op1_12_in11 = reg_0333;
    86: op1_12_in11 = reg_1001;
    74: op1_12_in11 = reg_0431;
    69: op1_12_in11 = reg_0106;
    49: op1_12_in11 = reg_0018;
    54: op1_12_in11 = reg_0065;
    75: op1_12_in11 = reg_0984;
    56: op1_12_in11 = reg_0311;
    50: op1_12_in11 = reg_0252;
    76: op1_12_in11 = reg_0334;
    68: op1_12_in11 = reg_0032;
    71: op1_12_in11 = reg_1290;
    87: op1_12_in11 = reg_0233;
    57: op1_12_in11 = reg_0165;
    77: op1_12_in11 = reg_0585;
    61: op1_12_in11 = reg_0725;
    58: op1_12_in11 = reg_0054;
    78: op1_12_in11 = reg_1216;
    70: op1_12_in11 = reg_1312;
    112: op1_12_in11 = reg_1312;
    59: op1_12_in11 = reg_0497;
    79: op1_12_in11 = reg_0067;
    51: op1_12_in11 = reg_0667;
    60: op1_12_in11 = reg_0057;
    88: op1_12_in11 = reg_0049;
    80: op1_12_in11 = reg_0073;
    62: op1_12_in11 = reg_0037;
    81: op1_12_in11 = reg_0280;
    52: op1_12_in11 = reg_0115;
    63: op1_12_in11 = reg_0272;
    82: op1_12_in11 = imem05_in[11:8];
    46: op1_12_in11 = reg_0486;
    83: op1_12_in11 = reg_0887;
    64: op1_12_in11 = reg_0928;
    129: op1_12_in11 = reg_0928;
    89: op1_12_in11 = reg_1077;
    84: op1_12_in11 = reg_0564;
    85: op1_12_in11 = reg_1516;
    65: op1_12_in11 = reg_0570;
    90: op1_12_in11 = reg_1339;
    48: op1_12_in11 = reg_0282;
    66: op1_12_in11 = reg_0194;
    91: op1_12_in11 = reg_0127;
    67: op1_12_in11 = reg_1094;
    92: op1_12_in11 = reg_0071;
    93: op1_12_in11 = reg_0225;
    94: op1_12_in11 = reg_0992;
    95: op1_12_in11 = reg_1231;
    96: op1_12_in11 = reg_0243;
    97: op1_12_in11 = reg_0269;
    99: op1_12_in11 = reg_0472;
    100: op1_12_in11 = reg_0215;
    101: op1_12_in11 = reg_1494;
    102: op1_12_in11 = reg_0158;
    103: op1_12_in11 = reg_0927;
    104: op1_12_in11 = reg_0712;
    105: op1_12_in11 = reg_0706;
    106: op1_12_in11 = reg_0206;
    47: op1_12_in11 = reg_0368;
    108: op1_12_in11 = reg_0557;
    109: op1_12_in11 = reg_1052;
    110: op1_12_in11 = reg_0370;
    111: op1_12_in11 = reg_0133;
    113: op1_12_in11 = reg_0973;
    114: op1_12_in11 = reg_0519;
    115: op1_12_in11 = reg_0276;
    116: op1_12_in11 = reg_0373;
    117: op1_12_in11 = reg_1235;
    119: op1_12_in11 = reg_0649;
    120: op1_12_in11 = reg_0701;
    122: op1_12_in11 = reg_1323;
    123: op1_12_in11 = reg_0168;
    124: op1_12_in11 = reg_0267;
    125: op1_12_in11 = reg_0954;
    44: op1_12_in11 = reg_0575;
    126: op1_12_in11 = reg_1432;
    127: op1_12_in11 = reg_0526;
    128: op1_12_in11 = reg_0116;
    130: op1_12_in11 = reg_0717;
    34: op1_12_in11 = reg_0053;
    default: op1_12_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv11 = 1;
    55: op1_12_inv11 = 1;
    74: op1_12_inv11 = 1;
    69: op1_12_inv11 = 1;
    54: op1_12_inv11 = 1;
    75: op1_12_inv11 = 1;
    56: op1_12_inv11 = 1;
    71: op1_12_inv11 = 1;
    87: op1_12_inv11 = 1;
    57: op1_12_inv11 = 1;
    77: op1_12_inv11 = 1;
    58: op1_12_inv11 = 1;
    78: op1_12_inv11 = 1;
    70: op1_12_inv11 = 1;
    59: op1_12_inv11 = 1;
    79: op1_12_inv11 = 1;
    51: op1_12_inv11 = 1;
    60: op1_12_inv11 = 1;
    81: op1_12_inv11 = 1;
    82: op1_12_inv11 = 1;
    83: op1_12_inv11 = 1;
    64: op1_12_inv11 = 1;
    89: op1_12_inv11 = 1;
    84: op1_12_inv11 = 1;
    90: op1_12_inv11 = 1;
    91: op1_12_inv11 = 1;
    67: op1_12_inv11 = 1;
    93: op1_12_inv11 = 1;
    94: op1_12_inv11 = 1;
    99: op1_12_inv11 = 1;
    100: op1_12_inv11 = 1;
    102: op1_12_inv11 = 1;
    103: op1_12_inv11 = 1;
    111: op1_12_inv11 = 1;
    113: op1_12_inv11 = 1;
    117: op1_12_inv11 = 1;
    118: op1_12_inv11 = 1;
    119: op1_12_inv11 = 1;
    120: op1_12_inv11 = 1;
    125: op1_12_inv11 = 1;
    126: op1_12_inv11 = 1;
    130: op1_12_inv11 = 1;
    34: op1_12_inv11 = 1;
    default: op1_12_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in12 = reg_0624;
    53: op1_12_in12 = reg_0041;
    55: op1_12_in12 = reg_0376;
    73: op1_12_in12 = reg_0565;
    86: op1_12_in12 = reg_0962;
    74: op1_12_in12 = reg_0409;
    69: op1_12_in12 = imem02_in[15:12];
    49: op1_12_in12 = reg_0017;
    54: op1_12_in12 = reg_0211;
    75: op1_12_in12 = reg_0718;
    56: op1_12_in12 = reg_0757;
    50: op1_12_in12 = imem07_in[3:0];
    76: op1_12_in12 = reg_1181;
    82: op1_12_in12 = reg_1181;
    84: op1_12_in12 = reg_1181;
    68: op1_12_in12 = reg_1339;
    71: op1_12_in12 = reg_1291;
    87: op1_12_in12 = reg_0049;
    57: op1_12_in12 = reg_1204;
    77: op1_12_in12 = reg_0617;
    61: op1_12_in12 = reg_0188;
    58: op1_12_in12 = reg_0970;
    78: op1_12_in12 = reg_1077;
    70: op1_12_in12 = reg_0975;
    59: op1_12_in12 = reg_0822;
    79: op1_12_in12 = reg_0023;
    51: op1_12_in12 = reg_0668;
    60: op1_12_in12 = imem01_in[7:4];
    88: op1_12_in12 = reg_0177;
    80: op1_12_in12 = imem01_in[15:12];
    62: op1_12_in12 = reg_0038;
    81: op1_12_in12 = reg_1515;
    52: op1_12_in12 = reg_0714;
    63: op1_12_in12 = reg_0939;
    46: op1_12_in12 = reg_0662;
    83: op1_12_in12 = reg_0057;
    64: op1_12_in12 = reg_0927;
    129: op1_12_in12 = reg_0927;
    89: op1_12_in12 = reg_0454;
    85: op1_12_in12 = reg_1518;
    65: op1_12_in12 = reg_0345;
    90: op1_12_in12 = reg_1203;
    48: op1_12_in12 = reg_0044;
    66: op1_12_in12 = reg_0619;
    116: op1_12_in12 = reg_0619;
    91: op1_12_in12 = reg_0496;
    67: op1_12_in12 = reg_0777;
    92: op1_12_in12 = reg_0203;
    93: op1_12_in12 = reg_0851;
    94: op1_12_in12 = reg_0831;
    95: op1_12_in12 = reg_0108;
    96: op1_12_in12 = reg_1346;
    97: op1_12_in12 = reg_0215;
    99: op1_12_in12 = reg_0495;
    100: op1_12_in12 = reg_0018;
    101: op1_12_in12 = reg_1516;
    102: op1_12_in12 = reg_0157;
    103: op1_12_in12 = reg_0722;
    104: op1_12_in12 = reg_0532;
    105: op1_12_in12 = reg_0216;
    106: op1_12_in12 = reg_0729;
    47: op1_12_in12 = reg_0835;
    108: op1_12_in12 = reg_0891;
    109: op1_12_in12 = reg_0293;
    110: op1_12_in12 = reg_1168;
    111: op1_12_in12 = reg_0712;
    112: op1_12_in12 = reg_0256;
    113: op1_12_in12 = reg_0876;
    114: op1_12_in12 = reg_1182;
    115: op1_12_in12 = reg_0588;
    117: op1_12_in12 = reg_0056;
    118: op1_12_in12 = reg_0070;
    119: op1_12_in12 = reg_0066;
    120: op1_12_in12 = reg_0182;
    122: op1_12_in12 = reg_0752;
    123: op1_12_in12 = reg_0632;
    124: op1_12_in12 = reg_1100;
    125: op1_12_in12 = reg_0627;
    44: op1_12_in12 = reg_0395;
    126: op1_12_in12 = reg_0229;
    127: op1_12_in12 = reg_1225;
    128: op1_12_in12 = reg_0374;
    130: op1_12_in12 = reg_0585;
    34: op1_12_in12 = reg_0086;
    default: op1_12_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv12 = 1;
    53: op1_12_inv12 = 1;
    69: op1_12_inv12 = 1;
    49: op1_12_inv12 = 1;
    54: op1_12_inv12 = 1;
    75: op1_12_inv12 = 1;
    77: op1_12_inv12 = 1;
    78: op1_12_inv12 = 1;
    79: op1_12_inv12 = 1;
    51: op1_12_inv12 = 1;
    60: op1_12_inv12 = 1;
    88: op1_12_inv12 = 1;
    62: op1_12_inv12 = 1;
    52: op1_12_inv12 = 1;
    82: op1_12_inv12 = 1;
    83: op1_12_inv12 = 1;
    64: op1_12_inv12 = 1;
    84: op1_12_inv12 = 1;
    85: op1_12_inv12 = 1;
    65: op1_12_inv12 = 1;
    91: op1_12_inv12 = 1;
    67: op1_12_inv12 = 1;
    93: op1_12_inv12 = 1;
    96: op1_12_inv12 = 1;
    100: op1_12_inv12 = 1;
    101: op1_12_inv12 = 1;
    102: op1_12_inv12 = 1;
    104: op1_12_inv12 = 1;
    106: op1_12_inv12 = 1;
    108: op1_12_inv12 = 1;
    109: op1_12_inv12 = 1;
    110: op1_12_inv12 = 1;
    111: op1_12_inv12 = 1;
    114: op1_12_inv12 = 1;
    115: op1_12_inv12 = 1;
    117: op1_12_inv12 = 1;
    118: op1_12_inv12 = 1;
    119: op1_12_inv12 = 1;
    120: op1_12_inv12 = 1;
    123: op1_12_inv12 = 1;
    125: op1_12_inv12 = 1;
    130: op1_12_inv12 = 1;
    default: op1_12_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in13 = reg_0323;
    53: op1_12_in13 = reg_0011;
    55: op1_12_in13 = reg_0177;
    73: op1_12_in13 = reg_1181;
    86: op1_12_in13 = reg_0145;
    74: op1_12_in13 = reg_0058;
    69: op1_12_in13 = reg_0138;
    49: op1_12_in13 = reg_0998;
    54: op1_12_in13 = reg_0209;
    75: op1_12_in13 = reg_0717;
    56: op1_12_in13 = reg_0234;
    50: op1_12_in13 = reg_0224;
    76: op1_12_in13 = reg_0118;
    68: op1_12_in13 = reg_1258;
    71: op1_12_in13 = reg_0260;
    87: op1_12_in13 = reg_0261;
    57: op1_12_in13 = reg_0271;
    77: op1_12_in13 = reg_0529;
    61: op1_12_in13 = reg_0389;
    58: op1_12_in13 = reg_0935;
    78: op1_12_in13 = reg_1082;
    70: op1_12_in13 = reg_1340;
    59: op1_12_in13 = reg_0474;
    79: op1_12_in13 = reg_0152;
    51: op1_12_in13 = reg_0605;
    60: op1_12_in13 = reg_1033;
    88: op1_12_in13 = reg_0962;
    80: op1_12_in13 = reg_1290;
    62: op1_12_in13 = reg_1036;
    81: op1_12_in13 = reg_0191;
    52: op1_12_in13 = reg_0617;
    63: op1_12_in13 = reg_0938;
    82: op1_12_in13 = reg_1180;
    46: op1_12_in13 = reg_0253;
    83: op1_12_in13 = reg_0166;
    64: op1_12_in13 = reg_0887;
    89: op1_12_in13 = reg_0582;
    84: op1_12_in13 = reg_1403;
    85: op1_12_in13 = reg_1314;
    101: op1_12_in13 = reg_1314;
    65: op1_12_in13 = reg_0296;
    90: op1_12_in13 = reg_0796;
    48: op1_12_in13 = reg_0012;
    66: op1_12_in13 = reg_0570;
    91: op1_12_in13 = imem02_in[3:0];
    67: op1_12_in13 = reg_0031;
    92: op1_12_in13 = reg_0985;
    93: op1_12_in13 = reg_1347;
    94: op1_12_in13 = reg_0066;
    95: op1_12_in13 = reg_1149;
    96: op1_12_in13 = reg_0344;
    97: op1_12_in13 = reg_0018;
    99: op1_12_in13 = reg_0776;
    100: op1_12_in13 = reg_1439;
    102: op1_12_in13 = reg_0489;
    103: op1_12_in13 = reg_0189;
    104: op1_12_in13 = reg_0390;
    105: op1_12_in13 = reg_0847;
    106: op1_12_in13 = reg_1064;
    47: op1_12_in13 = reg_0339;
    108: op1_12_in13 = reg_0556;
    109: op1_12_in13 = reg_1205;
    110: op1_12_in13 = reg_0793;
    111: op1_12_in13 = reg_1493;
    112: op1_12_in13 = reg_1146;
    113: op1_12_in13 = reg_0878;
    115: op1_12_in13 = reg_0561;
    116: op1_12_in13 = reg_0527;
    117: op1_12_in13 = reg_0712;
    118: op1_12_in13 = reg_1517;
    119: op1_12_in13 = reg_0173;
    120: op1_12_in13 = reg_0045;
    122: op1_12_in13 = reg_0827;
    123: op1_12_in13 = reg_0006;
    124: op1_12_in13 = reg_0635;
    125: op1_12_in13 = reg_0558;
    44: op1_12_in13 = reg_0748;
    126: op1_12_in13 = reg_0821;
    127: op1_12_in13 = reg_0119;
    128: op1_12_in13 = reg_0526;
    130: op1_12_in13 = reg_0526;
    129: op1_12_in13 = reg_0881;
    34: op1_12_in13 = reg_0518;
    default: op1_12_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_12_inv13 = 1;
    86: op1_12_inv13 = 1;
    74: op1_12_inv13 = 1;
    49: op1_12_inv13 = 1;
    54: op1_12_inv13 = 1;
    75: op1_12_inv13 = 1;
    56: op1_12_inv13 = 1;
    50: op1_12_inv13 = 1;
    57: op1_12_inv13 = 1;
    70: op1_12_inv13 = 1;
    59: op1_12_inv13 = 1;
    88: op1_12_inv13 = 1;
    62: op1_12_inv13 = 1;
    63: op1_12_inv13 = 1;
    46: op1_12_inv13 = 1;
    83: op1_12_inv13 = 1;
    64: op1_12_inv13 = 1;
    93: op1_12_inv13 = 1;
    94: op1_12_inv13 = 1;
    95: op1_12_inv13 = 1;
    97: op1_12_inv13 = 1;
    100: op1_12_inv13 = 1;
    101: op1_12_inv13 = 1;
    102: op1_12_inv13 = 1;
    103: op1_12_inv13 = 1;
    47: op1_12_inv13 = 1;
    110: op1_12_inv13 = 1;
    112: op1_12_inv13 = 1;
    113: op1_12_inv13 = 1;
    120: op1_12_inv13 = 1;
    44: op1_12_inv13 = 1;
    129: op1_12_inv13 = 1;
    default: op1_12_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in14 = reg_0165;
    53: op1_12_in14 = reg_0662;
    55: op1_12_in14 = reg_1000;
    73: op1_12_in14 = reg_0541;
    86: op1_12_in14 = reg_0144;
    88: op1_12_in14 = reg_0144;
    74: op1_12_in14 = reg_0786;
    69: op1_12_in14 = reg_0379;
    49: op1_12_in14 = reg_0703;
    54: op1_12_in14 = reg_0064;
    75: op1_12_in14 = reg_1302;
    56: op1_12_in14 = reg_0185;
    50: op1_12_in14 = reg_0299;
    76: op1_12_in14 = reg_0797;
    68: op1_12_in14 = reg_0466;
    71: op1_12_in14 = reg_0746;
    87: op1_12_in14 = reg_0378;
    57: op1_12_in14 = reg_0215;
    77: op1_12_in14 = reg_0570;
    130: op1_12_in14 = reg_0570;
    61: op1_12_in14 = reg_0072;
    58: op1_12_in14 = reg_0933;
    78: op1_12_in14 = reg_0412;
    90: op1_12_in14 = reg_0412;
    70: op1_12_in14 = reg_1215;
    59: op1_12_in14 = reg_0472;
    79: op1_12_in14 = reg_0018;
    51: op1_12_in14 = reg_0607;
    60: op1_12_in14 = reg_1031;
    80: op1_12_in14 = reg_0785;
    92: op1_12_in14 = reg_0785;
    62: op1_12_in14 = reg_1035;
    81: op1_12_in14 = reg_0233;
    52: op1_12_in14 = reg_0583;
    63: op1_12_in14 = reg_0070;
    82: op1_12_in14 = reg_1404;
    46: op1_12_in14 = reg_0605;
    83: op1_12_in14 = reg_1513;
    64: op1_12_in14 = reg_0886;
    89: op1_12_in14 = reg_0096;
    84: op1_12_in14 = reg_0939;
    85: op1_12_in14 = reg_0627;
    65: op1_12_in14 = reg_0295;
    66: op1_12_in14 = reg_0295;
    48: op1_12_in14 = reg_0013;
    91: op1_12_in14 = imem02_in[15:12];
    67: op1_12_in14 = reg_0030;
    93: op1_12_in14 = reg_0777;
    102: op1_12_in14 = reg_0777;
    94: op1_12_in14 = reg_0562;
    95: op1_12_in14 = reg_0348;
    96: op1_12_in14 = reg_0038;
    97: op1_12_in14 = reg_0022;
    99: op1_12_in14 = reg_1450;
    100: op1_12_in14 = reg_1414;
    101: op1_12_in14 = reg_0957;
    103: op1_12_in14 = reg_0435;
    104: op1_12_in14 = reg_1002;
    105: op1_12_in14 = reg_0312;
    106: op1_12_in14 = reg_0795;
    47: op1_12_in14 = reg_0208;
    108: op1_12_in14 = reg_0142;
    109: op1_12_in14 = reg_0155;
    110: op1_12_in14 = reg_1430;
    111: op1_12_in14 = reg_0822;
    112: op1_12_in14 = reg_0338;
    113: op1_12_in14 = reg_0897;
    115: op1_12_in14 = reg_0839;
    117: op1_12_in14 = reg_0839;
    116: op1_12_in14 = reg_0979;
    118: op1_12_in14 = reg_1314;
    119: op1_12_in14 = reg_0940;
    120: op1_12_in14 = reg_0630;
    122: op1_12_in14 = reg_1505;
    123: op1_12_in14 = reg_0049;
    124: op1_12_in14 = reg_0120;
    125: op1_12_in14 = reg_1231;
    44: op1_12_in14 = reg_0737;
    126: op1_12_in14 = reg_0476;
    127: op1_12_in14 = reg_0023;
    128: op1_12_in14 = reg_0571;
    129: op1_12_in14 = reg_0883;
    34: op1_12_in14 = reg_0124;
    default: op1_12_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv14 = 1;
    73: op1_12_inv14 = 1;
    74: op1_12_inv14 = 1;
    49: op1_12_inv14 = 1;
    54: op1_12_inv14 = 1;
    75: op1_12_inv14 = 1;
    56: op1_12_inv14 = 1;
    76: op1_12_inv14 = 1;
    68: op1_12_inv14 = 1;
    71: op1_12_inv14 = 1;
    78: op1_12_inv14 = 1;
    70: op1_12_inv14 = 1;
    60: op1_12_inv14 = 1;
    80: op1_12_inv14 = 1;
    81: op1_12_inv14 = 1;
    63: op1_12_inv14 = 1;
    46: op1_12_inv14 = 1;
    83: op1_12_inv14 = 1;
    64: op1_12_inv14 = 1;
    89: op1_12_inv14 = 1;
    85: op1_12_inv14 = 1;
    65: op1_12_inv14 = 1;
    48: op1_12_inv14 = 1;
    67: op1_12_inv14 = 1;
    92: op1_12_inv14 = 1;
    93: op1_12_inv14 = 1;
    95: op1_12_inv14 = 1;
    99: op1_12_inv14 = 1;
    100: op1_12_inv14 = 1;
    101: op1_12_inv14 = 1;
    102: op1_12_inv14 = 1;
    104: op1_12_inv14 = 1;
    105: op1_12_inv14 = 1;
    110: op1_12_inv14 = 1;
    111: op1_12_inv14 = 1;
    112: op1_12_inv14 = 1;
    118: op1_12_inv14 = 1;
    122: op1_12_inv14 = 1;
    124: op1_12_inv14 = 1;
    125: op1_12_inv14 = 1;
    44: op1_12_inv14 = 1;
    126: op1_12_inv14 = 1;
    127: op1_12_inv14 = 1;
    129: op1_12_inv14 = 1;
    34: op1_12_inv14 = 1;
    default: op1_12_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in15 = reg_0371;
    53: op1_12_in15 = reg_0820;
    55: op1_12_in15 = reg_0964;
    73: op1_12_in15 = reg_0539;
    86: op1_12_in15 = reg_1516;
    74: op1_12_in15 = reg_0785;
    69: op1_12_in15 = reg_0069;
    49: op1_12_in15 = reg_0674;
    54: op1_12_in15 = reg_0063;
    75: op1_12_in15 = reg_0636;
    56: op1_12_in15 = reg_0179;
    50: op1_12_in15 = reg_0170;
    76: op1_12_in15 = reg_0449;
    68: op1_12_in15 = reg_0552;
    71: op1_12_in15 = reg_0420;
    87: op1_12_in15 = reg_0541;
    57: op1_12_in15 = reg_1150;
    77: op1_12_in15 = reg_0289;
    61: op1_12_in15 = reg_0075;
    58: op1_12_in15 = reg_0125;
    78: op1_12_in15 = reg_0796;
    70: op1_12_in15 = reg_1077;
    59: op1_12_in15 = reg_0429;
    79: op1_12_in15 = reg_0034;
    51: op1_12_in15 = reg_0608;
    60: op1_12_in15 = reg_0257;
    88: op1_12_in15 = reg_0000;
    80: op1_12_in15 = reg_0549;
    62: op1_12_in15 = reg_0753;
    81: op1_12_in15 = reg_0699;
    52: op1_12_in15 = reg_0570;
    63: op1_12_in15 = reg_0418;
    82: op1_12_in15 = reg_0939;
    46: op1_12_in15 = reg_0472;
    83: op1_12_in15 = reg_0093;
    64: op1_12_in15 = reg_0189;
    129: op1_12_in15 = reg_0189;
    89: op1_12_in15 = reg_0065;
    84: op1_12_in15 = reg_0937;
    85: op1_12_in15 = reg_0329;
    108: op1_12_in15 = reg_0329;
    65: op1_12_in15 = reg_0067;
    90: op1_12_in15 = reg_0969;
    48: op1_12_in15 = reg_0662;
    66: op1_12_in15 = reg_0119;
    116: op1_12_in15 = reg_0119;
    91: op1_12_in15 = reg_1098;
    67: op1_12_in15 = reg_0366;
    92: op1_12_in15 = reg_1512;
    93: op1_12_in15 = reg_0779;
    94: op1_12_in15 = reg_0701;
    95: op1_12_in15 = reg_0252;
    96: op1_12_in15 = reg_1058;
    97: op1_12_in15 = reg_1170;
    99: op1_12_in15 = reg_0128;
    100: op1_12_in15 = reg_0994;
    101: op1_12_in15 = reg_0220;
    102: op1_12_in15 = reg_0030;
    103: op1_12_in15 = reg_0203;
    104: op1_12_in15 = reg_0256;
    105: op1_12_in15 = reg_0234;
    106: op1_12_in15 = reg_0906;
    47: op1_12_in15 = reg_0064;
    109: op1_12_in15 = reg_1418;
    110: op1_12_in15 = reg_0278;
    111: op1_12_in15 = reg_1207;
    112: op1_12_in15 = reg_0367;
    113: op1_12_in15 = reg_0560;
    115: op1_12_in15 = reg_0532;
    117: op1_12_in15 = reg_0390;
    118: op1_12_in15 = reg_1313;
    119: op1_12_in15 = reg_1070;
    120: op1_12_in15 = reg_1402;
    122: op1_12_in15 = reg_1504;
    123: op1_12_in15 = reg_0330;
    124: op1_12_in15 = reg_0550;
    125: op1_12_in15 = reg_0178;
    44: op1_12_in15 = reg_0347;
    126: op1_12_in15 = reg_0928;
    127: op1_12_in15 = reg_0518;
    128: op1_12_in15 = reg_0569;
    130: op1_12_in15 = reg_0323;
    default: op1_12_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv15 = 1;
    53: op1_12_inv15 = 1;
    86: op1_12_inv15 = 1;
    54: op1_12_inv15 = 1;
    56: op1_12_inv15 = 1;
    76: op1_12_inv15 = 1;
    71: op1_12_inv15 = 1;
    87: op1_12_inv15 = 1;
    77: op1_12_inv15 = 1;
    61: op1_12_inv15 = 1;
    60: op1_12_inv15 = 1;
    88: op1_12_inv15 = 1;
    80: op1_12_inv15 = 1;
    62: op1_12_inv15 = 1;
    52: op1_12_inv15 = 1;
    84: op1_12_inv15 = 1;
    65: op1_12_inv15 = 1;
    90: op1_12_inv15 = 1;
    48: op1_12_inv15 = 1;
    66: op1_12_inv15 = 1;
    91: op1_12_inv15 = 1;
    92: op1_12_inv15 = 1;
    93: op1_12_inv15 = 1;
    94: op1_12_inv15 = 1;
    95: op1_12_inv15 = 1;
    97: op1_12_inv15 = 1;
    101: op1_12_inv15 = 1;
    106: op1_12_inv15 = 1;
    47: op1_12_inv15 = 1;
    108: op1_12_inv15 = 1;
    110: op1_12_inv15 = 1;
    111: op1_12_inv15 = 1;
    112: op1_12_inv15 = 1;
    113: op1_12_inv15 = 1;
    115: op1_12_inv15 = 1;
    120: op1_12_inv15 = 1;
    123: op1_12_inv15 = 1;
    124: op1_12_inv15 = 1;
    125: op1_12_inv15 = 1;
    127: op1_12_inv15 = 1;
    129: op1_12_inv15 = 1;
    default: op1_12_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in16 = reg_1179;
    53: op1_12_in16 = reg_0606;
    55: op1_12_in16 = reg_0952;
    118: op1_12_in16 = reg_0952;
    73: op1_12_in16 = reg_0167;
    86: op1_12_in16 = reg_1314;
    74: op1_12_in16 = reg_1291;
    69: op1_12_in16 = reg_0280;
    49: op1_12_in16 = imem07_in[7:4];
    54: op1_12_in16 = reg_0391;
    75: op1_12_in16 = reg_0141;
    56: op1_12_in16 = reg_0180;
    50: op1_12_in16 = reg_0309;
    76: op1_12_in16 = reg_0151;
    68: op1_12_in16 = reg_1147;
    71: op1_12_in16 = reg_0438;
    87: op1_12_in16 = reg_0000;
    57: op1_12_in16 = reg_0229;
    77: op1_12_in16 = reg_1204;
    61: op1_12_in16 = reg_0267;
    58: op1_12_in16 = reg_0900;
    78: op1_12_in16 = reg_1233;
    70: op1_12_in16 = reg_0552;
    59: op1_12_in16 = reg_0380;
    79: op1_12_in16 = reg_0185;
    51: op1_12_in16 = reg_0253;
    60: op1_12_in16 = reg_0550;
    88: op1_12_in16 = reg_1003;
    80: op1_12_in16 = reg_0548;
    83: op1_12_in16 = reg_0548;
    62: op1_12_in16 = reg_0783;
    81: op1_12_in16 = reg_0227;
    52: op1_12_in16 = reg_0528;
    63: op1_12_in16 = reg_0896;
    82: op1_12_in16 = reg_0794;
    46: op1_12_in16 = reg_0054;
    64: op1_12_in16 = reg_0405;
    109: op1_12_in16 = reg_0405;
    89: op1_12_in16 = imem05_in[3:0];
    84: op1_12_in16 = reg_0300;
    85: op1_12_in16 = reg_1301;
    65: op1_12_in16 = reg_1150;
    90: op1_12_in16 = reg_0232;
    48: op1_12_in16 = reg_0666;
    66: op1_12_in16 = reg_0269;
    91: op1_12_in16 = reg_0008;
    67: op1_12_in16 = reg_0442;
    92: op1_12_in16 = reg_0093;
    93: op1_12_in16 = reg_0284;
    94: op1_12_in16 = reg_0182;
    95: op1_12_in16 = reg_0341;
    96: op1_12_in16 = reg_0193;
    97: op1_12_in16 = reg_0995;
    99: op1_12_in16 = reg_0127;
    100: op1_12_in16 = reg_0298;
    101: op1_12_in16 = reg_0246;
    102: op1_12_in16 = reg_0441;
    103: op1_12_in16 = reg_1290;
    104: op1_12_in16 = reg_0495;
    105: op1_12_in16 = reg_1494;
    106: op1_12_in16 = reg_0960;
    47: op1_12_in16 = reg_0062;
    108: op1_12_in16 = reg_1199;
    110: op1_12_in16 = reg_0333;
    111: op1_12_in16 = reg_0432;
    112: op1_12_in16 = reg_0833;
    113: op1_12_in16 = reg_1098;
    115: op1_12_in16 = reg_0497;
    116: op1_12_in16 = reg_0195;
    117: op1_12_in16 = reg_0494;
    119: op1_12_in16 = reg_1514;
    120: op1_12_in16 = reg_0792;
    122: op1_12_in16 = reg_1508;
    123: op1_12_in16 = reg_1000;
    124: op1_12_in16 = reg_0222;
    125: op1_12_in16 = reg_1208;
    44: op1_12_in16 = reg_0523;
    126: op1_12_in16 = reg_0886;
    127: op1_12_in16 = reg_0169;
    128: op1_12_in16 = reg_0522;
    129: op1_12_in16 = reg_0410;
    130: op1_12_in16 = reg_0977;
    default: op1_12_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv16 = 1;
    53: op1_12_inv16 = 1;
    69: op1_12_inv16 = 1;
    54: op1_12_inv16 = 1;
    56: op1_12_inv16 = 1;
    76: op1_12_inv16 = 1;
    68: op1_12_inv16 = 1;
    71: op1_12_inv16 = 1;
    87: op1_12_inv16 = 1;
    57: op1_12_inv16 = 1;
    77: op1_12_inv16 = 1;
    78: op1_12_inv16 = 1;
    59: op1_12_inv16 = 1;
    88: op1_12_inv16 = 1;
    80: op1_12_inv16 = 1;
    81: op1_12_inv16 = 1;
    63: op1_12_inv16 = 1;
    82: op1_12_inv16 = 1;
    65: op1_12_inv16 = 1;
    66: op1_12_inv16 = 1;
    91: op1_12_inv16 = 1;
    92: op1_12_inv16 = 1;
    97: op1_12_inv16 = 1;
    103: op1_12_inv16 = 1;
    104: op1_12_inv16 = 1;
    105: op1_12_inv16 = 1;
    106: op1_12_inv16 = 1;
    47: op1_12_inv16 = 1;
    108: op1_12_inv16 = 1;
    109: op1_12_inv16 = 1;
    112: op1_12_inv16 = 1;
    115: op1_12_inv16 = 1;
    118: op1_12_inv16 = 1;
    119: op1_12_inv16 = 1;
    120: op1_12_inv16 = 1;
    122: op1_12_inv16 = 1;
    44: op1_12_inv16 = 1;
    127: op1_12_inv16 = 1;
    129: op1_12_inv16 = 1;
    default: op1_12_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in17 = reg_0269;
    53: op1_12_in17 = reg_0607;
    55: op1_12_in17 = reg_0597;
    73: op1_12_in17 = reg_0477;
    86: op1_12_in17 = reg_0957;
    74: op1_12_in17 = reg_1255;
    69: op1_12_in17 = reg_1132;
    49: op1_12_in17 = reg_0169;
    54: op1_12_in17 = reg_0750;
    75: op1_12_in17 = reg_0585;
    56: op1_12_in17 = reg_1000;
    50: op1_12_in17 = reg_0851;
    76: op1_12_in17 = reg_0828;
    68: op1_12_in17 = reg_0414;
    71: op1_12_in17 = reg_0383;
    87: op1_12_in17 = reg_0891;
    57: op1_12_in17 = reg_1095;
    77: op1_12_in17 = reg_1441;
    61: op1_12_in17 = imem00_in[3:0];
    58: op1_12_in17 = reg_0708;
    78: op1_12_in17 = reg_0454;
    70: op1_12_in17 = reg_0407;
    59: op1_12_in17 = reg_0056;
    79: op1_12_in17 = reg_1439;
    51: op1_12_in17 = reg_0587;
    60: op1_12_in17 = reg_0238;
    88: op1_12_in17 = reg_0070;
    105: op1_12_in17 = reg_0070;
    80: op1_12_in17 = reg_0747;
    62: op1_12_in17 = reg_0730;
    81: op1_12_in17 = reg_0154;
    52: op1_12_in17 = reg_0419;
    63: op1_12_in17 = reg_0873;
    82: op1_12_in17 = reg_0450;
    46: op1_12_in17 = imem02_in[7:4];
    83: op1_12_in17 = reg_0242;
    64: op1_12_in17 = reg_0267;
    89: op1_12_in17 = imem05_in[7:4];
    84: op1_12_in17 = reg_0151;
    85: op1_12_in17 = reg_0178;
    65: op1_12_in17 = reg_0998;
    90: op1_12_in17 = reg_0698;
    48: op1_12_in17 = reg_0254;
    66: op1_12_in17 = reg_0214;
    91: op1_12_in17 = reg_1006;
    113: op1_12_in17 = reg_1006;
    67: op1_12_in17 = reg_0100;
    92: op1_12_in17 = reg_0610;
    93: op1_12_in17 = reg_0103;
    94: op1_12_in17 = reg_0630;
    95: op1_12_in17 = reg_1367;
    96: op1_12_in17 = reg_0795;
    97: op1_12_in17 = reg_0994;
    99: op1_12_in17 = reg_0105;
    100: op1_12_in17 = reg_0892;
    101: op1_12_in17 = reg_1301;
    102: op1_12_in17 = reg_0740;
    103: op1_12_in17 = reg_0553;
    104: op1_12_in17 = reg_1207;
    106: op1_12_in17 = reg_1420;
    47: op1_12_in17 = reg_0016;
    108: op1_12_in17 = reg_0107;
    109: op1_12_in17 = reg_0071;
    110: op1_12_in17 = reg_0395;
    111: op1_12_in17 = reg_0433;
    112: op1_12_in17 = reg_0702;
    115: op1_12_in17 = reg_0054;
    116: op1_12_in17 = reg_0977;
    117: op1_12_in17 = reg_1455;
    118: op1_12_in17 = reg_1300;
    119: op1_12_in17 = reg_0303;
    120: op1_12_in17 = reg_0197;
    122: op1_12_in17 = reg_0115;
    123: op1_12_in17 = reg_1063;
    124: op1_12_in17 = reg_0239;
    125: op1_12_in17 = reg_0025;
    44: op1_12_in17 = reg_0445;
    126: op1_12_in17 = reg_0202;
    127: op1_12_in17 = reg_0867;
    128: op1_12_in17 = reg_0213;
    129: op1_12_in17 = reg_0134;
    130: op1_12_in17 = reg_0394;
    default: op1_12_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_12_inv17 = 1;
    74: op1_12_inv17 = 1;
    69: op1_12_inv17 = 1;
    75: op1_12_inv17 = 1;
    56: op1_12_inv17 = 1;
    50: op1_12_inv17 = 1;
    87: op1_12_inv17 = 1;
    77: op1_12_inv17 = 1;
    58: op1_12_inv17 = 1;
    51: op1_12_inv17 = 1;
    88: op1_12_inv17 = 1;
    80: op1_12_inv17 = 1;
    81: op1_12_inv17 = 1;
    52: op1_12_inv17 = 1;
    63: op1_12_inv17 = 1;
    82: op1_12_inv17 = 1;
    46: op1_12_inv17 = 1;
    64: op1_12_inv17 = 1;
    89: op1_12_inv17 = 1;
    85: op1_12_inv17 = 1;
    48: op1_12_inv17 = 1;
    66: op1_12_inv17 = 1;
    91: op1_12_inv17 = 1;
    67: op1_12_inv17 = 1;
    92: op1_12_inv17 = 1;
    95: op1_12_inv17 = 1;
    96: op1_12_inv17 = 1;
    97: op1_12_inv17 = 1;
    99: op1_12_inv17 = 1;
    100: op1_12_inv17 = 1;
    101: op1_12_inv17 = 1;
    105: op1_12_inv17 = 1;
    108: op1_12_inv17 = 1;
    109: op1_12_inv17 = 1;
    110: op1_12_inv17 = 1;
    112: op1_12_inv17 = 1;
    115: op1_12_inv17 = 1;
    118: op1_12_inv17 = 1;
    119: op1_12_inv17 = 1;
    122: op1_12_inv17 = 1;
    123: op1_12_inv17 = 1;
    125: op1_12_inv17 = 1;
    126: op1_12_inv17 = 1;
    127: op1_12_inv17 = 1;
    128: op1_12_inv17 = 1;
    129: op1_12_inv17 = 1;
    default: op1_12_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in18 = imem07_in[7:4];
    53: op1_12_in18 = reg_1018;
    55: op1_12_in18 = reg_0559;
    73: op1_12_in18 = reg_0070;
    86: op1_12_in18 = reg_1208;
    74: op1_12_in18 = reg_1068;
    69: op1_12_in18 = reg_0758;
    49: op1_12_in18 = reg_0140;
    54: op1_12_in18 = reg_0832;
    75: op1_12_in18 = reg_0622;
    56: op1_12_in18 = reg_0952;
    50: op1_12_in18 = reg_0186;
    76: op1_12_in18 = reg_0014;
    68: op1_12_in18 = reg_0406;
    71: op1_12_in18 = reg_0724;
    87: op1_12_in18 = reg_0989;
    57: op1_12_in18 = imem07_in[3:0];
    77: op1_12_in18 = reg_0490;
    61: op1_12_in18 = imem01_in[15:12];
    58: op1_12_in18 = reg_0068;
    78: op1_12_in18 = reg_0451;
    70: op1_12_in18 = reg_0969;
    59: op1_12_in18 = reg_0897;
    79: op1_12_in18 = reg_0297;
    51: op1_12_in18 = reg_0981;
    60: op1_12_in18 = reg_0241;
    92: op1_12_in18 = reg_0241;
    88: op1_12_in18 = reg_0190;
    80: op1_12_in18 = reg_0222;
    62: op1_12_in18 = reg_0696;
    81: op1_12_in18 = reg_0444;
    52: op1_12_in18 = reg_0458;
    63: op1_12_in18 = reg_0243;
    82: op1_12_in18 = reg_0090;
    46: op1_12_in18 = reg_0934;
    83: op1_12_in18 = reg_1475;
    64: op1_12_in18 = reg_1100;
    89: op1_12_in18 = reg_0579;
    84: op1_12_in18 = reg_0828;
    85: op1_12_in18 = reg_0481;
    65: op1_12_in18 = reg_1183;
    66: op1_12_in18 = reg_1183;
    90: op1_12_in18 = reg_0304;
    48: op1_12_in18 = imem02_in[15:12];
    91: op1_12_in18 = reg_0999;
    67: op1_12_in18 = reg_0028;
    93: op1_12_in18 = reg_0114;
    94: op1_12_in18 = reg_1181;
    95: op1_12_in18 = reg_0493;
    96: op1_12_in18 = reg_0905;
    97: op1_12_in18 = reg_0298;
    99: op1_12_in18 = reg_1433;
    100: op1_12_in18 = reg_0310;
    101: op1_12_in18 = reg_1199;
    102: op1_12_in18 = reg_0413;
    103: op1_12_in18 = reg_0242;
    104: op1_12_in18 = reg_0433;
    105: op1_12_in18 = reg_1518;
    123: op1_12_in18 = reg_1518;
    106: op1_12_in18 = reg_0984;
    47: op1_12_in18 = reg_0033;
    108: op1_12_in18 = reg_0113;
    109: op1_12_in18 = reg_0059;
    110: op1_12_in18 = reg_0346;
    111: op1_12_in18 = reg_0496;
    112: op1_12_in18 = reg_0251;
    113: op1_12_in18 = reg_0759;
    115: op1_12_in18 = reg_0971;
    116: op1_12_in18 = reg_0212;
    117: op1_12_in18 = reg_0382;
    118: op1_12_in18 = reg_0048;
    119: op1_12_in18 = reg_0300;
    120: op1_12_in18 = reg_0240;
    122: op1_12_in18 = reg_0718;
    124: op1_12_in18 = reg_0830;
    125: op1_12_in18 = reg_0291;
    44: op1_12_in18 = reg_0648;
    126: op1_12_in18 = reg_0353;
    127: op1_12_in18 = reg_0225;
    128: op1_12_in18 = reg_0051;
    129: op1_12_in18 = reg_0238;
    130: op1_12_in18 = reg_1057;
    default: op1_12_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv18 = 1;
    53: op1_12_inv18 = 1;
    55: op1_12_inv18 = 1;
    73: op1_12_inv18 = 1;
    86: op1_12_inv18 = 1;
    69: op1_12_inv18 = 1;
    54: op1_12_inv18 = 1;
    75: op1_12_inv18 = 1;
    50: op1_12_inv18 = 1;
    87: op1_12_inv18 = 1;
    61: op1_12_inv18 = 1;
    58: op1_12_inv18 = 1;
    70: op1_12_inv18 = 1;
    80: op1_12_inv18 = 1;
    52: op1_12_inv18 = 1;
    82: op1_12_inv18 = 1;
    83: op1_12_inv18 = 1;
    89: op1_12_inv18 = 1;
    84: op1_12_inv18 = 1;
    90: op1_12_inv18 = 1;
    66: op1_12_inv18 = 1;
    91: op1_12_inv18 = 1;
    67: op1_12_inv18 = 1;
    92: op1_12_inv18 = 1;
    93: op1_12_inv18 = 1;
    94: op1_12_inv18 = 1;
    95: op1_12_inv18 = 1;
    96: op1_12_inv18 = 1;
    97: op1_12_inv18 = 1;
    101: op1_12_inv18 = 1;
    103: op1_12_inv18 = 1;
    105: op1_12_inv18 = 1;
    106: op1_12_inv18 = 1;
    47: op1_12_inv18 = 1;
    110: op1_12_inv18 = 1;
    111: op1_12_inv18 = 1;
    113: op1_12_inv18 = 1;
    116: op1_12_inv18 = 1;
    117: op1_12_inv18 = 1;
    119: op1_12_inv18 = 1;
    120: op1_12_inv18 = 1;
    122: op1_12_inv18 = 1;
    123: op1_12_inv18 = 1;
    126: op1_12_inv18 = 1;
    128: op1_12_inv18 = 1;
    default: op1_12_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in19 = imem07_in[15:12];
    57: op1_12_in19 = imem07_in[15:12];
    53: op1_12_in19 = reg_0561;
    48: op1_12_in19 = reg_0561;
    55: op1_12_in19 = reg_0505;
    73: op1_12_in19 = reg_1346;
    86: op1_12_in19 = reg_0885;
    74: op1_12_in19 = imem01_in[7:4];
    69: op1_12_in19 = reg_0630;
    49: op1_12_in19 = reg_0663;
    54: op1_12_in19 = reg_0700;
    75: op1_12_in19 = reg_0619;
    56: op1_12_in19 = reg_0246;
    50: op1_12_in19 = reg_0924;
    76: op1_12_in19 = reg_0751;
    68: op1_12_in19 = reg_0969;
    71: op1_12_in19 = reg_0896;
    87: op1_12_in19 = reg_0314;
    77: op1_12_in19 = reg_0162;
    61: op1_12_in19 = reg_0166;
    58: op1_12_in19 = reg_0217;
    78: op1_12_in19 = reg_0342;
    70: op1_12_in19 = reg_0797;
    59: op1_12_in19 = reg_0903;
    79: op1_12_in19 = reg_0156;
    51: op1_12_in19 = reg_0990;
    60: op1_12_in19 = reg_0553;
    88: op1_12_in19 = reg_0329;
    80: op1_12_in19 = reg_0239;
    62: op1_12_in19 = reg_0870;
    81: op1_12_in19 = reg_0707;
    52: op1_12_in19 = reg_0067;
    63: op1_12_in19 = reg_0240;
    82: op1_12_in19 = reg_1484;
    46: op1_12_in19 = reg_0105;
    83: op1_12_in19 = reg_0468;
    64: op1_12_in19 = reg_1254;
    89: op1_12_in19 = reg_0735;
    84: op1_12_in19 = reg_0466;
    85: op1_12_in19 = reg_0478;
    65: op1_12_in19 = imem07_in[3:0];
    90: op1_12_in19 = reg_0339;
    66: op1_12_in19 = reg_0667;
    91: op1_12_in19 = reg_0889;
    67: op1_12_in19 = reg_0361;
    92: op1_12_in19 = reg_0830;
    103: op1_12_in19 = reg_0830;
    93: op1_12_in19 = reg_0052;
    94: op1_12_in19 = reg_0872;
    95: op1_12_in19 = reg_0264;
    96: op1_12_in19 = reg_0960;
    97: op1_12_in19 = reg_0894;
    99: op1_12_in19 = reg_0306;
    100: op1_12_in19 = reg_0703;
    101: op1_12_in19 = reg_1092;
    102: op1_12_in19 = reg_0591;
    104: op1_12_in19 = reg_1455;
    105: op1_12_in19 = reg_0957;
    106: op1_12_in19 = reg_1326;
    47: op1_12_in19 = reg_0034;
    108: op1_12_in19 = reg_0448;
    109: op1_12_in19 = reg_1322;
    110: op1_12_in19 = reg_0272;
    111: op1_12_in19 = reg_0745;
    112: op1_12_in19 = reg_0066;
    113: op1_12_in19 = reg_1145;
    115: op1_12_in19 = reg_1458;
    116: op1_12_in19 = reg_0015;
    117: op1_12_in19 = reg_1140;
    118: op1_12_in19 = reg_1208;
    119: op1_12_in19 = reg_0301;
    120: op1_12_in19 = reg_1348;
    122: op1_12_in19 = reg_0194;
    123: op1_12_in19 = reg_1517;
    124: op1_12_in19 = reg_1473;
    125: op1_12_in19 = reg_0288;
    44: op1_12_in19 = reg_0601;
    126: op1_12_in19 = reg_0188;
    127: op1_12_in19 = reg_0457;
    128: op1_12_in19 = reg_1095;
    129: op1_12_in19 = reg_0577;
    130: op1_12_in19 = reg_0225;
    default: op1_12_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv19 = 1;
    73: op1_12_inv19 = 1;
    86: op1_12_inv19 = 1;
    69: op1_12_inv19 = 1;
    54: op1_12_inv19 = 1;
    75: op1_12_inv19 = 1;
    56: op1_12_inv19 = 1;
    50: op1_12_inv19 = 1;
    71: op1_12_inv19 = 1;
    87: op1_12_inv19 = 1;
    57: op1_12_inv19 = 1;
    58: op1_12_inv19 = 1;
    78: op1_12_inv19 = 1;
    70: op1_12_inv19 = 1;
    88: op1_12_inv19 = 1;
    80: op1_12_inv19 = 1;
    62: op1_12_inv19 = 1;
    81: op1_12_inv19 = 1;
    52: op1_12_inv19 = 1;
    63: op1_12_inv19 = 1;
    46: op1_12_inv19 = 1;
    64: op1_12_inv19 = 1;
    89: op1_12_inv19 = 1;
    84: op1_12_inv19 = 1;
    85: op1_12_inv19 = 1;
    90: op1_12_inv19 = 1;
    91: op1_12_inv19 = 1;
    67: op1_12_inv19 = 1;
    92: op1_12_inv19 = 1;
    94: op1_12_inv19 = 1;
    99: op1_12_inv19 = 1;
    100: op1_12_inv19 = 1;
    101: op1_12_inv19 = 1;
    102: op1_12_inv19 = 1;
    106: op1_12_inv19 = 1;
    47: op1_12_inv19 = 1;
    112: op1_12_inv19 = 1;
    113: op1_12_inv19 = 1;
    115: op1_12_inv19 = 1;
    117: op1_12_inv19 = 1;
    119: op1_12_inv19 = 1;
    120: op1_12_inv19 = 1;
    122: op1_12_inv19 = 1;
    123: op1_12_inv19 = 1;
    126: op1_12_inv19 = 1;
    127: op1_12_inv19 = 1;
    129: op1_12_inv19 = 1;
    130: op1_12_inv19 = 1;
    default: op1_12_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in20 = reg_1416;
    53: op1_12_in20 = imem02_in[3:0];
    55: op1_12_in20 = reg_0328;
    73: op1_12_in20 = reg_0631;
    86: op1_12_in20 = imem03_in[11:8];
    74: op1_12_in20 = imem01_in[15:12];
    69: op1_12_in20 = reg_0678;
    49: op1_12_in20 = reg_0366;
    54: op1_12_in20 = reg_1164;
    75: op1_12_in20 = reg_0526;
    56: op1_12_in20 = reg_0891;
    50: op1_12_in20 = reg_0489;
    76: op1_12_in20 = reg_0120;
    68: op1_12_in20 = reg_0471;
    71: op1_12_in20 = reg_0874;
    87: op1_12_in20 = reg_1314;
    57: op1_12_in20 = reg_0496;
    77: op1_12_in20 = reg_0851;
    61: op1_12_in20 = reg_0788;
    58: op1_12_in20 = reg_0325;
    78: op1_12_in20 = reg_0698;
    70: op1_12_in20 = imem04_in[7:4];
    59: op1_12_in20 = reg_0878;
    79: op1_12_in20 = reg_1094;
    51: op1_12_in20 = reg_0934;
    60: op1_12_in20 = reg_0982;
    88: op1_12_in20 = reg_1231;
    80: op1_12_in20 = reg_0896;
    62: op1_12_in20 = reg_0860;
    81: op1_12_in20 = reg_0145;
    52: op1_12_in20 = reg_0152;
    63: op1_12_in20 = imem05_in[3:0];
    82: op1_12_in20 = reg_0197;
    46: op1_12_in20 = reg_0294;
    83: op1_12_in20 = reg_0968;
    64: op1_12_in20 = reg_0259;
    89: op1_12_in20 = reg_0136;
    84: op1_12_in20 = reg_1437;
    85: op1_12_in20 = reg_0525;
    65: op1_12_in20 = reg_0297;
    90: op1_12_in20 = reg_1151;
    48: op1_12_in20 = reg_0475;
    66: op1_12_in20 = reg_0225;
    91: op1_12_in20 = reg_0235;
    67: op1_12_in20 = reg_0086;
    93: op1_12_in20 = reg_0086;
    92: op1_12_in20 = reg_0612;
    124: op1_12_in20 = reg_0612;
    94: op1_12_in20 = reg_1484;
    95: op1_12_in20 = reg_0694;
    96: op1_12_in20 = reg_1420;
    97: op1_12_in20 = reg_0219;
    99: op1_12_in20 = reg_1492;
    100: op1_12_in20 = reg_0299;
    101: op1_12_in20 = reg_0882;
    102: op1_12_in20 = reg_0137;
    103: op1_12_in20 = reg_0798;
    104: op1_12_in20 = reg_0126;
    105: op1_12_in20 = reg_0952;
    106: op1_12_in20 = reg_0720;
    47: op1_12_in20 = reg_0794;
    108: op1_12_in20 = reg_0425;
    125: op1_12_in20 = reg_0425;
    109: op1_12_in20 = reg_0723;
    110: op1_12_in20 = reg_0648;
    111: op1_12_in20 = reg_0711;
    112: op1_12_in20 = reg_0173;
    113: op1_12_in20 = reg_0154;
    115: op1_12_in20 = reg_0128;
    116: op1_12_in20 = imem07_in[3:0];
    117: op1_12_in20 = reg_0381;
    118: op1_12_in20 = reg_0108;
    119: op1_12_in20 = reg_0090;
    120: op1_12_in20 = reg_0730;
    122: op1_12_in20 = reg_0374;
    123: op1_12_in20 = reg_0104;
    44: op1_12_in20 = reg_0604;
    126: op1_12_in20 = reg_0431;
    127: op1_12_in20 = reg_0159;
    128: op1_12_in20 = reg_0994;
    129: op1_12_in20 = reg_0985;
    130: op1_12_in20 = reg_0157;
    default: op1_12_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv20 = 1;
    53: op1_12_inv20 = 1;
    55: op1_12_inv20 = 1;
    86: op1_12_inv20 = 1;
    74: op1_12_inv20 = 1;
    69: op1_12_inv20 = 1;
    49: op1_12_inv20 = 1;
    75: op1_12_inv20 = 1;
    56: op1_12_inv20 = 1;
    50: op1_12_inv20 = 1;
    76: op1_12_inv20 = 1;
    87: op1_12_inv20 = 1;
    57: op1_12_inv20 = 1;
    77: op1_12_inv20 = 1;
    70: op1_12_inv20 = 1;
    59: op1_12_inv20 = 1;
    51: op1_12_inv20 = 1;
    60: op1_12_inv20 = 1;
    88: op1_12_inv20 = 1;
    80: op1_12_inv20 = 1;
    81: op1_12_inv20 = 1;
    82: op1_12_inv20 = 1;
    46: op1_12_inv20 = 1;
    64: op1_12_inv20 = 1;
    89: op1_12_inv20 = 1;
    84: op1_12_inv20 = 1;
    85: op1_12_inv20 = 1;
    65: op1_12_inv20 = 1;
    90: op1_12_inv20 = 1;
    48: op1_12_inv20 = 1;
    67: op1_12_inv20 = 1;
    92: op1_12_inv20 = 1;
    94: op1_12_inv20 = 1;
    95: op1_12_inv20 = 1;
    96: op1_12_inv20 = 1;
    101: op1_12_inv20 = 1;
    106: op1_12_inv20 = 1;
    47: op1_12_inv20 = 1;
    108: op1_12_inv20 = 1;
    109: op1_12_inv20 = 1;
    113: op1_12_inv20 = 1;
    120: op1_12_inv20 = 1;
    125: op1_12_inv20 = 1;
    127: op1_12_inv20 = 1;
    129: op1_12_inv20 = 1;
    130: op1_12_inv20 = 1;
    default: op1_12_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in21 = reg_1315;
    53: op1_12_in21 = reg_0497;
    55: op1_12_in21 = reg_0840;
    73: op1_12_in21 = reg_0589;
    86: op1_12_in21 = imem04_in[15:12];
    70: op1_12_in21 = imem04_in[15:12];
    74: op1_12_in21 = reg_0548;
    69: op1_12_in21 = reg_0830;
    49: op1_12_in21 = reg_0592;
    102: op1_12_in21 = reg_0592;
    54: op1_12_in21 = reg_1163;
    75: op1_12_in21 = reg_0528;
    56: op1_12_in21 = reg_0481;
    50: op1_12_in21 = reg_0030;
    130: op1_12_in21 = reg_0030;
    76: op1_12_in21 = reg_1508;
    68: op1_12_in21 = reg_0454;
    71: op1_12_in21 = reg_0077;
    87: op1_12_in21 = reg_0246;
    57: op1_12_in21 = reg_0667;
    77: op1_12_in21 = reg_0159;
    61: op1_12_in21 = reg_1068;
    58: op1_12_in21 = reg_0280;
    78: op1_12_in21 = reg_0319;
    59: op1_12_in21 = reg_0879;
    79: op1_12_in21 = reg_0775;
    51: op1_12_in21 = reg_0380;
    60: op1_12_in21 = reg_0468;
    88: op1_12_in21 = reg_1199;
    80: op1_12_in21 = reg_0080;
    62: op1_12_in21 = reg_0859;
    81: op1_12_in21 = reg_0891;
    52: op1_12_in21 = reg_0214;
    63: op1_12_in21 = reg_0828;
    82: op1_12_in21 = reg_0492;
    46: op1_12_in21 = reg_0878;
    83: op1_12_in21 = reg_0434;
    64: op1_12_in21 = reg_0550;
    89: op1_12_in21 = reg_0333;
    84: op1_12_in21 = reg_0333;
    85: op1_12_in21 = reg_0348;
    65: op1_12_in21 = reg_1345;
    90: op1_12_in21 = reg_0096;
    48: op1_12_in21 = reg_0990;
    66: op1_12_in21 = reg_0157;
    91: op1_12_in21 = reg_0710;
    67: op1_12_in21 = reg_0518;
    92: op1_12_in21 = reg_0966;
    93: op1_12_in21 = reg_0521;
    94: op1_12_in21 = reg_0393;
    95: op1_12_in21 = reg_1203;
    96: op1_12_in21 = reg_0782;
    120: op1_12_in21 = reg_0782;
    97: op1_12_in21 = reg_1349;
    99: op1_12_in21 = reg_0695;
    111: op1_12_in21 = reg_0695;
    100: op1_12_in21 = reg_1350;
    101: op1_12_in21 = reg_0541;
    103: op1_12_in21 = reg_0967;
    104: op1_12_in21 = reg_0111;
    105: op1_12_in21 = reg_1231;
    106: op1_12_in21 = reg_1505;
    47: op1_12_in21 = reg_0347;
    108: op1_12_in21 = reg_1372;
    109: op1_12_in21 = reg_0277;
    110: op1_12_in21 = reg_0066;
    112: op1_12_in21 = reg_0491;
    113: op1_12_in21 = reg_0706;
    115: op1_12_in21 = reg_0126;
    116: op1_12_in21 = imem07_in[7:4];
    117: op1_12_in21 = reg_0473;
    118: op1_12_in21 = reg_0350;
    119: op1_12_in21 = reg_0873;
    122: op1_12_in21 = reg_0584;
    123: op1_12_in21 = reg_0882;
    124: op1_12_in21 = reg_1474;
    125: op1_12_in21 = reg_1144;
    44: op1_12_in21 = reg_0567;
    126: op1_12_in21 = reg_0435;
    127: op1_12_in21 = reg_0158;
    128: op1_12_in21 = reg_1055;
    129: op1_12_in21 = reg_0576;
    default: op1_12_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv21 = 1;
    69: op1_12_inv21 = 1;
    49: op1_12_inv21 = 1;
    54: op1_12_inv21 = 1;
    56: op1_12_inv21 = 1;
    50: op1_12_inv21 = 1;
    76: op1_12_inv21 = 1;
    68: op1_12_inv21 = 1;
    87: op1_12_inv21 = 1;
    57: op1_12_inv21 = 1;
    79: op1_12_inv21 = 1;
    60: op1_12_inv21 = 1;
    88: op1_12_inv21 = 1;
    80: op1_12_inv21 = 1;
    62: op1_12_inv21 = 1;
    52: op1_12_inv21 = 1;
    63: op1_12_inv21 = 1;
    83: op1_12_inv21 = 1;
    64: op1_12_inv21 = 1;
    89: op1_12_inv21 = 1;
    84: op1_12_inv21 = 1;
    65: op1_12_inv21 = 1;
    48: op1_12_inv21 = 1;
    91: op1_12_inv21 = 1;
    93: op1_12_inv21 = 1;
    96: op1_12_inv21 = 1;
    97: op1_12_inv21 = 1;
    99: op1_12_inv21 = 1;
    102: op1_12_inv21 = 1;
    106: op1_12_inv21 = 1;
    47: op1_12_inv21 = 1;
    110: op1_12_inv21 = 1;
    111: op1_12_inv21 = 1;
    113: op1_12_inv21 = 1;
    118: op1_12_inv21 = 1;
    119: op1_12_inv21 = 1;
    122: op1_12_inv21 = 1;
    124: op1_12_inv21 = 1;
    125: op1_12_inv21 = 1;
    126: op1_12_inv21 = 1;
    129: op1_12_inv21 = 1;
    default: op1_12_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in22 = reg_0187;
    53: op1_12_in22 = reg_0495;
    55: op1_12_in22 = reg_0537;
    73: op1_12_in22 = reg_0038;
    63: op1_12_in22 = reg_0038;
    86: op1_12_in22 = reg_0252;
    74: op1_12_in22 = reg_0742;
    69: op1_12_in22 = reg_0177;
    49: op1_12_in22 = reg_0114;
    54: op1_12_in22 = reg_0395;
    75: op1_12_in22 = reg_1228;
    56: op1_12_in22 = reg_0849;
    50: op1_12_in22 = reg_0285;
    76: op1_12_in22 = reg_0397;
    68: op1_12_in22 = reg_0904;
    90: op1_12_in22 = reg_0904;
    71: op1_12_in22 = reg_0079;
    87: op1_12_in22 = reg_1300;
    57: op1_12_in22 = reg_0668;
    77: op1_12_in22 = reg_0156;
    97: op1_12_in22 = reg_0156;
    61: op1_12_in22 = reg_0611;
    58: op1_12_in22 = reg_0758;
    78: op1_12_in22 = reg_0487;
    70: op1_12_in22 = reg_0320;
    59: op1_12_in22 = reg_0008;
    79: op1_12_in22 = reg_0665;
    51: op1_12_in22 = reg_0903;
    60: op1_12_in22 = reg_0469;
    124: op1_12_in22 = reg_0469;
    88: op1_12_in22 = reg_1208;
    80: op1_12_in22 = reg_0278;
    62: op1_12_in22 = reg_0109;
    81: op1_12_in22 = reg_1003;
    52: op1_12_in22 = reg_0223;
    82: op1_12_in22 = reg_0601;
    46: op1_12_in22 = reg_0009;
    83: op1_12_in22 = reg_1457;
    64: op1_12_in22 = reg_0548;
    89: op1_12_in22 = reg_0346;
    84: op1_12_in22 = reg_0795;
    85: op1_12_in22 = reg_0898;
    65: op1_12_in22 = reg_0924;
    48: op1_12_in22 = reg_0776;
    66: op1_12_in22 = reg_0139;
    91: op1_12_in22 = reg_0185;
    92: op1_12_in22 = reg_0967;
    94: op1_12_in22 = reg_0575;
    95: op1_12_in22 = reg_1200;
    96: op1_12_in22 = reg_1467;
    99: op1_12_in22 = reg_0024;
    100: op1_12_in22 = reg_0029;
    101: op1_12_in22 = reg_0025;
    102: op1_12_in22 = reg_0100;
    103: op1_12_in22 = reg_0147;
    104: op1_12_in22 = reg_0106;
    105: op1_12_in22 = reg_1093;
    106: op1_12_in22 = reg_0716;
    47: op1_12_in22 = reg_0831;
    108: op1_12_in22 = reg_0034;
    109: op1_12_in22 = imem01_in[15:12];
    110: op1_12_in22 = reg_0173;
    111: op1_12_in22 = reg_0294;
    112: op1_12_in22 = reg_0564;
    113: op1_12_in22 = reg_1425;
    115: op1_12_in22 = reg_0684;
    116: op1_12_in22 = imem07_in[15:12];
    117: op1_12_in22 = reg_0068;
    118: op1_12_in22 = reg_0378;
    119: op1_12_in22 = reg_0318;
    120: op1_12_in22 = reg_1437;
    122: op1_12_in22 = reg_0619;
    123: op1_12_in22 = reg_0673;
    125: op1_12_in22 = reg_1338;
    44: op1_12_in22 = reg_0566;
    126: op1_12_in22 = reg_1321;
    127: op1_12_in22 = reg_0775;
    128: op1_12_in22 = reg_0231;
    129: op1_12_in22 = reg_0401;
    130: op1_12_in22 = reg_0286;
    default: op1_12_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv22 = 1;
    74: op1_12_inv22 = 1;
    50: op1_12_inv22 = 1;
    71: op1_12_inv22 = 1;
    87: op1_12_inv22 = 1;
    61: op1_12_inv22 = 1;
    78: op1_12_inv22 = 1;
    70: op1_12_inv22 = 1;
    59: op1_12_inv22 = 1;
    51: op1_12_inv22 = 1;
    60: op1_12_inv22 = 1;
    80: op1_12_inv22 = 1;
    52: op1_12_inv22 = 1;
    63: op1_12_inv22 = 1;
    82: op1_12_inv22 = 1;
    46: op1_12_inv22 = 1;
    89: op1_12_inv22 = 1;
    85: op1_12_inv22 = 1;
    90: op1_12_inv22 = 1;
    92: op1_12_inv22 = 1;
    94: op1_12_inv22 = 1;
    95: op1_12_inv22 = 1;
    97: op1_12_inv22 = 1;
    100: op1_12_inv22 = 1;
    101: op1_12_inv22 = 1;
    102: op1_12_inv22 = 1;
    104: op1_12_inv22 = 1;
    106: op1_12_inv22 = 1;
    47: op1_12_inv22 = 1;
    109: op1_12_inv22 = 1;
    110: op1_12_inv22 = 1;
    112: op1_12_inv22 = 1;
    117: op1_12_inv22 = 1;
    118: op1_12_inv22 = 1;
    119: op1_12_inv22 = 1;
    120: op1_12_inv22 = 1;
    122: op1_12_inv22 = 1;
    125: op1_12_inv22 = 1;
    44: op1_12_inv22 = 1;
    128: op1_12_inv22 = 1;
    129: op1_12_inv22 = 1;
    130: op1_12_inv22 = 1;
    default: op1_12_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in23 = reg_0851;
    53: op1_12_in23 = reg_0496;
    55: op1_12_in23 = reg_0534;
    73: op1_12_in23 = reg_0039;
    86: op1_12_in23 = reg_0574;
    74: op1_12_in23 = reg_1474;
    69: op1_12_in23 = imem03_in[7:4];
    54: op1_12_in23 = reg_0392;
    75: op1_12_in23 = reg_0171;
    56: op1_12_in23 = reg_0823;
    50: op1_12_in23 = reg_0442;
    76: op1_12_in23 = reg_0172;
    68: op1_12_in23 = reg_0340;
    71: op1_12_in23 = reg_0292;
    87: op1_12_in23 = reg_1093;
    57: op1_12_in23 = reg_0225;
    77: op1_12_in23 = reg_0157;
    61: op1_12_in23 = reg_0602;
    82: op1_12_in23 = reg_0602;
    58: op1_12_in23 = reg_0756;
    78: op1_12_in23 = imem04_in[15:12];
    70: op1_12_in23 = reg_0342;
    59: op1_12_in23 = reg_0154;
    79: op1_12_in23 = reg_0661;
    51: op1_12_in23 = reg_0708;
    60: op1_12_in23 = reg_0930;
    88: op1_12_in23 = reg_0291;
    80: op1_12_in23 = reg_0043;
    62: op1_12_in23 = reg_0717;
    81: op1_12_in23 = reg_1184;
    52: op1_12_in23 = reg_0245;
    63: op1_12_in23 = reg_0974;
    46: op1_12_in23 = reg_0008;
    83: op1_12_in23 = reg_1456;
    64: op1_12_in23 = reg_0553;
    89: op1_12_in23 = reg_0733;
    84: op1_12_in23 = reg_0827;
    85: op1_12_in23 = reg_0263;
    65: op1_12_in23 = reg_0224;
    90: op1_12_in23 = reg_0420;
    48: op1_12_in23 = reg_0326;
    66: op1_12_in23 = reg_0031;
    91: op1_12_in23 = reg_0709;
    92: op1_12_in23 = reg_0439;
    94: op1_12_in23 = reg_1348;
    95: op1_12_in23 = reg_1233;
    96: op1_12_in23 = reg_0751;
    97: op1_12_in23 = reg_0158;
    99: op1_12_in23 = reg_0507;
    100: op1_12_in23 = reg_0030;
    101: op1_12_in23 = reg_0411;
    102: op1_12_in23 = reg_0002;
    103: op1_12_in23 = reg_0386;
    104: op1_12_in23 = reg_1433;
    105: op1_12_in23 = reg_1199;
    106: op1_12_in23 = reg_0622;
    47: op1_12_in23 = reg_0702;
    108: op1_12_in23 = reg_0164;
    109: op1_12_in23 = reg_0548;
    110: op1_12_in23 = reg_0302;
    111: op1_12_in23 = reg_1078;
    112: op1_12_in23 = reg_1180;
    113: op1_12_in23 = reg_0600;
    115: op1_12_in23 = reg_0473;
    116: op1_12_in23 = reg_0993;
    117: op1_12_in23 = reg_0217;
    118: op1_12_in23 = reg_0218;
    119: op1_12_in23 = reg_0450;
    120: op1_12_in23 = reg_1467;
    122: op1_12_in23 = reg_0345;
    123: op1_12_in23 = reg_0208;
    124: op1_12_in23 = reg_1457;
    125: op1_12_in23 = reg_0252;
    44: op1_12_in23 = reg_0334;
    126: op1_12_in23 = reg_0026;
    127: op1_12_in23 = reg_0366;
    128: op1_12_in23 = reg_0100;
    129: op1_12_in23 = reg_0013;
    130: op1_12_in23 = reg_0408;
    default: op1_12_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv23 = 1;
    55: op1_12_inv23 = 1;
    54: op1_12_inv23 = 1;
    75: op1_12_inv23 = 1;
    50: op1_12_inv23 = 1;
    68: op1_12_inv23 = 1;
    87: op1_12_inv23 = 1;
    57: op1_12_inv23 = 1;
    77: op1_12_inv23 = 1;
    59: op1_12_inv23 = 1;
    79: op1_12_inv23 = 1;
    51: op1_12_inv23 = 1;
    62: op1_12_inv23 = 1;
    81: op1_12_inv23 = 1;
    82: op1_12_inv23 = 1;
    46: op1_12_inv23 = 1;
    83: op1_12_inv23 = 1;
    64: op1_12_inv23 = 1;
    89: op1_12_inv23 = 1;
    85: op1_12_inv23 = 1;
    48: op1_12_inv23 = 1;
    66: op1_12_inv23 = 1;
    91: op1_12_inv23 = 1;
    92: op1_12_inv23 = 1;
    97: op1_12_inv23 = 1;
    100: op1_12_inv23 = 1;
    101: op1_12_inv23 = 1;
    102: op1_12_inv23 = 1;
    103: op1_12_inv23 = 1;
    104: op1_12_inv23 = 1;
    105: op1_12_inv23 = 1;
    106: op1_12_inv23 = 1;
    109: op1_12_inv23 = 1;
    110: op1_12_inv23 = 1;
    111: op1_12_inv23 = 1;
    112: op1_12_inv23 = 1;
    115: op1_12_inv23 = 1;
    116: op1_12_inv23 = 1;
    119: op1_12_inv23 = 1;
    126: op1_12_inv23 = 1;
    128: op1_12_inv23 = 1;
    129: op1_12_inv23 = 1;
    130: op1_12_inv23 = 1;
    default: op1_12_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in24 = reg_0031;
    53: op1_12_in24 = reg_0475;
    55: op1_12_in24 = reg_0493;
    73: op1_12_in24 = reg_0754;
    86: op1_12_in24 = reg_0414;
    74: op1_12_in24 = reg_0438;
    92: op1_12_in24 = reg_0438;
    69: op1_12_in24 = reg_1033;
    54: op1_12_in24 = reg_0564;
    75: op1_12_in24 = reg_0419;
    56: op1_12_in24 = reg_1143;
    50: op1_12_in24 = reg_0738;
    76: op1_12_in24 = reg_0636;
    68: op1_12_in24 = reg_0237;
    71: op1_12_in24 = reg_0010;
    87: op1_12_in24 = reg_0104;
    105: op1_12_in24 = reg_0104;
    57: op1_12_in24 = reg_0774;
    77: op1_12_in24 = reg_0489;
    97: op1_12_in24 = reg_0489;
    61: op1_12_in24 = reg_0547;
    58: op1_12_in24 = reg_0121;
    78: op1_12_in24 = reg_0117;
    70: op1_12_in24 = reg_0304;
    59: op1_12_in24 = reg_0024;
    79: op1_12_in24 = reg_0663;
    51: op1_12_in24 = reg_0294;
    60: op1_12_in24 = reg_0146;
    88: op1_12_in24 = reg_1384;
    80: op1_12_in24 = reg_0013;
    62: op1_12_in24 = reg_0585;
    81: op1_12_in24 = reg_1516;
    52: op1_12_in24 = reg_0867;
    63: op1_12_in24 = reg_0729;
    82: op1_12_in24 = reg_0631;
    46: op1_12_in24 = reg_0154;
    83: op1_12_in24 = reg_0148;
    64: op1_12_in24 = reg_0982;
    89: op1_12_in24 = reg_1164;
    84: op1_12_in24 = reg_0635;
    85: op1_12_in24 = reg_1372;
    65: op1_12_in24 = reg_0284;
    90: op1_12_in24 = reg_0019;
    48: op1_12_in24 = reg_0935;
    66: op1_12_in24 = reg_0665;
    91: op1_12_in24 = reg_0706;
    94: op1_12_in24 = reg_0602;
    95: op1_12_in24 = reg_0500;
    96: op1_12_in24 = reg_0827;
    99: op1_12_in24 = reg_0235;
    100: op1_12_in24 = reg_0437;
    101: op1_12_in24 = reg_0721;
    102: op1_12_in24 = reg_0087;
    103: op1_12_in24 = reg_0385;
    104: op1_12_in24 = reg_0684;
    106: op1_12_in24 = reg_0624;
    47: op1_12_in24 = reg_0445;
    108: op1_12_in24 = reg_0731;
    109: op1_12_in24 = reg_0239;
    110: op1_12_in24 = reg_0300;
    111: op1_12_in24 = reg_1006;
    112: op1_12_in24 = reg_1402;
    113: op1_12_in24 = reg_0312;
    115: op1_12_in24 = reg_0897;
    116: op1_12_in24 = reg_1315;
    117: op1_12_in24 = reg_0069;
    118: op1_12_in24 = reg_0443;
    119: op1_12_in24 = reg_0888;
    120: op1_12_in24 = reg_0115;
    122: op1_12_in24 = reg_1225;
    123: op1_12_in24 = reg_1216;
    124: op1_12_in24 = reg_1032;
    125: op1_12_in24 = imem04_in[15:12];
    44: op1_12_in24 = reg_0541;
    126: op1_12_in24 = reg_0966;
    127: op1_12_in24 = reg_0618;
    128: op1_12_in24 = reg_0219;
    129: op1_12_in24 = reg_0463;
    130: op1_12_in24 = reg_0137;
    default: op1_12_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv24 = 1;
    86: op1_12_inv24 = 1;
    54: op1_12_inv24 = 1;
    56: op1_12_inv24 = 1;
    71: op1_12_inv24 = 1;
    87: op1_12_inv24 = 1;
    61: op1_12_inv24 = 1;
    58: op1_12_inv24 = 1;
    70: op1_12_inv24 = 1;
    79: op1_12_inv24 = 1;
    51: op1_12_inv24 = 1;
    60: op1_12_inv24 = 1;
    88: op1_12_inv24 = 1;
    81: op1_12_inv24 = 1;
    82: op1_12_inv24 = 1;
    83: op1_12_inv24 = 1;
    64: op1_12_inv24 = 1;
    89: op1_12_inv24 = 1;
    48: op1_12_inv24 = 1;
    94: op1_12_inv24 = 1;
    96: op1_12_inv24 = 1;
    99: op1_12_inv24 = 1;
    101: op1_12_inv24 = 1;
    103: op1_12_inv24 = 1;
    105: op1_12_inv24 = 1;
    47: op1_12_inv24 = 1;
    109: op1_12_inv24 = 1;
    112: op1_12_inv24 = 1;
    113: op1_12_inv24 = 1;
    115: op1_12_inv24 = 1;
    116: op1_12_inv24 = 1;
    117: op1_12_inv24 = 1;
    118: op1_12_inv24 = 1;
    123: op1_12_inv24 = 1;
    125: op1_12_inv24 = 1;
    44: op1_12_inv24 = 1;
    127: op1_12_inv24 = 1;
    129: op1_12_inv24 = 1;
    default: op1_12_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in25 = reg_0465;
    53: op1_12_in25 = reg_0990;
    55: op1_12_in25 = reg_0464;
    73: op1_12_in25 = reg_0377;
    86: op1_12_in25 = reg_0598;
    74: op1_12_in25 = reg_0400;
    69: op1_12_in25 = reg_0638;
    54: op1_12_in25 = reg_0131;
    75: op1_12_in25 = reg_0165;
    56: op1_12_in25 = reg_0252;
    101: op1_12_in25 = reg_0252;
    50: op1_12_in25 = reg_0593;
    76: op1_12_in25 = reg_0194;
    68: op1_12_in25 = reg_0129;
    71: op1_12_in25 = reg_0013;
    87: op1_12_in25 = imem03_in[11:8];
    57: op1_12_in25 = reg_0103;
    77: op1_12_in25 = reg_0031;
    61: op1_12_in25 = reg_0550;
    58: op1_12_in25 = reg_0227;
    78: op1_12_in25 = reg_0095;
    70: op1_12_in25 = reg_0336;
    59: op1_12_in25 = reg_0276;
    79: op1_12_in25 = reg_0442;
    66: op1_12_in25 = reg_0442;
    51: op1_12_in25 = reg_0876;
    60: op1_12_in25 = reg_0403;
    88: op1_12_in25 = reg_1383;
    80: op1_12_in25 = reg_0184;
    62: op1_12_in25 = reg_0373;
    81: op1_12_in25 = reg_1517;
    52: op1_12_in25 = reg_0851;
    128: op1_12_in25 = reg_0851;
    63: op1_12_in25 = reg_0784;
    82: op1_12_in25 = reg_0828;
    46: op1_12_in25 = reg_0830;
    83: op1_12_in25 = reg_0257;
    64: op1_12_in25 = reg_0469;
    89: op1_12_in25 = reg_0996;
    84: op1_12_in25 = reg_0717;
    120: op1_12_in25 = reg_0717;
    85: op1_12_in25 = reg_1368;
    65: op1_12_in25 = reg_0437;
    90: op1_12_in25 = reg_0470;
    48: op1_12_in25 = reg_0127;
    91: op1_12_in25 = reg_0216;
    92: op1_12_in25 = reg_1456;
    94: op1_12_in25 = reg_0344;
    95: op1_12_in25 = reg_1147;
    96: op1_12_in25 = reg_0780;
    97: op1_12_in25 = reg_0030;
    99: op1_12_in25 = reg_0121;
    100: op1_12_in25 = reg_0413;
    103: op1_12_in25 = reg_0363;
    104: op1_12_in25 = reg_0327;
    105: op1_12_in25 = reg_0885;
    106: op1_12_in25 = reg_0979;
    47: op1_12_in25 = imem05_in[7:4];
    108: op1_12_in25 = reg_0694;
    109: op1_12_in25 = reg_0715;
    110: op1_12_in25 = reg_0197;
    119: op1_12_in25 = reg_0197;
    111: op1_12_in25 = reg_0024;
    112: op1_12_in25 = reg_1401;
    113: op1_12_in25 = reg_0962;
    115: op1_12_in25 = reg_0217;
    116: op1_12_in25 = reg_1440;
    117: op1_12_in25 = reg_1515;
    118: op1_12_in25 = reg_1339;
    122: op1_12_in25 = reg_0295;
    123: op1_12_in25 = reg_0493;
    124: op1_12_in25 = imem01_in[3:0];
    125: op1_12_in25 = reg_0535;
    44: op1_12_in25 = reg_0491;
    126: op1_12_in25 = imem01_in[7:4];
    127: op1_12_in25 = reg_0321;
    129: op1_12_in25 = reg_0549;
    130: op1_12_in25 = reg_0085;
    default: op1_12_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_12_inv25 = 1;
    55: op1_12_inv25 = 1;
    54: op1_12_inv25 = 1;
    56: op1_12_inv25 = 1;
    76: op1_12_inv25 = 1;
    68: op1_12_inv25 = 1;
    71: op1_12_inv25 = 1;
    87: op1_12_inv25 = 1;
    57: op1_12_inv25 = 1;
    58: op1_12_inv25 = 1;
    78: op1_12_inv25 = 1;
    59: op1_12_inv25 = 1;
    51: op1_12_inv25 = 1;
    80: op1_12_inv25 = 1;
    62: op1_12_inv25 = 1;
    81: op1_12_inv25 = 1;
    52: op1_12_inv25 = 1;
    63: op1_12_inv25 = 1;
    89: op1_12_inv25 = 1;
    84: op1_12_inv25 = 1;
    85: op1_12_inv25 = 1;
    66: op1_12_inv25 = 1;
    92: op1_12_inv25 = 1;
    95: op1_12_inv25 = 1;
    97: op1_12_inv25 = 1;
    101: op1_12_inv25 = 1;
    103: op1_12_inv25 = 1;
    47: op1_12_inv25 = 1;
    108: op1_12_inv25 = 1;
    109: op1_12_inv25 = 1;
    110: op1_12_inv25 = 1;
    113: op1_12_inv25 = 1;
    115: op1_12_inv25 = 1;
    118: op1_12_inv25 = 1;
    122: op1_12_inv25 = 1;
    125: op1_12_inv25 = 1;
    128: op1_12_inv25 = 1;
    129: op1_12_inv25 = 1;
    130: op1_12_inv25 = 1;
    default: op1_12_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in26 = reg_0284;
    53: op1_12_in26 = reg_0326;
    55: op1_12_in26 = imem04_in[7:4];
    73: op1_12_in26 = reg_1468;
    86: op1_12_in26 = reg_1041;
    74: op1_12_in26 = reg_0901;
    69: op1_12_in26 = reg_0261;
    54: op1_12_in26 = reg_0316;
    75: op1_12_in26 = reg_1179;
    56: op1_12_in26 = reg_0594;
    50: op1_12_in26 = reg_0028;
    127: op1_12_in26 = reg_0028;
    76: op1_12_in26 = reg_0141;
    68: op1_12_in26 = reg_0063;
    71: op1_12_in26 = reg_0446;
    87: op1_12_in26 = reg_0025;
    57: op1_12_in26 = reg_0321;
    77: op1_12_in26 = reg_0465;
    61: op1_12_in26 = reg_0259;
    58: op1_12_in26 = reg_0288;
    78: op1_12_in26 = reg_1488;
    70: op1_12_in26 = reg_0095;
    59: op1_12_in26 = reg_0280;
    79: op1_12_in26 = reg_0591;
    51: op1_12_in26 = reg_0879;
    60: op1_12_in26 = reg_0386;
    88: op1_12_in26 = reg_1372;
    80: op1_12_in26 = reg_1018;
    62: op1_12_in26 = reg_0528;
    81: op1_12_in26 = reg_0954;
    52: op1_12_in26 = reg_0921;
    63: op1_12_in26 = reg_0782;
    82: op1_12_in26 = reg_0038;
    46: op1_12_in26 = reg_0325;
    83: op1_12_in26 = reg_0727;
    64: op1_12_in26 = reg_0819;
    89: op1_12_in26 = reg_0649;
    84: op1_12_in26 = reg_1302;
    85: op1_12_in26 = reg_1339;
    65: op1_12_in26 = reg_0738;
    90: op1_12_in26 = reg_0736;
    48: op1_12_in26 = reg_0125;
    66: op1_12_in26 = reg_0621;
    91: op1_12_in26 = reg_0198;
    92: op1_12_in26 = reg_0149;
    94: op1_12_in26 = reg_0206;
    95: op1_12_in26 = reg_0421;
    96: op1_12_in26 = reg_1035;
    97: op1_12_in26 = reg_0665;
    99: op1_12_in26 = reg_0710;
    100: op1_12_in26 = reg_0620;
    101: op1_12_in26 = imem04_in[3:0];
    103: op1_12_in26 = reg_0595;
    104: op1_12_in26 = reg_0848;
    105: op1_12_in26 = reg_0427;
    106: op1_12_in26 = reg_1225;
    47: op1_12_in26 = reg_0567;
    108: op1_12_in26 = reg_0978;
    109: op1_12_in26 = reg_0968;
    110: op1_12_in26 = reg_0196;
    111: op1_12_in26 = reg_0009;
    112: op1_12_in26 = reg_0794;
    113: op1_12_in26 = reg_0048;
    115: op1_12_in26 = imem03_in[11:8];
    116: op1_12_in26 = reg_1345;
    117: op1_12_in26 = imem03_in[7:4];
    118: op1_12_in26 = reg_0699;
    119: op1_12_in26 = reg_0492;
    120: op1_12_in26 = reg_0714;
    122: op1_12_in26 = reg_0289;
    123: op1_12_in26 = imem04_in[15:12];
    124: op1_12_in26 = reg_0362;
    125: op1_12_in26 = reg_1083;
    44: op1_12_in26 = imem05_in[3:0];
    126: op1_12_in26 = imem01_in[15:12];
    128: op1_12_in26 = reg_1350;
    129: op1_12_in26 = reg_0550;
    default: op1_12_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv26 = 1;
    53: op1_12_inv26 = 1;
    73: op1_12_inv26 = 1;
    86: op1_12_inv26 = 1;
    69: op1_12_inv26 = 1;
    75: op1_12_inv26 = 1;
    50: op1_12_inv26 = 1;
    61: op1_12_inv26 = 1;
    70: op1_12_inv26 = 1;
    79: op1_12_inv26 = 1;
    60: op1_12_inv26 = 1;
    88: op1_12_inv26 = 1;
    82: op1_12_inv26 = 1;
    46: op1_12_inv26 = 1;
    83: op1_12_inv26 = 1;
    90: op1_12_inv26 = 1;
    48: op1_12_inv26 = 1;
    66: op1_12_inv26 = 1;
    91: op1_12_inv26 = 1;
    95: op1_12_inv26 = 1;
    100: op1_12_inv26 = 1;
    103: op1_12_inv26 = 1;
    104: op1_12_inv26 = 1;
    106: op1_12_inv26 = 1;
    111: op1_12_inv26 = 1;
    112: op1_12_inv26 = 1;
    113: op1_12_inv26 = 1;
    115: op1_12_inv26 = 1;
    118: op1_12_inv26 = 1;
    120: op1_12_inv26 = 1;
    122: op1_12_inv26 = 1;
    123: op1_12_inv26 = 1;
    44: op1_12_inv26 = 1;
    126: op1_12_inv26 = 1;
    127: op1_12_inv26 = 1;
    128: op1_12_inv26 = 1;
    default: op1_12_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in27 = reg_0740;
    53: op1_12_in27 = reg_0973;
    55: op1_12_in27 = reg_1082;
    73: op1_12_in27 = reg_0192;
    86: op1_12_in27 = reg_0537;
    74: op1_12_in27 = reg_0724;
    69: op1_12_in27 = reg_1314;
    54: op1_12_in27 = reg_0315;
    75: op1_12_in27 = reg_0152;
    56: op1_12_in27 = imem04_in[3:0];
    50: op1_12_in27 = reg_0085;
    76: op1_12_in27 = reg_0584;
    68: op1_12_in27 = reg_0061;
    71: op1_12_in27 = reg_0486;
    87: op1_12_in27 = reg_0032;
    57: op1_12_in27 = reg_0361;
    127: op1_12_in27 = reg_0361;
    77: op1_12_in27 = reg_0664;
    61: op1_12_in27 = reg_0743;
    58: op1_12_in27 = reg_0232;
    78: op1_12_in27 = reg_0470;
    70: op1_12_in27 = reg_0150;
    59: op1_12_in27 = reg_0218;
    79: op1_12_in27 = reg_0592;
    51: op1_12_in27 = reg_0839;
    60: op1_12_in27 = reg_0868;
    109: op1_12_in27 = reg_0868;
    88: op1_12_in27 = reg_0181;
    80: op1_12_in27 = reg_0138;
    62: op1_12_in27 = reg_0569;
    81: op1_12_in27 = reg_1301;
    52: op1_12_in27 = reg_0031;
    63: op1_12_in27 = reg_0906;
    94: op1_12_in27 = reg_0906;
    82: op1_12_in27 = reg_0039;
    46: op1_12_in27 = reg_0280;
    83: op1_12_in27 = reg_0874;
    64: op1_12_in27 = reg_0726;
    89: op1_12_in27 = reg_1104;
    84: op1_12_in27 = reg_0141;
    85: op1_12_in27 = reg_1257;
    65: op1_12_in27 = reg_0114;
    90: op1_12_in27 = reg_0205;
    48: op1_12_in27 = reg_0379;
    66: op1_12_in27 = reg_0620;
    91: op1_12_in27 = reg_0847;
    92: op1_12_in27 = reg_0383;
    95: op1_12_in27 = reg_0412;
    96: op1_12_in27 = reg_0110;
    97: op1_12_in27 = reg_0663;
    99: op1_12_in27 = reg_1448;
    100: op1_12_in27 = reg_0228;
    101: op1_12_in27 = imem04_in[11:8];
    118: op1_12_in27 = imem04_in[11:8];
    103: op1_12_in27 = reg_0079;
    104: op1_12_in27 = reg_0227;
    105: op1_12_in27 = reg_0443;
    106: op1_12_in27 = reg_0119;
    47: op1_12_in27 = reg_0333;
    108: op1_12_in27 = reg_0531;
    110: op1_12_in27 = reg_1348;
    111: op1_12_in27 = reg_0235;
    112: op1_12_in27 = reg_1373;
    113: op1_12_in27 = reg_0880;
    115: op1_12_in27 = imem03_in[15:12];
    116: op1_12_in27 = reg_0224;
    117: op1_12_in27 = reg_0479;
    119: op1_12_in27 = reg_0196;
    120: op1_12_in27 = reg_0373;
    122: op1_12_in27 = reg_0165;
    123: op1_12_in27 = reg_0462;
    124: op1_12_in27 = reg_0899;
    125: op1_12_in27 = reg_1198;
    44: op1_12_in27 = imem05_in[7:4];
    126: op1_12_in27 = reg_0463;
    128: op1_12_in27 = reg_0157;
    129: op1_12_in27 = reg_0612;
    default: op1_12_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_12_inv27 = 1;
    86: op1_12_inv27 = 1;
    74: op1_12_inv27 = 1;
    54: op1_12_inv27 = 1;
    75: op1_12_inv27 = 1;
    50: op1_12_inv27 = 1;
    68: op1_12_inv27 = 1;
    57: op1_12_inv27 = 1;
    77: op1_12_inv27 = 1;
    70: op1_12_inv27 = 1;
    80: op1_12_inv27 = 1;
    82: op1_12_inv27 = 1;
    46: op1_12_inv27 = 1;
    89: op1_12_inv27 = 1;
    84: op1_12_inv27 = 1;
    85: op1_12_inv27 = 1;
    48: op1_12_inv27 = 1;
    66: op1_12_inv27 = 1;
    91: op1_12_inv27 = 1;
    92: op1_12_inv27 = 1;
    96: op1_12_inv27 = 1;
    101: op1_12_inv27 = 1;
    103: op1_12_inv27 = 1;
    105: op1_12_inv27 = 1;
    47: op1_12_inv27 = 1;
    109: op1_12_inv27 = 1;
    110: op1_12_inv27 = 1;
    113: op1_12_inv27 = 1;
    115: op1_12_inv27 = 1;
    119: op1_12_inv27 = 1;
    125: op1_12_inv27 = 1;
    127: op1_12_inv27 = 1;
    129: op1_12_inv27 = 1;
    default: op1_12_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in28 = reg_0085;
    53: op1_12_in28 = reg_0106;
    55: op1_12_in28 = reg_0676;
    73: op1_12_in28 = reg_0906;
    86: op1_12_in28 = reg_0199;
    74: op1_12_in28 = reg_0895;
    69: op1_12_in28 = reg_1313;
    54: op1_12_in28 = reg_0539;
    75: op1_12_in28 = reg_0022;
    56: op1_12_in28 = reg_1203;
    76: op1_12_in28 = reg_0323;
    68: op1_12_in28 = reg_0021;
    71: op1_12_in28 = reg_0605;
    87: op1_12_in28 = reg_0535;
    57: op1_12_in28 = reg_0228;
    77: op1_12_in28 = reg_0284;
    61: op1_12_in28 = reg_0468;
    58: op1_12_in28 = imem03_in[3:0];
    78: op1_12_in28 = reg_0370;
    70: op1_12_in28 = reg_0209;
    59: op1_12_in28 = reg_0556;
    79: op1_12_in28 = reg_0321;
    51: op1_12_in28 = reg_0279;
    60: op1_12_in28 = reg_0077;
    88: op1_12_in28 = reg_1368;
    80: op1_12_in28 = reg_0056;
    62: op1_12_in28 = reg_0570;
    81: op1_12_in28 = reg_0178;
    52: op1_12_in28 = reg_0442;
    63: op1_12_in28 = reg_0730;
    82: op1_12_in28 = reg_0014;
    46: op1_12_in28 = reg_0312;
    83: op1_12_in28 = reg_0282;
    64: op1_12_in28 = reg_0148;
    89: op1_12_in28 = reg_1404;
    84: op1_12_in28 = reg_0619;
    85: op1_12_in28 = reg_1198;
    65: op1_12_in28 = reg_0051;
    90: op1_12_in28 = reg_0578;
    48: op1_12_in28 = reg_0007;
    66: op1_12_in28 = reg_0102;
    91: op1_12_in28 = reg_0180;
    92: op1_12_in28 = reg_0360;
    94: op1_12_in28 = reg_0377;
    95: op1_12_in28 = reg_0537;
    96: op1_12_in28 = reg_0716;
    97: op1_12_in28 = reg_0286;
    99: op1_12_in28 = reg_1425;
    100: op1_12_in28 = reg_0003;
    101: op1_12_in28 = reg_0467;
    103: op1_12_in28 = reg_0403;
    104: op1_12_in28 = reg_0759;
    111: op1_12_in28 = reg_0759;
    105: op1_12_in28 = imem04_in[3:0];
    106: op1_12_in28 = reg_0165;
    47: op1_12_in28 = reg_0940;
    108: op1_12_in28 = reg_0681;
    109: op1_12_in28 = reg_0384;
    110: op1_12_in28 = reg_1346;
    112: op1_12_in28 = reg_0603;
    113: op1_12_in28 = reg_0378;
    115: op1_12_in28 = reg_0750;
    116: op1_12_in28 = reg_0774;
    117: op1_12_in28 = reg_0049;
    118: op1_12_in28 = reg_0129;
    119: op1_12_in28 = reg_0243;
    120: op1_12_in28 = reg_0586;
    122: op1_12_in28 = reg_0583;
    123: op1_12_in28 = reg_0531;
    124: op1_12_in28 = reg_0080;
    125: op1_12_in28 = reg_1200;
    44: op1_12_in28 = reg_0888;
    126: op1_12_in28 = reg_1473;
    127: op1_12_in28 = reg_1182;
    128: op1_12_in28 = reg_0924;
    129: op1_12_in28 = reg_0715;
    default: op1_12_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_12_inv28 = 1;
    73: op1_12_inv28 = 1;
    74: op1_12_inv28 = 1;
    75: op1_12_inv28 = 1;
    56: op1_12_inv28 = 1;
    68: op1_12_inv28 = 1;
    61: op1_12_inv28 = 1;
    78: op1_12_inv28 = 1;
    59: op1_12_inv28 = 1;
    79: op1_12_inv28 = 1;
    51: op1_12_inv28 = 1;
    52: op1_12_inv28 = 1;
    63: op1_12_inv28 = 1;
    82: op1_12_inv28 = 1;
    83: op1_12_inv28 = 1;
    64: op1_12_inv28 = 1;
    89: op1_12_inv28 = 1;
    48: op1_12_inv28 = 1;
    66: op1_12_inv28 = 1;
    91: op1_12_inv28 = 1;
    92: op1_12_inv28 = 1;
    94: op1_12_inv28 = 1;
    96: op1_12_inv28 = 1;
    99: op1_12_inv28 = 1;
    101: op1_12_inv28 = 1;
    103: op1_12_inv28 = 1;
    47: op1_12_inv28 = 1;
    111: op1_12_inv28 = 1;
    112: op1_12_inv28 = 1;
    115: op1_12_inv28 = 1;
    123: op1_12_inv28 = 1;
    126: op1_12_inv28 = 1;
    127: op1_12_inv28 = 1;
    128: op1_12_inv28 = 1;
    default: op1_12_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_12_in29 = reg_0519;
    53: op1_12_in29 = reg_0105;
    55: op1_12_in29 = reg_0552;
    73: op1_12_in29 = reg_1326;
    86: op1_12_in29 = reg_0451;
    74: op1_12_in29 = reg_0896;
    69: op1_12_in29 = reg_0220;
    54: op1_12_in29 = reg_0939;
    47: op1_12_in29 = reg_0939;
    75: op1_12_in29 = reg_0868;
    56: op1_12_in29 = reg_1065;
    76: op1_12_in29 = reg_0289;
    68: op1_12_in29 = reg_0034;
    71: op1_12_in29 = reg_0590;
    87: op1_12_in29 = reg_1338;
    57: op1_12_in29 = reg_0003;
    77: op1_12_in29 = reg_0404;
    61: op1_12_in29 = reg_0968;
    58: op1_12_in29 = reg_1000;
    78: op1_12_in29 = reg_0675;
    70: op1_12_in29 = reg_0064;
    59: op1_12_in29 = reg_1149;
    79: op1_12_in29 = reg_0050;
    51: op1_12_in29 = reg_0314;
    91: op1_12_in29 = reg_0314;
    60: op1_12_in29 = reg_0290;
    88: op1_12_in29 = reg_0535;
    80: op1_12_in29 = reg_0532;
    62: op1_12_in29 = reg_0171;
    81: op1_12_in29 = reg_0104;
    52: op1_12_in29 = reg_0437;
    63: op1_12_in29 = reg_0696;
    82: op1_12_in29 = reg_0984;
    46: op1_12_in29 = reg_0757;
    83: op1_12_in29 = reg_0283;
    64: op1_12_in29 = reg_0092;
    89: op1_12_in29 = reg_0794;
    84: op1_12_in29 = reg_0617;
    85: op1_12_in29 = reg_0796;
    65: op1_12_in29 = reg_0002;
    90: op1_12_in29 = reg_0315;
    48: op1_12_in29 = reg_0006;
    66: op1_12_in29 = reg_0051;
    92: op1_12_in29 = reg_0595;
    94: op1_12_in29 = reg_1467;
    95: op1_12_in29 = reg_0097;
    96: op1_12_in29 = reg_0194;
    97: op1_12_in29 = reg_0740;
    99: op1_12_in29 = reg_0823;
    100: op1_12_in29 = reg_0085;
    101: op1_12_in29 = reg_0088;
    103: op1_12_in29 = reg_0634;
    104: op1_12_in29 = reg_0377;
    105: op1_12_in29 = reg_0694;
    106: op1_12_in29 = reg_0067;
    108: op1_12_in29 = reg_0407;
    109: op1_12_in29 = reg_0464;
    110: op1_12_in29 = reg_0603;
    111: op1_12_in29 = reg_0246;
    112: op1_12_in29 = reg_0263;
    113: op1_12_in29 = reg_0025;
    115: op1_12_in29 = reg_0759;
    116: op1_12_in29 = reg_0030;
    117: op1_12_in29 = reg_0573;
    118: op1_12_in29 = reg_0797;
    119: op1_12_in29 = reg_0602;
    120: op1_12_in29 = reg_0584;
    122: op1_12_in29 = reg_0754;
    123: op1_12_in29 = reg_0681;
    124: op1_12_in29 = reg_0043;
    125: op1_12_in29 = reg_0488;
    44: op1_12_in29 = reg_0303;
    126: op1_12_in29 = reg_0430;
    128: op1_12_in29 = reg_0665;
    129: op1_12_in29 = reg_0572;
    default: op1_12_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_12_inv29 = 1;
    55: op1_12_inv29 = 1;
    86: op1_12_inv29 = 1;
    74: op1_12_inv29 = 1;
    69: op1_12_inv29 = 1;
    75: op1_12_inv29 = 1;
    56: op1_12_inv29 = 1;
    76: op1_12_inv29 = 1;
    68: op1_12_inv29 = 1;
    87: op1_12_inv29 = 1;
    57: op1_12_inv29 = 1;
    77: op1_12_inv29 = 1;
    61: op1_12_inv29 = 1;
    58: op1_12_inv29 = 1;
    70: op1_12_inv29 = 1;
    51: op1_12_inv29 = 1;
    60: op1_12_inv29 = 1;
    62: op1_12_inv29 = 1;
    63: op1_12_inv29 = 1;
    82: op1_12_inv29 = 1;
    83: op1_12_inv29 = 1;
    64: op1_12_inv29 = 1;
    84: op1_12_inv29 = 1;
    66: op1_12_inv29 = 1;
    91: op1_12_inv29 = 1;
    92: op1_12_inv29 = 1;
    95: op1_12_inv29 = 1;
    96: op1_12_inv29 = 1;
    97: op1_12_inv29 = 1;
    99: op1_12_inv29 = 1;
    100: op1_12_inv29 = 1;
    105: op1_12_inv29 = 1;
    106: op1_12_inv29 = 1;
    109: op1_12_inv29 = 1;
    111: op1_12_inv29 = 1;
    112: op1_12_inv29 = 1;
    113: op1_12_inv29 = 1;
    116: op1_12_inv29 = 1;
    117: op1_12_inv29 = 1;
    118: op1_12_inv29 = 1;
    120: op1_12_inv29 = 1;
    122: op1_12_inv29 = 1;
    123: op1_12_inv29 = 1;
    124: op1_12_inv29 = 1;
    44: op1_12_inv29 = 1;
    126: op1_12_inv29 = 1;
    128: op1_12_inv29 = 1;
    129: op1_12_inv29 = 1;
    default: op1_12_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の30番目の入力
  always @ ( * ) begin
    case ( state )
    53: op1_12_in30 = reg_0307;
    55: op1_12_in30 = reg_0932;
    73: op1_12_in30 = reg_1334;
    86: op1_12_in30 = reg_0698;
    123: op1_12_in30 = reg_0698;
    74: op1_12_in30 = reg_0290;
    69: op1_12_in30 = reg_1300;
    54: op1_12_in30 = reg_0890;
    75: op1_12_in30 = reg_0997;
    56: op1_12_in30 = reg_0633;
    76: op1_12_in30 = reg_1179;
    68: op1_12_in30 = reg_0793;
    71: op1_12_in30 = reg_1260;
    87: op1_12_in30 = reg_1215;
    57: op1_12_in30 = reg_0053;
    65: op1_12_in30 = reg_0053;
    77: op1_12_in30 = reg_0415;
    61: op1_12_in30 = reg_0439;
    58: op1_12_in30 = reg_0965;
    78: op1_12_in30 = reg_0273;
    70: op1_12_in30 = reg_0799;
    59: op1_12_in30 = reg_0559;
    79: op1_12_in30 = reg_0023;
    51: op1_12_in30 = reg_0757;
    60: op1_12_in30 = reg_0277;
    88: op1_12_in30 = reg_0034;
    101: op1_12_in30 = reg_0034;
    80: op1_12_in30 = reg_0666;
    62: op1_12_in30 = reg_0371;
    81: op1_12_in30 = reg_0506;
    52: op1_12_in30 = reg_0621;
    63: op1_12_in30 = reg_0120;
    82: op1_12_in30 = reg_0466;
    90: op1_12_in30 = reg_0466;
    46: op1_12_in30 = reg_0707;
    83: op1_12_in30 = reg_0043;
    64: op1_12_in30 = reg_0874;
    89: op1_12_in30 = reg_0450;
    84: op1_12_in30 = reg_0345;
    85: op1_12_in30 = reg_0412;
    48: op1_12_in30 = reg_0327;
    91: op1_12_in30 = reg_0349;
    92: op1_12_in30 = reg_0335;
    94: op1_12_in30 = reg_0860;
    95: op1_12_in30 = reg_0061;
    96: op1_12_in30 = reg_0624;
    97: op1_12_in30 = reg_0228;
    99: op1_12_in30 = reg_0311;
    100: op1_12_in30 = reg_0123;
    103: op1_12_in30 = reg_0044;
    104: op1_12_in30 = reg_0525;
    105: op1_12_in30 = reg_0552;
    106: op1_12_in30 = reg_0015;
    47: op1_12_in30 = reg_0888;
    108: op1_12_in30 = reg_0598;
    109: op1_12_in30 = reg_0077;
    110: op1_12_in30 = reg_0828;
    111: op1_12_in30 = reg_0233;
    112: op1_12_in30 = reg_0193;
    113: op1_12_in30 = reg_0291;
    115: op1_12_in30 = reg_0246;
    116: op1_12_in30 = reg_0437;
    117: op1_12_in30 = reg_0597;
    118: op1_12_in30 = reg_0462;
    119: op1_12_in30 = reg_1346;
    120: op1_12_in30 = reg_0570;
    122: op1_12_in30 = reg_0195;
    124: op1_12_in30 = reg_0011;
    125: op1_12_in30 = reg_0537;
    44: op1_12_in30 = reg_0272;
    126: op1_12_in30 = reg_0899;
    128: op1_12_in30 = reg_0663;
    129: op1_12_in30 = reg_0819;
    default: op1_12_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_12_inv30 = 1;
    74: op1_12_inv30 = 1;
    69: op1_12_inv30 = 1;
    54: op1_12_inv30 = 1;
    76: op1_12_inv30 = 1;
    71: op1_12_inv30 = 1;
    58: op1_12_inv30 = 1;
    78: op1_12_inv30 = 1;
    59: op1_12_inv30 = 1;
    79: op1_12_inv30 = 1;
    51: op1_12_inv30 = 1;
    60: op1_12_inv30 = 1;
    88: op1_12_inv30 = 1;
    62: op1_12_inv30 = 1;
    82: op1_12_inv30 = 1;
    64: op1_12_inv30 = 1;
    65: op1_12_inv30 = 1;
    90: op1_12_inv30 = 1;
    92: op1_12_inv30 = 1;
    101: op1_12_inv30 = 1;
    110: op1_12_inv30 = 1;
    111: op1_12_inv30 = 1;
    119: op1_12_inv30 = 1;
    122: op1_12_inv30 = 1;
    129: op1_12_inv30 = 1;
    default: op1_12_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_12_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#12の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_12_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in00 = reg_0445;
    98: op1_13_in00 = reg_0445;
    53: op1_13_in00 = reg_0292;
    73: op1_13_in00 = reg_0720;
    86: op1_13_in00 = reg_0480;
    81: op1_13_in00 = reg_0480;
    55: op1_13_in00 = reg_0191;
    74: op1_13_in00 = imem04_in[11:8];
    69: op1_13_in00 = reg_0612;
    54: op1_13_in00 = reg_0902;
    49: op1_13_in00 = reg_0244;
    75: op1_13_in00 = reg_1078;
    56: op1_13_in00 = reg_0727;
    65: op1_13_in00 = reg_0727;
    50: op1_13_in00 = imem06_in[15:12];
    76: op1_13_in00 = reg_0575;
    71: op1_13_in00 = imem00_in[7:4];
    87: op1_13_in00 = reg_0255;
    68: op1_13_in00 = reg_0261;
    57: op1_13_in00 = reg_1182;
    77: op1_13_in00 = reg_0899;
    61: op1_13_in00 = reg_0580;
    58: op1_13_in00 = reg_0828;
    78: op1_13_in00 = reg_0219;
    79: op1_13_in00 = reg_0219;
    70: op1_13_in00 = reg_0281;
    59: op1_13_in00 = reg_0199;
    51: op1_13_in00 = reg_0264;
    60: op1_13_in00 = reg_1257;
    88: op1_13_in00 = reg_0326;
    80: op1_13_in00 = reg_0412;
    62: op1_13_in00 = reg_0018;
    63: op1_13_in00 = reg_0383;
    52: op1_13_in00 = reg_0925;
    82: op1_13_in00 = reg_0791;
    83: op1_13_in00 = reg_0449;
    119: op1_13_in00 = reg_0449;
    64: op1_13_in00 = reg_0077;
    89: op1_13_in00 = reg_0558;
    84: op1_13_in00 = reg_0983;
    46: op1_13_in00 = reg_0173;
    85: op1_13_in00 = reg_1041;
    90: op1_13_in00 = reg_1168;
    66: op1_13_in00 = reg_0047;
    48: op1_13_in00 = reg_0782;
    125: op1_13_in00 = reg_0782;
    91: op1_13_in00 = reg_1313;
    67: op1_13_in00 = reg_0161;
    92: op1_13_in00 = reg_0311;
    93: op1_13_in00 = reg_1207;
    33: op1_13_in00 = imem07_in[15:12];
    94: op1_13_in00 = reg_0869;
    95: op1_13_in00 = reg_0582;
    96: op1_13_in00 = reg_0569;
    28: op1_13_in00 = reg_0229;
    97: op1_13_in00 = reg_1244;
    99: op1_13_in00 = reg_0145;
    100: op1_13_in00 = reg_0638;
    101: op1_13_in00 = reg_0462;
    102: op1_13_in00 = reg_0248;
    116: op1_13_in00 = reg_0248;
    103: op1_13_in00 = reg_0011;
    104: op1_13_in00 = reg_0328;
    37: op1_13_in00 = reg_0441;
    105: op1_13_in00 = reg_0488;
    106: op1_13_in00 = imem07_in[11:8];
    107: op1_13_in00 = imem00_in[11:8];
    108: op1_13_in00 = reg_0537;
    109: op1_13_in00 = reg_0724;
    110: op1_13_in00 = reg_0039;
    111: op1_13_in00 = reg_0185;
    112: op1_13_in00 = reg_1058;
    113: op1_13_in00 = reg_0313;
    114: op1_13_in00 = reg_0958;
    115: op1_13_in00 = reg_1145;
    117: op1_13_in00 = reg_0180;
    47: op1_13_in00 = reg_0182;
    118: op1_13_in00 = reg_1233;
    120: op1_13_in00 = reg_0345;
    121: op1_13_in00 = reg_1080;
    122: op1_13_in00 = reg_0215;
    123: op1_13_in00 = reg_0835;
    124: op1_13_in00 = reg_0721;
    126: op1_13_in00 = reg_0162;
    44: op1_13_in00 = reg_0467;
    127: op1_13_in00 = reg_1469;
    128: op1_13_in00 = reg_1242;
    129: op1_13_in00 = reg_0430;
    130: op1_13_in00 = reg_0171;
    default: op1_13_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_13_inv00 = 1;
    55: op1_13_inv00 = 1;
    74: op1_13_inv00 = 1;
    54: op1_13_inv00 = 1;
    49: op1_13_inv00 = 1;
    56: op1_13_inv00 = 1;
    50: op1_13_inv00 = 1;
    71: op1_13_inv00 = 1;
    57: op1_13_inv00 = 1;
    78: op1_13_inv00 = 1;
    70: op1_13_inv00 = 1;
    60: op1_13_inv00 = 1;
    80: op1_13_inv00 = 1;
    81: op1_13_inv00 = 1;
    52: op1_13_inv00 = 1;
    82: op1_13_inv00 = 1;
    64: op1_13_inv00 = 1;
    89: op1_13_inv00 = 1;
    84: op1_13_inv00 = 1;
    46: op1_13_inv00 = 1;
    65: op1_13_inv00 = 1;
    66: op1_13_inv00 = 1;
    48: op1_13_inv00 = 1;
    91: op1_13_inv00 = 1;
    92: op1_13_inv00 = 1;
    93: op1_13_inv00 = 1;
    95: op1_13_inv00 = 1;
    28: op1_13_inv00 = 1;
    97: op1_13_inv00 = 1;
    99: op1_13_inv00 = 1;
    101: op1_13_inv00 = 1;
    104: op1_13_inv00 = 1;
    37: op1_13_inv00 = 1;
    107: op1_13_inv00 = 1;
    110: op1_13_inv00 = 1;
    113: op1_13_inv00 = 1;
    116: op1_13_inv00 = 1;
    117: op1_13_inv00 = 1;
    118: op1_13_inv00 = 1;
    122: op1_13_inv00 = 1;
    123: op1_13_inv00 = 1;
    124: op1_13_inv00 = 1;
    127: op1_13_inv00 = 1;
    130: op1_13_inv00 = 1;
    default: op1_13_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in01 = reg_0844;
    53: op1_13_in01 = reg_0278;
    73: op1_13_in01 = reg_0863;
    86: op1_13_in01 = reg_1325;
    55: op1_13_in01 = reg_0490;
    74: op1_13_in01 = reg_0675;
    69: op1_13_in01 = reg_0456;
    54: op1_13_in01 = reg_0077;
    49: op1_13_in01 = reg_0018;
    75: op1_13_in01 = reg_1242;
    56: op1_13_in01 = reg_0147;
    65: op1_13_in01 = reg_0147;
    50: op1_13_in01 = reg_0907;
    76: op1_13_in01 = reg_1346;
    71: op1_13_in01 = imem00_in[11:8];
    87: op1_13_in01 = reg_1132;
    68: op1_13_in01 = reg_0559;
    77: op1_13_in01 = reg_0901;
    61: op1_13_in01 = reg_0866;
    58: op1_13_in01 = reg_1164;
    90: op1_13_in01 = reg_1164;
    78: op1_13_in01 = reg_0445;
    70: op1_13_in01 = reg_0758;
    59: op1_13_in01 = reg_0305;
    79: op1_13_in01 = imem00_in[15:12];
    51: op1_13_in01 = reg_0619;
    60: op1_13_in01 = reg_1200;
    88: op1_13_in01 = reg_0168;
    80: op1_13_in01 = reg_0406;
    44: op1_13_in01 = reg_0406;
    62: op1_13_in01 = reg_0017;
    81: op1_13_in01 = reg_0573;
    63: op1_13_in01 = reg_0360;
    52: op1_13_in01 = reg_0193;
    82: op1_13_in01 = reg_0983;
    83: op1_13_in01 = reg_0984;
    125: op1_13_in01 = reg_0984;
    64: op1_13_in01 = reg_0043;
    89: op1_13_in01 = reg_1208;
    84: op1_13_in01 = reg_0640;
    46: op1_13_in01 = reg_0176;
    85: op1_13_in01 = reg_1077;
    66: op1_13_in01 = reg_0093;
    48: op1_13_in01 = reg_0784;
    91: op1_13_in01 = reg_0597;
    67: op1_13_in01 = reg_1151;
    92: op1_13_in01 = reg_0312;
    93: op1_13_in01 = reg_1455;
    33: op1_13_in01 = reg_0591;
    94: op1_13_in01 = reg_1501;
    95: op1_13_in01 = reg_0487;
    96: op1_13_in01 = reg_0296;
    28: op1_13_in01 = reg_0086;
    97: op1_13_in01 = reg_0672;
    98: op1_13_in01 = reg_1281;
    114: op1_13_in01 = reg_1281;
    99: op1_13_in01 = reg_0180;
    100: op1_13_in01 = reg_0725;
    107: op1_13_in01 = reg_0725;
    127: op1_13_in01 = reg_0725;
    101: op1_13_in01 = reg_1214;
    102: op1_13_in01 = reg_0669;
    103: op1_13_in01 = reg_0010;
    104: op1_13_in01 = reg_0049;
    37: op1_13_in01 = reg_0437;
    105: op1_13_in01 = reg_0500;
    118: op1_13_in01 = reg_0500;
    106: op1_13_in01 = reg_1096;
    108: op1_13_in01 = reg_1004;
    109: op1_13_in01 = reg_0403;
    110: op1_13_in01 = imem06_in[11:8];
    111: op1_13_in01 = reg_0847;
    112: op1_13_in01 = reg_0397;
    113: op1_13_in01 = reg_1139;
    115: op1_13_in01 = reg_0706;
    116: op1_13_in01 = reg_1278;
    117: op1_13_in01 = reg_0375;
    47: op1_13_in01 = reg_0045;
    119: op1_13_in01 = reg_0861;
    120: op1_13_in01 = reg_0979;
    121: op1_13_in01 = reg_0319;
    122: op1_13_in01 = reg_0213;
    123: op1_13_in01 = reg_1189;
    124: op1_13_in01 = reg_0659;
    126: op1_13_in01 = reg_1068;
    128: op1_13_in01 = reg_1099;
    129: op1_13_in01 = reg_0434;
    130: op1_13_in01 = reg_1079;
    default: op1_13_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv01 = 1;
    53: op1_13_inv01 = 1;
    55: op1_13_inv01 = 1;
    74: op1_13_inv01 = 1;
    54: op1_13_inv01 = 1;
    56: op1_13_inv01 = 1;
    76: op1_13_inv01 = 1;
    68: op1_13_inv01 = 1;
    77: op1_13_inv01 = 1;
    61: op1_13_inv01 = 1;
    70: op1_13_inv01 = 1;
    79: op1_13_inv01 = 1;
    80: op1_13_inv01 = 1;
    62: op1_13_inv01 = 1;
    81: op1_13_inv01 = 1;
    63: op1_13_inv01 = 1;
    52: op1_13_inv01 = 1;
    84: op1_13_inv01 = 1;
    65: op1_13_inv01 = 1;
    90: op1_13_inv01 = 1;
    48: op1_13_inv01 = 1;
    67: op1_13_inv01 = 1;
    93: op1_13_inv01 = 1;
    33: op1_13_inv01 = 1;
    94: op1_13_inv01 = 1;
    28: op1_13_inv01 = 1;
    97: op1_13_inv01 = 1;
    100: op1_13_inv01 = 1;
    103: op1_13_inv01 = 1;
    104: op1_13_inv01 = 1;
    105: op1_13_inv01 = 1;
    106: op1_13_inv01 = 1;
    108: op1_13_inv01 = 1;
    109: op1_13_inv01 = 1;
    110: op1_13_inv01 = 1;
    112: op1_13_inv01 = 1;
    113: op1_13_inv01 = 1;
    118: op1_13_inv01 = 1;
    119: op1_13_inv01 = 1;
    120: op1_13_inv01 = 1;
    122: op1_13_inv01 = 1;
    125: op1_13_inv01 = 1;
    44: op1_13_inv01 = 1;
    127: op1_13_inv01 = 1;
    128: op1_13_inv01 = 1;
    129: op1_13_inv01 = 1;
    default: op1_13_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in02 = imem00_in[7:4];
    53: op1_13_in02 = reg_0042;
    64: op1_13_in02 = reg_0042;
    73: op1_13_in02 = imem06_in[15:12];
    86: op1_13_in02 = reg_0425;
    55: op1_13_in02 = reg_0821;
    74: op1_13_in02 = reg_0587;
    69: op1_13_in02 = reg_0588;
    54: op1_13_in02 = reg_0290;
    49: op1_13_in02 = reg_0022;
    75: op1_13_in02 = reg_1241;
    56: op1_13_in02 = reg_0149;
    50: op1_13_in02 = reg_0906;
    76: op1_13_in02 = reg_0864;
    71: op1_13_in02 = reg_1027;
    87: op1_13_in02 = reg_1495;
    68: op1_13_in02 = reg_1233;
    77: op1_13_in02 = reg_0727;
    61: op1_13_in02 = reg_1278;
    84: op1_13_in02 = reg_1278;
    102: op1_13_in02 = reg_1278;
    58: op1_13_in02 = reg_0173;
    90: op1_13_in02 = reg_0173;
    78: op1_13_in02 = reg_0791;
    70: op1_13_in02 = reg_0732;
    59: op1_13_in02 = reg_0262;
    79: op1_13_in02 = reg_0907;
    51: op1_13_in02 = reg_0570;
    60: op1_13_in02 = reg_1082;
    88: op1_13_in02 = reg_0999;
    80: op1_13_in02 = reg_0407;
    62: op1_13_in02 = reg_1170;
    81: op1_13_in02 = reg_0348;
    63: op1_13_in02 = reg_0724;
    52: op1_13_in02 = reg_0192;
    82: op1_13_in02 = reg_1243;
    83: op1_13_in02 = imem06_in[11:8];
    89: op1_13_in02 = reg_0107;
    46: op1_13_in02 = reg_0648;
    85: op1_13_in02 = reg_0342;
    65: op1_13_in02 = reg_0091;
    66: op1_13_in02 = reg_0899;
    48: op1_13_in02 = reg_0753;
    91: op1_13_in02 = reg_0104;
    67: op1_13_in02 = reg_0147;
    92: op1_13_in02 = reg_0143;
    93: op1_13_in02 = reg_0128;
    33: op1_13_in02 = reg_0137;
    94: op1_13_in02 = reg_0372;
    95: op1_13_in02 = reg_0236;
    96: op1_13_in02 = reg_0171;
    28: op1_13_in02 = reg_0052;
    97: op1_13_in02 = reg_0616;
    98: op1_13_in02 = reg_1277;
    116: op1_13_in02 = reg_1277;
    99: op1_13_in02 = reg_1517;
    100: op1_13_in02 = reg_1281;
    101: op1_13_in02 = reg_1147;
    103: op1_13_in02 = reg_0662;
    104: op1_13_in02 = reg_0185;
    37: op1_13_in02 = imem07_in[7:4];
    105: op1_13_in02 = reg_1214;
    106: op1_13_in02 = reg_0394;
    107: op1_13_in02 = reg_0638;
    108: op1_13_in02 = reg_1143;
    109: op1_13_in02 = reg_0011;
    110: op1_13_in02 = reg_0269;
    111: op1_13_in02 = reg_0312;
    112: op1_13_in02 = reg_0925;
    113: op1_13_in02 = reg_1325;
    114: op1_13_in02 = reg_0804;
    115: op1_13_in02 = reg_1000;
    117: op1_13_in02 = reg_0070;
    47: op1_13_in02 = reg_0131;
    118: op1_13_in02 = reg_1040;
    119: op1_13_in02 = reg_0317;
    120: op1_13_in02 = reg_0323;
    121: op1_13_in02 = imem00_in[3:0];
    122: op1_13_in02 = reg_0015;
    123: op1_13_in02 = reg_1259;
    124: op1_13_in02 = reg_0008;
    125: op1_13_in02 = reg_0115;
    126: op1_13_in02 = reg_0456;
    44: op1_13_in02 = reg_0369;
    127: op1_13_in02 = reg_0806;
    128: op1_13_in02 = reg_1053;
    129: op1_13_in02 = reg_0146;
    130: op1_13_in02 = reg_0581;
    default: op1_13_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv02 = 1;
    74: op1_13_inv02 = 1;
    69: op1_13_inv02 = 1;
    75: op1_13_inv02 = 1;
    50: op1_13_inv02 = 1;
    71: op1_13_inv02 = 1;
    68: op1_13_inv02 = 1;
    77: op1_13_inv02 = 1;
    61: op1_13_inv02 = 1;
    58: op1_13_inv02 = 1;
    59: op1_13_inv02 = 1;
    79: op1_13_inv02 = 1;
    51: op1_13_inv02 = 1;
    60: op1_13_inv02 = 1;
    88: op1_13_inv02 = 1;
    80: op1_13_inv02 = 1;
    62: op1_13_inv02 = 1;
    82: op1_13_inv02 = 1;
    83: op1_13_inv02 = 1;
    89: op1_13_inv02 = 1;
    46: op1_13_inv02 = 1;
    66: op1_13_inv02 = 1;
    92: op1_13_inv02 = 1;
    33: op1_13_inv02 = 1;
    94: op1_13_inv02 = 1;
    95: op1_13_inv02 = 1;
    96: op1_13_inv02 = 1;
    97: op1_13_inv02 = 1;
    98: op1_13_inv02 = 1;
    99: op1_13_inv02 = 1;
    101: op1_13_inv02 = 1;
    104: op1_13_inv02 = 1;
    37: op1_13_inv02 = 1;
    107: op1_13_inv02 = 1;
    109: op1_13_inv02 = 1;
    110: op1_13_inv02 = 1;
    111: op1_13_inv02 = 1;
    116: op1_13_inv02 = 1;
    118: op1_13_inv02 = 1;
    119: op1_13_inv02 = 1;
    123: op1_13_inv02 = 1;
    124: op1_13_inv02 = 1;
    126: op1_13_inv02 = 1;
    129: op1_13_inv02 = 1;
    default: op1_13_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in03 = reg_1053;
    53: op1_13_in03 = reg_0012;
    73: op1_13_in03 = reg_0636;
    86: op1_13_in03 = reg_1369;
    55: op1_13_in03 = reg_1096;
    74: op1_13_in03 = reg_0736;
    69: op1_13_in03 = reg_0590;
    103: op1_13_in03 = reg_0590;
    54: op1_13_in03 = reg_0291;
    49: op1_13_in03 = reg_0394;
    75: op1_13_in03 = reg_0121;
    56: op1_13_in03 = reg_0363;
    50: op1_13_in03 = reg_0905;
    76: op1_13_in03 = reg_0458;
    71: op1_13_in03 = reg_0249;
    87: op1_13_in03 = reg_0706;
    68: op1_13_in03 = reg_0142;
    77: op1_13_in03 = reg_0895;
    61: op1_13_in03 = reg_0841;
    58: op1_13_in03 = reg_0565;
    78: op1_13_in03 = reg_1281;
    70: op1_13_in03 = reg_0677;
    59: op1_13_in03 = reg_0836;
    79: op1_13_in03 = reg_0804;
    51: op1_13_in03 = reg_0526;
    60: op1_13_in03 = reg_0798;
    88: op1_13_in03 = reg_0328;
    80: op1_13_in03 = reg_0471;
    62: op1_13_in03 = reg_0230;
    81: op1_13_in03 = reg_0427;
    63: op1_13_in03 = reg_0871;
    52: op1_13_in03 = reg_0960;
    82: op1_13_in03 = reg_0805;
    114: op1_13_in03 = reg_0805;
    116: op1_13_in03 = reg_0805;
    83: op1_13_in03 = reg_0268;
    64: op1_13_in03 = reg_0041;
    89: op1_13_in03 = reg_0350;
    84: op1_13_in03 = reg_1079;
    46: op1_13_in03 = reg_0649;
    85: op1_13_in03 = reg_0305;
    65: op1_13_in03 = reg_0080;
    90: op1_13_in03 = reg_0391;
    66: op1_13_in03 = imem01_in[3:0];
    48: op1_13_in03 = reg_0929;
    91: op1_13_in03 = reg_0448;
    67: op1_13_in03 = reg_0149;
    92: op1_13_in03 = reg_0180;
    93: op1_13_in03 = reg_0106;
    33: op1_13_in03 = reg_0028;
    94: op1_13_in03 = reg_0716;
    95: op1_13_in03 = reg_0536;
    96: op1_13_in03 = reg_0583;
    28: op1_13_in03 = reg_0053;
    97: op1_13_in03 = reg_0186;
    98: op1_13_in03 = reg_1279;
    100: op1_13_in03 = reg_1279;
    99: op1_13_in03 = reg_0627;
    101: op1_13_in03 = reg_0097;
    102: op1_13_in03 = reg_0748;
    104: op1_13_in03 = reg_0179;
    37: op1_13_in03 = reg_0623;
    105: op1_13_in03 = reg_1077;
    106: op1_13_in03 = reg_1414;
    107: op1_13_in03 = reg_1277;
    108: op1_13_in03 = reg_0062;
    109: op1_13_in03 = reg_0013;
    110: op1_13_in03 = reg_1064;
    111: op1_13_in03 = reg_0891;
    112: op1_13_in03 = reg_0974;
    113: op1_13_in03 = reg_0426;
    115: op1_13_in03 = reg_1425;
    117: op1_13_in03 = reg_1314;
    47: op1_13_in03 = reg_0937;
    118: op1_13_in03 = reg_0451;
    119: op1_13_in03 = reg_0206;
    120: op1_13_in03 = reg_0419;
    121: op1_13_in03 = reg_0248;
    122: op1_13_in03 = reg_0050;
    123: op1_13_in03 = reg_0708;
    124: op1_13_in03 = reg_0399;
    125: op1_13_in03 = reg_0110;
    126: op1_13_in03 = imem02_in[3:0];
    44: op1_13_in03 = reg_0904;
    127: op1_13_in03 = reg_0293;
    128: op1_13_in03 = reg_1453;
    129: op1_13_in03 = reg_1032;
    130: op1_13_in03 = reg_1242;
    default: op1_13_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv03 = 1;
    73: op1_13_inv03 = 1;
    86: op1_13_inv03 = 1;
    54: op1_13_inv03 = 1;
    56: op1_13_inv03 = 1;
    71: op1_13_inv03 = 1;
    87: op1_13_inv03 = 1;
    61: op1_13_inv03 = 1;
    78: op1_13_inv03 = 1;
    59: op1_13_inv03 = 1;
    51: op1_13_inv03 = 1;
    88: op1_13_inv03 = 1;
    81: op1_13_inv03 = 1;
    82: op1_13_inv03 = 1;
    83: op1_13_inv03 = 1;
    89: op1_13_inv03 = 1;
    46: op1_13_inv03 = 1;
    85: op1_13_inv03 = 1;
    65: op1_13_inv03 = 1;
    90: op1_13_inv03 = 1;
    48: op1_13_inv03 = 1;
    67: op1_13_inv03 = 1;
    95: op1_13_inv03 = 1;
    98: op1_13_inv03 = 1;
    99: op1_13_inv03 = 1;
    100: op1_13_inv03 = 1;
    101: op1_13_inv03 = 1;
    102: op1_13_inv03 = 1;
    104: op1_13_inv03 = 1;
    37: op1_13_inv03 = 1;
    105: op1_13_inv03 = 1;
    108: op1_13_inv03 = 1;
    109: op1_13_inv03 = 1;
    114: op1_13_inv03 = 1;
    115: op1_13_inv03 = 1;
    116: op1_13_inv03 = 1;
    117: op1_13_inv03 = 1;
    47: op1_13_inv03 = 1;
    119: op1_13_inv03 = 1;
    122: op1_13_inv03 = 1;
    126: op1_13_inv03 = 1;
    127: op1_13_inv03 = 1;
    128: op1_13_inv03 = 1;
    default: op1_13_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in04 = reg_1052;
    53: op1_13_in04 = reg_0679;
    73: op1_13_in04 = reg_0529;
    86: op1_13_in04 = imem04_in[3:0];
    55: op1_13_in04 = reg_0995;
    74: op1_13_in04 = reg_0579;
    69: op1_13_in04 = reg_0562;
    54: op1_13_in04 = reg_0043;
    49: op1_13_in04 = reg_0491;
    75: op1_13_in04 = reg_0805;
    56: op1_13_in04 = reg_0875;
    50: op1_13_in04 = reg_0120;
    76: op1_13_in04 = reg_1437;
    71: op1_13_in04 = reg_0460;
    127: op1_13_in04 = reg_0460;
    87: op1_13_in04 = reg_1447;
    68: op1_13_in04 = reg_0999;
    77: op1_13_in04 = reg_0290;
    65: op1_13_in04 = reg_0290;
    61: op1_13_in04 = reg_0523;
    114: op1_13_in04 = reg_0523;
    58: op1_13_in04 = reg_0745;
    78: op1_13_in04 = reg_1277;
    70: op1_13_in04 = reg_0121;
    59: op1_13_in04 = reg_0338;
    79: op1_13_in04 = reg_1470;
    51: op1_13_in04 = reg_0527;
    60: op1_13_in04 = reg_0797;
    88: op1_13_in04 = reg_0233;
    80: op1_13_in04 = imem04_in[7:4];
    62: op1_13_in04 = reg_0162;
    81: op1_13_in04 = reg_0898;
    63: op1_13_in04 = reg_0080;
    52: op1_13_in04 = reg_0141;
    94: op1_13_in04 = reg_0141;
    82: op1_13_in04 = reg_1471;
    83: op1_13_in04 = reg_0192;
    64: op1_13_in04 = reg_0222;
    89: op1_13_in04 = reg_0479;
    84: op1_13_in04 = reg_1490;
    46: op1_13_in04 = reg_0604;
    85: op1_13_in04 = reg_0319;
    90: op1_13_in04 = reg_1104;
    66: op1_13_in04 = reg_0078;
    48: op1_13_in04 = reg_0729;
    91: op1_13_in04 = reg_0350;
    67: op1_13_in04 = reg_0401;
    92: op1_13_in04 = reg_0891;
    93: op1_13_in04 = reg_0380;
    33: op1_13_in04 = reg_0228;
    95: op1_13_in04 = reg_0064;
    96: op1_13_in04 = reg_1179;
    28: op1_13_in04 = imem07_in[7:4];
    97: op1_13_in04 = reg_0249;
    98: op1_13_in04 = reg_0672;
    99: op1_13_in04 = reg_1301;
    100: op1_13_in04 = reg_1487;
    101: op1_13_in04 = reg_0232;
    102: op1_13_in04 = reg_1141;
    103: op1_13_in04 = reg_0533;
    104: op1_13_in04 = imem03_in[11:8];
    37: op1_13_in04 = reg_0102;
    105: op1_13_in04 = reg_0342;
    106: op1_13_in04 = reg_1055;
    107: op1_13_in04 = reg_0613;
    108: op1_13_in04 = reg_0862;
    109: op1_13_in04 = reg_0895;
    110: op1_13_in04 = reg_0397;
    111: op1_13_in04 = reg_0314;
    112: op1_13_in04 = reg_0860;
    113: op1_13_in04 = reg_0427;
    115: op1_13_in04 = reg_1517;
    116: op1_13_in04 = reg_0555;
    117: op1_13_in04 = reg_0957;
    47: op1_13_in04 = reg_0090;
    118: op1_13_in04 = reg_0097;
    119: op1_13_in04 = reg_1435;
    120: op1_13_in04 = reg_0289;
    121: op1_13_in04 = reg_0803;
    122: op1_13_in04 = reg_0124;
    123: op1_13_in04 = reg_0986;
    124: op1_13_in04 = reg_0666;
    125: op1_13_in04 = reg_0718;
    126: op1_13_in04 = reg_0138;
    44: op1_13_in04 = reg_0341;
    128: op1_13_in04 = reg_1230;
    129: op1_13_in04 = reg_1034;
    130: op1_13_in04 = reg_0926;
    default: op1_13_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv04 = 1;
    53: op1_13_inv04 = 1;
    73: op1_13_inv04 = 1;
    55: op1_13_inv04 = 1;
    74: op1_13_inv04 = 1;
    75: op1_13_inv04 = 1;
    50: op1_13_inv04 = 1;
    76: op1_13_inv04 = 1;
    71: op1_13_inv04 = 1;
    87: op1_13_inv04 = 1;
    61: op1_13_inv04 = 1;
    58: op1_13_inv04 = 1;
    70: op1_13_inv04 = 1;
    79: op1_13_inv04 = 1;
    51: op1_13_inv04 = 1;
    88: op1_13_inv04 = 1;
    80: op1_13_inv04 = 1;
    63: op1_13_inv04 = 1;
    82: op1_13_inv04 = 1;
    64: op1_13_inv04 = 1;
    89: op1_13_inv04 = 1;
    84: op1_13_inv04 = 1;
    46: op1_13_inv04 = 1;
    85: op1_13_inv04 = 1;
    65: op1_13_inv04 = 1;
    66: op1_13_inv04 = 1;
    48: op1_13_inv04 = 1;
    91: op1_13_inv04 = 1;
    67: op1_13_inv04 = 1;
    92: op1_13_inv04 = 1;
    93: op1_13_inv04 = 1;
    94: op1_13_inv04 = 1;
    95: op1_13_inv04 = 1;
    96: op1_13_inv04 = 1;
    28: op1_13_inv04 = 1;
    97: op1_13_inv04 = 1;
    98: op1_13_inv04 = 1;
    99: op1_13_inv04 = 1;
    100: op1_13_inv04 = 1;
    101: op1_13_inv04 = 1;
    102: op1_13_inv04 = 1;
    103: op1_13_inv04 = 1;
    106: op1_13_inv04 = 1;
    109: op1_13_inv04 = 1;
    110: op1_13_inv04 = 1;
    114: op1_13_inv04 = 1;
    115: op1_13_inv04 = 1;
    117: op1_13_inv04 = 1;
    120: op1_13_inv04 = 1;
    123: op1_13_inv04 = 1;
    124: op1_13_inv04 = 1;
    126: op1_13_inv04 = 1;
    130: op1_13_inv04 = 1;
    default: op1_13_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in05 = reg_0523;
    53: op1_13_in05 = reg_0446;
    64: op1_13_in05 = reg_0446;
    73: op1_13_in05 = reg_0345;
    86: op1_13_in05 = imem04_in[11:8];
    55: op1_13_in05 = imem07_in[7:4];
    74: op1_13_in05 = reg_1299;
    69: op1_13_in05 = reg_0473;
    54: op1_13_in05 = reg_0044;
    49: op1_13_in05 = reg_0224;
    75: op1_13_in05 = reg_0218;
    56: op1_13_in05 = reg_0078;
    50: op1_13_in05 = reg_0397;
    76: op1_13_in05 = reg_1435;
    71: op1_13_in05 = reg_0476;
    87: op1_13_in05 = reg_0177;
    68: op1_13_in05 = reg_0314;
    77: op1_13_in05 = reg_0283;
    61: op1_13_in05 = reg_1230;
    58: op1_13_in05 = reg_0937;
    78: op1_13_in05 = reg_1490;
    70: op1_13_in05 = reg_0707;
    59: op1_13_in05 = reg_0097;
    79: op1_13_in05 = reg_1454;
    51: op1_13_in05 = reg_0522;
    60: op1_13_in05 = reg_0795;
    88: op1_13_in05 = reg_0699;
    80: op1_13_in05 = reg_0320;
    62: op1_13_in05 = reg_0998;
    81: op1_13_in05 = reg_0696;
    63: op1_13_in05 = reg_0077;
    52: op1_13_in05 = reg_0636;
    82: op1_13_in05 = reg_1469;
    83: op1_13_in05 = reg_0720;
    89: op1_13_in05 = reg_0673;
    84: op1_13_in05 = reg_0615;
    46: op1_13_in05 = reg_0564;
    90: op1_13_in05 = reg_0564;
    85: op1_13_in05 = reg_1189;
    65: op1_13_in05 = reg_0222;
    66: op1_13_in05 = reg_0290;
    48: op1_13_in05 = imem06_in[7:4];
    91: op1_13_in05 = reg_0378;
    67: op1_13_in05 = reg_0874;
    92: op1_13_in05 = reg_0989;
    93: op1_13_in05 = reg_0381;
    33: op1_13_in05 = reg_0004;
    94: op1_13_in05 = reg_0586;
    95: op1_13_in05 = reg_0063;
    96: op1_13_in05 = reg_0270;
    97: op1_13_in05 = reg_0229;
    98: op1_13_in05 = reg_1491;
    99: op1_13_in05 = reg_0558;
    100: op1_13_in05 = reg_1027;
    116: op1_13_in05 = reg_1027;
    101: op1_13_in05 = reg_0061;
    102: op1_13_in05 = reg_1489;
    103: op1_13_in05 = imem02_in[11:8];
    104: op1_13_in05 = reg_0557;
    37: op1_13_in05 = reg_0103;
    105: op1_13_in05 = reg_0862;
    106: op1_13_in05 = reg_1315;
    107: op1_13_in05 = reg_0580;
    121: op1_13_in05 = reg_0580;
    108: op1_13_in05 = imem04_in[3:0];
    109: op1_13_in05 = reg_0008;
    110: op1_13_in05 = reg_0192;
    111: op1_13_in05 = reg_0957;
    112: op1_13_in05 = reg_0827;
    113: op1_13_in05 = reg_0443;
    114: op1_13_in05 = reg_0155;
    127: op1_13_in05 = reg_0155;
    115: op1_13_in05 = reg_1314;
    117: op1_13_in05 = reg_1208;
    47: op1_13_in05 = reg_0872;
    118: op1_13_in05 = reg_0033;
    119: op1_13_in05 = imem06_in[15:12];
    120: op1_13_in05 = reg_1202;
    122: op1_13_in05 = reg_0087;
    123: op1_13_in05 = reg_1168;
    124: op1_13_in05 = reg_0608;
    125: op1_13_in05 = reg_0714;
    126: op1_13_in05 = reg_1493;
    44: op1_13_in05 = reg_0199;
    128: op1_13_in05 = reg_1418;
    129: op1_13_in05 = reg_0360;
    130: op1_13_in05 = reg_1081;
    default: op1_13_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_13_inv05 = 1;
    55: op1_13_inv05 = 1;
    75: op1_13_inv05 = 1;
    56: op1_13_inv05 = 1;
    71: op1_13_inv05 = 1;
    87: op1_13_inv05 = 1;
    68: op1_13_inv05 = 1;
    61: op1_13_inv05 = 1;
    58: op1_13_inv05 = 1;
    78: op1_13_inv05 = 1;
    70: op1_13_inv05 = 1;
    51: op1_13_inv05 = 1;
    88: op1_13_inv05 = 1;
    82: op1_13_inv05 = 1;
    89: op1_13_inv05 = 1;
    90: op1_13_inv05 = 1;
    66: op1_13_inv05 = 1;
    48: op1_13_inv05 = 1;
    91: op1_13_inv05 = 1;
    67: op1_13_inv05 = 1;
    93: op1_13_inv05 = 1;
    96: op1_13_inv05 = 1;
    99: op1_13_inv05 = 1;
    100: op1_13_inv05 = 1;
    102: op1_13_inv05 = 1;
    37: op1_13_inv05 = 1;
    105: op1_13_inv05 = 1;
    107: op1_13_inv05 = 1;
    109: op1_13_inv05 = 1;
    110: op1_13_inv05 = 1;
    111: op1_13_inv05 = 1;
    114: op1_13_inv05 = 1;
    120: op1_13_inv05 = 1;
    125: op1_13_inv05 = 1;
    126: op1_13_inv05 = 1;
    129: op1_13_inv05 = 1;
    default: op1_13_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in06 = reg_0293;
    53: op1_13_in06 = reg_0254;
    73: op1_13_in06 = reg_1225;
    86: op1_13_in06 = reg_0531;
    55: op1_13_in06 = imem07_in[15:12];
    74: op1_13_in06 = reg_0833;
    69: op1_13_in06 = reg_0432;
    54: op1_13_in06 = reg_0662;
    49: op1_13_in06 = reg_0310;
    75: op1_13_in06 = reg_1230;
    100: op1_13_in06 = reg_1230;
    56: op1_13_in06 = reg_0282;
    50: op1_13_in06 = reg_0825;
    76: op1_13_in06 = reg_0192;
    71: op1_13_in06 = reg_0927;
    87: op1_13_in06 = reg_1033;
    68: op1_13_in06 = reg_1199;
    77: op1_13_in06 = reg_0043;
    61: op1_13_in06 = reg_0958;
    58: op1_13_in06 = reg_0449;
    78: op1_13_in06 = reg_1243;
    70: op1_13_in06 = imem03_in[7:4];
    59: op1_13_in06 = reg_0236;
    79: op1_13_in06 = reg_1459;
    82: op1_13_in06 = reg_1459;
    51: op1_13_in06 = reg_0459;
    114: op1_13_in06 = reg_0459;
    60: op1_13_in06 = reg_0370;
    88: op1_13_in06 = reg_0235;
    80: op1_13_in06 = reg_0837;
    62: op1_13_in06 = imem07_in[11:8];
    81: op1_13_in06 = reg_0534;
    63: op1_13_in06 = reg_0290;
    52: op1_13_in06 = reg_0263;
    83: op1_13_in06 = reg_0780;
    64: op1_13_in06 = reg_0699;
    89: op1_13_in06 = reg_0426;
    84: op1_13_in06 = reg_1470;
    46: op1_13_in06 = reg_0940;
    85: op1_13_in06 = reg_0016;
    65: op1_13_in06 = reg_0486;
    107: op1_13_in06 = reg_0486;
    90: op1_13_in06 = reg_0334;
    66: op1_13_in06 = reg_0088;
    48: op1_13_in06 = reg_0979;
    91: op1_13_in06 = reg_0673;
    67: op1_13_in06 = reg_0077;
    92: op1_13_in06 = reg_1517;
    93: op1_13_in06 = reg_0897;
    33: op1_13_in06 = reg_0001;
    94: op1_13_in06 = reg_0527;
    95: op1_13_in06 = reg_0633;
    96: op1_13_in06 = reg_0215;
    97: op1_13_in06 = reg_0886;
    98: op1_13_in06 = reg_0841;
    99: op1_13_in06 = reg_0880;
    101: op1_13_in06 = reg_0369;
    102: op1_13_in06 = reg_1491;
    103: op1_13_in06 = reg_0423;
    104: op1_13_in06 = reg_0600;
    37: op1_13_in06 = reg_0052;
    105: op1_13_in06 = reg_0336;
    106: op1_13_in06 = reg_0298;
    108: op1_13_in06 = reg_0904;
    109: op1_13_in06 = reg_0607;
    110: op1_13_in06 = reg_1437;
    111: op1_13_in06 = reg_1300;
    112: op1_13_in06 = reg_1179;
    113: op1_13_in06 = reg_1369;
    115: op1_13_in06 = reg_0350;
    116: op1_13_in06 = reg_1454;
    117: op1_13_in06 = reg_0104;
    47: op1_13_in06 = reg_0197;
    118: op1_13_in06 = reg_0061;
    119: op1_13_in06 = reg_0795;
    120: op1_13_in06 = reg_0017;
    121: op1_13_in06 = reg_0554;
    122: op1_13_in06 = imem07_in[7:4];
    123: op1_13_in06 = reg_0040;
    124: op1_13_in06 = reg_0839;
    125: op1_13_in06 = reg_0141;
    126: op1_13_in06 = reg_0822;
    44: op1_13_in06 = reg_0305;
    127: op1_13_in06 = reg_1406;
    128: op1_13_in06 = reg_0524;
    129: op1_13_in06 = reg_0363;
    130: op1_13_in06 = reg_0501;
    default: op1_13_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv06 = 1;
    74: op1_13_inv06 = 1;
    69: op1_13_inv06 = 1;
    54: op1_13_inv06 = 1;
    56: op1_13_inv06 = 1;
    76: op1_13_inv06 = 1;
    71: op1_13_inv06 = 1;
    87: op1_13_inv06 = 1;
    61: op1_13_inv06 = 1;
    58: op1_13_inv06 = 1;
    78: op1_13_inv06 = 1;
    79: op1_13_inv06 = 1;
    60: op1_13_inv06 = 1;
    80: op1_13_inv06 = 1;
    52: op1_13_inv06 = 1;
    83: op1_13_inv06 = 1;
    89: op1_13_inv06 = 1;
    84: op1_13_inv06 = 1;
    46: op1_13_inv06 = 1;
    90: op1_13_inv06 = 1;
    66: op1_13_inv06 = 1;
    48: op1_13_inv06 = 1;
    91: op1_13_inv06 = 1;
    67: op1_13_inv06 = 1;
    92: op1_13_inv06 = 1;
    96: op1_13_inv06 = 1;
    98: op1_13_inv06 = 1;
    99: op1_13_inv06 = 1;
    100: op1_13_inv06 = 1;
    101: op1_13_inv06 = 1;
    103: op1_13_inv06 = 1;
    104: op1_13_inv06 = 1;
    37: op1_13_inv06 = 1;
    105: op1_13_inv06 = 1;
    107: op1_13_inv06 = 1;
    108: op1_13_inv06 = 1;
    109: op1_13_inv06 = 1;
    110: op1_13_inv06 = 1;
    111: op1_13_inv06 = 1;
    114: op1_13_inv06 = 1;
    47: op1_13_inv06 = 1;
    122: op1_13_inv06 = 1;
    124: op1_13_inv06 = 1;
    125: op1_13_inv06 = 1;
    44: op1_13_inv06 = 1;
    130: op1_13_inv06 = 1;
    default: op1_13_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in07 = reg_1027;
    53: op1_13_in07 = reg_0629;
    73: op1_13_in07 = reg_0296;
    86: op1_13_in07 = reg_0297;
    55: op1_13_in07 = reg_0224;
    74: op1_13_in07 = reg_0136;
    69: op1_13_in07 = reg_0326;
    54: op1_13_in07 = reg_0606;
    49: op1_13_in07 = reg_0867;
    75: op1_13_in07 = reg_0155;
    56: op1_13_in07 = reg_0043;
    50: op1_13_in07 = reg_0827;
    76: op1_13_in07 = reg_1504;
    71: op1_13_in07 = reg_0883;
    87: op1_13_in07 = reg_0707;
    68: op1_13_in07 = reg_1092;
    77: op1_13_in07 = reg_0169;
    109: op1_13_in07 = reg_0169;
    61: op1_13_in07 = reg_1148;
    58: op1_13_in07 = reg_0204;
    78: op1_13_in07 = imem00_in[7:4];
    70: op1_13_in07 = reg_1033;
    59: op1_13_in07 = reg_0209;
    80: op1_13_in07 = reg_0209;
    79: op1_13_in07 = reg_0987;
    51: op1_13_in07 = reg_0271;
    60: op1_13_in07 = reg_0454;
    88: op1_13_in07 = reg_0261;
    62: op1_13_in07 = reg_0922;
    81: op1_13_in07 = reg_0341;
    63: op1_13_in07 = reg_0277;
    52: op1_13_in07 = reg_0622;
    82: op1_13_in07 = reg_1432;
    100: op1_13_in07 = reg_1432;
    83: op1_13_in07 = reg_0116;
    112: op1_13_in07 = reg_0116;
    64: op1_13_in07 = imem02_in[7:4];
    89: op1_13_in07 = reg_0411;
    84: op1_13_in07 = reg_0218;
    46: op1_13_in07 = reg_0939;
    85: op1_13_in07 = reg_0210;
    65: op1_13_in07 = reg_0605;
    90: op1_13_in07 = reg_0794;
    66: op1_13_in07 = reg_0291;
    48: op1_13_in07 = reg_0397;
    91: op1_13_in07 = reg_0348;
    115: op1_13_in07 = reg_0348;
    67: op1_13_in07 = reg_0012;
    92: op1_13_in07 = reg_1314;
    93: op1_13_in07 = reg_0800;
    33: op1_13_in07 = reg_0002;
    94: op1_13_in07 = reg_0289;
    95: op1_13_in07 = reg_1488;
    96: op1_13_in07 = imem07_in[7:4];
    97: op1_13_in07 = reg_0134;
    98: op1_13_in07 = reg_0580;
    99: op1_13_in07 = reg_0448;
    117: op1_13_in07 = reg_0448;
    101: op1_13_in07 = reg_1143;
    102: op1_13_in07 = reg_0805;
    103: op1_13_in07 = reg_1018;
    104: op1_13_in07 = reg_0191;
    37: op1_13_in07 = reg_0483;
    105: op1_13_in07 = reg_1502;
    106: op1_13_in07 = reg_0894;
    107: op1_13_in07 = reg_1052;
    108: op1_13_in07 = reg_1107;
    110: op1_13_in07 = reg_0751;
    111: op1_13_in07 = reg_0108;
    113: op1_13_in07 = reg_0535;
    114: op1_13_in07 = reg_0524;
    116: op1_13_in07 = reg_0353;
    47: op1_13_in07 = reg_0184;
    118: op1_13_in07 = reg_0369;
    119: op1_13_in07 = reg_0372;
    120: op1_13_in07 = reg_0051;
    121: op1_13_in07 = reg_1053;
    122: op1_13_in07 = reg_0994;
    123: op1_13_in07 = reg_0733;
    124: op1_13_in07 = reg_0533;
    126: op1_13_in07 = reg_0533;
    125: op1_13_in07 = reg_0373;
    44: op1_13_in07 = reg_0862;
    127: op1_13_in07 = reg_0821;
    128: op1_13_in07 = reg_0881;
    129: op1_13_in07 = reg_0901;
    130: op1_13_in07 = reg_0248;
    default: op1_13_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv07 = 1;
    73: op1_13_inv07 = 1;
    74: op1_13_inv07 = 1;
    54: op1_13_inv07 = 1;
    75: op1_13_inv07 = 1;
    68: op1_13_inv07 = 1;
    77: op1_13_inv07 = 1;
    59: op1_13_inv07 = 1;
    60: op1_13_inv07 = 1;
    80: op1_13_inv07 = 1;
    63: op1_13_inv07 = 1;
    82: op1_13_inv07 = 1;
    64: op1_13_inv07 = 1;
    84: op1_13_inv07 = 1;
    46: op1_13_inv07 = 1;
    85: op1_13_inv07 = 1;
    65: op1_13_inv07 = 1;
    48: op1_13_inv07 = 1;
    67: op1_13_inv07 = 1;
    93: op1_13_inv07 = 1;
    33: op1_13_inv07 = 1;
    94: op1_13_inv07 = 1;
    99: op1_13_inv07 = 1;
    102: op1_13_inv07 = 1;
    104: op1_13_inv07 = 1;
    106: op1_13_inv07 = 1;
    107: op1_13_inv07 = 1;
    108: op1_13_inv07 = 1;
    109: op1_13_inv07 = 1;
    110: op1_13_inv07 = 1;
    114: op1_13_inv07 = 1;
    47: op1_13_inv07 = 1;
    119: op1_13_inv07 = 1;
    120: op1_13_inv07 = 1;
    123: op1_13_inv07 = 1;
    124: op1_13_inv07 = 1;
    126: op1_13_inv07 = 1;
    44: op1_13_inv07 = 1;
    128: op1_13_inv07 = 1;
    129: op1_13_inv07 = 1;
    default: op1_13_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in08 = reg_1230;
    53: op1_13_in08 = reg_0606;
    73: op1_13_in08 = reg_0419;
    86: op1_13_in08 = reg_1198;
    55: op1_13_in08 = reg_0894;
    74: op1_13_in08 = reg_0877;
    69: op1_13_in08 = reg_0778;
    54: op1_13_in08 = reg_0922;
    49: op1_13_in08 = reg_0673;
    75: op1_13_in08 = reg_0883;
    56: op1_13_in08 = reg_0041;
    50: op1_13_in08 = reg_0116;
    76: op1_13_in08 = reg_0984;
    71: op1_13_in08 = reg_0353;
    87: op1_13_in08 = reg_1314;
    68: op1_13_in08 = reg_1208;
    77: op1_13_in08 = reg_0608;
    61: op1_13_in08 = reg_0887;
    58: op1_13_in08 = reg_0751;
    78: op1_13_in08 = reg_0804;
    70: op1_13_in08 = reg_0638;
    59: op1_13_in08 = reg_0035;
    95: op1_13_in08 = reg_0035;
    79: op1_13_in08 = reg_1201;
    51: op1_13_in08 = reg_0067;
    60: op1_13_in08 = reg_0932;
    88: op1_13_in08 = reg_0216;
    80: op1_13_in08 = reg_0470;
    62: op1_13_in08 = reg_0310;
    81: op1_13_in08 = reg_0493;
    63: op1_13_in08 = reg_0282;
    52: op1_13_in08 = reg_0529;
    82: op1_13_in08 = reg_1406;
    83: op1_13_in08 = reg_0109;
    64: op1_13_in08 = reg_1029;
    89: op1_13_in08 = imem04_in[15:12];
    84: op1_13_in08 = reg_1052;
    121: op1_13_in08 = reg_1052;
    46: op1_13_in08 = reg_0302;
    85: op1_13_in08 = reg_0708;
    65: op1_13_in08 = reg_0530;
    90: op1_13_in08 = reg_0873;
    66: op1_13_in08 = reg_0222;
    48: op1_13_in08 = reg_0396;
    91: op1_13_in08 = reg_0411;
    67: op1_13_in08 = reg_1140;
    92: op1_13_in08 = reg_0558;
    93: op1_13_in08 = reg_0327;
    33: op1_13_in08 = reg_0084;
    94: op1_13_in08 = reg_0583;
    96: op1_13_in08 = reg_0867;
    97: op1_13_in08 = reg_0075;
    98: op1_13_in08 = reg_1027;
    99: op1_13_in08 = reg_0541;
    100: op1_13_in08 = reg_0155;
    101: op1_13_in08 = reg_0487;
    102: op1_13_in08 = reg_0186;
    103: op1_13_in08 = reg_0839;
    104: op1_13_in08 = reg_0180;
    37: op1_13_in08 = reg_0484;
    105: op1_13_in08 = reg_0020;
    106: op1_13_in08 = reg_1056;
    107: op1_13_in08 = reg_0293;
    108: op1_13_in08 = reg_1502;
    109: op1_13_in08 = reg_0879;
    110: op1_13_in08 = reg_0869;
    111: op1_13_in08 = reg_0107;
    112: op1_13_in08 = reg_0110;
    113: op1_13_in08 = reg_0337;
    114: op1_13_in08 = reg_0821;
    115: op1_13_in08 = reg_0263;
    116: op1_13_in08 = reg_0351;
    117: op1_13_in08 = reg_0378;
    47: op1_13_in08 = reg_0130;
    118: op1_13_in08 = reg_0582;
    119: op1_13_in08 = reg_0929;
    120: op1_13_in08 = reg_0394;
    122: op1_13_in08 = reg_1060;
    123: op1_13_in08 = reg_0176;
    124: op1_13_in08 = reg_0495;
    125: op1_13_in08 = reg_0584;
    126: op1_13_in08 = reg_0472;
    44: op1_13_in08 = reg_0338;
    127: op1_13_in08 = reg_1405;
    128: op1_13_in08 = reg_0352;
    129: op1_13_in08 = reg_0079;
    130: op1_13_in08 = reg_0554;
    default: op1_13_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_13_inv08 = 1;
    69: op1_13_inv08 = 1;
    75: op1_13_inv08 = 1;
    50: op1_13_inv08 = 1;
    71: op1_13_inv08 = 1;
    87: op1_13_inv08 = 1;
    77: op1_13_inv08 = 1;
    61: op1_13_inv08 = 1;
    58: op1_13_inv08 = 1;
    78: op1_13_inv08 = 1;
    88: op1_13_inv08 = 1;
    62: op1_13_inv08 = 1;
    52: op1_13_inv08 = 1;
    64: op1_13_inv08 = 1;
    85: op1_13_inv08 = 1;
    90: op1_13_inv08 = 1;
    66: op1_13_inv08 = 1;
    48: op1_13_inv08 = 1;
    92: op1_13_inv08 = 1;
    93: op1_13_inv08 = 1;
    33: op1_13_inv08 = 1;
    94: op1_13_inv08 = 1;
    95: op1_13_inv08 = 1;
    97: op1_13_inv08 = 1;
    98: op1_13_inv08 = 1;
    102: op1_13_inv08 = 1;
    103: op1_13_inv08 = 1;
    37: op1_13_inv08 = 1;
    106: op1_13_inv08 = 1;
    109: op1_13_inv08 = 1;
    111: op1_13_inv08 = 1;
    112: op1_13_inv08 = 1;
    113: op1_13_inv08 = 1;
    115: op1_13_inv08 = 1;
    116: op1_13_inv08 = 1;
    117: op1_13_inv08 = 1;
    47: op1_13_inv08 = 1;
    122: op1_13_inv08 = 1;
    123: op1_13_inv08 = 1;
    124: op1_13_inv08 = 1;
    125: op1_13_inv08 = 1;
    44: op1_13_inv08 = 1;
    127: op1_13_inv08 = 1;
    128: op1_13_inv08 = 1;
    default: op1_13_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in09 = reg_0961;
    79: op1_13_in09 = reg_0961;
    53: op1_13_in09 = reg_0589;
    73: op1_13_in09 = reg_1202;
    86: op1_13_in09 = reg_1233;
    55: op1_13_in09 = reg_0867;
    74: op1_13_in09 = reg_0733;
    69: op1_13_in09 = reg_0970;
    124: op1_13_in09 = reg_0970;
    54: op1_13_in09 = reg_0563;
    49: op1_13_in09 = reg_0159;
    75: op1_13_in09 = reg_0886;
    61: op1_13_in09 = reg_0886;
    56: op1_13_in09 = reg_0010;
    50: op1_13_in09 = reg_0109;
    76: op1_13_in09 = reg_0116;
    71: op1_13_in09 = reg_0722;
    87: op1_13_in09 = reg_0957;
    68: op1_13_in09 = imem03_in[7:4];
    77: op1_13_in09 = reg_0561;
    58: op1_13_in09 = reg_0931;
    78: op1_13_in09 = reg_0803;
    70: op1_13_in09 = reg_1325;
    59: op1_13_in09 = reg_0793;
    51: op1_13_in09 = reg_0023;
    60: op1_13_in09 = reg_0470;
    95: op1_13_in09 = reg_0470;
    88: op1_13_in09 = reg_0962;
    80: op1_13_in09 = reg_0251;
    62: op1_13_in09 = reg_0703;
    81: op1_13_in09 = reg_1340;
    63: op1_13_in09 = reg_0278;
    52: op1_13_in09 = reg_0527;
    82: op1_13_in09 = reg_0821;
    83: op1_13_in09 = reg_1303;
    64: op1_13_in09 = reg_0976;
    89: op1_13_in09 = reg_1384;
    84: op1_13_in09 = reg_1459;
    46: op1_13_in09 = reg_0873;
    85: op1_13_in09 = reg_0175;
    65: op1_13_in09 = reg_1018;
    90: op1_13_in09 = reg_1485;
    66: op1_13_in09 = reg_0486;
    48: op1_13_in09 = reg_0720;
    91: op1_13_in09 = reg_0247;
    67: op1_13_in09 = reg_0605;
    92: op1_13_in09 = reg_0104;
    93: op1_13_in09 = reg_0227;
    94: op1_13_in09 = reg_0214;
    96: op1_13_in09 = reg_1439;
    97: op1_13_in09 = reg_0058;
    98: op1_13_in09 = reg_0249;
    99: op1_13_in09 = reg_0218;
    100: op1_13_in09 = reg_1418;
    101: op1_13_in09 = reg_0095;
    102: op1_13_in09 = reg_1454;
    103: op1_13_in09 = reg_0822;
    104: op1_13_in09 = reg_1313;
    105: op1_13_in09 = reg_1059;
    106: op1_13_in09 = reg_1350;
    107: op1_13_in09 = reg_0221;
    108: op1_13_in09 = reg_0021;
    109: op1_13_in09 = reg_0056;
    110: op1_13_in09 = reg_0752;
    111: op1_13_in09 = reg_0113;
    112: op1_13_in09 = reg_0718;
    113: op1_13_in09 = reg_0531;
    114: op1_13_in09 = reg_0388;
    115: op1_13_in09 = reg_1369;
    116: op1_13_in09 = reg_0440;
    117: op1_13_in09 = reg_0673;
    47: op1_13_in09 = reg_0275;
    118: op1_13_in09 = reg_0837;
    119: op1_13_in09 = reg_1064;
    120: op1_13_in09 = reg_0994;
    121: op1_13_in09 = reg_1027;
    122: op1_13_in09 = reg_0922;
    123: op1_13_in09 = reg_0340;
    125: op1_13_in09 = reg_0522;
    126: op1_13_in09 = reg_0631;
    44: op1_13_in09 = reg_0336;
    127: op1_13_in09 = reg_0928;
    128: op1_13_in09 = reg_0201;
    129: op1_13_in09 = reg_0402;
    130: op1_13_in09 = reg_0640;
    default: op1_13_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv09 = 1;
    53: op1_13_inv09 = 1;
    73: op1_13_inv09 = 1;
    86: op1_13_inv09 = 1;
    69: op1_13_inv09 = 1;
    54: op1_13_inv09 = 1;
    49: op1_13_inv09 = 1;
    75: op1_13_inv09 = 1;
    56: op1_13_inv09 = 1;
    76: op1_13_inv09 = 1;
    71: op1_13_inv09 = 1;
    87: op1_13_inv09 = 1;
    77: op1_13_inv09 = 1;
    58: op1_13_inv09 = 1;
    78: op1_13_inv09 = 1;
    70: op1_13_inv09 = 1;
    59: op1_13_inv09 = 1;
    51: op1_13_inv09 = 1;
    80: op1_13_inv09 = 1;
    62: op1_13_inv09 = 1;
    63: op1_13_inv09 = 1;
    52: op1_13_inv09 = 1;
    82: op1_13_inv09 = 1;
    83: op1_13_inv09 = 1;
    64: op1_13_inv09 = 1;
    89: op1_13_inv09 = 1;
    84: op1_13_inv09 = 1;
    65: op1_13_inv09 = 1;
    90: op1_13_inv09 = 1;
    48: op1_13_inv09 = 1;
    67: op1_13_inv09 = 1;
    92: op1_13_inv09 = 1;
    94: op1_13_inv09 = 1;
    95: op1_13_inv09 = 1;
    96: op1_13_inv09 = 1;
    99: op1_13_inv09 = 1;
    105: op1_13_inv09 = 1;
    106: op1_13_inv09 = 1;
    107: op1_13_inv09 = 1;
    108: op1_13_inv09 = 1;
    111: op1_13_inv09 = 1;
    112: op1_13_inv09 = 1;
    118: op1_13_inv09 = 1;
    119: op1_13_inv09 = 1;
    120: op1_13_inv09 = 1;
    123: op1_13_inv09 = 1;
    125: op1_13_inv09 = 1;
    126: op1_13_inv09 = 1;
    127: op1_13_inv09 = 1;
    128: op1_13_inv09 = 1;
    129: op1_13_inv09 = 1;
    default: op1_13_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in10 = reg_0460;
    53: op1_13_in10 = reg_0533;
    73: op1_13_in10 = reg_1179;
    86: op1_13_in10 = reg_0796;
    55: op1_13_in10 = reg_0297;
    74: op1_13_in10 = reg_0879;
    69: op1_13_in10 = reg_0972;
    54: op1_13_in10 = reg_0560;
    49: op1_13_in10 = reg_0158;
    106: op1_13_in10 = reg_0158;
    75: op1_13_in10 = reg_0351;
    56: op1_13_in10 = reg_0133;
    50: op1_13_in10 = reg_0619;
    76: op1_13_in10 = reg_0636;
    83: op1_13_in10 = reg_0636;
    71: op1_13_in10 = reg_0409;
    100: op1_13_in10 = reg_0409;
    87: op1_13_in10 = imem03_in[15:12];
    68: op1_13_in10 = reg_0840;
    77: op1_13_in10 = reg_0981;
    61: op1_13_in10 = reg_0416;
    116: op1_13_in10 = reg_0416;
    58: op1_13_in10 = reg_1105;
    78: op1_13_in10 = reg_1052;
    70: op1_13_in10 = reg_0143;
    59: op1_13_in10 = reg_1104;
    79: op1_13_in10 = reg_1432;
    98: op1_13_in10 = reg_1432;
    51: op1_13_in10 = reg_0046;
    60: op1_13_in10 = reg_0488;
    88: op1_13_in10 = reg_0891;
    80: op1_13_in10 = reg_0877;
    62: op1_13_in10 = reg_0775;
    81: op1_13_in10 = reg_1257;
    63: op1_13_in10 = reg_0662;
    66: op1_13_in10 = reg_0662;
    52: op1_13_in10 = reg_0296;
    82: op1_13_in10 = reg_1405;
    64: op1_13_in10 = reg_0605;
    89: op1_13_in10 = reg_1369;
    84: op1_13_in10 = reg_0821;
    46: op1_13_in10 = reg_0872;
    85: op1_13_in10 = reg_0578;
    65: op1_13_in10 = reg_0472;
    90: op1_13_in10 = reg_0492;
    48: op1_13_in10 = reg_0372;
    91: op1_13_in10 = reg_0181;
    67: op1_13_in10 = reg_0532;
    92: op1_13_in10 = reg_0378;
    93: op1_13_in10 = reg_1145;
    94: op1_13_in10 = reg_0998;
    95: op1_13_in10 = reg_0750;
    96: op1_13_in10 = reg_0324;
    97: op1_13_in10 = reg_0089;
    99: op1_13_in10 = reg_0673;
    101: op1_13_in10 = reg_0019;
    102: op1_13_in10 = reg_1453;
    103: op1_13_in10 = reg_1074;
    104: op1_13_in10 = reg_0957;
    105: op1_13_in10 = reg_0833;
    107: op1_13_in10 = reg_1201;
    108: op1_13_in10 = reg_0986;
    109: op1_13_in10 = reg_0588;
    110: op1_13_in10 = reg_0265;
    111: op1_13_in10 = reg_0541;
    112: op1_13_in10 = reg_0398;
    113: op1_13_in10 = reg_0552;
    114: op1_13_in10 = reg_0075;
    115: op1_13_in10 = reg_1368;
    117: op1_13_in10 = reg_0425;
    47: op1_13_in10 = reg_0929;
    118: op1_13_in10 = reg_0117;
    119: op1_13_in10 = reg_0161;
    120: op1_13_in10 = reg_0225;
    121: op1_13_in10 = reg_1230;
    122: op1_13_in10 = reg_0135;
    123: op1_13_in10 = reg_0562;
    124: op1_13_in10 = reg_1433;
    125: op1_13_in10 = reg_0132;
    126: op1_13_in10 = reg_0473;
    44: op1_13_in10 = reg_0097;
    127: op1_13_in10 = reg_0927;
    128: op1_13_in10 = reg_0057;
    129: op1_13_in10 = reg_0634;
    130: op1_13_in10 = reg_0293;
    default: op1_13_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv10 = 1;
    73: op1_13_inv10 = 1;
    86: op1_13_inv10 = 1;
    69: op1_13_inv10 = 1;
    49: op1_13_inv10 = 1;
    56: op1_13_inv10 = 1;
    50: op1_13_inv10 = 1;
    76: op1_13_inv10 = 1;
    87: op1_13_inv10 = 1;
    77: op1_13_inv10 = 1;
    61: op1_13_inv10 = 1;
    58: op1_13_inv10 = 1;
    78: op1_13_inv10 = 1;
    70: op1_13_inv10 = 1;
    59: op1_13_inv10 = 1;
    51: op1_13_inv10 = 1;
    60: op1_13_inv10 = 1;
    80: op1_13_inv10 = 1;
    62: op1_13_inv10 = 1;
    63: op1_13_inv10 = 1;
    83: op1_13_inv10 = 1;
    64: op1_13_inv10 = 1;
    46: op1_13_inv10 = 1;
    85: op1_13_inv10 = 1;
    48: op1_13_inv10 = 1;
    91: op1_13_inv10 = 1;
    67: op1_13_inv10 = 1;
    94: op1_13_inv10 = 1;
    96: op1_13_inv10 = 1;
    99: op1_13_inv10 = 1;
    102: op1_13_inv10 = 1;
    103: op1_13_inv10 = 1;
    107: op1_13_inv10 = 1;
    108: op1_13_inv10 = 1;
    109: op1_13_inv10 = 1;
    110: op1_13_inv10 = 1;
    111: op1_13_inv10 = 1;
    112: op1_13_inv10 = 1;
    113: op1_13_inv10 = 1;
    114: op1_13_inv10 = 1;
    115: op1_13_inv10 = 1;
    116: op1_13_inv10 = 1;
    47: op1_13_inv10 = 1;
    118: op1_13_inv10 = 1;
    120: op1_13_inv10 = 1;
    122: op1_13_inv10 = 1;
    126: op1_13_inv10 = 1;
    128: op1_13_inv10 = 1;
    129: op1_13_inv10 = 1;
    default: op1_13_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in11 = reg_0229;
    53: op1_13_in11 = imem02_in[11:8];
    73: op1_13_in11 = reg_0270;
    86: op1_13_in11 = reg_0598;
    55: op1_13_in11 = reg_0031;
    74: op1_13_in11 = reg_1164;
    69: op1_13_in11 = reg_0128;
    54: op1_13_in11 = reg_0531;
    49: op1_13_in11 = imem07_in[3:0];
    75: op1_13_in11 = reg_0188;
    56: op1_13_in11 = reg_0606;
    50: op1_13_in11 = reg_0570;
    76: op1_13_in11 = reg_0398;
    71: op1_13_in11 = reg_0410;
    87: op1_13_in11 = reg_0411;
    68: op1_13_in11 = reg_1282;
    77: op1_13_in11 = reg_0475;
    61: op1_13_in11 = imem01_in[3:0];
    58: op1_13_in11 = reg_0120;
    78: op1_13_in11 = reg_1028;
    70: op1_13_in11 = reg_0891;
    59: op1_13_in11 = reg_0749;
    79: op1_13_in11 = reg_0459;
    51: op1_13_in11 = reg_0215;
    60: op1_13_in11 = reg_0341;
    88: op1_13_in11 = reg_1517;
    80: op1_13_in11 = reg_0879;
    62: op1_13_in11 = reg_0366;
    81: op1_13_in11 = reg_1215;
    63: op1_13_in11 = reg_0820;
    52: op1_13_in11 = reg_0419;
    82: op1_13_in11 = reg_0476;
    83: op1_13_in11 = reg_0584;
    64: op1_13_in11 = reg_0533;
    89: op1_13_in11 = reg_1367;
    84: op1_13_in11 = reg_1405;
    46: op1_13_in11 = reg_0251;
    85: op1_13_in11 = reg_0832;
    105: op1_13_in11 = reg_0832;
    65: op1_13_in11 = reg_0973;
    90: op1_13_in11 = reg_0196;
    66: op1_13_in11 = reg_0699;
    48: op1_13_in11 = reg_0524;
    91: op1_13_in11 = reg_0088;
    67: op1_13_in11 = reg_0530;
    92: op1_13_in11 = reg_0313;
    93: op1_13_in11 = reg_0840;
    94: op1_13_in11 = reg_0394;
    95: op1_13_in11 = reg_0136;
    96: op1_13_in11 = reg_1010;
    97: op1_13_in11 = reg_0026;
    98: op1_13_in11 = reg_1418;
    99: op1_13_in11 = reg_0425;
    100: op1_13_in11 = reg_0387;
    101: op1_13_in11 = reg_1488;
    102: op1_13_in11 = reg_0987;
    103: op1_13_in11 = reg_0472;
    104: op1_13_in11 = reg_0220;
    106: op1_13_in11 = reg_0924;
    107: op1_13_in11 = reg_0961;
    108: op1_13_in11 = imem05_in[7:4];
    109: op1_13_in11 = reg_1493;
    110: op1_13_in11 = reg_0622;
    111: op1_13_in11 = reg_0673;
    112: op1_13_in11 = reg_0141;
    113: op1_13_in11 = reg_0281;
    114: op1_13_in11 = reg_1321;
    115: op1_13_in11 = reg_0731;
    116: op1_13_in11 = reg_0203;
    117: op1_13_in11 = reg_0443;
    47: op1_13_in11 = reg_0729;
    118: op1_13_in11 = reg_1502;
    119: op1_13_in11 = reg_0870;
    120: op1_13_in11 = reg_0309;
    121: op1_13_in11 = reg_1432;
    122: op1_13_in11 = reg_1056;
    123: op1_13_in11 = reg_0045;
    124: op1_13_in11 = reg_0876;
    125: op1_13_in11 = reg_0171;
    126: op1_13_in11 = reg_0829;
    44: op1_13_in11 = reg_0129;
    127: op1_13_in11 = reg_0073;
    128: op1_13_in11 = reg_0005;
    129: op1_13_in11 = reg_0041;
    130: op1_13_in11 = reg_0221;
    default: op1_13_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv11 = 1;
    73: op1_13_inv11 = 1;
    86: op1_13_inv11 = 1;
    55: op1_13_inv11 = 1;
    74: op1_13_inv11 = 1;
    54: op1_13_inv11 = 1;
    49: op1_13_inv11 = 1;
    71: op1_13_inv11 = 1;
    77: op1_13_inv11 = 1;
    61: op1_13_inv11 = 1;
    78: op1_13_inv11 = 1;
    60: op1_13_inv11 = 1;
    88: op1_13_inv11 = 1;
    63: op1_13_inv11 = 1;
    52: op1_13_inv11 = 1;
    82: op1_13_inv11 = 1;
    83: op1_13_inv11 = 1;
    64: op1_13_inv11 = 1;
    84: op1_13_inv11 = 1;
    46: op1_13_inv11 = 1;
    85: op1_13_inv11 = 1;
    66: op1_13_inv11 = 1;
    92: op1_13_inv11 = 1;
    94: op1_13_inv11 = 1;
    103: op1_13_inv11 = 1;
    104: op1_13_inv11 = 1;
    107: op1_13_inv11 = 1;
    109: op1_13_inv11 = 1;
    110: op1_13_inv11 = 1;
    112: op1_13_inv11 = 1;
    116: op1_13_inv11 = 1;
    117: op1_13_inv11 = 1;
    119: op1_13_inv11 = 1;
    123: op1_13_inv11 = 1;
    124: op1_13_inv11 = 1;
    126: op1_13_inv11 = 1;
    127: op1_13_inv11 = 1;
    default: op1_13_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in12 = reg_1405;
    121: op1_13_in12 = reg_1405;
    53: op1_13_in12 = reg_0497;
    73: op1_13_in12 = reg_0152;
    86: op1_13_in12 = reg_0471;
    55: op1_13_in12 = reg_0030;
    74: op1_13_in12 = reg_0996;
    69: op1_13_in12 = reg_0126;
    54: op1_13_in12 = reg_0256;
    49: op1_13_in12 = reg_0139;
    75: op1_13_in12 = reg_0405;
    56: op1_13_in12 = reg_0253;
    50: op1_13_in12 = reg_0459;
    107: op1_13_in12 = reg_0459;
    76: op1_13_in12 = reg_0374;
    71: op1_13_in12 = reg_0060;
    87: op1_13_in12 = reg_1369;
    68: op1_13_in12 = reg_1280;
    77: op1_13_in12 = reg_0474;
    61: op1_13_in12 = reg_0695;
    58: op1_13_in12 = reg_0866;
    78: op1_13_in12 = reg_1459;
    70: op1_13_in12 = reg_0789;
    59: op1_13_in12 = reg_0737;
    79: op1_13_in12 = reg_1406;
    51: op1_13_in12 = reg_0394;
    60: op1_13_in12 = reg_0305;
    88: op1_13_in12 = reg_0954;
    80: op1_13_in12 = reg_0168;
    62: op1_13_in12 = reg_0740;
    81: op1_13_in12 = reg_1083;
    63: op1_13_in12 = reg_0976;
    52: op1_13_in12 = reg_0460;
    82: op1_13_in12 = reg_0886;
    83: op1_13_in12 = reg_0528;
    64: op1_13_in12 = reg_0455;
    67: op1_13_in12 = reg_0455;
    89: op1_13_in12 = reg_0535;
    84: op1_13_in12 = reg_0189;
    46: op1_13_in12 = reg_0118;
    85: op1_13_in12 = reg_1164;
    105: op1_13_in12 = reg_1164;
    65: op1_13_in12 = reg_0972;
    90: op1_13_in12 = reg_0130;
    66: op1_13_in12 = reg_0612;
    48: op1_13_in12 = reg_0619;
    91: op1_13_in12 = reg_1077;
    92: op1_13_in12 = reg_1139;
    93: op1_13_in12 = reg_0889;
    94: op1_13_in12 = reg_0498;
    95: op1_13_in12 = reg_0395;
    96: op1_13_in12 = reg_0298;
    97: op1_13_in12 = reg_1253;
    98: op1_13_in12 = reg_0524;
    99: op1_13_in12 = reg_0427;
    100: op1_13_in12 = reg_0058;
    127: op1_13_in12 = reg_0058;
    101: op1_13_in12 = reg_0470;
    102: op1_13_in12 = reg_0155;
    103: op1_13_in12 = reg_0054;
    104: op1_13_in12 = reg_0350;
    106: op1_13_in12 = reg_0779;
    108: op1_13_in12 = imem05_in[11:8];
    109: op1_13_in12 = reg_1074;
    110: op1_13_in12 = reg_0569;
    111: op1_13_in12 = reg_0443;
    112: op1_13_in12 = reg_0585;
    113: op1_13_in12 = reg_0412;
    114: op1_13_in12 = reg_0917;
    128: op1_13_in12 = reg_0917;
    115: op1_13_in12 = reg_0797;
    116: op1_13_in12 = reg_0057;
    117: op1_13_in12 = imem04_in[11:8];
    47: op1_13_in12 = imem06_in[3:0];
    118: op1_13_in12 = reg_0035;
    119: op1_13_in12 = reg_0782;
    120: op1_13_in12 = reg_0489;
    122: op1_13_in12 = reg_0703;
    123: op1_13_in12 = reg_0792;
    124: op1_13_in12 = reg_0306;
    125: op1_13_in12 = reg_0289;
    126: op1_13_in12 = reg_1098;
    44: op1_13_in12 = reg_0065;
    129: op1_13_in12 = reg_0012;
    130: op1_13_in12 = reg_0249;
    default: op1_13_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv12 = 1;
    73: op1_13_inv12 = 1;
    55: op1_13_inv12 = 1;
    74: op1_13_inv12 = 1;
    75: op1_13_inv12 = 1;
    56: op1_13_inv12 = 1;
    50: op1_13_inv12 = 1;
    71: op1_13_inv12 = 1;
    68: op1_13_inv12 = 1;
    77: op1_13_inv12 = 1;
    61: op1_13_inv12 = 1;
    58: op1_13_inv12 = 1;
    70: op1_13_inv12 = 1;
    79: op1_13_inv12 = 1;
    60: op1_13_inv12 = 1;
    80: op1_13_inv12 = 1;
    62: op1_13_inv12 = 1;
    52: op1_13_inv12 = 1;
    82: op1_13_inv12 = 1;
    84: op1_13_inv12 = 1;
    85: op1_13_inv12 = 1;
    65: op1_13_inv12 = 1;
    91: op1_13_inv12 = 1;
    93: op1_13_inv12 = 1;
    99: op1_13_inv12 = 1;
    100: op1_13_inv12 = 1;
    101: op1_13_inv12 = 1;
    102: op1_13_inv12 = 1;
    105: op1_13_inv12 = 1;
    106: op1_13_inv12 = 1;
    107: op1_13_inv12 = 1;
    111: op1_13_inv12 = 1;
    113: op1_13_inv12 = 1;
    114: op1_13_inv12 = 1;
    116: op1_13_inv12 = 1;
    119: op1_13_inv12 = 1;
    121: op1_13_inv12 = 1;
    122: op1_13_inv12 = 1;
    123: op1_13_inv12 = 1;
    126: op1_13_inv12 = 1;
    44: op1_13_inv12 = 1;
    129: op1_13_inv12 = 1;
    default: op1_13_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in13 = reg_0883;
    79: op1_13_in13 = reg_0883;
    53: op1_13_in13 = reg_0989;
    73: op1_13_in13 = reg_0215;
    86: op1_13_in13 = reg_0537;
    55: op1_13_in13 = reg_0286;
    74: op1_13_in13 = reg_0567;
    69: op1_13_in13 = reg_0138;
    54: op1_13_in13 = reg_0473;
    67: op1_13_in13 = reg_0473;
    49: op1_13_in13 = reg_0774;
    75: op1_13_in13 = reg_0387;
    56: op1_13_in13 = reg_0981;
    50: op1_13_in13 = reg_0023;
    76: op1_13_in13 = reg_0585;
    71: op1_13_in13 = reg_0072;
    87: op1_13_in13 = reg_0088;
    89: op1_13_in13 = reg_0088;
    68: op1_13_in13 = reg_0488;
    77: op1_13_in13 = reg_0054;
    61: op1_13_in13 = reg_0166;
    58: op1_13_in13 = reg_0827;
    78: op1_13_in13 = reg_1227;
    70: op1_13_in13 = reg_0963;
    59: op1_13_in13 = reg_1168;
    51: op1_13_in13 = reg_0191;
    60: op1_13_in13 = reg_0368;
    88: op1_13_in13 = reg_0597;
    80: op1_13_in13 = reg_0174;
    62: op1_13_in13 = reg_0738;
    81: op1_13_in13 = reg_1082;
    63: op1_13_in13 = reg_0530;
    52: op1_13_in13 = reg_0270;
    82: op1_13_in13 = reg_0722;
    83: op1_13_in13 = reg_0244;
    64: op1_13_in13 = reg_1018;
    84: op1_13_in13 = reg_0410;
    46: op1_13_in13 = reg_0272;
    85: op1_13_in13 = reg_0700;
    65: op1_13_in13 = reg_0106;
    90: op1_13_in13 = reg_0602;
    66: op1_13_in13 = reg_0606;
    48: op1_13_in13 = reg_0526;
    91: op1_13_in13 = reg_1419;
    92: op1_13_in13 = reg_0467;
    93: op1_13_in13 = reg_0759;
    94: op1_13_in13 = reg_1315;
    95: op1_13_in13 = reg_1164;
    96: op1_13_in13 = reg_0299;
    97: op1_13_in13 = reg_0609;
    98: op1_13_in13 = reg_0928;
    121: op1_13_in13 = reg_0928;
    99: op1_13_in13 = imem04_in[3:0];
    100: op1_13_in13 = reg_0057;
    101: op1_13_in13 = reg_0708;
    102: op1_13_in13 = reg_1406;
    103: op1_13_in13 = reg_0973;
    104: op1_13_in13 = reg_0291;
    105: op1_13_in13 = reg_0066;
    106: op1_13_in13 = reg_0287;
    107: op1_13_in13 = reg_0524;
    108: op1_13_in13 = reg_0831;
    109: op1_13_in13 = imem02_in[15:12];
    110: op1_13_in13 = reg_0345;
    111: op1_13_in13 = reg_1339;
    112: op1_13_in13 = reg_0569;
    113: op1_13_in13 = reg_0406;
    114: op1_13_in13 = reg_0277;
    115: op1_13_in13 = reg_0978;
    116: op1_13_in13 = reg_0027;
    117: op1_13_in13 = reg_0032;
    47: op1_13_in13 = imem06_in[15:12];
    118: op1_13_in13 = reg_1298;
    119: op1_13_in13 = reg_1437;
    120: op1_13_in13 = reg_0029;
    122: op1_13_in13 = reg_0851;
    123: op1_13_in13 = reg_0266;
    124: op1_13_in13 = reg_0829;
    125: op1_13_in13 = reg_1202;
    126: op1_13_in13 = reg_0711;
    44: op1_13_in13 = reg_0019;
    127: op1_13_in13 = reg_1324;
    128: op1_13_in13 = imem01_in[3:0];
    129: op1_13_in13 = reg_0895;
    130: op1_13_in13 = reg_1230;
    default: op1_13_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv13 = 1;
    73: op1_13_inv13 = 1;
    86: op1_13_inv13 = 1;
    55: op1_13_inv13 = 1;
    69: op1_13_inv13 = 1;
    75: op1_13_inv13 = 1;
    56: op1_13_inv13 = 1;
    76: op1_13_inv13 = 1;
    71: op1_13_inv13 = 1;
    87: op1_13_inv13 = 1;
    68: op1_13_inv13 = 1;
    77: op1_13_inv13 = 1;
    58: op1_13_inv13 = 1;
    59: op1_13_inv13 = 1;
    79: op1_13_inv13 = 1;
    51: op1_13_inv13 = 1;
    88: op1_13_inv13 = 1;
    82: op1_13_inv13 = 1;
    83: op1_13_inv13 = 1;
    64: op1_13_inv13 = 1;
    89: op1_13_inv13 = 1;
    84: op1_13_inv13 = 1;
    46: op1_13_inv13 = 1;
    85: op1_13_inv13 = 1;
    90: op1_13_inv13 = 1;
    48: op1_13_inv13 = 1;
    91: op1_13_inv13 = 1;
    94: op1_13_inv13 = 1;
    95: op1_13_inv13 = 1;
    96: op1_13_inv13 = 1;
    98: op1_13_inv13 = 1;
    99: op1_13_inv13 = 1;
    100: op1_13_inv13 = 1;
    102: op1_13_inv13 = 1;
    104: op1_13_inv13 = 1;
    106: op1_13_inv13 = 1;
    108: op1_13_inv13 = 1;
    109: op1_13_inv13 = 1;
    110: op1_13_inv13 = 1;
    111: op1_13_inv13 = 1;
    112: op1_13_inv13 = 1;
    118: op1_13_inv13 = 1;
    120: op1_13_inv13 = 1;
    121: op1_13_inv13 = 1;
    122: op1_13_inv13 = 1;
    124: op1_13_inv13 = 1;
    127: op1_13_inv13 = 1;
    128: op1_13_inv13 = 1;
    129: op1_13_inv13 = 1;
    default: op1_13_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in14 = reg_0202;
    79: op1_13_in14 = reg_0202;
    98: op1_13_in14 = reg_0202;
    53: op1_13_in14 = reg_0436;
    73: op1_13_in14 = reg_0015;
    86: op1_13_in14 = reg_0199;
    113: op1_13_in14 = reg_0199;
    55: op1_13_in14 = reg_0366;
    106: op1_13_in14 = reg_0366;
    74: op1_13_in14 = reg_0565;
    69: op1_13_in14 = reg_0848;
    54: op1_13_in14 = reg_0429;
    49: op1_13_in14 = reg_0031;
    75: op1_13_in14 = reg_1324;
    100: op1_13_in14 = reg_1324;
    56: op1_13_in14 = reg_0472;
    67: op1_13_in14 = reg_0472;
    50: op1_13_in14 = reg_0213;
    76: op1_13_in14 = reg_1228;
    71: op1_13_in14 = reg_0175;
    87: op1_13_in14 = reg_0264;
    68: op1_13_in14 = reg_0696;
    77: op1_13_in14 = reg_0105;
    61: op1_13_in14 = reg_0576;
    58: op1_13_in14 = reg_0716;
    78: op1_13_in14 = reg_1229;
    70: op1_13_in14 = reg_0964;
    59: op1_13_in14 = reg_1169;
    51: op1_13_in14 = reg_1057;
    60: op1_13_in14 = reg_0236;
    88: op1_13_in14 = reg_1300;
    80: op1_13_in14 = reg_0646;
    62: op1_13_in14 = reg_0415;
    81: op1_13_in14 = reg_0406;
    63: op1_13_in14 = reg_0169;
    52: op1_13_in14 = reg_0269;
    82: op1_13_in14 = reg_0440;
    83: op1_13_in14 = reg_1204;
    64: op1_13_in14 = reg_0233;
    89: op1_13_in14 = reg_0034;
    84: op1_13_in14 = reg_0089;
    46: op1_13_in14 = reg_0207;
    85: op1_13_in14 = reg_0176;
    95: op1_13_in14 = reg_0176;
    65: op1_13_in14 = reg_0382;
    90: op1_13_in14 = reg_0797;
    66: op1_13_in14 = reg_0608;
    48: op1_13_in14 = reg_0528;
    91: op1_13_in14 = reg_0369;
    92: op1_13_in14 = reg_0208;
    93: op1_13_in14 = reg_0154;
    94: op1_13_in14 = reg_0922;
    96: op1_13_in14 = reg_0309;
    97: op1_13_in14 = reg_0241;
    99: op1_13_in14 = imem04_in[7:4];
    101: op1_13_in14 = reg_0833;
    102: op1_13_in14 = reg_0887;
    103: op1_13_in14 = reg_0112;
    104: op1_13_in14 = reg_1139;
    105: op1_13_in14 = reg_0491;
    107: op1_13_in14 = reg_0821;
    108: op1_13_in14 = reg_0701;
    109: op1_13_in14 = reg_1207;
    110: op1_13_in14 = reg_0522;
    111: op1_13_in14 = reg_1144;
    112: op1_13_in14 = reg_0979;
    114: op1_13_in14 = reg_0446;
    115: op1_13_in14 = reg_0531;
    116: op1_13_in14 = reg_0267;
    117: op1_13_in14 = reg_1368;
    47: op1_13_in14 = reg_0907;
    118: op1_13_in14 = reg_0315;
    119: op1_13_in14 = reg_0271;
    120: op1_13_in14 = reg_0030;
    121: op1_13_in14 = reg_0927;
    122: op1_13_in14 = reg_0457;
    123: op1_13_in14 = reg_1163;
    124: op1_13_in14 = reg_0897;
    125: op1_13_in14 = reg_0754;
    126: op1_13_in14 = reg_0294;
    44: op1_13_in14 = reg_0033;
    127: op1_13_in14 = reg_0026;
    128: op1_13_in14 = reg_0985;
    129: op1_13_in14 = reg_0662;
    130: op1_13_in14 = reg_1405;
    default: op1_13_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv14 = 1;
    73: op1_13_inv14 = 1;
    86: op1_13_inv14 = 1;
    49: op1_13_inv14 = 1;
    50: op1_13_inv14 = 1;
    71: op1_13_inv14 = 1;
    87: op1_13_inv14 = 1;
    70: op1_13_inv14 = 1;
    59: op1_13_inv14 = 1;
    51: op1_13_inv14 = 1;
    60: op1_13_inv14 = 1;
    88: op1_13_inv14 = 1;
    80: op1_13_inv14 = 1;
    62: op1_13_inv14 = 1;
    81: op1_13_inv14 = 1;
    82: op1_13_inv14 = 1;
    83: op1_13_inv14 = 1;
    89: op1_13_inv14 = 1;
    84: op1_13_inv14 = 1;
    46: op1_13_inv14 = 1;
    65: op1_13_inv14 = 1;
    90: op1_13_inv14 = 1;
    91: op1_13_inv14 = 1;
    67: op1_13_inv14 = 1;
    92: op1_13_inv14 = 1;
    94: op1_13_inv14 = 1;
    96: op1_13_inv14 = 1;
    97: op1_13_inv14 = 1;
    98: op1_13_inv14 = 1;
    100: op1_13_inv14 = 1;
    102: op1_13_inv14 = 1;
    107: op1_13_inv14 = 1;
    110: op1_13_inv14 = 1;
    111: op1_13_inv14 = 1;
    115: op1_13_inv14 = 1;
    47: op1_13_inv14 = 1;
    120: op1_13_inv14 = 1;
    122: op1_13_inv14 = 1;
    123: op1_13_inv14 = 1;
    127: op1_13_inv14 = 1;
    129: op1_13_inv14 = 1;
    130: op1_13_inv14 = 1;
    default: op1_13_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in15 = reg_0428;
    53: op1_13_in15 = reg_0054;
    73: op1_13_in15 = imem07_in[3:0];
    86: op1_13_in15 = reg_1004;
    55: op1_13_in15 = reg_0413;
    74: op1_13_in15 = reg_0334;
    69: op1_13_in15 = reg_0845;
    54: op1_13_in15 = reg_0127;
    49: op1_13_in15 = reg_0465;
    75: op1_13_in15 = reg_0122;
    56: op1_13_in15 = reg_1207;
    50: op1_13_in15 = reg_0457;
    76: op1_13_in15 = reg_0171;
    71: op1_13_in15 = reg_0553;
    87: op1_13_in15 = reg_1338;
    68: op1_13_in15 = reg_1372;
    111: op1_13_in15 = reg_1372;
    77: op1_13_in15 = reg_1433;
    61: op1_13_in15 = reg_0575;
    58: op1_13_in15 = reg_0637;
    78: op1_13_in15 = reg_1201;
    70: op1_13_in15 = reg_0627;
    59: op1_13_in15 = reg_0996;
    79: op1_13_in15 = reg_0353;
    51: op1_13_in15 = reg_1060;
    60: op1_13_in15 = reg_0799;
    88: op1_13_in15 = reg_1199;
    80: op1_13_in15 = reg_0649;
    62: op1_13_in15 = reg_0618;
    81: op1_13_in15 = reg_0471;
    63: op1_13_in15 = reg_0497;
    52: op1_13_in15 = reg_0067;
    82: op1_13_in15 = reg_0071;
    83: op1_13_in15 = reg_0215;
    64: op1_13_in15 = reg_0778;
    89: op1_13_in15 = reg_0531;
    84: op1_13_in15 = reg_0723;
    116: op1_13_in15 = reg_0723;
    46: op1_13_in15 = reg_0037;
    85: op1_13_in15 = reg_0648;
    65: op1_13_in15 = reg_0055;
    90: op1_13_in15 = reg_0449;
    66: op1_13_in15 = reg_0532;
    48: op1_13_in15 = reg_0529;
    91: op1_13_in15 = reg_0340;
    67: op1_13_in15 = reg_0436;
    92: op1_13_in15 = reg_0696;
    93: op1_13_in15 = reg_0573;
    94: op1_13_in15 = reg_0135;
    95: op1_13_in15 = reg_1403;
    96: op1_13_in15 = reg_1350;
    97: op1_13_in15 = reg_1457;
    98: op1_13_in15 = reg_0352;
    99: op1_13_in15 = reg_0263;
    100: op1_13_in15 = reg_1031;
    101: op1_13_in15 = reg_0466;
    102: op1_13_in15 = reg_0202;
    107: op1_13_in15 = reg_0202;
    103: op1_13_in15 = reg_0684;
    104: op1_13_in15 = reg_0790;
    105: op1_13_in15 = reg_1181;
    106: op1_13_in15 = reg_0739;
    108: op1_13_in15 = reg_0566;
    109: op1_13_in15 = reg_1451;
    110: op1_13_in15 = reg_0295;
    112: op1_13_in15 = reg_0119;
    113: op1_13_in15 = reg_0097;
    114: op1_13_in15 = reg_0874;
    115: op1_13_in15 = reg_0574;
    117: op1_13_in15 = reg_1367;
    47: op1_13_in15 = reg_0905;
    118: op1_13_in15 = reg_0538;
    119: op1_13_in15 = reg_1467;
    120: op1_13_in15 = reg_0661;
    121: op1_13_in15 = reg_0883;
    130: op1_13_in15 = reg_0883;
    122: op1_13_in15 = reg_0139;
    123: op1_13_in15 = reg_0477;
    124: op1_13_in15 = reg_0632;
    125: op1_13_in15 = reg_0977;
    126: op1_13_in15 = reg_0007;
    44: op1_13_in15 = reg_0392;
    127: op1_13_in15 = reg_0383;
    128: op1_13_in15 = reg_0013;
    129: op1_13_in15 = reg_0056;
    default: op1_13_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv15 = 1;
    73: op1_13_inv15 = 1;
    69: op1_13_inv15 = 1;
    54: op1_13_inv15 = 1;
    49: op1_13_inv15 = 1;
    68: op1_13_inv15 = 1;
    61: op1_13_inv15 = 1;
    58: op1_13_inv15 = 1;
    78: op1_13_inv15 = 1;
    51: op1_13_inv15 = 1;
    63: op1_13_inv15 = 1;
    52: op1_13_inv15 = 1;
    64: op1_13_inv15 = 1;
    85: op1_13_inv15 = 1;
    65: op1_13_inv15 = 1;
    48: op1_13_inv15 = 1;
    91: op1_13_inv15 = 1;
    92: op1_13_inv15 = 1;
    93: op1_13_inv15 = 1;
    94: op1_13_inv15 = 1;
    95: op1_13_inv15 = 1;
    96: op1_13_inv15 = 1;
    98: op1_13_inv15 = 1;
    99: op1_13_inv15 = 1;
    102: op1_13_inv15 = 1;
    103: op1_13_inv15 = 1;
    104: op1_13_inv15 = 1;
    107: op1_13_inv15 = 1;
    108: op1_13_inv15 = 1;
    109: op1_13_inv15 = 1;
    110: op1_13_inv15 = 1;
    111: op1_13_inv15 = 1;
    112: op1_13_inv15 = 1;
    114: op1_13_inv15 = 1;
    116: op1_13_inv15 = 1;
    47: op1_13_inv15 = 1;
    122: op1_13_inv15 = 1;
    123: op1_13_inv15 = 1;
    124: op1_13_inv15 = 1;
    125: op1_13_inv15 = 1;
    44: op1_13_inv15 = 1;
    129: op1_13_inv15 = 1;
    default: op1_13_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in16 = reg_0440;
    53: op1_13_in16 = reg_0776;
    73: op1_13_in16 = reg_0065;
    86: op1_13_in16 = reg_0262;
    55: op1_13_in16 = reg_0621;
    74: op1_13_in16 = reg_1181;
    69: op1_13_in16 = reg_0846;
    54: op1_13_in16 = reg_0105;
    49: op1_13_in16 = reg_0741;
    75: op1_13_in16 = reg_0917;
    56: op1_13_in16 = reg_0934;
    50: op1_13_in16 = reg_0230;
    76: op1_13_in16 = reg_1204;
    71: op1_13_in16 = reg_0259;
    61: op1_13_in16 = reg_0259;
    87: op1_13_in16 = reg_0978;
    68: op1_13_in16 = reg_1369;
    77: op1_13_in16 = reg_0839;
    58: op1_13_in16 = imem06_in[15:12];
    78: op1_13_in16 = reg_0961;
    70: op1_13_in16 = reg_0048;
    124: op1_13_in16 = reg_0048;
    59: op1_13_in16 = reg_0346;
    79: op1_13_in16 = reg_0201;
    51: op1_13_in16 = reg_0993;
    60: op1_13_in16 = reg_0332;
    88: op1_13_in16 = reg_0178;
    80: op1_13_in16 = imem05_in[11:8];
    62: op1_13_in16 = reg_0620;
    81: op1_13_in16 = reg_0837;
    63: op1_13_in16 = reg_0981;
    52: op1_13_in16 = imem07_in[7:4];
    82: op1_13_in16 = reg_0963;
    83: op1_13_in16 = reg_0214;
    64: op1_13_in16 = reg_0973;
    89: op1_13_in16 = reg_0552;
    84: op1_13_in16 = reg_1100;
    46: op1_13_in16 = reg_0040;
    85: op1_13_in16 = reg_0391;
    65: op1_13_in16 = reg_0294;
    90: op1_13_in16 = reg_0207;
    66: op1_13_in16 = reg_0588;
    48: op1_13_in16 = reg_0527;
    91: op1_13_in16 = reg_0304;
    67: op1_13_in16 = reg_0054;
    92: op1_13_in16 = reg_0264;
    93: op1_13_in16 = reg_0600;
    94: op1_13_in16 = reg_0225;
    95: op1_13_in16 = reg_1401;
    96: op1_13_in16 = reg_0924;
    97: op1_13_in16 = reg_0091;
    98: op1_13_in16 = reg_0435;
    99: op1_13_in16 = reg_1372;
    100: op1_13_in16 = reg_0355;
    101: op1_13_in16 = reg_0278;
    102: op1_13_in16 = reg_0188;
    103: op1_13_in16 = reg_0631;
    104: op1_13_in16 = reg_0427;
    105: op1_13_in16 = reg_0697;
    108: op1_13_in16 = reg_0697;
    106: op1_13_in16 = reg_0137;
    107: op1_13_in16 = reg_0058;
    109: op1_13_in16 = reg_0126;
    110: op1_13_in16 = reg_0583;
    111: op1_13_in16 = imem04_in[3:0];
    112: op1_13_in16 = imem07_in[11:8];
    113: op1_13_in16 = reg_0698;
    114: op1_13_in16 = reg_0930;
    115: op1_13_in16 = reg_1215;
    116: op1_13_in16 = imem01_in[7:4];
    117: op1_13_in16 = reg_0493;
    47: op1_13_in16 = reg_0730;
    118: op1_13_in16 = reg_0579;
    119: op1_13_in16 = reg_0752;
    120: op1_13_in16 = reg_0663;
    121: op1_13_in16 = reg_0431;
    122: op1_13_in16 = reg_0031;
    123: op1_13_in16 = reg_0090;
    125: op1_13_in16 = reg_0023;
    126: op1_13_in16 = reg_1006;
    44: op1_13_in16 = reg_0745;
    127: op1_13_in16 = reg_0183;
    128: op1_13_in16 = reg_0463;
    129: op1_13_in16 = reg_0608;
    130: op1_13_in16 = reg_0886;
    default: op1_13_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv16 = 1;
    86: op1_13_inv16 = 1;
    69: op1_13_inv16 = 1;
    49: op1_13_inv16 = 1;
    75: op1_13_inv16 = 1;
    56: op1_13_inv16 = 1;
    71: op1_13_inv16 = 1;
    68: op1_13_inv16 = 1;
    77: op1_13_inv16 = 1;
    58: op1_13_inv16 = 1;
    78: op1_13_inv16 = 1;
    70: op1_13_inv16 = 1;
    79: op1_13_inv16 = 1;
    80: op1_13_inv16 = 1;
    63: op1_13_inv16 = 1;
    52: op1_13_inv16 = 1;
    82: op1_13_inv16 = 1;
    83: op1_13_inv16 = 1;
    90: op1_13_inv16 = 1;
    48: op1_13_inv16 = 1;
    91: op1_13_inv16 = 1;
    94: op1_13_inv16 = 1;
    95: op1_13_inv16 = 1;
    97: op1_13_inv16 = 1;
    98: op1_13_inv16 = 1;
    99: op1_13_inv16 = 1;
    101: op1_13_inv16 = 1;
    105: op1_13_inv16 = 1;
    106: op1_13_inv16 = 1;
    108: op1_13_inv16 = 1;
    109: op1_13_inv16 = 1;
    110: op1_13_inv16 = 1;
    112: op1_13_inv16 = 1;
    115: op1_13_inv16 = 1;
    121: op1_13_inv16 = 1;
    122: op1_13_inv16 = 1;
    124: op1_13_inv16 = 1;
    125: op1_13_inv16 = 1;
    126: op1_13_inv16 = 1;
    44: op1_13_inv16 = 1;
    130: op1_13_inv16 = 1;
    default: op1_13_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in17 = reg_0134;
    53: op1_13_in17 = reg_0326;
    73: op1_13_in17 = reg_1441;
    86: op1_13_in17 = reg_0836;
    55: op1_13_in17 = reg_0114;
    120: op1_13_in17 = reg_0114;
    74: op1_13_in17 = reg_1401;
    69: op1_13_in17 = reg_0024;
    54: op1_13_in17 = reg_0876;
    65: op1_13_in17 = reg_0876;
    49: op1_13_in17 = reg_0103;
    75: op1_13_in17 = reg_0822;
    56: op1_13_in17 = reg_0106;
    50: op1_13_in17 = reg_0135;
    76: op1_13_in17 = reg_1179;
    119: op1_13_in17 = reg_1179;
    71: op1_13_in17 = reg_0548;
    87: op1_13_in17 = reg_1083;
    68: op1_13_in17 = reg_0252;
    77: op1_13_in17 = reg_0708;
    61: op1_13_in17 = reg_0258;
    58: op1_13_in17 = reg_0622;
    78: op1_13_in17 = reg_1417;
    70: op1_13_in17 = reg_1093;
    59: op1_13_in17 = reg_0392;
    79: op1_13_in17 = reg_0428;
    51: op1_13_in17 = reg_0704;
    60: op1_13_in17 = reg_0736;
    88: op1_13_in17 = reg_0480;
    80: op1_13_in17 = imem05_in[15:12];
    62: op1_13_in17 = reg_0050;
    81: op1_13_in17 = reg_0719;
    63: op1_13_in17 = reg_0256;
    66: op1_13_in17 = reg_0256;
    52: op1_13_in17 = imem07_in[11:8];
    82: op1_13_in17 = reg_0553;
    83: op1_13_in17 = reg_1170;
    64: op1_13_in17 = reg_0128;
    89: op1_13_in17 = reg_1214;
    117: op1_13_in17 = reg_1214;
    84: op1_13_in17 = reg_0335;
    46: op1_13_in17 = reg_0752;
    85: op1_13_in17 = reg_0566;
    90: op1_13_in17 = reg_0206;
    48: op1_13_in17 = reg_0295;
    91: op1_13_in17 = reg_0305;
    67: op1_13_in17 = reg_0971;
    92: op1_13_in17 = reg_1203;
    93: op1_13_in17 = reg_0312;
    94: op1_13_in17 = reg_0309;
    95: op1_13_in17 = reg_0794;
    123: op1_13_in17 = reg_0794;
    96: op1_13_in17 = reg_0923;
    97: op1_13_in17 = reg_0724;
    98: op1_13_in17 = reg_0416;
    99: op1_13_in17 = reg_0181;
    100: op1_13_in17 = reg_0550;
    114: op1_13_in17 = reg_0550;
    101: op1_13_in17 = reg_0251;
    102: op1_13_in17 = reg_0201;
    103: op1_13_in17 = reg_0379;
    104: op1_13_in17 = imem04_in[7:4];
    105: op1_13_in17 = reg_0940;
    106: op1_13_in17 = reg_0102;
    107: op1_13_in17 = reg_0027;
    108: op1_13_in17 = reg_1404;
    109: op1_13_in17 = reg_0382;
    110: op1_13_in17 = reg_0213;
    111: op1_13_in17 = reg_1082;
    112: op1_13_in17 = reg_1097;
    113: op1_13_in17 = reg_0420;
    115: op1_13_in17 = reg_0500;
    116: op1_13_in17 = imem01_in[11:8];
    47: op1_13_in17 = reg_0396;
    118: op1_13_in17 = reg_0833;
    44: op1_13_in17 = reg_0833;
    121: op1_13_in17 = reg_0435;
    122: op1_13_in17 = reg_0665;
    124: op1_13_in17 = reg_0444;
    125: op1_13_in17 = reg_0215;
    126: op1_13_in17 = reg_0217;
    127: op1_13_in17 = reg_0577;
    128: op1_13_in17 = reg_0549;
    129: op1_13_in17 = reg_0934;
    130: op1_13_in17 = reg_0202;
    default: op1_13_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    49: op1_13_inv17 = 1;
    75: op1_13_inv17 = 1;
    56: op1_13_inv17 = 1;
    71: op1_13_inv17 = 1;
    68: op1_13_inv17 = 1;
    58: op1_13_inv17 = 1;
    78: op1_13_inv17 = 1;
    70: op1_13_inv17 = 1;
    88: op1_13_inv17 = 1;
    62: op1_13_inv17 = 1;
    81: op1_13_inv17 = 1;
    52: op1_13_inv17 = 1;
    84: op1_13_inv17 = 1;
    85: op1_13_inv17 = 1;
    90: op1_13_inv17 = 1;
    66: op1_13_inv17 = 1;
    67: op1_13_inv17 = 1;
    93: op1_13_inv17 = 1;
    107: op1_13_inv17 = 1;
    108: op1_13_inv17 = 1;
    112: op1_13_inv17 = 1;
    113: op1_13_inv17 = 1;
    114: op1_13_inv17 = 1;
    116: op1_13_inv17 = 1;
    121: op1_13_inv17 = 1;
    122: op1_13_inv17 = 1;
    123: op1_13_inv17 = 1;
    124: op1_13_inv17 = 1;
    126: op1_13_inv17 = 1;
    44: op1_13_inv17 = 1;
    127: op1_13_inv17 = 1;
    130: op1_13_inv17 = 1;
    default: op1_13_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in18 = reg_0203;
    79: op1_13_in18 = reg_0203;
    53: op1_13_in18 = reg_0379;
    73: op1_13_in18 = reg_1439;
    86: op1_13_in18 = reg_0338;
    55: op1_13_in18 = reg_0051;
    62: op1_13_in18 = reg_0051;
    74: op1_13_in18 = imem05_in[7:4];
    69: op1_13_in18 = reg_0757;
    54: op1_13_in18 = reg_0848;
    77: op1_13_in18 = reg_0848;
    49: op1_13_in18 = reg_0228;
    75: op1_13_in18 = reg_0785;
    56: op1_13_in18 = reg_0105;
    50: op1_13_in18 = reg_0490;
    76: op1_13_in18 = reg_0067;
    71: op1_13_in18 = reg_0610;
    87: op1_13_in18 = reg_1233;
    68: op1_13_in18 = reg_0462;
    61: op1_13_in18 = reg_0241;
    58: op1_13_in18 = reg_0526;
    78: op1_13_in18 = reg_0524;
    70: op1_13_in18 = reg_1226;
    59: op1_13_in18 = reg_0174;
    44: op1_13_in18 = reg_0174;
    51: op1_13_in18 = reg_0867;
    60: op1_13_in18 = reg_0737;
    88: op1_13_in18 = reg_0288;
    80: op1_13_in18 = reg_0697;
    81: op1_13_in18 = reg_0835;
    63: op1_13_in18 = reg_0475;
    52: op1_13_in18 = reg_1055;
    82: op1_13_in18 = reg_0163;
    83: op1_13_in18 = imem07_in[11:8];
    64: op1_13_in18 = reg_0380;
    89: op1_13_in18 = reg_1147;
    84: op1_13_in18 = reg_1256;
    46: op1_13_in18 = reg_0193;
    85: op1_13_in18 = reg_0131;
    65: op1_13_in18 = reg_0755;
    90: op1_13_in18 = reg_0753;
    66: op1_13_in18 = reg_1260;
    48: op1_13_in18 = reg_0171;
    91: op1_13_in18 = reg_0836;
    67: op1_13_in18 = reg_0972;
    92: op1_13_in18 = reg_0796;
    93: op1_13_in18 = reg_1517;
    94: op1_13_in18 = reg_0851;
    95: op1_13_in18 = reg_0450;
    96: op1_13_in18 = reg_1094;
    97: op1_13_in18 = reg_0042;
    98: op1_13_in18 = reg_0057;
    99: op1_13_in18 = reg_1369;
    100: op1_13_in18 = reg_0746;
    101: op1_13_in18 = reg_0491;
    102: op1_13_in18 = reg_0134;
    103: op1_13_in18 = reg_1392;
    104: op1_13_in18 = reg_0032;
    105: op1_13_in18 = reg_0937;
    106: op1_13_in18 = reg_0050;
    107: op1_13_in18 = imem01_in[11:8];
    108: op1_13_in18 = reg_1514;
    109: op1_13_in18 = reg_1492;
    110: op1_13_in18 = reg_0017;
    111: op1_13_in18 = reg_0414;
    112: op1_13_in18 = reg_1096;
    113: op1_13_in18 = reg_1502;
    114: op1_13_in18 = reg_0747;
    115: op1_13_in18 = reg_1082;
    116: op1_13_in18 = reg_0982;
    117: op1_13_in18 = reg_0421;
    47: op1_13_in18 = reg_0826;
    118: op1_13_in18 = reg_0278;
    119: op1_13_in18 = reg_0115;
    120: op1_13_in18 = reg_0361;
    121: op1_13_in18 = reg_0416;
    122: op1_13_in18 = reg_0442;
    123: op1_13_in18 = reg_0151;
    124: op1_13_in18 = reg_0507;
    125: op1_13_in18 = reg_0213;
    126: op1_13_in18 = reg_0009;
    127: op1_13_in18 = reg_1152;
    128: op1_13_in18 = reg_0609;
    129: op1_13_in18 = reg_0055;
    130: op1_13_in18 = reg_0351;
    default: op1_13_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv18 = 1;
    73: op1_13_inv18 = 1;
    86: op1_13_inv18 = 1;
    55: op1_13_inv18 = 1;
    54: op1_13_inv18 = 1;
    75: op1_13_inv18 = 1;
    56: op1_13_inv18 = 1;
    50: op1_13_inv18 = 1;
    71: op1_13_inv18 = 1;
    87: op1_13_inv18 = 1;
    68: op1_13_inv18 = 1;
    58: op1_13_inv18 = 1;
    78: op1_13_inv18 = 1;
    59: op1_13_inv18 = 1;
    88: op1_13_inv18 = 1;
    81: op1_13_inv18 = 1;
    63: op1_13_inv18 = 1;
    64: op1_13_inv18 = 1;
    46: op1_13_inv18 = 1;
    66: op1_13_inv18 = 1;
    94: op1_13_inv18 = 1;
    95: op1_13_inv18 = 1;
    96: op1_13_inv18 = 1;
    98: op1_13_inv18 = 1;
    100: op1_13_inv18 = 1;
    107: op1_13_inv18 = 1;
    109: op1_13_inv18 = 1;
    110: op1_13_inv18 = 1;
    112: op1_13_inv18 = 1;
    113: op1_13_inv18 = 1;
    114: op1_13_inv18 = 1;
    116: op1_13_inv18 = 1;
    47: op1_13_inv18 = 1;
    118: op1_13_inv18 = 1;
    119: op1_13_inv18 = 1;
    121: op1_13_inv18 = 1;
    123: op1_13_inv18 = 1;
    124: op1_13_inv18 = 1;
    44: op1_13_inv18 = 1;
    127: op1_13_inv18 = 1;
    130: op1_13_inv18 = 1;
    default: op1_13_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in19 = reg_0060;
    53: op1_13_in19 = reg_0897;
    73: op1_13_in19 = reg_1416;
    86: op1_13_in19 = reg_1237;
    55: op1_13_in19 = reg_0003;
    49: op1_13_in19 = reg_0003;
    74: op1_13_in19 = reg_0090;
    69: op1_13_in19 = reg_0755;
    54: op1_13_in19 = reg_0846;
    75: op1_13_in19 = reg_0335;
    56: op1_13_in19 = reg_0379;
    50: op1_13_in19 = reg_0491;
    76: op1_13_in19 = reg_0046;
    71: op1_13_in19 = reg_0149;
    87: op1_13_in19 = reg_0500;
    68: op1_13_in19 = reg_0574;
    77: op1_13_in19 = reg_0008;
    61: op1_13_in19 = reg_1152;
    58: op1_13_in19 = reg_0568;
    78: op1_13_in19 = reg_0886;
    70: op1_13_in19 = reg_0107;
    59: op1_13_in19 = reg_0045;
    79: op1_13_in19 = reg_0072;
    51: op1_13_in19 = reg_0673;
    60: op1_13_in19 = reg_0700;
    88: op1_13_in19 = imem04_in[11:8];
    80: op1_13_in19 = reg_1070;
    62: op1_13_in19 = reg_0052;
    81: op1_13_in19 = reg_0336;
    63: op1_13_in19 = reg_0433;
    52: op1_13_in19 = reg_1056;
    82: op1_13_in19 = reg_0547;
    83: op1_13_in19 = imem07_in[15:12];
    64: op1_13_in19 = reg_0900;
    89: op1_13_in19 = reg_0033;
    84: op1_13_in19 = reg_0742;
    46: op1_13_in19 = reg_0160;
    85: op1_13_in19 = reg_0938;
    65: op1_13_in19 = reg_0732;
    90: op1_13_in19 = reg_0195;
    66: op1_13_in19 = reg_0631;
    48: op1_13_in19 = reg_0023;
    91: op1_13_in19 = reg_1189;
    67: op1_13_in19 = reg_0106;
    92: op1_13_in19 = reg_0421;
    93: op1_13_in19 = reg_0314;
    94: op1_13_in19 = reg_1350;
    95: op1_13_in19 = reg_0477;
    96: op1_13_in19 = reg_0779;
    97: op1_13_in19 = reg_1068;
    98: op1_13_in19 = reg_0026;
    99: op1_13_in19 = reg_0264;
    100: op1_13_in19 = reg_0612;
    101: op1_13_in19 = reg_0131;
    102: op1_13_in19 = reg_1321;
    103: op1_13_in19 = reg_1006;
    104: op1_13_in19 = reg_0263;
    105: op1_13_in19 = reg_0418;
    106: op1_13_in19 = reg_0002;
    107: op1_13_in19 = reg_0788;
    108: op1_13_in19 = reg_0301;
    109: op1_13_in19 = reg_0024;
    110: op1_13_in19 = reg_1170;
    111: op1_13_in19 = reg_1419;
    112: op1_13_in19 = reg_0963;
    113: op1_13_in19 = reg_0021;
    114: op1_13_in19 = reg_0239;
    115: op1_13_in19 = reg_0796;
    116: op1_13_in19 = reg_0549;
    117: op1_13_in19 = reg_0406;
    47: op1_13_in19 = reg_0110;
    118: op1_13_in19 = reg_0333;
    119: op1_13_in19 = reg_0116;
    120: op1_13_in19 = reg_0226;
    121: op1_13_in19 = reg_0405;
    122: op1_13_in19 = reg_0593;
    123: op1_13_in19 = reg_0207;
    124: op1_13_in19 = reg_1033;
    125: op1_13_in19 = reg_0017;
    126: op1_13_in19 = reg_0006;
    44: op1_13_in19 = reg_0445;
    127: op1_13_in19 = reg_0078;
    128: op1_13_in19 = reg_0242;
    129: op1_13_in19 = reg_0898;
    130: op1_13_in19 = reg_0188;
    default: op1_13_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv19 = 1;
    73: op1_13_inv19 = 1;
    55: op1_13_inv19 = 1;
    49: op1_13_inv19 = 1;
    50: op1_13_inv19 = 1;
    76: op1_13_inv19 = 1;
    71: op1_13_inv19 = 1;
    87: op1_13_inv19 = 1;
    68: op1_13_inv19 = 1;
    77: op1_13_inv19 = 1;
    78: op1_13_inv19 = 1;
    59: op1_13_inv19 = 1;
    60: op1_13_inv19 = 1;
    80: op1_13_inv19 = 1;
    63: op1_13_inv19 = 1;
    52: op1_13_inv19 = 1;
    84: op1_13_inv19 = 1;
    46: op1_13_inv19 = 1;
    65: op1_13_inv19 = 1;
    90: op1_13_inv19 = 1;
    66: op1_13_inv19 = 1;
    48: op1_13_inv19 = 1;
    91: op1_13_inv19 = 1;
    67: op1_13_inv19 = 1;
    92: op1_13_inv19 = 1;
    94: op1_13_inv19 = 1;
    96: op1_13_inv19 = 1;
    98: op1_13_inv19 = 1;
    99: op1_13_inv19 = 1;
    100: op1_13_inv19 = 1;
    102: op1_13_inv19 = 1;
    104: op1_13_inv19 = 1;
    105: op1_13_inv19 = 1;
    106: op1_13_inv19 = 1;
    108: op1_13_inv19 = 1;
    109: op1_13_inv19 = 1;
    111: op1_13_inv19 = 1;
    113: op1_13_inv19 = 1;
    114: op1_13_inv19 = 1;
    117: op1_13_inv19 = 1;
    47: op1_13_inv19 = 1;
    119: op1_13_inv19 = 1;
    120: op1_13_inv19 = 1;
    121: op1_13_inv19 = 1;
    126: op1_13_inv19 = 1;
    44: op1_13_inv19 = 1;
    127: op1_13_inv19 = 1;
    128: op1_13_inv19 = 1;
    default: op1_13_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in20 = reg_0057;
    53: op1_13_in20 = reg_0900;
    73: op1_13_in20 = reg_0025;
    86: op1_13_in20 = reg_0904;
    55: op1_13_in20 = reg_0086;
    74: op1_13_in20 = reg_0873;
    69: op1_13_in20 = reg_0675;
    54: op1_13_in20 = reg_0007;
    49: op1_13_in20 = reg_0001;
    75: op1_13_in20 = reg_0175;
    56: op1_13_in20 = reg_0380;
    50: op1_13_in20 = imem07_in[11:8];
    76: op1_13_in20 = reg_0962;
    71: op1_13_in20 = reg_0896;
    87: op1_13_in20 = reg_0471;
    68: op1_13_in20 = reg_1065;
    77: op1_13_in20 = reg_0006;
    109: op1_13_in20 = reg_0006;
    61: op1_13_in20 = reg_0982;
    58: op1_13_in20 = reg_0571;
    78: op1_13_in20 = reg_0351;
    70: op1_13_in20 = reg_0504;
    59: op1_13_in20 = reg_0538;
    79: op1_13_in20 = reg_1321;
    51: op1_13_in20 = reg_0779;
    60: op1_13_in20 = reg_0649;
    88: op1_13_in20 = reg_0341;
    80: op1_13_in20 = reg_0937;
    95: op1_13_in20 = reg_0937;
    62: op1_13_in20 = reg_0084;
    81: op1_13_in20 = reg_1503;
    63: op1_13_in20 = reg_0326;
    52: op1_13_in20 = reg_0159;
    82: op1_13_in20 = reg_0612;
    83: op1_13_in20 = reg_0187;
    64: op1_13_in20 = reg_0705;
    89: op1_13_in20 = reg_1419;
    84: op1_13_in20 = reg_1456;
    46: op1_13_in20 = reg_0906;
    85: op1_13_in20 = reg_0450;
    65: op1_13_in20 = reg_0525;
    90: op1_13_in20 = reg_1058;
    66: op1_13_in20 = reg_0475;
    48: op1_13_in20 = reg_0152;
    91: op1_13_in20 = reg_0211;
    67: op1_13_in20 = reg_0056;
    92: op1_13_in20 = reg_0414;
    93: op1_13_in20 = reg_0954;
    94: op1_13_in20 = reg_1347;
    96: op1_13_in20 = reg_0775;
    97: op1_13_in20 = reg_0934;
    98: op1_13_in20 = reg_1152;
    99: op1_13_in20 = reg_0164;
    100: op1_13_in20 = reg_0438;
    101: op1_13_in20 = reg_0938;
    102: op1_13_in20 = reg_1322;
    103: op1_13_in20 = reg_0217;
    104: op1_13_in20 = reg_1372;
    105: op1_13_in20 = reg_0302;
    106: op1_13_in20 = reg_0085;
    107: op1_13_in20 = reg_0446;
    108: op1_13_in20 = reg_0575;
    110: op1_13_in20 = imem07_in[15:12];
    111: op1_13_in20 = reg_0862;
    112: op1_13_in20 = reg_0324;
    113: op1_13_in20 = reg_0035;
    114: op1_13_in20 = reg_0715;
    115: op1_13_in20 = reg_0598;
    116: op1_13_in20 = reg_0819;
    117: op1_13_in20 = reg_0969;
    47: op1_13_in20 = reg_0585;
    118: op1_13_in20 = reg_0733;
    119: op1_13_in20 = reg_0714;
    121: op1_13_in20 = reg_0134;
    122: op1_13_in20 = reg_1351;
    123: op1_13_in20 = reg_1431;
    124: op1_13_in20 = reg_0312;
    125: op1_13_in20 = reg_0034;
    126: op1_13_in20 = reg_0952;
    44: op1_13_in20 = reg_0603;
    127: op1_13_in20 = reg_0163;
    128: op1_13_in20 = reg_0241;
    129: op1_13_in20 = reg_0778;
    130: op1_13_in20 = reg_0410;
    default: op1_13_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_13_inv20 = 1;
    55: op1_13_inv20 = 1;
    69: op1_13_inv20 = 1;
    49: op1_13_inv20 = 1;
    75: op1_13_inv20 = 1;
    68: op1_13_inv20 = 1;
    77: op1_13_inv20 = 1;
    61: op1_13_inv20 = 1;
    78: op1_13_inv20 = 1;
    79: op1_13_inv20 = 1;
    60: op1_13_inv20 = 1;
    88: op1_13_inv20 = 1;
    80: op1_13_inv20 = 1;
    62: op1_13_inv20 = 1;
    52: op1_13_inv20 = 1;
    64: op1_13_inv20 = 1;
    84: op1_13_inv20 = 1;
    46: op1_13_inv20 = 1;
    65: op1_13_inv20 = 1;
    91: op1_13_inv20 = 1;
    67: op1_13_inv20 = 1;
    92: op1_13_inv20 = 1;
    93: op1_13_inv20 = 1;
    97: op1_13_inv20 = 1;
    99: op1_13_inv20 = 1;
    100: op1_13_inv20 = 1;
    102: op1_13_inv20 = 1;
    103: op1_13_inv20 = 1;
    108: op1_13_inv20 = 1;
    110: op1_13_inv20 = 1;
    111: op1_13_inv20 = 1;
    114: op1_13_inv20 = 1;
    115: op1_13_inv20 = 1;
    47: op1_13_inv20 = 1;
    118: op1_13_inv20 = 1;
    121: op1_13_inv20 = 1;
    122: op1_13_inv20 = 1;
    123: op1_13_inv20 = 1;
    124: op1_13_inv20 = 1;
    126: op1_13_inv20 = 1;
    44: op1_13_inv20 = 1;
    129: op1_13_inv20 = 1;
    default: op1_13_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in21 = reg_1034;
    75: op1_13_in21 = reg_1034;
    53: op1_13_in21 = reg_0024;
    73: op1_13_in21 = reg_0922;
    86: op1_13_in21 = reg_0117;
    74: op1_13_in21 = reg_0576;
    69: op1_13_in21 = reg_0707;
    54: op1_13_in21 = reg_0154;
    49: op1_13_in21 = reg_0002;
    56: op1_13_in21 = reg_0900;
    50: op1_13_in21 = reg_0224;
    76: op1_13_in21 = reg_0672;
    71: op1_13_in21 = reg_0079;
    87: op1_13_in21 = reg_0599;
    115: op1_13_in21 = reg_0599;
    68: op1_13_in21 = reg_1082;
    77: op1_13_in21 = reg_0801;
    61: op1_13_in21 = reg_0968;
    58: op1_13_in21 = reg_0171;
    78: op1_13_in21 = reg_0189;
    70: op1_13_in21 = reg_0480;
    59: op1_13_in21 = reg_0541;
    79: op1_13_in21 = reg_0057;
    51: op1_13_in21 = reg_0775;
    60: op1_13_in21 = reg_0131;
    88: op1_13_in21 = reg_0032;
    80: op1_13_in21 = reg_0090;
    62: op1_13_in21 = reg_0521;
    81: op1_13_in21 = reg_0748;
    63: op1_13_in21 = reg_0379;
    52: op1_13_in21 = reg_0156;
    82: op1_13_in21 = reg_0726;
    83: op1_13_in21 = reg_0297;
    64: op1_13_in21 = reg_0153;
    89: op1_13_in21 = reg_0836;
    84: op1_13_in21 = reg_0080;
    46: op1_13_in21 = imem06_in[3:0];
    85: op1_13_in21 = reg_0937;
    101: op1_13_in21 = reg_0937;
    65: op1_13_in21 = reg_0734;
    90: op1_13_in21 = reg_0397;
    66: op1_13_in21 = reg_1207;
    48: op1_13_in21 = reg_0213;
    91: op1_13_in21 = reg_0932;
    67: op1_13_in21 = reg_0695;
    92: op1_13_in21 = reg_0406;
    93: op1_13_in21 = reg_0957;
    94: op1_13_in21 = reg_0924;
    95: op1_13_in21 = reg_0196;
    96: op1_13_in21 = reg_0665;
    97: op1_13_in21 = reg_1343;
    98: op1_13_in21 = reg_1032;
    99: op1_13_in21 = reg_0694;
    100: op1_13_in21 = reg_0149;
    102: op1_13_in21 = reg_0089;
    103: op1_13_in21 = reg_0168;
    104: op1_13_in21 = reg_0797;
    105: op1_13_in21 = reg_0318;
    106: op1_13_in21 = reg_0519;
    107: op1_13_in21 = reg_0401;
    108: op1_13_in21 = reg_1348;
    109: op1_13_in21 = reg_0235;
    110: op1_13_in21 = reg_0893;
    111: op1_13_in21 = reg_0209;
    112: op1_13_in21 = reg_0225;
    113: op1_13_in21 = reg_0370;
    114: op1_13_in21 = reg_0438;
    116: op1_13_in21 = reg_0438;
    117: op1_13_in21 = reg_0320;
    47: op1_13_in21 = reg_0296;
    118: op1_13_in21 = reg_0272;
    119: op1_13_in21 = reg_1303;
    121: op1_13_in21 = reg_1255;
    122: op1_13_in21 = reg_0053;
    123: op1_13_in21 = reg_1299;
    124: op1_13_in21 = reg_0000;
    125: op1_13_in21 = reg_0461;
    126: op1_13_in21 = imem03_in[11:8];
    44: op1_13_in21 = reg_0066;
    127: op1_13_in21 = reg_0548;
    128: op1_13_in21 = reg_0830;
    129: op1_13_in21 = reg_0973;
    130: op1_13_in21 = reg_0071;
    default: op1_13_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv21 = 1;
    86: op1_13_inv21 = 1;
    74: op1_13_inv21 = 1;
    69: op1_13_inv21 = 1;
    54: op1_13_inv21 = 1;
    49: op1_13_inv21 = 1;
    56: op1_13_inv21 = 1;
    50: op1_13_inv21 = 1;
    76: op1_13_inv21 = 1;
    68: op1_13_inv21 = 1;
    77: op1_13_inv21 = 1;
    61: op1_13_inv21 = 1;
    58: op1_13_inv21 = 1;
    51: op1_13_inv21 = 1;
    62: op1_13_inv21 = 1;
    63: op1_13_inv21 = 1;
    52: op1_13_inv21 = 1;
    82: op1_13_inv21 = 1;
    83: op1_13_inv21 = 1;
    85: op1_13_inv21 = 1;
    90: op1_13_inv21 = 1;
    94: op1_13_inv21 = 1;
    95: op1_13_inv21 = 1;
    96: op1_13_inv21 = 1;
    103: op1_13_inv21 = 1;
    105: op1_13_inv21 = 1;
    106: op1_13_inv21 = 1;
    107: op1_13_inv21 = 1;
    112: op1_13_inv21 = 1;
    113: op1_13_inv21 = 1;
    114: op1_13_inv21 = 1;
    115: op1_13_inv21 = 1;
    119: op1_13_inv21 = 1;
    121: op1_13_inv21 = 1;
    122: op1_13_inv21 = 1;
    123: op1_13_inv21 = 1;
    125: op1_13_inv21 = 1;
    126: op1_13_inv21 = 1;
    44: op1_13_inv21 = 1;
    127: op1_13_inv21 = 1;
    128: op1_13_inv21 = 1;
    130: op1_13_inv21 = 1;
    default: op1_13_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in22 = reg_0788;
    53: op1_13_in22 = reg_0227;
    73: op1_13_in22 = reg_1351;
    86: op1_13_in22 = reg_0020;
    74: op1_13_in22 = reg_0275;
    69: op1_13_in22 = imem03_in[11:8];
    54: op1_13_in22 = reg_0755;
    49: op1_13_in22 = reg_0053;
    75: op1_13_in22 = reg_1254;
    56: op1_13_in22 = reg_0294;
    50: op1_13_in22 = reg_0310;
    76: op1_13_in22 = reg_0135;
    71: op1_13_in22 = reg_0278;
    87: op1_13_in22 = reg_1041;
    92: op1_13_in22 = reg_1041;
    68: op1_13_in22 = reg_0466;
    77: op1_13_in22 = reg_0802;
    61: op1_13_in22 = reg_0930;
    58: op1_13_in22 = reg_1170;
    78: op1_13_in22 = reg_0410;
    70: op1_13_in22 = reg_0734;
    59: op1_13_in22 = reg_0539;
    79: op1_13_in22 = reg_1324;
    51: op1_13_in22 = reg_0661;
    60: op1_13_in22 = reg_0541;
    88: op1_13_in22 = reg_0088;
    80: op1_13_in22 = reg_0576;
    85: op1_13_in22 = reg_0576;
    81: op1_13_in22 = reg_0272;
    63: op1_13_in22 = reg_0381;
    52: op1_13_in22 = reg_0777;
    82: op1_13_in22 = reg_0400;
    83: op1_13_in22 = reg_1345;
    64: op1_13_in22 = reg_0009;
    89: op1_13_in22 = reg_0337;
    84: op1_13_in22 = reg_0078;
    46: op1_13_in22 = reg_0398;
    65: op1_13_in22 = reg_0216;
    90: op1_13_in22 = reg_0863;
    66: op1_13_in22 = reg_0935;
    48: op1_13_in22 = reg_0022;
    91: op1_13_in22 = reg_0210;
    67: op1_13_in22 = reg_0800;
    93: op1_13_in22 = reg_0190;
    94: op1_13_in22 = reg_0923;
    95: op1_13_in22 = reg_1348;
    96: op1_13_in22 = reg_0442;
    97: op1_13_in22 = reg_0433;
    98: op1_13_in22 = reg_0282;
    99: op1_13_in22 = reg_0297;
    100: op1_13_in22 = reg_0868;
    101: op1_13_in22 = reg_1486;
    102: op1_13_in22 = reg_0917;
    103: op1_13_in22 = reg_0759;
    104: op1_13_in22 = reg_0488;
    105: op1_13_in22 = reg_0130;
    107: op1_13_in22 = reg_0047;
    108: op1_13_in22 = reg_0344;
    109: op1_13_in22 = reg_0185;
    110: op1_13_in22 = reg_1416;
    111: op1_13_in22 = reg_0579;
    112: op1_13_in22 = reg_0457;
    113: op1_13_in22 = reg_0204;
    114: op1_13_in22 = reg_1457;
    115: op1_13_in22 = reg_0454;
    116: op1_13_in22 = reg_0148;
    117: op1_13_in22 = reg_0452;
    47: op1_13_in22 = reg_0295;
    118: op1_13_in22 = reg_0205;
    119: op1_13_in22 = reg_1228;
    121: op1_13_in22 = reg_0577;
    122: op1_13_in22 = reg_0519;
    123: op1_13_in22 = reg_0795;
    124: op1_13_in22 = reg_0789;
    125: op1_13_in22 = reg_0246;
    126: op1_13_in22 = reg_1009;
    44: op1_13_in22 = reg_0131;
    127: op1_13_in22 = reg_0610;
    128: op1_13_in22 = reg_0468;
    129: op1_13_in22 = reg_1451;
    130: op1_13_in22 = reg_0073;
    default: op1_13_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv22 = 1;
    69: op1_13_inv22 = 1;
    54: op1_13_inv22 = 1;
    56: op1_13_inv22 = 1;
    50: op1_13_inv22 = 1;
    87: op1_13_inv22 = 1;
    68: op1_13_inv22 = 1;
    77: op1_13_inv22 = 1;
    61: op1_13_inv22 = 1;
    78: op1_13_inv22 = 1;
    70: op1_13_inv22 = 1;
    59: op1_13_inv22 = 1;
    79: op1_13_inv22 = 1;
    60: op1_13_inv22 = 1;
    88: op1_13_inv22 = 1;
    80: op1_13_inv22 = 1;
    63: op1_13_inv22 = 1;
    52: op1_13_inv22 = 1;
    82: op1_13_inv22 = 1;
    64: op1_13_inv22 = 1;
    84: op1_13_inv22 = 1;
    46: op1_13_inv22 = 1;
    91: op1_13_inv22 = 1;
    93: op1_13_inv22 = 1;
    97: op1_13_inv22 = 1;
    98: op1_13_inv22 = 1;
    100: op1_13_inv22 = 1;
    101: op1_13_inv22 = 1;
    102: op1_13_inv22 = 1;
    103: op1_13_inv22 = 1;
    104: op1_13_inv22 = 1;
    105: op1_13_inv22 = 1;
    108: op1_13_inv22 = 1;
    112: op1_13_inv22 = 1;
    115: op1_13_inv22 = 1;
    116: op1_13_inv22 = 1;
    47: op1_13_inv22 = 1;
    118: op1_13_inv22 = 1;
    124: op1_13_inv22 = 1;
    125: op1_13_inv22 = 1;
    126: op1_13_inv22 = 1;
    128: op1_13_inv22 = 1;
    default: op1_13_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in23 = reg_1070;
    53: op1_13_in23 = reg_0375;
    73: op1_13_in23 = reg_0245;
    86: op1_13_in23 = reg_0579;
    74: op1_13_in23 = reg_0196;
    69: op1_13_in23 = imem03_in[15:12];
    54: op1_13_in23 = reg_0732;
    49: op1_13_in23 = reg_0521;
    122: op1_13_in23 = reg_0521;
    75: op1_13_in23 = reg_1256;
    56: op1_13_in23 = reg_0845;
    50: op1_13_in23 = reg_0159;
    76: op1_13_in23 = reg_0851;
    71: op1_13_in23 = reg_0744;
    87: op1_13_in23 = reg_0199;
    92: op1_13_in23 = reg_0199;
    68: op1_13_in23 = reg_0464;
    77: op1_13_in23 = reg_0800;
    61: op1_13_in23 = reg_0727;
    58: op1_13_in23 = reg_0229;
    78: op1_13_in23 = reg_0057;
    70: op1_13_in23 = reg_0426;
    59: op1_13_in23 = reg_0418;
    79: op1_13_in23 = reg_0335;
    51: op1_13_in23 = reg_0739;
    60: op1_13_in23 = reg_0937;
    88: op1_13_in23 = reg_0252;
    80: op1_13_in23 = reg_0197;
    85: op1_13_in23 = reg_0197;
    81: op1_13_in23 = reg_0736;
    63: op1_13_in23 = reg_0878;
    52: op1_13_in23 = reg_0030;
    82: op1_13_in23 = reg_0385;
    83: op1_13_in23 = reg_1094;
    94: op1_13_in23 = reg_1094;
    64: op1_13_in23 = reg_0007;
    89: op1_13_in23 = reg_1151;
    84: op1_13_in23 = reg_0077;
    46: op1_13_in23 = reg_0115;
    65: op1_13_in23 = reg_0707;
    90: op1_13_in23 = reg_1501;
    66: op1_13_in23 = reg_0128;
    129: op1_13_in23 = reg_0128;
    48: op1_13_in23 = reg_0191;
    91: op1_13_in23 = reg_0035;
    67: op1_13_in23 = reg_1132;
    93: op1_13_in23 = reg_0178;
    95: op1_13_in23 = reg_0344;
    105: op1_13_in23 = reg_0344;
    96: op1_13_in23 = reg_0738;
    97: op1_13_in23 = reg_1451;
    98: op1_13_in23 = reg_1255;
    99: op1_13_in23 = reg_0574;
    100: op1_13_in23 = reg_0092;
    101: op1_13_in23 = reg_1485;
    102: op1_13_in23 = reg_0183;
    111: op1_13_in23 = reg_0183;
    103: op1_13_in23 = reg_0377;
    104: op1_13_in23 = reg_0796;
    107: op1_13_in23 = reg_0553;
    108: op1_13_in23 = reg_0799;
    109: op1_13_in23 = reg_0154;
    110: op1_13_in23 = reg_0994;
    112: op1_13_in23 = reg_1350;
    113: op1_13_in23 = reg_0315;
    114: op1_13_in23 = reg_1456;
    115: op1_13_in23 = reg_1419;
    117: op1_13_in23 = reg_1419;
    116: op1_13_in23 = reg_0384;
    47: op1_13_in23 = reg_0419;
    118: op1_13_in23 = reg_1268;
    119: op1_13_in23 = reg_1202;
    121: op1_13_in23 = reg_1290;
    123: op1_13_in23 = imem06_in[3:0];
    124: op1_13_in23 = reg_1495;
    125: op1_13_in23 = reg_0791;
    126: op1_13_in23 = reg_1033;
    44: op1_13_in23 = reg_0331;
    127: op1_13_in23 = reg_0609;
    128: op1_13_in23 = reg_0469;
    130: op1_13_in23 = reg_0089;
    default: op1_13_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_13_inv23 = 1;
    69: op1_13_inv23 = 1;
    75: op1_13_inv23 = 1;
    56: op1_13_inv23 = 1;
    76: op1_13_inv23 = 1;
    71: op1_13_inv23 = 1;
    87: op1_13_inv23 = 1;
    68: op1_13_inv23 = 1;
    58: op1_13_inv23 = 1;
    70: op1_13_inv23 = 1;
    59: op1_13_inv23 = 1;
    88: op1_13_inv23 = 1;
    80: op1_13_inv23 = 1;
    81: op1_13_inv23 = 1;
    63: op1_13_inv23 = 1;
    52: op1_13_inv23 = 1;
    82: op1_13_inv23 = 1;
    89: op1_13_inv23 = 1;
    84: op1_13_inv23 = 1;
    46: op1_13_inv23 = 1;
    65: op1_13_inv23 = 1;
    48: op1_13_inv23 = 1;
    67: op1_13_inv23 = 1;
    92: op1_13_inv23 = 1;
    98: op1_13_inv23 = 1;
    100: op1_13_inv23 = 1;
    107: op1_13_inv23 = 1;
    108: op1_13_inv23 = 1;
    109: op1_13_inv23 = 1;
    110: op1_13_inv23 = 1;
    111: op1_13_inv23 = 1;
    113: op1_13_inv23 = 1;
    116: op1_13_inv23 = 1;
    117: op1_13_inv23 = 1;
    118: op1_13_inv23 = 1;
    119: op1_13_inv23 = 1;
    121: op1_13_inv23 = 1;
    123: op1_13_inv23 = 1;
    124: op1_13_inv23 = 1;
    126: op1_13_inv23 = 1;
    44: op1_13_inv23 = 1;
    127: op1_13_inv23 = 1;
    128: op1_13_inv23 = 1;
    130: op1_13_inv23 = 1;
    default: op1_13_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in24 = reg_0166;
    53: op1_13_in24 = reg_0378;
    73: op1_13_in24 = reg_0703;
    86: op1_13_in24 = reg_0750;
    74: op1_13_in24 = reg_1346;
    69: op1_13_in24 = reg_0376;
    54: op1_13_in24 = imem03_in[3:0];
    49: op1_13_in24 = reg_0483;
    75: op1_13_in24 = reg_0550;
    56: op1_13_in24 = reg_0006;
    50: op1_13_in24 = reg_0156;
    76: op1_13_in24 = reg_0224;
    71: op1_13_in24 = reg_0997;
    87: op1_13_in24 = reg_1065;
    68: op1_13_in24 = reg_1147;
    77: op1_13_in24 = reg_1515;
    61: op1_13_in24 = reg_0402;
    58: op1_13_in24 = reg_0496;
    78: op1_13_in24 = reg_0122;
    70: op1_13_in24 = reg_0898;
    59: op1_13_in24 = reg_0300;
    79: op1_13_in24 = reg_0446;
    51: op1_13_in24 = reg_0621;
    60: op1_13_in24 = reg_0938;
    88: op1_13_in24 = reg_0552;
    80: op1_13_in24 = reg_0275;
    101: op1_13_in24 = reg_0275;
    81: op1_13_in24 = reg_0579;
    63: op1_13_in24 = reg_0829;
    52: op1_13_in24 = reg_0661;
    82: op1_13_in24 = reg_0042;
    83: op1_13_in24 = reg_0777;
    94: op1_13_in24 = reg_0777;
    64: op1_13_in24 = reg_0802;
    89: op1_13_in24 = reg_1189;
    84: op1_13_in24 = reg_0292;
    46: op1_13_in24 = reg_0619;
    85: op1_13_in24 = reg_0118;
    65: op1_13_in24 = reg_0706;
    90: op1_13_in24 = reg_0716;
    66: op1_13_in24 = reg_0112;
    48: op1_13_in24 = reg_0994;
    91: op1_13_in24 = reg_1299;
    67: op1_13_in24 = imem03_in[15:12];
    92: op1_13_in24 = reg_1077;
    93: op1_13_in24 = reg_0107;
    95: op1_13_in24 = reg_0589;
    96: op1_13_in24 = reg_0103;
    97: op1_13_in24 = reg_0128;
    98: op1_13_in24 = reg_0576;
    99: op1_13_in24 = reg_1215;
    100: op1_13_in24 = reg_0257;
    102: op1_13_in24 = reg_0788;
    103: op1_13_in24 = imem03_in[7:4];
    104: op1_13_in24 = reg_0414;
    105: op1_13_in24 = reg_0039;
    107: op1_13_in24 = reg_0258;
    108: op1_13_in24 = reg_0603;
    109: op1_13_in24 = reg_1063;
    110: op1_13_in24 = reg_0219;
    111: op1_13_in24 = reg_1431;
    112: op1_13_in24 = reg_0223;
    113: op1_13_in24 = reg_0832;
    114: op1_13_in24 = reg_0386;
    115: op1_13_in24 = reg_0836;
    116: op1_13_in24 = reg_0362;
    117: op1_13_in24 = reg_1143;
    47: op1_13_in24 = reg_0244;
    118: op1_13_in24 = reg_0251;
    119: op1_13_in24 = reg_0215;
    121: op1_13_in24 = reg_0553;
    122: op1_13_in24 = reg_0484;
    123: op1_13_in24 = reg_0929;
    124: op1_13_in24 = reg_0556;
    125: op1_13_in24 = reg_0867;
    126: op1_13_in24 = reg_1001;
    44: op1_13_in24 = reg_0318;
    127: op1_13_in24 = reg_0241;
    128: op1_13_in24 = reg_0968;
    129: op1_13_in24 = reg_0127;
    130: op1_13_in24 = reg_0027;
    default: op1_13_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv24 = 1;
    73: op1_13_inv24 = 1;
    86: op1_13_inv24 = 1;
    69: op1_13_inv24 = 1;
    54: op1_13_inv24 = 1;
    50: op1_13_inv24 = 1;
    76: op1_13_inv24 = 1;
    71: op1_13_inv24 = 1;
    87: op1_13_inv24 = 1;
    58: op1_13_inv24 = 1;
    78: op1_13_inv24 = 1;
    70: op1_13_inv24 = 1;
    88: op1_13_inv24 = 1;
    81: op1_13_inv24 = 1;
    63: op1_13_inv24 = 1;
    52: op1_13_inv24 = 1;
    83: op1_13_inv24 = 1;
    89: op1_13_inv24 = 1;
    84: op1_13_inv24 = 1;
    46: op1_13_inv24 = 1;
    66: op1_13_inv24 = 1;
    48: op1_13_inv24 = 1;
    67: op1_13_inv24 = 1;
    92: op1_13_inv24 = 1;
    93: op1_13_inv24 = 1;
    94: op1_13_inv24 = 1;
    95: op1_13_inv24 = 1;
    98: op1_13_inv24 = 1;
    101: op1_13_inv24 = 1;
    102: op1_13_inv24 = 1;
    103: op1_13_inv24 = 1;
    104: op1_13_inv24 = 1;
    112: op1_13_inv24 = 1;
    114: op1_13_inv24 = 1;
    116: op1_13_inv24 = 1;
    117: op1_13_inv24 = 1;
    119: op1_13_inv24 = 1;
    121: op1_13_inv24 = 1;
    122: op1_13_inv24 = 1;
    126: op1_13_inv24 = 1;
    44: op1_13_inv24 = 1;
    129: op1_13_inv24 = 1;
    130: op1_13_inv24 = 1;
    default: op1_13_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in25 = reg_0258;
    53: op1_13_in25 = imem03_in[3:0];
    73: op1_13_in25 = reg_0299;
    86: op1_13_in25 = reg_1269;
    74: op1_13_in25 = reg_0631;
    69: op1_13_in25 = reg_1003;
    54: op1_13_in25 = reg_0709;
    75: op1_13_in25 = reg_0787;
    56: op1_13_in25 = reg_0154;
    50: op1_13_in25 = reg_0779;
    76: op1_13_in25 = reg_0031;
    71: op1_13_in25 = reg_0184;
    59: op1_13_in25 = reg_0184;
    87: op1_13_in25 = reg_0451;
    68: op1_13_in25 = reg_0407;
    104: op1_13_in25 = reg_0407;
    77: op1_13_in25 = reg_1132;
    61: op1_13_in25 = reg_0384;
    58: op1_13_in25 = reg_0225;
    110: op1_13_in25 = reg_0225;
    78: op1_13_in25 = reg_0446;
    70: op1_13_in25 = reg_1384;
    79: op1_13_in25 = reg_1255;
    51: op1_13_in25 = reg_0591;
    60: op1_13_in25 = reg_0301;
    88: op1_13_in25 = reg_1200;
    80: op1_13_in25 = reg_0130;
    81: op1_13_in25 = reg_0174;
    118: op1_13_in25 = reg_0174;
    63: op1_13_in25 = reg_0024;
    52: op1_13_in25 = reg_0285;
    82: op1_13_in25 = reg_0486;
    83: op1_13_in25 = reg_0774;
    64: op1_13_in25 = reg_0311;
    89: op1_13_in25 = reg_0236;
    84: op1_13_in25 = imem01_in[11:8];
    46: op1_13_in25 = reg_0617;
    85: op1_13_in25 = reg_0602;
    65: op1_13_in25 = reg_1033;
    90: op1_13_in25 = reg_0718;
    66: op1_13_in25 = reg_0106;
    48: op1_13_in25 = reg_0993;
    91: op1_13_in25 = reg_0333;
    67: op1_13_in25 = reg_0375;
    92: op1_13_in25 = reg_0337;
    93: op1_13_in25 = reg_0288;
    94: op1_13_in25 = reg_0775;
    95: op1_13_in25 = reg_0799;
    96: op1_13_in25 = reg_0228;
    97: op1_13_in25 = reg_0111;
    98: op1_13_in25 = reg_0930;
    99: op1_13_in25 = reg_0537;
    100: op1_13_in25 = reg_0499;
    101: op1_13_in25 = reg_1348;
    102: op1_13_in25 = reg_0282;
    103: op1_13_in25 = reg_0732;
    105: op1_13_in25 = imem06_in[11:8];
    107: op1_13_in25 = reg_0547;
    108: op1_13_in25 = reg_0014;
    109: op1_13_in25 = reg_0557;
    111: op1_13_in25 = reg_0702;
    113: op1_13_in25 = reg_0702;
    112: op1_13_in25 = reg_0661;
    114: op1_13_in25 = reg_0385;
    115: op1_13_in25 = reg_1312;
    116: op1_13_in25 = reg_0875;
    117: op1_13_in25 = reg_0062;
    47: op1_13_in25 = reg_0458;
    119: op1_13_in25 = reg_0214;
    121: op1_13_in25 = reg_0463;
    122: op1_13_in25 = reg_1182;
    123: op1_13_in25 = reg_0669;
    124: op1_13_in25 = reg_1184;
    125: op1_13_in25 = reg_0498;
    126: op1_13_in25 = reg_0191;
    44: op1_13_in25 = reg_0492;
    127: op1_13_in25 = reg_1474;
    128: op1_13_in25 = reg_0439;
    129: op1_13_in25 = reg_0802;
    130: op1_13_in25 = reg_0238;
    default: op1_13_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv25 = 1;
    53: op1_13_inv25 = 1;
    73: op1_13_inv25 = 1;
    86: op1_13_inv25 = 1;
    69: op1_13_inv25 = 1;
    54: op1_13_inv25 = 1;
    75: op1_13_inv25 = 1;
    50: op1_13_inv25 = 1;
    68: op1_13_inv25 = 1;
    58: op1_13_inv25 = 1;
    78: op1_13_inv25 = 1;
    79: op1_13_inv25 = 1;
    60: op1_13_inv25 = 1;
    80: op1_13_inv25 = 1;
    63: op1_13_inv25 = 1;
    52: op1_13_inv25 = 1;
    82: op1_13_inv25 = 1;
    64: op1_13_inv25 = 1;
    46: op1_13_inv25 = 1;
    66: op1_13_inv25 = 1;
    91: op1_13_inv25 = 1;
    92: op1_13_inv25 = 1;
    93: op1_13_inv25 = 1;
    94: op1_13_inv25 = 1;
    96: op1_13_inv25 = 1;
    97: op1_13_inv25 = 1;
    98: op1_13_inv25 = 1;
    99: op1_13_inv25 = 1;
    102: op1_13_inv25 = 1;
    105: op1_13_inv25 = 1;
    110: op1_13_inv25 = 1;
    111: op1_13_inv25 = 1;
    115: op1_13_inv25 = 1;
    118: op1_13_inv25 = 1;
    119: op1_13_inv25 = 1;
    126: op1_13_inv25 = 1;
    44: op1_13_inv25 = 1;
    127: op1_13_inv25 = 1;
    129: op1_13_inv25 = 1;
    default: op1_13_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in26 = reg_0463;
    53: op1_13_in26 = imem03_in[11:8];
    73: op1_13_in26 = reg_0740;
    86: op1_13_in26 = reg_0272;
    74: op1_13_in26 = reg_0151;
    60: op1_13_in26 = reg_0151;
    69: op1_13_in26 = reg_1301;
    54: op1_13_in26 = reg_0378;
    75: op1_13_in26 = reg_0222;
    56: op1_13_in26 = reg_0830;
    107: op1_13_in26 = reg_0830;
    50: op1_13_in26 = reg_0029;
    76: op1_13_in26 = reg_0029;
    71: op1_13_in26 = reg_1029;
    87: op1_13_in26 = reg_0698;
    68: op1_13_in26 = reg_0797;
    77: op1_13_in26 = reg_1495;
    61: op1_13_in26 = reg_0047;
    58: op1_13_in26 = reg_0245;
    78: op1_13_in26 = reg_1290;
    70: op1_13_in26 = reg_1383;
    59: op1_13_in26 = reg_0240;
    80: op1_13_in26 = reg_0240;
    79: op1_13_in26 = reg_1254;
    102: op1_13_in26 = reg_1254;
    51: op1_13_in26 = reg_0137;
    88: op1_13_in26 = reg_0488;
    81: op1_13_in26 = reg_0167;
    63: op1_13_in26 = reg_0280;
    52: op1_13_in26 = reg_0741;
    82: op1_13_in26 = reg_0607;
    83: op1_13_in26 = reg_0030;
    64: op1_13_in26 = reg_0756;
    89: op1_13_in26 = imem05_in[3:0];
    84: op1_13_in26 = reg_0011;
    46: op1_13_in26 = reg_0584;
    85: op1_13_in26 = reg_1346;
    65: op1_13_in26 = reg_0559;
    90: op1_13_in26 = reg_0637;
    66: op1_13_in26 = reg_0381;
    48: op1_13_in26 = reg_0995;
    91: op1_13_in26 = reg_1169;
    67: op1_13_in26 = reg_0143;
    126: op1_13_in26 = reg_0143;
    92: op1_13_in26 = reg_1151;
    93: op1_13_in26 = reg_1282;
    94: op1_13_in26 = reg_0031;
    95: op1_13_in26 = reg_0729;
    96: op1_13_in26 = reg_0050;
    97: op1_13_in26 = reg_0829;
    98: op1_13_in26 = reg_0239;
    99: op1_13_in26 = reg_0451;
    100: op1_13_in26 = reg_0475;
    101: op1_13_in26 = reg_0799;
    103: op1_13_in26 = reg_0600;
    104: op1_13_in26 = reg_0199;
    105: op1_13_in26 = imem06_in[15:12];
    108: op1_13_in26 = reg_0670;
    109: op1_13_in26 = reg_1001;
    110: op1_13_in26 = reg_0851;
    111: op1_13_in26 = reg_1268;
    112: op1_13_in26 = reg_0285;
    113: op1_13_in26 = reg_0992;
    114: op1_13_in26 = reg_0360;
    115: op1_13_in26 = reg_0096;
    116: op1_13_in26 = reg_0292;
    117: op1_13_in26 = reg_0835;
    47: op1_13_in26 = reg_0212;
    118: op1_13_in26 = reg_0562;
    119: op1_13_in26 = reg_0017;
    121: op1_13_in26 = reg_0743;
    123: op1_13_in26 = reg_0782;
    124: op1_13_in26 = reg_0070;
    125: op1_13_in26 = reg_0994;
    44: op1_13_in26 = imem05_in[15:12];
    127: op1_13_in26 = reg_0430;
    128: op1_13_in26 = reg_0434;
    129: op1_13_in26 = reg_0279;
    130: op1_13_in26 = reg_0320;
    default: op1_13_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv26 = 1;
    53: op1_13_inv26 = 1;
    54: op1_13_inv26 = 1;
    75: op1_13_inv26 = 1;
    71: op1_13_inv26 = 1;
    68: op1_13_inv26 = 1;
    77: op1_13_inv26 = 1;
    70: op1_13_inv26 = 1;
    51: op1_13_inv26 = 1;
    60: op1_13_inv26 = 1;
    80: op1_13_inv26 = 1;
    84: op1_13_inv26 = 1;
    46: op1_13_inv26 = 1;
    85: op1_13_inv26 = 1;
    65: op1_13_inv26 = 1;
    66: op1_13_inv26 = 1;
    48: op1_13_inv26 = 1;
    67: op1_13_inv26 = 1;
    92: op1_13_inv26 = 1;
    93: op1_13_inv26 = 1;
    94: op1_13_inv26 = 1;
    95: op1_13_inv26 = 1;
    96: op1_13_inv26 = 1;
    97: op1_13_inv26 = 1;
    99: op1_13_inv26 = 1;
    102: op1_13_inv26 = 1;
    103: op1_13_inv26 = 1;
    105: op1_13_inv26 = 1;
    111: op1_13_inv26 = 1;
    112: op1_13_inv26 = 1;
    113: op1_13_inv26 = 1;
    116: op1_13_inv26 = 1;
    117: op1_13_inv26 = 1;
    47: op1_13_inv26 = 1;
    118: op1_13_inv26 = 1;
    119: op1_13_inv26 = 1;
    121: op1_13_inv26 = 1;
    123: op1_13_inv26 = 1;
    125: op1_13_inv26 = 1;
    44: op1_13_inv26 = 1;
    130: op1_13_inv26 = 1;
    default: op1_13_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in27 = reg_0420;
    53: op1_13_in27 = reg_0049;
    73: op1_13_in27 = reg_0415;
    86: op1_13_in27 = reg_0700;
    74: op1_13_in27 = reg_0828;
    69: op1_13_in27 = reg_0107;
    54: op1_13_in27 = reg_0177;
    75: op1_13_in27 = reg_0830;
    56: op1_13_in27 = reg_0024;
    50: op1_13_in27 = reg_0030;
    76: op1_13_in27 = reg_0665;
    83: op1_13_in27 = reg_0665;
    71: op1_13_in27 = reg_0532;
    87: op1_13_in27 = reg_0304;
    68: op1_13_in27 = reg_0936;
    77: op1_13_in27 = reg_0999;
    61: op1_13_in27 = reg_0093;
    58: op1_13_in27 = reg_0674;
    78: op1_13_in27 = reg_0788;
    70: op1_13_in27 = reg_1372;
    59: op1_13_in27 = reg_0274;
    79: op1_13_in27 = reg_0258;
    51: op1_13_in27 = reg_0100;
    60: op1_13_in27 = reg_0206;
    88: op1_13_in27 = reg_0500;
    80: op1_13_in27 = reg_0631;
    81: op1_13_in27 = reg_1402;
    63: op1_13_in27 = reg_1132;
    52: op1_13_in27 = reg_0623;
    82: op1_13_in27 = reg_0846;
    64: op1_13_in27 = reg_0677;
    89: op1_13_in27 = reg_0205;
    84: op1_13_in27 = reg_0457;
    46: op1_13_in27 = reg_0571;
    85: op1_13_in27 = reg_0799;
    65: op1_13_in27 = reg_1301;
    90: op1_13_in27 = reg_0398;
    66: op1_13_in27 = reg_0876;
    48: op1_13_in27 = reg_0703;
    91: op1_13_in27 = reg_0992;
    67: op1_13_in27 = reg_0964;
    92: op1_13_in27 = reg_1189;
    93: op1_13_in27 = reg_1280;
    94: op1_13_in27 = reg_0465;
    95: op1_13_in27 = reg_0195;
    96: op1_13_in27 = reg_0001;
    97: op1_13_in27 = reg_0379;
    98: op1_13_in27 = reg_0241;
    99: op1_13_in27 = reg_1419;
    100: op1_13_in27 = reg_0626;
    101: op1_13_in27 = reg_0603;
    102: op1_13_in27 = reg_0166;
    103: op1_13_in27 = reg_1495;
    104: op1_13_in27 = reg_1004;
    105: op1_13_in27 = reg_0755;
    107: op1_13_in27 = reg_0798;
    108: op1_13_in27 = imem06_in[3:0];
    109: op1_13_in27 = reg_0311;
    110: op1_13_in27 = reg_1350;
    111: op1_13_in27 = reg_0251;
    112: op1_13_in27 = reg_0286;
    113: op1_13_in27 = reg_0831;
    114: op1_13_in27 = reg_0875;
    115: op1_13_in27 = reg_0904;
    116: op1_13_in27 = reg_0728;
    117: op1_13_in27 = reg_1312;
    47: op1_13_in27 = reg_0215;
    118: op1_13_in27 = reg_0173;
    119: op1_13_in27 = reg_0050;
    121: op1_13_in27 = reg_0238;
    123: op1_13_in27 = reg_0751;
    124: op1_13_in27 = reg_1092;
    125: op1_13_in27 = imem07_in[15:12];
    126: op1_13_in27 = reg_0142;
    44: op1_13_in27 = reg_0070;
    127: op1_13_in27 = reg_0438;
    128: op1_13_in27 = reg_1457;
    129: op1_13_in27 = reg_0707;
    130: op1_13_in27 = reg_0047;
    default: op1_13_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv27 = 1;
    53: op1_13_inv27 = 1;
    73: op1_13_inv27 = 1;
    54: op1_13_inv27 = 1;
    75: op1_13_inv27 = 1;
    56: op1_13_inv27 = 1;
    50: op1_13_inv27 = 1;
    68: op1_13_inv27 = 1;
    77: op1_13_inv27 = 1;
    61: op1_13_inv27 = 1;
    79: op1_13_inv27 = 1;
    60: op1_13_inv27 = 1;
    88: op1_13_inv27 = 1;
    81: op1_13_inv27 = 1;
    52: op1_13_inv27 = 1;
    82: op1_13_inv27 = 1;
    83: op1_13_inv27 = 1;
    90: op1_13_inv27 = 1;
    66: op1_13_inv27 = 1;
    95: op1_13_inv27 = 1;
    97: op1_13_inv27 = 1;
    98: op1_13_inv27 = 1;
    100: op1_13_inv27 = 1;
    102: op1_13_inv27 = 1;
    104: op1_13_inv27 = 1;
    105: op1_13_inv27 = 1;
    107: op1_13_inv27 = 1;
    109: op1_13_inv27 = 1;
    110: op1_13_inv27 = 1;
    112: op1_13_inv27 = 1;
    113: op1_13_inv27 = 1;
    114: op1_13_inv27 = 1;
    115: op1_13_inv27 = 1;
    116: op1_13_inv27 = 1;
    118: op1_13_inv27 = 1;
    123: op1_13_inv27 = 1;
    124: op1_13_inv27 = 1;
    125: op1_13_inv27 = 1;
    126: op1_13_inv27 = 1;
    129: op1_13_inv27 = 1;
    default: op1_13_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in28 = reg_0241;
    53: op1_13_in28 = reg_0232;
    77: op1_13_in28 = reg_0232;
    104: op1_13_in28 = reg_0232;
    129: op1_13_in28 = reg_0232;
    73: op1_13_in28 = reg_0618;
    86: op1_13_in28 = reg_0648;
    74: op1_13_in28 = reg_0377;
    69: op1_13_in28 = reg_0104;
    54: op1_13_in28 = reg_0049;
    75: op1_13_in28 = reg_0798;
    56: op1_13_in28 = reg_0801;
    50: op1_13_in28 = reg_0663;
    76: op1_13_in28 = reg_0740;
    71: op1_13_in28 = reg_0533;
    87: op1_13_in28 = reg_0932;
    68: op1_13_in28 = reg_0451;
    61: op1_13_in28 = reg_0724;
    58: op1_13_in28 = reg_0791;
    78: op1_13_in28 = reg_1255;
    70: op1_13_in28 = reg_1368;
    59: op1_13_in28 = reg_0039;
    79: op1_13_in28 = reg_1473;
    51: op1_13_in28 = reg_0321;
    60: op1_13_in28 = reg_0752;
    88: op1_13_in28 = reg_1214;
    80: op1_13_in28 = reg_0151;
    81: op1_13_in28 = reg_0183;
    63: op1_13_in28 = reg_0312;
    52: op1_13_in28 = reg_0103;
    82: op1_13_in28 = reg_1344;
    83: op1_13_in28 = reg_0287;
    64: op1_13_in28 = reg_0678;
    89: op1_13_in28 = reg_0578;
    84: op1_13_in28 = reg_0590;
    46: op1_13_in28 = reg_0269;
    85: op1_13_in28 = reg_0207;
    65: op1_13_in28 = reg_0479;
    90: op1_13_in28 = reg_0373;
    66: op1_13_in28 = reg_0878;
    48: op1_13_in28 = reg_0892;
    91: op1_13_in28 = reg_0831;
    67: op1_13_in28 = reg_0962;
    92: op1_13_in28 = reg_0117;
    93: op1_13_in28 = imem04_in[7:4];
    94: op1_13_in28 = reg_0665;
    95: op1_13_in28 = reg_0825;
    96: op1_13_in28 = reg_0053;
    97: op1_13_in28 = reg_1492;
    98: op1_13_in28 = reg_1475;
    99: op1_13_in28 = reg_0719;
    100: op1_13_in28 = reg_0607;
    101: op1_13_in28 = reg_0828;
    102: op1_13_in28 = reg_1512;
    103: op1_13_in28 = reg_1313;
    105: op1_13_in28 = reg_0870;
    107: op1_13_in28 = reg_0572;
    108: op1_13_in28 = imem06_in[11:8];
    109: op1_13_in28 = reg_0234;
    110: op1_13_in28 = reg_1347;
    111: op1_13_in28 = reg_0174;
    112: op1_13_in28 = reg_0441;
    113: op1_13_in28 = reg_0173;
    114: op1_13_in28 = reg_0464;
    115: op1_13_in28 = reg_0540;
    116: op1_13_in28 = reg_1068;
    117: op1_13_in28 = reg_1146;
    47: op1_13_in28 = reg_0921;
    118: op1_13_in28 = reg_0391;
    119: op1_13_in28 = reg_1095;
    121: op1_13_in28 = reg_1474;
    123: op1_13_in28 = reg_0720;
    124: op1_13_in28 = reg_1208;
    125: op1_13_in28 = reg_1056;
    126: op1_13_in28 = reg_1199;
    44: op1_13_in28 = reg_0890;
    127: op1_13_in28 = reg_0149;
    128: op1_13_in28 = reg_1456;
    130: op1_13_in28 = imem01_in[7:4];
    default: op1_13_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_13_inv28 = 1;
    53: op1_13_inv28 = 1;
    54: op1_13_inv28 = 1;
    71: op1_13_inv28 = 1;
    87: op1_13_inv28 = 1;
    77: op1_13_inv28 = 1;
    78: op1_13_inv28 = 1;
    70: op1_13_inv28 = 1;
    80: op1_13_inv28 = 1;
    81: op1_13_inv28 = 1;
    52: op1_13_inv28 = 1;
    46: op1_13_inv28 = 1;
    85: op1_13_inv28 = 1;
    65: op1_13_inv28 = 1;
    90: op1_13_inv28 = 1;
    48: op1_13_inv28 = 1;
    91: op1_13_inv28 = 1;
    67: op1_13_inv28 = 1;
    94: op1_13_inv28 = 1;
    95: op1_13_inv28 = 1;
    96: op1_13_inv28 = 1;
    100: op1_13_inv28 = 1;
    101: op1_13_inv28 = 1;
    103: op1_13_inv28 = 1;
    105: op1_13_inv28 = 1;
    108: op1_13_inv28 = 1;
    109: op1_13_inv28 = 1;
    111: op1_13_inv28 = 1;
    115: op1_13_inv28 = 1;
    116: op1_13_inv28 = 1;
    117: op1_13_inv28 = 1;
    47: op1_13_inv28 = 1;
    118: op1_13_inv28 = 1;
    121: op1_13_inv28 = 1;
    128: op1_13_inv28 = 1;
    default: op1_13_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in29 = reg_1475;
    53: op1_13_in29 = reg_0233;
    73: op1_13_in29 = reg_0620;
    86: op1_13_in29 = reg_0174;
    91: op1_13_in29 = reg_0174;
    74: op1_13_in29 = reg_0795;
    69: op1_13_in29 = reg_0504;
    54: op1_13_in29 = reg_0180;
    75: op1_13_in29 = reg_0612;
    56: op1_13_in29 = reg_0325;
    50: op1_13_in29 = reg_0664;
    76: op1_13_in29 = reg_0404;
    71: op1_13_in29 = reg_0169;
    87: op1_13_in29 = reg_0117;
    68: op1_13_in29 = reg_0320;
    77: op1_13_in29 = reg_1149;
    61: op1_13_in29 = reg_0278;
    58: op1_13_in29 = reg_0779;
    78: op1_13_in29 = imem01_in[3:0];
    70: op1_13_in29 = reg_1339;
    59: op1_13_in29 = reg_1035;
    79: op1_13_in29 = reg_1474;
    51: op1_13_in29 = reg_0053;
    60: op1_13_in29 = reg_0907;
    88: op1_13_in29 = reg_1147;
    80: op1_13_in29 = reg_0828;
    81: op1_13_in29 = reg_0301;
    63: op1_13_in29 = reg_0525;
    52: op1_13_in29 = reg_0051;
    82: op1_13_in29 = reg_0256;
    83: op1_13_in29 = reg_0286;
    64: op1_13_in29 = reg_0706;
    89: op1_13_in29 = reg_0733;
    84: op1_13_in29 = reg_1235;
    46: op1_13_in29 = reg_0046;
    85: op1_13_in29 = reg_0669;
    65: op1_13_in29 = reg_0411;
    90: op1_13_in29 = reg_0586;
    66: op1_13_in29 = reg_0846;
    48: op1_13_in29 = reg_0310;
    67: op1_13_in29 = reg_0220;
    92: op1_13_in29 = reg_0536;
    93: op1_13_in29 = reg_0034;
    94: op1_13_in29 = reg_0366;
    95: op1_13_in29 = reg_0908;
    96: op1_13_in29 = reg_0521;
    97: op1_13_in29 = reg_1098;
    98: op1_13_in29 = reg_0715;
    121: op1_13_in29 = reg_0715;
    99: op1_13_in29 = reg_0339;
    100: op1_13_in29 = reg_0845;
    101: op1_13_in29 = reg_0038;
    102: op1_13_in29 = reg_0093;
    103: op1_13_in29 = reg_0627;
    104: op1_13_in29 = reg_0340;
    105: op1_13_in29 = reg_1209;
    107: op1_13_in29 = reg_0146;
    108: op1_13_in29 = reg_0270;
    109: op1_13_in29 = reg_1516;
    110: op1_13_in29 = reg_0157;
    111: op1_13_in29 = reg_0392;
    112: op1_13_in29 = reg_0739;
    113: op1_13_in29 = reg_1104;
    114: op1_13_in29 = reg_0043;
    115: op1_13_in29 = reg_0579;
    116: op1_13_in29 = reg_0659;
    117: op1_13_in29 = reg_0932;
    47: op1_13_in29 = reg_0135;
    118: op1_13_in29 = reg_0630;
    119: op1_13_in29 = reg_0993;
    123: op1_13_in29 = reg_1323;
    124: op1_13_in29 = reg_0884;
    125: op1_13_in29 = reg_0703;
    126: op1_13_in29 = reg_0107;
    44: op1_13_in29 = reg_0895;
    127: op1_13_in29 = reg_0148;
    128: op1_13_in29 = reg_0269;
    129: op1_13_in29 = reg_1003;
    130: op1_13_in29 = reg_0902;
    default: op1_13_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv29 = 1;
    86: op1_13_inv29 = 1;
    74: op1_13_inv29 = 1;
    69: op1_13_inv29 = 1;
    54: op1_13_inv29 = 1;
    56: op1_13_inv29 = 1;
    71: op1_13_inv29 = 1;
    87: op1_13_inv29 = 1;
    77: op1_13_inv29 = 1;
    61: op1_13_inv29 = 1;
    58: op1_13_inv29 = 1;
    70: op1_13_inv29 = 1;
    59: op1_13_inv29 = 1;
    79: op1_13_inv29 = 1;
    63: op1_13_inv29 = 1;
    52: op1_13_inv29 = 1;
    82: op1_13_inv29 = 1;
    64: op1_13_inv29 = 1;
    89: op1_13_inv29 = 1;
    46: op1_13_inv29 = 1;
    66: op1_13_inv29 = 1;
    91: op1_13_inv29 = 1;
    92: op1_13_inv29 = 1;
    93: op1_13_inv29 = 1;
    94: op1_13_inv29 = 1;
    95: op1_13_inv29 = 1;
    96: op1_13_inv29 = 1;
    100: op1_13_inv29 = 1;
    102: op1_13_inv29 = 1;
    104: op1_13_inv29 = 1;
    105: op1_13_inv29 = 1;
    107: op1_13_inv29 = 1;
    108: op1_13_inv29 = 1;
    109: op1_13_inv29 = 1;
    110: op1_13_inv29 = 1;
    111: op1_13_inv29 = 1;
    115: op1_13_inv29 = 1;
    118: op1_13_inv29 = 1;
    119: op1_13_inv29 = 1;
    121: op1_13_inv29 = 1;
    124: op1_13_inv29 = 1;
    127: op1_13_inv29 = 1;
    129: op1_13_inv29 = 1;
    default: op1_13_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_13_in30 = reg_1474;
    53: op1_13_in30 = reg_0178;
    73: op1_13_in30 = reg_0065;
    92: op1_13_in30 = reg_0065;
    86: op1_13_in30 = reg_0392;
    74: op1_13_in30 = reg_0192;
    69: op1_13_in30 = reg_0831;
    54: op1_13_in30 = reg_0963;
    75: op1_13_in30 = reg_0439;
    79: op1_13_in30 = reg_0439;
    56: op1_13_in30 = reg_0675;
    50: op1_13_in30 = reg_0287;
    76: op1_13_in30 = reg_0591;
    71: op1_13_in30 = reg_0475;
    87: op1_13_in30 = reg_0633;
    68: op1_13_in30 = imem04_in[3:0];
    65: op1_13_in30 = imem04_in[3:0];
    77: op1_13_in30 = reg_0199;
    61: op1_13_in30 = reg_0043;
    58: op1_13_in30 = reg_0030;
    78: op1_13_in30 = imem01_in[15:12];
    70: op1_13_in30 = reg_1198;
    59: op1_13_in30 = reg_0754;
    51: op1_13_in30 = reg_0087;
    60: op1_13_in30 = reg_0859;
    88: op1_13_in30 = reg_0421;
    80: op1_13_in30 = reg_0984;
    81: op1_13_in30 = reg_1486;
    63: op1_13_in30 = reg_0734;
    52: op1_13_in30 = reg_0086;
    82: op1_13_in30 = reg_0822;
    83: op1_13_in30 = reg_0050;
    64: op1_13_in30 = reg_0143;
    89: op1_13_in30 = reg_1168;
    84: op1_13_in30 = reg_0845;
    46: op1_13_in30 = reg_0152;
    85: op1_13_in30 = reg_0795;
    90: op1_13_in30 = reg_0270;
    66: op1_13_in30 = imem02_in[15:12];
    48: op1_13_in30 = reg_0867;
    91: op1_13_in30 = reg_0604;
    67: op1_13_in30 = reg_0882;
    93: op1_13_in30 = reg_0731;
    94: op1_13_in30 = reg_0740;
    95: op1_13_in30 = reg_0870;
    96: op1_13_in30 = reg_0484;
    97: op1_13_in30 = reg_0801;
    98: op1_13_in30 = reg_0967;
    99: op1_13_in30 = reg_0904;
    100: op1_13_in30 = reg_0455;
    101: op1_13_in30 = reg_0635;
    102: op1_13_in30 = reg_0746;
    103: op1_13_in30 = reg_1226;
    104: op1_13_in30 = reg_0338;
    105: op1_13_in30 = reg_0316;
    107: op1_13_in30 = reg_0363;
    108: op1_13_in30 = reg_0397;
    109: op1_13_in30 = reg_1093;
    110: op1_13_in30 = reg_0366;
    111: op1_13_in30 = reg_0391;
    112: op1_13_in30 = reg_0741;
    113: op1_13_in30 = reg_0564;
    114: op1_13_in30 = reg_0042;
    115: op1_13_in30 = reg_0702;
    116: op1_13_in30 = reg_0608;
    117: op1_13_in30 = reg_0117;
    47: op1_13_in30 = reg_0252;
    118: op1_13_in30 = reg_1403;
    119: op1_13_in30 = reg_1440;
    121: op1_13_in30 = reg_0469;
    123: op1_13_in30 = reg_0752;
    124: op1_13_in30 = reg_0638;
    125: op1_13_in30 = reg_0851;
    126: op1_13_in30 = reg_0313;
    44: op1_13_in30 = reg_0303;
    127: op1_13_in30 = reg_1032;
    128: op1_13_in30 = reg_0679;
    129: op1_13_in30 = reg_0557;
    130: op1_13_in30 = reg_0401;
    default: op1_13_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_13_inv30 = 1;
    74: op1_13_inv30 = 1;
    69: op1_13_inv30 = 1;
    54: op1_13_inv30 = 1;
    75: op1_13_inv30 = 1;
    56: op1_13_inv30 = 1;
    71: op1_13_inv30 = 1;
    77: op1_13_inv30 = 1;
    61: op1_13_inv30 = 1;
    58: op1_13_inv30 = 1;
    78: op1_13_inv30 = 1;
    59: op1_13_inv30 = 1;
    79: op1_13_inv30 = 1;
    60: op1_13_inv30 = 1;
    81: op1_13_inv30 = 1;
    63: op1_13_inv30 = 1;
    52: op1_13_inv30 = 1;
    89: op1_13_inv30 = 1;
    46: op1_13_inv30 = 1;
    85: op1_13_inv30 = 1;
    65: op1_13_inv30 = 1;
    91: op1_13_inv30 = 1;
    93: op1_13_inv30 = 1;
    94: op1_13_inv30 = 1;
    95: op1_13_inv30 = 1;
    96: op1_13_inv30 = 1;
    100: op1_13_inv30 = 1;
    103: op1_13_inv30 = 1;
    107: op1_13_inv30 = 1;
    109: op1_13_inv30 = 1;
    110: op1_13_inv30 = 1;
    111: op1_13_inv30 = 1;
    113: op1_13_inv30 = 1;
    115: op1_13_inv30 = 1;
    116: op1_13_inv30 = 1;
    117: op1_13_inv30 = 1;
    47: op1_13_inv30 = 1;
    119: op1_13_inv30 = 1;
    121: op1_13_inv30 = 1;
    124: op1_13_inv30 = 1;
    126: op1_13_inv30 = 1;
    128: op1_13_inv30 = 1;
    129: op1_13_inv30 = 1;
    130: op1_13_inv30 = 1;
    default: op1_13_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_13_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#13の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_13_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in00 = reg_0616;
    53: op1_14_in00 = reg_0833;
    73: op1_14_in00 = reg_0580;
    55: op1_14_in00 = reg_0729;
    86: op1_14_in00 = reg_0261;
    74: op1_14_in00 = reg_0974;
    54: op1_14_in00 = reg_0342;
    75: op1_14_in00 = reg_0021;
    49: op1_14_in00 = reg_0193;
    69: op1_14_in00 = reg_0013;
    56: op1_14_in00 = reg_0220;
    50: op1_14_in00 = reg_0171;
    76: op1_14_in00 = reg_0554;
    71: op1_14_in00 = reg_0554;
    85: op1_14_in00 = reg_0554;
    87: op1_14_in00 = reg_1132;
    57: op1_14_in00 = reg_0670;
    68: op1_14_in00 = reg_0255;
    77: op1_14_in00 = reg_1147;
    61: op1_14_in00 = reg_0791;
    91: op1_14_in00 = reg_0791;
    78: op1_14_in00 = reg_0020;
    58: op1_14_in00 = reg_0092;
    70: op1_14_in00 = reg_0142;
    59: op1_14_in00 = reg_0340;
    79: op1_14_in00 = reg_0207;
    51: op1_14_in00 = reg_0746;
    60: op1_14_in00 = reg_0144;
    80: op1_14_in00 = reg_0458;
    88: op1_14_in00 = reg_0577;
    62: op1_14_in00 = reg_0629;
    81: op1_14_in00 = reg_1485;
    82: op1_14_in00 = reg_1074;
    52: op1_14_in00 = reg_0635;
    63: op1_14_in00 = reg_0230;
    64: op1_14_in00 = reg_0789;
    83: op1_14_in00 = reg_1510;
    89: op1_14_in00 = reg_0448;
    84: op1_14_in00 = reg_0996;
    65: op1_14_in00 = reg_0907;
    90: op1_14_in00 = reg_0573;
    66: op1_14_in00 = reg_0609;
    48: op1_14_in00 = reg_0541;
    46: op1_14_in00 = reg_0112;
    67: op1_14_in00 = reg_0064;
    92: op1_14_in00 = reg_1505;
    93: op1_14_in00 = reg_0694;
    33: op1_14_in00 = imem07_in[11:8];
    94: op1_14_in00 = reg_1278;
    95: op1_14_in00 = reg_1323;
    96: op1_14_in00 = reg_1182;
    97: op1_14_in00 = reg_1006;
    98: op1_14_in00 = reg_0438;
    99: op1_14_in00 = reg_1107;
    28: op1_14_in00 = imem07_in[15:12];
    100: op1_14_in00 = reg_0254;
    101: op1_14_in00 = reg_1058;
    102: op1_14_in00 = reg_0238;
    103: op1_14_in00 = reg_1208;
    109: op1_14_in00 = reg_1208;
    104: op1_14_in00 = reg_0339;
    105: op1_14_in00 = reg_1420;
    106: op1_14_in00 = imem00_in[7:4];
    107: op1_14_in00 = reg_0899;
    37: op1_14_in00 = reg_0224;
    108: op1_14_in00 = reg_1334;
    110: op1_14_in00 = imem00_in[3:0];
    111: op1_14_in00 = reg_0630;
    112: op1_14_in00 = reg_0669;
    113: op1_14_in00 = reg_0334;
    114: op1_14_in00 = reg_0895;
    115: op1_14_in00 = reg_0395;
    116: op1_14_in00 = reg_0561;
    117: op1_14_in00 = reg_0536;
    118: op1_14_in00 = reg_0938;
    119: op1_14_in00 = reg_0299;
    47: op1_14_in00 = reg_0540;
    120: op1_14_in00 = reg_1244;
    121: op1_14_in00 = reg_0147;
    122: op1_14_in00 = imem00_in[15:12];
    123: op1_14_in00 = reg_0714;
    124: op1_14_in00 = reg_0750;
    125: op1_14_in00 = reg_0159;
    126: op1_14_in00 = reg_0426;
    127: op1_14_in00 = reg_0234;
    128: op1_14_in00 = reg_0963;
    129: op1_14_in00 = reg_0312;
    130: op1_14_in00 = reg_0423;
    default: op1_14_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_14_inv00 = 1;
    73: op1_14_inv00 = 1;
    55: op1_14_inv00 = 1;
    74: op1_14_inv00 = 1;
    54: op1_14_inv00 = 1;
    49: op1_14_inv00 = 1;
    69: op1_14_inv00 = 1;
    56: op1_14_inv00 = 1;
    76: op1_14_inv00 = 1;
    71: op1_14_inv00 = 1;
    87: op1_14_inv00 = 1;
    57: op1_14_inv00 = 1;
    78: op1_14_inv00 = 1;
    58: op1_14_inv00 = 1;
    70: op1_14_inv00 = 1;
    59: op1_14_inv00 = 1;
    79: op1_14_inv00 = 1;
    51: op1_14_inv00 = 1;
    62: op1_14_inv00 = 1;
    81: op1_14_inv00 = 1;
    82: op1_14_inv00 = 1;
    52: op1_14_inv00 = 1;
    63: op1_14_inv00 = 1;
    64: op1_14_inv00 = 1;
    83: op1_14_inv00 = 1;
    84: op1_14_inv00 = 1;
    65: op1_14_inv00 = 1;
    67: op1_14_inv00 = 1;
    92: op1_14_inv00 = 1;
    93: op1_14_inv00 = 1;
    95: op1_14_inv00 = 1;
    100: op1_14_inv00 = 1;
    101: op1_14_inv00 = 1;
    102: op1_14_inv00 = 1;
    37: op1_14_inv00 = 1;
    108: op1_14_inv00 = 1;
    110: op1_14_inv00 = 1;
    111: op1_14_inv00 = 1;
    113: op1_14_inv00 = 1;
    114: op1_14_inv00 = 1;
    115: op1_14_inv00 = 1;
    116: op1_14_inv00 = 1;
    118: op1_14_inv00 = 1;
    123: op1_14_inv00 = 1;
    124: op1_14_inv00 = 1;
    125: op1_14_inv00 = 1;
    126: op1_14_inv00 = 1;
    128: op1_14_inv00 = 1;
    130: op1_14_inv00 = 1;
    default: op1_14_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in01 = reg_0445;
    53: op1_14_in01 = reg_0832;
    73: op1_14_in01 = reg_0791;
    55: op1_14_in01 = reg_0869;
    108: op1_14_in01 = reg_0869;
    86: op1_14_in01 = reg_0823;
    74: op1_14_in01 = reg_0536;
    54: op1_14_in01 = reg_0488;
    75: op1_14_in01 = reg_0204;
    49: op1_14_in01 = reg_0931;
    69: op1_14_in01 = reg_0446;
    56: op1_14_in01 = reg_0891;
    50: op1_14_in01 = reg_0460;
    76: op1_14_in01 = reg_1510;
    71: op1_14_in01 = reg_0555;
    87: op1_14_in01 = reg_0559;
    57: op1_14_in01 = reg_0637;
    52: op1_14_in01 = reg_0637;
    68: op1_14_in01 = reg_0497;
    77: op1_14_in01 = reg_0412;
    61: op1_14_in01 = reg_1079;
    78: op1_14_in01 = reg_0736;
    58: op1_14_in01 = reg_0899;
    70: op1_14_in01 = reg_1000;
    64: op1_14_in01 = reg_1000;
    59: op1_14_in01 = reg_0305;
    79: op1_14_in01 = reg_0040;
    51: op1_14_in01 = reg_0743;
    60: op1_14_in01 = reg_0957;
    80: op1_14_in01 = reg_0905;
    88: op1_14_in01 = reg_0120;
    62: op1_14_in01 = imem07_in[11:8];
    81: op1_14_in01 = reg_0602;
    82: op1_14_in01 = reg_0474;
    63: op1_14_in01 = reg_1055;
    83: op1_14_in01 = reg_0868;
    89: op1_14_in01 = reg_1149;
    84: op1_14_in01 = imem05_in[3:0];
    85: op1_14_in01 = imem00_in[3:0];
    65: op1_14_in01 = reg_0696;
    90: op1_14_in01 = reg_0049;
    66: op1_14_in01 = reg_0967;
    48: op1_14_in01 = reg_0539;
    91: op1_14_in01 = reg_1243;
    46: op1_14_in01 = reg_0106;
    67: op1_14_in01 = reg_0034;
    92: op1_14_in01 = reg_0172;
    93: op1_14_in01 = reg_1203;
    33: op1_14_in01 = reg_0100;
    94: op1_14_in01 = reg_0803;
    95: op1_14_in01 = reg_0372;
    97: op1_14_in01 = reg_0009;
    98: op1_14_in01 = reg_0148;
    99: op1_14_in01 = reg_0021;
    100: op1_14_in01 = reg_1074;
    101: op1_14_in01 = reg_1334;
    102: op1_14_in01 = reg_0830;
    103: op1_14_in01 = reg_0458;
    104: op1_14_in01 = reg_0336;
    105: op1_14_in01 = reg_0265;
    106: op1_14_in01 = reg_0248;
    107: op1_14_in01 = reg_0292;
    37: op1_14_in01 = reg_0170;
    109: op1_14_in01 = reg_0884;
    110: op1_14_in01 = reg_0958;
    111: op1_14_in01 = reg_0697;
    112: op1_14_in01 = reg_1242;
    113: op1_14_in01 = reg_1402;
    114: op1_14_in01 = imem02_in[15:12];
    115: op1_14_in01 = reg_0648;
    116: op1_14_in01 = reg_0975;
    117: op1_14_in01 = reg_0064;
    118: op1_14_in01 = reg_0937;
    119: op1_14_in01 = reg_0140;
    47: op1_14_in01 = reg_0541;
    120: op1_14_in01 = reg_0926;
    121: op1_14_in01 = reg_0146;
    122: op1_14_in01 = reg_0866;
    123: op1_14_in01 = reg_1303;
    124: op1_14_in01 = reg_0025;
    125: op1_14_in01 = reg_0661;
    126: op1_14_in01 = reg_1216;
    127: op1_14_in01 = reg_0375;
    128: op1_14_in01 = reg_0363;
    129: op1_14_in01 = reg_0144;
    130: op1_14_in01 = reg_0254;
    default: op1_14_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    75: op1_14_inv01 = 1;
    71: op1_14_inv01 = 1;
    57: op1_14_inv01 = 1;
    68: op1_14_inv01 = 1;
    77: op1_14_inv01 = 1;
    78: op1_14_inv01 = 1;
    58: op1_14_inv01 = 1;
    70: op1_14_inv01 = 1;
    59: op1_14_inv01 = 1;
    79: op1_14_inv01 = 1;
    51: op1_14_inv01 = 1;
    80: op1_14_inv01 = 1;
    88: op1_14_inv01 = 1;
    62: op1_14_inv01 = 1;
    81: op1_14_inv01 = 1;
    63: op1_14_inv01 = 1;
    64: op1_14_inv01 = 1;
    89: op1_14_inv01 = 1;
    84: op1_14_inv01 = 1;
    65: op1_14_inv01 = 1;
    48: op1_14_inv01 = 1;
    91: op1_14_inv01 = 1;
    46: op1_14_inv01 = 1;
    92: op1_14_inv01 = 1;
    95: op1_14_inv01 = 1;
    97: op1_14_inv01 = 1;
    99: op1_14_inv01 = 1;
    101: op1_14_inv01 = 1;
    102: op1_14_inv01 = 1;
    106: op1_14_inv01 = 1;
    37: op1_14_inv01 = 1;
    108: op1_14_inv01 = 1;
    110: op1_14_inv01 = 1;
    113: op1_14_inv01 = 1;
    114: op1_14_inv01 = 1;
    115: op1_14_inv01 = 1;
    117: op1_14_inv01 = 1;
    118: op1_14_inv01 = 1;
    119: op1_14_inv01 = 1;
    121: op1_14_inv01 = 1;
    122: op1_14_inv01 = 1;
    125: op1_14_inv01 = 1;
    127: op1_14_inv01 = 1;
    128: op1_14_inv01 = 1;
    default: op1_14_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in02 = reg_1277;
    53: op1_14_in02 = imem05_in[11:8];
    73: op1_14_in02 = reg_1078;
    55: op1_14_in02 = reg_0141;
    123: op1_14_in02 = reg_0141;
    86: op1_14_in02 = reg_0989;
    74: op1_14_in02 = reg_0397;
    54: op1_14_in02 = reg_0836;
    75: op1_14_in02 = reg_0877;
    49: op1_14_in02 = reg_0133;
    69: op1_14_in02 = reg_0699;
    87: op1_14_in02 = reg_0699;
    56: op1_14_in02 = reg_1199;
    50: op1_14_in02 = reg_0268;
    76: op1_14_in02 = reg_1080;
    61: op1_14_in02 = reg_1080;
    71: op1_14_in02 = reg_0748;
    120: op1_14_in02 = reg_0748;
    57: op1_14_in02 = reg_0263;
    68: op1_14_in02 = reg_0981;
    77: op1_14_in02 = reg_0406;
    78: op1_14_in02 = reg_0579;
    58: op1_14_in02 = reg_0290;
    98: op1_14_in02 = reg_0290;
    70: op1_14_in02 = reg_1003;
    59: op1_14_in02 = reg_0319;
    79: op1_14_in02 = reg_0014;
    51: op1_14_in02 = reg_0982;
    60: op1_14_in02 = reg_0597;
    80: op1_14_in02 = reg_1334;
    88: op1_14_in02 = reg_1071;
    62: op1_14_in02 = reg_0245;
    81: op1_14_in02 = reg_0797;
    82: op1_14_in02 = reg_0971;
    52: op1_14_in02 = reg_0586;
    63: op1_14_in02 = reg_1183;
    64: op1_14_in02 = reg_1001;
    83: op1_14_in02 = reg_0616;
    89: op1_14_in02 = reg_0481;
    84: op1_14_in02 = reg_0604;
    85: op1_14_in02 = reg_0907;
    65: op1_14_in02 = reg_0194;
    90: op1_14_in02 = reg_1448;
    66: op1_14_in02 = reg_0726;
    48: op1_14_in02 = reg_0302;
    91: op1_14_in02 = reg_0445;
    46: op1_14_in02 = reg_0380;
    67: op1_14_in02 = reg_0799;
    92: op1_14_in02 = reg_0372;
    93: op1_14_in02 = reg_1233;
    33: op1_14_in02 = reg_0518;
    94: op1_14_in02 = reg_0615;
    95: op1_14_in02 = reg_0717;
    97: op1_14_in02 = reg_0227;
    99: op1_14_in02 = reg_0370;
    100: op1_14_in02 = reg_0432;
    101: op1_14_in02 = reg_1420;
    102: op1_14_in02 = reg_0439;
    103: op1_14_in02 = reg_0707;
    104: op1_14_in02 = reg_1237;
    105: op1_14_in02 = reg_1302;
    106: op1_14_in02 = reg_0725;
    107: op1_14_in02 = reg_0080;
    37: op1_14_in02 = reg_0298;
    108: op1_14_in02 = reg_0827;
    109: op1_14_in02 = reg_1149;
    110: op1_14_in02 = reg_1101;
    111: op1_14_in02 = reg_1402;
    112: op1_14_in02 = reg_0843;
    113: op1_14_in02 = reg_0939;
    114: op1_14_in02 = reg_0668;
    115: op1_14_in02 = reg_1181;
    116: op1_14_in02 = reg_1493;
    130: op1_14_in02 = reg_1493;
    117: op1_14_in02 = reg_1502;
    118: op1_14_in02 = reg_1514;
    119: op1_14_in02 = reg_0309;
    47: op1_14_in02 = reg_0418;
    121: op1_14_in02 = reg_1511;
    122: op1_14_in02 = reg_1081;
    124: op1_14_in02 = reg_0425;
    125: op1_14_in02 = reg_0286;
    126: op1_14_in02 = reg_0129;
    127: op1_14_in02 = reg_1494;
    129: op1_14_in02 = reg_1494;
    128: op1_14_in02 = reg_0901;
    default: op1_14_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv02 = 1;
    73: op1_14_inv02 = 1;
    54: op1_14_inv02 = 1;
    75: op1_14_inv02 = 1;
    69: op1_14_inv02 = 1;
    56: op1_14_inv02 = 1;
    76: op1_14_inv02 = 1;
    71: op1_14_inv02 = 1;
    87: op1_14_inv02 = 1;
    77: op1_14_inv02 = 1;
    78: op1_14_inv02 = 1;
    58: op1_14_inv02 = 1;
    59: op1_14_inv02 = 1;
    88: op1_14_inv02 = 1;
    62: op1_14_inv02 = 1;
    82: op1_14_inv02 = 1;
    83: op1_14_inv02 = 1;
    84: op1_14_inv02 = 1;
    85: op1_14_inv02 = 1;
    66: op1_14_inv02 = 1;
    48: op1_14_inv02 = 1;
    93: op1_14_inv02 = 1;
    94: op1_14_inv02 = 1;
    95: op1_14_inv02 = 1;
    97: op1_14_inv02 = 1;
    98: op1_14_inv02 = 1;
    99: op1_14_inv02 = 1;
    100: op1_14_inv02 = 1;
    102: op1_14_inv02 = 1;
    103: op1_14_inv02 = 1;
    105: op1_14_inv02 = 1;
    37: op1_14_inv02 = 1;
    109: op1_14_inv02 = 1;
    110: op1_14_inv02 = 1;
    113: op1_14_inv02 = 1;
    114: op1_14_inv02 = 1;
    116: op1_14_inv02 = 1;
    119: op1_14_inv02 = 1;
    47: op1_14_inv02 = 1;
    120: op1_14_inv02 = 1;
    122: op1_14_inv02 = 1;
    123: op1_14_inv02 = 1;
    124: op1_14_inv02 = 1;
    125: op1_14_inv02 = 1;
    127: op1_14_inv02 = 1;
    129: op1_14_inv02 = 1;
    130: op1_14_inv02 = 1;
    default: op1_14_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in03 = reg_0841;
    53: op1_14_in03 = reg_0174;
    73: op1_14_in03 = imem00_in[15:12];
    55: op1_14_in03 = reg_0399;
    86: op1_14_in03 = reg_1314;
    74: op1_14_in03 = reg_0869;
    54: op1_14_in03 = reg_0719;
    75: op1_14_in03 = reg_1164;
    49: op1_14_in03 = reg_0141;
    69: op1_14_in03 = reg_1140;
    56: op1_14_in03 = reg_0178;
    50: op1_14_in03 = reg_0230;
    76: op1_14_in03 = reg_0350;
    71: op1_14_in03 = reg_0445;
    87: op1_14_in03 = reg_0444;
    57: op1_14_in03 = reg_0568;
    123: op1_14_in03 = reg_0568;
    68: op1_14_in03 = reg_0256;
    77: op1_14_in03 = reg_0094;
    61: op1_14_in03 = reg_0155;
    78: op1_14_in03 = reg_1431;
    58: op1_14_in03 = reg_0088;
    70: op1_14_in03 = reg_0314;
    59: op1_14_in03 = reg_0862;
    79: op1_14_in03 = reg_1435;
    51: op1_14_in03 = reg_0819;
    60: op1_14_in03 = imem03_in[11:8];
    80: op1_14_in03 = reg_1323;
    88: op1_14_in03 = imem02_in[3:0];
    62: op1_14_in03 = reg_0489;
    81: op1_14_in03 = reg_0039;
    82: op1_14_in03 = reg_0973;
    52: op1_14_in03 = reg_0526;
    63: op1_14_in03 = reg_0186;
    64: op1_14_in03 = reg_0962;
    83: op1_14_in03 = reg_1281;
    89: op1_14_in03 = reg_0025;
    84: op1_14_in03 = reg_0392;
    85: op1_14_in03 = reg_0615;
    65: op1_14_in03 = reg_0374;
    108: op1_14_in03 = reg_0374;
    90: op1_14_in03 = reg_1033;
    66: op1_14_in03 = reg_0400;
    128: op1_14_in03 = reg_0400;
    48: op1_14_in03 = reg_0300;
    91: op1_14_in03 = reg_1490;
    122: op1_14_in03 = reg_1490;
    46: op1_14_in03 = reg_0900;
    67: op1_14_in03 = reg_0737;
    92: op1_14_in03 = reg_0109;
    93: op1_14_in03 = reg_1082;
    33: op1_14_in03 = reg_0521;
    94: op1_14_in03 = reg_0554;
    112: op1_14_in03 = reg_0554;
    95: op1_14_in03 = reg_0637;
    97: op1_14_in03 = reg_0006;
    98: op1_14_in03 = reg_0464;
    99: op1_14_in03 = reg_0315;
    100: op1_14_in03 = reg_0436;
    101: op1_14_in03 = reg_0696;
    102: op1_14_in03 = reg_0438;
    103: op1_14_in03 = reg_1009;
    104: op1_14_in03 = reg_0536;
    105: op1_14_in03 = reg_0584;
    106: op1_14_in03 = reg_1491;
    107: op1_14_in03 = reg_0079;
    37: op1_14_in03 = reg_0299;
    109: op1_14_in03 = reg_0707;
    110: op1_14_in03 = reg_1277;
    111: op1_14_in03 = reg_1404;
    113: op1_14_in03 = reg_0792;
    114: op1_14_in03 = reg_0889;
    115: op1_14_in03 = reg_1401;
    116: op1_14_in03 = reg_0532;
    117: op1_14_in03 = reg_0210;
    118: op1_14_in03 = reg_0303;
    119: op1_14_in03 = reg_0139;
    47: op1_14_in03 = reg_0873;
    120: op1_14_in03 = reg_1489;
    121: op1_14_in03 = reg_0384;
    124: op1_14_in03 = reg_0208;
    125: op1_14_in03 = reg_0739;
    126: op1_14_in03 = reg_0337;
    127: op1_14_in03 = reg_1184;
    129: op1_14_in03 = reg_0556;
    130: op1_14_in03 = reg_0744;
    default: op1_14_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv03 = 1;
    55: op1_14_inv03 = 1;
    74: op1_14_inv03 = 1;
    75: op1_14_inv03 = 1;
    69: op1_14_inv03 = 1;
    56: op1_14_inv03 = 1;
    50: op1_14_inv03 = 1;
    71: op1_14_inv03 = 1;
    87: op1_14_inv03 = 1;
    68: op1_14_inv03 = 1;
    77: op1_14_inv03 = 1;
    61: op1_14_inv03 = 1;
    78: op1_14_inv03 = 1;
    70: op1_14_inv03 = 1;
    60: op1_14_inv03 = 1;
    62: op1_14_inv03 = 1;
    82: op1_14_inv03 = 1;
    63: op1_14_inv03 = 1;
    64: op1_14_inv03 = 1;
    89: op1_14_inv03 = 1;
    85: op1_14_inv03 = 1;
    65: op1_14_inv03 = 1;
    66: op1_14_inv03 = 1;
    91: op1_14_inv03 = 1;
    67: op1_14_inv03 = 1;
    93: op1_14_inv03 = 1;
    33: op1_14_inv03 = 1;
    94: op1_14_inv03 = 1;
    95: op1_14_inv03 = 1;
    99: op1_14_inv03 = 1;
    101: op1_14_inv03 = 1;
    102: op1_14_inv03 = 1;
    103: op1_14_inv03 = 1;
    104: op1_14_inv03 = 1;
    37: op1_14_inv03 = 1;
    111: op1_14_inv03 = 1;
    113: op1_14_inv03 = 1;
    114: op1_14_inv03 = 1;
    115: op1_14_inv03 = 1;
    119: op1_14_inv03 = 1;
    47: op1_14_inv03 = 1;
    120: op1_14_inv03 = 1;
    121: op1_14_inv03 = 1;
    122: op1_14_inv03 = 1;
    123: op1_14_inv03 = 1;
    125: op1_14_inv03 = 1;
    128: op1_14_inv03 = 1;
    130: op1_14_inv03 = 1;
    default: op1_14_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in04 = imem00_in[15:12];
    53: op1_14_in04 = reg_0996;
    73: op1_14_in04 = reg_0350;
    55: op1_14_in04 = reg_0115;
    86: op1_14_in04 = reg_0246;
    74: op1_14_in04 = reg_1323;
    54: op1_14_in04 = reg_0129;
    75: op1_14_in04 = reg_1163;
    49: op1_14_in04 = reg_0822;
    116: op1_14_in04 = reg_0822;
    69: op1_14_in04 = reg_1029;
    56: op1_14_in04 = reg_0104;
    50: op1_14_in04 = imem07_in[11:8];
    76: op1_14_in04 = reg_1028;
    71: op1_14_in04 = reg_0824;
    87: op1_14_in04 = reg_1425;
    57: op1_14_in04 = reg_0171;
    68: op1_14_in04 = reg_1207;
    77: op1_14_in04 = reg_0452;
    61: op1_14_in04 = reg_0172;
    78: op1_14_in04 = reg_0832;
    58: op1_14_in04 = reg_0012;
    70: op1_14_in04 = reg_0952;
    59: op1_14_in04 = reg_0835;
    79: op1_14_in04 = reg_0908;
    51: op1_14_in04 = reg_0439;
    60: op1_14_in04 = reg_1093;
    80: op1_14_in04 = imem06_in[11:8];
    88: op1_14_in04 = reg_0530;
    62: op1_14_in04 = reg_0224;
    119: op1_14_in04 = reg_0224;
    81: op1_14_in04 = reg_0014;
    82: op1_14_in04 = reg_1450;
    52: op1_14_in04 = reg_0295;
    63: op1_14_in04 = reg_0667;
    64: op1_14_in04 = reg_1301;
    83: op1_14_in04 = reg_1278;
    89: op1_14_in04 = reg_0427;
    84: op1_14_in04 = reg_0491;
    85: op1_14_in04 = reg_0580;
    65: op1_14_in04 = reg_0584;
    90: op1_14_in04 = reg_1001;
    66: op1_14_in04 = reg_0384;
    48: op1_14_in04 = reg_0184;
    91: op1_14_in04 = reg_0615;
    46: op1_14_in04 = reg_0705;
    67: op1_14_in04 = reg_0702;
    92: op1_14_in04 = reg_0714;
    93: op1_14_in04 = reg_0340;
    33: op1_14_in04 = reg_0483;
    94: op1_14_in04 = reg_0640;
    95: op1_14_in04 = reg_0585;
    108: op1_14_in04 = reg_0585;
    97: op1_14_in04 = reg_0504;
    98: op1_14_in04 = reg_0335;
    99: op1_14_in04 = reg_0735;
    100: op1_14_in04 = reg_0971;
    101: op1_14_in04 = reg_1326;
    102: op1_14_in04 = reg_1456;
    103: op1_14_in04 = reg_0348;
    104: op1_14_in04 = reg_1503;
    105: op1_14_in04 = reg_0622;
    106: op1_14_in04 = reg_1053;
    107: op1_14_in04 = reg_0403;
    37: op1_14_in04 = reg_0159;
    109: op1_14_in04 = reg_1009;
    110: op1_14_in04 = reg_0501;
    111: op1_14_in04 = reg_0940;
    112: op1_14_in04 = reg_0486;
    113: op1_14_in04 = reg_0888;
    114: op1_14_in04 = reg_0423;
    115: op1_14_in04 = reg_0477;
    117: op1_14_in04 = reg_0035;
    118: op1_14_in04 = reg_0450;
    47: op1_14_in04 = reg_0168;
    120: op1_14_in04 = reg_0804;
    121: op1_14_in04 = reg_0360;
    122: op1_14_in04 = reg_0841;
    123: op1_14_in04 = reg_0571;
    124: op1_14_in04 = imem04_in[7:4];
    125: op1_14_in04 = reg_0413;
    126: op1_14_in04 = reg_1257;
    127: op1_14_in04 = reg_0964;
    128: op1_14_in04 = reg_0292;
    129: op1_14_in04 = reg_0070;
    130: op1_14_in04 = reg_0532;
    default: op1_14_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_14_inv04 = 1;
    56: op1_14_inv04 = 1;
    79: op1_14_inv04 = 1;
    51: op1_14_inv04 = 1;
    60: op1_14_inv04 = 1;
    88: op1_14_inv04 = 1;
    62: op1_14_inv04 = 1;
    81: op1_14_inv04 = 1;
    82: op1_14_inv04 = 1;
    83: op1_14_inv04 = 1;
    89: op1_14_inv04 = 1;
    65: op1_14_inv04 = 1;
    48: op1_14_inv04 = 1;
    46: op1_14_inv04 = 1;
    67: op1_14_inv04 = 1;
    93: op1_14_inv04 = 1;
    94: op1_14_inv04 = 1;
    95: op1_14_inv04 = 1;
    99: op1_14_inv04 = 1;
    101: op1_14_inv04 = 1;
    103: op1_14_inv04 = 1;
    105: op1_14_inv04 = 1;
    106: op1_14_inv04 = 1;
    107: op1_14_inv04 = 1;
    37: op1_14_inv04 = 1;
    108: op1_14_inv04 = 1;
    109: op1_14_inv04 = 1;
    110: op1_14_inv04 = 1;
    111: op1_14_inv04 = 1;
    113: op1_14_inv04 = 1;
    115: op1_14_inv04 = 1;
    116: op1_14_inv04 = 1;
    119: op1_14_inv04 = 1;
    47: op1_14_inv04 = 1;
    120: op1_14_inv04 = 1;
    124: op1_14_inv04 = 1;
    125: op1_14_inv04 = 1;
    127: op1_14_inv04 = 1;
    128: op1_14_inv04 = 1;
    129: op1_14_inv04 = 1;
    default: op1_14_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in05 = reg_0523;
    120: op1_14_in05 = reg_0523;
    53: op1_14_in05 = reg_0992;
    73: op1_14_in05 = reg_1230;
    55: op1_14_in05 = reg_0116;
    86: op1_14_in05 = reg_1300;
    70: op1_14_in05 = reg_1300;
    74: op1_14_in05 = reg_0752;
    54: op1_14_in05 = reg_0034;
    75: op1_14_in05 = reg_0066;
    49: op1_14_in05 = reg_0827;
    69: op1_14_in05 = reg_1018;
    56: op1_14_in05 = reg_0479;
    50: op1_14_in05 = reg_0994;
    76: op1_14_in05 = reg_0887;
    71: op1_14_in05 = reg_1278;
    87: op1_14_in05 = reg_0707;
    57: op1_14_in05 = reg_0371;
    68: op1_14_in05 = reg_0970;
    77: op1_14_in05 = reg_0537;
    61: op1_14_in05 = reg_1227;
    78: op1_14_in05 = reg_0702;
    58: op1_14_in05 = reg_0010;
    59: op1_14_in05 = reg_0020;
    79: op1_14_in05 = reg_0960;
    51: op1_14_in05 = reg_0438;
    60: op1_14_in05 = reg_0113;
    80: op1_14_in05 = imem06_in[15:12];
    88: op1_14_in05 = reg_0934;
    62: op1_14_in05 = reg_1094;
    119: op1_14_in05 = reg_1094;
    81: op1_14_in05 = reg_0751;
    82: op1_14_in05 = reg_0112;
    52: op1_14_in05 = reg_0419;
    63: op1_14_in05 = reg_0922;
    64: op1_14_in05 = reg_1231;
    83: op1_14_in05 = reg_1490;
    89: op1_14_in05 = reg_0443;
    84: op1_14_in05 = reg_1104;
    85: op1_14_in05 = reg_1053;
    65: op1_14_in05 = reg_0244;
    90: op1_14_in05 = reg_0783;
    66: op1_14_in05 = reg_0365;
    48: op1_14_in05 = reg_0118;
    91: op1_14_in05 = reg_1052;
    46: op1_14_in05 = reg_0307;
    67: op1_14_in05 = reg_0833;
    92: op1_14_in05 = reg_0529;
    93: op1_14_in05 = reg_0262;
    94: op1_14_in05 = reg_0293;
    95: op1_14_in05 = reg_0526;
    97: op1_14_in05 = reg_1000;
    98: op1_14_in05 = reg_0013;
    99: op1_14_in05 = reg_0136;
    100: op1_14_in05 = reg_0972;
    101: op1_14_in05 = imem06_in[11:8];
    102: op1_14_in05 = reg_1511;
    103: op1_14_in05 = reg_0425;
    104: op1_14_in05 = reg_0035;
    105: op1_14_in05 = reg_1228;
    106: op1_14_in05 = reg_0221;
    107: op1_14_in05 = reg_0634;
    128: op1_14_in05 = reg_0634;
    37: op1_14_in05 = reg_0156;
    108: op1_14_in05 = reg_0568;
    109: op1_14_in05 = reg_0218;
    110: op1_14_in05 = reg_0613;
    111: op1_14_in05 = reg_0938;
    112: op1_14_in05 = reg_1028;
    113: op1_14_in05 = reg_0601;
    114: op1_14_in05 = reg_0056;
    115: op1_14_in05 = reg_0888;
    116: op1_14_in05 = reg_0390;
    117: op1_14_in05 = reg_1168;
    118: op1_14_in05 = reg_0197;
    47: op1_14_in05 = reg_0192;
    121: op1_14_in05 = reg_0901;
    122: op1_14_in05 = reg_0616;
    123: op1_14_in05 = reg_0569;
    124: op1_14_in05 = reg_0252;
    125: op1_14_in05 = reg_0620;
    126: op1_14_in05 = reg_0531;
    127: op1_14_in05 = reg_1314;
    129: op1_14_in05 = reg_0349;
    130: op1_14_in05 = reg_0533;
    default: op1_14_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_14_inv05 = 1;
    73: op1_14_inv05 = 1;
    86: op1_14_inv05 = 1;
    74: op1_14_inv05 = 1;
    75: op1_14_inv05 = 1;
    69: op1_14_inv05 = 1;
    50: op1_14_inv05 = 1;
    87: op1_14_inv05 = 1;
    68: op1_14_inv05 = 1;
    61: op1_14_inv05 = 1;
    78: op1_14_inv05 = 1;
    58: op1_14_inv05 = 1;
    70: op1_14_inv05 = 1;
    59: op1_14_inv05 = 1;
    80: op1_14_inv05 = 1;
    88: op1_14_inv05 = 1;
    62: op1_14_inv05 = 1;
    82: op1_14_inv05 = 1;
    63: op1_14_inv05 = 1;
    64: op1_14_inv05 = 1;
    83: op1_14_inv05 = 1;
    89: op1_14_inv05 = 1;
    85: op1_14_inv05 = 1;
    90: op1_14_inv05 = 1;
    66: op1_14_inv05 = 1;
    91: op1_14_inv05 = 1;
    46: op1_14_inv05 = 1;
    92: op1_14_inv05 = 1;
    97: op1_14_inv05 = 1;
    98: op1_14_inv05 = 1;
    99: op1_14_inv05 = 1;
    102: op1_14_inv05 = 1;
    106: op1_14_inv05 = 1;
    107: op1_14_inv05 = 1;
    37: op1_14_inv05 = 1;
    108: op1_14_inv05 = 1;
    110: op1_14_inv05 = 1;
    111: op1_14_inv05 = 1;
    113: op1_14_inv05 = 1;
    114: op1_14_inv05 = 1;
    115: op1_14_inv05 = 1;
    116: op1_14_inv05 = 1;
    117: op1_14_inv05 = 1;
    118: op1_14_inv05 = 1;
    119: op1_14_inv05 = 1;
    120: op1_14_inv05 = 1;
    123: op1_14_inv05 = 1;
    125: op1_14_inv05 = 1;
    127: op1_14_inv05 = 1;
    default: op1_14_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in06 = reg_1229;
    53: op1_14_in06 = reg_0182;
    73: op1_14_in06 = reg_0987;
    55: op1_14_in06 = reg_0716;
    86: op1_14_in06 = reg_1226;
    74: op1_14_in06 = imem06_in[11:8];
    81: op1_14_in06 = imem06_in[11:8];
    54: op1_14_in06 = reg_0175;
    75: op1_14_in06 = reg_0333;
    49: op1_14_in06 = reg_0115;
    80: op1_14_in06 = reg_0115;
    69: op1_14_in06 = reg_0254;
    56: op1_14_in06 = reg_0840;
    50: op1_14_in06 = reg_0226;
    76: op1_14_in06 = reg_0188;
    71: op1_14_in06 = reg_1080;
    87: op1_14_in06 = reg_0541;
    57: op1_14_in06 = reg_0067;
    68: op1_14_in06 = reg_0973;
    77: op1_14_in06 = reg_0596;
    61: op1_14_in06 = reg_1201;
    78: op1_14_in06 = reg_0992;
    58: op1_14_in06 = reg_0486;
    70: op1_14_in06 = reg_0558;
    59: op1_14_in06 = reg_0033;
    79: op1_14_in06 = reg_1323;
    51: op1_14_in06 = reg_0402;
    60: op1_14_in06 = reg_0478;
    88: op1_14_in06 = reg_0981;
    62: op1_14_in06 = reg_0777;
    82: op1_14_in06 = reg_0379;
    52: op1_14_in06 = reg_0459;
    63: op1_14_in06 = reg_0310;
    64: op1_14_in06 = reg_1208;
    83: op1_14_in06 = reg_1244;
    89: op1_14_in06 = reg_1384;
    84: op1_14_in06 = reg_0630;
    85: op1_14_in06 = reg_1052;
    65: op1_14_in06 = reg_1202;
    90: op1_14_in06 = reg_0600;
    66: op1_14_in06 = reg_0047;
    48: op1_14_in06 = reg_0275;
    91: op1_14_in06 = reg_0293;
    46: op1_14_in06 = reg_0876;
    67: op1_14_in06 = reg_1259;
    92: op1_14_in06 = reg_0323;
    93: op1_14_in06 = reg_0904;
    94: op1_14_in06 = reg_1027;
    122: op1_14_in06 = reg_1027;
    95: op1_14_in06 = reg_0583;
    123: op1_14_in06 = reg_0583;
    97: op1_14_in06 = reg_0154;
    98: op1_14_in06 = reg_0895;
    99: op1_14_in06 = reg_0205;
    100: op1_14_in06 = reg_0127;
    101: op1_14_in06 = reg_0619;
    102: op1_14_in06 = reg_0362;
    103: op1_14_in06 = imem04_in[7:4];
    104: op1_14_in06 = reg_0708;
    105: op1_14_in06 = reg_1225;
    106: op1_14_in06 = reg_0883;
    107: op1_14_in06 = reg_1002;
    37: op1_14_in06 = reg_0031;
    108: op1_14_in06 = reg_0571;
    109: op1_14_in06 = reg_1325;
    110: op1_14_in06 = reg_0615;
    111: op1_14_in06 = reg_0197;
    112: op1_14_in06 = reg_0221;
    113: op1_14_in06 = reg_0274;
    114: op1_14_in06 = reg_0712;
    115: op1_14_in06 = reg_0601;
    118: op1_14_in06 = reg_0601;
    116: op1_14_in06 = reg_0433;
    117: op1_14_in06 = reg_0040;
    119: op1_14_in06 = reg_0661;
    47: op1_14_in06 = reg_0729;
    120: op1_14_in06 = reg_1230;
    121: op1_14_in06 = reg_0162;
    124: op1_14_in06 = reg_1216;
    125: op1_14_in06 = reg_0593;
    126: op1_14_in06 = reg_0297;
    127: op1_14_in06 = reg_0957;
    128: op1_14_in06 = reg_1068;
    129: op1_14_in06 = reg_1314;
    130: op1_14_in06 = reg_0326;
    default: op1_14_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv06 = 1;
    74: op1_14_inv06 = 1;
    54: op1_14_inv06 = 1;
    49: op1_14_inv06 = 1;
    69: op1_14_inv06 = 1;
    56: op1_14_inv06 = 1;
    76: op1_14_inv06 = 1;
    71: op1_14_inv06 = 1;
    57: op1_14_inv06 = 1;
    68: op1_14_inv06 = 1;
    77: op1_14_inv06 = 1;
    78: op1_14_inv06 = 1;
    70: op1_14_inv06 = 1;
    79: op1_14_inv06 = 1;
    51: op1_14_inv06 = 1;
    60: op1_14_inv06 = 1;
    88: op1_14_inv06 = 1;
    62: op1_14_inv06 = 1;
    63: op1_14_inv06 = 1;
    64: op1_14_inv06 = 1;
    89: op1_14_inv06 = 1;
    85: op1_14_inv06 = 1;
    65: op1_14_inv06 = 1;
    90: op1_14_inv06 = 1;
    46: op1_14_inv06 = 1;
    67: op1_14_inv06 = 1;
    97: op1_14_inv06 = 1;
    98: op1_14_inv06 = 1;
    99: op1_14_inv06 = 1;
    100: op1_14_inv06 = 1;
    101: op1_14_inv06 = 1;
    102: op1_14_inv06 = 1;
    103: op1_14_inv06 = 1;
    105: op1_14_inv06 = 1;
    106: op1_14_inv06 = 1;
    107: op1_14_inv06 = 1;
    109: op1_14_inv06 = 1;
    110: op1_14_inv06 = 1;
    111: op1_14_inv06 = 1;
    114: op1_14_inv06 = 1;
    118: op1_14_inv06 = 1;
    120: op1_14_inv06 = 1;
    122: op1_14_inv06 = 1;
    123: op1_14_inv06 = 1;
    124: op1_14_inv06 = 1;
    127: op1_14_inv06 = 1;
    128: op1_14_inv06 = 1;
    129: op1_14_inv06 = 1;
    default: op1_14_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in07 = reg_0987;
    53: op1_14_in07 = reg_0317;
    73: op1_14_in07 = reg_1205;
    120: op1_14_in07 = reg_1205;
    55: op1_14_in07 = reg_0718;
    49: op1_14_in07 = reg_0718;
    86: op1_14_in07 = reg_0882;
    74: op1_14_in07 = reg_0984;
    54: op1_14_in07 = reg_0831;
    75: op1_14_in07 = reg_0045;
    69: op1_14_in07 = reg_0326;
    56: op1_14_in07 = reg_0426;
    50: op1_14_in07 = reg_0186;
    76: op1_14_in07 = reg_0201;
    71: op1_14_in07 = reg_0841;
    87: op1_14_in07 = reg_0000;
    57: op1_14_in07 = reg_0215;
    68: op1_14_in07 = reg_0935;
    77: op1_14_in07 = reg_0369;
    61: op1_14_in07 = reg_0203;
    78: op1_14_in07 = reg_0131;
    58: op1_14_in07 = reg_0742;
    70: op1_14_in07 = reg_1231;
    59: op1_14_in07 = reg_0792;
    79: op1_14_in07 = reg_0752;
    51: op1_14_in07 = reg_0384;
    60: op1_14_in07 = reg_0840;
    80: op1_14_in07 = reg_0716;
    88: op1_14_in07 = reg_0432;
    62: op1_14_in07 = reg_0031;
    81: op1_14_in07 = reg_1435;
    82: op1_14_in07 = reg_0802;
    52: op1_14_in07 = reg_0213;
    63: op1_14_in07 = reg_0297;
    64: op1_14_in07 = reg_0104;
    83: op1_14_in07 = reg_1242;
    89: op1_14_in07 = reg_0088;
    84: op1_14_in07 = reg_1404;
    85: op1_14_in07 = reg_0523;
    65: op1_14_in07 = reg_0191;
    90: op1_14_in07 = reg_0143;
    66: op1_14_in07 = reg_0092;
    48: op1_14_in07 = reg_0039;
    91: op1_14_in07 = reg_1028;
    46: op1_14_in07 = reg_0878;
    67: op1_14_in07 = reg_0996;
    92: op1_14_in07 = reg_0165;
    93: op1_14_in07 = reg_0420;
    94: op1_14_in07 = reg_0485;
    122: op1_14_in07 = reg_0485;
    95: op1_14_in07 = reg_1202;
    97: op1_14_in07 = reg_1447;
    98: op1_14_in07 = reg_0668;
    99: op1_14_in07 = reg_0701;
    100: op1_14_in07 = reg_0105;
    101: op1_14_in07 = reg_0132;
    102: op1_14_in07 = reg_0091;
    103: op1_14_in07 = reg_0493;
    104: op1_14_in07 = reg_0367;
    105: op1_14_in07 = reg_0308;
    106: op1_14_in07 = reg_0886;
    107: op1_14_in07 = reg_0626;
    37: op1_14_in07 = reg_0465;
    108: op1_14_in07 = reg_1225;
    109: op1_14_in07 = reg_1280;
    110: op1_14_in07 = reg_0616;
    111: op1_14_in07 = reg_0492;
    112: op1_14_in07 = reg_0249;
    113: op1_14_in07 = reg_0130;
    114: op1_14_in07 = reg_0532;
    115: op1_14_in07 = reg_0274;
    116: op1_14_in07 = reg_0429;
    117: op1_14_in07 = reg_0793;
    118: op1_14_in07 = reg_0449;
    119: op1_14_in07 = reg_0664;
    47: op1_14_in07 = imem06_in[7:4];
    121: op1_14_in07 = reg_0041;
    123: op1_14_in07 = reg_0067;
    124: op1_14_in07 = reg_0032;
    125: op1_14_in07 = reg_0592;
    126: op1_14_in07 = reg_1214;
    127: op1_14_in07 = reg_0329;
    128: op1_14_in07 = reg_0895;
    129: op1_14_in07 = reg_0756;
    130: op1_14_in07 = reg_0970;
    default: op1_14_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv07 = 1;
    73: op1_14_inv07 = 1;
    86: op1_14_inv07 = 1;
    54: op1_14_inv07 = 1;
    87: op1_14_inv07 = 1;
    68: op1_14_inv07 = 1;
    61: op1_14_inv07 = 1;
    78: op1_14_inv07 = 1;
    70: op1_14_inv07 = 1;
    59: op1_14_inv07 = 1;
    51: op1_14_inv07 = 1;
    60: op1_14_inv07 = 1;
    88: op1_14_inv07 = 1;
    81: op1_14_inv07 = 1;
    82: op1_14_inv07 = 1;
    63: op1_14_inv07 = 1;
    83: op1_14_inv07 = 1;
    89: op1_14_inv07 = 1;
    85: op1_14_inv07 = 1;
    90: op1_14_inv07 = 1;
    91: op1_14_inv07 = 1;
    67: op1_14_inv07 = 1;
    95: op1_14_inv07 = 1;
    98: op1_14_inv07 = 1;
    100: op1_14_inv07 = 1;
    102: op1_14_inv07 = 1;
    103: op1_14_inv07 = 1;
    104: op1_14_inv07 = 1;
    105: op1_14_inv07 = 1;
    37: op1_14_inv07 = 1;
    111: op1_14_inv07 = 1;
    114: op1_14_inv07 = 1;
    116: op1_14_inv07 = 1;
    118: op1_14_inv07 = 1;
    47: op1_14_inv07 = 1;
    120: op1_14_inv07 = 1;
    122: op1_14_inv07 = 1;
    123: op1_14_inv07 = 1;
    124: op1_14_inv07 = 1;
    130: op1_14_inv07 = 1;
    default: op1_14_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in08 = reg_0460;
    73: op1_14_in08 = reg_0460;
    53: op1_14_in08 = reg_0541;
    55: op1_14_in08 = reg_0619;
    86: op1_14_in08 = reg_0480;
    74: op1_14_in08 = reg_0669;
    54: op1_14_in08 = reg_1163;
    75: op1_14_in08 = reg_0940;
    49: op1_14_in08 = reg_0714;
    69: op1_14_in08 = reg_0106;
    56: op1_14_in08 = reg_1065;
    50: op1_14_in08 = reg_0921;
    76: op1_14_in08 = reg_0134;
    71: op1_14_in08 = imem00_in[3:0];
    87: op1_14_in08 = reg_1184;
    57: op1_14_in08 = reg_1170;
    68: op1_14_in08 = reg_0125;
    77: op1_14_in08 = reg_0340;
    61: op1_14_in08 = reg_0492;
    78: op1_14_in08 = imem05_in[7:4];
    117: op1_14_in08 = imem05_in[7:4];
    58: op1_14_in08 = reg_1098;
    70: op1_14_in08 = reg_1208;
    59: op1_14_in08 = reg_0631;
    79: op1_14_in08 = reg_0161;
    51: op1_14_in08 = reg_0360;
    60: op1_14_in08 = reg_0330;
    80: op1_14_in08 = reg_0617;
    88: op1_14_in08 = reg_0629;
    62: op1_14_in08 = reg_0287;
    81: op1_14_in08 = reg_0795;
    82: op1_14_in08 = reg_0325;
    52: op1_14_in08 = reg_0457;
    63: op1_14_in08 = reg_0157;
    64: op1_14_in08 = reg_0507;
    83: op1_14_in08 = reg_1470;
    89: op1_14_in08 = reg_0034;
    84: op1_14_in08 = reg_1514;
    85: op1_14_in08 = reg_0293;
    65: op1_14_in08 = reg_0162;
    90: op1_14_in08 = reg_0375;
    66: op1_14_in08 = reg_0093;
    48: op1_14_in08 = reg_0014;
    113: op1_14_in08 = reg_0014;
    91: op1_14_in08 = reg_1027;
    46: op1_14_in08 = reg_0009;
    67: op1_14_in08 = reg_0346;
    92: op1_14_in08 = reg_1202;
    108: op1_14_in08 = reg_1202;
    93: op1_14_in08 = reg_0470;
    94: op1_14_in08 = reg_1206;
    95: op1_14_in08 = reg_0269;
    97: op1_14_in08 = reg_0311;
    98: op1_14_in08 = reg_0846;
    99: op1_14_in08 = reg_0167;
    100: op1_14_in08 = reg_0381;
    101: op1_14_in08 = reg_0171;
    102: op1_14_in08 = reg_0662;
    103: op1_14_in08 = reg_1233;
    104: op1_14_in08 = reg_0702;
    105: op1_14_in08 = reg_0583;
    106: op1_14_in08 = reg_0428;
    107: op1_14_in08 = reg_0423;
    37: op1_14_in08 = reg_0664;
    109: op1_14_in08 = reg_0427;
    110: op1_14_in08 = reg_0640;
    111: op1_14_in08 = reg_0601;
    112: op1_14_in08 = reg_1230;
    114: op1_14_in08 = reg_0970;
    115: op1_14_in08 = reg_0196;
    116: op1_14_in08 = reg_0054;
    118: op1_14_in08 = reg_0317;
    119: op1_14_in08 = reg_0408;
    47: op1_14_in08 = reg_0141;
    120: op1_14_in08 = reg_0459;
    121: op1_14_in08 = reg_0012;
    122: op1_14_in08 = reg_1227;
    123: op1_14_in08 = reg_0518;
    124: op1_14_in08 = reg_0534;
    125: op1_14_in08 = reg_0103;
    126: op1_14_in08 = reg_0598;
    127: op1_14_in08 = reg_1231;
    128: op1_14_in08 = reg_0659;
    129: op1_14_in08 = reg_0329;
    130: op1_14_in08 = reg_1455;
    default: op1_14_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_14_inv08 = 1;
    75: op1_14_inv08 = 1;
    50: op1_14_inv08 = 1;
    76: op1_14_inv08 = 1;
    71: op1_14_inv08 = 1;
    87: op1_14_inv08 = 1;
    77: op1_14_inv08 = 1;
    61: op1_14_inv08 = 1;
    78: op1_14_inv08 = 1;
    59: op1_14_inv08 = 1;
    79: op1_14_inv08 = 1;
    51: op1_14_inv08 = 1;
    60: op1_14_inv08 = 1;
    88: op1_14_inv08 = 1;
    62: op1_14_inv08 = 1;
    82: op1_14_inv08 = 1;
    64: op1_14_inv08 = 1;
    65: op1_14_inv08 = 1;
    90: op1_14_inv08 = 1;
    66: op1_14_inv08 = 1;
    48: op1_14_inv08 = 1;
    67: op1_14_inv08 = 1;
    92: op1_14_inv08 = 1;
    93: op1_14_inv08 = 1;
    99: op1_14_inv08 = 1;
    100: op1_14_inv08 = 1;
    104: op1_14_inv08 = 1;
    106: op1_14_inv08 = 1;
    37: op1_14_inv08 = 1;
    110: op1_14_inv08 = 1;
    111: op1_14_inv08 = 1;
    113: op1_14_inv08 = 1;
    114: op1_14_inv08 = 1;
    116: op1_14_inv08 = 1;
    117: op1_14_inv08 = 1;
    120: op1_14_inv08 = 1;
    121: op1_14_inv08 = 1;
    123: op1_14_inv08 = 1;
    124: op1_14_inv08 = 1;
    125: op1_14_inv08 = 1;
    126: op1_14_inv08 = 1;
    130: op1_14_inv08 = 1;
    default: op1_14_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in09 = reg_0524;
    53: op1_14_in09 = reg_0539;
    73: op1_14_in09 = reg_0155;
    55: op1_14_in09 = reg_0213;
    86: op1_14_in09 = reg_0481;
    74: op1_14_in09 = reg_0109;
    54: op1_14_in09 = reg_0646;
    75: op1_14_in09 = reg_0938;
    49: op1_14_in09 = reg_0263;
    69: op1_14_in09 = reg_0876;
    56: op1_14_in09 = reg_0421;
    50: op1_14_in09 = reg_0924;
    76: op1_14_in09 = reg_0027;
    71: op1_14_in09 = reg_0250;
    87: op1_14_in09 = reg_1314;
    57: op1_14_in09 = reg_0230;
    68: op1_14_in09 = reg_0711;
    77: op1_14_in09 = reg_0305;
    61: op1_14_in09 = reg_0883;
    78: op1_14_in09 = reg_0697;
    58: op1_14_in09 = reg_0607;
    70: op1_14_in09 = reg_0107;
    59: op1_14_in09 = reg_0578;
    79: op1_14_in09 = reg_0116;
    51: op1_14_in09 = reg_0047;
    60: op1_14_in09 = reg_1282;
    80: op1_14_in09 = reg_0526;
    88: op1_14_in09 = reg_1032;
    62: op1_14_in09 = reg_0739;
    81: op1_14_in09 = reg_1426;
    82: op1_14_in09 = reg_0889;
    52: op1_14_in09 = reg_1095;
    63: op1_14_in09 = reg_0923;
    64: op1_14_in09 = reg_0478;
    83: op1_14_in09 = reg_1052;
    89: op1_14_in09 = reg_1257;
    84: op1_14_in09 = reg_0300;
    85: op1_14_in09 = reg_0249;
    65: op1_14_in09 = reg_0821;
    90: op1_14_in09 = reg_0377;
    66: op1_14_in09 = reg_0901;
    48: op1_14_in09 = reg_0784;
    91: op1_14_in09 = reg_1229;
    46: op1_14_in09 = reg_0154;
    67: op1_14_in09 = reg_0174;
    92: op1_14_in09 = reg_0023;
    93: op1_14_in09 = imem05_in[7:4];
    94: op1_14_in09 = reg_1405;
    95: op1_14_in09 = reg_0018;
    97: op1_14_in09 = reg_1518;
    98: op1_14_in09 = reg_0456;
    99: op1_14_in09 = reg_1403;
    100: op1_14_in09 = reg_0829;
    101: op1_14_in09 = reg_0165;
    102: op1_14_in09 = reg_0989;
    103: op1_14_in09 = reg_1082;
    104: op1_14_in09 = reg_0184;
    105: op1_14_in09 = reg_0371;
    106: op1_14_in09 = reg_0388;
    107: op1_14_in09 = reg_1493;
    37: op1_14_in09 = reg_0366;
    108: op1_14_in09 = reg_0215;
    109: op1_14_in09 = reg_0577;
    110: op1_14_in09 = reg_1053;
    111: op1_14_in09 = reg_0393;
    115: op1_14_in09 = reg_0393;
    112: op1_14_in09 = reg_0459;
    113: op1_14_in09 = reg_1035;
    114: op1_14_in09 = reg_0972;
    116: op1_14_in09 = reg_0326;
    117: op1_14_in09 = imem05_in[11:8];
    118: op1_14_in09 = imem06_in[3:0];
    119: op1_14_in09 = reg_0415;
    47: op1_14_in09 = reg_0720;
    120: op1_14_in09 = reg_0887;
    121: op1_14_in09 = reg_0011;
    122: op1_14_in09 = reg_1205;
    123: op1_14_in09 = reg_0124;
    124: op1_14_in09 = reg_0181;
    125: op1_14_in09 = reg_0321;
    126: op1_14_in09 = reg_0454;
    127: op1_14_in09 = reg_1226;
    128: op1_14_in09 = reg_0606;
    129: op1_14_in09 = reg_1093;
    130: op1_14_in09 = reg_0127;
    default: op1_14_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    75: op1_14_inv09 = 1;
    69: op1_14_inv09 = 1;
    50: op1_14_inv09 = 1;
    76: op1_14_inv09 = 1;
    58: op1_14_inv09 = 1;
    79: op1_14_inv09 = 1;
    80: op1_14_inv09 = 1;
    88: op1_14_inv09 = 1;
    82: op1_14_inv09 = 1;
    89: op1_14_inv09 = 1;
    84: op1_14_inv09 = 1;
    85: op1_14_inv09 = 1;
    65: op1_14_inv09 = 1;
    66: op1_14_inv09 = 1;
    48: op1_14_inv09 = 1;
    91: op1_14_inv09 = 1;
    95: op1_14_inv09 = 1;
    97: op1_14_inv09 = 1;
    98: op1_14_inv09 = 1;
    102: op1_14_inv09 = 1;
    103: op1_14_inv09 = 1;
    104: op1_14_inv09 = 1;
    105: op1_14_inv09 = 1;
    108: op1_14_inv09 = 1;
    113: op1_14_inv09 = 1;
    116: op1_14_inv09 = 1;
    118: op1_14_inv09 = 1;
    119: op1_14_inv09 = 1;
    47: op1_14_inv09 = 1;
    120: op1_14_inv09 = 1;
    122: op1_14_inv09 = 1;
    123: op1_14_inv09 = 1;
    125: op1_14_inv09 = 1;
    128: op1_14_inv09 = 1;
    default: op1_14_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in10 = reg_1405;
    53: op1_14_in10 = reg_0937;
    73: op1_14_in10 = reg_1418;
    55: op1_14_in10 = reg_0230;
    86: op1_14_in10 = imem03_in[3:0];
    74: op1_14_in10 = reg_0717;
    54: op1_14_in10 = reg_0648;
    75: op1_14_in10 = reg_0302;
    49: op1_14_in10 = reg_0264;
    69: op1_14_in10 = reg_0009;
    56: op1_14_in10 = reg_0414;
    50: op1_14_in10 = reg_0489;
    76: op1_14_in10 = reg_1100;
    71: op1_14_in10 = reg_0293;
    87: op1_14_in10 = reg_0957;
    57: op1_14_in10 = reg_0490;
    68: op1_14_in10 = reg_0153;
    77: op1_14_in10 = reg_0487;
    61: op1_14_in10 = reg_0886;
    78: op1_14_in10 = reg_1402;
    58: op1_14_in10 = reg_1018;
    70: op1_14_in10 = reg_0113;
    59: op1_14_in10 = reg_0750;
    79: op1_14_in10 = reg_0110;
    51: op1_14_in10 = reg_0078;
    60: op1_14_in10 = reg_0790;
    80: op1_14_in10 = reg_0529;
    88: op1_14_in10 = reg_1098;
    62: op1_14_in10 = reg_0404;
    81: op1_14_in10 = reg_1209;
    82: op1_14_in10 = reg_0235;
    52: op1_14_in10 = reg_0995;
    63: op1_14_in10 = reg_0139;
    64: op1_14_in10 = reg_0348;
    83: op1_14_in10 = reg_0250;
    89: op1_14_in10 = reg_1203;
    84: op1_14_in10 = reg_1373;
    85: op1_14_in10 = reg_1206;
    91: op1_14_in10 = reg_1206;
    65: op1_14_in10 = reg_1056;
    90: op1_14_in10 = reg_1003;
    66: op1_14_in10 = imem01_in[15:12];
    48: op1_14_in10 = reg_0752;
    46: op1_14_in10 = reg_0829;
    67: op1_14_in10 = reg_0650;
    92: op1_14_in10 = reg_0046;
    93: op1_14_in10 = reg_1299;
    94: op1_14_in10 = reg_0927;
    110: op1_14_in10 = reg_0927;
    95: op1_14_in10 = reg_0993;
    97: op1_14_in10 = reg_0048;
    98: op1_14_in10 = reg_0608;
    99: op1_14_in10 = reg_0183;
    100: op1_14_in10 = reg_0897;
    101: op1_14_in10 = reg_1170;
    102: op1_14_in10 = reg_0530;
    103: op1_14_in10 = reg_0537;
    104: op1_14_in10 = reg_0700;
    105: op1_14_in10 = reg_0195;
    106: op1_14_in10 = reg_0075;
    107: op1_14_in10 = reg_0390;
    37: op1_14_in10 = imem07_in[11:8];
    108: op1_14_in10 = reg_0017;
    109: op1_14_in10 = reg_0263;
    111: op1_14_in10 = reg_0130;
    112: op1_14_in10 = reg_0524;
    113: op1_14_in10 = reg_0905;
    114: op1_14_in10 = reg_0128;
    115: op1_14_in10 = reg_0243;
    116: op1_14_in10 = reg_0970;
    117: op1_14_in10 = reg_0735;
    118: op1_14_in10 = reg_0825;
    119: op1_14_in10 = reg_0413;
    47: op1_14_in10 = reg_0671;
    120: op1_14_in10 = reg_0883;
    121: op1_14_in10 = reg_0166;
    122: op1_14_in10 = reg_1406;
    123: op1_14_in10 = reg_0246;
    124: op1_14_in10 = reg_1368;
    125: op1_14_in10 = reg_1351;
    126: op1_14_in10 = reg_1004;
    127: op1_14_in10 = reg_0178;
    128: op1_14_in10 = reg_0845;
    129: op1_14_in10 = reg_1092;
    130: op1_14_in10 = reg_0106;
    default: op1_14_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv10 = 1;
    73: op1_14_inv10 = 1;
    86: op1_14_inv10 = 1;
    74: op1_14_inv10 = 1;
    75: op1_14_inv10 = 1;
    49: op1_14_inv10 = 1;
    69: op1_14_inv10 = 1;
    56: op1_14_inv10 = 1;
    71: op1_14_inv10 = 1;
    87: op1_14_inv10 = 1;
    57: op1_14_inv10 = 1;
    68: op1_14_inv10 = 1;
    77: op1_14_inv10 = 1;
    61: op1_14_inv10 = 1;
    78: op1_14_inv10 = 1;
    58: op1_14_inv10 = 1;
    70: op1_14_inv10 = 1;
    51: op1_14_inv10 = 1;
    60: op1_14_inv10 = 1;
    80: op1_14_inv10 = 1;
    88: op1_14_inv10 = 1;
    62: op1_14_inv10 = 1;
    52: op1_14_inv10 = 1;
    63: op1_14_inv10 = 1;
    89: op1_14_inv10 = 1;
    84: op1_14_inv10 = 1;
    65: op1_14_inv10 = 1;
    90: op1_14_inv10 = 1;
    66: op1_14_inv10 = 1;
    48: op1_14_inv10 = 1;
    91: op1_14_inv10 = 1;
    93: op1_14_inv10 = 1;
    94: op1_14_inv10 = 1;
    95: op1_14_inv10 = 1;
    97: op1_14_inv10 = 1;
    98: op1_14_inv10 = 1;
    99: op1_14_inv10 = 1;
    101: op1_14_inv10 = 1;
    102: op1_14_inv10 = 1;
    105: op1_14_inv10 = 1;
    110: op1_14_inv10 = 1;
    116: op1_14_inv10 = 1;
    118: op1_14_inv10 = 1;
    119: op1_14_inv10 = 1;
    120: op1_14_inv10 = 1;
    121: op1_14_inv10 = 1;
    122: op1_14_inv10 = 1;
    123: op1_14_inv10 = 1;
    127: op1_14_inv10 = 1;
    128: op1_14_inv10 = 1;
    130: op1_14_inv10 = 1;
    default: op1_14_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in11 = reg_1393;
    110: op1_14_in11 = reg_1393;
    112: op1_14_in11 = reg_1393;
    53: op1_14_in11 = reg_0938;
    73: op1_14_in11 = reg_1406;
    55: op1_14_in11 = reg_0191;
    86: op1_14_in11 = imem03_in[11:8];
    74: op1_14_in11 = reg_0637;
    54: op1_14_in11 = reg_0567;
    75: op1_14_in11 = reg_1486;
    49: op1_14_in11 = reg_0619;
    69: op1_14_in11 = reg_0848;
    56: op1_14_in11 = reg_0407;
    50: op1_14_in11 = reg_0465;
    76: op1_14_in11 = reg_1256;
    71: op1_14_in11 = reg_1229;
    87: op1_14_in11 = reg_0952;
    57: op1_14_in11 = reg_0821;
    68: op1_14_in11 = reg_0294;
    77: op1_14_in11 = reg_0862;
    61: op1_14_in11 = reg_0638;
    78: op1_14_in11 = reg_1070;
    58: op1_14_in11 = reg_0588;
    70: op1_14_in11 = reg_0104;
    59: op1_14_in11 = reg_0733;
    79: op1_14_in11 = reg_1302;
    51: op1_14_in11 = reg_0290;
    60: op1_14_in11 = reg_0425;
    80: op1_14_in11 = reg_0295;
    88: op1_14_in11 = reg_0800;
    62: op1_14_in11 = reg_0621;
    81: op1_14_in11 = reg_0160;
    82: op1_14_in11 = imem03_in[3:0];
    52: op1_14_in11 = reg_0704;
    63: op1_14_in11 = reg_0224;
    64: op1_14_in11 = reg_0247;
    83: op1_14_in11 = reg_0293;
    89: op1_14_in11 = reg_1214;
    84: op1_14_in11 = reg_0037;
    85: op1_14_in11 = reg_1417;
    65: op1_14_in11 = reg_0994;
    90: op1_14_in11 = reg_1184;
    66: op1_14_in11 = reg_0078;
    48: op1_14_in11 = reg_0751;
    91: op1_14_in11 = reg_0524;
    46: op1_14_in11 = reg_0024;
    67: op1_14_in11 = reg_0333;
    92: op1_14_in11 = reg_0212;
    93: op1_14_in11 = reg_0832;
    94: op1_14_in11 = reg_0027;
    95: op1_14_in11 = reg_0995;
    97: op1_14_in11 = reg_0025;
    98: op1_14_in11 = reg_0055;
    99: op1_14_in11 = reg_0477;
    100: op1_14_in11 = reg_1515;
    101: op1_14_in11 = imem07_in[11:8];
    102: op1_14_in11 = reg_0879;
    103: op1_14_in11 = reg_1004;
    104: op1_14_in11 = reg_1104;
    105: op1_14_in11 = reg_0977;
    106: op1_14_in11 = reg_0060;
    107: op1_14_in11 = reg_1458;
    37: op1_14_in11 = reg_0404;
    108: op1_14_in11 = reg_0963;
    109: op1_14_in11 = reg_1372;
    111: op1_14_in11 = reg_1348;
    113: op1_14_in11 = reg_0730;
    114: op1_14_in11 = reg_0629;
    130: op1_14_in11 = reg_0629;
    115: op1_14_in11 = reg_0240;
    116: op1_14_in11 = reg_1451;
    117: op1_14_in11 = reg_0466;
    118: op1_14_in11 = reg_0372;
    119: op1_14_in11 = reg_0623;
    47: op1_14_in11 = reg_0634;
    120: op1_14_in11 = reg_0201;
    121: op1_14_in11 = reg_0447;
    122: op1_14_in11 = reg_0476;
    123: op1_14_in11 = reg_0791;
    124: op1_14_in11 = reg_1367;
    125: op1_14_in11 = reg_0998;
    126: op1_14_in11 = reg_0451;
    127: op1_14_in11 = reg_0108;
    128: op1_14_in11 = reg_0846;
    129: op1_14_in11 = reg_0178;
    default: op1_14_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_14_inv11 = 1;
    55: op1_14_inv11 = 1;
    86: op1_14_inv11 = 1;
    74: op1_14_inv11 = 1;
    54: op1_14_inv11 = 1;
    49: op1_14_inv11 = 1;
    69: op1_14_inv11 = 1;
    77: op1_14_inv11 = 1;
    61: op1_14_inv11 = 1;
    78: op1_14_inv11 = 1;
    58: op1_14_inv11 = 1;
    59: op1_14_inv11 = 1;
    79: op1_14_inv11 = 1;
    51: op1_14_inv11 = 1;
    88: op1_14_inv11 = 1;
    62: op1_14_inv11 = 1;
    81: op1_14_inv11 = 1;
    82: op1_14_inv11 = 1;
    63: op1_14_inv11 = 1;
    65: op1_14_inv11 = 1;
    91: op1_14_inv11 = 1;
    97: op1_14_inv11 = 1;
    99: op1_14_inv11 = 1;
    100: op1_14_inv11 = 1;
    106: op1_14_inv11 = 1;
    37: op1_14_inv11 = 1;
    108: op1_14_inv11 = 1;
    110: op1_14_inv11 = 1;
    111: op1_14_inv11 = 1;
    113: op1_14_inv11 = 1;
    114: op1_14_inv11 = 1;
    117: op1_14_inv11 = 1;
    47: op1_14_inv11 = 1;
    123: op1_14_inv11 = 1;
    126: op1_14_inv11 = 1;
    default: op1_14_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in12 = reg_0887;
    53: op1_14_in12 = reg_0163;
    73: op1_14_in12 = reg_1393;
    55: op1_14_in12 = reg_0162;
    86: op1_14_in12 = reg_1282;
    74: op1_14_in12 = reg_0529;
    54: op1_14_in12 = reg_0066;
    75: op1_14_in12 = reg_0576;
    49: op1_14_in12 = reg_0617;
    69: op1_14_in12 = reg_0802;
    56: op1_14_in12 = reg_0452;
    126: op1_14_in12 = reg_0452;
    50: op1_14_in12 = reg_0030;
    76: op1_14_in12 = imem01_in[7:4];
    71: op1_14_in12 = reg_1205;
    87: op1_14_in12 = reg_0190;
    57: op1_14_in12 = imem07_in[11:8];
    68: op1_14_in12 = reg_0531;
    77: op1_14_in12 = reg_0097;
    61: op1_14_in12 = reg_0409;
    78: op1_14_in12 = reg_0939;
    58: op1_14_in12 = reg_0590;
    70: op1_14_in12 = reg_0479;
    59: op1_14_in12 = reg_0833;
    79: op1_14_in12 = reg_0636;
    51: op1_14_in12 = reg_0043;
    60: op1_14_in12 = reg_0247;
    80: op1_14_in12 = reg_0022;
    88: op1_14_in12 = imem03_in[7:4];
    62: op1_14_in12 = reg_0593;
    81: op1_14_in12 = reg_1505;
    82: op1_14_in12 = reg_1448;
    52: op1_14_in12 = reg_0310;
    63: op1_14_in12 = reg_0665;
    64: op1_14_in12 = reg_1082;
    89: op1_14_in12 = reg_1082;
    83: op1_14_in12 = reg_1028;
    84: op1_14_in12 = reg_1064;
    85: op1_14_in12 = reg_0155;
    65: op1_14_in12 = reg_0993;
    90: op1_14_in12 = reg_0964;
    66: op1_14_in12 = reg_0290;
    48: op1_14_in12 = reg_0194;
    91: op1_14_in12 = reg_0928;
    46: op1_14_in12 = reg_0069;
    67: op1_14_in12 = reg_0182;
    92: op1_14_in12 = reg_0213;
    93: op1_14_in12 = reg_0702;
    94: op1_14_in12 = reg_0871;
    95: op1_14_in12 = reg_1414;
    97: op1_14_in12 = reg_1369;
    98: op1_14_in12 = reg_1343;
    99: op1_14_in12 = reg_0418;
    100: op1_14_in12 = reg_0154;
    101: op1_14_in12 = reg_0226;
    102: op1_14_in12 = reg_0497;
    103: op1_14_in12 = reg_0320;
    104: op1_14_in12 = reg_1404;
    105: op1_14_in12 = reg_0067;
    106: op1_14_in12 = reg_0058;
    107: op1_14_in12 = reg_0111;
    37: op1_14_in12 = reg_0415;
    108: op1_14_in12 = reg_1183;
    109: op1_14_in12 = reg_0088;
    124: op1_14_in12 = reg_0088;
    110: op1_14_in12 = reg_0405;
    111: op1_14_in12 = reg_0603;
    112: op1_14_in12 = reg_0387;
    113: op1_14_in12 = reg_1326;
    114: op1_14_in12 = reg_0496;
    130: op1_14_in12 = reg_0496;
    115: op1_14_in12 = reg_0575;
    116: op1_14_in12 = reg_0382;
    117: op1_14_in12 = reg_0278;
    118: op1_14_in12 = reg_0669;
    119: op1_14_in12 = reg_0591;
    47: op1_14_in12 = reg_0635;
    120: op1_14_in12 = reg_0428;
    121: op1_14_in12 = reg_0877;
    122: op1_14_in12 = reg_0188;
    123: op1_14_in12 = reg_1055;
    125: op1_14_in12 = reg_0002;
    127: op1_14_in12 = reg_0104;
    128: op1_14_in12 = reg_0056;
    129: op1_14_in12 = reg_1208;
    default: op1_14_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_14_inv12 = 1;
    55: op1_14_inv12 = 1;
    86: op1_14_inv12 = 1;
    74: op1_14_inv12 = 1;
    54: op1_14_inv12 = 1;
    49: op1_14_inv12 = 1;
    69: op1_14_inv12 = 1;
    50: op1_14_inv12 = 1;
    57: op1_14_inv12 = 1;
    68: op1_14_inv12 = 1;
    61: op1_14_inv12 = 1;
    78: op1_14_inv12 = 1;
    58: op1_14_inv12 = 1;
    70: op1_14_inv12 = 1;
    62: op1_14_inv12 = 1;
    82: op1_14_inv12 = 1;
    63: op1_14_inv12 = 1;
    83: op1_14_inv12 = 1;
    84: op1_14_inv12 = 1;
    85: op1_14_inv12 = 1;
    65: op1_14_inv12 = 1;
    92: op1_14_inv12 = 1;
    94: op1_14_inv12 = 1;
    103: op1_14_inv12 = 1;
    106: op1_14_inv12 = 1;
    107: op1_14_inv12 = 1;
    109: op1_14_inv12 = 1;
    114: op1_14_inv12 = 1;
    115: op1_14_inv12 = 1;
    118: op1_14_inv12 = 1;
    122: op1_14_inv12 = 1;
    125: op1_14_inv12 = 1;
    127: op1_14_inv12 = 1;
    129: op1_14_inv12 = 1;
    default: op1_14_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in13 = reg_0202;
    53: op1_14_in13 = reg_0896;
    73: op1_14_in13 = reg_0881;
    55: op1_14_in13 = reg_1096;
    86: op1_14_in13 = reg_0425;
    74: op1_14_in13 = reg_0345;
    54: op1_14_in13 = reg_0538;
    75: op1_14_in13 = reg_0197;
    49: op1_14_in13 = reg_0528;
    69: op1_14_in13 = reg_0311;
    56: op1_14_in13 = reg_0305;
    50: op1_14_in13 = reg_0286;
    76: op1_14_in13 = reg_0743;
    71: op1_14_in13 = reg_0460;
    87: op1_14_in13 = reg_0246;
    57: op1_14_in13 = reg_0461;
    68: op1_14_in13 = reg_0839;
    77: op1_14_in13 = reg_0117;
    61: op1_14_in13 = reg_0351;
    91: op1_14_in13 = reg_0351;
    78: op1_14_in13 = reg_0938;
    58: op1_14_in13 = reg_0587;
    70: op1_14_in13 = reg_0525;
    59: op1_14_in13 = reg_0168;
    79: op1_14_in13 = reg_0373;
    51: op1_14_in13 = reg_0042;
    60: op1_14_in13 = reg_0698;
    80: op1_14_in13 = reg_0017;
    92: op1_14_in13 = reg_0017;
    88: op1_14_in13 = reg_1063;
    82: op1_14_in13 = reg_1063;
    62: op1_14_in13 = reg_0051;
    81: op1_14_in13 = reg_0172;
    52: op1_14_in13 = reg_0297;
    63: op1_14_in13 = reg_0591;
    64: op1_14_in13 = reg_0552;
    83: op1_14_in13 = reg_1418;
    85: op1_14_in13 = reg_1418;
    89: op1_14_in13 = reg_0342;
    126: op1_14_in13 = reg_0342;
    84: op1_14_in13 = reg_1426;
    65: op1_14_in13 = reg_0998;
    90: op1_14_in13 = reg_1518;
    66: op1_14_in13 = reg_0012;
    48: op1_14_in13 = reg_0195;
    46: op1_14_in13 = reg_0325;
    67: op1_14_in13 = imem05_in[3:0];
    93: op1_14_in13 = reg_1268;
    94: op1_14_in13 = reg_1152;
    95: op1_14_in13 = reg_1416;
    97: op1_14_in13 = reg_0462;
    98: op1_14_in13 = reg_0822;
    99: op1_14_in13 = reg_0301;
    100: op1_14_in13 = reg_0049;
    101: op1_14_in13 = reg_0324;
    102: op1_14_in13 = reg_1002;
    103: op1_14_in13 = reg_0368;
    104: op1_14_in13 = reg_0940;
    105: op1_14_in13 = reg_0023;
    106: op1_14_in13 = reg_1322;
    107: op1_14_in13 = reg_0382;
    37: op1_14_in13 = reg_0137;
    108: op1_14_in13 = reg_1415;
    109: op1_14_in13 = reg_0694;
    110: op1_14_in13 = reg_0026;
    111: op1_14_in13 = reg_0038;
    112: op1_14_in13 = reg_0075;
    113: op1_14_in13 = reg_0720;
    114: op1_14_in13 = reg_1140;
    115: op1_14_in13 = reg_0207;
    116: op1_14_in13 = reg_0629;
    117: op1_14_in13 = reg_0272;
    118: op1_14_in13 = reg_0397;
    119: op1_14_in13 = reg_0592;
    47: op1_14_in13 = reg_0624;
    120: op1_14_in13 = reg_0005;
    121: op1_14_in13 = reg_0399;
    122: op1_14_in13 = reg_0722;
    123: op1_14_in13 = reg_0219;
    124: op1_14_in13 = reg_0319;
    125: op1_14_in13 = reg_0053;
    127: op1_14_in13 = reg_0884;
    129: op1_14_in13 = reg_0884;
    128: op1_14_in13 = reg_0608;
    130: op1_14_in13 = reg_0473;
    default: op1_14_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_14_inv13 = 1;
    86: op1_14_inv13 = 1;
    74: op1_14_inv13 = 1;
    54: op1_14_inv13 = 1;
    69: op1_14_inv13 = 1;
    56: op1_14_inv13 = 1;
    50: op1_14_inv13 = 1;
    68: op1_14_inv13 = 1;
    77: op1_14_inv13 = 1;
    61: op1_14_inv13 = 1;
    79: op1_14_inv13 = 1;
    80: op1_14_inv13 = 1;
    88: op1_14_inv13 = 1;
    62: op1_14_inv13 = 1;
    81: op1_14_inv13 = 1;
    82: op1_14_inv13 = 1;
    83: op1_14_inv13 = 1;
    85: op1_14_inv13 = 1;
    65: op1_14_inv13 = 1;
    90: op1_14_inv13 = 1;
    48: op1_14_inv13 = 1;
    91: op1_14_inv13 = 1;
    46: op1_14_inv13 = 1;
    67: op1_14_inv13 = 1;
    92: op1_14_inv13 = 1;
    95: op1_14_inv13 = 1;
    97: op1_14_inv13 = 1;
    98: op1_14_inv13 = 1;
    101: op1_14_inv13 = 1;
    103: op1_14_inv13 = 1;
    105: op1_14_inv13 = 1;
    106: op1_14_inv13 = 1;
    107: op1_14_inv13 = 1;
    37: op1_14_inv13 = 1;
    109: op1_14_inv13 = 1;
    110: op1_14_inv13 = 1;
    111: op1_14_inv13 = 1;
    114: op1_14_inv13 = 1;
    119: op1_14_inv13 = 1;
    47: op1_14_inv13 = 1;
    120: op1_14_inv13 = 1;
    121: op1_14_inv13 = 1;
    122: op1_14_inv13 = 1;
    126: op1_14_inv13 = 1;
    127: op1_14_inv13 = 1;
    128: op1_14_inv13 = 1;
    default: op1_14_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in14 = reg_0353;
    53: op1_14_in14 = reg_0130;
    73: op1_14_in14 = reg_0201;
    122: op1_14_in14 = reg_0201;
    55: op1_14_in14 = imem07_in[15:12];
    86: op1_14_in14 = reg_0443;
    74: op1_14_in14 = reg_1225;
    54: op1_14_in14 = reg_0940;
    75: op1_14_in14 = reg_0243;
    49: op1_14_in14 = reg_0132;
    69: op1_14_in14 = reg_0756;
    56: op1_14_in14 = reg_0319;
    50: op1_14_in14 = reg_0441;
    76: op1_14_in14 = reg_1473;
    71: op1_14_in14 = reg_1417;
    87: op1_14_in14 = reg_1092;
    57: op1_14_in14 = reg_0629;
    65: op1_14_in14 = reg_0629;
    68: op1_14_in14 = reg_0069;
    77: op1_14_in14 = reg_0020;
    61: op1_14_in14 = reg_0352;
    78: op1_14_in14 = reg_0183;
    58: op1_14_in14 = reg_0561;
    70: op1_14_in14 = reg_0734;
    59: op1_14_in14 = reg_1164;
    79: op1_14_in14 = reg_0586;
    47: op1_14_in14 = reg_0586;
    51: op1_14_in14 = reg_0553;
    60: op1_14_in14 = reg_1144;
    80: op1_14_in14 = reg_0391;
    88: op1_14_in14 = reg_0378;
    62: op1_14_in14 = reg_0003;
    63: op1_14_in14 = reg_0003;
    81: op1_14_in14 = reg_0115;
    82: op1_14_in14 = reg_1425;
    52: op1_14_in14 = reg_0673;
    64: op1_14_in14 = reg_0407;
    83: op1_14_in14 = reg_0883;
    85: op1_14_in14 = reg_0883;
    89: op1_14_in14 = reg_0340;
    84: op1_14_in14 = reg_0264;
    90: op1_14_in14 = reg_1093;
    66: op1_14_in14 = reg_0662;
    48: op1_14_in14 = imem06_in[3:0];
    91: op1_14_in14 = reg_0428;
    46: op1_14_in14 = reg_0279;
    67: op1_14_in14 = reg_0540;
    92: op1_14_in14 = imem07_in[3:0];
    95: op1_14_in14 = imem07_in[3:0];
    93: op1_14_in14 = reg_0996;
    94: op1_14_in14 = reg_0282;
    97: op1_14_in14 = reg_0297;
    98: op1_14_in14 = reg_1260;
    99: op1_14_in14 = reg_0318;
    100: op1_14_in14 = reg_1494;
    101: op1_14_in14 = reg_0394;
    102: op1_14_in14 = reg_0256;
    103: op1_14_in14 = reg_0862;
    104: op1_14_in14 = reg_0939;
    105: op1_14_in14 = reg_0215;
    106: op1_14_in14 = reg_1032;
    107: op1_14_in14 = reg_0496;
    116: op1_14_in14 = reg_0496;
    37: op1_14_in14 = reg_0228;
    108: op1_14_in14 = reg_0298;
    109: op1_14_in14 = reg_0471;
    110: op1_14_in14 = reg_0027;
    111: op1_14_in14 = reg_0014;
    112: op1_14_in14 = reg_0059;
    113: op1_14_in14 = reg_1179;
    114: op1_14_in14 = reg_0628;
    115: op1_14_in14 = imem05_in[11:8];
    117: op1_14_in14 = reg_1268;
    118: op1_14_in14 = reg_0782;
    119: op1_14_in14 = reg_0321;
    120: op1_14_in14 = reg_1090;
    121: op1_14_in14 = reg_0276;
    123: op1_14_in14 = reg_0703;
    124: op1_14_in14 = reg_0552;
    125: op1_14_in14 = reg_1182;
    126: op1_14_in14 = reg_0097;
    127: op1_14_in14 = reg_0458;
    128: op1_14_in14 = reg_0588;
    129: op1_14_in14 = reg_0448;
    130: op1_14_in14 = reg_0829;
    default: op1_14_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_14_inv14 = 1;
    55: op1_14_inv14 = 1;
    54: op1_14_inv14 = 1;
    69: op1_14_inv14 = 1;
    76: op1_14_inv14 = 1;
    71: op1_14_inv14 = 1;
    57: op1_14_inv14 = 1;
    68: op1_14_inv14 = 1;
    77: op1_14_inv14 = 1;
    61: op1_14_inv14 = 1;
    58: op1_14_inv14 = 1;
    59: op1_14_inv14 = 1;
    79: op1_14_inv14 = 1;
    51: op1_14_inv14 = 1;
    80: op1_14_inv14 = 1;
    88: op1_14_inv14 = 1;
    62: op1_14_inv14 = 1;
    89: op1_14_inv14 = 1;
    84: op1_14_inv14 = 1;
    65: op1_14_inv14 = 1;
    90: op1_14_inv14 = 1;
    66: op1_14_inv14 = 1;
    67: op1_14_inv14 = 1;
    94: op1_14_inv14 = 1;
    102: op1_14_inv14 = 1;
    104: op1_14_inv14 = 1;
    37: op1_14_inv14 = 1;
    108: op1_14_inv14 = 1;
    109: op1_14_inv14 = 1;
    111: op1_14_inv14 = 1;
    113: op1_14_inv14 = 1;
    114: op1_14_inv14 = 1;
    115: op1_14_inv14 = 1;
    116: op1_14_inv14 = 1;
    117: op1_14_inv14 = 1;
    121: op1_14_inv14 = 1;
    122: op1_14_inv14 = 1;
    123: op1_14_inv14 = 1;
    124: op1_14_inv14 = 1;
    126: op1_14_inv14 = 1;
    128: op1_14_inv14 = 1;
    default: op1_14_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in15 = reg_0352;
    53: op1_14_in15 = reg_0240;
    73: op1_14_in15 = reg_0440;
    55: op1_14_in15 = reg_0225;
    95: op1_14_in15 = reg_0225;
    86: op1_14_in15 = reg_1383;
    74: op1_14_in15 = reg_0323;
    54: op1_14_in15 = reg_0938;
    104: op1_14_in15 = reg_0938;
    75: op1_14_in15 = reg_0799;
    49: op1_14_in15 = reg_0244;
    69: op1_14_in15 = reg_0706;
    56: op1_14_in15 = reg_0487;
    50: op1_14_in15 = reg_0740;
    76: op1_14_in15 = reg_0572;
    71: op1_14_in15 = reg_0524;
    87: op1_14_in15 = reg_1208;
    57: op1_14_in15 = reg_0224;
    68: op1_14_in15 = reg_0802;
    77: op1_14_in15 = reg_0370;
    61: op1_14_in15 = reg_0075;
    78: op1_14_in15 = reg_0477;
    58: op1_14_in15 = imem02_in[3:0];
    51: op1_14_in15 = imem02_in[3:0];
    70: op1_14_in15 = reg_0573;
    59: op1_14_in15 = reg_1169;
    79: op1_14_in15 = reg_0622;
    60: op1_14_in15 = reg_1143;
    80: op1_14_in15 = reg_1440;
    88: op1_14_in15 = reg_0962;
    62: op1_14_in15 = reg_0521;
    81: op1_14_in15 = reg_0110;
    82: op1_14_in15 = reg_1033;
    52: op1_14_in15 = reg_0674;
    63: op1_14_in15 = reg_0053;
    64: op1_14_in15 = reg_0598;
    83: op1_14_in15 = reg_0428;
    122: op1_14_in15 = reg_0428;
    89: op1_14_in15 = reg_0338;
    84: op1_14_in15 = reg_1508;
    85: op1_14_in15 = reg_0886;
    65: op1_14_in15 = reg_0673;
    90: op1_14_in15 = reg_0885;
    66: op1_14_in15 = reg_0606;
    48: op1_14_in15 = reg_0908;
    91: op1_14_in15 = reg_0416;
    46: op1_14_in15 = reg_0311;
    67: op1_14_in15 = reg_0541;
    92: op1_14_in15 = reg_0498;
    93: op1_14_in15 = reg_0391;
    94: op1_14_in15 = reg_0355;
    97: op1_14_in15 = reg_1198;
    98: op1_14_in15 = reg_0971;
    99: op1_14_in15 = reg_1485;
    100: op1_14_in15 = reg_0558;
    101: op1_14_in15 = reg_1010;
    102: op1_14_in15 = reg_0382;
    103: op1_14_in15 = reg_0835;
    105: op1_14_in15 = reg_0213;
    106: op1_14_in15 = reg_1152;
    107: op1_14_in15 = reg_0381;
    37: op1_14_in15 = reg_0003;
    108: op1_14_in15 = reg_0310;
    109: op1_14_in15 = reg_1040;
    110: op1_14_in15 = reg_0723;
    111: op1_14_in15 = reg_0670;
    112: op1_14_in15 = reg_0089;
    113: op1_14_in15 = reg_0345;
    114: op1_14_in15 = reg_0876;
    115: op1_14_in15 = reg_0270;
    116: op1_14_in15 = reg_0684;
    117: op1_14_in15 = reg_0604;
    118: op1_14_in15 = reg_0984;
    119: op1_14_in15 = reg_0028;
    47: op1_14_in15 = reg_0568;
    120: op1_14_in15 = reg_0871;
    121: op1_14_in15 = reg_0822;
    123: op1_14_in15 = reg_0140;
    124: op1_14_in15 = reg_1203;
    126: op1_14_in15 = reg_0061;
    127: op1_14_in15 = reg_0831;
    128: op1_14_in15 = reg_0975;
    129: op1_14_in15 = reg_0458;
    130: op1_14_in15 = reg_0897;
    default: op1_14_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv15 = 1;
    55: op1_14_inv15 = 1;
    86: op1_14_inv15 = 1;
    54: op1_14_inv15 = 1;
    75: op1_14_inv15 = 1;
    69: op1_14_inv15 = 1;
    76: op1_14_inv15 = 1;
    87: op1_14_inv15 = 1;
    68: op1_14_inv15 = 1;
    78: op1_14_inv15 = 1;
    58: op1_14_inv15 = 1;
    59: op1_14_inv15 = 1;
    62: op1_14_inv15 = 1;
    82: op1_14_inv15 = 1;
    63: op1_14_inv15 = 1;
    83: op1_14_inv15 = 1;
    84: op1_14_inv15 = 1;
    85: op1_14_inv15 = 1;
    65: op1_14_inv15 = 1;
    90: op1_14_inv15 = 1;
    66: op1_14_inv15 = 1;
    48: op1_14_inv15 = 1;
    46: op1_14_inv15 = 1;
    67: op1_14_inv15 = 1;
    93: op1_14_inv15 = 1;
    94: op1_14_inv15 = 1;
    97: op1_14_inv15 = 1;
    99: op1_14_inv15 = 1;
    100: op1_14_inv15 = 1;
    102: op1_14_inv15 = 1;
    37: op1_14_inv15 = 1;
    111: op1_14_inv15 = 1;
    112: op1_14_inv15 = 1;
    118: op1_14_inv15 = 1;
    119: op1_14_inv15 = 1;
    122: op1_14_inv15 = 1;
    124: op1_14_inv15 = 1;
    126: op1_14_inv15 = 1;
    127: op1_14_inv15 = 1;
    129: op1_14_inv15 = 1;
    130: op1_14_inv15 = 1;
    default: op1_14_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in16 = reg_0188;
    53: op1_14_in16 = reg_0449;
    73: op1_14_in16 = reg_0071;
    122: op1_14_in16 = reg_0071;
    55: op1_14_in16 = reg_0224;
    86: op1_14_in16 = reg_0208;
    74: op1_14_in16 = reg_0583;
    54: op1_14_in16 = reg_0896;
    75: op1_14_in16 = reg_0040;
    49: op1_14_in16 = reg_0191;
    69: op1_14_in16 = reg_0704;
    56: op1_14_in16 = reg_0094;
    50: op1_14_in16 = reg_0623;
    76: op1_14_in16 = reg_0966;
    71: op1_14_in16 = reg_0189;
    87: op1_14_in16 = reg_0107;
    57: op1_14_in16 = reg_0245;
    68: op1_14_in16 = reg_0313;
    77: op1_14_in16 = reg_0273;
    61: op1_14_in16 = imem01_in[15:12];
    78: op1_14_in16 = reg_0090;
    58: op1_14_in16 = reg_0822;
    70: op1_14_in16 = reg_0443;
    59: op1_14_in16 = reg_0992;
    79: op1_14_in16 = reg_1204;
    51: op1_14_in16 = imem02_in[11:8];
    60: op1_14_in16 = imem04_in[3:0];
    80: op1_14_in16 = reg_0491;
    88: op1_14_in16 = reg_0145;
    62: op1_14_in16 = reg_1182;
    81: op1_14_in16 = reg_0714;
    82: op1_14_in16 = reg_0144;
    52: op1_14_in16 = reg_0159;
    63: op1_14_in16 = reg_0086;
    64: op1_14_in16 = reg_0369;
    83: op1_14_in16 = reg_0203;
    89: op1_14_in16 = reg_0096;
    84: op1_14_in16 = reg_0397;
    85: op1_14_in16 = reg_0722;
    65: op1_14_in16 = reg_0299;
    90: op1_14_in16 = reg_0884;
    66: op1_14_in16 = reg_0474;
    48: op1_14_in16 = reg_0905;
    91: op1_14_in16 = reg_0405;
    46: op1_14_in16 = reg_0756;
    67: op1_14_in16 = reg_0939;
    92: op1_14_in16 = reg_0461;
    93: op1_14_in16 = reg_0566;
    94: op1_14_in16 = reg_0550;
    95: op1_14_in16 = reg_0775;
    97: op1_14_in16 = reg_1215;
    98: op1_14_in16 = reg_1458;
    99: op1_14_in16 = reg_0196;
    100: op1_14_in16 = reg_1092;
    101: op1_14_in16 = reg_1414;
    102: op1_14_in16 = reg_0631;
    103: op1_14_in16 = reg_0338;
    104: op1_14_in16 = reg_0266;
    105: op1_14_in16 = imem07_in[7:4];
    106: op1_14_in16 = reg_0576;
    107: op1_14_in16 = reg_0307;
    114: op1_14_in16 = reg_0307;
    37: op1_14_in16 = reg_0001;
    108: op1_14_in16 = reg_0921;
    109: op1_14_in16 = reg_1065;
    110: op1_14_in16 = imem01_in[7:4];
    111: op1_14_in16 = reg_0269;
    112: op1_14_in16 = reg_0267;
    113: op1_14_in16 = reg_0371;
    115: op1_14_in16 = imem06_in[3:0];
    116: op1_14_in16 = reg_0381;
    117: op1_14_in16 = reg_0173;
    118: op1_14_in16 = reg_0860;
    119: op1_14_in16 = reg_1351;
    47: op1_14_in16 = reg_0522;
    120: op1_14_in16 = reg_0874;
    121: op1_14_in16 = reg_1074;
    123: op1_14_in16 = reg_0923;
    124: op1_14_in16 = reg_0574;
    126: op1_14_in16 = reg_0268;
    127: op1_14_in16 = reg_0638;
    128: op1_14_in16 = reg_0712;
    129: op1_14_in16 = reg_0218;
    130: op1_14_in16 = reg_0802;
    default: op1_14_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv16 = 1;
    54: op1_14_inv16 = 1;
    75: op1_14_inv16 = 1;
    49: op1_14_inv16 = 1;
    69: op1_14_inv16 = 1;
    57: op1_14_inv16 = 1;
    68: op1_14_inv16 = 1;
    58: op1_14_inv16 = 1;
    70: op1_14_inv16 = 1;
    59: op1_14_inv16 = 1;
    88: op1_14_inv16 = 1;
    62: op1_14_inv16 = 1;
    81: op1_14_inv16 = 1;
    82: op1_14_inv16 = 1;
    52: op1_14_inv16 = 1;
    63: op1_14_inv16 = 1;
    83: op1_14_inv16 = 1;
    89: op1_14_inv16 = 1;
    66: op1_14_inv16 = 1;
    48: op1_14_inv16 = 1;
    91: op1_14_inv16 = 1;
    67: op1_14_inv16 = 1;
    93: op1_14_inv16 = 1;
    94: op1_14_inv16 = 1;
    97: op1_14_inv16 = 1;
    99: op1_14_inv16 = 1;
    100: op1_14_inv16 = 1;
    102: op1_14_inv16 = 1;
    103: op1_14_inv16 = 1;
    105: op1_14_inv16 = 1;
    109: op1_14_inv16 = 1;
    111: op1_14_inv16 = 1;
    115: op1_14_inv16 = 1;
    116: op1_14_inv16 = 1;
    117: op1_14_inv16 = 1;
    118: op1_14_inv16 = 1;
    119: op1_14_inv16 = 1;
    120: op1_14_inv16 = 1;
    124: op1_14_inv16 = 1;
    126: op1_14_inv16 = 1;
    127: op1_14_inv16 = 1;
    128: op1_14_inv16 = 1;
    default: op1_14_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in17 = reg_0722;
    53: op1_14_in17 = reg_0206;
    73: op1_14_in17 = reg_0122;
    55: op1_14_in17 = reg_0892;
    86: op1_14_in17 = reg_1372;
    74: op1_14_in17 = reg_1179;
    54: op1_14_in17 = reg_0890;
    75: op1_14_in17 = reg_0039;
    49: op1_14_in17 = reg_0998;
    69: op1_14_in17 = imem03_in[7:4];
    56: op1_14_in17 = reg_0095;
    50: op1_14_in17 = reg_0114;
    76: op1_14_in17 = reg_0968;
    71: op1_14_in17 = reg_0416;
    87: op1_14_in17 = imem03_in[3:0];
    57: op1_14_in17 = reg_0704;
    68: op1_14_in17 = reg_0757;
    77: op1_14_in17 = reg_1268;
    61: op1_14_in17 = reg_0611;
    78: op1_14_in17 = reg_1486;
    58: op1_14_in17 = reg_0495;
    70: op1_14_in17 = reg_0694;
    59: op1_14_in17 = reg_0646;
    79: op1_14_in17 = imem07_in[11:8];
    51: op1_14_in17 = reg_0608;
    60: op1_14_in17 = imem04_in[11:8];
    80: op1_14_in17 = reg_0310;
    88: op1_14_in17 = reg_0234;
    81: op1_14_in17 = reg_0373;
    82: op1_14_in17 = reg_0965;
    52: op1_14_in17 = reg_0921;
    63: op1_14_in17 = reg_0087;
    64: op1_14_in17 = reg_0904;
    83: op1_14_in17 = reg_1255;
    89: op1_14_in17 = reg_0470;
    84: op1_14_in17 = reg_1334;
    85: op1_14_in17 = reg_0387;
    65: op1_14_in17 = reg_0170;
    90: op1_14_in17 = reg_0350;
    100: op1_14_in17 = reg_0350;
    66: op1_14_in17 = reg_0472;
    48: op1_14_in17 = reg_0396;
    91: op1_14_in17 = reg_0388;
    46: op1_14_in17 = reg_0121;
    67: op1_14_in17 = reg_0938;
    92: op1_14_in17 = reg_0786;
    93: op1_14_in17 = reg_1402;
    94: op1_14_in17 = reg_0830;
    95: op1_14_in17 = reg_0284;
    97: op1_14_in17 = reg_0500;
    98: op1_14_in17 = reg_1450;
    99: op1_14_in17 = reg_0243;
    101: op1_14_in17 = reg_0478;
    102: op1_14_in17 = reg_1492;
    103: op1_14_in17 = reg_0209;
    104: op1_14_in17 = reg_1514;
    105: op1_14_in17 = reg_0461;
    106: op1_14_in17 = reg_0401;
    107: op1_14_in17 = reg_0560;
    37: op1_14_in17 = reg_0484;
    108: op1_14_in17 = reg_0224;
    109: op1_14_in17 = reg_0342;
    110: op1_14_in17 = imem01_in[15:12];
    111: op1_14_in17 = reg_0161;
    112: op1_14_in17 = reg_0635;
    113: op1_14_in17 = reg_0226;
    114: op1_14_in17 = reg_0473;
    115: op1_14_in17 = imem06_in[11:8];
    116: op1_14_in17 = reg_0802;
    117: op1_14_in17 = reg_0391;
    118: op1_14_in17 = reg_1501;
    119: op1_14_in17 = reg_1439;
    47: op1_14_in17 = reg_0289;
    120: op1_14_in17 = reg_0930;
    121: op1_14_in17 = reg_0533;
    122: op1_14_in17 = reg_0059;
    123: op1_14_in17 = reg_0139;
    124: op1_14_in17 = reg_0412;
    126: op1_14_in17 = reg_0368;
    127: op1_14_in17 = reg_0427;
    128: op1_14_in17 = reg_0532;
    129: op1_14_in17 = reg_0673;
    130: op1_14_in17 = reg_0227;
    default: op1_14_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv17 = 1;
    53: op1_14_inv17 = 1;
    74: op1_14_inv17 = 1;
    49: op1_14_inv17 = 1;
    76: op1_14_inv17 = 1;
    71: op1_14_inv17 = 1;
    87: op1_14_inv17 = 1;
    57: op1_14_inv17 = 1;
    77: op1_14_inv17 = 1;
    61: op1_14_inv17 = 1;
    70: op1_14_inv17 = 1;
    59: op1_14_inv17 = 1;
    60: op1_14_inv17 = 1;
    80: op1_14_inv17 = 1;
    88: op1_14_inv17 = 1;
    52: op1_14_inv17 = 1;
    63: op1_14_inv17 = 1;
    64: op1_14_inv17 = 1;
    83: op1_14_inv17 = 1;
    85: op1_14_inv17 = 1;
    65: op1_14_inv17 = 1;
    66: op1_14_inv17 = 1;
    48: op1_14_inv17 = 1;
    99: op1_14_inv17 = 1;
    103: op1_14_inv17 = 1;
    104: op1_14_inv17 = 1;
    105: op1_14_inv17 = 1;
    108: op1_14_inv17 = 1;
    111: op1_14_inv17 = 1;
    112: op1_14_inv17 = 1;
    114: op1_14_inv17 = 1;
    116: op1_14_inv17 = 1;
    117: op1_14_inv17 = 1;
    118: op1_14_inv17 = 1;
    120: op1_14_inv17 = 1;
    123: op1_14_inv17 = 1;
    124: op1_14_inv17 = 1;
    126: op1_14_inv17 = 1;
    127: op1_14_inv17 = 1;
    default: op1_14_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in18 = reg_0440;
    53: op1_14_in18 = reg_0974;
    73: op1_14_in18 = reg_1100;
    55: op1_14_in18 = reg_0673;
    86: op1_14_in18 = reg_1368;
    74: op1_14_in18 = reg_0270;
    47: op1_14_in18 = reg_0270;
    54: op1_14_in18 = reg_0130;
    75: op1_14_in18 = reg_0458;
    49: op1_14_in18 = reg_0867;
    57: op1_14_in18 = reg_0867;
    69: op1_14_in18 = reg_0640;
    56: op1_14_in18 = reg_0181;
    50: op1_14_in18 = reg_0361;
    76: op1_14_in18 = reg_1456;
    71: op1_14_in18 = reg_0072;
    91: op1_14_in18 = reg_0072;
    87: op1_14_in18 = reg_0480;
    68: op1_14_in18 = reg_0191;
    77: op1_14_in18 = reg_0992;
    61: op1_14_in18 = reg_0746;
    78: op1_14_in18 = reg_0576;
    58: op1_14_in18 = reg_0436;
    70: op1_14_in18 = reg_0493;
    59: op1_14_in18 = reg_1212;
    79: op1_14_in18 = reg_0186;
    51: op1_14_in18 = reg_1018;
    60: op1_14_in18 = reg_1257;
    80: op1_14_in18 = reg_0187;
    88: op1_14_in18 = reg_0375;
    81: op1_14_in18 = reg_0617;
    82: op1_14_in18 = reg_0349;
    52: op1_14_in18 = reg_0774;
    63: op1_14_in18 = reg_0520;
    64: op1_14_in18 = reg_0341;
    83: op1_14_in18 = reg_0093;
    120: op1_14_in18 = reg_0093;
    89: op1_14_in18 = imem05_in[3:0];
    84: op1_14_in18 = reg_0720;
    48: op1_14_in18 = reg_0720;
    85: op1_14_in18 = reg_0071;
    65: op1_14_in18 = reg_1345;
    90: op1_14_in18 = reg_0291;
    66: op1_14_in18 = reg_0494;
    46: op1_14_in18 = reg_0706;
    67: op1_14_in18 = reg_0477;
    92: op1_14_in18 = reg_0703;
    93: op1_14_in18 = reg_0938;
    94: op1_14_in18 = reg_0148;
    95: op1_14_in18 = reg_0441;
    97: op1_14_in18 = reg_0796;
    98: op1_14_in18 = reg_0126;
    99: op1_14_in18 = reg_0589;
    100: op1_14_in18 = reg_1280;
    101: op1_14_in18 = reg_1060;
    102: op1_14_in18 = reg_0802;
    103: op1_14_in18 = reg_0536;
    104: op1_14_in18 = reg_0601;
    105: op1_14_in18 = reg_1055;
    106: op1_14_in18 = reg_0047;
    107: op1_14_in18 = reg_0801;
    108: op1_14_in18 = reg_0287;
    109: op1_14_in18 = reg_0232;
    110: op1_14_in18 = reg_1290;
    111: op1_14_in18 = reg_1504;
    112: op1_14_in18 = reg_0871;
    113: op1_14_in18 = reg_0324;
    114: op1_14_in18 = reg_0829;
    115: op1_14_in18 = reg_0161;
    116: op1_14_in18 = reg_1098;
    117: op1_14_in18 = reg_0045;
    118: op1_14_in18 = reg_0780;
    119: op1_14_in18 = reg_0235;
    121: op1_14_in18 = reg_0900;
    128: op1_14_in18 = reg_0900;
    122: op1_14_in18 = reg_1321;
    123: op1_14_in18 = reg_0031;
    124: op1_14_in18 = reg_0407;
    126: op1_14_in18 = reg_0096;
    127: op1_14_in18 = reg_1369;
    129: op1_14_in18 = reg_0348;
    130: op1_14_in18 = reg_0104;
    default: op1_14_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv18 = 1;
    53: op1_14_inv18 = 1;
    86: op1_14_inv18 = 1;
    74: op1_14_inv18 = 1;
    56: op1_14_inv18 = 1;
    71: op1_14_inv18 = 1;
    77: op1_14_inv18 = 1;
    58: op1_14_inv18 = 1;
    70: op1_14_inv18 = 1;
    59: op1_14_inv18 = 1;
    51: op1_14_inv18 = 1;
    60: op1_14_inv18 = 1;
    88: op1_14_inv18 = 1;
    82: op1_14_inv18 = 1;
    63: op1_14_inv18 = 1;
    83: op1_14_inv18 = 1;
    84: op1_14_inv18 = 1;
    90: op1_14_inv18 = 1;
    48: op1_14_inv18 = 1;
    91: op1_14_inv18 = 1;
    67: op1_14_inv18 = 1;
    92: op1_14_inv18 = 1;
    93: op1_14_inv18 = 1;
    94: op1_14_inv18 = 1;
    95: op1_14_inv18 = 1;
    97: op1_14_inv18 = 1;
    98: op1_14_inv18 = 1;
    101: op1_14_inv18 = 1;
    102: op1_14_inv18 = 1;
    103: op1_14_inv18 = 1;
    107: op1_14_inv18 = 1;
    109: op1_14_inv18 = 1;
    111: op1_14_inv18 = 1;
    112: op1_14_inv18 = 1;
    114: op1_14_inv18 = 1;
    116: op1_14_inv18 = 1;
    118: op1_14_inv18 = 1;
    47: op1_14_inv18 = 1;
    120: op1_14_inv18 = 1;
    123: op1_14_inv18 = 1;
    124: op1_14_inv18 = 1;
    126: op1_14_inv18 = 1;
    127: op1_14_inv18 = 1;
    default: op1_14_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in19 = reg_0071;
    53: op1_14_in19 = reg_1035;
    73: op1_14_in19 = reg_0785;
    55: op1_14_in19 = reg_0156;
    86: op1_14_in19 = imem04_in[11:8];
    74: op1_14_in19 = reg_0046;
    54: op1_14_in19 = reg_0960;
    75: op1_14_in19 = reg_0399;
    49: op1_14_in19 = reg_0851;
    80: op1_14_in19 = reg_0851;
    69: op1_14_in19 = reg_0638;
    56: op1_14_in19 = reg_0064;
    50: op1_14_in19 = reg_0228;
    76: op1_14_in19 = reg_0365;
    71: op1_14_in19 = reg_0059;
    87: op1_14_in19 = reg_1139;
    57: op1_14_in19 = reg_0299;
    68: op1_14_in19 = reg_0227;
    77: op1_14_in19 = imem05_in[15:12];
    61: op1_14_in19 = reg_1151;
    78: op1_14_in19 = reg_0197;
    58: op1_14_in19 = reg_0970;
    70: op1_14_in19 = reg_1339;
    59: op1_14_in19 = reg_0131;
    79: op1_14_in19 = reg_0225;
    51: op1_14_in19 = reg_0589;
    60: op1_14_in19 = reg_0798;
    88: op1_14_in19 = reg_1516;
    81: op1_14_in19 = reg_0526;
    82: op1_14_in19 = reg_0957;
    52: op1_14_in19 = reg_0030;
    63: op1_14_in19 = reg_0484;
    64: op1_14_in19 = reg_0305;
    83: op1_14_in19 = reg_0549;
    89: op1_14_in19 = reg_1299;
    84: op1_14_in19 = reg_0780;
    85: op1_14_in19 = reg_0203;
    65: op1_14_in19 = reg_0489;
    90: op1_14_in19 = reg_0288;
    66: op1_14_in19 = reg_0054;
    48: op1_14_in19 = reg_0371;
    91: op1_14_in19 = reg_0057;
    46: op1_14_in19 = reg_0378;
    67: op1_14_in19 = reg_0367;
    92: op1_14_in19 = reg_0366;
    93: op1_14_in19 = reg_0418;
    94: op1_14_in19 = reg_0146;
    95: op1_14_in19 = reg_0408;
    97: op1_14_in19 = reg_0094;
    98: op1_14_in19 = reg_0112;
    99: op1_14_in19 = reg_0603;
    104: op1_14_in19 = reg_0603;
    100: op1_14_in19 = reg_0427;
    101: op1_14_in19 = reg_0140;
    102: op1_14_in19 = reg_1091;
    103: op1_14_in19 = reg_1502;
    105: op1_14_in19 = reg_0667;
    106: op1_14_in19 = reg_0553;
    110: op1_14_in19 = reg_0553;
    107: op1_14_in19 = reg_0695;
    108: op1_14_in19 = reg_0442;
    109: op1_14_in19 = reg_0582;
    111: op1_14_in19 = reg_0109;
    112: op1_14_in19 = reg_1152;
    113: op1_14_in19 = reg_1183;
    114: op1_14_in19 = reg_0745;
    115: op1_14_in19 = reg_1209;
    116: op1_14_in19 = reg_0294;
    117: op1_14_in19 = reg_1402;
    118: op1_14_in19 = reg_0714;
    119: op1_14_in19 = reg_0002;
    47: op1_14_in19 = reg_0269;
    120: op1_14_in19 = reg_0743;
    121: op1_14_in19 = reg_0878;
    122: op1_14_in19 = reg_0122;
    123: op1_14_in19 = reg_0287;
    124: op1_14_in19 = reg_0097;
    126: op1_14_in19 = reg_0904;
    127: op1_14_in19 = reg_0181;
    128: op1_14_in19 = reg_0429;
    129: op1_14_in19 = reg_1216;
    130: op1_14_in19 = reg_0049;
    default: op1_14_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv19 = 1;
    74: op1_14_inv19 = 1;
    54: op1_14_inv19 = 1;
    49: op1_14_inv19 = 1;
    69: op1_14_inv19 = 1;
    50: op1_14_inv19 = 1;
    76: op1_14_inv19 = 1;
    71: op1_14_inv19 = 1;
    68: op1_14_inv19 = 1;
    77: op1_14_inv19 = 1;
    61: op1_14_inv19 = 1;
    70: op1_14_inv19 = 1;
    88: op1_14_inv19 = 1;
    81: op1_14_inv19 = 1;
    82: op1_14_inv19 = 1;
    52: op1_14_inv19 = 1;
    65: op1_14_inv19 = 1;
    90: op1_14_inv19 = 1;
    66: op1_14_inv19 = 1;
    91: op1_14_inv19 = 1;
    67: op1_14_inv19 = 1;
    93: op1_14_inv19 = 1;
    95: op1_14_inv19 = 1;
    97: op1_14_inv19 = 1;
    98: op1_14_inv19 = 1;
    101: op1_14_inv19 = 1;
    102: op1_14_inv19 = 1;
    104: op1_14_inv19 = 1;
    107: op1_14_inv19 = 1;
    108: op1_14_inv19 = 1;
    109: op1_14_inv19 = 1;
    111: op1_14_inv19 = 1;
    112: op1_14_inv19 = 1;
    113: op1_14_inv19 = 1;
    47: op1_14_inv19 = 1;
    120: op1_14_inv19 = 1;
    122: op1_14_inv19 = 1;
    123: op1_14_inv19 = 1;
    124: op1_14_inv19 = 1;
    126: op1_14_inv19 = 1;
    127: op1_14_inv19 = 1;
    128: op1_14_inv19 = 1;
    130: op1_14_inv19 = 1;
    default: op1_14_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in20 = reg_1321;
    53: op1_14_in20 = reg_0979;
    73: op1_14_in20 = reg_0335;
    55: op1_14_in20 = reg_0921;
    86: op1_14_in20 = reg_1083;
    74: op1_14_in20 = reg_0212;
    54: op1_14_in20 = reg_0859;
    75: op1_14_in20 = reg_1064;
    49: op1_14_in20 = reg_0156;
    69: op1_14_in20 = reg_1325;
    56: op1_14_in20 = reg_0033;
    50: op1_14_in20 = reg_0001;
    76: op1_14_in20 = reg_0092;
    71: op1_14_in20 = reg_1322;
    87: op1_14_in20 = reg_0443;
    57: op1_14_in20 = reg_0187;
    68: op1_14_in20 = reg_0154;
    77: op1_14_in20 = reg_0794;
    61: op1_14_in20 = reg_0968;
    78: op1_14_in20 = reg_1373;
    58: op1_14_in20 = reg_0055;
    70: op1_14_in20 = reg_1338;
    59: op1_14_in20 = reg_0182;
    79: op1_14_in20 = reg_0309;
    51: op1_14_in20 = reg_0473;
    60: op1_14_in20 = reg_0932;
    80: op1_14_in20 = reg_1350;
    88: op1_14_in20 = reg_1314;
    81: op1_14_in20 = reg_0568;
    82: op1_14_in20 = reg_0246;
    52: op1_14_in20 = reg_0287;
    64: op1_14_in20 = reg_0319;
    83: op1_14_in20 = reg_0787;
    89: op1_14_in20 = reg_0251;
    84: op1_14_in20 = reg_0115;
    48: op1_14_in20 = reg_0115;
    85: op1_14_in20 = reg_0075;
    65: op1_14_in20 = reg_0030;
    90: op1_14_in20 = reg_1144;
    66: op1_14_in20 = reg_0970;
    91: op1_14_in20 = reg_1324;
    46: op1_14_in20 = reg_0232;
    67: op1_14_in20 = reg_0090;
    92: op1_14_in20 = reg_0741;
    93: op1_14_in20 = reg_0873;
    94: op1_14_in20 = reg_0403;
    95: op1_14_in20 = reg_0623;
    97: op1_14_in20 = reg_1147;
    98: op1_14_in20 = reg_0631;
    99: op1_14_in20 = reg_0120;
    122: op1_14_in20 = reg_0120;
    100: op1_14_in20 = imem04_in[3:0];
    101: op1_14_in20 = reg_0170;
    102: op1_14_in20 = reg_0479;
    103: op1_14_in20 = reg_0210;
    104: op1_14_in20 = imem06_in[3:0];
    105: op1_14_in20 = reg_0703;
    106: op1_14_in20 = reg_0548;
    112: op1_14_in20 = reg_0548;
    107: op1_14_in20 = imem02_in[11:8];
    108: op1_14_in20 = reg_0137;
    109: op1_14_in20 = reg_0262;
    110: op1_14_in20 = reg_0550;
    111: op1_14_in20 = reg_0717;
    113: op1_14_in20 = imem07_in[3:0];
    114: op1_14_in20 = reg_0379;
    115: op1_14_in20 = reg_0960;
    116: op1_14_in20 = reg_0217;
    117: op1_14_in20 = reg_0938;
    118: op1_14_in20 = reg_0637;
    119: op1_14_in20 = reg_1182;
    47: op1_14_in20 = reg_0213;
    120: op1_14_in20 = reg_0830;
    121: op1_14_in20 = reg_0711;
    123: op1_14_in20 = reg_0285;
    124: op1_14_in20 = reg_1419;
    126: op1_14_in20 = reg_0650;
    127: op1_14_in20 = reg_1339;
    128: op1_14_in20 = reg_0971;
    129: op1_14_in20 = reg_0034;
    130: op1_14_in20 = reg_0709;
    default: op1_14_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv20 = 1;
    86: op1_14_inv20 = 1;
    75: op1_14_inv20 = 1;
    57: op1_14_inv20 = 1;
    77: op1_14_inv20 = 1;
    61: op1_14_inv20 = 1;
    70: op1_14_inv20 = 1;
    79: op1_14_inv20 = 1;
    51: op1_14_inv20 = 1;
    81: op1_14_inv20 = 1;
    82: op1_14_inv20 = 1;
    52: op1_14_inv20 = 1;
    64: op1_14_inv20 = 1;
    89: op1_14_inv20 = 1;
    84: op1_14_inv20 = 1;
    65: op1_14_inv20 = 1;
    48: op1_14_inv20 = 1;
    91: op1_14_inv20 = 1;
    93: op1_14_inv20 = 1;
    99: op1_14_inv20 = 1;
    102: op1_14_inv20 = 1;
    107: op1_14_inv20 = 1;
    108: op1_14_inv20 = 1;
    109: op1_14_inv20 = 1;
    111: op1_14_inv20 = 1;
    113: op1_14_inv20 = 1;
    114: op1_14_inv20 = 1;
    117: op1_14_inv20 = 1;
    118: op1_14_inv20 = 1;
    47: op1_14_inv20 = 1;
    120: op1_14_inv20 = 1;
    122: op1_14_inv20 = 1;
    123: op1_14_inv20 = 1;
    127: op1_14_inv20 = 1;
    default: op1_14_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in21 = reg_0089;
    53: op1_14_in21 = reg_0907;
    73: op1_14_in21 = reg_0372;
    55: op1_14_in21 = reg_0169;
    86: op1_14_in21 = reg_0552;
    74: op1_14_in21 = reg_0022;
    54: op1_14_in21 = reg_0115;
    75: op1_14_in21 = reg_0120;
    49: op1_14_in21 = imem07_in[7:4];
    69: op1_14_in21 = reg_0789;
    56: op1_14_in21 = reg_0792;
    50: op1_14_in21 = reg_0052;
    76: op1_14_in21 = reg_0724;
    71: op1_14_in21 = reg_0723;
    87: op1_14_in21 = imem04_in[15:12];
    100: op1_14_in21 = imem04_in[15:12];
    57: op1_14_in21 = reg_0170;
    68: op1_14_in21 = reg_0377;
    77: op1_14_in21 = reg_0303;
    61: op1_14_in21 = reg_0430;
    78: op1_14_in21 = reg_0601;
    58: op1_14_in21 = reg_0897;
    70: op1_14_in21 = reg_0577;
    59: op1_14_in21 = reg_0315;
    79: op1_14_in21 = reg_0297;
    51: op1_14_in21 = reg_0474;
    60: op1_14_in21 = reg_0451;
    80: op1_14_in21 = reg_1347;
    101: op1_14_in21 = reg_1347;
    88: op1_14_in21 = reg_0597;
    81: op1_14_in21 = reg_0165;
    82: op1_14_in21 = reg_0329;
    52: op1_14_in21 = reg_0285;
    64: op1_14_in21 = reg_0262;
    83: op1_14_in21 = reg_0241;
    89: op1_14_in21 = reg_0833;
    84: op1_14_in21 = reg_0373;
    85: op1_14_in21 = reg_0917;
    65: op1_14_in21 = reg_0284;
    90: op1_14_in21 = reg_1372;
    66: op1_14_in21 = reg_0105;
    48: op1_14_in21 = reg_0671;
    91: op1_14_in21 = reg_1322;
    46: op1_14_in21 = reg_0049;
    67: op1_14_in21 = reg_0197;
    92: op1_14_in21 = reg_0408;
    93: op1_14_in21 = reg_0872;
    94: op1_14_in21 = reg_0385;
    95: op1_14_in21 = reg_0618;
    97: op1_14_in21 = reg_0599;
    98: op1_14_in21 = reg_0380;
    99: op1_14_in21 = reg_0397;
    102: op1_14_in21 = reg_0999;
    103: op1_14_in21 = reg_0986;
    104: op1_14_in21 = reg_1467;
    105: op1_14_in21 = reg_0457;
    106: op1_14_in21 = reg_0609;
    110: op1_14_in21 = reg_0609;
    107: op1_14_in21 = reg_0024;
    108: op1_14_in21 = reg_0087;
    109: op1_14_in21 = reg_0487;
    111: op1_14_in21 = reg_0636;
    112: op1_14_in21 = reg_1474;
    113: op1_14_in21 = reg_0922;
    114: op1_14_in21 = reg_0802;
    115: op1_14_in21 = reg_0974;
    116: op1_14_in21 = reg_0235;
    117: op1_14_in21 = reg_0937;
    118: op1_14_in21 = reg_0619;
    47: op1_14_in21 = imem07_in[15:12];
    120: op1_14_in21 = reg_0798;
    121: op1_14_in21 = reg_0824;
    122: op1_14_in21 = reg_0902;
    123: op1_14_in21 = reg_0739;
    124: op1_14_in21 = reg_0268;
    126: op1_14_in21 = reg_0445;
    127: op1_14_in21 = imem04_in[3:0];
    128: op1_14_in21 = reg_1450;
    129: op1_14_in21 = reg_0493;
    130: op1_14_in21 = reg_0507;
    default: op1_14_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv21 = 1;
    73: op1_14_inv21 = 1;
    55: op1_14_inv21 = 1;
    75: op1_14_inv21 = 1;
    69: op1_14_inv21 = 1;
    56: op1_14_inv21 = 1;
    50: op1_14_inv21 = 1;
    76: op1_14_inv21 = 1;
    87: op1_14_inv21 = 1;
    57: op1_14_inv21 = 1;
    68: op1_14_inv21 = 1;
    61: op1_14_inv21 = 1;
    58: op1_14_inv21 = 1;
    59: op1_14_inv21 = 1;
    79: op1_14_inv21 = 1;
    60: op1_14_inv21 = 1;
    88: op1_14_inv21 = 1;
    83: op1_14_inv21 = 1;
    65: op1_14_inv21 = 1;
    48: op1_14_inv21 = 1;
    92: op1_14_inv21 = 1;
    95: op1_14_inv21 = 1;
    97: op1_14_inv21 = 1;
    98: op1_14_inv21 = 1;
    99: op1_14_inv21 = 1;
    100: op1_14_inv21 = 1;
    101: op1_14_inv21 = 1;
    102: op1_14_inv21 = 1;
    105: op1_14_inv21 = 1;
    106: op1_14_inv21 = 1;
    111: op1_14_inv21 = 1;
    112: op1_14_inv21 = 1;
    113: op1_14_inv21 = 1;
    116: op1_14_inv21 = 1;
    117: op1_14_inv21 = 1;
    121: op1_14_inv21 = 1;
    122: op1_14_inv21 = 1;
    123: op1_14_inv21 = 1;
    124: op1_14_inv21 = 1;
    129: op1_14_inv21 = 1;
    130: op1_14_inv21 = 1;
    default: op1_14_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in22 = reg_0027;
    53: op1_14_in22 = reg_0730;
    73: op1_14_in22 = reg_0166;
    55: op1_14_in22 = reg_0779;
    49: op1_14_in22 = reg_0779;
    86: op1_14_in22 = reg_0488;
    74: op1_14_in22 = imem07_in[7:4];
    54: op1_14_in22 = reg_0110;
    75: op1_14_in22 = reg_0907;
    69: op1_14_in22 = reg_0142;
    56: op1_14_in22 = reg_0794;
    50: op1_14_in22 = reg_0518;
    76: op1_14_in22 = reg_0896;
    71: op1_14_in22 = reg_1291;
    87: op1_14_in22 = reg_1312;
    57: op1_14_in22 = reg_0159;
    80: op1_14_in22 = reg_0159;
    68: op1_14_in22 = reg_0557;
    77: op1_14_in22 = reg_0300;
    61: op1_14_in22 = reg_0728;
    78: op1_14_in22 = reg_0130;
    58: op1_14_in22 = reg_0711;
    70: op1_14_in22 = reg_1077;
    59: op1_14_in22 = reg_0539;
    79: op1_14_in22 = reg_0223;
    51: op1_14_in22 = reg_0989;
    60: op1_14_in22 = reg_0487;
    64: op1_14_in22 = reg_0487;
    88: op1_14_in22 = reg_0350;
    81: op1_14_in22 = reg_0271;
    82: op1_14_in22 = reg_1231;
    52: op1_14_in22 = reg_0740;
    83: op1_14_in22 = reg_0968;
    89: op1_14_in22 = reg_1431;
    84: op1_14_in22 = reg_0622;
    85: op1_14_in22 = reg_0679;
    65: op1_14_in22 = reg_0285;
    90: op1_14_in22 = reg_0264;
    66: op1_14_in22 = reg_0380;
    48: op1_14_in22 = reg_0669;
    91: op1_14_in22 = reg_0653;
    46: op1_14_in22 = reg_0600;
    67: op1_14_in22 = reg_0207;
    92: op1_14_in22 = reg_0623;
    93: op1_14_in22 = reg_0196;
    94: op1_14_in22 = reg_0363;
    95: op1_14_in22 = reg_0100;
    97: op1_14_in22 = reg_0537;
    98: op1_14_in22 = reg_0473;
    99: op1_14_in22 = reg_0925;
    100: op1_14_in22 = reg_1368;
    101: op1_14_in22 = reg_0156;
    47: op1_14_in22 = reg_0156;
    102: op1_14_in22 = imem03_in[11:8];
    103: op1_14_in22 = reg_0604;
    104: op1_14_in22 = reg_0860;
    115: op1_14_in22 = reg_0860;
    105: op1_14_in22 = reg_0774;
    106: op1_14_in22 = reg_0242;
    107: op1_14_in22 = reg_0068;
    121: op1_14_in22 = reg_0068;
    108: op1_14_in22 = reg_0124;
    109: op1_14_in22 = reg_0719;
    110: op1_14_in22 = reg_1473;
    111: op1_14_in22 = reg_0398;
    112: op1_14_in22 = reg_0715;
    113: op1_14_in22 = reg_0135;
    114: op1_14_in22 = reg_1078;
    116: op1_14_in22 = reg_0677;
    117: op1_14_in22 = reg_0303;
    118: op1_14_in22 = reg_0571;
    120: op1_14_in22 = reg_0819;
    122: op1_14_in22 = reg_0787;
    123: op1_14_in22 = reg_0102;
    124: op1_14_in22 = reg_0862;
    126: op1_14_in22 = reg_1402;
    127: op1_14_in22 = imem04_in[7:4];
    128: op1_14_in22 = reg_0106;
    129: op1_14_in22 = reg_0535;
    130: op1_14_in22 = reg_0177;
    default: op1_14_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv22 = 1;
    86: op1_14_inv22 = 1;
    75: op1_14_inv22 = 1;
    49: op1_14_inv22 = 1;
    69: op1_14_inv22 = 1;
    56: op1_14_inv22 = 1;
    71: op1_14_inv22 = 1;
    87: op1_14_inv22 = 1;
    57: op1_14_inv22 = 1;
    59: op1_14_inv22 = 1;
    51: op1_14_inv22 = 1;
    60: op1_14_inv22 = 1;
    81: op1_14_inv22 = 1;
    52: op1_14_inv22 = 1;
    64: op1_14_inv22 = 1;
    83: op1_14_inv22 = 1;
    85: op1_14_inv22 = 1;
    65: op1_14_inv22 = 1;
    66: op1_14_inv22 = 1;
    95: op1_14_inv22 = 1;
    97: op1_14_inv22 = 1;
    99: op1_14_inv22 = 1;
    100: op1_14_inv22 = 1;
    104: op1_14_inv22 = 1;
    106: op1_14_inv22 = 1;
    107: op1_14_inv22 = 1;
    110: op1_14_inv22 = 1;
    112: op1_14_inv22 = 1;
    114: op1_14_inv22 = 1;
    118: op1_14_inv22 = 1;
    120: op1_14_inv22 = 1;
    121: op1_14_inv22 = 1;
    122: op1_14_inv22 = 1;
    127: op1_14_inv22 = 1;
    130: op1_14_inv22 = 1;
    default: op1_14_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in23 = reg_0005;
    53: op1_14_in23 = reg_0870;
    99: op1_14_in23 = reg_0870;
    73: op1_14_in23 = reg_1473;
    55: op1_14_in23 = reg_0664;
    86: op1_14_in23 = reg_0796;
    74: op1_14_in23 = reg_0490;
    54: op1_14_in23 = reg_0109;
    75: op1_14_in23 = reg_1420;
    49: op1_14_in23 = reg_0465;
    69: op1_14_in23 = reg_1003;
    56: op1_14_in23 = reg_1059;
    50: op1_14_in23 = reg_0520;
    76: op1_14_in23 = reg_0079;
    71: op1_14_in23 = reg_0930;
    87: op1_14_in23 = reg_0032;
    57: op1_14_in23 = reg_0156;
    68: op1_14_in23 = reg_1033;
    77: op1_14_in23 = reg_1486;
    61: op1_14_in23 = reg_0401;
    78: op1_14_in23 = reg_0243;
    93: op1_14_in23 = reg_0243;
    58: op1_14_in23 = reg_0008;
    70: op1_14_in23 = reg_1065;
    59: op1_14_in23 = reg_0183;
    79: op1_14_in23 = reg_1094;
    51: op1_14_in23 = reg_0981;
    60: op1_14_in23 = reg_0837;
    80: op1_14_in23 = reg_0157;
    88: op1_14_in23 = reg_1139;
    81: op1_14_in23 = reg_0034;
    82: op1_14_in23 = reg_1199;
    52: op1_14_in23 = reg_0621;
    65: op1_14_in23 = reg_0621;
    64: op1_14_in23 = reg_0237;
    83: op1_14_in23 = reg_0430;
    89: op1_14_in23 = reg_1169;
    126: op1_14_in23 = reg_1169;
    84: op1_14_in23 = reg_0619;
    85: op1_14_in23 = reg_0161;
    90: op1_14_in23 = reg_0252;
    66: op1_14_in23 = reg_0381;
    48: op1_14_in23 = reg_0634;
    91: op1_14_in23 = reg_0677;
    46: op1_14_in23 = reg_0179;
    67: op1_14_in23 = imem06_in[3:0];
    92: op1_14_in23 = reg_0228;
    94: op1_14_in23 = reg_0901;
    95: op1_14_in23 = reg_0518;
    97: op1_14_in23 = reg_0199;
    98: op1_14_in23 = reg_0829;
    100: op1_14_in23 = reg_0493;
    101: op1_14_in23 = reg_0923;
    102: op1_14_in23 = reg_0185;
    103: op1_14_in23 = reg_1104;
    104: op1_14_in23 = reg_1501;
    105: op1_14_in23 = reg_0665;
    106: op1_14_in23 = reg_1474;
    107: op1_14_in23 = reg_0009;
    121: op1_14_in23 = reg_0009;
    109: op1_14_in23 = reg_1146;
    110: op1_14_in23 = reg_0612;
    111: op1_14_in23 = reg_0527;
    112: op1_14_in23 = reg_0469;
    113: op1_14_in23 = reg_1440;
    114: op1_14_in23 = reg_0217;
    115: op1_14_in23 = reg_0863;
    116: op1_14_in23 = reg_0759;
    117: op1_14_in23 = reg_0090;
    118: op1_14_in23 = reg_0570;
    47: op1_14_in23 = reg_0140;
    120: op1_14_in23 = reg_0438;
    122: op1_14_in23 = reg_0609;
    123: op1_14_in23 = reg_0114;
    124: op1_14_in23 = reg_0719;
    127: op1_14_in23 = imem04_in[11:8];
    128: op1_14_in23 = reg_1433;
    129: op1_14_in23 = reg_0694;
    130: op1_14_in23 = reg_0600;
    default: op1_14_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv23 = 1;
    55: op1_14_inv23 = 1;
    74: op1_14_inv23 = 1;
    75: op1_14_inv23 = 1;
    49: op1_14_inv23 = 1;
    50: op1_14_inv23 = 1;
    87: op1_14_inv23 = 1;
    57: op1_14_inv23 = 1;
    68: op1_14_inv23 = 1;
    61: op1_14_inv23 = 1;
    79: op1_14_inv23 = 1;
    51: op1_14_inv23 = 1;
    80: op1_14_inv23 = 1;
    88: op1_14_inv23 = 1;
    82: op1_14_inv23 = 1;
    52: op1_14_inv23 = 1;
    64: op1_14_inv23 = 1;
    84: op1_14_inv23 = 1;
    85: op1_14_inv23 = 1;
    48: op1_14_inv23 = 1;
    91: op1_14_inv23 = 1;
    46: op1_14_inv23 = 1;
    92: op1_14_inv23 = 1;
    95: op1_14_inv23 = 1;
    97: op1_14_inv23 = 1;
    100: op1_14_inv23 = 1;
    101: op1_14_inv23 = 1;
    102: op1_14_inv23 = 1;
    105: op1_14_inv23 = 1;
    106: op1_14_inv23 = 1;
    107: op1_14_inv23 = 1;
    109: op1_14_inv23 = 1;
    112: op1_14_inv23 = 1;
    113: op1_14_inv23 = 1;
    116: op1_14_inv23 = 1;
    117: op1_14_inv23 = 1;
    118: op1_14_inv23 = 1;
    120: op1_14_inv23 = 1;
    127: op1_14_inv23 = 1;
    130: op1_14_inv23 = 1;
    default: op1_14_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in24 = reg_0917;
    53: op1_14_in24 = reg_0141;
    73: op1_14_in24 = reg_0612;
    55: op1_14_in24 = reg_0287;
    86: op1_14_in24 = reg_0598;
    74: op1_14_in24 = reg_0491;
    54: op1_14_in24 = reg_0264;
    75: op1_14_in24 = reg_0860;
    49: op1_14_in24 = reg_0665;
    69: op1_14_in24 = reg_0349;
    56: op1_14_in24 = reg_0833;
    76: op1_14_in24 = reg_0277;
    71: op1_14_in24 = reg_0553;
    87: op1_14_in24 = reg_1369;
    57: op1_14_in24 = reg_0140;
    68: op1_14_in24 = reg_0638;
    77: op1_14_in24 = reg_1484;
    61: op1_14_in24 = reg_0386;
    78: op1_14_in24 = reg_1348;
    58: op1_14_in24 = reg_0829;
    70: op1_14_in24 = reg_0466;
    59: op1_14_in24 = reg_0477;
    79: op1_14_in24 = reg_0779;
    101: op1_14_in24 = reg_0779;
    51: op1_14_in24 = reg_0432;
    60: op1_14_in24 = reg_0836;
    80: op1_14_in24 = reg_0441;
    88: op1_14_in24 = reg_0288;
    81: op1_14_in24 = reg_0461;
    82: op1_14_in24 = reg_0481;
    52: op1_14_in24 = reg_0618;
    64: op1_14_in24 = reg_0016;
    83: op1_14_in24 = reg_0362;
    89: op1_14_in24 = reg_0996;
    84: op1_14_in24 = reg_0569;
    85: op1_14_in24 = reg_1511;
    65: op1_14_in24 = reg_0591;
    90: op1_14_in24 = reg_0462;
    66: op1_14_in24 = reg_0056;
    48: op1_14_in24 = reg_0635;
    91: op1_14_in24 = reg_1513;
    46: op1_14_in24 = imem03_in[11:8];
    67: op1_14_in24 = imem06_in[11:8];
    92: op1_14_in24 = reg_0050;
    93: op1_14_in24 = reg_0602;
    94: op1_14_in24 = reg_0078;
    97: op1_14_in24 = reg_0454;
    98: op1_14_in24 = reg_1098;
    99: op1_14_in24 = reg_0782;
    100: op1_14_in24 = reg_0088;
    102: op1_14_in24 = reg_1063;
    103: op1_14_in24 = reg_0182;
    104: op1_14_in24 = reg_0714;
    105: op1_14_in24 = reg_0663;
    106: op1_14_in24 = reg_0468;
    107: op1_14_in24 = reg_0168;
    109: op1_14_in24 = reg_1189;
    110: op1_14_in24 = reg_0469;
    111: op1_14_in24 = reg_0568;
    112: op1_14_in24 = reg_0968;
    113: op1_14_in24 = reg_1094;
    114: op1_14_in24 = reg_0069;
    115: op1_14_in24 = reg_0265;
    116: op1_14_in24 = reg_0233;
    117: op1_14_in24 = reg_0794;
    118: op1_14_in24 = reg_1225;
    47: op1_14_in24 = reg_0031;
    120: op1_14_in24 = reg_1457;
    121: op1_14_in24 = reg_0632;
    122: op1_14_in24 = reg_0238;
    123: op1_14_in24 = reg_0028;
    124: op1_14_in24 = reg_0904;
    126: op1_14_in24 = reg_1163;
    127: op1_14_in24 = reg_0164;
    128: op1_14_in24 = reg_0876;
    129: op1_14_in24 = reg_1258;
    130: op1_14_in24 = reg_0312;
    default: op1_14_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_14_inv24 = 1;
    55: op1_14_inv24 = 1;
    86: op1_14_inv24 = 1;
    71: op1_14_inv24 = 1;
    87: op1_14_inv24 = 1;
    57: op1_14_inv24 = 1;
    68: op1_14_inv24 = 1;
    78: op1_14_inv24 = 1;
    51: op1_14_inv24 = 1;
    60: op1_14_inv24 = 1;
    82: op1_14_inv24 = 1;
    64: op1_14_inv24 = 1;
    83: op1_14_inv24 = 1;
    89: op1_14_inv24 = 1;
    90: op1_14_inv24 = 1;
    91: op1_14_inv24 = 1;
    67: op1_14_inv24 = 1;
    92: op1_14_inv24 = 1;
    93: op1_14_inv24 = 1;
    98: op1_14_inv24 = 1;
    102: op1_14_inv24 = 1;
    105: op1_14_inv24 = 1;
    114: op1_14_inv24 = 1;
    117: op1_14_inv24 = 1;
    118: op1_14_inv24 = 1;
    122: op1_14_inv24 = 1;
    126: op1_14_inv24 = 1;
    127: op1_14_inv24 = 1;
    128: op1_14_inv24 = 1;
    default: op1_14_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in25 = reg_1100;
    53: op1_14_in25 = reg_0374;
    73: op1_14_in25 = reg_0715;
    55: op1_14_in25 = reg_0442;
    86: op1_14_in25 = reg_1041;
    74: op1_14_in25 = reg_0298;
    54: op1_14_in25 = reg_0568;
    75: op1_14_in25 = reg_0720;
    49: op1_14_in25 = reg_0741;
    69: op1_14_in25 = reg_1199;
    56: op1_14_in25 = reg_0832;
    76: op1_14_in25 = reg_0679;
    71: op1_14_in25 = reg_0260;
    87: op1_14_in25 = reg_1368;
    57: op1_14_in25 = reg_0777;
    68: op1_14_in25 = reg_0000;
    77: op1_14_in25 = reg_0864;
    61: op1_14_in25 = reg_0092;
    78: op1_14_in25 = reg_0589;
    58: op1_14_in25 = reg_0068;
    70: op1_14_in25 = reg_0676;
    59: op1_14_in25 = reg_0872;
    79: op1_14_in25 = reg_0287;
    105: op1_14_in25 = reg_0287;
    51: op1_14_in25 = reg_0970;
    60: op1_14_in25 = reg_0096;
    80: op1_14_in25 = reg_0740;
    88: op1_14_in25 = reg_1282;
    81: op1_14_in25 = reg_1315;
    82: op1_14_in25 = reg_0790;
    52: op1_14_in25 = reg_0593;
    64: op1_14_in25 = reg_0020;
    83: op1_14_in25 = reg_0091;
    89: op1_14_in25 = reg_0648;
    84: op1_14_in25 = reg_0570;
    85: op1_14_in25 = reg_0609;
    65: op1_14_in25 = reg_0592;
    90: op1_14_in25 = reg_1083;
    66: op1_14_in25 = reg_0878;
    48: op1_14_in25 = reg_0586;
    91: op1_14_in25 = reg_0258;
    46: op1_14_in25 = reg_0627;
    67: op1_14_in25 = reg_0195;
    92: op1_14_in25 = reg_0002;
    93: op1_14_in25 = reg_1346;
    94: op1_14_in25 = reg_0896;
    97: op1_14_in25 = reg_1419;
    98: op1_14_in25 = imem03_in[11:8];
    99: op1_14_in25 = reg_0714;
    100: op1_14_in25 = reg_0034;
    101: op1_14_in25 = reg_0665;
    102: op1_14_in25 = reg_0177;
    103: op1_14_in25 = reg_0045;
    104: op1_14_in25 = reg_1303;
    106: op1_14_in25 = reg_0966;
    107: op1_14_in25 = reg_0750;
    109: op1_14_in25 = reg_0064;
    110: op1_14_in25 = reg_1452;
    111: op1_14_in25 = reg_0569;
    112: op1_14_in25 = reg_0148;
    113: op1_14_in25 = reg_0774;
    114: op1_14_in25 = reg_0279;
    115: op1_14_in25 = reg_0716;
    116: op1_14_in25 = reg_0220;
    117: op1_14_in25 = reg_0492;
    118: op1_14_in25 = reg_0296;
    47: op1_14_in25 = reg_0284;
    120: op1_14_in25 = reg_0726;
    121: op1_14_in25 = reg_0328;
    122: op1_14_in25 = reg_1457;
    123: op1_14_in25 = reg_0520;
    124: op1_14_in25 = reg_0209;
    126: op1_14_in25 = reg_0393;
    127: op1_14_in25 = reg_1383;
    128: op1_14_in25 = reg_0473;
    129: op1_14_in25 = reg_1203;
    130: op1_14_in25 = reg_0234;
    default: op1_14_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_14_inv25 = 1;
    55: op1_14_inv25 = 1;
    54: op1_14_inv25 = 1;
    69: op1_14_inv25 = 1;
    76: op1_14_inv25 = 1;
    71: op1_14_inv25 = 1;
    87: op1_14_inv25 = 1;
    57: op1_14_inv25 = 1;
    68: op1_14_inv25 = 1;
    77: op1_14_inv25 = 1;
    58: op1_14_inv25 = 1;
    70: op1_14_inv25 = 1;
    79: op1_14_inv25 = 1;
    51: op1_14_inv25 = 1;
    80: op1_14_inv25 = 1;
    81: op1_14_inv25 = 1;
    52: op1_14_inv25 = 1;
    64: op1_14_inv25 = 1;
    89: op1_14_inv25 = 1;
    85: op1_14_inv25 = 1;
    65: op1_14_inv25 = 1;
    90: op1_14_inv25 = 1;
    66: op1_14_inv25 = 1;
    48: op1_14_inv25 = 1;
    91: op1_14_inv25 = 1;
    67: op1_14_inv25 = 1;
    93: op1_14_inv25 = 1;
    94: op1_14_inv25 = 1;
    98: op1_14_inv25 = 1;
    99: op1_14_inv25 = 1;
    102: op1_14_inv25 = 1;
    104: op1_14_inv25 = 1;
    106: op1_14_inv25 = 1;
    110: op1_14_inv25 = 1;
    111: op1_14_inv25 = 1;
    112: op1_14_inv25 = 1;
    117: op1_14_inv25 = 1;
    123: op1_14_inv25 = 1;
    124: op1_14_inv25 = 1;
    127: op1_14_inv25 = 1;
    129: op1_14_inv25 = 1;
    default: op1_14_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in26 = reg_0785;
    53: op1_14_in26 = reg_0822;
    73: op1_14_in26 = reg_0967;
    55: op1_14_in26 = reg_0739;
    86: op1_14_in26 = reg_0199;
    74: op1_14_in26 = reg_1351;
    54: op1_14_in26 = reg_0529;
    75: op1_14_in26 = reg_0161;
    49: op1_14_in26 = reg_0738;
    69: op1_14_in26 = reg_0113;
    56: op1_14_in26 = reg_1169;
    76: op1_14_in26 = reg_1493;
    71: op1_14_in26 = reg_0610;
    87: op1_14_in26 = reg_0535;
    57: op1_14_in26 = reg_0779;
    68: op1_14_in26 = reg_0180;
    77: op1_14_in26 = reg_0151;
    61: op1_14_in26 = reg_0724;
    78: op1_14_in26 = reg_0797;
    58: op1_14_in26 = reg_0801;
    70: op1_14_in26 = reg_0396;
    59: op1_14_in26 = reg_0196;
    79: op1_14_in26 = reg_0620;
    51: op1_14_in26 = reg_0971;
    60: op1_14_in26 = reg_0064;
    124: op1_14_in26 = reg_0064;
    80: op1_14_in26 = reg_0623;
    88: op1_14_in26 = reg_0790;
    81: op1_14_in26 = reg_0922;
    82: op1_14_in26 = reg_0443;
    52: op1_14_in26 = reg_0137;
    64: op1_14_in26 = reg_0792;
    83: op1_14_in26 = reg_0875;
    112: op1_14_in26 = reg_0875;
    89: op1_14_in26 = reg_0604;
    84: op1_14_in26 = reg_0419;
    85: op1_14_in26 = reg_0238;
    65: op1_14_in26 = reg_0100;
    90: op1_14_in26 = reg_0488;
    66: op1_14_in26 = imem02_in[7:4];
    48: op1_14_in26 = reg_0132;
    91: op1_14_in26 = reg_0549;
    46: op1_14_in26 = reg_0220;
    67: op1_14_in26 = reg_0268;
    92: op1_14_in26 = reg_0084;
    93: op1_14_in26 = reg_0603;
    94: op1_14_in26 = imem02_in[3:0];
    97: op1_14_in26 = reg_0837;
    98: op1_14_in26 = reg_0507;
    99: op1_14_in26 = reg_0636;
    100: op1_14_in26 = reg_0552;
    101: op1_14_in26 = reg_0661;
    113: op1_14_in26 = reg_0661;
    102: op1_14_in26 = reg_0891;
    103: op1_14_in26 = reg_0566;
    104: op1_14_in26 = reg_0374;
    105: op1_14_in26 = reg_0593;
    106: op1_14_in26 = reg_0438;
    107: op1_14_in26 = reg_1145;
    109: op1_14_in26 = reg_0016;
    110: op1_14_in26 = reg_1457;
    111: op1_14_in26 = reg_0570;
    114: op1_14_in26 = reg_0479;
    115: op1_14_in26 = reg_0622;
    116: op1_14_in26 = reg_1425;
    117: op1_14_in26 = reg_0275;
    118: op1_14_in26 = reg_0165;
    47: op1_14_in26 = reg_0366;
    120: op1_14_in26 = reg_0146;
    121: op1_14_in26 = reg_0750;
    122: op1_14_in26 = reg_0726;
    126: op1_14_in26 = reg_0130;
    127: op1_14_in26 = reg_0328;
    128: op1_14_in26 = reg_1098;
    129: op1_14_in26 = reg_1215;
    130: op1_14_in26 = reg_0965;
    default: op1_14_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv26 = 1;
    53: op1_14_inv26 = 1;
    73: op1_14_inv26 = 1;
    74: op1_14_inv26 = 1;
    54: op1_14_inv26 = 1;
    69: op1_14_inv26 = 1;
    56: op1_14_inv26 = 1;
    76: op1_14_inv26 = 1;
    71: op1_14_inv26 = 1;
    87: op1_14_inv26 = 1;
    68: op1_14_inv26 = 1;
    77: op1_14_inv26 = 1;
    61: op1_14_inv26 = 1;
    78: op1_14_inv26 = 1;
    70: op1_14_inv26 = 1;
    59: op1_14_inv26 = 1;
    79: op1_14_inv26 = 1;
    60: op1_14_inv26 = 1;
    80: op1_14_inv26 = 1;
    81: op1_14_inv26 = 1;
    52: op1_14_inv26 = 1;
    83: op1_14_inv26 = 1;
    65: op1_14_inv26 = 1;
    90: op1_14_inv26 = 1;
    66: op1_14_inv26 = 1;
    48: op1_14_inv26 = 1;
    67: op1_14_inv26 = 1;
    94: op1_14_inv26 = 1;
    97: op1_14_inv26 = 1;
    100: op1_14_inv26 = 1;
    101: op1_14_inv26 = 1;
    103: op1_14_inv26 = 1;
    107: op1_14_inv26 = 1;
    110: op1_14_inv26 = 1;
    111: op1_14_inv26 = 1;
    113: op1_14_inv26 = 1;
    115: op1_14_inv26 = 1;
    116: op1_14_inv26 = 1;
    117: op1_14_inv26 = 1;
    118: op1_14_inv26 = 1;
    47: op1_14_inv26 = 1;
    121: op1_14_inv26 = 1;
    124: op1_14_inv26 = 1;
    126: op1_14_inv26 = 1;
    127: op1_14_inv26 = 1;
    128: op1_14_inv26 = 1;
    130: op1_14_inv26 = 1;
    default: op1_14_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in27 = reg_0372;
    53: op1_14_in27 = reg_0115;
    73: op1_14_in27 = reg_0439;
    55: op1_14_in27 = reg_0738;
    86: op1_14_in27 = reg_1004;
    74: op1_14_in27 = reg_0187;
    54: op1_14_in27 = reg_0132;
    75: op1_14_in27 = reg_0669;
    49: op1_14_in27 = reg_0103;
    69: op1_14_in27 = reg_0885;
    56: op1_14_in27 = reg_0347;
    76: op1_14_in27 = reg_0457;
    71: op1_14_in27 = reg_0420;
    87: op1_14_in27 = reg_0264;
    57: op1_14_in27 = reg_0029;
    68: op1_14_in27 = reg_0559;
    77: op1_14_in27 = reg_0861;
    61: op1_14_in27 = reg_0278;
    78: op1_14_in27 = reg_0449;
    58: op1_14_in27 = reg_0276;
    70: op1_14_in27 = reg_0464;
    59: op1_14_in27 = reg_0130;
    79: op1_14_in27 = reg_0114;
    51: op1_14_in27 = reg_0972;
    60: op1_14_in27 = reg_0063;
    80: op1_14_in27 = reg_0620;
    88: op1_14_in27 = reg_1383;
    81: op1_14_in27 = reg_0892;
    82: op1_14_in27 = reg_0488;
    52: op1_14_in27 = reg_0592;
    64: op1_14_in27 = reg_0578;
    83: op1_14_in27 = reg_0896;
    89: op1_14_in27 = reg_0986;
    109: op1_14_in27 = reg_0986;
    84: op1_14_in27 = reg_0270;
    85: op1_14_in27 = reg_0820;
    65: op1_14_in27 = reg_0228;
    90: op1_14_in27 = reg_0681;
    129: op1_14_in27 = reg_0681;
    66: op1_14_in27 = reg_0695;
    48: op1_14_in27 = reg_0171;
    91: op1_14_in27 = reg_0747;
    46: op1_14_in27 = reg_0557;
    67: op1_14_in27 = reg_0905;
    93: op1_14_in27 = reg_0268;
    94: op1_14_in27 = imem02_in[7:4];
    97: op1_14_in27 = reg_0096;
    98: op1_14_in27 = reg_0840;
    121: op1_14_in27 = reg_0840;
    99: op1_14_in27 = reg_0637;
    100: op1_14_in27 = reg_0281;
    101: op1_14_in27 = reg_0286;
    113: op1_14_in27 = reg_0286;
    102: op1_14_in27 = reg_0142;
    103: op1_14_in27 = reg_0564;
    104: op1_14_in27 = reg_0345;
    105: op1_14_in27 = reg_0483;
    106: op1_14_in27 = reg_0146;
    110: op1_14_in27 = reg_0146;
    107: op1_14_in27 = reg_0198;
    111: op1_14_in27 = reg_1225;
    112: op1_14_in27 = reg_0335;
    114: op1_14_in27 = imem03_in[3:0];
    115: op1_14_in27 = reg_0570;
    116: op1_14_in27 = reg_0216;
    117: op1_14_in27 = reg_0196;
    118: op1_14_in27 = reg_1204;
    47: op1_14_in27 = reg_0437;
    120: op1_14_in27 = reg_0362;
    122: op1_14_in27 = reg_0384;
    124: op1_14_in27 = reg_0020;
    126: op1_14_in27 = reg_0240;
    127: op1_14_in27 = reg_0797;
    128: op1_14_in27 = reg_0632;
    130: op1_14_in27 = reg_0964;
    default: op1_14_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv27 = 1;
    53: op1_14_inv27 = 1;
    55: op1_14_inv27 = 1;
    86: op1_14_inv27 = 1;
    74: op1_14_inv27 = 1;
    54: op1_14_inv27 = 1;
    75: op1_14_inv27 = 1;
    49: op1_14_inv27 = 1;
    69: op1_14_inv27 = 1;
    76: op1_14_inv27 = 1;
    57: op1_14_inv27 = 1;
    70: op1_14_inv27 = 1;
    59: op1_14_inv27 = 1;
    79: op1_14_inv27 = 1;
    60: op1_14_inv27 = 1;
    81: op1_14_inv27 = 1;
    89: op1_14_inv27 = 1;
    84: op1_14_inv27 = 1;
    66: op1_14_inv27 = 1;
    46: op1_14_inv27 = 1;
    67: op1_14_inv27 = 1;
    93: op1_14_inv27 = 1;
    97: op1_14_inv27 = 1;
    98: op1_14_inv27 = 1;
    99: op1_14_inv27 = 1;
    100: op1_14_inv27 = 1;
    102: op1_14_inv27 = 1;
    103: op1_14_inv27 = 1;
    109: op1_14_inv27 = 1;
    110: op1_14_inv27 = 1;
    111: op1_14_inv27 = 1;
    113: op1_14_inv27 = 1;
    114: op1_14_inv27 = 1;
    47: op1_14_inv27 = 1;
    121: op1_14_inv27 = 1;
    126: op1_14_inv27 = 1;
    129: op1_14_inv27 = 1;
    default: op1_14_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in28 = reg_1290;
    53: op1_14_in28 = reg_0670;
    73: op1_14_in28 = reg_0146;
    55: op1_14_in28 = reg_0404;
    86: op1_14_in28 = reg_0837;
    74: op1_14_in28 = reg_0225;
    54: op1_14_in28 = reg_0295;
    75: op1_14_in28 = reg_0716;
    49: op1_14_in28 = reg_0100;
    69: op1_14_in28 = reg_0880;
    56: op1_14_in28 = reg_0646;
    76: op1_14_in28 = reg_0590;
    71: op1_14_in28 = reg_0241;
    87: op1_14_in28 = reg_0252;
    82: op1_14_in28 = reg_0252;
    57: op1_14_in28 = reg_0663;
    68: op1_14_in28 = reg_1001;
    77: op1_14_in28 = reg_0751;
    61: op1_14_in28 = reg_0042;
    78: op1_14_in28 = reg_0828;
    58: op1_14_in28 = reg_0313;
    66: op1_14_in28 = reg_0313;
    70: op1_14_in28 = imem04_in[15:12];
    59: op1_14_in28 = reg_0243;
    79: op1_14_in28 = reg_0028;
    51: op1_14_in28 = reg_0111;
    60: op1_14_in28 = reg_0792;
    80: op1_14_in28 = reg_0592;
    88: op1_14_in28 = reg_0263;
    81: op1_14_in28 = reg_1350;
    52: op1_14_in28 = reg_0085;
    65: op1_14_in28 = reg_0085;
    64: op1_14_in28 = reg_0251;
    83: op1_14_in28 = reg_1139;
    89: op1_14_in28 = reg_0196;
    84: op1_14_in28 = reg_1170;
    85: op1_14_in28 = reg_1473;
    90: op1_14_in28 = reg_1233;
    48: op1_14_in28 = reg_0023;
    91: op1_14_in28 = reg_0238;
    46: op1_14_in28 = reg_0113;
    67: op1_14_in28 = reg_0960;
    93: op1_14_in28 = reg_0396;
    94: op1_14_in28 = reg_1235;
    97: op1_14_in28 = reg_0420;
    98: op1_14_in28 = reg_0889;
    99: op1_14_in28 = reg_0570;
    100: op1_14_in28 = reg_0414;
    101: op1_14_in28 = reg_0366;
    102: op1_14_in28 = reg_1516;
    130: op1_14_in28 = reg_1516;
    103: op1_14_in28 = reg_0131;
    104: op1_14_in28 = reg_0979;
    115: op1_14_in28 = reg_0979;
    106: op1_14_in28 = reg_0290;
    107: op1_14_in28 = reg_0145;
    109: op1_14_in28 = reg_0346;
    110: op1_14_in28 = reg_0292;
    111: op1_14_in28 = reg_0171;
    112: op1_14_in28 = reg_0728;
    113: op1_14_in28 = reg_0103;
    114: op1_14_in28 = reg_1145;
    116: op1_14_in28 = reg_0312;
    117: op1_14_in28 = reg_0393;
    118: op1_14_in28 = reg_0067;
    47: op1_14_in28 = reg_0415;
    120: op1_14_in28 = reg_0365;
    121: op1_14_in28 = reg_0573;
    122: op1_14_in28 = reg_0077;
    124: op1_14_in28 = imem05_in[7:4];
    126: op1_14_in28 = reg_0575;
    127: op1_14_in28 = reg_0297;
    128: op1_14_in28 = reg_0377;
    129: op1_14_in28 = reg_1077;
    default: op1_14_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    74: op1_14_inv28 = 1;
    49: op1_14_inv28 = 1;
    69: op1_14_inv28 = 1;
    76: op1_14_inv28 = 1;
    57: op1_14_inv28 = 1;
    68: op1_14_inv28 = 1;
    77: op1_14_inv28 = 1;
    61: op1_14_inv28 = 1;
    51: op1_14_inv28 = 1;
    82: op1_14_inv28 = 1;
    52: op1_14_inv28 = 1;
    83: op1_14_inv28 = 1;
    84: op1_14_inv28 = 1;
    85: op1_14_inv28 = 1;
    65: op1_14_inv28 = 1;
    91: op1_14_inv28 = 1;
    94: op1_14_inv28 = 1;
    98: op1_14_inv28 = 1;
    99: op1_14_inv28 = 1;
    103: op1_14_inv28 = 1;
    107: op1_14_inv28 = 1;
    112: op1_14_inv28 = 1;
    114: op1_14_inv28 = 1;
    116: op1_14_inv28 = 1;
    117: op1_14_inv28 = 1;
    118: op1_14_inv28 = 1;
    47: op1_14_inv28 = 1;
    120: op1_14_inv28 = 1;
    122: op1_14_inv28 = 1;
    124: op1_14_inv28 = 1;
    126: op1_14_inv28 = 1;
    127: op1_14_inv28 = 1;
    128: op1_14_inv28 = 1;
    129: op1_14_inv28 = 1;
    default: op1_14_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in29 = reg_0258;
    53: op1_14_in29 = reg_0636;
    73: op1_14_in29 = reg_0360;
    55: op1_14_in29 = reg_0592;
    86: op1_14_in29 = reg_0836;
    74: op1_14_in29 = reg_0297;
    54: op1_14_in29 = reg_0461;
    75: op1_14_in29 = reg_1302;
    49: op1_14_in29 = reg_0004;
    69: op1_14_in29 = reg_0884;
    56: op1_14_in29 = reg_0648;
    76: op1_14_in29 = reg_0256;
    71: op1_14_in29 = reg_0984;
    87: op1_14_in29 = reg_1198;
    57: op1_14_in29 = reg_0284;
    68: op1_14_in29 = reg_0597;
    77: op1_14_in29 = reg_0268;
    61: op1_14_in29 = reg_0457;
    78: op1_14_in29 = reg_0207;
    58: op1_14_in29 = reg_0756;
    70: op1_14_in29 = reg_0451;
    129: op1_14_in29 = reg_0451;
    59: op1_14_in29 = reg_0864;
    79: op1_14_in29 = reg_0050;
    80: op1_14_in29 = reg_0050;
    51: op1_14_in29 = reg_0897;
    60: op1_14_in29 = reg_0391;
    88: op1_14_in29 = reg_0181;
    81: op1_14_in29 = reg_1347;
    82: op1_14_in29 = reg_1338;
    52: op1_14_in29 = reg_0520;
    64: op1_14_in29 = reg_0702;
    83: op1_14_in29 = reg_1029;
    89: op1_14_in29 = reg_0130;
    84: op1_14_in29 = reg_0490;
    85: op1_14_in29 = reg_0966;
    90: op1_14_in29 = reg_0796;
    66: op1_14_in29 = reg_0198;
    48: op1_14_in29 = reg_0152;
    118: op1_14_in29 = reg_0152;
    91: op1_14_in29 = reg_0241;
    46: op1_14_in29 = reg_0425;
    67: op1_14_in29 = reg_0925;
    93: op1_14_in29 = reg_0931;
    94: op1_14_in29 = reg_0399;
    97: op1_14_in29 = reg_0020;
    98: op1_14_in29 = reg_0328;
    99: op1_14_in29 = reg_0979;
    100: op1_14_in29 = reg_0412;
    101: op1_14_in29 = reg_0738;
    102: op1_14_in29 = reg_0314;
    103: op1_14_in29 = reg_1070;
    104: op1_14_in29 = reg_0296;
    106: op1_14_in29 = reg_0899;
    107: op1_14_in29 = reg_0143;
    109: op1_14_in29 = reg_0700;
    110: op1_14_in29 = reg_0728;
    111: op1_14_in29 = reg_0215;
    112: op1_14_in29 = reg_0043;
    113: op1_14_in29 = reg_0114;
    47: op1_14_in29 = reg_0114;
    114: op1_14_in29 = reg_0573;
    115: op1_14_in29 = reg_1225;
    116: op1_14_in29 = reg_0375;
    117: op1_14_in29 = reg_0602;
    120: op1_14_in29 = reg_0400;
    121: op1_14_in29 = reg_0179;
    122: op1_14_in29 = reg_0257;
    124: op1_14_in29 = reg_0646;
    126: op1_14_in29 = reg_1346;
    127: op1_14_in29 = reg_0681;
    128: op1_14_in29 = reg_0220;
    130: op1_14_in29 = reg_1208;
    default: op1_14_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv29 = 1;
    53: op1_14_inv29 = 1;
    74: op1_14_inv29 = 1;
    75: op1_14_inv29 = 1;
    49: op1_14_inv29 = 1;
    76: op1_14_inv29 = 1;
    71: op1_14_inv29 = 1;
    57: op1_14_inv29 = 1;
    68: op1_14_inv29 = 1;
    60: op1_14_inv29 = 1;
    81: op1_14_inv29 = 1;
    52: op1_14_inv29 = 1;
    64: op1_14_inv29 = 1;
    83: op1_14_inv29 = 1;
    91: op1_14_inv29 = 1;
    67: op1_14_inv29 = 1;
    99: op1_14_inv29 = 1;
    100: op1_14_inv29 = 1;
    103: op1_14_inv29 = 1;
    104: op1_14_inv29 = 1;
    107: op1_14_inv29 = 1;
    109: op1_14_inv29 = 1;
    110: op1_14_inv29 = 1;
    112: op1_14_inv29 = 1;
    116: op1_14_inv29 = 1;
    117: op1_14_inv29 = 1;
    47: op1_14_inv29 = 1;
    122: op1_14_inv29 = 1;
    129: op1_14_inv29 = 1;
    130: op1_14_inv29 = 1;
    default: op1_14_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_14_in30 = reg_0239;
    53: op1_14_in30 = reg_0527;
    73: op1_14_in30 = reg_0899;
    55: op1_14_in30 = reg_0100;
    86: op1_14_in30 = reg_0719;
    74: op1_14_in30 = reg_1349;
    54: op1_14_in30 = imem06_in[3:0];
    75: op1_14_in30 = reg_0374;
    49: op1_14_in30 = reg_0001;
    69: op1_14_in30 = reg_0480;
    56: op1_14_in30 = imem05_in[11:8];
    76: op1_14_in30 = reg_0473;
    71: op1_14_in30 = reg_0967;
    85: op1_14_in30 = reg_0967;
    87: op1_14_in30 = reg_1200;
    57: op1_14_in30 = reg_0441;
    68: op1_14_in30 = imem03_in[7:4];
    77: op1_14_in30 = reg_0730;
    61: op1_14_in30 = imem02_in[11:8];
    78: op1_14_in30 = reg_0206;
    58: op1_14_in30 = reg_0573;
    70: op1_14_in30 = reg_0452;
    100: op1_14_in30 = reg_0452;
    59: op1_14_in30 = reg_0205;
    79: op1_14_in30 = reg_0051;
    51: op1_14_in30 = reg_0898;
    60: op1_14_in30 = reg_1269;
    80: op1_14_in30 = reg_0123;
    88: op1_14_in30 = reg_0535;
    81: op1_14_in30 = reg_0924;
    82: op1_14_in30 = reg_1257;
    64: op1_14_in30 = reg_1259;
    83: op1_14_in30 = reg_0399;
    89: op1_14_in30 = reg_0631;
    84: op1_14_in30 = reg_1440;
    90: op1_14_in30 = reg_1147;
    66: op1_14_in30 = reg_0710;
    48: op1_14_in30 = reg_0017;
    91: op1_14_in30 = reg_0798;
    46: op1_14_in30 = reg_0443;
    67: op1_14_in30 = reg_0752;
    93: op1_14_in30 = reg_0905;
    94: op1_14_in30 = reg_0845;
    97: op1_14_in30 = reg_0210;
    98: op1_14_in30 = reg_0235;
    99: op1_14_in30 = reg_0323;
    101: op1_14_in30 = reg_0408;
    102: op1_14_in30 = reg_0954;
    103: op1_14_in30 = reg_0302;
    104: op1_14_in30 = reg_1204;
    106: op1_14_in30 = reg_0901;
    107: op1_14_in30 = reg_0964;
    109: op1_14_in30 = reg_0649;
    110: op1_14_in30 = reg_0042;
    111: op1_14_in30 = reg_0214;
    112: op1_14_in30 = reg_0662;
    114: op1_14_in30 = reg_1033;
    115: op1_14_in30 = reg_0308;
    116: op1_14_in30 = reg_0556;
    117: op1_14_in30 = reg_0729;
    118: op1_14_in30 = reg_0215;
    47: op1_14_in30 = reg_0321;
    120: op1_14_in30 = reg_0403;
    121: op1_14_in30 = reg_0709;
    122: op1_14_in30 = reg_0162;
    124: op1_14_in30 = reg_0040;
    126: op1_14_in30 = reg_0151;
    127: op1_14_in30 = reg_0094;
    128: op1_14_in30 = reg_0600;
    129: op1_14_in30 = reg_0097;
    130: op1_14_in30 = reg_0108;
    default: op1_14_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_14_inv30 = 1;
    55: op1_14_inv30 = 1;
    74: op1_14_inv30 = 1;
    54: op1_14_inv30 = 1;
    49: op1_14_inv30 = 1;
    57: op1_14_inv30 = 1;
    68: op1_14_inv30 = 1;
    61: op1_14_inv30 = 1;
    78: op1_14_inv30 = 1;
    58: op1_14_inv30 = 1;
    79: op1_14_inv30 = 1;
    51: op1_14_inv30 = 1;
    80: op1_14_inv30 = 1;
    81: op1_14_inv30 = 1;
    83: op1_14_inv30 = 1;
    89: op1_14_inv30 = 1;
    85: op1_14_inv30 = 1;
    90: op1_14_inv30 = 1;
    66: op1_14_inv30 = 1;
    93: op1_14_inv30 = 1;
    94: op1_14_inv30 = 1;
    97: op1_14_inv30 = 1;
    98: op1_14_inv30 = 1;
    100: op1_14_inv30 = 1;
    101: op1_14_inv30 = 1;
    104: op1_14_inv30 = 1;
    106: op1_14_inv30 = 1;
    110: op1_14_inv30 = 1;
    111: op1_14_inv30 = 1;
    114: op1_14_inv30 = 1;
    116: op1_14_inv30 = 1;
    47: op1_14_inv30 = 1;
    120: op1_14_inv30 = 1;
    124: op1_14_inv30 = 1;
    126: op1_14_inv30 = 1;
    128: op1_14_inv30 = 1;
    130: op1_14_inv30 = 1;
    default: op1_14_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_14_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#14の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_14_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の0番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in00 = reg_0613;
    73: op1_15_in00 = reg_1259;
    53: op1_15_in00 = reg_0555;
    63: op1_15_in00 = reg_0555;
    84: op1_15_in00 = reg_0555;
    55: op1_15_in00 = reg_0571;
    86: op1_15_in00 = reg_1447;
    74: op1_15_in00 = imem00_in[11:8];
    54: op1_15_in00 = reg_0430;
    75: op1_15_in00 = reg_0318;
    90: op1_15_in00 = reg_0318;
    69: op1_15_in00 = reg_0278;
    56: op1_15_in00 = reg_0715;
    49: op1_15_in00 = reg_0527;
    76: op1_15_in00 = reg_1207;
    87: op1_15_in00 = reg_0541;
    57: op1_15_in00 = reg_0257;
    50: op1_15_in00 = reg_0871;
    68: op1_15_in00 = reg_0880;
    71: op1_15_in00 = reg_0554;
    79: op1_15_in00 = reg_0554;
    77: op1_15_in00 = imem06_in[7:4];
    78: op1_15_in00 = reg_0040;
    52: op1_15_in00 = reg_0040;
    61: op1_15_in00 = reg_0219;
    58: op1_15_in00 = reg_1258;
    70: op1_15_in00 = reg_0216;
    59: op1_15_in00 = reg_0147;
    51: op1_15_in00 = reg_0588;
    60: op1_15_in00 = reg_0023;
    88: op1_15_in00 = reg_0088;
    80: op1_15_in00 = reg_0797;
    62: op1_15_in00 = reg_0962;
    81: op1_15_in00 = reg_1475;
    82: op1_15_in00 = reg_0978;
    83: op1_15_in00 = reg_0253;
    64: op1_15_in00 = reg_0629;
    89: op1_15_in00 = reg_1093;
    102: op1_15_in00 = reg_1093;
    85: op1_15_in00 = reg_0462;
    65: op1_15_in00 = reg_0283;
    66: op1_15_in00 = reg_1350;
    91: op1_15_in00 = reg_0411;
    46: op1_15_in00 = reg_0792;
    48: op1_15_in00 = reg_0282;
    67: op1_15_in00 = reg_0580;
    92: op1_15_in00 = reg_0362;
    93: op1_15_in00 = reg_0397;
    94: op1_15_in00 = reg_0532;
    95: op1_15_in00 = reg_0983;
    96: op1_15_in00 = imem00_in[7:4];
    97: op1_15_in00 = imem05_in[11:8];
    98: op1_15_in00 = reg_0185;
    99: op1_15_in00 = reg_0244;
    100: op1_15_in00 = reg_0342;
    33: op1_15_in00 = imem07_in[7:4];
    101: op1_15_in00 = reg_0907;
    103: op1_15_in00 = reg_0090;
    104: op1_15_in00 = reg_1244;
    105: op1_15_in00 = imem00_in[15:12];
    119: op1_15_in00 = imem00_in[15:12];
    106: op1_15_in00 = reg_0175;
    107: op1_15_in00 = reg_0070;
    108: op1_15_in00 = reg_0866;
    109: op1_15_in00 = reg_0392;
    37: op1_15_in00 = reg_0225;
    28: op1_15_in00 = reg_0085;
    110: op1_15_in00 = imem02_in[7:4];
    111: op1_15_in00 = reg_0213;
    118: op1_15_in00 = reg_0213;
    112: op1_15_in00 = reg_0456;
    113: op1_15_in00 = imem00_in[3:0];
    114: op1_15_in00 = reg_0000;
    115: op1_15_in00 = reg_0119;
    116: op1_15_in00 = reg_1184;
    117: op1_15_in00 = reg_1035;
    47: op1_15_in00 = reg_0649;
    120: op1_15_in00 = reg_0166;
    121: op1_15_in00 = reg_1063;
    122: op1_15_in00 = reg_0634;
    123: op1_15_in00 = reg_0843;
    124: op1_15_in00 = reg_0445;
    125: op1_15_in00 = reg_1469;
    126: op1_15_in00 = reg_1030;
    127: op1_15_in00 = reg_0014;
    128: op1_15_in00 = reg_0311;
    129: op1_15_in00 = reg_0033;
    130: op1_15_in00 = reg_0559;
    default: op1_15_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の0番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv00 = 1;
    54: op1_15_inv00 = 1;
    75: op1_15_inv00 = 1;
    69: op1_15_inv00 = 1;
    49: op1_15_inv00 = 1;
    87: op1_15_inv00 = 1;
    57: op1_15_inv00 = 1;
    50: op1_15_inv00 = 1;
    71: op1_15_inv00 = 1;
    78: op1_15_inv00 = 1;
    61: op1_15_inv00 = 1;
    58: op1_15_inv00 = 1;
    70: op1_15_inv00 = 1;
    59: op1_15_inv00 = 1;
    88: op1_15_inv00 = 1;
    80: op1_15_inv00 = 1;
    62: op1_15_inv00 = 1;
    83: op1_15_inv00 = 1;
    64: op1_15_inv00 = 1;
    89: op1_15_inv00 = 1;
    90: op1_15_inv00 = 1;
    91: op1_15_inv00 = 1;
    46: op1_15_inv00 = 1;
    48: op1_15_inv00 = 1;
    94: op1_15_inv00 = 1;
    95: op1_15_inv00 = 1;
    99: op1_15_inv00 = 1;
    33: op1_15_inv00 = 1;
    101: op1_15_inv00 = 1;
    103: op1_15_inv00 = 1;
    106: op1_15_inv00 = 1;
    107: op1_15_inv00 = 1;
    108: op1_15_inv00 = 1;
    109: op1_15_inv00 = 1;
    28: op1_15_inv00 = 1;
    113: op1_15_inv00 = 1;
    114: op1_15_inv00 = 1;
    115: op1_15_inv00 = 1;
    117: op1_15_inv00 = 1;
    119: op1_15_inv00 = 1;
    121: op1_15_inv00 = 1;
    122: op1_15_inv00 = 1;
    125: op1_15_inv00 = 1;
    126: op1_15_inv00 = 1;
    127: op1_15_inv00 = 1;
    128: op1_15_inv00 = 1;
    129: op1_15_inv00 = 1;
    default: op1_15_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の1番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in01 = reg_0615;
    61: op1_15_in01 = reg_0615;
    73: op1_15_in01 = reg_0700;
    53: op1_15_in01 = reg_0580;
    71: op1_15_in01 = reg_0580;
    55: op1_15_in01 = reg_0528;
    86: op1_15_in01 = reg_0049;
    74: op1_15_in01 = reg_1277;
    54: op1_15_in01 = reg_0362;
    75: op1_15_in01 = reg_1485;
    69: op1_15_in01 = reg_0486;
    56: op1_15_in01 = reg_0438;
    49: op1_15_in01 = reg_0132;
    76: op1_15_in01 = reg_0973;
    87: op1_15_in01 = reg_0143;
    57: op1_15_in01 = reg_0238;
    50: op1_15_in01 = reg_0875;
    68: op1_15_in01 = imem03_in[7:4];
    77: op1_15_in01 = imem06_in[11:8];
    78: op1_15_in01 = reg_0014;
    58: op1_15_in01 = reg_0577;
    70: op1_15_in01 = reg_0378;
    59: op1_15_in01 = reg_0149;
    79: op1_15_in01 = imem00_in[3:0];
    125: op1_15_in01 = imem00_in[3:0];
    51: op1_15_in01 = reg_0561;
    60: op1_15_in01 = reg_1170;
    99: op1_15_in01 = reg_1170;
    88: op1_15_in01 = reg_0252;
    80: op1_15_in01 = reg_0861;
    62: op1_15_in01 = reg_0597;
    81: op1_15_in01 = reg_0572;
    82: op1_15_in01 = reg_1203;
    63: op1_15_in01 = reg_0613;
    52: op1_15_in01 = reg_0974;
    83: op1_15_in01 = reg_0456;
    64: op1_15_in01 = reg_0186;
    89: op1_15_in01 = reg_1208;
    84: op1_15_in01 = imem00_in[15:12];
    85: op1_15_in01 = reg_0796;
    65: op1_15_in01 = reg_0010;
    90: op1_15_in01 = reg_1484;
    66: op1_15_in01 = reg_0923;
    91: op1_15_in01 = reg_1372;
    46: op1_15_in01 = reg_0793;
    48: op1_15_in01 = reg_0044;
    67: op1_15_in01 = reg_0669;
    92: op1_15_in01 = reg_0363;
    93: op1_15_in01 = reg_0925;
    94: op1_15_in01 = reg_0970;
    95: op1_15_in01 = imem00_in[7:4];
    123: op1_15_in01 = imem00_in[7:4];
    96: op1_15_in01 = reg_0866;
    97: op1_15_in01 = reg_0750;
    98: op1_15_in01 = reg_0444;
    100: op1_15_in01 = reg_0835;
    33: op1_15_in01 = reg_0593;
    101: op1_15_in01 = reg_0555;
    102: op1_15_in01 = reg_1199;
    103: op1_15_in01 = reg_1373;
    104: op1_15_in01 = reg_0319;
    105: op1_15_in01 = reg_1101;
    106: op1_15_in01 = reg_0335;
    107: op1_15_in01 = reg_1517;
    108: op1_15_in01 = reg_0725;
    109: op1_15_in01 = reg_0045;
    37: op1_15_in01 = reg_0704;
    28: op1_15_in01 = reg_0050;
    110: op1_15_in01 = reg_0659;
    111: op1_15_in01 = reg_0084;
    112: op1_15_in01 = reg_0138;
    113: op1_15_in01 = reg_1242;
    114: op1_15_in01 = reg_0891;
    115: op1_15_in01 = reg_1202;
    116: op1_15_in01 = reg_0142;
    117: op1_15_in01 = reg_0870;
    118: op1_15_in01 = reg_0015;
    119: op1_15_in01 = reg_0581;
    47: op1_15_in01 = imem05_in[7:4];
    120: op1_15_in01 = reg_0447;
    121: op1_15_in01 = reg_0847;
    122: op1_15_in01 = reg_0889;
    124: op1_15_in01 = reg_0272;
    126: op1_15_in01 = reg_0825;
    127: op1_15_in01 = reg_0039;
    128: op1_15_in01 = reg_0191;
    129: op1_15_in01 = reg_0262;
    130: op1_15_in01 = reg_0790;
    default: op1_15_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の1番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv01 = 1;
    73: op1_15_inv01 = 1;
    53: op1_15_inv01 = 1;
    54: op1_15_inv01 = 1;
    56: op1_15_inv01 = 1;
    49: op1_15_inv01 = 1;
    76: op1_15_inv01 = 1;
    57: op1_15_inv01 = 1;
    50: op1_15_inv01 = 1;
    77: op1_15_inv01 = 1;
    78: op1_15_inv01 = 1;
    61: op1_15_inv01 = 1;
    58: op1_15_inv01 = 1;
    62: op1_15_inv01 = 1;
    81: op1_15_inv01 = 1;
    82: op1_15_inv01 = 1;
    52: op1_15_inv01 = 1;
    64: op1_15_inv01 = 1;
    84: op1_15_inv01 = 1;
    65: op1_15_inv01 = 1;
    90: op1_15_inv01 = 1;
    66: op1_15_inv01 = 1;
    48: op1_15_inv01 = 1;
    92: op1_15_inv01 = 1;
    94: op1_15_inv01 = 1;
    95: op1_15_inv01 = 1;
    97: op1_15_inv01 = 1;
    98: op1_15_inv01 = 1;
    99: op1_15_inv01 = 1;
    33: op1_15_inv01 = 1;
    103: op1_15_inv01 = 1;
    104: op1_15_inv01 = 1;
    105: op1_15_inv01 = 1;
    107: op1_15_inv01 = 1;
    109: op1_15_inv01 = 1;
    110: op1_15_inv01 = 1;
    111: op1_15_inv01 = 1;
    115: op1_15_inv01 = 1;
    117: op1_15_inv01 = 1;
    119: op1_15_inv01 = 1;
    121: op1_15_inv01 = 1;
    122: op1_15_inv01 = 1;
    123: op1_15_inv01 = 1;
    125: op1_15_inv01 = 1;
    126: op1_15_inv01 = 1;
    127: op1_15_inv01 = 1;
    128: op1_15_inv01 = 1;
    129: op1_15_inv01 = 1;
    130: op1_15_inv01 = 1;
    default: op1_15_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の2番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in02 = reg_1281;
    71: op1_15_in02 = reg_1281;
    63: op1_15_in02 = reg_1281;
    67: op1_15_in02 = reg_1281;
    96: op1_15_in02 = reg_1281;
    105: op1_15_in02 = reg_1281;
    73: op1_15_in02 = reg_0392;
    46: op1_15_in02 = reg_0392;
    53: op1_15_in02 = reg_1099;
    55: op1_15_in02 = reg_0527;
    86: op1_15_in02 = reg_0847;
    74: op1_15_in02 = reg_1079;
    95: op1_15_in02 = reg_1079;
    54: op1_15_in02 = reg_0047;
    75: op1_15_in02 = reg_0197;
    90: op1_15_in02 = reg_0197;
    69: op1_15_in02 = reg_0699;
    56: op1_15_in02 = reg_0727;
    49: op1_15_in02 = reg_0289;
    76: op1_15_in02 = reg_0972;
    87: op1_15_in02 = reg_0180;
    57: op1_15_in02 = reg_1152;
    50: op1_15_in02 = reg_0080;
    68: op1_15_in02 = imem03_in[11:8];
    77: op1_15_in02 = reg_0192;
    78: op1_15_in02 = reg_0780;
    61: op1_15_in02 = reg_1080;
    58: op1_15_in02 = reg_1214;
    70: op1_15_in02 = reg_1425;
    59: op1_15_in02 = reg_0402;
    79: op1_15_in02 = reg_0866;
    113: op1_15_in02 = reg_0866;
    51: op1_15_in02 = reg_0532;
    60: op1_15_in02 = reg_0491;
    88: op1_15_in02 = reg_0488;
    80: op1_15_in02 = reg_0317;
    62: op1_15_in02 = reg_0178;
    81: op1_15_in02 = reg_0967;
    82: op1_15_in02 = reg_0574;
    52: op1_15_in02 = reg_0751;
    83: op1_15_in02 = reg_0934;
    64: op1_15_in02 = reg_0667;
    89: op1_15_in02 = reg_0350;
    84: op1_15_in02 = reg_0791;
    85: op1_15_in02 = reg_0599;
    65: op1_15_in02 = reg_1029;
    66: op1_15_in02 = reg_0223;
    91: op1_15_in02 = reg_1368;
    48: op1_15_in02 = reg_0012;
    92: op1_15_in02 = reg_0092;
    93: op1_15_in02 = imem06_in[7:4];
    94: op1_15_in02 = reg_0127;
    97: op1_15_in02 = reg_0266;
    98: op1_15_in02 = reg_0706;
    99: op1_15_in02 = reg_1415;
    100: op1_15_in02 = reg_0932;
    33: op1_15_in02 = reg_0003;
    101: op1_15_in02 = reg_0961;
    102: op1_15_in02 = reg_0108;
    103: op1_15_in02 = reg_1346;
    104: op1_15_in02 = imem00_in[3:0];
    106: op1_15_in02 = reg_0078;
    107: op1_15_in02 = reg_0627;
    108: op1_15_in02 = reg_1489;
    109: op1_15_in02 = reg_0564;
    37: op1_15_in02 = reg_0309;
    28: op1_15_in02 = imem07_in[11:8];
    110: op1_15_in02 = reg_0626;
    111: op1_15_in02 = reg_0668;
    112: op1_15_in02 = reg_0561;
    114: op1_15_in02 = reg_0556;
    115: op1_15_in02 = reg_0977;
    116: op1_15_in02 = reg_1516;
    117: op1_15_in02 = reg_1504;
    118: op1_15_in02 = reg_0022;
    119: op1_15_in02 = reg_1470;
    47: op1_15_in02 = reg_0565;
    120: op1_15_in02 = reg_1071;
    121: op1_15_in02 = reg_0143;
    128: op1_15_in02 = reg_0143;
    122: op1_15_in02 = reg_0322;
    123: op1_15_in02 = reg_0725;
    124: op1_15_in02 = reg_0251;
    125: op1_15_in02 = reg_1141;
    126: op1_15_in02 = reg_0753;
    127: op1_15_in02 = reg_0729;
    129: op1_15_in02 = reg_0835;
    130: op1_15_in02 = reg_0348;
    default: op1_15_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の2番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv02 = 1;
    53: op1_15_inv02 = 1;
    86: op1_15_inv02 = 1;
    74: op1_15_inv02 = 1;
    54: op1_15_inv02 = 1;
    76: op1_15_inv02 = 1;
    87: op1_15_inv02 = 1;
    50: op1_15_inv02 = 1;
    68: op1_15_inv02 = 1;
    71: op1_15_inv02 = 1;
    61: op1_15_inv02 = 1;
    58: op1_15_inv02 = 1;
    60: op1_15_inv02 = 1;
    88: op1_15_inv02 = 1;
    81: op1_15_inv02 = 1;
    63: op1_15_inv02 = 1;
    52: op1_15_inv02 = 1;
    83: op1_15_inv02 = 1;
    89: op1_15_inv02 = 1;
    84: op1_15_inv02 = 1;
    66: op1_15_inv02 = 1;
    91: op1_15_inv02 = 1;
    48: op1_15_inv02 = 1;
    67: op1_15_inv02 = 1;
    93: op1_15_inv02 = 1;
    94: op1_15_inv02 = 1;
    95: op1_15_inv02 = 1;
    97: op1_15_inv02 = 1;
    98: op1_15_inv02 = 1;
    99: op1_15_inv02 = 1;
    100: op1_15_inv02 = 1;
    102: op1_15_inv02 = 1;
    103: op1_15_inv02 = 1;
    104: op1_15_inv02 = 1;
    105: op1_15_inv02 = 1;
    111: op1_15_inv02 = 1;
    112: op1_15_inv02 = 1;
    116: op1_15_inv02 = 1;
    118: op1_15_inv02 = 1;
    47: op1_15_inv02 = 1;
    120: op1_15_inv02 = 1;
    122: op1_15_inv02 = 1;
    123: op1_15_inv02 = 1;
    126: op1_15_inv02 = 1;
    127: op1_15_inv02 = 1;
    128: op1_15_inv02 = 1;
    129: op1_15_inv02 = 1;
    default: op1_15_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の3番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in03 = reg_1277;
    63: op1_15_in03 = reg_1277;
    73: op1_15_in03 = reg_0174;
    53: op1_15_in03 = reg_1081;
    55: op1_15_in03 = reg_0419;
    86: op1_15_in03 = reg_0789;
    74: op1_15_in03 = reg_1491;
    54: op1_15_in03 = reg_0078;
    75: op1_15_in03 = reg_0275;
    69: op1_15_in03 = reg_0532;
    56: op1_15_in03 = reg_0146;
    49: op1_15_in03 = reg_0119;
    76: op1_15_in03 = reg_0126;
    94: op1_15_in03 = reg_0126;
    87: op1_15_in03 = reg_0142;
    57: op1_15_in03 = reg_0715;
    50: op1_15_in03 = reg_0277;
    68: op1_15_in03 = reg_0790;
    71: op1_15_in03 = imem00_in[7:4];
    104: op1_15_in03 = imem00_in[7:4];
    77: op1_15_in03 = reg_0264;
    78: op1_15_in03 = reg_0795;
    61: op1_15_in03 = reg_1241;
    58: op1_15_in03 = reg_1216;
    70: op1_15_in03 = reg_0640;
    59: op1_15_in03 = reg_0384;
    79: op1_15_in03 = reg_1510;
    51: op1_15_in03 = reg_0475;
    60: op1_15_in03 = reg_1057;
    88: op1_15_in03 = reg_1147;
    80: op1_15_in03 = reg_0038;
    62: op1_15_in03 = reg_0505;
    81: op1_15_in03 = reg_0968;
    82: op1_15_in03 = reg_1083;
    52: op1_15_in03 = reg_0866;
    83: op1_15_in03 = reg_0055;
    64: op1_15_in03 = reg_0922;
    89: op1_15_in03 = reg_0313;
    84: op1_15_in03 = reg_0907;
    85: op1_15_in03 = reg_0305;
    65: op1_15_in03 = reg_0976;
    90: op1_15_in03 = reg_0130;
    66: op1_15_in03 = reg_1094;
    91: op1_15_in03 = reg_0088;
    46: op1_15_in03 = reg_0393;
    48: op1_15_in03 = reg_0553;
    67: op1_15_in03 = reg_0843;
    92: op1_15_in03 = reg_0175;
    93: op1_15_in03 = reg_0860;
    95: op1_15_in03 = reg_0804;
    96: op1_15_in03 = reg_1278;
    123: op1_15_in03 = reg_1278;
    97: op1_15_in03 = reg_0604;
    98: op1_15_in03 = reg_1033;
    99: op1_15_in03 = reg_1055;
    100: op1_15_in03 = reg_0536;
    33: op1_15_in03 = reg_0001;
    101: op1_15_in03 = reg_1432;
    102: op1_15_in03 = reg_0113;
    103: op1_15_in03 = reg_0799;
    105: op1_15_in03 = reg_0501;
    106: op1_15_in03 = reg_0079;
    107: op1_15_in03 = reg_0952;
    108: op1_15_in03 = reg_0293;
    109: op1_15_in03 = reg_0266;
    37: op1_15_in03 = reg_0298;
    110: op1_15_in03 = reg_0846;
    111: op1_15_in03 = reg_1096;
    112: op1_15_in03 = reg_0839;
    113: op1_15_in03 = reg_1099;
    114: op1_15_in03 = reg_1184;
    115: op1_15_in03 = reg_0067;
    116: op1_15_in03 = reg_1518;
    117: op1_15_in03 = reg_0265;
    118: op1_15_in03 = reg_0017;
    119: op1_15_in03 = reg_0638;
    47: op1_15_in03 = reg_0540;
    120: op1_15_in03 = reg_0662;
    121: op1_15_in03 = reg_0314;
    122: op1_15_in03 = reg_0845;
    124: op1_15_in03 = reg_0996;
    125: op1_15_in03 = reg_1490;
    126: op1_15_in03 = reg_1323;
    127: op1_15_in03 = reg_0397;
    128: op1_15_in03 = reg_1494;
    129: op1_15_in03 = reg_0096;
    130: op1_15_in03 = reg_0368;
    default: op1_15_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の3番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_15_inv03 = 1;
    53: op1_15_inv03 = 1;
    74: op1_15_inv03 = 1;
    54: op1_15_inv03 = 1;
    69: op1_15_inv03 = 1;
    87: op1_15_inv03 = 1;
    57: op1_15_inv03 = 1;
    77: op1_15_inv03 = 1;
    78: op1_15_inv03 = 1;
    70: op1_15_inv03 = 1;
    79: op1_15_inv03 = 1;
    82: op1_15_inv03 = 1;
    64: op1_15_inv03 = 1;
    85: op1_15_inv03 = 1;
    48: op1_15_inv03 = 1;
    67: op1_15_inv03 = 1;
    92: op1_15_inv03 = 1;
    93: op1_15_inv03 = 1;
    100: op1_15_inv03 = 1;
    33: op1_15_inv03 = 1;
    102: op1_15_inv03 = 1;
    104: op1_15_inv03 = 1;
    105: op1_15_inv03 = 1;
    37: op1_15_inv03 = 1;
    110: op1_15_inv03 = 1;
    111: op1_15_inv03 = 1;
    114: op1_15_inv03 = 1;
    117: op1_15_inv03 = 1;
    119: op1_15_inv03 = 1;
    47: op1_15_inv03 = 1;
    121: op1_15_inv03 = 1;
    122: op1_15_inv03 = 1;
    123: op1_15_inv03 = 1;
    125: op1_15_inv03 = 1;
    129: op1_15_inv03 = 1;
    130: op1_15_inv03 = 1;
    default: op1_15_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の4番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in04 = reg_1081;
    73: op1_15_in04 = reg_0646;
    53: op1_15_in04 = reg_0293;
    55: op1_15_in04 = reg_0289;
    86: op1_15_in04 = reg_0375;
    74: op1_15_in04 = reg_0562;
    54: op1_15_in04 = reg_0291;
    75: op1_15_in04 = reg_0240;
    69: op1_15_in04 = reg_0253;
    56: op1_15_in04 = reg_0383;
    49: op1_15_in04 = reg_0023;
    76: op1_15_in04 = reg_0112;
    87: op1_15_in04 = reg_0314;
    57: op1_15_in04 = reg_0968;
    50: op1_15_in04 = reg_0282;
    68: op1_15_in04 = reg_1280;
    71: op1_15_in04 = reg_1230;
    77: op1_15_in04 = reg_0827;
    78: op1_15_in04 = reg_1426;
    61: op1_15_in04 = reg_1028;
    58: op1_15_in04 = reg_1203;
    70: op1_15_in04 = reg_1325;
    59: op1_15_in04 = reg_0385;
    79: op1_15_in04 = reg_0868;
    51: op1_15_in04 = reg_0981;
    60: op1_15_in04 = reg_1055;
    88: op1_15_in04 = reg_0969;
    80: op1_15_in04 = reg_0014;
    62: op1_15_in04 = reg_0479;
    81: op1_15_in04 = reg_0149;
    82: op1_15_in04 = reg_0199;
    63: op1_15_in04 = reg_1080;
    52: op1_15_in04 = reg_0860;
    83: op1_15_in04 = reg_1074;
    64: op1_15_in04 = reg_0225;
    89: op1_15_in04 = reg_0341;
    84: op1_15_in04 = reg_0640;
    85: op1_15_in04 = reg_0319;
    65: op1_15_in04 = reg_0605;
    90: op1_15_in04 = reg_0861;
    66: op1_15_in04 = reg_0779;
    91: op1_15_in04 = reg_0264;
    46: op1_15_in04 = reg_0832;
    48: op1_15_in04 = reg_0255;
    67: op1_15_in04 = reg_1242;
    92: op1_15_in04 = reg_0080;
    93: op1_15_in04 = reg_0752;
    94: op1_15_in04 = reg_0111;
    95: op1_15_in04 = reg_0907;
    96: op1_15_in04 = reg_0153;
    97: op1_15_in04 = reg_0491;
    98: op1_15_in04 = reg_0783;
    99: op1_15_in04 = reg_0310;
    100: op1_15_in04 = reg_0063;
    33: op1_15_in04 = reg_0084;
    101: op1_15_in04 = reg_1418;
    102: op1_15_in04 = reg_0882;
    103: op1_15_in04 = reg_0603;
    104: op1_15_in04 = reg_0725;
    105: op1_15_in04 = reg_0580;
    125: op1_15_in04 = reg_0580;
    106: op1_15_in04 = reg_0896;
    107: op1_15_in04 = reg_0190;
    108: op1_15_in04 = reg_1201;
    109: op1_15_in04 = reg_0303;
    37: op1_15_in04 = reg_0299;
    110: op1_15_in04 = reg_0423;
    111: op1_15_in04 = reg_1416;
    112: op1_15_in04 = reg_0744;
    113: op1_15_in04 = reg_0803;
    114: op1_15_in04 = reg_0627;
    121: op1_15_in04 = reg_0627;
    115: op1_15_in04 = reg_0215;
    116: op1_15_in04 = reg_0954;
    117: op1_15_in04 = reg_1302;
    118: op1_15_in04 = reg_0246;
    119: op1_15_in04 = reg_0613;
    47: op1_15_in04 = reg_0418;
    120: op1_15_in04 = reg_0666;
    122: op1_15_in04 = reg_0666;
    123: op1_15_in04 = reg_1277;
    124: op1_15_in04 = reg_1104;
    126: op1_15_in04 = reg_0115;
    127: op1_15_in04 = reg_1334;
    128: op1_15_in04 = reg_0965;
    129: op1_15_in04 = reg_0117;
    130: op1_15_in04 = imem04_in[7:4];
    default: op1_15_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の4番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv04 = 1;
    55: op1_15_inv04 = 1;
    86: op1_15_inv04 = 1;
    69: op1_15_inv04 = 1;
    49: op1_15_inv04 = 1;
    50: op1_15_inv04 = 1;
    71: op1_15_inv04 = 1;
    77: op1_15_inv04 = 1;
    70: op1_15_inv04 = 1;
    51: op1_15_inv04 = 1;
    60: op1_15_inv04 = 1;
    88: op1_15_inv04 = 1;
    80: op1_15_inv04 = 1;
    62: op1_15_inv04 = 1;
    63: op1_15_inv04 = 1;
    52: op1_15_inv04 = 1;
    83: op1_15_inv04 = 1;
    64: op1_15_inv04 = 1;
    89: op1_15_inv04 = 1;
    90: op1_15_inv04 = 1;
    94: op1_15_inv04 = 1;
    96: op1_15_inv04 = 1;
    97: op1_15_inv04 = 1;
    98: op1_15_inv04 = 1;
    33: op1_15_inv04 = 1;
    102: op1_15_inv04 = 1;
    105: op1_15_inv04 = 1;
    108: op1_15_inv04 = 1;
    37: op1_15_inv04 = 1;
    112: op1_15_inv04 = 1;
    113: op1_15_inv04 = 1;
    114: op1_15_inv04 = 1;
    115: op1_15_inv04 = 1;
    116: op1_15_inv04 = 1;
    117: op1_15_inv04 = 1;
    118: op1_15_inv04 = 1;
    120: op1_15_inv04 = 1;
    123: op1_15_inv04 = 1;
    124: op1_15_inv04 = 1;
    125: op1_15_inv04 = 1;
    127: op1_15_inv04 = 1;
    129: op1_15_inv04 = 1;
    default: op1_15_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の5番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in05 = imem00_in[11:8];
    73: op1_15_in05 = reg_0648;
    53: op1_15_in05 = reg_0987;
    55: op1_15_in05 = imem06_in[11:8];
    90: op1_15_in05 = imem06_in[11:8];
    86: op1_15_in05 = reg_0142;
    74: op1_15_in05 = reg_1469;
    54: op1_15_in05 = reg_0277;
    75: op1_15_in05 = reg_0631;
    69: op1_15_in05 = reg_1018;
    56: op1_15_in05 = reg_0362;
    59: op1_15_in05 = reg_0362;
    49: op1_15_in05 = reg_0457;
    76: op1_15_in05 = imem02_in[15:12];
    87: op1_15_in05 = reg_1314;
    57: op1_15_in05 = reg_0430;
    50: op1_15_in05 = reg_0255;
    68: op1_15_in05 = reg_0348;
    71: op1_15_in05 = reg_1432;
    77: op1_15_in05 = reg_1065;
    78: op1_15_in05 = reg_1209;
    61: op1_15_in05 = reg_0459;
    58: op1_15_in05 = reg_1077;
    70: op1_15_in05 = reg_0891;
    79: op1_15_in05 = reg_1079;
    51: op1_15_in05 = reg_0970;
    60: op1_15_in05 = reg_1183;
    88: op1_15_in05 = reg_0097;
    80: op1_15_in05 = reg_1105;
    62: op1_15_in05 = reg_0247;
    81: op1_15_in05 = reg_0401;
    82: op1_15_in05 = reg_0320;
    63: op1_15_in05 = reg_1243;
    52: op1_15_in05 = reg_0822;
    83: op1_15_in05 = reg_0436;
    64: op1_15_in05 = reg_1347;
    89: op1_15_in05 = reg_0032;
    84: op1_15_in05 = reg_1487;
    85: op1_15_in05 = reg_0262;
    65: op1_15_in05 = reg_0254;
    66: op1_15_in05 = reg_0284;
    91: op1_15_in05 = reg_0978;
    46: op1_15_in05 = reg_0523;
    48: op1_15_in05 = reg_0606;
    67: op1_15_in05 = reg_0805;
    113: op1_15_in05 = reg_0805;
    92: op1_15_in05 = reg_0734;
    93: op1_15_in05 = reg_1501;
    94: op1_15_in05 = reg_0628;
    95: op1_15_in05 = reg_0554;
    125: op1_15_in05 = reg_0554;
    96: op1_15_in05 = reg_0186;
    97: op1_15_in05 = reg_0045;
    98: op1_15_in05 = reg_0312;
    99: op1_15_in05 = reg_0139;
    100: op1_15_in05 = reg_0210;
    33: op1_15_in05 = reg_0519;
    101: op1_15_in05 = reg_0928;
    102: op1_15_in05 = reg_0884;
    103: op1_15_in05 = reg_0037;
    104: op1_15_in05 = reg_1281;
    105: op1_15_in05 = reg_0153;
    106: op1_15_in05 = reg_0162;
    107: op1_15_in05 = reg_1199;
    108: op1_15_in05 = reg_0961;
    109: op1_15_in05 = reg_0300;
    37: op1_15_in05 = reg_0674;
    110: op1_15_in05 = reg_0138;
    111: op1_15_in05 = reg_0478;
    112: op1_15_in05 = reg_0429;
    114: op1_15_in05 = reg_0957;
    115: op1_15_in05 = reg_0213;
    116: op1_15_in05 = reg_1300;
    117: op1_15_in05 = reg_0194;
    118: op1_15_in05 = reg_0995;
    119: op1_15_in05 = reg_0486;
    47: op1_15_in05 = reg_0895;
    120: op1_15_in05 = reg_0455;
    121: op1_15_in05 = reg_0541;
    122: op1_15_in05 = reg_0056;
    123: op1_15_in05 = reg_0803;
    124: op1_15_in05 = reg_1402;
    126: op1_15_in05 = reg_0622;
    127: op1_15_in05 = reg_0925;
    128: op1_15_in05 = reg_1517;
    129: op1_15_in05 = reg_0095;
    130: op1_15_in05 = imem04_in[11:8];
    default: op1_15_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の5番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv05 = 1;
    73: op1_15_inv05 = 1;
    55: op1_15_inv05 = 1;
    74: op1_15_inv05 = 1;
    75: op1_15_inv05 = 1;
    49: op1_15_inv05 = 1;
    76: op1_15_inv05 = 1;
    87: op1_15_inv05 = 1;
    57: op1_15_inv05 = 1;
    68: op1_15_inv05 = 1;
    77: op1_15_inv05 = 1;
    61: op1_15_inv05 = 1;
    58: op1_15_inv05 = 1;
    70: op1_15_inv05 = 1;
    51: op1_15_inv05 = 1;
    81: op1_15_inv05 = 1;
    84: op1_15_inv05 = 1;
    66: op1_15_inv05 = 1;
    46: op1_15_inv05 = 1;
    92: op1_15_inv05 = 1;
    93: op1_15_inv05 = 1;
    94: op1_15_inv05 = 1;
    95: op1_15_inv05 = 1;
    97: op1_15_inv05 = 1;
    33: op1_15_inv05 = 1;
    101: op1_15_inv05 = 1;
    102: op1_15_inv05 = 1;
    104: op1_15_inv05 = 1;
    106: op1_15_inv05 = 1;
    107: op1_15_inv05 = 1;
    37: op1_15_inv05 = 1;
    110: op1_15_inv05 = 1;
    111: op1_15_inv05 = 1;
    113: op1_15_inv05 = 1;
    114: op1_15_inv05 = 1;
    115: op1_15_inv05 = 1;
    117: op1_15_inv05 = 1;
    118: op1_15_inv05 = 1;
    47: op1_15_inv05 = 1;
    120: op1_15_inv05 = 1;
    121: op1_15_inv05 = 1;
    123: op1_15_inv05 = 1;
    124: op1_15_inv05 = 1;
    125: op1_15_inv05 = 1;
    126: op1_15_inv05 = 1;
    127: op1_15_inv05 = 1;
    129: op1_15_inv05 = 1;
    130: op1_15_inv05 = 1;
    default: op1_15_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の6番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in06 = reg_1469;
    73: op1_15_in06 = reg_0567;
    53: op1_15_in06 = imem00_in[7:4];
    55: op1_15_in06 = reg_0271;
    86: op1_15_in06 = reg_0952;
    74: op1_15_in06 = reg_0218;
    54: op1_15_in06 = reg_0041;
    75: op1_15_in06 = reg_0799;
    69: op1_15_in06 = reg_0589;
    56: op1_15_in06 = reg_0363;
    49: op1_15_in06 = reg_0490;
    76: op1_15_in06 = reg_0381;
    87: op1_15_in06 = reg_0178;
    107: op1_15_in06 = reg_0178;
    57: op1_15_in06 = reg_0384;
    81: op1_15_in06 = reg_0384;
    50: op1_15_in06 = imem02_in[3:0];
    68: op1_15_in06 = reg_0411;
    71: op1_15_in06 = reg_0476;
    77: op1_15_in06 = reg_0110;
    78: op1_15_in06 = reg_1334;
    61: op1_15_in06 = reg_0961;
    58: op1_15_in06 = reg_0797;
    70: op1_15_in06 = reg_0261;
    59: op1_15_in06 = reg_0360;
    79: op1_15_in06 = reg_1080;
    51: op1_15_in06 = reg_0973;
    60: op1_15_in06 = reg_0170;
    88: op1_15_in06 = reg_0319;
    80: op1_15_in06 = reg_0195;
    62: op1_15_in06 = reg_0694;
    82: op1_15_in06 = reg_0862;
    85: op1_15_in06 = reg_0862;
    63: op1_15_in06 = reg_1242;
    52: op1_15_in06 = reg_0718;
    83: op1_15_in06 = reg_0326;
    64: op1_15_in06 = reg_0159;
    89: op1_15_in06 = reg_0264;
    84: op1_15_in06 = reg_1491;
    65: op1_15_in06 = reg_0497;
    90: op1_15_in06 = reg_1508;
    66: op1_15_in06 = reg_0620;
    91: op1_15_in06 = reg_0552;
    46: op1_15_in06 = reg_0648;
    48: op1_15_in06 = reg_0605;
    67: op1_15_in06 = reg_0221;
    92: op1_15_in06 = reg_0044;
    93: op1_15_in06 = reg_0115;
    94: op1_15_in06 = reg_1492;
    95: op1_15_in06 = reg_0523;
    96: op1_15_in06 = reg_1053;
    97: op1_15_in06 = reg_0697;
    98: op1_15_in06 = reg_0143;
    99: op1_15_in06 = reg_0030;
    100: op1_15_in06 = imem05_in[11:8];
    101: op1_15_in06 = reg_0431;
    102: op1_15_in06 = imem04_in[11:8];
    103: op1_15_in06 = reg_0014;
    104: op1_15_in06 = reg_0748;
    105: op1_15_in06 = reg_1459;
    106: op1_15_in06 = reg_0402;
    108: op1_15_in06 = reg_0459;
    109: op1_15_in06 = reg_0872;
    37: op1_15_in06 = reg_0156;
    110: op1_15_in06 = reg_0133;
    111: op1_15_in06 = reg_0667;
    112: op1_15_in06 = reg_0436;
    113: op1_15_in06 = reg_0554;
    114: op1_15_in06 = reg_0048;
    115: op1_15_in06 = reg_1170;
    116: op1_15_in06 = reg_1301;
    117: op1_15_in06 = reg_0141;
    118: op1_15_in06 = reg_1095;
    119: op1_15_in06 = reg_0186;
    47: op1_15_in06 = reg_0302;
    120: op1_15_in06 = reg_1493;
    121: op1_15_in06 = reg_1009;
    122: op1_15_in06 = reg_0276;
    123: op1_15_in06 = reg_0555;
    124: op1_15_in06 = reg_1404;
    125: op1_15_in06 = reg_1417;
    126: op1_15_in06 = reg_0528;
    127: op1_15_in06 = reg_0870;
    128: op1_15_in06 = reg_0349;
    129: op1_15_in06 = reg_0210;
    130: op1_15_in06 = reg_1367;
    default: op1_15_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の6番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv06 = 1;
    53: op1_15_inv06 = 1;
    86: op1_15_inv06 = 1;
    69: op1_15_inv06 = 1;
    56: op1_15_inv06 = 1;
    76: op1_15_inv06 = 1;
    87: op1_15_inv06 = 1;
    57: op1_15_inv06 = 1;
    50: op1_15_inv06 = 1;
    68: op1_15_inv06 = 1;
    71: op1_15_inv06 = 1;
    79: op1_15_inv06 = 1;
    51: op1_15_inv06 = 1;
    80: op1_15_inv06 = 1;
    81: op1_15_inv06 = 1;
    83: op1_15_inv06 = 1;
    89: op1_15_inv06 = 1;
    90: op1_15_inv06 = 1;
    66: op1_15_inv06 = 1;
    91: op1_15_inv06 = 1;
    46: op1_15_inv06 = 1;
    48: op1_15_inv06 = 1;
    67: op1_15_inv06 = 1;
    93: op1_15_inv06 = 1;
    95: op1_15_inv06 = 1;
    100: op1_15_inv06 = 1;
    103: op1_15_inv06 = 1;
    104: op1_15_inv06 = 1;
    105: op1_15_inv06 = 1;
    106: op1_15_inv06 = 1;
    108: op1_15_inv06 = 1;
    37: op1_15_inv06 = 1;
    111: op1_15_inv06 = 1;
    112: op1_15_inv06 = 1;
    113: op1_15_inv06 = 1;
    114: op1_15_inv06 = 1;
    117: op1_15_inv06 = 1;
    118: op1_15_inv06 = 1;
    120: op1_15_inv06 = 1;
    121: op1_15_inv06 = 1;
    124: op1_15_inv06 = 1;
    125: op1_15_inv06 = 1;
    128: op1_15_inv06 = 1;
    129: op1_15_inv06 = 1;
    default: op1_15_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の7番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in07 = reg_1470;
    73: op1_15_in07 = reg_0564;
    53: op1_15_in07 = reg_0928;
    108: op1_15_in07 = reg_0928;
    55: op1_15_in07 = reg_0067;
    86: op1_15_in07 = reg_0246;
    74: op1_15_in07 = reg_1027;
    54: op1_15_in07 = reg_0486;
    75: op1_15_in07 = reg_0037;
    69: op1_15_in07 = reg_0934;
    56: op1_15_in07 = reg_0093;
    49: op1_15_in07 = reg_0226;
    76: op1_15_in07 = reg_0307;
    87: op1_15_in07 = reg_0107;
    57: op1_15_in07 = reg_0385;
    50: op1_15_in07 = reg_0975;
    68: op1_15_in07 = reg_0534;
    71: op1_15_in07 = reg_0886;
    77: op1_15_in07 = reg_1302;
    78: op1_15_in07 = reg_0669;
    61: op1_15_in07 = reg_0959;
    58: op1_15_in07 = reg_0340;
    70: op1_15_in07 = reg_1000;
    59: op1_15_in07 = reg_0724;
    79: op1_15_in07 = reg_1078;
    51: op1_15_in07 = reg_0972;
    60: op1_15_in07 = reg_0297;
    88: op1_15_in07 = reg_0862;
    80: op1_15_in07 = reg_1468;
    62: op1_15_in07 = reg_0536;
    81: op1_15_in07 = reg_0363;
    82: op1_15_in07 = reg_0470;
    129: op1_15_in07 = reg_0470;
    63: op1_15_in07 = reg_1053;
    52: op1_15_in07 = reg_0635;
    83: op1_15_in07 = reg_0973;
    64: op1_15_in07 = reg_0923;
    89: op1_15_in07 = reg_1233;
    84: op1_15_in07 = reg_0841;
    85: op1_15_in07 = reg_1237;
    65: op1_15_in07 = reg_0256;
    90: op1_15_in07 = reg_0984;
    66: op1_15_in07 = reg_0591;
    91: op1_15_in07 = reg_1215;
    46: op1_15_in07 = reg_0601;
    48: op1_15_in07 = imem02_in[11:8];
    67: op1_15_in07 = reg_0961;
    92: op1_15_in07 = reg_0662;
    93: op1_15_in07 = reg_0109;
    94: op1_15_in07 = reg_1392;
    95: op1_15_in07 = reg_1454;
    96: op1_15_in07 = reg_0250;
    113: op1_15_in07 = reg_0250;
    97: op1_15_in07 = reg_1401;
    98: op1_15_in07 = reg_0144;
    99: op1_15_in07 = reg_0665;
    100: op1_15_in07 = reg_0793;
    101: op1_15_in07 = reg_0440;
    102: op1_15_in07 = imem04_in[15:12];
    103: op1_15_in07 = imem06_in[15:12];
    104: op1_15_in07 = reg_1490;
    105: op1_15_in07 = reg_0229;
    106: op1_15_in07 = reg_0044;
    107: op1_15_in07 = reg_0104;
    109: op1_15_in07 = reg_0736;
    37: op1_15_in07 = reg_0140;
    110: op1_15_in07 = reg_0898;
    111: op1_15_in07 = reg_0786;
    112: op1_15_in07 = reg_0776;
    114: op1_15_in07 = reg_1093;
    115: op1_15_in07 = reg_0995;
    116: op1_15_in07 = reg_1226;
    117: op1_15_in07 = reg_0569;
    126: op1_15_in07 = reg_0569;
    118: op1_15_in07 = reg_1055;
    119: op1_15_in07 = reg_0555;
    47: op1_15_in07 = reg_0090;
    120: op1_15_in07 = reg_0532;
    121: op1_15_in07 = reg_1368;
    122: op1_15_in07 = reg_0608;
    123: op1_15_in07 = reg_0640;
    124: op1_15_in07 = reg_1070;
    125: op1_15_in07 = reg_1393;
    127: op1_15_in07 = reg_0271;
    128: op1_15_in07 = reg_0885;
    130: op1_15_in07 = reg_0236;
    default: op1_15_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の7番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_15_inv07 = 1;
    74: op1_15_inv07 = 1;
    69: op1_15_inv07 = 1;
    56: op1_15_inv07 = 1;
    49: op1_15_inv07 = 1;
    87: op1_15_inv07 = 1;
    57: op1_15_inv07 = 1;
    50: op1_15_inv07 = 1;
    68: op1_15_inv07 = 1;
    80: op1_15_inv07 = 1;
    82: op1_15_inv07 = 1;
    64: op1_15_inv07 = 1;
    89: op1_15_inv07 = 1;
    84: op1_15_inv07 = 1;
    85: op1_15_inv07 = 1;
    66: op1_15_inv07 = 1;
    91: op1_15_inv07 = 1;
    48: op1_15_inv07 = 1;
    92: op1_15_inv07 = 1;
    95: op1_15_inv07 = 1;
    96: op1_15_inv07 = 1;
    98: op1_15_inv07 = 1;
    102: op1_15_inv07 = 1;
    105: op1_15_inv07 = 1;
    108: op1_15_inv07 = 1;
    109: op1_15_inv07 = 1;
    37: op1_15_inv07 = 1;
    117: op1_15_inv07 = 1;
    118: op1_15_inv07 = 1;
    119: op1_15_inv07 = 1;
    47: op1_15_inv07 = 1;
    120: op1_15_inv07 = 1;
    121: op1_15_inv07 = 1;
    125: op1_15_inv07 = 1;
    126: op1_15_inv07 = 1;
    130: op1_15_inv07 = 1;
    default: op1_15_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の8番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in08 = reg_1053;
    73: op1_15_in08 = reg_0334;
    53: op1_15_in08 = reg_0926;
    55: op1_15_in08 = reg_0215;
    86: op1_15_in08 = reg_1301;
    74: op1_15_in08 = reg_1453;
    95: op1_15_in08 = reg_1453;
    54: op1_15_in08 = reg_0662;
    75: op1_15_in08 = reg_0039;
    69: op1_15_in08 = reg_0056;
    56: op1_15_in08 = reg_0724;
    49: op1_15_in08 = reg_0893;
    76: op1_15_in08 = reg_0294;
    87: op1_15_in08 = imem03_in[7:4];
    57: op1_15_in08 = reg_0093;
    50: op1_15_in08 = reg_0563;
    68: op1_15_in08 = reg_1203;
    71: op1_15_in08 = reg_0073;
    77: op1_15_in08 = reg_0637;
    93: op1_15_in08 = reg_0637;
    78: op1_15_in08 = reg_0718;
    61: op1_15_in08 = reg_0135;
    58: op1_15_in08 = reg_0837;
    70: op1_15_in08 = reg_1001;
    59: op1_15_in08 = reg_0278;
    79: op1_15_in08 = reg_1491;
    51: op1_15_in08 = reg_0934;
    60: op1_15_in08 = reg_0159;
    88: op1_15_in08 = reg_0835;
    80: op1_15_in08 = reg_1467;
    90: op1_15_in08 = reg_1467;
    62: op1_15_in08 = reg_0493;
    130: op1_15_in08 = reg_0493;
    81: op1_15_in08 = reg_0896;
    82: op1_15_in08 = reg_0204;
    63: op1_15_in08 = reg_0136;
    52: op1_15_in08 = reg_0264;
    83: op1_15_in08 = reg_1455;
    64: op1_15_in08 = reg_0284;
    89: op1_15_in08 = reg_0421;
    84: op1_15_in08 = reg_0615;
    85: op1_15_in08 = reg_0211;
    65: op1_15_in08 = reg_0472;
    110: op1_15_in08 = reg_0472;
    66: op1_15_in08 = reg_0137;
    91: op1_15_in08 = reg_0681;
    46: op1_15_in08 = reg_0604;
    48: op1_15_in08 = imem02_in[15:12];
    67: op1_15_in08 = imem00_in[11:8];
    92: op1_15_in08 = reg_0879;
    94: op1_15_in08 = reg_1091;
    96: op1_15_in08 = reg_0221;
    97: op1_15_in08 = reg_0418;
    98: op1_15_in08 = reg_1495;
    99: op1_15_in08 = reg_0663;
    100: op1_15_in08 = reg_0832;
    101: op1_15_in08 = reg_0409;
    102: op1_15_in08 = reg_1146;
    103: op1_15_in08 = reg_0784;
    104: op1_15_in08 = reg_0186;
    105: op1_15_in08 = reg_1417;
    106: op1_15_in08 = imem01_in[3:0];
    107: op1_15_in08 = reg_0880;
    108: op1_15_in08 = reg_0202;
    109: op1_15_in08 = reg_0274;
    37: op1_15_in08 = reg_0286;
    111: op1_15_in08 = reg_1349;
    112: op1_15_in08 = reg_0307;
    113: op1_15_in08 = reg_1459;
    114: op1_15_in08 = reg_0178;
    116: op1_15_in08 = reg_0178;
    115: op1_15_in08 = imem07_in[3:0];
    117: op1_15_in08 = reg_0570;
    118: op1_15_in08 = reg_1060;
    119: op1_15_in08 = reg_0523;
    47: op1_15_in08 = reg_0873;
    120: op1_15_in08 = reg_0105;
    121: op1_15_in08 = reg_0088;
    122: op1_15_in08 = reg_0561;
    123: op1_15_in08 = reg_1052;
    124: op1_15_in08 = reg_0938;
    125: op1_15_in08 = reg_0416;
    126: op1_15_in08 = reg_0345;
    127: op1_15_in08 = reg_0869;
    128: op1_15_in08 = reg_0882;
    129: op1_15_in08 = imem05_in[7:4];
    default: op1_15_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の8番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_15_inv08 = 1;
    55: op1_15_inv08 = 1;
    86: op1_15_inv08 = 1;
    74: op1_15_inv08 = 1;
    75: op1_15_inv08 = 1;
    69: op1_15_inv08 = 1;
    87: op1_15_inv08 = 1;
    50: op1_15_inv08 = 1;
    71: op1_15_inv08 = 1;
    59: op1_15_inv08 = 1;
    60: op1_15_inv08 = 1;
    88: op1_15_inv08 = 1;
    63: op1_15_inv08 = 1;
    52: op1_15_inv08 = 1;
    64: op1_15_inv08 = 1;
    89: op1_15_inv08 = 1;
    66: op1_15_inv08 = 1;
    91: op1_15_inv08 = 1;
    48: op1_15_inv08 = 1;
    93: op1_15_inv08 = 1;
    102: op1_15_inv08 = 1;
    108: op1_15_inv08 = 1;
    109: op1_15_inv08 = 1;
    110: op1_15_inv08 = 1;
    113: op1_15_inv08 = 1;
    115: op1_15_inv08 = 1;
    116: op1_15_inv08 = 1;
    117: op1_15_inv08 = 1;
    47: op1_15_inv08 = 1;
    123: op1_15_inv08 = 1;
    124: op1_15_inv08 = 1;
    125: op1_15_inv08 = 1;
    127: op1_15_inv08 = 1;
    128: op1_15_inv08 = 1;
    129: op1_15_inv08 = 1;
    130: op1_15_inv08 = 1;
    default: op1_15_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の9番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in09 = reg_0523;
    123: op1_15_in09 = reg_0523;
    73: op1_15_in09 = reg_1403;
    53: op1_15_in09 = reg_0887;
    55: op1_15_in09 = reg_0490;
    86: op1_15_in09 = reg_0558;
    74: op1_15_in09 = reg_1206;
    54: op1_15_in09 = imem02_in[7:4];
    75: op1_15_in09 = reg_0193;
    69: op1_15_in09 = reg_0381;
    56: op1_15_in09 = reg_0901;
    49: op1_15_in09 = reg_0867;
    76: op1_15_in09 = reg_0845;
    87: op1_15_in09 = reg_0291;
    57: op1_15_in09 = reg_0899;
    50: op1_15_in09 = reg_0472;
    68: op1_15_in09 = reg_1198;
    71: op1_15_in09 = reg_0075;
    77: op1_15_in09 = reg_0374;
    78: op1_15_in09 = reg_1303;
    61: op1_15_in09 = reg_0926;
    58: op1_15_in09 = reg_0337;
    70: op1_15_in09 = reg_1300;
    59: op1_15_in09 = reg_0254;
    122: op1_15_in09 = reg_0254;
    79: op1_15_in09 = reg_1242;
    51: op1_15_in09 = reg_0933;
    60: op1_15_in09 = reg_0156;
    88: op1_15_in09 = reg_0338;
    80: op1_15_in09 = reg_1064;
    62: op1_15_in09 = reg_0574;
    81: op1_15_in09 = reg_0290;
    82: op1_15_in09 = reg_0702;
    63: op1_15_in09 = reg_0249;
    95: op1_15_in09 = reg_0249;
    52: op1_15_in09 = reg_0568;
    83: op1_15_in09 = reg_0128;
    64: op1_15_in09 = reg_0441;
    89: op1_15_in09 = reg_0599;
    84: op1_15_in09 = reg_0806;
    85: op1_15_in09 = reg_0117;
    65: op1_15_in09 = reg_0970;
    90: op1_15_in09 = reg_0869;
    66: op1_15_in09 = reg_0100;
    91: op1_15_in09 = reg_0421;
    46: op1_15_in09 = reg_0566;
    48: op1_15_in09 = reg_0588;
    67: op1_15_in09 = reg_0476;
    92: op1_15_in09 = imem02_in[3:0];
    93: op1_15_in09 = reg_0398;
    94: op1_15_in09 = reg_0279;
    96: op1_15_in09 = reg_0485;
    97: op1_15_in09 = reg_0302;
    98: op1_15_in09 = reg_0965;
    99: op1_15_in09 = reg_0415;
    100: op1_15_in09 = reg_0347;
    101: op1_15_in09 = reg_0073;
    102: op1_15_in09 = reg_0181;
    103: op1_15_in09 = reg_1030;
    104: op1_15_in09 = reg_1028;
    105: op1_15_in09 = reg_1418;
    106: op1_15_in09 = reg_0662;
    107: op1_15_in09 = reg_1009;
    108: op1_15_in09 = reg_0352;
    109: op1_15_in09 = reg_0196;
    37: op1_15_in09 = imem07_in[7:4];
    110: op1_15_in09 = reg_0973;
    111: op1_15_in09 = reg_0923;
    112: op1_15_in09 = reg_0473;
    113: op1_15_in09 = reg_1406;
    114: op1_15_in09 = reg_0467;
    115: op1_15_in09 = reg_0394;
    116: op1_15_in09 = reg_0885;
    117: op1_15_in09 = reg_0295;
    118: op1_15_in09 = reg_0298;
    119: op1_15_in09 = reg_1454;
    47: op1_15_in09 = reg_0130;
    120: op1_15_in09 = reg_0382;
    121: op1_15_in09 = reg_1258;
    124: op1_15_in09 = reg_0937;
    125: op1_15_in09 = reg_0072;
    126: op1_15_in09 = reg_0583;
    127: op1_15_in09 = reg_0827;
    128: op1_15_in09 = reg_0884;
    129: op1_15_in09 = reg_0708;
    130: op1_15_in09 = reg_0088;
    default: op1_15_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の9番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv09 = 1;
    73: op1_15_inv09 = 1;
    53: op1_15_inv09 = 1;
    86: op1_15_inv09 = 1;
    74: op1_15_inv09 = 1;
    54: op1_15_inv09 = 1;
    69: op1_15_inv09 = 1;
    76: op1_15_inv09 = 1;
    50: op1_15_inv09 = 1;
    77: op1_15_inv09 = 1;
    58: op1_15_inv09 = 1;
    70: op1_15_inv09 = 1;
    79: op1_15_inv09 = 1;
    88: op1_15_inv09 = 1;
    80: op1_15_inv09 = 1;
    81: op1_15_inv09 = 1;
    82: op1_15_inv09 = 1;
    63: op1_15_inv09 = 1;
    89: op1_15_inv09 = 1;
    84: op1_15_inv09 = 1;
    85: op1_15_inv09 = 1;
    90: op1_15_inv09 = 1;
    91: op1_15_inv09 = 1;
    67: op1_15_inv09 = 1;
    92: op1_15_inv09 = 1;
    93: op1_15_inv09 = 1;
    94: op1_15_inv09 = 1;
    95: op1_15_inv09 = 1;
    96: op1_15_inv09 = 1;
    99: op1_15_inv09 = 1;
    101: op1_15_inv09 = 1;
    104: op1_15_inv09 = 1;
    105: op1_15_inv09 = 1;
    106: op1_15_inv09 = 1;
    109: op1_15_inv09 = 1;
    110: op1_15_inv09 = 1;
    111: op1_15_inv09 = 1;
    115: op1_15_inv09 = 1;
    116: op1_15_inv09 = 1;
    118: op1_15_inv09 = 1;
    120: op1_15_inv09 = 1;
    123: op1_15_inv09 = 1;
    124: op1_15_inv09 = 1;
    125: op1_15_inv09 = 1;
    128: op1_15_inv09 = 1;
    default: op1_15_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の10番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in10 = reg_0293;
    73: op1_15_in10 = reg_1404;
    53: op1_15_in10 = reg_0886;
    55: op1_15_in10 = imem07_in[15:12];
    86: op1_15_in10 = reg_0506;
    74: op1_15_in10 = reg_0961;
    54: op1_15_in10 = imem02_in[11:8];
    75: op1_15_in10 = reg_0466;
    69: op1_15_in10 = reg_0712;
    56: op1_15_in10 = reg_0078;
    49: op1_15_in10 = reg_0170;
    76: op1_15_in10 = reg_1515;
    87: op1_15_in10 = reg_0313;
    57: op1_15_in10 = reg_0871;
    50: op1_15_in10 = reg_0989;
    68: op1_15_in10 = reg_0552;
    71: op1_15_in10 = reg_0057;
    77: op1_15_in10 = reg_0585;
    78: op1_15_in10 = reg_0194;
    61: op1_15_in10 = reg_0881;
    119: op1_15_in10 = reg_0881;
    58: op1_15_in10 = reg_0339;
    70: op1_15_in10 = reg_1199;
    59: op1_15_in10 = reg_0632;
    79: op1_15_in10 = reg_1469;
    51: op1_15_in10 = reg_0127;
    60: op1_15_in10 = reg_0924;
    88: op1_15_in10 = reg_1189;
    80: op1_15_in10 = reg_0906;
    103: op1_15_in10 = reg_0906;
    62: op1_15_in10 = reg_1082;
    81: op1_15_in10 = reg_0043;
    82: op1_15_in10 = reg_0395;
    63: op1_15_in10 = reg_0959;
    52: op1_15_in10 = reg_0569;
    83: op1_15_in10 = reg_0839;
    64: op1_15_in10 = reg_0366;
    89: op1_15_in10 = reg_1041;
    91: op1_15_in10 = reg_1041;
    84: op1_15_in10 = reg_0803;
    85: op1_15_in10 = reg_0016;
    65: op1_15_in10 = reg_0935;
    90: op1_15_in10 = reg_0780;
    127: op1_15_in10 = reg_0780;
    66: op1_15_in10 = reg_0114;
    46: op1_15_in10 = reg_0045;
    48: op1_15_in10 = reg_0589;
    67: op1_15_in10 = reg_0351;
    92: op1_15_in10 = reg_0845;
    93: op1_15_in10 = reg_0622;
    94: op1_15_in10 = reg_0507;
    95: op1_15_in10 = reg_0476;
    96: op1_15_in10 = reg_1229;
    97: op1_15_in10 = reg_0300;
    98: op1_15_in10 = reg_0964;
    99: op1_15_in10 = reg_0620;
    100: op1_15_in10 = reg_0733;
    101: op1_15_in10 = reg_1324;
    102: op1_15_in10 = reg_0088;
    104: op1_15_in10 = reg_0221;
    123: op1_15_in10 = reg_0221;
    105: op1_15_in10 = reg_0353;
    106: op1_15_in10 = reg_0322;
    107: op1_15_in10 = reg_0790;
    108: op1_15_in10 = reg_0440;
    109: op1_15_in10 = reg_0575;
    37: op1_15_in10 = imem07_in[11:8];
    110: op1_15_in10 = reg_0111;
    111: op1_15_in10 = reg_0777;
    112: op1_15_in10 = reg_1492;
    113: op1_15_in10 = reg_0072;
    114: op1_15_in10 = reg_1383;
    115: op1_15_in10 = reg_0084;
    116: op1_15_in10 = reg_1149;
    117: op1_15_in10 = reg_0171;
    118: op1_15_in10 = reg_0703;
    47: op1_15_in10 = imem06_in[7:4];
    120: op1_15_in10 = reg_0878;
    121: op1_15_in10 = reg_1083;
    122: op1_15_in10 = reg_0532;
    124: op1_15_in10 = reg_0418;
    125: op1_15_in10 = reg_1321;
    126: op1_15_in10 = reg_0023;
    128: op1_15_in10 = reg_0291;
    129: op1_15_in10 = reg_0538;
    130: op1_15_in10 = reg_0328;
    default: op1_15_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の10番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_15_inv10 = 1;
    53: op1_15_inv10 = 1;
    55: op1_15_inv10 = 1;
    86: op1_15_inv10 = 1;
    74: op1_15_inv10 = 1;
    54: op1_15_inv10 = 1;
    49: op1_15_inv10 = 1;
    50: op1_15_inv10 = 1;
    68: op1_15_inv10 = 1;
    71: op1_15_inv10 = 1;
    61: op1_15_inv10 = 1;
    59: op1_15_inv10 = 1;
    60: op1_15_inv10 = 1;
    62: op1_15_inv10 = 1;
    81: op1_15_inv10 = 1;
    82: op1_15_inv10 = 1;
    63: op1_15_inv10 = 1;
    83: op1_15_inv10 = 1;
    64: op1_15_inv10 = 1;
    89: op1_15_inv10 = 1;
    85: op1_15_inv10 = 1;
    92: op1_15_inv10 = 1;
    93: op1_15_inv10 = 1;
    94: op1_15_inv10 = 1;
    95: op1_15_inv10 = 1;
    96: op1_15_inv10 = 1;
    97: op1_15_inv10 = 1;
    98: op1_15_inv10 = 1;
    100: op1_15_inv10 = 1;
    103: op1_15_inv10 = 1;
    104: op1_15_inv10 = 1;
    105: op1_15_inv10 = 1;
    106: op1_15_inv10 = 1;
    110: op1_15_inv10 = 1;
    112: op1_15_inv10 = 1;
    113: op1_15_inv10 = 1;
    115: op1_15_inv10 = 1;
    116: op1_15_inv10 = 1;
    119: op1_15_inv10 = 1;
    47: op1_15_inv10 = 1;
    121: op1_15_inv10 = 1;
    123: op1_15_inv10 = 1;
    126: op1_15_inv10 = 1;
    128: op1_15_inv10 = 1;
    default: op1_15_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の11番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in11 = reg_0460;
    73: op1_15_in11 = reg_0872;
    53: op1_15_in11 = reg_0638;
    55: op1_15_in11 = reg_0324;
    86: op1_15_in11 = reg_1282;
    128: op1_15_in11 = reg_1282;
    74: op1_15_in11 = reg_1418;
    96: op1_15_in11 = reg_1418;
    54: op1_15_in11 = reg_0455;
    75: op1_15_in11 = reg_1436;
    69: op1_15_in11 = reg_0009;
    56: op1_15_in11 = reg_0291;
    49: op1_15_in11 = reg_0309;
    76: op1_15_in11 = reg_0216;
    87: op1_15_in11 = reg_1280;
    57: op1_15_in11 = reg_0868;
    50: op1_15_in11 = reg_0776;
    68: op1_15_in11 = reg_0412;
    71: op1_15_in11 = reg_0026;
    77: op1_15_in11 = reg_0617;
    78: op1_15_in11 = reg_0586;
    61: op1_15_in11 = reg_0640;
    58: op1_15_in11 = reg_0336;
    70: op1_15_in11 = reg_0505;
    59: op1_15_in11 = reg_1029;
    79: op1_15_in11 = reg_1470;
    51: op1_15_in11 = reg_0380;
    120: op1_15_in11 = reg_0380;
    60: op1_15_in11 = reg_0223;
    88: op1_15_in11 = reg_0904;
    80: op1_15_in11 = reg_0120;
    62: op1_15_in11 = reg_0676;
    81: op1_15_in11 = reg_1492;
    82: op1_15_in11 = reg_1163;
    63: op1_15_in11 = reg_0135;
    52: op1_15_in11 = reg_0527;
    83: op1_15_in11 = reg_0824;
    64: op1_15_in11 = reg_0408;
    89: op1_15_in11 = reg_0342;
    84: op1_15_in11 = reg_1471;
    85: op1_15_in11 = reg_0370;
    65: op1_15_in11 = reg_0903;
    90: op1_15_in11 = reg_0109;
    66: op1_15_in11 = reg_0004;
    91: op1_15_in11 = reg_1065;
    46: op1_15_in11 = reg_0316;
    48: op1_15_in11 = reg_0562;
    67: op1_15_in11 = reg_0060;
    92: op1_15_in11 = reg_1018;
    93: op1_15_in11 = reg_0624;
    94: op1_15_in11 = reg_0999;
    95: op1_15_in11 = reg_0881;
    97: op1_15_in11 = reg_0318;
    98: op1_15_in11 = reg_0190;
    99: op1_15_in11 = reg_0114;
    100: op1_15_in11 = reg_0992;
    101: op1_15_in11 = reg_0089;
    102: op1_15_in11 = reg_0034;
    103: op1_15_in11 = reg_0908;
    47: op1_15_in11 = reg_0908;
    104: op1_15_in11 = reg_1453;
    105: op1_15_in11 = reg_0722;
    106: op1_15_in11 = reg_0659;
    107: op1_15_in11 = reg_0411;
    108: op1_15_in11 = reg_0072;
    109: op1_15_in11 = imem06_in[7:4];
    37: op1_15_in11 = reg_0085;
    110: op1_15_in11 = reg_0382;
    111: op1_15_in11 = reg_0465;
    112: op1_15_in11 = reg_0294;
    113: op1_15_in11 = reg_0871;
    114: op1_15_in11 = reg_0208;
    115: op1_15_in11 = reg_1010;
    116: op1_15_in11 = reg_1325;
    117: op1_15_in11 = reg_0023;
    118: op1_15_in11 = reg_0170;
    119: op1_15_in11 = reg_0886;
    121: op1_15_in11 = reg_1203;
    122: op1_15_in11 = reg_0494;
    123: op1_15_in11 = reg_1230;
    124: op1_15_in11 = reg_0090;
    125: op1_15_in11 = reg_0267;
    126: op1_15_in11 = reg_0046;
    127: op1_15_in11 = reg_0718;
    129: op1_15_in11 = reg_0251;
    130: op1_15_in11 = reg_0797;
    default: op1_15_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の11番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_15_inv11 = 1;
    86: op1_15_inv11 = 1;
    74: op1_15_inv11 = 1;
    54: op1_15_inv11 = 1;
    69: op1_15_inv11 = 1;
    56: op1_15_inv11 = 1;
    49: op1_15_inv11 = 1;
    76: op1_15_inv11 = 1;
    87: op1_15_inv11 = 1;
    68: op1_15_inv11 = 1;
    71: op1_15_inv11 = 1;
    61: op1_15_inv11 = 1;
    58: op1_15_inv11 = 1;
    79: op1_15_inv11 = 1;
    60: op1_15_inv11 = 1;
    62: op1_15_inv11 = 1;
    81: op1_15_inv11 = 1;
    63: op1_15_inv11 = 1;
    83: op1_15_inv11 = 1;
    64: op1_15_inv11 = 1;
    89: op1_15_inv11 = 1;
    84: op1_15_inv11 = 1;
    85: op1_15_inv11 = 1;
    65: op1_15_inv11 = 1;
    66: op1_15_inv11 = 1;
    46: op1_15_inv11 = 1;
    48: op1_15_inv11 = 1;
    67: op1_15_inv11 = 1;
    92: op1_15_inv11 = 1;
    93: op1_15_inv11 = 1;
    94: op1_15_inv11 = 1;
    95: op1_15_inv11 = 1;
    98: op1_15_inv11 = 1;
    99: op1_15_inv11 = 1;
    101: op1_15_inv11 = 1;
    103: op1_15_inv11 = 1;
    104: op1_15_inv11 = 1;
    105: op1_15_inv11 = 1;
    108: op1_15_inv11 = 1;
    110: op1_15_inv11 = 1;
    113: op1_15_inv11 = 1;
    114: op1_15_inv11 = 1;
    115: op1_15_inv11 = 1;
    116: op1_15_inv11 = 1;
    117: op1_15_inv11 = 1;
    119: op1_15_inv11 = 1;
    120: op1_15_inv11 = 1;
    121: op1_15_inv11 = 1;
    123: op1_15_inv11 = 1;
    124: op1_15_inv11 = 1;
    128: op1_15_inv11 = 1;
    129: op1_15_inv11 = 1;
    default: op1_15_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の12番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in12 = reg_1405;
    73: op1_15_in12 = imem05_in[7:4];
    53: op1_15_in12 = reg_0201;
    55: op1_15_in12 = reg_0867;
    86: op1_15_in12 = reg_0427;
    74: op1_15_in12 = reg_1406;
    54: op1_15_in12 = reg_0981;
    75: op1_15_in12 = reg_0730;
    69: op1_15_in12 = reg_0845;
    56: op1_15_in12 = reg_0283;
    49: op1_15_in12 = reg_0157;
    76: op1_15_in12 = reg_1447;
    87: op1_15_in12 = reg_0443;
    57: op1_15_in12 = reg_0278;
    50: op1_15_in12 = reg_0971;
    68: op1_15_in12 = reg_0969;
    71: op1_15_in12 = reg_0005;
    77: op1_15_in12 = reg_0527;
    78: op1_15_in12 = reg_0584;
    61: op1_15_in12 = reg_0075;
    58: op1_15_in12 = reg_0097;
    70: op1_15_in12 = reg_0831;
    59: op1_15_in12 = imem02_in[11:8];
    79: op1_15_in12 = reg_0250;
    51: op1_15_in12 = reg_0138;
    60: op1_15_in12 = reg_0663;
    88: op1_15_in12 = reg_0063;
    80: op1_15_in12 = reg_1209;
    62: op1_15_in12 = reg_0552;
    81: op1_15_in12 = reg_1139;
    82: op1_15_in12 = reg_0996;
    63: op1_15_in12 = reg_0725;
    52: op1_15_in12 = reg_0323;
    83: op1_15_in12 = reg_0876;
    64: op1_15_in12 = reg_0413;
    89: op1_15_in12 = reg_1419;
    84: op1_15_in12 = reg_1053;
    85: op1_15_in12 = reg_0735;
    65: op1_15_in12 = reg_0900;
    90: op1_15_in12 = reg_0717;
    91: op1_15_in12 = reg_0061;
    46: op1_15_in12 = reg_0541;
    48: op1_15_in12 = reg_0531;
    67: op1_15_in12 = reg_1321;
    92: op1_15_in12 = reg_1343;
    93: op1_15_in12 = reg_0528;
    94: op1_15_in12 = reg_0573;
    95: op1_15_in12 = reg_0886;
    96: op1_15_in12 = reg_0927;
    97: op1_15_in12 = reg_0243;
    98: op1_15_in12 = reg_1092;
    99: op1_15_in12 = reg_0521;
    100: op1_15_in12 = reg_0066;
    101: op1_15_in12 = imem01_in[11:8];
    102: op1_15_in12 = reg_0164;
    103: op1_15_in12 = reg_0316;
    104: op1_15_in12 = reg_0134;
    105: op1_15_in12 = reg_0134;
    106: op1_15_in12 = reg_0846;
    107: op1_15_in12 = reg_0129;
    108: op1_15_in12 = reg_0267;
    109: op1_15_in12 = imem06_in[11:8];
    110: op1_15_in12 = reg_0380;
    111: op1_15_in12 = reg_0442;
    112: op1_15_in12 = reg_0903;
    113: op1_15_in12 = reg_1290;
    114: op1_15_in12 = reg_1215;
    115: op1_15_in12 = reg_0310;
    116: op1_15_in12 = reg_0534;
    117: op1_15_in12 = reg_0215;
    126: op1_15_in12 = reg_0215;
    118: op1_15_in12 = reg_0457;
    119: op1_15_in12 = reg_0352;
    47: op1_15_in12 = reg_0696;
    120: op1_15_in12 = reg_0560;
    121: op1_15_in12 = reg_0574;
    122: op1_15_in12 = reg_0429;
    123: op1_15_in12 = reg_1229;
    124: op1_15_in12 = reg_0039;
    125: op1_15_in12 = reg_0917;
    127: op1_15_in12 = reg_1303;
    128: op1_15_in12 = imem04_in[11:8];
    129: op1_15_in12 = reg_0992;
    130: op1_15_in12 = reg_1203;
    default: op1_15_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の12番目の入力反転
  always @ ( * ) begin
    case ( state )
    55: op1_15_inv12 = 1;
    49: op1_15_inv12 = 1;
    76: op1_15_inv12 = 1;
    87: op1_15_inv12 = 1;
    77: op1_15_inv12 = 1;
    78: op1_15_inv12 = 1;
    61: op1_15_inv12 = 1;
    58: op1_15_inv12 = 1;
    79: op1_15_inv12 = 1;
    60: op1_15_inv12 = 1;
    62: op1_15_inv12 = 1;
    82: op1_15_inv12 = 1;
    63: op1_15_inv12 = 1;
    52: op1_15_inv12 = 1;
    64: op1_15_inv12 = 1;
    65: op1_15_inv12 = 1;
    67: op1_15_inv12 = 1;
    92: op1_15_inv12 = 1;
    94: op1_15_inv12 = 1;
    95: op1_15_inv12 = 1;
    96: op1_15_inv12 = 1;
    97: op1_15_inv12 = 1;
    102: op1_15_inv12 = 1;
    103: op1_15_inv12 = 1;
    106: op1_15_inv12 = 1;
    107: op1_15_inv12 = 1;
    109: op1_15_inv12 = 1;
    110: op1_15_inv12 = 1;
    111: op1_15_inv12 = 1;
    115: op1_15_inv12 = 1;
    47: op1_15_inv12 = 1;
    120: op1_15_inv12 = 1;
    121: op1_15_inv12 = 1;
    124: op1_15_inv12 = 1;
    125: op1_15_inv12 = 1;
    127: op1_15_inv12 = 1;
    128: op1_15_inv12 = 1;
    129: op1_15_inv12 = 1;
    default: op1_15_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の13番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in13 = reg_0202;
    73: op1_15_in13 = reg_0275;
    53: op1_15_in13 = reg_0410;
    55: op1_15_in13 = reg_0923;
    86: op1_15_in13 = reg_0696;
    74: op1_15_in13 = reg_0928;
    54: op1_15_in13 = reg_0473;
    75: op1_15_in13 = reg_0316;
    69: op1_15_in13 = reg_0846;
    56: op1_15_in13 = reg_0486;
    49: op1_15_in13 = imem07_in[15:12];
    76: op1_15_in13 = reg_0185;
    87: op1_15_in13 = reg_0341;
    57: op1_15_in13 = reg_0042;
    50: op1_15_in13 = reg_0626;
    68: op1_15_in13 = reg_0370;
    71: op1_15_in13 = reg_0917;
    77: op1_15_in13 = reg_0568;
    78: op1_15_in13 = reg_0619;
    61: op1_15_in13 = reg_0122;
    58: op1_15_in13 = reg_0237;
    70: op1_15_in13 = reg_0330;
    59: op1_15_in13 = imem02_in[15:12];
    79: op1_15_in13 = reg_1027;
    51: op1_15_in13 = reg_0712;
    60: op1_15_in13 = reg_0287;
    88: op1_15_in13 = reg_0095;
    80: op1_15_in13 = reg_0860;
    103: op1_15_in13 = reg_0860;
    62: op1_15_in13 = imem04_in[11:8];
    81: op1_15_in13 = reg_0184;
    82: op1_15_in13 = reg_0648;
    63: op1_15_in13 = reg_0201;
    52: op1_15_in13 = reg_0289;
    83: op1_15_in13 = reg_0897;
    64: op1_15_in13 = reg_0620;
    89: op1_15_in13 = reg_0339;
    84: op1_15_in13 = reg_0250;
    85: op1_15_in13 = reg_1430;
    65: op1_15_in13 = reg_0306;
    90: op1_15_in13 = reg_1303;
    91: op1_15_in13 = reg_0304;
    46: op1_15_in13 = reg_0167;
    48: op1_15_in13 = reg_0495;
    67: op1_15_in13 = reg_0057;
    92: op1_15_in13 = reg_0256;
    93: op1_15_in13 = reg_0419;
    94: op1_15_in13 = reg_1449;
    95: op1_15_in13 = reg_0388;
    96: op1_15_in13 = reg_0722;
    97: op1_15_in13 = reg_0603;
    98: op1_15_in13 = reg_0178;
    100: op1_15_in13 = reg_0604;
    101: op1_15_in13 = reg_1032;
    102: op1_15_in13 = reg_0199;
    104: op1_15_in13 = reg_0073;
    105: op1_15_in13 = reg_0389;
    106: op1_15_in13 = reg_0423;
    107: op1_15_in13 = reg_0898;
    108: op1_15_in13 = reg_1254;
    109: op1_15_in13 = reg_0826;
    110: op1_15_in13 = reg_0560;
    111: op1_15_in13 = reg_0593;
    112: op1_15_in13 = reg_0068;
    113: op1_15_in13 = reg_0576;
    114: op1_15_in13 = reg_0681;
    115: op1_15_in13 = reg_0851;
    116: op1_15_in13 = reg_0531;
    117: op1_15_in13 = reg_0213;
    118: op1_15_in13 = reg_1350;
    119: op1_15_in13 = reg_0440;
    47: op1_15_in13 = reg_0960;
    120: op1_15_in13 = reg_1492;
    121: op1_15_in13 = reg_0281;
    122: op1_15_in13 = reg_0382;
    123: op1_15_in13 = reg_1432;
    124: op1_15_in13 = imem06_in[7:4];
    125: op1_15_in13 = reg_0635;
    126: op1_15_in13 = imem07_in[3:0];
    127: op1_15_in13 = reg_0584;
    128: op1_15_in13 = reg_1384;
    129: op1_15_in13 = reg_1059;
    130: op1_15_in13 = reg_0488;
    default: op1_15_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の13番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_15_inv13 = 1;
    53: op1_15_inv13 = 1;
    55: op1_15_inv13 = 1;
    74: op1_15_inv13 = 1;
    54: op1_15_inv13 = 1;
    75: op1_15_inv13 = 1;
    69: op1_15_inv13 = 1;
    56: op1_15_inv13 = 1;
    87: op1_15_inv13 = 1;
    77: op1_15_inv13 = 1;
    78: op1_15_inv13 = 1;
    58: op1_15_inv13 = 1;
    70: op1_15_inv13 = 1;
    59: op1_15_inv13 = 1;
    88: op1_15_inv13 = 1;
    80: op1_15_inv13 = 1;
    81: op1_15_inv13 = 1;
    82: op1_15_inv13 = 1;
    64: op1_15_inv13 = 1;
    65: op1_15_inv13 = 1;
    90: op1_15_inv13 = 1;
    48: op1_15_inv13 = 1;
    67: op1_15_inv13 = 1;
    92: op1_15_inv13 = 1;
    93: op1_15_inv13 = 1;
    95: op1_15_inv13 = 1;
    97: op1_15_inv13 = 1;
    98: op1_15_inv13 = 1;
    100: op1_15_inv13 = 1;
    101: op1_15_inv13 = 1;
    104: op1_15_inv13 = 1;
    105: op1_15_inv13 = 1;
    108: op1_15_inv13 = 1;
    112: op1_15_inv13 = 1;
    113: op1_15_inv13 = 1;
    114: op1_15_inv13 = 1;
    115: op1_15_inv13 = 1;
    116: op1_15_inv13 = 1;
    47: op1_15_inv13 = 1;
    120: op1_15_inv13 = 1;
    122: op1_15_inv13 = 1;
    124: op1_15_inv13 = 1;
    125: op1_15_inv13 = 1;
    129: op1_15_inv13 = 1;
    130: op1_15_inv13 = 1;
    default: op1_15_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の14番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in14 = reg_0189;
    73: op1_15_in14 = reg_0393;
    53: op1_15_in14 = reg_0058;
    55: op1_15_in14 = reg_0489;
    86: op1_15_in14 = reg_0975;
    74: op1_15_in14 = reg_0431;
    54: op1_15_in14 = reg_0991;
    75: op1_15_in14 = imem06_in[3:0];
    69: op1_15_in14 = reg_0327;
    56: op1_15_in14 = reg_0662;
    49: op1_15_in14 = reg_0030;
    76: op1_15_in14 = reg_0789;
    87: op1_15_in14 = reg_0535;
    57: op1_15_in14 = reg_0041;
    50: op1_15_in14 = reg_0379;
    68: op1_15_in14 = reg_0932;
    71: op1_15_in14 = reg_1100;
    77: op1_15_in14 = reg_0571;
    78: op1_15_in14 = reg_0529;
    61: op1_15_in14 = imem00_in[3:0];
    58: op1_15_in14 = reg_0117;
    70: op1_15_in14 = reg_1282;
    59: op1_15_in14 = reg_0256;
    79: op1_15_in14 = reg_1453;
    51: op1_15_in14 = reg_0708;
    60: op1_15_in14 = reg_0741;
    88: op1_15_in14 = reg_0470;
    80: op1_15_in14 = reg_0869;
    62: op1_15_in14 = reg_0406;
    81: op1_15_in14 = reg_0976;
    82: op1_15_in14 = reg_0649;
    63: op1_15_in14 = reg_0428;
    96: op1_15_in14 = reg_0428;
    52: op1_15_in14 = reg_0459;
    83: op1_15_in14 = reg_0294;
    64: op1_15_in14 = reg_0004;
    89: op1_15_in14 = reg_0096;
    84: op1_15_in14 = reg_0987;
    85: op1_15_in14 = reg_0833;
    65: op1_15_in14 = reg_0877;
    90: op1_15_in14 = reg_0194;
    91: op1_15_in14 = reg_0339;
    46: op1_15_in14 = reg_0163;
    48: op1_15_in14 = reg_0990;
    67: op1_15_in14 = reg_0005;
    92: op1_15_in14 = reg_0054;
    93: op1_15_in14 = reg_0119;
    94: op1_15_in14 = reg_1447;
    95: op1_15_in14 = reg_0387;
    97: op1_15_in14 = reg_0317;
    98: op1_15_in14 = reg_0541;
    100: op1_15_in14 = reg_0045;
    101: op1_15_in14 = reg_1512;
    102: op1_15_in14 = reg_0454;
    103: op1_15_in14 = reg_0720;
    104: op1_15_in14 = reg_0060;
    105: op1_15_in14 = reg_0980;
    106: op1_15_in14 = reg_0056;
    107: op1_15_in14 = reg_0577;
    108: op1_15_in14 = reg_1256;
    109: op1_15_in14 = reg_0784;
    110: op1_15_in14 = reg_1098;
    120: op1_15_in14 = reg_1098;
    111: op1_15_in14 = reg_0592;
    112: op1_15_in14 = reg_0227;
    113: op1_15_in14 = reg_0743;
    114: op1_15_in14 = reg_0268;
    115: op1_15_in14 = reg_0457;
    116: op1_15_in14 = reg_0574;
    117: op1_15_in14 = imem07_in[3:0];
    118: op1_15_in14 = reg_1347;
    119: op1_15_in14 = reg_0134;
    47: op1_15_in14 = reg_0716;
    121: op1_15_in14 = reg_0500;
    122: op1_15_in14 = reg_1140;
    123: op1_15_in14 = reg_1418;
    124: op1_15_in14 = reg_0905;
    125: op1_15_in14 = reg_0985;
    126: op1_15_in14 = imem07_in[7:4];
    127: op1_15_in14 = reg_0527;
    128: op1_15_in14 = reg_1372;
    129: op1_15_in14 = reg_0793;
    130: op1_15_in14 = reg_0681;
    default: op1_15_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の14番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv14 = 1;
    53: op1_15_inv14 = 1;
    55: op1_15_inv14 = 1;
    56: op1_15_inv14 = 1;
    49: op1_15_inv14 = 1;
    76: op1_15_inv14 = 1;
    87: op1_15_inv14 = 1;
    50: op1_15_inv14 = 1;
    77: op1_15_inv14 = 1;
    79: op1_15_inv14 = 1;
    62: op1_15_inv14 = 1;
    82: op1_15_inv14 = 1;
    63: op1_15_inv14 = 1;
    52: op1_15_inv14 = 1;
    83: op1_15_inv14 = 1;
    89: op1_15_inv14 = 1;
    85: op1_15_inv14 = 1;
    90: op1_15_inv14 = 1;
    92: op1_15_inv14 = 1;
    95: op1_15_inv14 = 1;
    100: op1_15_inv14 = 1;
    101: op1_15_inv14 = 1;
    102: op1_15_inv14 = 1;
    103: op1_15_inv14 = 1;
    104: op1_15_inv14 = 1;
    105: op1_15_inv14 = 1;
    107: op1_15_inv14 = 1;
    109: op1_15_inv14 = 1;
    112: op1_15_inv14 = 1;
    115: op1_15_inv14 = 1;
    116: op1_15_inv14 = 1;
    118: op1_15_inv14 = 1;
    121: op1_15_inv14 = 1;
    125: op1_15_inv14 = 1;
    128: op1_15_inv14 = 1;
    default: op1_15_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の15番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in15 = reg_0428;
    73: op1_15_in15 = reg_0602;
    53: op1_15_in15 = reg_0089;
    55: op1_15_in15 = reg_0140;
    86: op1_15_in15 = reg_0534;
    74: op1_15_in15 = reg_0060;
    95: op1_15_in15 = reg_0060;
    54: op1_15_in15 = reg_0432;
    48: op1_15_in15 = reg_0432;
    75: op1_15_in15 = reg_0859;
    69: op1_15_in15 = reg_0632;
    56: op1_15_in15 = reg_0742;
    49: op1_15_in15 = reg_0366;
    76: op1_15_in15 = reg_1517;
    87: op1_15_in15 = reg_0264;
    57: op1_15_in15 = reg_0012;
    50: op1_15_in15 = reg_0381;
    68: op1_15_in15 = reg_0451;
    71: op1_15_in15 = reg_0611;
    77: op1_15_in15 = reg_0979;
    78: op1_15_in15 = reg_0527;
    61: op1_15_in15 = imem01_in[3:0];
    58: op1_15_in15 = reg_0211;
    70: op1_15_in15 = reg_1280;
    59: op1_15_in15 = reg_0474;
    79: op1_15_in15 = reg_1227;
    51: op1_15_in15 = reg_0711;
    60: op1_15_in15 = reg_0593;
    88: op1_15_in15 = reg_0251;
    80: op1_15_in15 = reg_1501;
    62: op1_15_in15 = reg_0969;
    81: op1_15_in15 = reg_0607;
    82: op1_15_in15 = reg_0182;
    63: op1_15_in15 = reg_0435;
    96: op1_15_in15 = reg_0435;
    52: op1_15_in15 = reg_0269;
    83: op1_15_in15 = reg_0327;
    64: op1_15_in15 = reg_0002;
    89: op1_15_in15 = reg_0020;
    84: op1_15_in15 = reg_0927;
    85: op1_15_in15 = reg_0832;
    65: op1_15_in15 = reg_0009;
    90: op1_15_in15 = reg_0141;
    91: op1_15_in15 = reg_0336;
    46: op1_15_in15 = reg_0873;
    67: op1_15_in15 = reg_0723;
    92: op1_15_in15 = reg_0127;
    93: op1_15_in15 = reg_0165;
    94: op1_15_in15 = reg_0216;
    97: op1_15_in15 = reg_0206;
    98: op1_15_in15 = reg_1009;
    100: op1_15_in15 = reg_0630;
    101: op1_15_in15 = reg_0553;
    102: op1_15_in15 = reg_0061;
    103: op1_15_in15 = reg_0869;
    109: op1_15_in15 = reg_0869;
    104: op1_15_in15 = reg_0372;
    105: op1_15_in15 = reg_1253;
    106: op1_15_in15 = reg_0276;
    107: op1_15_in15 = reg_1257;
    108: op1_15_in15 = reg_0093;
    110: op1_15_in15 = reg_0007;
    111: op1_15_in15 = reg_0103;
    112: op1_15_in15 = reg_0989;
    113: op1_15_in15 = reg_0798;
    114: op1_15_in15 = reg_1151;
    115: op1_15_in15 = reg_1345;
    116: op1_15_in15 = reg_1237;
    117: op1_15_in15 = imem07_in[7:4];
    118: op1_15_in15 = reg_0921;
    119: op1_15_in15 = reg_0389;
    47: op1_15_in15 = reg_0568;
    120: op1_15_in15 = reg_0801;
    121: op1_15_in15 = reg_0094;
    122: op1_15_in15 = reg_0829;
    123: op1_15_in15 = reg_0821;
    124: op1_15_in15 = reg_0133;
    125: op1_15_in15 = reg_1290;
    126: op1_15_in15 = reg_1183;
    127: op1_15_in15 = reg_0570;
    128: op1_15_in15 = reg_1338;
    129: op1_15_in15 = reg_0173;
    130: op1_15_in15 = reg_1233;
    default: op1_15_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の15番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv15 = 1;
    73: op1_15_inv15 = 1;
    55: op1_15_inv15 = 1;
    86: op1_15_inv15 = 1;
    74: op1_15_inv15 = 1;
    54: op1_15_inv15 = 1;
    75: op1_15_inv15 = 1;
    76: op1_15_inv15 = 1;
    87: op1_15_inv15 = 1;
    57: op1_15_inv15 = 1;
    68: op1_15_inv15 = 1;
    77: op1_15_inv15 = 1;
    59: op1_15_inv15 = 1;
    79: op1_15_inv15 = 1;
    51: op1_15_inv15 = 1;
    88: op1_15_inv15 = 1;
    62: op1_15_inv15 = 1;
    81: op1_15_inv15 = 1;
    52: op1_15_inv15 = 1;
    83: op1_15_inv15 = 1;
    64: op1_15_inv15 = 1;
    89: op1_15_inv15 = 1;
    84: op1_15_inv15 = 1;
    85: op1_15_inv15 = 1;
    65: op1_15_inv15 = 1;
    48: op1_15_inv15 = 1;
    92: op1_15_inv15 = 1;
    101: op1_15_inv15 = 1;
    102: op1_15_inv15 = 1;
    103: op1_15_inv15 = 1;
    104: op1_15_inv15 = 1;
    108: op1_15_inv15 = 1;
    109: op1_15_inv15 = 1;
    110: op1_15_inv15 = 1;
    111: op1_15_inv15 = 1;
    112: op1_15_inv15 = 1;
    113: op1_15_inv15 = 1;
    114: op1_15_inv15 = 1;
    117: op1_15_inv15 = 1;
    118: op1_15_inv15 = 1;
    119: op1_15_inv15 = 1;
    47: op1_15_inv15 = 1;
    120: op1_15_inv15 = 1;
    121: op1_15_inv15 = 1;
    123: op1_15_inv15 = 1;
    124: op1_15_inv15 = 1;
    126: op1_15_inv15 = 1;
    127: op1_15_inv15 = 1;
    128: op1_15_inv15 = 1;
    default: op1_15_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の16番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in16 = reg_0388;
    73: op1_15_in16 = reg_0797;
    53: op1_15_in16 = reg_0005;
    55: op1_15_in16 = reg_0779;
    86: op1_15_in16 = reg_0032;
    74: op1_15_in16 = reg_0059;
    54: op1_15_in16 = reg_0054;
    75: op1_15_in16 = reg_0718;
    69: op1_15_in16 = reg_0800;
    120: op1_15_in16 = reg_0800;
    56: op1_15_in16 = reg_0255;
    49: op1_15_in16 = reg_0738;
    76: op1_15_in16 = reg_0048;
    87: op1_15_in16 = reg_1083;
    57: op1_15_in16 = reg_0222;
    50: op1_15_in16 = reg_0153;
    68: op1_15_in16 = reg_0339;
    71: op1_15_in16 = reg_1291;
    67: op1_15_in16 = reg_1291;
    77: op1_15_in16 = reg_0522;
    78: op1_15_in16 = reg_0571;
    61: op1_15_in16 = imem01_in[15:12];
    58: op1_15_in16 = reg_0792;
    70: op1_15_in16 = reg_0348;
    59: op1_15_in16 = reg_0436;
    79: op1_15_in16 = reg_1205;
    51: op1_15_in16 = reg_0306;
    60: op1_15_in16 = reg_0100;
    88: op1_15_in16 = reg_0702;
    80: op1_15_in16 = imem06_in[15:12];
    62: op1_15_in16 = reg_0936;
    81: op1_15_in16 = reg_0253;
    82: op1_15_in16 = reg_0697;
    63: op1_15_in16 = reg_0409;
    52: op1_15_in16 = reg_0271;
    83: op1_15_in16 = reg_0008;
    64: op1_15_in16 = reg_0053;
    89: op1_15_in16 = reg_1163;
    84: op1_15_in16 = reg_1393;
    85: op1_15_in16 = reg_0273;
    65: op1_15_in16 = reg_0802;
    90: op1_15_in16 = reg_0619;
    91: op1_15_in16 = reg_1151;
    46: op1_15_in16 = reg_0196;
    48: op1_15_in16 = reg_0433;
    92: op1_15_in16 = reg_0106;
    93: op1_15_in16 = reg_0269;
    94: op1_15_in16 = reg_0311;
    95: op1_15_in16 = reg_0917;
    96: op1_15_in16 = reg_0387;
    97: op1_15_in16 = reg_0040;
    98: op1_15_in16 = imem04_in[7:4];
    100: op1_15_in16 = reg_1180;
    101: op1_15_in16 = reg_0550;
    102: op1_15_in16 = reg_0369;
    103: op1_15_in16 = reg_1323;
    104: op1_15_in16 = reg_1255;
    105: op1_15_in16 = reg_1152;
    106: op1_15_in16 = reg_0133;
    107: op1_15_in16 = reg_1258;
    108: op1_15_in16 = reg_0463;
    109: op1_15_in16 = reg_0109;
    110: op1_15_in16 = reg_1006;
    111: op1_15_in16 = reg_0228;
    112: op1_15_in16 = reg_0759;
    113: op1_15_in16 = reg_0820;
    114: op1_15_in16 = reg_0536;
    115: op1_15_in16 = reg_0159;
    116: op1_15_in16 = reg_1503;
    117: op1_15_in16 = imem07_in[15:12];
    118: op1_15_in16 = reg_0489;
    119: op1_15_in16 = reg_0577;
    47: op1_15_in16 = reg_0171;
    121: op1_15_in16 = reg_0414;
    122: op1_15_in16 = reg_0801;
    123: op1_15_in16 = reg_0202;
    124: op1_15_in16 = reg_0870;
    125: op1_15_in16 = reg_0576;
    126: op1_15_in16 = reg_0478;
    127: op1_15_in16 = reg_0132;
    128: op1_15_in16 = reg_0699;
    129: op1_15_in16 = reg_0391;
    130: op1_15_in16 = reg_0094;
    default: op1_15_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の16番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv16 = 1;
    53: op1_15_inv16 = 1;
    55: op1_15_inv16 = 1;
    49: op1_15_inv16 = 1;
    76: op1_15_inv16 = 1;
    57: op1_15_inv16 = 1;
    68: op1_15_inv16 = 1;
    71: op1_15_inv16 = 1;
    77: op1_15_inv16 = 1;
    78: op1_15_inv16 = 1;
    61: op1_15_inv16 = 1;
    58: op1_15_inv16 = 1;
    59: op1_15_inv16 = 1;
    51: op1_15_inv16 = 1;
    60: op1_15_inv16 = 1;
    88: op1_15_inv16 = 1;
    80: op1_15_inv16 = 1;
    62: op1_15_inv16 = 1;
    81: op1_15_inv16 = 1;
    63: op1_15_inv16 = 1;
    89: op1_15_inv16 = 1;
    90: op1_15_inv16 = 1;
    91: op1_15_inv16 = 1;
    46: op1_15_inv16 = 1;
    67: op1_15_inv16 = 1;
    93: op1_15_inv16 = 1;
    95: op1_15_inv16 = 1;
    98: op1_15_inv16 = 1;
    103: op1_15_inv16 = 1;
    106: op1_15_inv16 = 1;
    107: op1_15_inv16 = 1;
    108: op1_15_inv16 = 1;
    109: op1_15_inv16 = 1;
    114: op1_15_inv16 = 1;
    115: op1_15_inv16 = 1;
    116: op1_15_inv16 = 1;
    119: op1_15_inv16 = 1;
    47: op1_15_inv16 = 1;
    126: op1_15_inv16 = 1;
    129: op1_15_inv16 = 1;
    default: op1_15_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の17番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in17 = reg_0073;
    73: op1_15_in17 = reg_0828;
    53: op1_15_in17 = reg_0610;
    55: op1_15_in17 = reg_0442;
    86: op1_15_in17 = reg_0181;
    74: op1_15_in17 = reg_1321;
    54: op1_15_in17 = reg_0776;
    75: op1_15_in17 = reg_0373;
    69: op1_15_in17 = reg_0279;
    56: op1_15_in17 = reg_0976;
    49: op1_15_in17 = reg_0623;
    76: op1_15_in17 = reg_1301;
    87: op1_15_in17 = reg_1198;
    107: op1_15_in17 = reg_1198;
    57: op1_15_in17 = reg_0446;
    50: op1_15_in17 = reg_0877;
    68: op1_15_in17 = reg_0064;
    71: op1_15_in17 = reg_1256;
    77: op1_15_in17 = reg_0171;
    78: op1_15_in17 = reg_0345;
    61: op1_15_in17 = reg_1290;
    119: op1_15_in17 = reg_1290;
    58: op1_15_in17 = reg_1104;
    70: op1_15_in17 = reg_0411;
    59: op1_15_in17 = reg_0127;
    79: op1_15_in17 = reg_1406;
    51: op1_15_in17 = reg_0878;
    60: op1_15_in17 = reg_0114;
    88: op1_15_in17 = reg_0332;
    80: op1_15_in17 = reg_0716;
    62: op1_15_in17 = reg_0369;
    81: op1_15_in17 = reg_1074;
    82: op1_15_in17 = reg_1401;
    63: op1_15_in17 = reg_0353;
    52: op1_15_in17 = reg_0213;
    83: op1_15_in17 = reg_1392;
    64: op1_15_in17 = reg_0085;
    89: op1_15_in17 = reg_0562;
    84: op1_15_in17 = reg_0202;
    85: op1_15_in17 = reg_0879;
    65: op1_15_in17 = reg_0281;
    90: op1_15_in17 = reg_0529;
    91: op1_15_in17 = reg_1189;
    46: op1_15_in17 = reg_0274;
    48: op1_15_in17 = reg_0429;
    67: op1_15_in17 = reg_1071;
    92: op1_15_in17 = reg_0684;
    93: op1_15_in17 = reg_0015;
    94: op1_15_in17 = reg_1184;
    95: op1_15_in17 = reg_1291;
    96: op1_15_in17 = reg_0075;
    97: op1_15_in17 = reg_0039;
    98: op1_15_in17 = reg_1312;
    100: op1_15_in17 = reg_1402;
    101: op1_15_in17 = reg_0798;
    102: op1_15_in17 = reg_0062;
    103: op1_15_in17 = reg_1501;
    104: op1_15_in17 = reg_1254;
    105: op1_15_in17 = reg_0463;
    106: op1_15_in17 = reg_0712;
    108: op1_15_in17 = reg_1473;
    113: op1_15_in17 = reg_1473;
    109: op1_15_in17 = reg_0717;
    110: op1_15_in17 = reg_0009;
    111: op1_15_in17 = reg_0051;
    112: op1_15_in17 = reg_0573;
    114: op1_15_in17 = reg_0538;
    115: op1_15_in17 = reg_0156;
    116: op1_15_in17 = reg_1488;
    117: op1_15_in17 = reg_1096;
    118: op1_15_in17 = reg_0777;
    47: op1_15_in17 = reg_0271;
    120: op1_15_in17 = reg_0168;
    121: op1_15_in17 = reg_0406;
    122: op1_15_in17 = reg_0903;
    123: op1_15_in17 = reg_0409;
    124: op1_15_in17 = reg_0265;
    125: op1_15_in17 = reg_0549;
    126: op1_15_in17 = reg_0219;
    127: op1_15_in17 = reg_0295;
    128: op1_15_in17 = reg_0164;
    129: op1_15_in17 = reg_0491;
    130: op1_15_in17 = reg_0421;
    default: op1_15_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の17番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_15_inv17 = 1;
    53: op1_15_inv17 = 1;
    86: op1_15_inv17 = 1;
    74: op1_15_inv17 = 1;
    54: op1_15_inv17 = 1;
    69: op1_15_inv17 = 1;
    56: op1_15_inv17 = 1;
    49: op1_15_inv17 = 1;
    76: op1_15_inv17 = 1;
    87: op1_15_inv17 = 1;
    57: op1_15_inv17 = 1;
    50: op1_15_inv17 = 1;
    68: op1_15_inv17 = 1;
    77: op1_15_inv17 = 1;
    61: op1_15_inv17 = 1;
    70: op1_15_inv17 = 1;
    59: op1_15_inv17 = 1;
    79: op1_15_inv17 = 1;
    88: op1_15_inv17 = 1;
    81: op1_15_inv17 = 1;
    63: op1_15_inv17 = 1;
    64: op1_15_inv17 = 1;
    89: op1_15_inv17 = 1;
    84: op1_15_inv17 = 1;
    85: op1_15_inv17 = 1;
    65: op1_15_inv17 = 1;
    90: op1_15_inv17 = 1;
    67: op1_15_inv17 = 1;
    92: op1_15_inv17 = 1;
    94: op1_15_inv17 = 1;
    97: op1_15_inv17 = 1;
    98: op1_15_inv17 = 1;
    103: op1_15_inv17 = 1;
    105: op1_15_inv17 = 1;
    106: op1_15_inv17 = 1;
    107: op1_15_inv17 = 1;
    110: op1_15_inv17 = 1;
    111: op1_15_inv17 = 1;
    113: op1_15_inv17 = 1;
    114: op1_15_inv17 = 1;
    115: op1_15_inv17 = 1;
    117: op1_15_inv17 = 1;
    118: op1_15_inv17 = 1;
    119: op1_15_inv17 = 1;
    47: op1_15_inv17 = 1;
    120: op1_15_inv17 = 1;
    123: op1_15_inv17 = 1;
    127: op1_15_inv17 = 1;
    128: op1_15_inv17 = 1;
    129: op1_15_inv17 = 1;
    130: op1_15_inv17 = 1;
    default: op1_15_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の18番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in18 = reg_0075;
    73: op1_15_in18 = reg_0207;
    53: op1_15_in18 = reg_0786;
    55: op1_15_in18 = reg_0050;
    86: op1_15_in18 = imem04_in[15:12];
    74: op1_15_in18 = reg_1324;
    54: op1_15_in18 = reg_0971;
    75: op1_15_in18 = reg_0529;
    69: op1_15_in18 = reg_0755;
    56: op1_15_in18 = reg_0563;
    49: op1_15_in18 = reg_0620;
    76: op1_15_in18 = reg_0113;
    87: op1_15_in18 = reg_1233;
    57: op1_15_in18 = reg_0744;
    106: op1_15_in18 = reg_0744;
    50: op1_15_in18 = reg_0024;
    68: op1_15_in18 = reg_0035;
    71: op1_15_in18 = reg_1068;
    77: op1_15_in18 = reg_0371;
    78: op1_15_in18 = reg_0979;
    61: op1_15_in18 = reg_1256;
    58: op1_15_in18 = reg_1168;
    70: op1_15_in18 = reg_0898;
    59: op1_15_in18 = reg_0112;
    79: op1_15_in18 = reg_0881;
    51: op1_15_in18 = reg_0839;
    60: op1_15_in18 = reg_0086;
    88: op1_15_in18 = reg_0996;
    80: op1_15_in18 = reg_0585;
    62: op1_15_in18 = reg_0305;
    81: op1_15_in18 = reg_0776;
    82: op1_15_in18 = reg_0938;
    63: op1_15_in18 = reg_1322;
    52: op1_15_in18 = reg_0457;
    83: op1_15_in18 = reg_0848;
    64: op1_15_in18 = reg_0087;
    89: op1_15_in18 = reg_0173;
    84: op1_15_in18 = reg_0435;
    85: op1_15_in18 = imem05_in[11:8];
    65: op1_15_in18 = reg_0276;
    90: op1_15_in18 = reg_0570;
    91: op1_15_in18 = reg_0211;
    46: op1_15_in18 = reg_0151;
    48: op1_15_in18 = reg_0127;
    67: op1_15_in18 = reg_0548;
    92: op1_15_in18 = reg_0628;
    93: op1_15_in18 = reg_1351;
    94: op1_15_in18 = reg_0142;
    95: op1_15_in18 = reg_1032;
    96: op1_15_in18 = reg_0089;
    97: op1_15_in18 = reg_0265;
    98: op1_15_in18 = reg_0319;
    100: op1_15_in18 = reg_1070;
    101: op1_15_in18 = reg_0967;
    102: op1_15_in18 = reg_0262;
    103: op1_15_in18 = reg_1504;
    104: op1_15_in18 = reg_0093;
    105: op1_15_in18 = reg_0163;
    107: op1_15_in18 = reg_0574;
    108: op1_15_in18 = reg_1474;
    109: op1_15_in18 = reg_1302;
    110: op1_15_in18 = reg_0732;
    111: op1_15_in18 = reg_0052;
    112: op1_15_in18 = reg_0234;
    113: op1_15_in18 = reg_0612;
    114: op1_15_in18 = reg_0338;
    115: op1_15_in18 = reg_0921;
    116: op1_15_in18 = reg_0540;
    117: op1_15_in18 = reg_0051;
    118: op1_15_in18 = reg_0774;
    119: op1_15_in18 = reg_0902;
    47: op1_15_in18 = reg_0230;
    120: op1_15_in18 = reg_0006;
    121: op1_15_in18 = reg_1065;
    122: op1_15_in18 = reg_0824;
    123: op1_15_in18 = reg_0388;
    124: op1_15_in18 = reg_0115;
    125: op1_15_in18 = reg_0743;
    126: op1_15_in18 = reg_0225;
    127: op1_15_in18 = reg_0419;
    128: op1_15_in18 = reg_0088;
    129: op1_15_in18 = reg_0167;
    130: op1_15_in18 = reg_0969;
    default: op1_15_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の18番目の入力反転
  always @ ( * ) begin
    case ( state )
    73: op1_15_inv18 = 1;
    55: op1_15_inv18 = 1;
    69: op1_15_inv18 = 1;
    49: op1_15_inv18 = 1;
    76: op1_15_inv18 = 1;
    87: op1_15_inv18 = 1;
    50: op1_15_inv18 = 1;
    71: op1_15_inv18 = 1;
    78: op1_15_inv18 = 1;
    61: op1_15_inv18 = 1;
    51: op1_15_inv18 = 1;
    60: op1_15_inv18 = 1;
    88: op1_15_inv18 = 1;
    62: op1_15_inv18 = 1;
    83: op1_15_inv18 = 1;
    89: op1_15_inv18 = 1;
    84: op1_15_inv18 = 1;
    65: op1_15_inv18 = 1;
    91: op1_15_inv18 = 1;
    46: op1_15_inv18 = 1;
    48: op1_15_inv18 = 1;
    67: op1_15_inv18 = 1;
    92: op1_15_inv18 = 1;
    96: op1_15_inv18 = 1;
    97: op1_15_inv18 = 1;
    103: op1_15_inv18 = 1;
    105: op1_15_inv18 = 1;
    108: op1_15_inv18 = 1;
    109: op1_15_inv18 = 1;
    110: op1_15_inv18 = 1;
    111: op1_15_inv18 = 1;
    114: op1_15_inv18 = 1;
    115: op1_15_inv18 = 1;
    116: op1_15_inv18 = 1;
    118: op1_15_inv18 = 1;
    119: op1_15_inv18 = 1;
    120: op1_15_inv18 = 1;
    121: op1_15_inv18 = 1;
    122: op1_15_inv18 = 1;
    123: op1_15_inv18 = 1;
    125: op1_15_inv18 = 1;
    127: op1_15_inv18 = 1;
    128: op1_15_inv18 = 1;
    129: op1_15_inv18 = 1;
    default: op1_15_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の19番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in19 = reg_0060;
    73: op1_15_in19 = reg_0040;
    53: op1_15_in19 = reg_0335;
    86: op1_15_in19 = reg_1257;
    74: op1_15_in19 = reg_0089;
    54: op1_15_in19 = reg_0933;
    75: op1_15_in19 = reg_1228;
    90: op1_15_in19 = reg_1228;
    69: op1_15_in19 = reg_0732;
    56: op1_15_in19 = reg_0561;
    49: op1_15_in19 = reg_0103;
    76: op1_15_in19 = reg_0880;
    87: op1_15_in19 = reg_1214;
    57: op1_15_in19 = reg_0255;
    122: op1_15_in19 = reg_0255;
    50: op1_15_in19 = reg_0800;
    68: op1_15_in19 = reg_0034;
    71: op1_15_in19 = reg_0420;
    67: op1_15_in19 = reg_0420;
    77: op1_15_in19 = reg_1170;
    78: op1_15_in19 = reg_0296;
    61: op1_15_in19 = reg_1068;
    58: op1_15_in19 = reg_1164;
    85: op1_15_in19 = reg_1164;
    70: op1_15_in19 = reg_0696;
    59: op1_15_in19 = reg_0106;
    79: op1_15_in19 = reg_0883;
    51: op1_15_in19 = reg_0006;
    60: op1_15_in19 = reg_0084;
    88: op1_15_in19 = reg_0174;
    80: op1_15_in19 = reg_0622;
    62: op1_15_in19 = reg_0835;
    81: op1_15_in19 = reg_0971;
    82: op1_15_in19 = reg_1486;
    63: op1_15_in19 = reg_0005;
    52: op1_15_in19 = imem07_in[15:12];
    47: op1_15_in19 = imem07_in[15:12];
    83: op1_15_in19 = reg_1078;
    89: op1_15_in19 = reg_0491;
    84: op1_15_in19 = reg_0387;
    123: op1_15_in19 = reg_0387;
    65: op1_15_in19 = reg_0758;
    91: op1_15_in19 = reg_0117;
    46: op1_15_in19 = reg_0204;
    48: op1_15_in19 = reg_0111;
    92: op1_15_in19 = reg_0897;
    93: op1_15_in19 = imem07_in[3:0];
    94: op1_15_in19 = reg_0957;
    95: op1_15_in19 = reg_1253;
    96: op1_15_in19 = reg_0734;
    97: op1_15_in19 = reg_0825;
    98: op1_15_in19 = reg_0467;
    100: op1_15_in19 = reg_0939;
    101: op1_15_in19 = reg_0819;
    102: op1_15_in19 = reg_1189;
    103: op1_15_in19 = reg_1179;
    104: op1_15_in19 = reg_0830;
    105: op1_15_in19 = reg_0331;
    106: op1_15_in19 = reg_0497;
    107: op1_15_in19 = reg_0094;
    108: op1_15_in19 = reg_0715;
    109: op1_15_in19 = reg_0398;
    110: op1_15_in19 = reg_0444;
    111: op1_15_in19 = reg_0053;
    112: op1_15_in19 = reg_0789;
    113: op1_15_in19 = reg_1475;
    114: op1_15_in19 = reg_0136;
    115: op1_15_in19 = reg_0777;
    116: op1_15_in19 = imem05_in[7:4];
    117: op1_15_in19 = reg_1095;
    118: op1_15_in19 = reg_0465;
    119: op1_15_in19 = reg_0930;
    120: op1_15_in19 = reg_0328;
    121: op1_15_in19 = reg_0454;
    124: op1_15_in19 = reg_0585;
    125: op1_15_in19 = reg_0609;
    126: op1_15_in19 = reg_0299;
    127: op1_15_in19 = reg_0308;
    128: op1_15_in19 = reg_1258;
    129: op1_15_in19 = reg_1181;
    130: op1_15_in19 = reg_1041;
    default: op1_15_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の19番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv19 = 1;
    73: op1_15_inv19 = 1;
    86: op1_15_inv19 = 1;
    74: op1_15_inv19 = 1;
    54: op1_15_inv19 = 1;
    75: op1_15_inv19 = 1;
    49: op1_15_inv19 = 1;
    50: op1_15_inv19 = 1;
    68: op1_15_inv19 = 1;
    78: op1_15_inv19 = 1;
    70: op1_15_inv19 = 1;
    51: op1_15_inv19 = 1;
    88: op1_15_inv19 = 1;
    62: op1_15_inv19 = 1;
    81: op1_15_inv19 = 1;
    63: op1_15_inv19 = 1;
    83: op1_15_inv19 = 1;
    89: op1_15_inv19 = 1;
    48: op1_15_inv19 = 1;
    94: op1_15_inv19 = 1;
    101: op1_15_inv19 = 1;
    105: op1_15_inv19 = 1;
    107: op1_15_inv19 = 1;
    113: op1_15_inv19 = 1;
    114: op1_15_inv19 = 1;
    116: op1_15_inv19 = 1;
    117: op1_15_inv19 = 1;
    118: op1_15_inv19 = 1;
    47: op1_15_inv19 = 1;
    123: op1_15_inv19 = 1;
    124: op1_15_inv19 = 1;
    127: op1_15_inv19 = 1;
    128: op1_15_inv19 = 1;
    default: op1_15_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の20番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in20 = reg_1321;
    73: op1_15_in20 = reg_0466;
    53: op1_15_in20 = reg_1033;
    86: op1_15_in20 = reg_1258;
    74: op1_15_in20 = reg_1100;
    54: op1_15_in20 = reg_0106;
    75: op1_15_in20 = reg_0419;
    69: op1_15_in20 = reg_0191;
    56: op1_15_in20 = reg_0981;
    49: op1_15_in20 = reg_0050;
    76: op1_15_in20 = reg_0478;
    87: op1_15_in20 = reg_0421;
    57: op1_15_in20 = reg_0253;
    50: op1_15_in20 = reg_0313;
    68: op1_15_in20 = reg_1298;
    71: op1_15_in20 = reg_0984;
    77: op1_15_in20 = reg_1441;
    78: op1_15_in20 = reg_0289;
    61: op1_15_in20 = reg_0611;
    58: op1_15_in20 = reg_1169;
    85: op1_15_in20 = reg_1169;
    70: op1_15_in20 = reg_1312;
    59: op1_15_in20 = reg_0153;
    79: op1_15_in20 = reg_0352;
    51: op1_15_in20 = reg_0830;
    60: op1_15_in20 = reg_0124;
    88: op1_15_in20 = reg_1104;
    80: op1_15_in20 = reg_0979;
    62: op1_15_in20 = reg_0065;
    81: op1_15_in20 = reg_1458;
    82: op1_15_in20 = reg_0118;
    63: op1_15_in20 = imem01_in[15:12];
    52: op1_15_in20 = reg_0245;
    83: op1_15_in20 = reg_0312;
    89: op1_15_in20 = reg_0566;
    84: op1_15_in20 = reg_0058;
    65: op1_15_in20 = reg_0216;
    90: op1_15_in20 = reg_1225;
    91: op1_15_in20 = reg_0064;
    46: op1_15_in20 = reg_0038;
    48: op1_15_in20 = reg_0381;
    67: op1_15_in20 = reg_0238;
    92: op1_15_in20 = reg_0802;
    93: op1_15_in20 = imem07_in[11:8];
    94: op1_15_in20 = reg_0108;
    95: op1_15_in20 = reg_0963;
    120: op1_15_in20 = reg_0963;
    96: op1_15_in20 = reg_0239;
    97: op1_15_in20 = reg_0905;
    98: op1_15_in20 = reg_1383;
    100: op1_15_in20 = reg_0794;
    101: op1_15_in20 = reg_1457;
    102: op1_15_in20 = reg_0904;
    103: op1_15_in20 = reg_1508;
    104: op1_15_in20 = reg_1474;
    113: op1_15_in20 = reg_1474;
    105: op1_15_in20 = reg_0610;
    106: op1_15_in20 = reg_0256;
    107: op1_15_in20 = reg_0407;
    108: op1_15_in20 = reg_0819;
    109: op1_15_in20 = reg_0624;
    110: op1_15_in20 = reg_0573;
    112: op1_15_in20 = reg_0314;
    114: op1_15_in20 = reg_0700;
    115: op1_15_in20 = reg_0031;
    116: op1_15_in20 = reg_1059;
    117: op1_15_in20 = reg_1010;
    118: op1_15_in20 = reg_0441;
    119: op1_15_in20 = reg_0047;
    47: op1_15_in20 = reg_0224;
    121: op1_15_in20 = reg_0033;
    122: op1_15_in20 = imem03_in[15:12];
    123: op1_15_in20 = reg_0057;
    124: op1_15_in20 = reg_1228;
    125: op1_15_in20 = reg_0798;
    126: op1_15_in20 = reg_0140;
    127: op1_15_in20 = reg_1204;
    128: op1_15_in20 = reg_0978;
    129: op1_15_in20 = reg_1403;
    130: op1_15_in20 = reg_1040;
    default: op1_15_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の20番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv20 = 1;
    73: op1_15_inv20 = 1;
    86: op1_15_inv20 = 1;
    54: op1_15_inv20 = 1;
    75: op1_15_inv20 = 1;
    69: op1_15_inv20 = 1;
    56: op1_15_inv20 = 1;
    57: op1_15_inv20 = 1;
    78: op1_15_inv20 = 1;
    59: op1_15_inv20 = 1;
    79: op1_15_inv20 = 1;
    60: op1_15_inv20 = 1;
    88: op1_15_inv20 = 1;
    80: op1_15_inv20 = 1;
    62: op1_15_inv20 = 1;
    82: op1_15_inv20 = 1;
    63: op1_15_inv20 = 1;
    52: op1_15_inv20 = 1;
    89: op1_15_inv20 = 1;
    84: op1_15_inv20 = 1;
    85: op1_15_inv20 = 1;
    48: op1_15_inv20 = 1;
    92: op1_15_inv20 = 1;
    95: op1_15_inv20 = 1;
    96: op1_15_inv20 = 1;
    97: op1_15_inv20 = 1;
    98: op1_15_inv20 = 1;
    101: op1_15_inv20 = 1;
    102: op1_15_inv20 = 1;
    104: op1_15_inv20 = 1;
    105: op1_15_inv20 = 1;
    106: op1_15_inv20 = 1;
    107: op1_15_inv20 = 1;
    112: op1_15_inv20 = 1;
    115: op1_15_inv20 = 1;
    116: op1_15_inv20 = 1;
    117: op1_15_inv20 = 1;
    119: op1_15_inv20 = 1;
    121: op1_15_inv20 = 1;
    122: op1_15_inv20 = 1;
    124: op1_15_inv20 = 1;
    127: op1_15_inv20 = 1;
    128: op1_15_inv20 = 1;
    129: op1_15_inv20 = 1;
    default: op1_15_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の21番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in21 = reg_0057;
    73: op1_15_in21 = reg_0906;
    53: op1_15_in21 = reg_0788;
    86: op1_15_in21 = reg_0462;
    128: op1_15_in21 = reg_0462;
    74: op1_15_in21 = reg_1032;
    54: op1_15_in21 = reg_0105;
    75: op1_15_in21 = reg_0015;
    69: op1_15_in21 = reg_0677;
    56: op1_15_in21 = reg_1139;
    49: op1_15_in21 = reg_0521;
    76: op1_15_in21 = reg_0411;
    87: op1_15_in21 = reg_1041;
    57: op1_15_in21 = reg_0456;
    50: op1_15_in21 = reg_0525;
    68: op1_15_in21 = reg_0392;
    71: op1_15_in21 = reg_0609;
    77: op1_15_in21 = reg_1183;
    78: op1_15_in21 = reg_1179;
    61: op1_15_in21 = reg_0576;
    58: op1_15_in21 = reg_0176;
    70: op1_15_in21 = reg_0341;
    59: op1_15_in21 = reg_0878;
    79: op1_15_in21 = reg_0073;
    51: op1_15_in21 = reg_0217;
    88: op1_15_in21 = reg_0131;
    80: op1_15_in21 = reg_0271;
    62: op1_15_in21 = reg_0211;
    81: op1_15_in21 = reg_1433;
    82: op1_15_in21 = reg_0458;
    63: op1_15_in21 = reg_0549;
    52: op1_15_in21 = reg_0851;
    47: op1_15_in21 = reg_0851;
    83: op1_15_in21 = reg_1495;
    89: op1_15_in21 = reg_0450;
    100: op1_15_in21 = reg_0450;
    84: op1_15_in21 = reg_0723;
    85: op1_15_in21 = reg_0182;
    65: op1_15_in21 = reg_0218;
    90: op1_15_in21 = reg_0522;
    91: op1_15_in21 = reg_0016;
    46: op1_15_in21 = reg_0783;
    48: op1_15_in21 = reg_0138;
    67: op1_15_in21 = reg_1152;
    92: op1_15_in21 = reg_0007;
    93: op1_15_in21 = reg_1095;
    94: op1_15_in21 = reg_0880;
    95: op1_15_in21 = reg_0163;
    96: op1_15_in21 = reg_0238;
    97: op1_15_in21 = reg_0960;
    98: op1_15_in21 = reg_1369;
    101: op1_15_in21 = reg_0726;
    102: op1_15_in21 = reg_0932;
    103: op1_15_in21 = reg_0115;
    104: op1_15_in21 = reg_0468;
    105: op1_15_in21 = reg_0787;
    106: op1_15_in21 = reg_1207;
    107: op1_15_in21 = reg_0471;
    108: op1_15_in21 = reg_0439;
    109: op1_15_in21 = reg_0568;
    110: op1_15_in21 = reg_0706;
    112: op1_15_in21 = reg_1231;
    113: op1_15_in21 = reg_0819;
    114: op1_15_in21 = reg_0334;
    115: op1_15_in21 = reg_0441;
    116: op1_15_in21 = reg_0395;
    117: op1_15_in21 = reg_0478;
    118: op1_15_in21 = reg_0437;
    119: op1_15_in21 = reg_0331;
    120: op1_15_in21 = reg_0999;
    121: op1_15_in21 = reg_0096;
    122: op1_15_in21 = reg_0989;
    123: op1_15_in21 = reg_1324;
    124: op1_15_in21 = reg_1204;
    125: op1_15_in21 = reg_0820;
    126: op1_15_in21 = reg_0309;
    127: op1_15_in21 = reg_0371;
    129: op1_15_in21 = reg_0792;
    130: op1_15_in21 = reg_1065;
    default: op1_15_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の21番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_15_inv21 = 1;
    86: op1_15_inv21 = 1;
    74: op1_15_inv21 = 1;
    54: op1_15_inv21 = 1;
    76: op1_15_inv21 = 1;
    87: op1_15_inv21 = 1;
    57: op1_15_inv21 = 1;
    68: op1_15_inv21 = 1;
    78: op1_15_inv21 = 1;
    61: op1_15_inv21 = 1;
    58: op1_15_inv21 = 1;
    59: op1_15_inv21 = 1;
    79: op1_15_inv21 = 1;
    51: op1_15_inv21 = 1;
    88: op1_15_inv21 = 1;
    62: op1_15_inv21 = 1;
    82: op1_15_inv21 = 1;
    52: op1_15_inv21 = 1;
    83: op1_15_inv21 = 1;
    89: op1_15_inv21 = 1;
    85: op1_15_inv21 = 1;
    65: op1_15_inv21 = 1;
    92: op1_15_inv21 = 1;
    96: op1_15_inv21 = 1;
    98: op1_15_inv21 = 1;
    100: op1_15_inv21 = 1;
    101: op1_15_inv21 = 1;
    102: op1_15_inv21 = 1;
    104: op1_15_inv21 = 1;
    105: op1_15_inv21 = 1;
    106: op1_15_inv21 = 1;
    110: op1_15_inv21 = 1;
    114: op1_15_inv21 = 1;
    47: op1_15_inv21 = 1;
    127: op1_15_inv21 = 1;
    128: op1_15_inv21 = 1;
    129: op1_15_inv21 = 1;
    default: op1_15_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の22番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in22 = reg_1100;
    73: op1_15_in22 = reg_0905;
    53: op1_15_in22 = reg_0787;
    86: op1_15_in22 = reg_0531;
    74: op1_15_in22 = reg_0728;
    54: op1_15_in22 = reg_0897;
    75: op1_15_in22 = reg_0962;
    69: op1_15_in22 = reg_0216;
    56: op1_15_in22 = reg_0497;
    76: op1_15_in22 = reg_1372;
    87: op1_15_in22 = reg_0199;
    57: op1_15_in22 = reg_0563;
    50: op1_15_in22 = reg_0707;
    68: op1_15_in22 = reg_0646;
    71: op1_15_in22 = imem01_in[3:0];
    77: op1_15_in22 = reg_0186;
    47: op1_15_in22 = reg_0186;
    78: op1_15_in22 = reg_0023;
    80: op1_15_in22 = reg_0023;
    61: op1_15_in22 = reg_0984;
    58: op1_15_in22 = reg_0346;
    70: op1_15_in22 = reg_0181;
    59: op1_15_in22 = reg_0848;
    79: op1_15_in22 = reg_1321;
    51: op1_15_in22 = reg_0280;
    88: op1_15_in22 = reg_0334;
    62: op1_15_in22 = reg_0035;
    81: op1_15_in22 = reg_0876;
    82: op1_15_in22 = reg_0466;
    63: op1_15_in22 = reg_0982;
    52: op1_15_in22 = reg_0921;
    83: op1_15_in22 = reg_0288;
    89: op1_15_in22 = reg_0418;
    84: op1_15_in22 = reg_1512;
    85: op1_15_in22 = reg_0564;
    65: op1_15_in22 = reg_0235;
    90: op1_15_in22 = reg_0419;
    91: op1_15_in22 = reg_1488;
    46: op1_15_in22 = reg_0192;
    48: op1_15_in22 = reg_0008;
    67: op1_15_in22 = reg_0553;
    92: op1_15_in22 = imem03_in[3:0];
    120: op1_15_in22 = imem03_in[3:0];
    93: op1_15_in22 = reg_0394;
    94: op1_15_in22 = reg_0448;
    95: op1_15_in22 = reg_0550;
    96: op1_15_in22 = reg_0241;
    97: op1_15_in22 = reg_0782;
    98: op1_15_in22 = reg_0034;
    100: op1_15_in22 = reg_0318;
    101: op1_15_in22 = reg_0146;
    102: op1_15_in22 = reg_0633;
    103: op1_15_in22 = reg_0109;
    104: op1_15_in22 = reg_0149;
    105: op1_15_in22 = reg_0238;
    106: op1_15_in22 = reg_0432;
    107: op1_15_in22 = reg_0537;
    108: op1_15_in22 = reg_0148;
    109: op1_15_in22 = reg_0571;
    110: op1_15_in22 = reg_0999;
    112: op1_15_in22 = reg_0107;
    113: op1_15_in22 = reg_0868;
    114: op1_15_in22 = reg_1180;
    115: op1_15_in22 = reg_0404;
    116: op1_15_in22 = reg_0831;
    117: op1_15_in22 = reg_1060;
    118: op1_15_in22 = reg_0740;
    119: op1_15_in22 = reg_1474;
    125: op1_15_in22 = reg_1474;
    121: op1_15_in22 = reg_0210;
    122: op1_15_in22 = reg_0732;
    123: op1_15_in22 = reg_0723;
    124: op1_15_in22 = reg_0754;
    126: op1_15_in22 = reg_1350;
    127: op1_15_in22 = reg_0067;
    128: op1_15_in22 = reg_1200;
    129: op1_15_in22 = reg_1163;
    130: op1_15_in22 = reg_0451;
    default: op1_15_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の22番目の入力反転
  always @ ( * ) begin
    case ( state )
    53: op1_15_inv22 = 1;
    74: op1_15_inv22 = 1;
    54: op1_15_inv22 = 1;
    69: op1_15_inv22 = 1;
    76: op1_15_inv22 = 1;
    87: op1_15_inv22 = 1;
    57: op1_15_inv22 = 1;
    61: op1_15_inv22 = 1;
    58: op1_15_inv22 = 1;
    70: op1_15_inv22 = 1;
    51: op1_15_inv22 = 1;
    88: op1_15_inv22 = 1;
    62: op1_15_inv22 = 1;
    81: op1_15_inv22 = 1;
    82: op1_15_inv22 = 1;
    52: op1_15_inv22 = 1;
    89: op1_15_inv22 = 1;
    65: op1_15_inv22 = 1;
    91: op1_15_inv22 = 1;
    94: op1_15_inv22 = 1;
    96: op1_15_inv22 = 1;
    100: op1_15_inv22 = 1;
    101: op1_15_inv22 = 1;
    103: op1_15_inv22 = 1;
    104: op1_15_inv22 = 1;
    105: op1_15_inv22 = 1;
    107: op1_15_inv22 = 1;
    109: op1_15_inv22 = 1;
    110: op1_15_inv22 = 1;
    112: op1_15_inv22 = 1;
    114: op1_15_inv22 = 1;
    115: op1_15_inv22 = 1;
    47: op1_15_inv22 = 1;
    121: op1_15_inv22 = 1;
    123: op1_15_inv22 = 1;
    126: op1_15_inv22 = 1;
    127: op1_15_inv22 = 1;
    130: op1_15_inv22 = 1;
    default: op1_15_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の23番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in23 = reg_0372;
    73: op1_15_in23 = reg_1326;
    53: op1_15_in23 = reg_0547;
    86: op1_15_in23 = reg_0500;
    74: op1_15_in23 = imem01_in[7:4];
    71: op1_15_in23 = imem01_in[7:4];
    54: op1_15_in23 = reg_0306;
    75: op1_15_in23 = reg_0324;
    69: op1_15_in23 = reg_1064;
    56: op1_15_in23 = imem02_in[11:8];
    76: op1_15_in23 = reg_0181;
    87: op1_15_in23 = reg_1077;
    57: op1_15_in23 = reg_0530;
    50: op1_15_in23 = reg_0180;
    68: op1_15_in23 = reg_0131;
    77: op1_15_in23 = reg_0894;
    78: op1_15_in23 = reg_0152;
    61: op1_15_in23 = reg_0743;
    58: op1_15_in23 = reg_0648;
    70: op1_15_in23 = reg_1367;
    59: op1_15_in23 = reg_0154;
    120: op1_15_in23 = reg_0154;
    79: op1_15_in23 = reg_0005;
    51: op1_15_in23 = reg_0121;
    88: op1_15_in23 = reg_0697;
    80: op1_15_in23 = reg_0046;
    62: op1_15_in23 = reg_0794;
    81: op1_15_in23 = reg_0712;
    82: op1_15_in23 = reg_0120;
    63: op1_15_in23 = reg_0363;
    52: op1_15_in23 = reg_0924;
    83: op1_15_in23 = imem03_in[11:8];
    89: op1_15_in23 = reg_0873;
    84: op1_15_in23 = reg_0093;
    85: op1_15_in23 = reg_0938;
    65: op1_15_in23 = imem03_in[3:0];
    90: op1_15_in23 = reg_0119;
    91: op1_15_in23 = reg_0210;
    102: op1_15_in23 = reg_0210;
    46: op1_15_in23 = reg_0925;
    48: op1_15_in23 = reg_0279;
    67: op1_15_in23 = reg_0982;
    92: op1_15_in23 = reg_0840;
    93: op1_15_in23 = reg_1183;
    94: op1_15_in23 = reg_1282;
    95: op1_15_in23 = reg_0609;
    96: op1_15_in23 = reg_0572;
    97: op1_15_in23 = reg_0717;
    98: op1_15_in23 = reg_1258;
    100: op1_15_in23 = reg_0828;
    101: op1_15_in23 = reg_1513;
    103: op1_15_in23 = reg_0636;
    104: op1_15_in23 = reg_1511;
    113: op1_15_in23 = reg_1511;
    105: op1_15_in23 = reg_0612;
    106: op1_15_in23 = reg_0436;
    107: op1_15_in23 = reg_1040;
    108: op1_15_in23 = reg_0146;
    109: op1_15_in23 = reg_0323;
    110: op1_15_in23 = reg_0216;
    112: op1_15_in23 = reg_0882;
    114: op1_15_in23 = reg_1404;
    115: op1_15_in23 = reg_0620;
    116: op1_15_in23 = reg_0392;
    117: op1_15_in23 = reg_0892;
    118: op1_15_in23 = reg_0404;
    119: op1_15_in23 = reg_0819;
    47: op1_15_in23 = reg_0139;
    121: op1_15_in23 = reg_0278;
    122: op1_15_in23 = reg_0179;
    123: op1_15_in23 = reg_0383;
    124: op1_15_in23 = reg_0195;
    125: op1_15_in23 = reg_0439;
    126: op1_15_in23 = reg_0156;
    127: op1_15_in23 = reg_0498;
    128: op1_15_in23 = reg_0796;
    129: op1_15_in23 = reg_0418;
    130: op1_15_in23 = reg_0097;
    default: op1_15_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の23番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_15_inv23 = 1;
    54: op1_15_inv23 = 1;
    69: op1_15_inv23 = 1;
    56: op1_15_inv23 = 1;
    76: op1_15_inv23 = 1;
    87: op1_15_inv23 = 1;
    78: op1_15_inv23 = 1;
    70: op1_15_inv23 = 1;
    59: op1_15_inv23 = 1;
    79: op1_15_inv23 = 1;
    62: op1_15_inv23 = 1;
    81: op1_15_inv23 = 1;
    63: op1_15_inv23 = 1;
    85: op1_15_inv23 = 1;
    67: op1_15_inv23 = 1;
    92: op1_15_inv23 = 1;
    94: op1_15_inv23 = 1;
    95: op1_15_inv23 = 1;
    98: op1_15_inv23 = 1;
    101: op1_15_inv23 = 1;
    102: op1_15_inv23 = 1;
    104: op1_15_inv23 = 1;
    107: op1_15_inv23 = 1;
    110: op1_15_inv23 = 1;
    112: op1_15_inv23 = 1;
    113: op1_15_inv23 = 1;
    114: op1_15_inv23 = 1;
    116: op1_15_inv23 = 1;
    47: op1_15_inv23 = 1;
    120: op1_15_inv23 = 1;
    122: op1_15_inv23 = 1;
    123: op1_15_inv23 = 1;
    125: op1_15_inv23 = 1;
    126: op1_15_inv23 = 1;
    127: op1_15_inv23 = 1;
    130: op1_15_inv23 = 1;
    default: op1_15_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の24番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in24 = reg_0788;
    123: op1_15_in24 = reg_0788;
    73: op1_15_in24 = reg_0860;
    53: op1_15_in24 = reg_0548;
    86: op1_15_in24 = reg_1147;
    128: op1_15_in24 = reg_1147;
    74: op1_15_in24 = reg_0239;
    54: op1_15_in24 = reg_0154;
    75: op1_15_in24 = imem07_in[15:12];
    69: op1_15_in24 = reg_1149;
    56: op1_15_in24 = reg_0970;
    76: op1_15_in24 = reg_1368;
    87: op1_15_in24 = reg_1004;
    57: op1_15_in24 = reg_1140;
    50: op1_15_in24 = reg_0178;
    68: op1_15_in24 = reg_0567;
    71: op1_15_in24 = imem01_in[15:12];
    77: op1_15_in24 = reg_0135;
    117: op1_15_in24 = reg_0135;
    78: op1_15_in24 = reg_0015;
    61: op1_15_in24 = reg_1151;
    58: op1_15_in24 = reg_0131;
    70: op1_15_in24 = reg_1257;
    59: op1_15_in24 = reg_0279;
    79: op1_15_in24 = reg_0917;
    51: op1_15_in24 = reg_0198;
    88: op1_15_in24 = reg_1401;
    80: op1_15_in24 = reg_0560;
    62: op1_15_in24 = reg_0393;
    81: op1_15_in24 = reg_0307;
    82: op1_15_in24 = reg_1209;
    63: op1_15_in24 = reg_0724;
    52: op1_15_in24 = reg_0465;
    83: op1_15_in24 = reg_0216;
    89: op1_15_in24 = reg_1484;
    84: op1_15_in24 = reg_0550;
    85: op1_15_in24 = reg_0090;
    65: op1_15_in24 = reg_1139;
    90: op1_15_in24 = reg_0165;
    91: op1_15_in24 = reg_0266;
    46: op1_15_in24 = reg_0161;
    48: op1_15_in24 = reg_0314;
    67: op1_15_in24 = reg_0572;
    105: op1_15_in24 = reg_0572;
    92: op1_15_in24 = reg_0999;
    93: op1_15_in24 = reg_0868;
    94: op1_15_in24 = reg_0426;
    95: op1_15_in24 = reg_0242;
    96: op1_15_in24 = reg_0147;
    97: op1_15_in24 = reg_0373;
    98: op1_15_in24 = reg_0574;
    100: op1_15_in24 = imem06_in[3:0];
    101: op1_15_in24 = reg_0092;
    102: op1_15_in24 = reg_1430;
    103: op1_15_in24 = reg_0529;
    104: op1_15_in24 = reg_0386;
    106: op1_15_in24 = reg_0776;
    107: op1_15_in24 = reg_1077;
    108: op1_15_in24 = reg_0400;
    109: op1_15_in24 = reg_0295;
    110: op1_15_in24 = reg_1033;
    122: op1_15_in24 = reg_1033;
    112: op1_15_in24 = reg_0880;
    113: op1_15_in24 = reg_0875;
    114: op1_15_in24 = reg_0477;
    115: op1_15_in24 = reg_0361;
    116: op1_15_in24 = reg_0391;
    118: op1_15_in24 = reg_0415;
    119: op1_15_in24 = reg_0430;
    47: op1_15_in24 = reg_0774;
    120: op1_15_in24 = reg_1000;
    121: op1_15_in24 = reg_0315;
    124: op1_15_in24 = reg_0215;
    125: op1_15_in24 = reg_1456;
    126: op1_15_in24 = reg_0775;
    127: op1_15_in24 = reg_1010;
    129: op1_15_in24 = reg_0130;
    130: op1_15_in24 = reg_0487;
    default: op1_15_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の24番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv24 = 1;
    73: op1_15_inv24 = 1;
    86: op1_15_inv24 = 1;
    69: op1_15_inv24 = 1;
    68: op1_15_inv24 = 1;
    71: op1_15_inv24 = 1;
    78: op1_15_inv24 = 1;
    61: op1_15_inv24 = 1;
    70: op1_15_inv24 = 1;
    59: op1_15_inv24 = 1;
    80: op1_15_inv24 = 1;
    62: op1_15_inv24 = 1;
    81: op1_15_inv24 = 1;
    63: op1_15_inv24 = 1;
    52: op1_15_inv24 = 1;
    83: op1_15_inv24 = 1;
    65: op1_15_inv24 = 1;
    46: op1_15_inv24 = 1;
    48: op1_15_inv24 = 1;
    67: op1_15_inv24 = 1;
    92: op1_15_inv24 = 1;
    94: op1_15_inv24 = 1;
    97: op1_15_inv24 = 1;
    98: op1_15_inv24 = 1;
    101: op1_15_inv24 = 1;
    102: op1_15_inv24 = 1;
    105: op1_15_inv24 = 1;
    108: op1_15_inv24 = 1;
    109: op1_15_inv24 = 1;
    110: op1_15_inv24 = 1;
    112: op1_15_inv24 = 1;
    113: op1_15_inv24 = 1;
    114: op1_15_inv24 = 1;
    119: op1_15_inv24 = 1;
    47: op1_15_inv24 = 1;
    120: op1_15_inv24 = 1;
    122: op1_15_inv24 = 1;
    123: op1_15_inv24 = 1;
    126: op1_15_inv24 = 1;
    128: op1_15_inv24 = 1;
    default: op1_15_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の25番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in25 = reg_1291;
    73: op1_15_in25 = reg_0115;
    53: op1_15_in25 = reg_0166;
    86: op1_15_in25 = reg_0969;
    74: op1_15_in25 = reg_0819;
    54: op1_15_in25 = reg_0830;
    75: op1_15_in25 = reg_0667;
    69: op1_15_in25 = reg_0177;
    56: op1_15_in25 = reg_0626;
    76: op1_15_in25 = reg_1257;
    87: op1_15_in25 = reg_0452;
    57: op1_15_in25 = reg_1139;
    50: op1_15_in25 = reg_0999;
    68: op1_15_in25 = reg_0564;
    71: op1_15_in25 = reg_0439;
    77: op1_15_in25 = reg_0674;
    78: op1_15_in25 = imem07_in[7:4];
    61: op1_15_in25 = reg_0930;
    67: op1_15_in25 = reg_0930;
    58: op1_15_in25 = reg_0567;
    70: op1_15_in25 = reg_1258;
    59: op1_15_in25 = reg_0276;
    79: op1_15_in25 = reg_1100;
    51: op1_15_in25 = reg_0710;
    88: op1_15_in25 = reg_1070;
    80: op1_15_in25 = imem07_in[15:12];
    62: op1_15_in25 = reg_0736;
    81: op1_15_in25 = reg_0531;
    82: op1_15_in25 = reg_0869;
    63: op1_15_in25 = reg_0282;
    52: op1_15_in25 = reg_0286;
    83: op1_15_in25 = reg_0198;
    89: op1_15_in25 = reg_0197;
    84: op1_15_in25 = reg_0548;
    85: op1_15_in25 = reg_1486;
    65: op1_15_in25 = reg_0145;
    90: op1_15_in25 = reg_1202;
    91: op1_15_in25 = reg_0367;
    46: op1_15_in25 = reg_0906;
    48: op1_15_in25 = reg_0677;
    92: op1_15_in25 = reg_0261;
    93: op1_15_in25 = reg_1440;
    94: op1_15_in25 = reg_1146;
    95: op1_15_in25 = reg_0239;
    96: op1_15_in25 = reg_0149;
    125: op1_15_in25 = reg_0149;
    97: op1_15_in25 = reg_0622;
    98: op1_15_in25 = reg_0681;
    100: op1_15_in25 = reg_1064;
    101: op1_15_in25 = reg_0464;
    102: op1_15_in25 = reg_0136;
    103: op1_15_in25 = reg_0345;
    104: op1_15_in25 = reg_0595;
    105: op1_15_in25 = reg_1511;
    106: op1_15_in25 = reg_0778;
    107: op1_15_in25 = reg_0320;
    108: op1_15_in25 = reg_0896;
    109: op1_15_in25 = reg_0152;
    110: op1_15_in25 = reg_0311;
    112: op1_15_in25 = reg_1009;
    113: op1_15_in25 = reg_0400;
    114: op1_15_in25 = reg_0937;
    115: op1_15_in25 = reg_0519;
    116: op1_15_in25 = reg_0303;
    117: op1_15_in25 = reg_0703;
    118: op1_15_in25 = reg_0413;
    119: op1_15_in25 = reg_1452;
    47: op1_15_in25 = reg_0739;
    120: op1_15_in25 = reg_0216;
    121: op1_15_in25 = imem05_in[3:0];
    122: op1_15_in25 = reg_1001;
    123: op1_15_in25 = reg_1254;
    124: op1_15_in25 = reg_0018;
    126: op1_15_in25 = reg_0285;
    127: op1_15_in25 = reg_0922;
    128: op1_15_in25 = reg_1041;
    129: op1_15_in25 = reg_0602;
    130: op1_15_in25 = reg_1340;
    default: op1_15_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の25番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv25 = 1;
    73: op1_15_inv25 = 1;
    86: op1_15_inv25 = 1;
    74: op1_15_inv25 = 1;
    75: op1_15_inv25 = 1;
    56: op1_15_inv25 = 1;
    57: op1_15_inv25 = 1;
    61: op1_15_inv25 = 1;
    59: op1_15_inv25 = 1;
    79: op1_15_inv25 = 1;
    51: op1_15_inv25 = 1;
    88: op1_15_inv25 = 1;
    80: op1_15_inv25 = 1;
    62: op1_15_inv25 = 1;
    63: op1_15_inv25 = 1;
    52: op1_15_inv25 = 1;
    89: op1_15_inv25 = 1;
    84: op1_15_inv25 = 1;
    85: op1_15_inv25 = 1;
    90: op1_15_inv25 = 1;
    91: op1_15_inv25 = 1;
    46: op1_15_inv25 = 1;
    67: op1_15_inv25 = 1;
    92: op1_15_inv25 = 1;
    95: op1_15_inv25 = 1;
    101: op1_15_inv25 = 1;
    102: op1_15_inv25 = 1;
    103: op1_15_inv25 = 1;
    105: op1_15_inv25 = 1;
    108: op1_15_inv25 = 1;
    112: op1_15_inv25 = 1;
    113: op1_15_inv25 = 1;
    116: op1_15_inv25 = 1;
    47: op1_15_inv25 = 1;
    120: op1_15_inv25 = 1;
    121: op1_15_inv25 = 1;
    124: op1_15_inv25 = 1;
    125: op1_15_inv25 = 1;
    126: op1_15_inv25 = 1;
    128: op1_15_inv25 = 1;
    129: op1_15_inv25 = 1;
    default: op1_15_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の26番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in26 = reg_1068;
    73: op1_15_in26 = reg_0637;
    53: op1_15_in26 = reg_0242;
    86: op1_15_in26 = reg_0599;
    74: op1_15_in26 = reg_0438;
    54: op1_15_in26 = reg_0325;
    75: op1_15_in26 = reg_0309;
    69: op1_15_in26 = imem03_in[7:4];
    56: op1_15_in26 = reg_0128;
    76: op1_15_in26 = reg_1216;
    87: op1_15_in26 = reg_0061;
    107: op1_15_in26 = reg_0061;
    57: op1_15_in26 = reg_0474;
    50: op1_15_in26 = reg_0142;
    68: op1_15_in26 = reg_0275;
    71: op1_15_in26 = reg_0430;
    77: op1_15_in26 = reg_0187;
    78: op1_15_in26 = imem07_in[11:8];
    61: op1_15_in26 = reg_0403;
    58: op1_15_in26 = reg_0566;
    70: op1_15_in26 = reg_1203;
    59: op1_15_in26 = reg_1132;
    79: op1_15_in26 = imem01_in[3:0];
    51: op1_15_in26 = reg_0444;
    88: op1_15_in26 = reg_0450;
    80: op1_15_in26 = reg_0391;
    62: op1_15_in26 = reg_0273;
    81: op1_15_in26 = reg_0800;
    82: op1_15_in26 = reg_0752;
    63: op1_15_in26 = reg_0012;
    52: op1_15_in26 = reg_0740;
    83: op1_15_in26 = reg_0143;
    65: op1_15_in26 = reg_0143;
    89: op1_15_in26 = reg_0274;
    84: op1_15_in26 = reg_0746;
    85: op1_15_in26 = reg_0601;
    90: op1_15_in26 = reg_0023;
    91: op1_15_in26 = reg_0833;
    46: op1_15_in26 = imem06_in[7:4];
    48: op1_15_in26 = reg_0630;
    67: op1_15_in26 = reg_0149;
    92: op1_15_in26 = reg_0216;
    93: op1_15_in26 = reg_0703;
    127: op1_15_in26 = reg_0703;
    94: op1_15_in26 = reg_0237;
    95: op1_15_in26 = reg_0572;
    96: op1_15_in26 = reg_0360;
    97: op1_15_in26 = reg_0527;
    98: op1_15_in26 = reg_0094;
    100: op1_15_in26 = reg_0908;
    101: op1_15_in26 = reg_0400;
    102: op1_15_in26 = reg_0702;
    121: op1_15_in26 = reg_0702;
    103: op1_15_in26 = reg_0979;
    104: op1_15_in26 = reg_0724;
    105: op1_15_in26 = reg_0384;
    106: op1_15_in26 = reg_1433;
    108: op1_15_in26 = imem02_in[3:0];
    109: op1_15_in26 = imem07_in[3:0];
    110: op1_15_in26 = reg_0891;
    112: op1_15_in26 = reg_0313;
    113: op1_15_in26 = reg_0078;
    114: op1_15_in26 = reg_0873;
    115: op1_15_in26 = reg_0518;
    116: op1_15_in26 = reg_0240;
    117: op1_15_in26 = reg_0170;
    118: op1_15_in26 = reg_0102;
    119: op1_15_in26 = reg_1456;
    47: op1_15_in26 = reg_0404;
    120: op1_15_in26 = reg_0600;
    122: op1_15_in26 = reg_0600;
    123: op1_15_in26 = reg_0874;
    124: op1_15_in26 = reg_0022;
    125: op1_15_in26 = reg_1032;
    126: op1_15_in26 = reg_0437;
    128: op1_15_in26 = reg_1065;
    129: op1_15_in26 = reg_0589;
    130: op1_15_in26 = reg_1237;
    default: op1_15_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の26番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv26 = 1;
    73: op1_15_inv26 = 1;
    53: op1_15_inv26 = 1;
    54: op1_15_inv26 = 1;
    76: op1_15_inv26 = 1;
    68: op1_15_inv26 = 1;
    71: op1_15_inv26 = 1;
    77: op1_15_inv26 = 1;
    78: op1_15_inv26 = 1;
    70: op1_15_inv26 = 1;
    79: op1_15_inv26 = 1;
    51: op1_15_inv26 = 1;
    82: op1_15_inv26 = 1;
    63: op1_15_inv26 = 1;
    83: op1_15_inv26 = 1;
    89: op1_15_inv26 = 1;
    84: op1_15_inv26 = 1;
    65: op1_15_inv26 = 1;
    91: op1_15_inv26 = 1;
    48: op1_15_inv26 = 1;
    67: op1_15_inv26 = 1;
    95: op1_15_inv26 = 1;
    96: op1_15_inv26 = 1;
    98: op1_15_inv26 = 1;
    100: op1_15_inv26 = 1;
    103: op1_15_inv26 = 1;
    107: op1_15_inv26 = 1;
    108: op1_15_inv26 = 1;
    109: op1_15_inv26 = 1;
    114: op1_15_inv26 = 1;
    117: op1_15_inv26 = 1;
    47: op1_15_inv26 = 1;
    123: op1_15_inv26 = 1;
    124: op1_15_inv26 = 1;
    125: op1_15_inv26 = 1;
    127: op1_15_inv26 = 1;
    128: op1_15_inv26 = 1;
    129: op1_15_inv26 = 1;
    default: op1_15_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の27番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in27 = reg_0550;
    73: op1_15_in27 = reg_0622;
    53: op1_15_in27 = reg_0239;
    86: op1_15_in27 = reg_1065;
    74: op1_15_in27 = reg_0383;
    54: op1_15_in27 = reg_0279;
    75: op1_15_in27 = reg_0157;
    69: op1_15_in27 = reg_1139;
    56: op1_15_in27 = reg_0112;
    76: op1_15_in27 = reg_1198;
    70: op1_15_in27 = reg_1198;
    87: op1_15_in27 = reg_0836;
    57: op1_15_in27 = reg_0429;
    50: op1_15_in27 = reg_0246;
    68: op1_15_in27 = reg_1373;
    71: op1_15_in27 = reg_0149;
    77: op1_15_in27 = reg_0297;
    94: op1_15_in27 = reg_0297;
    78: op1_15_in27 = reg_0198;
    61: op1_15_in27 = reg_0047;
    58: op1_15_in27 = reg_1181;
    59: op1_15_in27 = reg_0755;
    79: op1_15_in27 = reg_0448;
    51: op1_15_in27 = reg_0698;
    88: op1_15_in27 = reg_0302;
    80: op1_15_in27 = reg_0491;
    62: op1_15_in27 = reg_0833;
    81: op1_15_in27 = reg_1515;
    82: op1_15_in27 = reg_1505;
    63: op1_15_in27 = reg_0530;
    52: op1_15_in27 = reg_0408;
    83: op1_15_in27 = reg_0964;
    89: op1_15_in27 = reg_0118;
    84: op1_15_in27 = reg_0820;
    85: op1_15_in27 = reg_0240;
    65: op1_15_in27 = reg_0559;
    90: op1_15_in27 = reg_0046;
    91: op1_15_in27 = reg_0702;
    46: op1_15_in27 = reg_0860;
    48: op1_15_in27 = reg_0444;
    67: op1_15_in27 = reg_0148;
    119: op1_15_in27 = reg_0148;
    92: op1_15_in27 = reg_1001;
    93: op1_15_in27 = reg_0309;
    95: op1_15_in27 = reg_1457;
    96: op1_15_in27 = reg_0875;
    97: op1_15_in27 = reg_0568;
    98: op1_15_in27 = reg_1040;
    100: op1_15_in27 = reg_0316;
    101: op1_15_in27 = reg_1071;
    102: op1_15_in27 = reg_0346;
    103: op1_15_in27 = reg_0119;
    104: op1_15_in27 = reg_0403;
    105: op1_15_in27 = reg_0385;
    106: op1_15_in27 = reg_1140;
    107: op1_15_in27 = reg_0487;
    108: op1_15_in27 = imem02_in[7:4];
    109: op1_15_in27 = imem07_in[11:8];
    110: op1_15_in27 = reg_0556;
    112: op1_15_in27 = reg_1325;
    113: op1_15_in27 = reg_0257;
    114: op1_15_in27 = reg_0492;
    115: op1_15_in27 = reg_0483;
    116: op1_15_in27 = reg_1348;
    117: op1_15_in27 = reg_0457;
    118: op1_15_in27 = reg_0321;
    47: op1_15_in27 = reg_0415;
    120: op1_15_in27 = reg_0891;
    121: op1_15_in27 = reg_1164;
    122: op1_15_in27 = reg_0143;
    123: op1_15_in27 = reg_0576;
    124: op1_15_in27 = reg_0017;
    125: op1_15_in27 = reg_1511;
    126: op1_15_in27 = reg_0620;
    127: op1_15_in27 = reg_0225;
    128: op1_15_in27 = reg_0835;
    129: op1_15_in27 = reg_0014;
    130: op1_15_in27 = reg_0117;
    default: op1_15_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の27番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv27 = 1;
    53: op1_15_inv27 = 1;
    87: op1_15_inv27 = 1;
    57: op1_15_inv27 = 1;
    50: op1_15_inv27 = 1;
    68: op1_15_inv27 = 1;
    71: op1_15_inv27 = 1;
    77: op1_15_inv27 = 1;
    78: op1_15_inv27 = 1;
    61: op1_15_inv27 = 1;
    79: op1_15_inv27 = 1;
    51: op1_15_inv27 = 1;
    88: op1_15_inv27 = 1;
    62: op1_15_inv27 = 1;
    82: op1_15_inv27 = 1;
    90: op1_15_inv27 = 1;
    92: op1_15_inv27 = 1;
    93: op1_15_inv27 = 1;
    97: op1_15_inv27 = 1;
    98: op1_15_inv27 = 1;
    102: op1_15_inv27 = 1;
    104: op1_15_inv27 = 1;
    106: op1_15_inv27 = 1;
    107: op1_15_inv27 = 1;
    108: op1_15_inv27 = 1;
    112: op1_15_inv27 = 1;
    113: op1_15_inv27 = 1;
    118: op1_15_inv27 = 1;
    47: op1_15_inv27 = 1;
    121: op1_15_inv27 = 1;
    125: op1_15_inv27 = 1;
    128: op1_15_inv27 = 1;
    default: op1_15_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の28番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in28 = reg_0747;
    73: op1_15_in28 = reg_0323;
    53: op1_15_in28 = reg_0746;
    86: op1_15_in28 = reg_0320;
    98: op1_15_in28 = reg_0320;
    74: op1_15_in28 = reg_0360;
    54: op1_15_in28 = reg_0312;
    75: op1_15_in28 = reg_0924;
    69: op1_15_in28 = reg_0144;
    56: op1_15_in28 = reg_0105;
    76: op1_15_in28 = reg_1147;
    87: op1_15_in28 = reg_0117;
    57: op1_15_in28 = reg_0436;
    50: op1_15_in28 = reg_0891;
    68: op1_15_in28 = reg_0274;
    71: op1_15_in28 = reg_0400;
    125: op1_15_in28 = reg_0400;
    77: op1_15_in28 = reg_1347;
    78: op1_15_in28 = reg_1056;
    61: op1_15_in28 = reg_0724;
    58: op1_15_in28 = reg_0316;
    70: op1_15_in28 = reg_0412;
    59: op1_15_in28 = reg_0525;
    79: op1_15_in28 = reg_1254;
    51: op1_15_in28 = reg_0178;
    88: op1_15_in28 = reg_0275;
    80: op1_15_in28 = reg_0461;
    62: op1_15_in28 = reg_1168;
    81: op1_15_in28 = reg_0191;
    82: op1_15_in28 = reg_0780;
    63: op1_15_in28 = reg_1018;
    52: op1_15_in28 = reg_0413;
    83: op1_15_in28 = reg_1517;
    89: op1_15_in28 = reg_0151;
    84: op1_15_in28 = reg_0715;
    85: op1_15_in28 = reg_0014;
    65: op1_15_in28 = reg_1000;
    90: op1_15_in28 = reg_0215;
    91: op1_15_in28 = reg_0466;
    46: op1_15_in28 = reg_0720;
    48: op1_15_in28 = reg_0709;
    67: op1_15_in28 = reg_0401;
    92: op1_15_in28 = reg_0783;
    93: op1_15_in28 = reg_0457;
    94: op1_15_in28 = reg_1214;
    95: op1_15_in28 = reg_0726;
    96: op1_15_in28 = reg_0335;
    97: op1_15_in28 = reg_0289;
    100: op1_15_in28 = reg_0271;
    101: op1_15_in28 = reg_0668;
    102: op1_15_in28 = reg_1164;
    103: op1_15_in28 = reg_0023;
    104: op1_15_in28 = reg_0043;
    105: op1_15_in28 = reg_0362;
    106: op1_15_in28 = reg_0878;
    107: op1_15_in28 = reg_0368;
    108: op1_15_in28 = imem02_in[15:12];
    109: op1_15_in28 = reg_0226;
    110: op1_15_in28 = reg_1184;
    112: op1_15_in28 = reg_0790;
    113: op1_15_in28 = reg_0634;
    114: op1_15_in28 = reg_0601;
    116: op1_15_in28 = reg_0602;
    117: op1_15_in28 = reg_1350;
    118: op1_15_in28 = reg_0228;
    119: op1_15_in28 = reg_0146;
    47: op1_15_in28 = reg_0137;
    120: op1_15_in28 = reg_0965;
    121: op1_15_in28 = reg_0251;
    122: op1_15_in28 = reg_0234;
    123: op1_15_in28 = reg_0548;
    124: op1_15_in28 = reg_0791;
    126: op1_15_in28 = reg_0028;
    127: op1_15_in28 = reg_0299;
    128: op1_15_in28 = reg_1340;
    129: op1_15_in28 = reg_0039;
    130: op1_15_in28 = reg_0209;
    default: op1_15_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の28番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv28 = 1;
    73: op1_15_inv28 = 1;
    53: op1_15_inv28 = 1;
    86: op1_15_inv28 = 1;
    54: op1_15_inv28 = 1;
    76: op1_15_inv28 = 1;
    87: op1_15_inv28 = 1;
    57: op1_15_inv28 = 1;
    50: op1_15_inv28 = 1;
    68: op1_15_inv28 = 1;
    71: op1_15_inv28 = 1;
    78: op1_15_inv28 = 1;
    61: op1_15_inv28 = 1;
    70: op1_15_inv28 = 1;
    59: op1_15_inv28 = 1;
    79: op1_15_inv28 = 1;
    88: op1_15_inv28 = 1;
    81: op1_15_inv28 = 1;
    63: op1_15_inv28 = 1;
    84: op1_15_inv28 = 1;
    85: op1_15_inv28 = 1;
    65: op1_15_inv28 = 1;
    90: op1_15_inv28 = 1;
    46: op1_15_inv28 = 1;
    92: op1_15_inv28 = 1;
    93: op1_15_inv28 = 1;
    94: op1_15_inv28 = 1;
    97: op1_15_inv28 = 1;
    98: op1_15_inv28 = 1;
    100: op1_15_inv28 = 1;
    102: op1_15_inv28 = 1;
    105: op1_15_inv28 = 1;
    107: op1_15_inv28 = 1;
    108: op1_15_inv28 = 1;
    110: op1_15_inv28 = 1;
    112: op1_15_inv28 = 1;
    113: op1_15_inv28 = 1;
    119: op1_15_inv28 = 1;
    47: op1_15_inv28 = 1;
    120: op1_15_inv28 = 1;
    122: op1_15_inv28 = 1;
    123: op1_15_inv28 = 1;
    125: op1_15_inv28 = 1;
    126: op1_15_inv28 = 1;
    127: op1_15_inv28 = 1;
    129: op1_15_inv28 = 1;
    default: op1_15_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の29番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in29 = imem01_in[7:4];
    73: op1_15_in29 = reg_0119;
    53: op1_15_in29 = reg_0747;
    86: op1_15_in29 = reg_0369;
    74: op1_15_in29 = reg_0091;
    54: op1_15_in29 = reg_0313;
    75: op1_15_in29 = reg_0031;
    69: op1_15_in29 = reg_0962;
    56: op1_15_in29 = reg_0379;
    76: op1_15_in29 = reg_0421;
    87: op1_15_in29 = reg_0420;
    57: op1_15_in29 = reg_0326;
    50: op1_15_in29 = reg_0559;
    68: op1_15_in29 = reg_0130;
    71: op1_15_in29 = reg_0384;
    67: op1_15_in29 = reg_0384;
    77: op1_15_in29 = reg_0156;
    78: op1_15_in29 = reg_0324;
    61: op1_15_in29 = reg_0902;
    58: op1_15_in29 = reg_0540;
    70: op1_15_in29 = reg_0798;
    59: op1_15_in29 = reg_0573;
    79: op1_15_in29 = reg_0787;
    51: op1_15_in29 = reg_0177;
    88: op1_15_in29 = reg_0601;
    80: op1_15_in29 = reg_1183;
    62: op1_15_in29 = reg_1169;
    81: op1_15_in29 = reg_0889;
    82: op1_15_in29 = reg_0115;
    63: op1_15_in29 = reg_1207;
    52: op1_15_in29 = reg_0137;
    83: op1_15_in29 = reg_0190;
    89: op1_15_in29 = reg_0037;
    84: op1_15_in29 = reg_0572;
    85: op1_15_in29 = reg_1437;
    65: op1_15_in29 = reg_0954;
    90: op1_15_in29 = reg_0490;
    91: op1_15_in29 = reg_0278;
    46: op1_15_in29 = reg_0827;
    48: op1_15_in29 = reg_0378;
    92: op1_15_in29 = reg_0234;
    93: op1_15_in29 = reg_1350;
    94: op1_15_in29 = reg_1065;
    95: op1_15_in29 = reg_0146;
    96: op1_15_in29 = reg_0079;
    97: op1_15_in29 = reg_1202;
    98: op1_15_in29 = reg_0262;
    100: op1_15_in29 = reg_1467;
    101: op1_15_in29 = reg_0530;
    102: op1_15_in29 = reg_0167;
    103: op1_15_in29 = reg_0214;
    104: op1_15_in29 = reg_0042;
    105: op1_15_in29 = reg_0162;
    106: op1_15_in29 = reg_0560;
    107: op1_15_in29 = reg_0862;
    108: op1_15_in29 = reg_0254;
    109: op1_15_in29 = reg_0394;
    110: op1_15_in29 = reg_1517;
    112: op1_15_in29 = reg_0936;
    113: op1_15_in29 = reg_0043;
    114: op1_15_in29 = reg_0196;
    116: op1_15_in29 = reg_0828;
    117: op1_15_in29 = reg_0923;
    118: op1_15_in29 = reg_0001;
    119: op1_15_in29 = reg_0290;
    47: op1_15_in29 = reg_0228;
    120: op1_15_in29 = reg_0070;
    121: op1_15_in29 = reg_0700;
    122: op1_15_in29 = reg_0505;
    123: op1_15_in29 = reg_0819;
    124: op1_15_in29 = reg_1010;
    125: op1_15_in29 = reg_0896;
    126: op1_15_in29 = reg_0235;
    127: op1_15_in29 = reg_0159;
    128: op1_15_in29 = reg_1151;
    129: op1_15_in29 = reg_1299;
    130: op1_15_in29 = reg_0064;
    default: op1_15_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の29番目の入力反転
  always @ ( * ) begin
    case ( state )
    72: op1_15_inv29 = 1;
    53: op1_15_inv29 = 1;
    86: op1_15_inv29 = 1;
    74: op1_15_inv29 = 1;
    54: op1_15_inv29 = 1;
    75: op1_15_inv29 = 1;
    56: op1_15_inv29 = 1;
    76: op1_15_inv29 = 1;
    87: op1_15_inv29 = 1;
    50: op1_15_inv29 = 1;
    68: op1_15_inv29 = 1;
    77: op1_15_inv29 = 1;
    78: op1_15_inv29 = 1;
    70: op1_15_inv29 = 1;
    79: op1_15_inv29 = 1;
    62: op1_15_inv29 = 1;
    81: op1_15_inv29 = 1;
    82: op1_15_inv29 = 1;
    89: op1_15_inv29 = 1;
    84: op1_15_inv29 = 1;
    85: op1_15_inv29 = 1;
    91: op1_15_inv29 = 1;
    92: op1_15_inv29 = 1;
    95: op1_15_inv29 = 1;
    96: op1_15_inv29 = 1;
    98: op1_15_inv29 = 1;
    102: op1_15_inv29 = 1;
    104: op1_15_inv29 = 1;
    110: op1_15_inv29 = 1;
    112: op1_15_inv29 = 1;
    116: op1_15_inv29 = 1;
    117: op1_15_inv29 = 1;
    119: op1_15_inv29 = 1;
    120: op1_15_inv29 = 1;
    121: op1_15_inv29 = 1;
    124: op1_15_inv29 = 1;
    125: op1_15_inv29 = 1;
    126: op1_15_inv29 = 1;
    129: op1_15_inv29 = 1;
    default: op1_15_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の30番目の入力
  always @ ( * ) begin
    case ( state )
    72: op1_15_in30 = imem01_in[11:8];
    73: op1_15_in30 = reg_0269;
    53: op1_15_in30 = imem01_in[15:12];
    86: op1_15_in30 = reg_0262;
    74: op1_15_in30 = reg_0899;
    54: op1_15_in30 = reg_0755;
    75: op1_15_in30 = reg_0663;
    69: op1_15_in30 = reg_0627;
    120: op1_15_in30 = reg_0627;
    56: op1_15_in30 = reg_0900;
    76: op1_15_in30 = reg_0471;
    87: op1_15_in30 = reg_0633;
    57: op1_15_in30 = reg_0106;
    50: op1_15_in30 = reg_0557;
    68: op1_15_in30 = reg_0602;
    71: op1_15_in30 = reg_0386;
    77: op1_15_in30 = reg_0924;
    78: op1_15_in30 = reg_1440;
    61: op1_15_in30 = reg_0013;
    58: op1_15_in30 = reg_0541;
    70: op1_15_in30 = reg_1419;
    59: op1_15_in30 = reg_0677;
    79: op1_15_in30 = reg_0222;
    51: op1_15_in30 = reg_0964;
    88: op1_15_in30 = reg_0243;
    80: op1_15_in30 = reg_0245;
    62: op1_15_in30 = reg_0697;
    81: op1_15_in30 = reg_0233;
    82: op1_15_in30 = reg_0716;
    63: op1_15_in30 = reg_0429;
    52: op1_15_in30 = reg_0103;
    83: op1_15_in30 = reg_1300;
    89: op1_15_in30 = reg_0753;
    84: op1_15_in30 = reg_0968;
    85: op1_15_in30 = reg_0192;
    65: op1_15_in30 = reg_0597;
    90: op1_15_in30 = reg_1439;
    91: op1_15_in30 = reg_0347;
    46: op1_15_in30 = reg_0714;
    48: op1_15_in30 = reg_0376;
    67: op1_15_in30 = reg_0385;
    92: op1_15_in30 = reg_0180;
    93: op1_15_in30 = reg_1349;
    94: op1_15_in30 = reg_1004;
    95: op1_15_in30 = reg_0402;
    96: op1_15_in30 = reg_0896;
    97: op1_15_in30 = reg_1179;
    98: op1_15_in30 = reg_0096;
    100: op1_15_in30 = reg_0720;
    101: op1_15_in30 = imem02_in[7:4];
    102: op1_15_in30 = reg_1180;
    103: op1_15_in30 = reg_0015;
    104: op1_15_in30 = reg_0044;
    105: op1_15_in30 = reg_0728;
    106: op1_15_in30 = reg_0695;
    107: op1_15_in30 = reg_0337;
    108: op1_15_in30 = reg_0455;
    109: op1_15_in30 = reg_1010;
    110: op1_15_in30 = reg_0957;
    112: op1_15_in30 = reg_0328;
    113: op1_15_in30 = reg_0042;
    114: op1_15_in30 = reg_0575;
    116: op1_15_in30 = reg_0565;
    117: op1_15_in30 = reg_0740;
    118: op1_15_in30 = reg_0053;
    126: op1_15_in30 = reg_0053;
    119: op1_15_in30 = reg_0868;
    47: op1_15_in30 = reg_0521;
    121: op1_15_in30 = reg_0648;
    122: op1_15_in30 = reg_0756;
    123: op1_15_in30 = reg_0149;
    124: op1_15_in30 = reg_0667;
    125: op1_15_in30 = reg_0447;
    127: op1_15_in30 = reg_0158;
    128: op1_15_in30 = reg_1237;
    129: op1_15_in30 = reg_0669;
    130: op1_15_in30 = reg_1503;
    default: op1_15_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の30番目の入力反転
  always @ ( * ) begin
    case ( state )
    86: op1_15_inv30 = 1;
    54: op1_15_inv30 = 1;
    75: op1_15_inv30 = 1;
    57: op1_15_inv30 = 1;
    50: op1_15_inv30 = 1;
    68: op1_15_inv30 = 1;
    77: op1_15_inv30 = 1;
    78: op1_15_inv30 = 1;
    61: op1_15_inv30 = 1;
    58: op1_15_inv30 = 1;
    70: op1_15_inv30 = 1;
    59: op1_15_inv30 = 1;
    79: op1_15_inv30 = 1;
    82: op1_15_inv30 = 1;
    83: op1_15_inv30 = 1;
    89: op1_15_inv30 = 1;
    90: op1_15_inv30 = 1;
    92: op1_15_inv30 = 1;
    93: op1_15_inv30 = 1;
    95: op1_15_inv30 = 1;
    97: op1_15_inv30 = 1;
    101: op1_15_inv30 = 1;
    102: op1_15_inv30 = 1;
    105: op1_15_inv30 = 1;
    106: op1_15_inv30 = 1;
    107: op1_15_inv30 = 1;
    108: op1_15_inv30 = 1;
    110: op1_15_inv30 = 1;
    112: op1_15_inv30 = 1;
    114: op1_15_inv30 = 1;
    123: op1_15_inv30 = 1;
    125: op1_15_inv30 = 1;
    127: op1_15_inv30 = 1;
    default: op1_15_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_15_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#15の31番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_15_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の0番目の入力
  always @ ( * ) begin
    case ( state )
    21: op2_00_in00 = reg_0049;
    36: op2_00_in00 = reg_0625;
    46: op2_00_in00 = reg_0865;
    53: op2_00_in00 = reg_0394;
    87: op2_00_in00 = reg_0394;
    59: op2_00_in00 = reg_0298;
    68: op2_00_in00 = reg_0988;
    77: op2_00_in00 = reg_0498;
    69: op2_00_in00 = reg_0226;
    79: op2_00_in00 = reg_0226;
    88: op2_00_in00 = reg_1483;
    74: op2_00_in00 = reg_0611;
    73: op2_00_in00 = reg_1002;
    70: op2_00_in00 = reg_0324;
    89: op2_00_in00 = reg_0757;
    75: op2_00_in00 = reg_1153;
    76: op2_00_in00 = reg_0539;
    61: op2_00_in00 = reg_0639;
    72: op2_00_in00 = reg_0150;
    78: op2_00_in00 = reg_0563;
    80: op2_00_in00 = reg_0422;
    81: op2_00_in00 = reg_0745;
    90: op2_00_in00 = reg_0248;
    82: op2_00_in00 = reg_0355;
    83: op2_00_in00 = reg_1353;
    84: op2_00_in00 = reg_1125;
    65: op2_00_in00 = reg_0193;
    105: op2_00_in00 = reg_0193;
    131: op2_00_in00 = reg_0193;
    85: op2_00_in00 = reg_1101;
    91: op2_00_in00 = reg_1288;
    86: op2_00_in00 = reg_0668;
    92: op2_00_in00 = reg_0036;
    93: op2_00_in00 = reg_0721;
    96: op2_00_in00 = reg_0721;
    94: op2_00_in00 = reg_1413;
    95: op2_00_in00 = reg_0074;
    101: op2_00_in00 = reg_0074;
    111: op2_00_in00 = reg_0074;
    113: op2_00_in00 = reg_0074;
    117: op2_00_in00 = reg_0074;
    129: op2_00_in00 = reg_0074;
    97: op2_00_in00 = reg_0758;
    103: op2_00_in00 = reg_0758;
    107: op2_00_in00 = reg_0758;
    110: op2_00_in00 = reg_0758;
    98: op2_00_in00 = reg_0843;
    99: op2_00_in00 = reg_1049;
    102: op2_00_in00 = reg_1049;
    100: op2_00_in00 = reg_0658;
    104: op2_00_in00 = reg_0658;
    109: op2_00_in00 = reg_0658;
    123: op2_00_in00 = reg_0658;
    106: op2_00_in00 = reg_0660;
    115: op2_00_in00 = reg_0660;
    121: op2_00_in00 = reg_0660;
    127: op2_00_in00 = reg_0660;
    108: op2_00_in00 = reg_0614;
    112: op2_00_in00 = reg_0516;
    122: op2_00_in00 = reg_0516;
    114: op2_00_in00 = reg_0772;
    116: op2_00_in00 = reg_0515;
    118: op2_00_in00 = reg_0771;
    130: op2_00_in00 = reg_0771;
    119: op2_00_in00 = reg_0259;
    120: op2_00_in00 = reg_0511;
    124: op2_00_in00 = reg_0211;
    125: op2_00_in00 = reg_0517;
    126: op2_00_in00 = reg_0446;
    128: op2_00_in00 = reg_0770;
    132: op2_00_in00 = reg_0641;
    default: op2_00_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の1番目の入力
  always @ ( * ) begin
    case ( state )
    21: op2_00_in01 = reg_0265;
    36: op2_00_in01 = reg_0694;
    46: op2_00_in01 = reg_0781;
    53: op2_00_in01 = reg_1138;
    59: op2_00_in01 = reg_0988;
    88: op2_00_in01 = reg_0988;
    73: op2_00_in01 = reg_0988;
    68: op2_00_in01 = reg_0485;
    77: op2_00_in01 = reg_1091;
    69: op2_00_in01 = reg_1054;
    74: op2_00_in01 = reg_0931;
    87: op2_00_in01 = reg_1114;
    70: op2_00_in01 = reg_0164;
    89: op2_00_in01 = reg_0200;
    75: op2_00_in01 = reg_1185;
    76: op2_00_in01 = reg_0367;
    61: op2_00_in01 = reg_1232;
    72: op2_00_in01 = reg_0721;
    78: op2_00_in01 = reg_0581;
    79: op2_00_in01 = reg_0936;
    80: op2_00_in01 = reg_1097;
    81: op2_00_in01 = reg_1130;
    90: op2_00_in01 = reg_1165;
    82: op2_00_in01 = reg_1043;
    83: op2_00_in01 = reg_0668;
    84: op2_00_in01 = reg_0725;
    86: op2_00_in01 = reg_0725;
    65: op2_00_in01 = reg_0641;
    85: op2_00_in01 = reg_0826;
    91: op2_00_in01 = reg_1387;
    92: op2_00_in01 = reg_1398;
    93: op2_00_in01 = reg_0900;
    94: op2_00_in01 = reg_1089;
    95: op2_00_in01 = reg_0226;
    117: op2_00_in01 = reg_0226;
    96: op2_00_in01 = reg_0606;
    108: op2_00_in01 = reg_0606;
    97: op2_00_in01 = reg_0074;
    103: op2_00_in01 = reg_0074;
    107: op2_00_in01 = reg_0074;
    115: op2_00_in01 = reg_0074;
    121: op2_00_in01 = reg_0074;
    125: op2_00_in01 = reg_0074;
    127: op2_00_in01 = reg_0074;
    98: op2_00_in01 = reg_0036;
    106: op2_00_in01 = reg_0036;
    110: op2_00_in01 = reg_0036;
    99: op2_00_in01 = reg_0642;
    100: op2_00_in01 = reg_0659;
    101: op2_00_in01 = reg_0266;
    102: op2_00_in01 = reg_0756;
    104: op2_00_in01 = reg_0516;
    109: op2_00_in01 = reg_0516;
    105: op2_00_in01 = reg_0515;
    126: op2_00_in01 = reg_0515;
    131: op2_00_in01 = reg_0515;
    111: op2_00_in01 = reg_0761;
    113: op2_00_in01 = reg_0761;
    112: op2_00_in01 = reg_0660;
    124: op2_00_in01 = reg_0660;
    114: op2_00_in01 = reg_0517;
    122: op2_00_in01 = reg_0517;
    116: op2_00_in01 = reg_1016;
    118: op2_00_in01 = reg_0772;
    123: op2_00_in01 = reg_0772;
    130: op2_00_in01 = reg_0772;
    119: op2_00_in01 = reg_0446;
    120: op2_00_in01 = reg_0512;
    128: op2_00_in01 = reg_0658;
    129: op2_00_in01 = reg_0099;
    132: op2_00_in01 = reg_0920;
    default: op2_00_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の2番目の入力
  always @ ( * ) begin
    case ( state )
    21: op2_00_in02 = reg_0322;
    36: op2_00_in02 = reg_0594;
    46: op2_00_in02 = reg_0594;
    53: op2_00_in02 = reg_1054;
    59: op2_00_in02 = reg_1142;
    61: op2_00_in02 = reg_1142;
    68: op2_00_in02 = reg_0049;
    77: op2_00_in02 = reg_0783;
    69: op2_00_in02 = reg_0230;
    90: op2_00_in02 = reg_0230;
    88: op2_00_in02 = reg_0725;
    74: op2_00_in02 = reg_0985;
    87: op2_00_in02 = reg_0498;
    73: op2_00_in02 = reg_0990;
    70: op2_00_in02 = reg_1002;
    89: op2_00_in02 = reg_1428;
    75: op2_00_in02 = reg_0977;
    76: op2_00_in02 = reg_1152;
    72: op2_00_in02 = reg_0749;
    78: op2_00_in02 = reg_1236;
    79: op2_00_in02 = reg_0825;
    80: op2_00_in02 = reg_1460;
    81: op2_00_in02 = reg_0447;
    82: op2_00_in02 = reg_0324;
    83: op2_00_in02 = reg_0036;
    94: op2_00_in02 = reg_0036;
    96: op2_00_in02 = reg_0036;
    108: op2_00_in02 = reg_0036;
    112: op2_00_in02 = reg_0036;
    114: op2_00_in02 = reg_0036;
    122: op2_00_in02 = reg_0036;
    124: op2_00_in02 = reg_0036;
    84: op2_00_in02 = reg_0834;
    65: op2_00_in02 = reg_0642;
    85: op2_00_in02 = reg_1332;
    91: op2_00_in02 = reg_0074;
    86: op2_00_in02 = reg_1376;
    92: op2_00_in02 = reg_0081;
    98: op2_00_in02 = reg_0081;
    106: op2_00_in02 = reg_0081;
    110: op2_00_in02 = reg_0081;
    93: op2_00_in02 = reg_1016;
    95: op2_00_in02 = reg_0082;
    101: op2_00_in02 = reg_0082;
    111: op2_00_in02 = reg_0082;
    113: op2_00_in02 = reg_0082;
    117: op2_00_in02 = reg_0082;
    129: op2_00_in02 = reg_0082;
    97: op2_00_in02 = reg_0423;
    99: op2_00_in02 = reg_0606;
    102: op2_00_in02 = reg_0606;
    100: op2_00_in02 = reg_0758;
    116: op2_00_in02 = reg_0758;
    103: op2_00_in02 = reg_0857;
    104: op2_00_in02 = reg_1017;
    105: op2_00_in02 = reg_0756;
    107: op2_00_in02 = reg_0761;
    109: op2_00_in02 = reg_0660;
    118: op2_00_in02 = reg_0660;
    130: op2_00_in02 = reg_0660;
    115: op2_00_in02 = reg_0226;
    119: op2_00_in02 = reg_0515;
    120: op2_00_in02 = reg_0513;
    121: op2_00_in02 = reg_0231;
    123: op2_00_in02 = reg_0773;
    125: op2_00_in02 = reg_0099;
    127: op2_00_in02 = reg_0099;
    126: op2_00_in02 = reg_0772;
    128: op2_00_in02 = reg_0516;
    131: op2_00_in02 = reg_0516;
    132: op2_00_in02 = reg_0659;
    default: op2_00_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の3番目の入力
  always @ ( * ) begin
    case ( state )
    21: op2_00_in03 = reg_0200;
    36: op2_00_in03 = reg_0447;
    77: op2_00_in03 = reg_0447;
    46: op2_00_in03 = reg_0344;
    53: op2_00_in03 = reg_0988;
    59: op2_00_in03 = reg_0694;
    68: op2_00_in03 = reg_0726;
    69: op2_00_in03 = reg_0581;
    88: op2_00_in03 = reg_0230;
    74: op2_00_in03 = reg_0367;
    87: op2_00_in03 = reg_1217;
    73: op2_00_in03 = reg_0062;
    70: op2_00_in03 = reg_0989;
    89: op2_00_in03 = reg_1178;
    75: op2_00_in03 = reg_0990;
    76: op2_00_in03 = reg_0560;
    61: op2_00_in03 = reg_1061;
    72: op2_00_in03 = reg_1106;
    78: op2_00_in03 = reg_0179;
    79: op2_00_in03 = reg_0941;
    80: op2_00_in03 = reg_0499;
    81: op2_00_in03 = reg_1141;
    90: op2_00_in03 = reg_1341;
    82: op2_00_in03 = reg_1156;
    83: op2_00_in03 = reg_1157;
    84: op2_00_in03 = reg_1162;
    65: op2_00_in03 = reg_0838;
    85: op2_00_in03 = reg_1042;
    91: op2_00_in03 = reg_1130;
    86: op2_00_in03 = reg_1009;
    92: op2_00_in03 = reg_0643;
    93: op2_00_in03 = reg_1060;
    94: op2_00_in03 = reg_0081;
    108: op2_00_in03 = reg_0081;
    112: op2_00_in03 = reg_0081;
    114: op2_00_in03 = reg_0081;
    122: op2_00_in03 = reg_0081;
    124: op2_00_in03 = reg_0081;
    95: op2_00_in03 = reg_0654;
    101: op2_00_in03 = reg_0654;
    96: op2_00_in03 = reg_0856;
    97: op2_00_in03 = reg_0082;
    107: op2_00_in03 = reg_0082;
    115: op2_00_in03 = reg_0082;
    121: op2_00_in03 = reg_0082;
    125: op2_00_in03 = reg_0082;
    127: op2_00_in03 = reg_0082;
    98: op2_00_in03 = reg_0354;
    106: op2_00_in03 = reg_0354;
    110: op2_00_in03 = reg_0354;
    99: op2_00_in03 = reg_0074;
    109: op2_00_in03 = reg_0074;
    123: op2_00_in03 = reg_0074;
    100: op2_00_in03 = reg_0036;
    102: op2_00_in03 = reg_0036;
    104: op2_00_in03 = reg_0036;
    116: op2_00_in03 = reg_0036;
    118: op2_00_in03 = reg_0036;
    130: op2_00_in03 = reg_0036;
    103: op2_00_in03 = reg_0226;
    105: op2_00_in03 = reg_0606;
    132: op2_00_in03 = reg_0606;
    111: op2_00_in03 = reg_0355;
    113: op2_00_in03 = reg_0355;
    117: op2_00_in03 = reg_0355;
    129: op2_00_in03 = reg_0355;
    119: op2_00_in03 = reg_0516;
    120: op2_00_in03 = reg_0770;
    126: op2_00_in03 = reg_0773;
    128: op2_00_in03 = reg_0517;
    131: op2_00_in03 = reg_0517;
    default: op2_00_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の4番目の入力
  always @ ( * ) begin
    case ( state )
    21: op2_00_in04 = reg_0266;
    36: op2_00_in04 = reg_0248;
    46: op2_00_in04 = reg_0394;
    68: op2_00_in04 = reg_1062;
    77: op2_00_in04 = reg_1001;
    69: op2_00_in04 = reg_1138;
    88: op2_00_in04 = reg_1270;
    87: op2_00_in04 = reg_1496;
    73: op2_00_in04 = reg_0991;
    70: op2_00_in04 = reg_0447;
    89: op2_00_in04 = reg_0344;
    75: op2_00_in04 = reg_1072;
    76: op2_00_in04 = reg_1075;
    61: op2_00_in04 = reg_0074;
    93: op2_00_in04 = reg_0074;
    105: op2_00_in04 = reg_0074;
    131: op2_00_in04 = reg_0074;
    72: op2_00_in04 = reg_1234;
    79: op2_00_in04 = reg_0826;
    80: op2_00_in04 = reg_1125;
    81: op2_00_in04 = reg_1304;
    90: op2_00_in04 = reg_1342;
    82: op2_00_in04 = reg_1061;
    83: op2_00_in04 = reg_1158;
    84: op2_00_in04 = reg_0503;
    65: op2_00_in04 = reg_0643;
    85: op2_00_in04 = reg_1374;
    91: op2_00_in04 = reg_0781;
    86: op2_00_in04 = reg_0852;
    92: op2_00_in04 = reg_0354;
    94: op2_00_in04 = reg_0354;
    122: op2_00_in04 = reg_0354;
    95: op2_00_in04 = reg_0658;
    120: op2_00_in04 = reg_0658;
    97: op2_00_in04 = reg_0654;
    107: op2_00_in04 = reg_0654;
    98: op2_00_in04 = reg_0076;
    106: op2_00_in04 = reg_0076;
    100: op2_00_in04 = reg_0081;
    104: op2_00_in04 = reg_0081;
    130: op2_00_in04 = reg_0081;
    101: op2_00_in04 = reg_0760;
    113: op2_00_in04 = reg_0760;
    103: op2_00_in04 = reg_0082;
    108: op2_00_in04 = reg_0482;
    109: op2_00_in04 = reg_0761;
    111: op2_00_in04 = reg_0129;
    112: op2_00_in04 = reg_0808;
    114: op2_00_in04 = reg_0099;
    115: op2_00_in04 = reg_0811;
    117: op2_00_in04 = reg_0324;
    129: op2_00_in04 = reg_0324;
    118: op2_00_in04 = reg_0359;
    119: op2_00_in04 = reg_0517;
    121: op2_00_in04 = reg_0355;
    125: op2_00_in04 = reg_0355;
    127: op2_00_in04 = reg_0355;
    123: op2_00_in04 = reg_0545;
    124: op2_00_in04 = reg_0101;
    126: op2_00_in04 = reg_0036;
    128: op2_00_in04 = reg_0036;
    132: op2_00_in04 = reg_0036;
    default: op2_00_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の5番目の入力
  always @ ( * ) begin
    case ( state )
    77: op2_00_in05 = reg_0847;
    87: op2_00_in05 = reg_1084;
    81: op2_00_in05 = reg_0759;
    92: op2_00_in05 = reg_0767;
    93: op2_00_in05 = reg_0902;
    94: op2_00_in05 = reg_0657;
    106: op2_00_in05 = reg_0687;
    119: op2_00_in05 = reg_0074;
    120: op2_00_in05 = reg_1016;
    132: op2_00_in05 = reg_0081;
    default: op2_00_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の6番目の入力
  always @ ( * ) begin
    case ( state )
    93: op2_00_in06 = reg_0512;
    120: op2_00_in06 = reg_0758;
    132: op2_00_in06 = reg_0693;
    default: op2_00_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の7番目の入力
  always @ ( * ) begin
    case ( state )
    120: op2_00_in07 = reg_0036;
    default: op2_00_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#0のバイアス入力
  always @ ( * ) begin
    case ( state )
    21: op2_00_bias = 80;
    36: op2_00_bias = 67;
    46: op2_00_bias = 64;
    53: op2_00_bias = 57;
    59: op2_00_bias = 55;
    68: op2_00_bias = 66;
    77: op2_00_bias = 86;
    69: op2_00_bias = 62;
    88: op2_00_bias = 63;
    74: op2_00_bias = 55;
    87: op2_00_bias = 81;
    73: op2_00_bias = 83;
    70: op2_00_bias = 57;
    89: op2_00_bias = 70;
    75: op2_00_bias = 65;
    76: op2_00_bias = 71;
    61: op2_00_bias = 61;
    72: op2_00_bias = 79;
    78: op2_00_bias = 73;
    79: op2_00_bias = 74;
    80: op2_00_bias = 65;
    81: op2_00_bias = 82;
    90: op2_00_bias = 75;
    82: op2_00_bias = 71;
    83: op2_00_bias = 68;
    84: op2_00_bias = 62;
    65: op2_00_bias = 66;
    85: op2_00_bias = 56;
    91: op2_00_bias = 64;
    86: op2_00_bias = 70;
    92: op2_00_bias = 80;
    93: op2_00_bias = 83;
    94: op2_00_bias = 86;
    95: op2_00_bias = 67;
    96: op2_00_bias = 45;
    97: op2_00_bias = 75;
    98: op2_00_bias = 68;
    99: op2_00_bias = 54;
    100: op2_00_bias = 72;
    101: op2_00_bias = 64;
    102: op2_00_bias = 55;
    103: op2_00_bias = 69;
    104: op2_00_bias = 71;
    105: op2_00_bias = 64;
    106: op2_00_bias = 86;
    107: op2_00_bias = 84;
    108: op2_00_bias = 74;
    109: op2_00_bias = 70;
    110: op2_00_bias = 63;
    111: op2_00_bias = 74;
    112: op2_00_bias = 61;
    113: op2_00_bias = 63;
    114: op2_00_bias = 57;
    115: op2_00_bias = 72;
    116: op2_00_bias = 69;
    117: op2_00_bias = 75;
    118: op2_00_bias = 69;
    119: op2_00_bias = 73;
    120: op2_00_bias = 107;
    121: op2_00_bias = 61;
    122: op2_00_bias = 78;
    123: op2_00_bias = 56;
    124: op2_00_bias = 61;
    125: op2_00_bias = 78;
    126: op2_00_bias = 65;
    127: op2_00_bias = 78;
    128: op2_00_bias = 65;
    129: op2_00_bias = 72;
    130: op2_00_bias = 84;
    131: op2_00_bias = 83;
    132: op2_00_bias = 76;
    default: op2_00_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#1の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_01_in00 = reg_1140;
    74: op2_01_in00 = reg_0839;
    73: op2_01_in00 = reg_0259;
    75: op2_01_in00 = reg_0129;
    95: op2_01_in00 = reg_0129;
    76: op2_01_in00 = reg_0745;
    88: op2_01_in00 = reg_0678;
    77: op2_01_in00 = reg_0226;
    93: op2_01_in00 = reg_0226;
    72: op2_01_in00 = reg_0209;
    78: op2_01_in00 = reg_1108;
    89: op2_01_in00 = reg_1075;
    79: op2_01_in00 = reg_0603;
    80: op2_01_in00 = reg_0668;
    81: op2_01_in00 = reg_0639;
    90: op2_01_in00 = reg_0499;
    82: op2_01_in00 = reg_0502;
    83: op2_01_in00 = reg_1236;
    84: op2_01_in00 = reg_1007;
    85: op2_01_in00 = reg_1128;
    91: op2_01_in00 = reg_0729;
    86: op2_01_in00 = reg_0503;
    92: op2_01_in00 = reg_0076;
    94: op2_01_in00 = reg_0076;
    110: op2_01_in00 = reg_0076;
    122: op2_01_in00 = reg_0076;
    124: op2_01_in00 = reg_0076;
    96: op2_01_in00 = reg_0081;
    102: op2_01_in00 = reg_0081;
    116: op2_01_in00 = reg_0081;
    118: op2_01_in00 = reg_0081;
    120: op2_01_in00 = reg_0081;
    126: op2_01_in00 = reg_0081;
    128: op2_01_in00 = reg_0081;
    97: op2_01_in00 = reg_0760;
    107: op2_01_in00 = reg_0760;
    98: op2_01_in00 = reg_0083;
    106: op2_01_in00 = reg_0083;
    99: op2_01_in00 = reg_0834;
    100: op2_01_in00 = reg_0354;
    104: op2_01_in00 = reg_0354;
    108: op2_01_in00 = reg_0354;
    112: op2_01_in00 = reg_0354;
    114: op2_01_in00 = reg_0354;
    101: op2_01_in00 = reg_0625;
    111: op2_01_in00 = reg_0625;
    113: op2_01_in00 = reg_0625;
    117: op2_01_in00 = reg_0625;
    129: op2_01_in00 = reg_0625;
    103: op2_01_in00 = reg_0654;
    105: op2_01_in00 = reg_0761;
    109: op2_01_in00 = reg_0082;
    115: op2_01_in00 = reg_0355;
    119: op2_01_in00 = reg_0543;
    121: op2_01_in00 = reg_0324;
    125: op2_01_in00 = reg_0324;
    123: op2_01_in00 = reg_0231;
    127: op2_01_in00 = reg_0546;
    130: op2_01_in00 = reg_0101;
    132: op2_01_in00 = reg_0101;
    131: op2_01_in00 = reg_0099;
    default: op2_01_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_01_in01 = reg_1045;
    74: op2_01_in01 = reg_0986;
    73: op2_01_in01 = reg_0792;
    75: op2_01_in01 = reg_1110;
    76: op2_01_in01 = reg_0179;
    72: op2_01_in01 = reg_0179;
    80: op2_01_in01 = reg_0179;
    88: op2_01_in01 = reg_1446;
    77: op2_01_in01 = reg_1004;
    78: op2_01_in01 = reg_0933;
    89: op2_01_in01 = reg_1429;
    79: op2_01_in01 = reg_1104;
    81: op2_01_in01 = reg_1131;
    90: op2_01_in01 = reg_0354;
    96: op2_01_in01 = reg_0354;
    102: op2_01_in01 = reg_0354;
    116: op2_01_in01 = reg_0354;
    118: op2_01_in01 = reg_0354;
    120: op2_01_in01 = reg_0354;
    82: op2_01_in01 = reg_0376;
    83: op2_01_in01 = reg_1354;
    84: op2_01_in01 = reg_0729;
    85: op2_01_in01 = reg_1044;
    91: op2_01_in01 = reg_0226;
    86: op2_01_in01 = reg_0871;
    92: op2_01_in01 = reg_1048;
    93: op2_01_in01 = reg_0082;
    99: op2_01_in01 = reg_0082;
    105: op2_01_in01 = reg_0082;
    119: op2_01_in01 = reg_0082;
    123: op2_01_in01 = reg_0082;
    131: op2_01_in01 = reg_0082;
    94: op2_01_in01 = reg_0083;
    110: op2_01_in01 = reg_0083;
    122: op2_01_in01 = reg_0083;
    124: op2_01_in01 = reg_0083;
    95: op2_01_in01 = reg_0625;
    97: op2_01_in01 = reg_0625;
    107: op2_01_in01 = reg_0625;
    121: op2_01_in01 = reg_0625;
    125: op2_01_in01 = reg_0625;
    127: op2_01_in01 = reg_0625;
    98: op2_01_in01 = reg_0358;
    106: op2_01_in01 = reg_0358;
    100: op2_01_in01 = reg_0076;
    104: op2_01_in01 = reg_0076;
    108: op2_01_in01 = reg_0076;
    112: op2_01_in01 = reg_0076;
    114: op2_01_in01 = reg_0076;
    130: op2_01_in01 = reg_0076;
    132: op2_01_in01 = reg_0076;
    101: op2_01_in01 = reg_0356;
    111: op2_01_in01 = reg_0356;
    113: op2_01_in01 = reg_0356;
    117: op2_01_in01 = reg_0356;
    129: op2_01_in01 = reg_0356;
    103: op2_01_in01 = reg_0760;
    109: op2_01_in01 = reg_0355;
    115: op2_01_in01 = reg_0324;
    126: op2_01_in01 = reg_0101;
    128: op2_01_in01 = reg_0101;
    default: op2_01_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_01_in02 = reg_0834;
    74: op2_01_in02 = reg_1062;
    73: op2_01_in02 = reg_0888;
    75: op2_01_in02 = reg_0904;
    76: op2_01_in02 = reg_1236;
    88: op2_01_in02 = reg_1352;
    77: op2_01_in02 = reg_1099;
    72: op2_01_in02 = reg_0634;
    78: op2_01_in02 = reg_1423;
    89: op2_01_in02 = reg_0628;
    79: op2_01_in02 = reg_1041;
    80: op2_01_in02 = reg_0248;
    81: op2_01_in02 = reg_1305;
    90: op2_01_in02 = reg_0081;
    82: op2_01_in02 = reg_1333;
    83: op2_01_in02 = reg_0639;
    84: op2_01_in02 = reg_0753;
    85: op2_01_in02 = reg_1375;
    91: op2_01_in02 = reg_1388;
    86: op2_01_in02 = reg_1377;
    92: op2_01_in02 = reg_0083;
    100: op2_01_in02 = reg_0083;
    104: op2_01_in02 = reg_0083;
    108: op2_01_in02 = reg_0083;
    112: op2_01_in02 = reg_0083;
    114: op2_01_in02 = reg_0083;
    130: op2_01_in02 = reg_0083;
    132: op2_01_in02 = reg_0083;
    93: op2_01_in02 = reg_0903;
    94: op2_01_in02 = reg_0358;
    110: op2_01_in02 = reg_0358;
    122: op2_01_in02 = reg_0358;
    124: op2_01_in02 = reg_0358;
    95: op2_01_in02 = reg_0356;
    97: op2_01_in02 = reg_0356;
    107: op2_01_in02 = reg_0356;
    121: op2_01_in02 = reg_0356;
    125: op2_01_in02 = reg_0356;
    127: op2_01_in02 = reg_0356;
    96: op2_01_in02 = reg_0076;
    102: op2_01_in02 = reg_0076;
    116: op2_01_in02 = reg_0076;
    118: op2_01_in02 = reg_0076;
    120: op2_01_in02 = reg_0076;
    126: op2_01_in02 = reg_0076;
    98: op2_01_in02 = reg_0764;
    106: op2_01_in02 = reg_0764;
    99: op2_01_in02 = reg_0654;
    105: op2_01_in02 = reg_0654;
    101: op2_01_in02 = reg_0645;
    111: op2_01_in02 = reg_0645;
    113: op2_01_in02 = reg_0645;
    117: op2_01_in02 = reg_0645;
    103: op2_01_in02 = reg_0625;
    109: op2_01_in02 = reg_0760;
    115: op2_01_in02 = reg_0763;
    119: op2_01_in02 = reg_0355;
    123: op2_01_in02 = reg_0355;
    131: op2_01_in02 = reg_0355;
    128: op2_01_in02 = reg_0956;
    129: op2_01_in02 = reg_0510;
    default: op2_01_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_01_in03 = reg_1476;
    74: op2_01_in03 = reg_0179;
    73: op2_01_in03 = reg_0446;
    75: op2_01_in03 = reg_1066;
    76: op2_01_in03 = reg_0985;
    88: op2_01_in03 = reg_1088;
    77: op2_01_in03 = reg_0603;
    72: op2_01_in03 = reg_0467;
    78: op2_01_in03 = reg_1040;
    89: op2_01_in03 = reg_1188;
    79: op2_01_in03 = reg_1095;
    82: op2_01_in03 = reg_1095;
    80: op2_01_in03 = reg_1126;
    81: op2_01_in03 = reg_0500;
    90: op2_01_in03 = reg_1166;
    83: op2_01_in03 = reg_0076;
    128: op2_01_in03 = reg_0076;
    84: op2_01_in03 = reg_1043;
    85: op2_01_in03 = reg_1058;
    91: op2_01_in03 = reg_1037;
    86: op2_01_in03 = reg_0652;
    92: op2_01_in03 = reg_0358;
    100: op2_01_in03 = reg_0358;
    104: op2_01_in03 = reg_0358;
    112: op2_01_in03 = reg_0358;
    114: op2_01_in03 = reg_0358;
    130: op2_01_in03 = reg_0358;
    132: op2_01_in03 = reg_0358;
    93: op2_01_in03 = reg_0929;
    94: op2_01_in03 = reg_0376;
    110: op2_01_in03 = reg_0376;
    95: op2_01_in03 = reg_0645;
    97: op2_01_in03 = reg_0645;
    107: op2_01_in03 = reg_0645;
    96: op2_01_in03 = reg_0083;
    116: op2_01_in03 = reg_0083;
    118: op2_01_in03 = reg_0083;
    120: op2_01_in03 = reg_0083;
    126: op2_01_in03 = reg_0083;
    98: op2_01_in03 = reg_0510;
    125: op2_01_in03 = reg_0510;
    127: op2_01_in03 = reg_0510;
    99: op2_01_in03 = reg_0760;
    105: op2_01_in03 = reg_0760;
    101: op2_01_in03 = reg_0949;
    102: op2_01_in03 = reg_1019;
    103: op2_01_in03 = reg_0356;
    115: op2_01_in03 = reg_0356;
    106: op2_01_in03 = reg_1021;
    108: op2_01_in03 = reg_0951;
    109: op2_01_in03 = reg_0625;
    111: op2_01_in03 = reg_0766;
    113: op2_01_in03 = reg_0647;
    117: op2_01_in03 = reg_0647;
    119: op2_01_in03 = reg_0231;
    121: op2_01_in03 = reg_1025;
    122: op2_01_in03 = reg_0687;
    124: op2_01_in03 = reg_0687;
    123: op2_01_in03 = reg_0324;
    131: op2_01_in03 = reg_0324;
    129: op2_01_in03 = reg_0539;
    default: op2_01_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_01_in04 = reg_1218;
    74: op2_01_in04 = reg_1209;
    75: op2_01_in04 = reg_1213;
    76: op2_01_in04 = reg_1237;
    77: op2_01_in04 = reg_1238;
    72: op2_01_in04 = reg_0633;
    78: op2_01_in04 = reg_1058;
    89: op2_01_in04 = reg_0656;
    81: op2_01_in04 = reg_1306;
    90: op2_01_in04 = reg_0763;
    105: op2_01_in04 = reg_0763;
    82: op2_01_in04 = reg_0850;
    83: op2_01_in04 = reg_1355;
    84: op2_01_in04 = reg_0652;
    85: op2_01_in04 = reg_0625;
    123: op2_01_in04 = reg_0625;
    131: op2_01_in04 = reg_0625;
    86: op2_01_in04 = reg_1378;
    92: op2_01_in04 = reg_1399;
    93: op2_01_in04 = reg_0423;
    94: op2_01_in04 = reg_0510;
    95: op2_01_in04 = reg_0766;
    97: op2_01_in04 = reg_0766;
    101: op2_01_in04 = reg_0766;
    107: op2_01_in04 = reg_0766;
    96: op2_01_in04 = reg_0358;
    108: op2_01_in04 = reg_0358;
    116: op2_01_in04 = reg_0358;
    118: op2_01_in04 = reg_0358;
    98: op2_01_in04 = reg_0503;
    99: op2_01_in04 = reg_0677;
    100: op2_01_in04 = reg_0769;
    102: op2_01_in04 = reg_0083;
    128: op2_01_in04 = reg_0083;
    103: op2_01_in04 = reg_0645;
    115: op2_01_in04 = reg_0645;
    104: op2_01_in04 = reg_0376;
    112: op2_01_in04 = reg_0376;
    114: op2_01_in04 = reg_0376;
    106: op2_01_in04 = reg_0771;
    109: op2_01_in04 = reg_0356;
    110: op2_01_in04 = reg_0098;
    111: op2_01_in04 = reg_0517;
    113: op2_01_in04 = reg_0511;
    117: op2_01_in04 = reg_0812;
    119: op2_01_in04 = reg_0324;
    121: op2_01_in04 = reg_0101;
    122: op2_01_in04 = reg_0359;
    124: op2_01_in04 = reg_0690;
    127: op2_01_in04 = reg_0692;
    129: op2_01_in04 = reg_0816;
    130: op2_01_in04 = reg_0687;
    132: op2_01_in04 = reg_0687;
    default: op2_01_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の5番目の入力
  always @ ( * ) begin
    case ( state )
    75: op2_01_in05 = reg_0498;
    78: op2_01_in05 = reg_1059;
    104: op2_01_in05 = reg_0770;
    114: op2_01_in05 = reg_0810;
    115: op2_01_in05 = reg_0543;
    119: op2_01_in05 = reg_0424;
    123: op2_01_in05 = reg_0356;
    131: op2_01_in05 = reg_0551;
    132: op2_01_in05 = reg_0359;
    default: op2_01_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の6番目の入力
  always @ ( * ) begin
    case ( state )
    123: op2_01_in06 = reg_0510;
    default: op2_01_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の7番目の入力
  always @ ( * ) begin
    case ( state )
    123: op2_01_in07 = reg_0546;
    default: op2_01_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#1の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_01_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#1のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_01_bias = 68;
    74: op2_01_bias = 72;
    73: op2_01_bias = 59;
    75: op2_01_bias = 89;
    76: op2_01_bias = 83;
    88: op2_01_bias = 58;
    77: op2_01_bias = 70;
    72: op2_01_bias = 70;
    78: op2_01_bias = 90;
    89: op2_01_bias = 72;
    79: op2_01_bias = 61;
    80: op2_01_bias = 55;
    81: op2_01_bias = 67;
    90: op2_01_bias = 71;
    82: op2_01_bias = 72;
    83: op2_01_bias = 71;
    84: op2_01_bias = 75;
    85: op2_01_bias = 84;
    91: op2_01_bias = 64;
    86: op2_01_bias = 78;
    92: op2_01_bias = 79;
    93: op2_01_bias = 72;
    94: op2_01_bias = 78;
    95: op2_01_bias = 81;
    96: op2_01_bias = 72;
    97: op2_01_bias = 77;
    98: op2_01_bias = 84;
    99: op2_01_bias = 84;
    100: op2_01_bias = 69;
    101: op2_01_bias = 68;
    102: op2_01_bias = 73;
    103: op2_01_bias = 64;
    104: op2_01_bias = 80;
    105: op2_01_bias = 72;
    106: op2_01_bias = 79;
    107: op2_01_bias = 78;
    108: op2_01_bias = 66;
    109: op2_01_bias = 78;
    110: op2_01_bias = 68;
    111: op2_01_bias = 63;
    112: op2_01_bias = 62;
    113: op2_01_bias = 72;
    114: op2_01_bias = 64;
    115: op2_01_bias = 73;
    116: op2_01_bias = 71;
    117: op2_01_bias = 56;
    118: op2_01_bias = 72;
    119: op2_01_bias = 84;
    120: op2_01_bias = 57;
    121: op2_01_bias = 60;
    122: op2_01_bias = 84;
    123: op2_01_bias = 119;
    124: op2_01_bias = 74;
    125: op2_01_bias = 64;
    126: op2_01_bias = 72;
    127: op2_01_bias = 63;
    128: op2_01_bias = 72;
    129: op2_01_bias = 68;
    130: op2_01_bias = 68;
    131: op2_01_bias = 83;
    132: op2_01_bias = 89;
    default: op2_01_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#2の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_02_in00 = reg_1477;
    74: op2_02_in00 = reg_1107;
    73: op2_02_in00 = reg_0533;
    75: op2_02_in00 = reg_0989;
    76: op2_02_in00 = reg_0164;
    88: op2_02_in00 = reg_1109;
    77: op2_02_in00 = reg_0129;
    78: op2_02_in00 = reg_1110;
    89: op2_02_in00 = reg_0758;
    79: op2_02_in00 = reg_1073;
    80: op2_02_in00 = reg_0935;
    81: op2_02_in00 = reg_1039;
    90: op2_02_in00 = reg_0539;
    125: op2_02_in00 = reg_0539;
    127: op2_02_in00 = reg_0539;
    82: op2_02_in00 = reg_0535;
    84: op2_02_in00 = reg_0535;
    83: op2_02_in00 = reg_0826;
    91: op2_02_in00 = reg_0909;
    86: op2_02_in00 = reg_0926;
    92: op2_02_in00 = reg_0764;
    96: op2_02_in00 = reg_0764;
    93: op2_02_in00 = reg_0062;
    94: op2_02_in00 = reg_0503;
    122: op2_02_in00 = reg_0503;
    95: op2_02_in00 = reg_0511;
    97: op2_02_in00 = reg_0511;
    101: op2_02_in00 = reg_0511;
    107: op2_02_in00 = reg_0511;
    111: op2_02_in00 = reg_0511;
    117: op2_02_in00 = reg_0511;
    98: op2_02_in00 = reg_0538;
    99: op2_02_in00 = reg_0356;
    105: op2_02_in00 = reg_0356;
    131: op2_02_in00 = reg_0356;
    100: op2_02_in00 = reg_0376;
    102: op2_02_in00 = reg_0358;
    120: op2_02_in00 = reg_0358;
    126: op2_02_in00 = reg_0358;
    128: op2_02_in00 = reg_0358;
    103: op2_02_in00 = reg_0766;
    104: op2_02_in00 = reg_0510;
    106: op2_02_in00 = reg_0510;
    110: op2_02_in00 = reg_0510;
    112: op2_02_in00 = reg_0510;
    114: op2_02_in00 = reg_0510;
    121: op2_02_in00 = reg_0510;
    108: op2_02_in00 = reg_0687;
    116: op2_02_in00 = reg_0687;
    118: op2_02_in00 = reg_0687;
    109: op2_02_in00 = reg_0645;
    113: op2_02_in00 = reg_0512;
    115: op2_02_in00 = reg_0647;
    123: op2_02_in00 = reg_0647;
    119: op2_02_in00 = reg_0625;
    124: op2_02_in00 = reg_0359;
    130: op2_02_in00 = reg_0359;
    129: op2_02_in00 = reg_0651;
    132: op2_02_in00 = reg_0364;
    default: op2_02_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_02_in01 = reg_1442;
    74: op2_02_in01 = reg_0794;
    73: op2_02_in01 = reg_0983;
    75: op2_02_in01 = reg_0982;
    76: op2_02_in01 = reg_1188;
    88: op2_02_in01 = reg_1374;
    77: op2_02_in01 = reg_1239;
    78: op2_02_in01 = reg_1060;
    89: op2_02_in01 = reg_1076;
    79: op2_02_in01 = reg_1122;
    80: op2_02_in01 = reg_0867;
    81: op2_02_in01 = reg_1328;
    90: op2_02_in01 = reg_0538;
    82: op2_02_in01 = reg_1352;
    83: op2_02_in01 = reg_1159;
    84: op2_02_in01 = reg_0782;
    91: op2_02_in01 = reg_0644;
    86: op2_02_in01 = reg_1379;
    92: op2_02_in01 = reg_0641;
    93: op2_02_in01 = reg_0682;
    94: op2_02_in01 = reg_0705;
    95: op2_02_in01 = reg_0512;
    101: op2_02_in01 = reg_0512;
    107: op2_02_in01 = reg_0512;
    111: op2_02_in01 = reg_0512;
    117: op2_02_in01 = reg_0512;
    96: op2_02_in01 = reg_0510;
    100: op2_02_in01 = reg_0510;
    108: op2_02_in01 = reg_0510;
    116: op2_02_in01 = reg_0510;
    118: op2_02_in01 = reg_0510;
    131: op2_02_in01 = reg_0510;
    97: op2_02_in01 = reg_0915;
    98: op2_02_in01 = reg_0150;
    99: op2_02_in01 = reg_0645;
    105: op2_02_in01 = reg_0645;
    102: op2_02_in01 = reg_0376;
    103: op2_02_in01 = reg_0511;
    115: op2_02_in01 = reg_0511;
    122: op2_02_in01 = reg_0511;
    132: op2_02_in01 = reg_0511;
    104: op2_02_in01 = reg_0503;
    106: op2_02_in01 = reg_0503;
    110: op2_02_in01 = reg_0503;
    112: op2_02_in01 = reg_0503;
    114: op2_02_in01 = reg_0503;
    124: op2_02_in01 = reg_0503;
    130: op2_02_in01 = reg_0503;
    109: op2_02_in01 = reg_0766;
    113: op2_02_in01 = reg_0513;
    119: op2_02_in01 = reg_0356;
    120: op2_02_in01 = reg_0687;
    126: op2_02_in01 = reg_0687;
    128: op2_02_in01 = reg_0687;
    121: op2_02_in01 = reg_0647;
    123: op2_02_in01 = reg_0651;
    125: op2_02_in01 = reg_0651;
    127: op2_02_in01 = reg_0651;
    129: op2_02_in01 = reg_0919;
    default: op2_02_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_02_in02 = reg_0611;
    89: op2_02_in02 = reg_0611;
    74: op2_02_in02 = reg_0959;
    73: op2_02_in02 = reg_0793;
    75: op2_02_in02 = reg_1235;
    76: op2_02_in02 = reg_1421;
    88: op2_02_in02 = reg_1195;
    77: op2_02_in02 = reg_1039;
    78: op2_02_in02 = reg_0635;
    79: op2_02_in02 = reg_1054;
    80: op2_02_in02 = reg_1461;
    81: op2_02_in02 = reg_0825;
    90: op2_02_in02 = reg_0762;
    82: op2_02_in02 = reg_0193;
    86: op2_02_in02 = reg_0193;
    83: op2_02_in02 = reg_1356;
    84: op2_02_in02 = reg_0784;
    91: op2_02_in02 = reg_0082;
    92: op2_02_in02 = reg_0510;
    102: op2_02_in02 = reg_0510;
    93: op2_02_in02 = reg_0958;
    94: op2_02_in02 = reg_0150;
    122: op2_02_in02 = reg_0150;
    132: op2_02_in02 = reg_0150;
    95: op2_02_in02 = reg_0513;
    101: op2_02_in02 = reg_0513;
    107: op2_02_in02 = reg_0513;
    111: op2_02_in02 = reg_0513;
    117: op2_02_in02 = reg_0513;
    96: op2_02_in02 = reg_0503;
    100: op2_02_in02 = reg_0503;
    116: op2_02_in02 = reg_0503;
    118: op2_02_in02 = reg_0503;
    97: op2_02_in02 = reg_0512;
    103: op2_02_in02 = reg_0512;
    115: op2_02_in02 = reg_0512;
    123: op2_02_in02 = reg_0512;
    125: op2_02_in02 = reg_0512;
    127: op2_02_in02 = reg_0512;
    129: op2_02_in02 = reg_0512;
    98: op2_02_in02 = reg_0259;
    99: op2_02_in02 = reg_0766;
    105: op2_02_in02 = reg_0766;
    104: op2_02_in02 = reg_0705;
    106: op2_02_in02 = reg_0705;
    110: op2_02_in02 = reg_0705;
    112: op2_02_in02 = reg_0705;
    108: op2_02_in02 = reg_1022;
    109: op2_02_in02 = reg_0511;
    124: op2_02_in02 = reg_0511;
    130: op2_02_in02 = reg_0511;
    113: op2_02_in02 = reg_1015;
    114: op2_02_in02 = reg_0651;
    119: op2_02_in02 = reg_0645;
    120: op2_02_in02 = reg_0359;
    126: op2_02_in02 = reg_0359;
    128: op2_02_in02 = reg_0359;
    121: op2_02_in02 = reg_1026;
    131: op2_02_in02 = reg_0539;
    default: op2_02_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_02_in03 = reg_0467;
    74: op2_02_in03 = reg_0450;
    73: op2_02_in03 = reg_1037;
    75: op2_02_in03 = reg_0793;
    76: op2_02_in03 = reg_1108;
    91: op2_02_in03 = reg_1108;
    88: op2_02_in03 = reg_1067;
    77: op2_02_in03 = reg_1111;
    78: op2_02_in03 = reg_0538;
    131: op2_02_in03 = reg_0538;
    89: op2_02_in03 = reg_0614;
    79: op2_02_in03 = reg_1123;
    80: op2_02_in03 = reg_0376;
    81: op2_02_in03 = reg_1329;
    90: op2_02_in03 = reg_0581;
    82: op2_02_in03 = reg_1096;
    86: op2_02_in03 = reg_1096;
    83: op2_02_in03 = reg_1160;
    84: op2_02_in03 = reg_0829;
    92: op2_02_in03 = reg_0503;
    102: op2_02_in03 = reg_0503;
    108: op2_02_in03 = reg_0503;
    126: op2_02_in03 = reg_0503;
    128: op2_02_in03 = reg_0503;
    93: op2_02_in03 = reg_1017;
    94: op2_02_in03 = reg_0259;
    123: op2_02_in03 = reg_0259;
    125: op2_02_in03 = reg_0259;
    95: op2_02_in03 = reg_0634;
    96: op2_02_in03 = reg_0948;
    97: op2_02_in03 = reg_0513;
    103: op2_02_in03 = reg_0513;
    115: op2_02_in03 = reg_0513;
    122: op2_02_in03 = reg_0513;
    98: op2_02_in03 = reg_0446;
    99: op2_02_in03 = reg_0511;
    100: op2_02_in03 = reg_0705;
    101: op2_02_in03 = reg_0514;
    104: op2_02_in03 = reg_0150;
    110: op2_02_in03 = reg_0150;
    112: op2_02_in03 = reg_0150;
    114: op2_02_in03 = reg_0150;
    124: op2_02_in03 = reg_0150;
    130: op2_02_in03 = reg_0150;
    105: op2_02_in03 = reg_0950;
    106: op2_02_in03 = reg_0768;
    107: op2_02_in03 = reg_0193;
    109: op2_02_in03 = reg_0512;
    111: op2_02_in03 = reg_1015;
    113: op2_02_in03 = reg_0515;
    116: op2_02_in03 = reg_0651;
    118: op2_02_in03 = reg_0651;
    117: op2_02_in03 = reg_0770;
    119: op2_02_in03 = reg_1024;
    120: op2_02_in03 = reg_0858;
    127: op2_02_in03 = reg_0955;
    129: op2_02_in03 = reg_0643;
    132: op2_02_in03 = reg_0209;
    default: op2_02_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_02_in04 = reg_1190;
    74: op2_02_in04 = reg_1184;
    73: op2_02_in04 = reg_1066;
    75: op2_02_in04 = reg_1073;
    76: op2_02_in04 = reg_0422;
    88: op2_02_in04 = reg_0853;
    78: op2_02_in04 = reg_0670;
    89: op2_02_in04 = reg_1133;
    80: op2_02_in04 = reg_1098;
    81: op2_02_in04 = reg_0760;
    90: op2_02_in04 = reg_1357;
    82: op2_02_in04 = reg_1097;
    83: op2_02_in04 = reg_0651;
    84: op2_02_in04 = reg_0871;
    91: op2_02_in04 = reg_1389;
    86: op2_02_in04 = reg_1380;
    92: op2_02_in04 = reg_0913;
    93: op2_02_in04 = reg_1036;
    94: op2_02_in04 = reg_0446;
    123: op2_02_in04 = reg_0446;
    129: op2_02_in04 = reg_0446;
    95: op2_02_in04 = reg_0728;
    96: op2_02_in04 = reg_0538;
    97: op2_02_in04 = reg_0657;
    98: op2_02_in04 = reg_0515;
    107: op2_02_in04 = reg_0515;
    111: op2_02_in04 = reg_0515;
    99: op2_02_in04 = reg_0512;
    100: op2_02_in04 = reg_0150;
    116: op2_02_in04 = reg_0150;
    118: op2_02_in04 = reg_0150;
    101: op2_02_in04 = reg_0516;
    102: op2_02_in04 = reg_0705;
    103: op2_02_in04 = reg_0514;
    104: op2_02_in04 = reg_0259;
    110: op2_02_in04 = reg_0259;
    127: op2_02_in04 = reg_0259;
    105: op2_02_in04 = reg_0511;
    126: op2_02_in04 = reg_0511;
    109: op2_02_in04 = reg_0772;
    112: op2_02_in04 = reg_0809;
    113: op2_02_in04 = reg_0688;
    114: op2_02_in04 = reg_0542;
    115: op2_02_in04 = reg_0770;
    117: op2_02_in04 = reg_0813;
    119: op2_02_in04 = reg_0647;
    120: op2_02_in04 = reg_0503;
    122: op2_02_in04 = reg_0193;
    124: op2_02_in04 = reg_0691;
    130: op2_02_in04 = reg_0513;
    131: op2_02_in04 = reg_0818;
    132: op2_02_in04 = reg_0417;
    default: op2_02_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の5番目の入力
  always @ ( * ) begin
    case ( state )
    78: op2_02_in05 = reg_0499;
    89: op2_02_in05 = reg_0684;
    90: op2_02_in05 = reg_0357;
    82: op2_02_in05 = reg_0682;
    92: op2_02_in05 = reg_0768;
    95: op2_02_in05 = reg_0659;
    96: op2_02_in05 = reg_0514;
    97: op2_02_in05 = reg_0658;
    99: op2_02_in05 = reg_0513;
    105: op2_02_in05 = reg_0512;
    111: op2_02_in05 = reg_0807;
    116: op2_02_in05 = reg_0544;
    120: op2_02_in05 = reg_0689;
    123: op2_02_in05 = reg_0515;
    127: op2_02_in05 = reg_0814;
    129: op2_02_in05 = reg_0817;
    130: op2_02_in05 = reg_0364;
    default: op2_02_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の6番目の入力
  always @ ( * ) begin
    case ( state )
    97: op2_02_in06 = reg_0659;
    99: op2_02_in06 = reg_0514;
    default: op2_02_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#2の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_02_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#2のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_02_bias = 62;
    74: op2_02_bias = 74;
    73: op2_02_bias = 64;
    75: op2_02_bias = 62;
    76: op2_02_bias = 77;
    88: op2_02_bias = 79;
    77: op2_02_bias = 62;
    78: op2_02_bias = 72;
    89: op2_02_bias = 87;
    79: op2_02_bias = 67;
    80: op2_02_bias = 71;
    81: op2_02_bias = 69;
    90: op2_02_bias = 85;
    82: op2_02_bias = 84;
    83: op2_02_bias = 69;
    84: op2_02_bias = 70;
    91: op2_02_bias = 69;
    86: op2_02_bias = 64;
    92: op2_02_bias = 78;
    93: op2_02_bias = 66;
    94: op2_02_bias = 79;
    95: op2_02_bias = 81;
    96: op2_02_bias = 79;
    97: op2_02_bias = 85;
    98: op2_02_bias = 64;
    99: op2_02_bias = 118;
    100: op2_02_bias = 66;
    101: op2_02_bias = 71;
    102: op2_02_bias = 70;
    103: op2_02_bias = 74;
    104: op2_02_bias = 71;
    105: op2_02_bias = 98;
    106: op2_02_bias = 64;
    107: op2_02_bias = 72;
    108: op2_02_bias = 51;
    109: op2_02_bias = 65;
    110: op2_02_bias = 67;
    111: op2_02_bias = 84;
    112: op2_02_bias = 71;
    113: op2_02_bias = 69;
    114: op2_02_bias = 63;
    115: op2_02_bias = 58;
    116: op2_02_bias = 81;
    117: op2_02_bias = 67;
    118: op2_02_bias = 80;
    119: op2_02_bias = 69;
    120: op2_02_bias = 97;
    121: op2_02_bias = 57;
    122: op2_02_bias = 71;
    123: op2_02_bias = 86;
    124: op2_02_bias = 61;
    125: op2_02_bias = 51;
    126: op2_02_bias = 87;
    127: op2_02_bias = 69;
    128: op2_02_bias = 54;
    129: op2_02_bias = 72;
    130: op2_02_bias = 78;
    131: op2_02_bias = 67;
    132: op2_02_bias = 64;
    default: op2_02_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#3の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_03_in00 = reg_1292;
    74: op2_03_in00 = reg_0538;
    92: op2_03_in00 = reg_0538;
    75: op2_03_in00 = reg_0259;
    100: op2_03_in00 = reg_0259;
    106: op2_03_in00 = reg_0259;
    112: op2_03_in00 = reg_0259;
    114: op2_03_in00 = reg_0259;
    116: op2_03_in00 = reg_0259;
    76: op2_03_in00 = reg_0615;
    88: op2_03_in00 = reg_1146;
    77: op2_03_in00 = reg_0982;
    78: op2_03_in00 = reg_0535;
    89: op2_03_in00 = reg_1099;
    79: op2_03_in00 = reg_0556;
    80: op2_03_in00 = reg_1327;
    81: op2_03_in00 = reg_1330;
    90: op2_03_in00 = reg_1142;
    83: op2_03_in00 = reg_1288;
    84: op2_03_in00 = reg_0193;
    91: op2_03_in00 = reg_0356;
    86: op2_03_in00 = reg_1161;
    93: op2_03_in00 = reg_0625;
    94: op2_03_in00 = reg_0914;
    96: op2_03_in00 = reg_0768;
    102: op2_03_in00 = reg_0768;
    105: op2_03_in00 = reg_0513;
    109: op2_03_in00 = reg_0513;
    124: op2_03_in00 = reg_0513;
    108: op2_03_in00 = reg_0705;
    121: op2_03_in00 = reg_0705;
    110: op2_03_in00 = reg_0770;
    120: op2_03_in00 = reg_0651;
    126: op2_03_in00 = reg_0150;
    128: op2_03_in00 = reg_0511;
    131: op2_03_in00 = reg_0512;
    default: op2_03_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_03_in01 = reg_1115;
    74: op2_03_in01 = reg_1090;
    75: op2_03_in01 = reg_1186;
    76: op2_03_in01 = reg_1189;
    88: op2_03_in01 = reg_1328;
    77: op2_03_in01 = reg_1438;
    78: op2_03_in01 = reg_1113;
    89: op2_03_in01 = reg_1271;
    79: op2_03_in01 = reg_1063;
    80: op2_03_in01 = reg_1007;
    81: op2_03_in01 = reg_1155;
    90: op2_03_in01 = reg_0654;
    83: op2_03_in01 = reg_1130;
    84: op2_03_in01 = reg_0893;
    91: op2_03_in01 = reg_1390;
    86: op2_03_in01 = reg_1381;
    92: op2_03_in01 = reg_0642;
    93: op2_03_in01 = reg_0356;
    94: op2_03_in01 = reg_0533;
    96: op2_03_in01 = reg_0259;
    102: op2_03_in01 = reg_0259;
    131: op2_03_in01 = reg_0259;
    100: op2_03_in01 = reg_0657;
    105: op2_03_in01 = reg_0514;
    106: op2_03_in01 = reg_0770;
    112: op2_03_in01 = reg_0770;
    108: op2_03_in01 = reg_0150;
    128: op2_03_in01 = reg_0150;
    109: op2_03_in01 = reg_0446;
    110: op2_03_in01 = reg_0771;
    114: op2_03_in01 = reg_0193;
    116: op2_03_in01 = reg_0193;
    124: op2_03_in01 = reg_0193;
    120: op2_03_in01 = reg_0916;
    121: op2_03_in01 = reg_0581;
    126: op2_03_in01 = reg_0513;
    default: op2_03_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_03_in02 = reg_1122;
    74: op2_03_in02 = reg_1210;
    75: op2_03_in02 = reg_0932;
    76: op2_03_in02 = reg_1422;
    88: op2_03_in02 = reg_1196;
    77: op2_03_in02 = reg_1240;
    78: op2_03_in02 = reg_1424;
    89: op2_03_in02 = reg_0129;
    79: op2_03_in02 = reg_1006;
    80: op2_03_in02 = reg_1283;
    81: op2_03_in02 = reg_0826;
    90: op2_03_in02 = reg_1014;
    83: op2_03_in02 = reg_0745;
    84: op2_03_in02 = reg_0926;
    91: op2_03_in02 = reg_0670;
    86: op2_03_in02 = reg_1131;
    92: op2_03_in02 = reg_0150;
    120: op2_03_in02 = reg_0150;
    93: op2_03_in02 = reg_1055;
    94: op2_03_in02 = reg_0642;
    96: op2_03_in02 = reg_0446;
    102: op2_03_in02 = reg_0446;
    100: op2_03_in02 = reg_0515;
    109: op2_03_in02 = reg_0515;
    105: op2_03_in02 = reg_1049;
    106: op2_03_in02 = reg_0658;
    112: op2_03_in02 = reg_0658;
    114: op2_03_in02 = reg_0658;
    116: op2_03_in02 = reg_0658;
    108: op2_03_in02 = reg_1023;
    110: op2_03_in02 = reg_0614;
    121: op2_03_in02 = reg_0259;
    124: op2_03_in02 = reg_0641;
    126: op2_03_in02 = reg_0193;
    128: op2_03_in02 = reg_0513;
    131: op2_03_in02 = reg_0453;
    default: op2_03_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_03_in03 = reg_0749;
    74: op2_03_in03 = reg_0150;
    75: op2_03_in03 = reg_1187;
    76: op2_03_in03 = reg_0538;
    88: op2_03_in03 = reg_1245;
    77: op2_03_in03 = reg_0793;
    78: op2_03_in03 = reg_1434;
    89: op2_03_in03 = reg_0676;
    79: op2_03_in03 = reg_1422;
    80: op2_03_in03 = reg_0539;
    81: op2_03_in03 = reg_1054;
    90: op2_03_in03 = reg_1358;
    83: op2_03_in03 = reg_1161;
    84: op2_03_in03 = reg_1096;
    91: op2_03_in03 = reg_0784;
    86: op2_03_in03 = reg_1382;
    92: op2_03_in03 = reg_0947;
    93: op2_03_in03 = reg_1407;
    94: op2_03_in03 = reg_0843;
    96: op2_03_in03 = reg_0533;
    100: op2_03_in03 = reg_0614;
    112: op2_03_in03 = reg_0614;
    102: op2_03_in03 = reg_0515;
    105: op2_03_in03 = reg_1016;
    106: op2_03_in03 = reg_0516;
    114: op2_03_in03 = reg_0516;
    116: op2_03_in03 = reg_0516;
    124: op2_03_in03 = reg_0516;
    108: op2_03_in03 = reg_0259;
    109: op2_03_in03 = reg_0756;
    110: op2_03_in03 = reg_1017;
    120: op2_03_in03 = reg_0535;
    121: op2_03_in03 = reg_0446;
    131: op2_03_in03 = reg_0446;
    126: op2_03_in03 = reg_0953;
    128: op2_03_in03 = reg_0193;
    default: op2_03_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_03_in04 = reg_1085;
    74: op2_03_in04 = reg_1067;
    75: op2_03_in04 = reg_0603;
    76: op2_03_in04 = reg_1076;
    77: op2_03_in04 = reg_0644;
    78: op2_03_in04 = reg_0645;
    89: op2_03_in04 = reg_0890;
    79: op2_03_in04 = reg_0500;
    80: op2_03_in04 = reg_0501;
    81: op2_03_in04 = reg_0076;
    84: op2_03_in04 = reg_0356;
    91: op2_03_in04 = reg_0765;
    92: op2_03_in04 = reg_1049;
    93: op2_03_in04 = reg_0513;
    94: op2_03_in04 = reg_0855;
    96: op2_03_in04 = reg_0642;
    100: op2_03_in04 = reg_0843;
    102: op2_03_in04 = reg_0614;
    105: op2_03_in04 = reg_1020;
    108: op2_03_in04 = reg_0770;
    110: op2_03_in04 = reg_0773;
    112: op2_03_in04 = reg_0758;
    116: op2_03_in04 = reg_0517;
    120: op2_03_in04 = reg_0193;
    121: op2_03_in04 = reg_0515;
    126: op2_03_in04 = reg_0641;
    default: op2_03_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の5番目の入力
  always @ ( * ) begin
    case ( state )
    89: op2_03_in05 = reg_1272;
    92: op2_03_in05 = reg_1400;
    102: op2_03_in05 = reg_0660;
    120: op2_03_in05 = reg_0771;
    126: op2_03_in05 = reg_0211;
    default: op2_03_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の6番目の入力
  always @ ( * ) begin
    case ( state )
    120: op2_03_in06 = reg_0772;
    default: op2_03_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#3の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_03_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#3のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_03_bias = 84;
    74: op2_03_bias = 70;
    75: op2_03_bias = 75;
    76: op2_03_bias = 83;
    88: op2_03_bias = 51;
    77: op2_03_bias = 65;
    78: op2_03_bias = 65;
    89: op2_03_bias = 101;
    79: op2_03_bias = 62;
    80: op2_03_bias = 63;
    81: op2_03_bias = 68;
    90: op2_03_bias = 63;
    83: op2_03_bias = 64;
    84: op2_03_bias = 60;
    91: op2_03_bias = 76;
    86: op2_03_bias = 65;
    92: op2_03_bias = 90;
    93: op2_03_bias = 65;
    94: op2_03_bias = 64;
    96: op2_03_bias = 70;
    100: op2_03_bias = 70;
    102: op2_03_bias = 74;
    105: op2_03_bias = 64;
    106: op2_03_bias = 50;
    108: op2_03_bias = 61;
    109: op2_03_bias = 51;
    110: op2_03_bias = 63;
    112: op2_03_bias = 82;
    114: op2_03_bias = 61;
    116: op2_03_bias = 73;
    120: op2_03_bias = 102;
    121: op2_03_bias = 74;
    124: op2_03_bias = 66;
    126: op2_03_bias = 86;
    128: op2_03_bias = 53;
    131: op2_03_bias = 50;
    default: op2_03_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#4の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_04_in00 = reg_1293;
    74: op2_04_in00 = reg_0164;
    75: op2_04_in00 = reg_0446;
    88: op2_04_in00 = reg_0150;
    77: op2_04_in00 = reg_1072;
    78: op2_04_in00 = reg_1154;
    89: op2_04_in00 = reg_1319;
    79: op2_04_in00 = reg_0259;
    92: op2_04_in00 = reg_0259;
    80: op2_04_in00 = reg_0538;
    81: op2_04_in00 = reg_1056;
    90: op2_04_in00 = reg_0760;
    91: op2_04_in00 = reg_0129;
    93: op2_04_in00 = reg_1408;
    128: op2_04_in00 = reg_0515;
    default: op2_04_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_04_in01 = reg_1307;
    74: op2_04_in01 = reg_1211;
    75: op2_04_in01 = reg_1434;
    88: op2_04_in01 = reg_1197;
    77: op2_04_in01 = reg_0230;
    78: op2_04_in01 = reg_0935;
    89: op2_04_in01 = reg_1273;
    79: op2_04_in01 = reg_1124;
    80: op2_04_in01 = reg_1462;
    81: op2_04_in01 = reg_1331;
    90: op2_04_in01 = reg_0164;
    91: op2_04_in01 = reg_1391;
    92: op2_04_in01 = reg_0446;
    93: op2_04_in01 = reg_1409;
    128: op2_04_in01 = reg_0918;
    default: op2_04_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_04_in02 = reg_1039;
    74: op2_04_in02 = reg_0209;
    75: op2_04_in02 = reg_1056;
    88: op2_04_in02 = reg_1123;
    77: op2_04_in02 = reg_1101;
    78: op2_04_in02 = reg_0671;
    89: op2_04_in02 = reg_0749;
    79: op2_04_in02 = reg_1111;
    80: op2_04_in02 = reg_1463;
    81: op2_04_in02 = reg_1008;
    90: op2_04_in02 = reg_1359;
    91: op2_04_in02 = reg_0890;
    92: op2_04_in02 = reg_0533;
    93: op2_04_in02 = reg_0645;
    128: op2_04_in02 = reg_0211;
    default: op2_04_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_04_in03 = reg_1478;
    74: op2_04_in03 = reg_1108;
    75: op2_04_in03 = reg_0533;
    88: op2_04_in03 = reg_1210;
    77: op2_04_in03 = reg_1073;
    78: op2_04_in03 = reg_0745;
    89: op2_04_in03 = reg_1274;
    79: op2_04_in03 = reg_1096;
    80: op2_04_in03 = reg_0581;
    81: op2_04_in03 = reg_1332;
    90: op2_04_in03 = reg_0935;
    91: op2_04_in03 = reg_0993;
    92: op2_04_in03 = reg_1050;
    93: op2_04_in03 = reg_0766;
    128: op2_04_in03 = reg_0343;
    default: op2_04_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_04_in04 = reg_0653;
    75: op2_04_in04 = reg_0211;
    88: op2_04_in04 = reg_1211;
    77: op2_04_in04 = reg_1112;
    78: op2_04_in04 = reg_0980;
    89: op2_04_in04 = reg_1102;
    79: op2_04_in04 = reg_0680;
    80: op2_04_in04 = reg_1127;
    81: op2_04_in04 = reg_0647;
    90: op2_04_in04 = reg_0083;
    91: op2_04_in04 = reg_0511;
    92: op2_04_in04 = reg_0865;
    93: op2_04_in04 = reg_1410;
    128: op2_04_in04 = reg_0668;
    default: op2_04_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の5番目の入力
  always @ ( * ) begin
    case ( state )
    75: op2_04_in05 = reg_1074;
    88: op2_04_in05 = reg_1246;
    89: op2_04_in05 = reg_0508;
    128: op2_04_in05 = reg_0815;
    default: op2_04_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#4の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_04_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#4のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_04_bias = 73;
    74: op2_04_bias = 60;
    75: op2_04_bias = 79;
    88: op2_04_bias = 86;
    77: op2_04_bias = 71;
    78: op2_04_bias = 65;
    89: op2_04_bias = 70;
    79: op2_04_bias = 70;
    80: op2_04_bias = 76;
    81: op2_04_bias = 69;
    90: op2_04_bias = 56;
    91: op2_04_bias = 56;
    92: op2_04_bias = 71;
    93: op2_04_bias = 77;
    128: op2_04_bias = 88;
    default: op2_04_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#5の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in00 = reg_0638;
    74: op2_05_in00 = reg_0721;
    88: op2_05_in00 = reg_1090;
    77: op2_05_in00 = reg_0594;
    89: op2_05_in00 = reg_1320;
    80: op2_05_in00 = reg_0535;
    81: op2_05_in00 = reg_1422;
    90: op2_05_in00 = reg_1360;
    91: op2_05_in00 = reg_0994;
    93: op2_05_in00 = reg_0511;
    default: op2_05_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in01 = reg_1030;
    74: op2_05_in01 = reg_1038;
    88: op2_05_in01 = reg_1247;
    77: op2_05_in01 = reg_0259;
    89: op2_05_in01 = reg_1275;
    80: op2_05_in01 = reg_1284;
    81: op2_05_in01 = reg_0909;
    90: op2_05_in01 = reg_1054;
    91: op2_05_in01 = reg_0509;
    93: op2_05_in01 = reg_1411;
    default: op2_05_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in02 = reg_1171;
    74: op2_05_in02 = reg_0960;
    88: op2_05_in02 = reg_0825;
    77: op2_05_in02 = reg_1102;
    89: op2_05_in02 = reg_0625;
    80: op2_05_in02 = reg_1464;
    81: op2_05_in02 = reg_0259;
    90: op2_05_in02 = reg_0655;
    91: op2_05_in02 = reg_0645;
    93: op2_05_in02 = reg_0888;
    default: op2_05_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in03 = reg_1443;
    74: op2_05_in03 = reg_0843;
    88: op2_05_in03 = reg_0721;
    77: op2_05_in03 = reg_0193;
    89: op2_05_in03 = reg_0793;
    80: op2_05_in03 = reg_1285;
    81: op2_05_in03 = reg_1042;
    90: op2_05_in03 = reg_0647;
    91: op2_05_in03 = reg_1007;
    93: op2_05_in03 = reg_0926;
    default: op2_05_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in04 = reg_0625;
    74: op2_05_in04 = reg_1109;
    88: op2_05_in04 = reg_1119;
    77: op2_05_in04 = reg_0823;
    89: op2_05_in04 = reg_1072;
    80: op2_05_in04 = reg_1128;
    81: op2_05_in04 = reg_0604;
    90: op2_05_in04 = reg_1361;
    91: op2_05_in04 = reg_1013;
    93: op2_05_in04 = reg_0686;
    default: op2_05_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の5番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in05 = reg_1172;
    89: op2_05_in05 = reg_1134;
    80: op2_05_in05 = reg_0354;
    81: op2_05_in05 = reg_0036;
    default: op2_05_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の6番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in06 = reg_1479;
    default: op2_05_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の7番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in07 = reg_1219;
    default: op2_05_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の8番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_in08 = reg_1086;
    default: op2_05_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#5の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_05_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#5のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_05_bias = 131;
    74: op2_05_bias = 74;
    88: op2_05_bias = 78;
    77: op2_05_bias = 77;
    89: op2_05_bias = 84;
    80: op2_05_bias = 70;
    81: op2_05_bias = 73;
    90: op2_05_bias = 69;
    91: op2_05_bias = 75;
    93: op2_05_bias = 70;
    default: op2_05_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#6の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_06_in00 = reg_1143;
    88: op2_06_in00 = reg_1316;
    77: op2_06_in00 = reg_1213;
    89: op2_06_in00 = reg_0728;
    80: op2_06_in00 = reg_1286;
    90: op2_06_in00 = reg_1238;
    91: op2_06_in00 = reg_0888;
    93: op2_06_in00 = reg_0634;
    default: op2_06_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_06_in01 = reg_0322;
    88: op2_06_in01 = reg_0910;
    77: op2_06_in01 = reg_0606;
    89: op2_06_in01 = reg_0911;
    80: op2_06_in01 = reg_1287;
    90: op2_06_in01 = reg_1362;
    91: op2_06_in01 = reg_0995;
    93: op2_06_in01 = reg_1051;
    default: op2_06_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_06_in02 = reg_0782;
    88: op2_06_in02 = reg_0826;
    90: op2_06_in02 = reg_0826;
    77: op2_06_in02 = reg_1005;
    89: op2_06_in02 = reg_1012;
    80: op2_06_in02 = reg_1465;
    91: op2_06_in02 = reg_1044;
    93: op2_06_in02 = reg_1059;
    default: op2_06_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_06_in03 = reg_1480;
    88: op2_06_in03 = reg_1248;
    77: op2_06_in03 = reg_0890;
    89: op2_06_in03 = reg_0782;
    80: op2_06_in03 = reg_1288;
    90: op2_06_in03 = reg_1363;
    91: op2_06_in03 = reg_0838;
    93: op2_06_in03 = reg_1412;
    default: op2_06_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_06_in04 = reg_1173;
    88: op2_06_in04 = reg_0761;
    89: op2_06_in04 = reg_1112;
    80: op2_06_in04 = reg_1058;
    90: op2_06_in04 = reg_1008;
    91: op2_06_in04 = reg_0766;
    93: op2_06_in04 = reg_1061;
    default: op2_06_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の5番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_06_in05 = reg_1191;
    89: op2_06_in05 = reg_0606;
    80: op2_06_in05 = reg_0502;
    90: op2_06_in05 = reg_0358;
    default: op2_06_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の6番目の入力
  always @ ( * ) begin
    case ( state )
    89: op2_06_in06 = reg_1135;
    default: op2_06_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#6の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_06_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#6のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_06_bias = 67;
    88: op2_06_bias = 75;
    77: op2_06_bias = 68;
    89: op2_06_bias = 107;
    80: op2_06_bias = 76;
    90: op2_06_bias = 87;
    91: op2_06_bias = 58;
    93: op2_06_bias = 78;
    default: op2_06_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#7の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_07_in00 = reg_0676;
    88: op2_07_in00 = reg_1249;
    89: op2_07_in00 = reg_0670;
    80: op2_07_in00 = reg_0563;
    90: op2_07_in00 = reg_0259;
    91: op2_07_in00 = reg_0998;
    default: op2_07_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_07_in01 = reg_1174;
    88: op2_07_in01 = reg_1011;
    89: op2_07_in01 = reg_0713;
    80: op2_07_in01 = reg_1129;
    90: op2_07_in01 = reg_1364;
    91: op2_07_in01 = reg_1150;
    default: op2_07_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_07_in02 = reg_1125;
    88: op2_07_in02 = reg_1332;
    89: op2_07_in02 = reg_1118;
    80: op2_07_in02 = reg_1466;
    90: op2_07_in02 = reg_1067;
    91: op2_07_in02 = reg_0634;
    default: op2_07_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_07_in03 = reg_1175;
    88: op2_07_in03 = reg_0843;
    89: op2_07_in03 = reg_1276;
    80: op2_07_in03 = reg_1289;
    90: op2_07_in03 = reg_0446;
    91: op2_07_in03 = reg_1059;
    default: op2_07_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_07_in04 = reg_0942;
    88: op2_07_in04 = reg_0762;
    89: op2_07_in04 = reg_0671;
    80: op2_07_in04 = reg_1213;
    90: op2_07_in04 = reg_1167;
    91: op2_07_in04 = reg_1394;
    default: op2_07_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の5番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_07_in05 = reg_1220;
    89: op2_07_in05 = reg_1136;
    80: op2_07_in05 = reg_0355;
    90: op2_07_in05 = reg_0510;
    default: op2_07_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#7の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_07_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#7のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_07_bias = 87;
    88: op2_07_bias = 53;
    89: op2_07_bias = 69;
    80: op2_07_bias = 78;
    90: op2_07_bias = 92;
    91: op2_07_bias = 63;
    default: op2_07_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#8の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_08_in00 = reg_1144;
    88: op2_08_in00 = reg_0705;
    89: op2_08_in00 = reg_0074;
    90: op2_08_in00 = reg_0650;
    91: op2_08_in00 = reg_1395;
    default: op2_08_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_08_in01 = reg_1116;
    88: op2_08_in01 = reg_1120;
    89: op2_08_in01 = reg_1295;
    90: op2_08_in01 = reg_1327;
    91: op2_08_in01 = reg_1396;
    default: op2_08_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_08_in02 = reg_1007;
    89: op2_08_in02 = reg_1007;
    88: op2_08_in02 = reg_0503;
    90: op2_08_in02 = reg_0503;
    91: op2_08_in02 = reg_0556;
    default: op2_08_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_08_in03 = reg_1497;
    88: op2_08_in03 = reg_1250;
    89: op2_08_in03 = reg_0645;
    90: op2_08_in03 = reg_0850;
    91: op2_08_in03 = reg_0946;
    default: op2_08_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の4番目の入力
  always @ ( * ) begin
    case ( state )
    88: op2_08_in04 = reg_1153;
    89: op2_08_in04 = reg_1296;
    90: op2_08_in04 = reg_1365;
    91: op2_08_in04 = reg_0606;
    default: op2_08_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の5番目の入力
  always @ ( * ) begin
    case ( state )
    88: op2_08_in05 = reg_0683;
    91: op2_08_in05 = reg_1397;
    default: op2_08_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#8の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_08_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#8のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_08_bias = 59;
    88: op2_08_bias = 82;
    89: op2_08_bias = 82;
    90: op2_08_bias = 73;
    91: op2_08_bias = 83;
    default: op2_08_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#9の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_09_in00 = reg_1481;
    88: op2_09_in00 = reg_1294;
    89: op2_09_in00 = reg_0912;
    90: op2_09_in00 = reg_1366;
    default: op2_09_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_09_in01 = reg_1117;
    88: op2_09_in01 = reg_1251;
    89: op2_09_in01 = reg_1297;
    90: op2_09_in01 = reg_0705;
    default: op2_09_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_09_in02 = reg_1043;
    89: op2_09_in02 = reg_1043;
    88: op2_09_in02 = reg_0871;
    90: op2_09_in02 = reg_0355;
    default: op2_09_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_09_in03 = reg_1498;
    88: op2_09_in03 = reg_0977;
    89: op2_09_in03 = reg_1046;
    90: op2_09_in03 = reg_0682;
    default: op2_09_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_09_in04 = reg_1221;
    88: op2_09_in04 = reg_1121;
    89: op2_09_in04 = reg_1137;
    default: op2_09_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の5番目の入力
  always @ ( * ) begin
    case ( state )
    88: op2_09_in05 = reg_0654;
    89: op2_09_in05 = reg_0082;
    default: op2_09_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#9の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_09_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#9のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_09_bias = 85;
    88: op2_09_bias = 78;
    89: op2_09_bias = 72;
    90: op2_09_bias = 53;
    default: op2_09_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#10の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_10_in00 = reg_1482;
    88: op2_10_in00 = reg_1317;
    89: op2_10_in00 = reg_0226;
    90: op2_10_in00 = reg_0502;
    default: op2_10_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_10_in01 = reg_1176;
    88: op2_10_in01 = reg_1252;
    89: op2_10_in01 = reg_1308;
    90: op2_10_in01 = reg_1015;
    default: op2_10_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_10_in02 = reg_0893;
    88: op2_10_in02 = reg_1427;
    89: op2_10_in02 = reg_0888;
    90: op2_10_in02 = reg_0150;
    default: op2_10_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_10_in03 = reg_1222;
    88: op2_10_in03 = reg_0652;
    89: op2_10_in03 = reg_1013;
    90: op2_10_in03 = reg_0376;
    default: op2_10_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_10_in04 = reg_1499;
    88: op2_10_in04 = reg_1187;
    89: op2_10_in04 = reg_1309;
    90: op2_10_in04 = reg_0731;
    default: op2_10_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の5番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_10_in05 = reg_1087;
    88: op2_10_in05 = reg_1089;
    default: op2_10_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#10の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_10_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#10のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_10_bias = 94;
    88: op2_10_bias = 92;
    89: op2_10_bias = 68;
    90: op2_10_bias = 73;
    default: op2_10_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#11の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_11_in00 = reg_0677;
    88: op2_11_in00 = reg_1318;
    89: op2_11_in00 = reg_1310;
    90: op2_11_in00 = reg_1127;
    default: op2_11_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_11_in01 = reg_1444;
    88: op2_11_in01 = reg_1138;
    89: op2_11_in01 = reg_1044;
    90: op2_11_in01 = reg_1057;
    default: op2_11_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_11_in02 = reg_1044;
    88: op2_11_in02 = reg_0926;
    90: op2_11_in02 = reg_0926;
    89: op2_11_in02 = reg_1311;
    default: op2_11_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_11_in03 = reg_0634;
    88: op2_11_in03 = reg_0533;
    89: op2_11_in03 = reg_0603;
    90: op2_11_in03 = reg_1148;
    default: op2_11_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_11_in04 = reg_1500;
    88: op2_11_in04 = reg_0266;
    89: op2_11_in04 = reg_0509;
    90: op2_11_in04 = reg_1370;
    default: op2_11_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の5番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_11_in05 = reg_0200;
    default: op2_11_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#11の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_11_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#11のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_11_bias = 84;
    88: op2_11_bias = 48;
    89: op2_11_bias = 61;
    90: op2_11_bias = 66;
    default: op2_11_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#12の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_12_in00 = reg_1177;
    88: op2_12_in00 = reg_0732;
    89: op2_12_in00 = reg_1232;
    90: op2_12_in00 = reg_1061;
    default: op2_12_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_12_in01 = reg_1192;
    88: op2_12_in01 = reg_0193;
    89: op2_12_in01 = reg_1335;
    90: op2_12_in01 = reg_1113;
    default: op2_12_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_12_in02 = reg_1058;
    88: op2_12_in02 = reg_0367;
    89: op2_12_in02 = reg_0634;
    90: op2_12_in02 = reg_0732;
    default: op2_12_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_12_in03 = reg_1002;
    88: op2_12_in03 = reg_1261;
    89: op2_12_in03 = reg_0945;
    90: op2_12_in03 = reg_0036;
    default: op2_12_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_12_in04 = reg_0628;
    89: op2_12_in04 = reg_1073;
    90: op2_12_in04 = reg_0764;
    default: op2_12_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の5番目の入力
  always @ ( * ) begin
    case ( state )
    89: op2_12_in05 = reg_0685;
    default: op2_12_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#12の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_12_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#12のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_12_bias = 79;
    88: op2_12_bias = 63;
    89: op2_12_bias = 83;
    90: op2_12_bias = 65;
    default: op2_12_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#13の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_13_in00 = reg_1118;
    88: op2_13_in00 = reg_0756;
    89: op2_13_in00 = reg_1111;
    90: op2_13_in00 = reg_1236;
    default: op2_13_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_13_in01 = reg_1193;
    88: op2_13_in01 = reg_1262;
    89: op2_13_in01 = reg_1223;
    90: op2_13_in01 = reg_0639;
    default: op2_13_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_13_in02 = reg_1445;
    88: op2_13_in02 = reg_1009;
    89: op2_13_in02 = reg_1059;
    90: op2_13_in02 = reg_0533;
    default: op2_13_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_13_in03 = reg_1423;
    88: op2_13_in03 = reg_0944;
    89: op2_13_in03 = reg_0556;
    90: op2_13_in03 = reg_0076;
    default: op2_13_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_13_in04 = reg_0062;
    88: op2_13_in04 = reg_1263;
    89: op2_13_in04 = reg_1336;
    90: op2_13_in04 = reg_1371;
    default: op2_13_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の5番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_13_in05 = reg_1223;
    88: op2_13_in05 = reg_0081;
    default: op2_13_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#13の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_13_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#13のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_13_bias = 93;
    88: op2_13_bias = 85;
    89: op2_13_bias = 62;
    90: op2_13_bias = 69;
    default: op2_13_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#14の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_14_in00 = reg_0792;
    88: op2_14_in00 = reg_0985;
    89: op2_14_in00 = reg_1337;
    90: op2_14_in00 = reg_1385;
    default: op2_14_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_14_in01 = reg_1194;
    88: op2_14_in01 = reg_1264;
    89: op2_14_in01 = reg_1213;
    90: op2_14_in01 = reg_1386;
    default: op2_14_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_14_in02 = reg_1213;
    88: op2_14_in02 = reg_1161;
    89: op2_14_in02 = reg_1162;
    90: op2_14_in02 = reg_0721;
    default: op2_14_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_14_in03 = reg_1010;
    88: op2_14_in03 = reg_0164;
    89: op2_14_in03 = reg_1060;
    90: op2_14_in03 = reg_0867;
    default: op2_14_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_14_in04 = reg_1224;
    88: op2_14_in04 = reg_1265;
    89: op2_14_in04 = reg_0265;
    default: op2_14_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の5番目の入力
  always @ ( * ) begin
    case ( state )
    88: op2_14_in05 = reg_1266;
    default: op2_14_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#14の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_14_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#14のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_14_bias = 70;
    88: op2_14_bias = 79;
    89: op2_14_bias = 69;
    90: op2_14_bias = 60;
    default: op2_14_bias = 0;
    endcase
  end // always @ ( * )

  // OP2#15の0番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_15_in00 = reg_1145;
    88: op2_15_in00 = reg_1185;
    90: op2_15_in00 = reg_0651;
    default: op2_15_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の1番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_15_in01 = reg_0931;
    88: op2_15_in01 = reg_1472;
    90: op2_15_in01 = reg_1158;
    default: op2_15_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の2番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_15_in02 = reg_1162;
    88: op2_15_in02 = reg_1131;
    90: op2_15_in02 = reg_0843;
    default: op2_15_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の3番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_15_in03 = reg_0943;
    88: op2_15_in03 = reg_1152;
    90: op2_15_in03 = reg_1047;
    default: op2_15_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の4番目の入力
  always @ ( * ) begin
    case ( state )
    87: op2_15_in04 = reg_0888;
    88: op2_15_in04 = reg_1267;
    90: op2_15_in04 = reg_0854;
    default: op2_15_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の5番目の入力
  always @ ( * ) begin
    case ( state )
    88: op2_15_in05 = reg_0655;
    default: op2_15_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の15番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in15 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の16番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in16 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の17番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in17 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の18番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in18 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の19番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in19 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の20番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in20 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の21番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in21 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の22番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in22 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の23番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in23 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の24番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in24 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の25番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in25 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の26番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in26 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の27番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in27 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の28番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in28 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の29番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in29 = 0;
    endcase
  end // always @ ( * )

  // OP2#15の30番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_15_in30 = 0;
    endcase
  end // always @ ( * )

  // OP2#15のバイアス入力
  always @ ( * ) begin
    case ( state )
    87: op2_15_bias = 84;
    88: op2_15_bias = 93;
    90: op2_15_bias = 75;
    default: op2_15_bias = 0;
    endcase
  end // always @ ( * )

  // REG#0の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0000 <= imem03_in[3:0];
    21: reg_0000 <= imem03_in[3:0];
    40: reg_0000 <= imem03_in[3:0];
    58: reg_0000 <= imem03_in[3:0];
    endcase
  end

  // REG#1の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0001 <= imem07_in[3:0];
    30: reg_0001 <= imem07_in[3:0];
    endcase
  end

  // REG#2の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0002 <= imem07_in[7:4];
    30: reg_0002 <= imem07_in[7:4];
    127: reg_0002 <= imem07_in[7:4];
    endcase
  end

  // REG#3の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0003 <= imem07_in[15:12];
    31: reg_0003 <= imem07_in[15:12];
    111: reg_0003 <= imem07_in[15:12];
    endcase
  end

  // REG#4の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0004 <= imem07_in[11:8];
    31: reg_0004 <= imem07_in[11:8];
    119: reg_0004 <= imem07_in[11:8];
    127: reg_0004 <= imem07_in[11:8];
    endcase
  end

  // REG#5の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0005 <= imem00_in[3:0];
    43: reg_0005 <= imem00_in[3:0];
    130: reg_0005 <= imem00_in[3:0];
    endcase
  end

  // REG#6の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0006 <= imem02_in[15:12];
    65: reg_0006 <= imem02_in[15:12];
    82: reg_0006 <= imem02_in[15:12];
    endcase
  end

  // REG#7の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0007 <= imem02_in[7:4];
    66: reg_0007 <= imem02_in[7:4];
    107: reg_0007 <= imem02_in[7:4];
    endcase
  end

  // REG#8の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0008 <= imem02_in[11:8];
    66: reg_0008 <= imem02_in[11:8];
    108: reg_0008 <= imem02_in[11:8];
    111: reg_0008 <= imem02_in[11:8];
    116: reg_0008 <= imem02_in[11:8];
    118: reg_0008 <= imem02_in[11:8];
    126: reg_0008 <= imem02_in[11:8];
    131: reg_0008 <= imem02_in[11:8];
    endcase
  end

  // REG#9の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0009 <= imem02_in[3:0];
    67: reg_0009 <= imem02_in[3:0];
    83: reg_0009 <= imem02_in[3:0];
    129: reg_0009 <= imem02_in[3:0];
    endcase
  end

  // REG#10の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0010 <= imem01_in[11:8];
    105: reg_0010 <= imem01_in[11:8];
    107: reg_0010 <= imem01_in[11:8];
    109: reg_0010 <= imem01_in[11:8];
    114: reg_0010 <= imem01_in[11:8];
    129: reg_0010 <= imem01_in[11:8];
    131: reg_0010 <= imem01_in[11:8];
    endcase
  end

  // REG#11の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0011 <= imem01_in[7:4];
    106: reg_0011 <= imem01_in[7:4];
    111: reg_0011 <= imem01_in[7:4];
    114: reg_0011 <= imem01_in[7:4];
    endcase
  end

  // REG#12の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0012 <= imem01_in[3:0];
    106: reg_0012 <= imem01_in[3:0];
    114: reg_0012 <= imem01_in[3:0];
    endcase
  end

  // REG#13の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0013 <= imem01_in[15:12];
    106: reg_0013 <= imem01_in[15:12];
    111: reg_0013 <= imem01_in[15:12];
    116: reg_0013 <= op2_01_out;
    118: reg_0013 <= op2_01_out;
    126: reg_0013 <= imem01_in[15:12];
    132: reg_0013 <= op2_01_out;
    endcase
  end

  // REG#14の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0014 <= imem05_in[3:0];
    115: reg_0014 <= imem05_in[3:0];
    endcase
  end

  // REG#15の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0015 <= imem06_in[3:0];
    123: reg_0015 <= op2_00_out;
    endcase
  end

  // REG#16の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0016 <= imem04_in[7:4];
    124: reg_0016 <= imem04_in[7:4];
    endcase
  end

  // REG#17の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0017 <= imem06_in[15:12];
    endcase
  end

  // REG#18の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0018 <= imem06_in[7:4];
    131: reg_0018 <= imem06_in[7:4];
    endcase
  end

  // REG#19の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0019 <= imem04_in[3:0];
    endcase
  end

  // REG#20の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0020 <= imem04_in[15:12];
    endcase
  end

  // REG#21の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0021 <= imem04_in[11:8];
    131: reg_0021 <= imem04_in[11:8];
    endcase
  end

  // REG#22の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0022 <= imem06_in[11:8];
    endcase
  end

  // REG#23の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0023 <= imem06_in[7:4];
    13: reg_0023 <= imem06_in[7:4];
    endcase
  end

  // REG#24の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0024 <= imem02_in[3:0];
    17: reg_0024 <= imem02_in[3:0];
    endcase
  end

  // REG#25の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0025 <= imem03_in[3:0];
    21: reg_0025 <= imem07_in[11:8];
    23: reg_0025 <= imem03_in[3:0];
    62: reg_0025 <= imem07_in[11:8];
    86: reg_0025 <= imem03_in[3:0];
    129: reg_0025 <= imem07_in[11:8];
    endcase
  end

  // REG#26の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0026 <= imem00_in[11:8];
    22: reg_0026 <= imem00_in[11:8];
    130: reg_0026 <= imem00_in[11:8];
    endcase
  end

  // REG#27の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0027 <= imem00_in[15:12];
    22: reg_0027 <= imem00_in[15:12];
    endcase
  end

  // REG#28の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0028 <= imem07_in[7:4];
    23: reg_0028 <= imem07_in[7:4];
    endcase
  end

  // REG#29の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0029 <= imem07_in[11:8];
    24: reg_0029 <= imem07_in[11:8];
    27: reg_0029 <= imem07_in[11:8];
    128: reg_0029 <= imem07_in[11:8];
    endcase
  end

  // REG#30の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0030 <= imem07_in[15:12];
    24: reg_0030 <= imem07_in[15:12];
    27: reg_0030 <= imem07_in[15:12];
    endcase
  end

  // REG#31の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0031 <= imem07_in[3:0];
    24: reg_0031 <= imem07_in[3:0];
    27: reg_0031 <= imem07_in[3:0];
    endcase
  end

  // REG#32の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0032 <= imem04_in[3:0];
    65: reg_0032 <= imem04_in[3:0];
    113: reg_0032 <= imem04_in[3:0];
    128: reg_0032 <= imem04_in[3:0];
    endcase
  end

  // REG#33の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0033 <= imem04_in[7:4];
    70: reg_0033 <= imem04_in[7:4];
    79: reg_0033 <= imem04_in[7:4];
    endcase
  end

  // REG#34の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0034 <= imem04_in[15:12];
    72: reg_0034 <= imem07_in[3:0];
    74: reg_0034 <= imem07_in[3:0];
    78: reg_0034 <= imem07_in[3:0];
    86: reg_0034 <= imem04_in[15:12];
    122: reg_0034 <= imem07_in[3:0];
    124: reg_0034 <= imem07_in[3:0];
    127: reg_0034 <= imem04_in[15:12];
    endcase
  end

  // REG#35の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0035 <= imem04_in[11:8];
    73: reg_0035 <= imem04_in[11:8];
    130: reg_0035 <= imem04_in[11:8];
    endcase
  end

  // REG#36の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0036 <= op1_00_out;
    82: reg_0036 <= op1_00_out;
    84: reg_0036 <= op1_00_out;
    91: reg_0036 <= op1_00_out;
    93: reg_0036 <= op1_00_out;
    95: reg_0036 <= op1_00_out;
    97: reg_0036 <= op1_00_out;
    99: reg_0036 <= op1_00_out;
    101: reg_0036 <= op1_00_out;
    103: reg_0036 <= op1_00_out;
    105: reg_0036 <= op1_00_out;
    107: reg_0036 <= op1_00_out;
    109: reg_0036 <= op1_00_out;
    111: reg_0036 <= op1_00_out;
    113: reg_0036 <= op1_00_out;
    115: reg_0036 <= op1_00_out;
    117: reg_0036 <= op1_00_out;
    119: reg_0036 <= op1_00_out;
    121: reg_0036 <= op1_00_out;
    123: reg_0036 <= op1_00_out;
    125: reg_0036 <= op1_00_out;
    127: reg_0036 <= op1_00_out;
    129: reg_0036 <= op1_00_out;
    131: reg_0036 <= op1_00_out;
    endcase
  end

  // REG#37の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0037 <= imem05_in[3:0];
    111: reg_0037 <= op2_00_out;
    endcase
  end

  // REG#38の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0038 <= imem05_in[7:4];
    113: reg_0038 <= imem05_in[7:4];
    124: reg_0038 <= imem05_in[7:4];
    126: reg_0038 <= imem05_in[7:4];
    129: reg_0038 <= imem05_in[7:4];
    endcase
  end

  // REG#39の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0039 <= imem05_in[15:12];
    115: reg_0039 <= imem05_in[15:12];
    endcase
  end

  // REG#40の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0040 <= imem05_in[11:8];
    116: reg_0040 <= imem05_in[11:8];
    119: reg_0040 <= imem05_in[11:8];
    endcase
  end

  // REG#41の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0041 <= imem01_in[15:12];
    endcase
  end

  // REG#42の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0042 <= imem01_in[7:4];
    endcase
  end

  // REG#43の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0043 <= imem01_in[3:0];
    endcase
  end

  // REG#44の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0044 <= imem01_in[11:8];
    endcase
  end

  // REG#45の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0045 <= imem05_in[11:8];
    13: reg_0045 <= imem05_in[11:8];
    55: reg_0045 <= imem05_in[11:8];
    78: reg_0045 <= imem05_in[11:8];
    81: reg_0045 <= imem05_in[11:8];
    endcase
  end

  // REG#46の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0046 <= imem06_in[11:8];
    13: reg_0046 <= imem06_in[11:8];
    endcase
  end

  // REG#47の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0047 <= imem01_in[7:4];
    17: reg_0047 <= imem01_in[7:4];
    22: reg_0047 <= imem01_in[7:4];
    44: reg_0047 <= imem01_in[7:4];
    69: reg_0047 <= imem01_in[7:4];
    128: reg_0047 <= imem01_in[7:4];
    endcase
  end

  // REG#48の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0048 <= imem03_in[7:4];
    21: reg_0048 <= imem03_in[7:4];
    40: reg_0048 <= imem03_in[7:4];
    60: reg_0048 <= imem03_in[7:4];
    120: reg_0048 <= imem03_in[7:4];
    126: reg_0048 <= imem03_in[7:4];
    128: reg_0048 <= imem03_in[7:4];
    130: reg_0048 <= imem03_in[7:4];
    endcase
  end

  // REG#49の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0049 <= imem03_in[11:8];
    20: reg_0049 <= op1_00_out;
    23: reg_0049 <= imem03_in[11:8];
    61: reg_0049 <= op1_00_out;
    70: reg_0049 <= imem03_in[11:8];
    102: reg_0049 <= imem03_in[11:8];
    endcase
  end

  // REG#50の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0050 <= imem07_in[3:0];
    31: reg_0050 <= imem07_in[3:0];
    115: reg_0050 <= imem07_in[3:0];
    121: reg_0050 <= imem07_in[3:0];
    125: reg_0050 <= imem07_in[3:0];
    endcase
  end

  // REG#51の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0051 <= imem07_in[7:4];
    31: reg_0051 <= imem07_in[7:4];
    116: reg_0051 <= imem07_in[7:4];
    123: reg_0051 <= imem07_in[7:4];
    130: reg_0051 <= imem07_in[7:4];
    endcase
  end

  // REG#52の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0052 <= imem07_in[11:8];
    30: reg_0052 <= imem07_in[11:8];
    endcase
  end

  // REG#53の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0053 <= imem07_in[15:12];
    30: reg_0053 <= imem07_in[15:12];
    endcase
  end

  // REG#54の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0054 <= imem02_in[3:0];
    38: reg_0054 <= imem02_in[3:0];
    127: reg_0054 <= imem02_in[3:0];
    endcase
  end

  // REG#55の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0055 <= imem02_in[15:12];
    44: reg_0055 <= imem02_in[15:12];
    71: reg_0055 <= imem02_in[15:12];
    endcase
  end

  // REG#56の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0056 <= imem02_in[7:4];
    44: reg_0056 <= imem02_in[7:4];
    72: reg_0056 <= imem02_in[7:4];
    endcase
  end

  // REG#57の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0057 <= imem00_in[7:4];
    62: reg_0057 <= imem00_in[7:4];
    endcase
  end

  // REG#58の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0058 <= imem00_in[15:12];
    63: reg_0058 <= imem00_in[15:12];
    131: reg_0058 <= imem00_in[15:12];
    endcase
  end

  // REG#59の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0059 <= imem00_in[11:8];
    63: reg_0059 <= imem00_in[11:8];
    124: reg_0059 <= imem00_in[11:8];
    126: reg_0059 <= imem00_in[11:8];
    endcase
  end

  // REG#60の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0060 <= imem00_in[3:0];
    63: reg_0060 <= imem00_in[3:0];
    endcase
  end

  // REG#61の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0061 <= imem04_in[15:12];
    70: reg_0061 <= imem04_in[15:12];
    79: reg_0061 <= imem04_in[15:12];
    endcase
  end

  // REG#62の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0062 <= imem04_in[11:8];
    72: reg_0062 <= op1_03_out;
    74: reg_0062 <= op1_03_out;
    89: reg_0062 <= imem04_in[11:8];
    92: reg_0062 <= op1_03_out;
    95: reg_0062 <= imem04_in[11:8];
    endcase
  end

  // REG#63の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0063 <= imem04_in[7:4];
    75: reg_0063 <= imem04_in[7:4];
    130: reg_0063 <= imem04_in[7:4];
    endcase
  end

  // REG#64の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0064 <= imem04_in[3:0];
    75: reg_0064 <= imem04_in[3:0];
    endcase
  end

  // REG#65の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0065 <= imem04_in[11:8];
    13: reg_0065 <= imem04_in[11:8];
    71: reg_0065 <= imem07_in[7:4];
    75: reg_0065 <= imem04_in[11:8];
    endcase
  end

  // REG#66の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0066 <= imem05_in[3:0];
    13: reg_0066 <= imem05_in[3:0];
    56: reg_0066 <= imem05_in[3:0];
    83: reg_0066 <= imem05_in[3:0];
    127: reg_0066 <= imem05_in[3:0];
    endcase
  end

  // REG#67の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0067 <= imem06_in[3:0];
    13: reg_0067 <= imem06_in[3:0];
    endcase
  end

  // REG#68の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0068 <= imem02_in[7:4];
    17: reg_0068 <= imem02_in[7:4];
    endcase
  end

  // REG#69の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0069 <= imem02_in[15:12];
    17: reg_0069 <= imem02_in[15:12];
    endcase
  end

  // REG#70の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0070 <= imem03_in[3:0];
    21: reg_0070 <= imem05_in[7:4];
    28: reg_0070 <= imem05_in[7:4];
    75: reg_0070 <= imem03_in[3:0];
    endcase
  end

  // REG#71の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0071 <= imem00_in[3:0];
    64: reg_0071 <= imem00_in[3:0];
    endcase
  end

  // REG#72の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0072 <= imem00_in[7:4];
    63: reg_0072 <= imem00_in[7:4];
    endcase
  end

  // REG#73の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0073 <= imem00_in[11:8];
    64: reg_0073 <= imem00_in[11:8];
    endcase
  end

  // REG#74の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0074 <= op1_00_out;
    62: reg_0074 <= op1_00_out;
    90: reg_0074 <= op1_00_out;
    92: reg_0074 <= op1_00_out;
    94: reg_0074 <= op1_00_out;
    96: reg_0074 <= op1_00_out;
    98: reg_0074 <= op1_00_out;
    100: reg_0074 <= op1_00_out;
    102: reg_0074 <= op1_00_out;
    104: reg_0074 <= op1_00_out;
    106: reg_0074 <= op1_00_out;
    108: reg_0074 <= op1_00_out;
    110: reg_0074 <= op1_00_out;
    112: reg_0074 <= op1_00_out;
    114: reg_0074 <= op1_00_out;
    116: reg_0074 <= op1_00_out;
    118: reg_0074 <= op1_00_out;
    120: reg_0074 <= op1_00_out;
    122: reg_0074 <= op1_00_out;
    124: reg_0074 <= op1_00_out;
    126: reg_0074 <= op1_00_out;
    128: reg_0074 <= op1_00_out;
    130: reg_0074 <= op1_00_out;
    endcase
  end

  // REG#75の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0075 <= imem00_in[15:12];
    64: reg_0075 <= imem00_in[15:12];
    129: reg_0075 <= imem00_in[15:12];
    endcase
  end

  // REG#76の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0076 <= op1_03_out;
    82: reg_0076 <= op1_03_out;
    84: reg_0076 <= op1_03_out;
    91: reg_0076 <= op1_03_out;
    93: reg_0076 <= op1_03_out;
    95: reg_0076 <= op1_03_out;
    97: reg_0076 <= op1_03_out;
    99: reg_0076 <= op1_03_out;
    101: reg_0076 <= op1_03_out;
    103: reg_0076 <= op1_03_out;
    105: reg_0076 <= op1_03_out;
    107: reg_0076 <= op1_03_out;
    109: reg_0076 <= op1_03_out;
    111: reg_0076 <= op1_03_out;
    113: reg_0076 <= op1_03_out;
    115: reg_0076 <= op1_03_out;
    117: reg_0076 <= op1_03_out;
    119: reg_0076 <= op1_03_out;
    121: reg_0076 <= op1_03_out;
    123: reg_0076 <= op1_03_out;
    125: reg_0076 <= op1_03_out;
    127: reg_0076 <= op1_03_out;
    129: reg_0076 <= op1_03_out;
    131: reg_0076 <= op1_03_out;
    endcase
  end

  // REG#77の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0077 <= imem01_in[11:8];
    86: reg_0077 <= imem01_in[11:8];
    endcase
  end

  // REG#78の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0078 <= imem01_in[7:4];
    86: reg_0078 <= imem01_in[7:4];
    126: reg_0078 <= imem01_in[7:4];
    endcase
  end

  // REG#79の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0079 <= imem01_in[15:12];
    86: reg_0079 <= imem01_in[15:12];
    endcase
  end

  // REG#80の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0080 <= imem01_in[3:0];
    86: reg_0080 <= imem01_in[3:0];
    endcase
  end

  // REG#81の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0081 <= op1_01_out;
    89: reg_0081 <= op1_01_out;
    91: reg_0081 <= op1_01_out;
    93: reg_0081 <= op1_01_out;
    95: reg_0081 <= op1_01_out;
    97: reg_0081 <= op1_01_out;
    99: reg_0081 <= op1_01_out;
    101: reg_0081 <= op1_01_out;
    103: reg_0081 <= op1_01_out;
    105: reg_0081 <= op1_01_out;
    107: reg_0081 <= op1_01_out;
    109: reg_0081 <= op1_01_out;
    111: reg_0081 <= op1_01_out;
    113: reg_0081 <= op1_01_out;
    115: reg_0081 <= op1_01_out;
    117: reg_0081 <= op1_01_out;
    119: reg_0081 <= op1_01_out;
    121: reg_0081 <= op1_01_out;
    123: reg_0081 <= op1_01_out;
    125: reg_0081 <= op1_01_out;
    127: reg_0081 <= op1_01_out;
    129: reg_0081 <= op1_01_out;
    131: reg_0081 <= op1_01_out;
    endcase
  end

  // REG#82の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0082 <= op1_02_out;
    90: reg_0082 <= op1_02_out;
    92: reg_0082 <= op1_02_out;
    94: reg_0082 <= op1_02_out;
    96: reg_0082 <= op1_02_out;
    98: reg_0082 <= op1_02_out;
    100: reg_0082 <= op1_02_out;
    102: reg_0082 <= op1_02_out;
    104: reg_0082 <= op1_02_out;
    106: reg_0082 <= op1_02_out;
    108: reg_0082 <= op1_02_out;
    110: reg_0082 <= op1_02_out;
    112: reg_0082 <= op1_02_out;
    114: reg_0082 <= op1_02_out;
    116: reg_0082 <= op1_02_out;
    118: reg_0082 <= op1_02_out;
    120: reg_0082 <= op1_02_out;
    122: reg_0082 <= op1_02_out;
    124: reg_0082 <= op1_02_out;
    126: reg_0082 <= op1_02_out;
    128: reg_0082 <= op1_02_out;
    130: reg_0082 <= op1_02_out;
    endcase
  end

  // REG#83の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0083 <= op1_04_out;
    91: reg_0083 <= op1_04_out;
    93: reg_0083 <= op1_04_out;
    95: reg_0083 <= op1_04_out;
    97: reg_0083 <= op1_04_out;
    99: reg_0083 <= op1_04_out;
    101: reg_0083 <= op1_04_out;
    103: reg_0083 <= op1_04_out;
    105: reg_0083 <= op1_04_out;
    107: reg_0083 <= op1_04_out;
    109: reg_0083 <= op1_04_out;
    111: reg_0083 <= op1_04_out;
    113: reg_0083 <= op1_04_out;
    115: reg_0083 <= op1_04_out;
    117: reg_0083 <= op1_04_out;
    119: reg_0083 <= op1_04_out;
    121: reg_0083 <= op1_04_out;
    123: reg_0083 <= op1_04_out;
    125: reg_0083 <= op1_04_out;
    127: reg_0083 <= op1_04_out;
    129: reg_0083 <= op1_04_out;
    131: reg_0083 <= op1_04_out;
    endcase
  end

  // REG#84の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0084 <= imem07_in[11:8];
    110: reg_0084 <= imem07_in[11:8];
    113: reg_0084 <= imem07_in[11:8];
    endcase
  end

  // REG#85の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0085 <= imem07_in[3:0];
    119: reg_0085 <= imem07_in[3:0];
    endcase
  end

  // REG#86の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0086 <= imem07_in[7:4];
    119: reg_0086 <= imem07_in[7:4];
    endcase
  end

  // REG#87の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0087 <= imem07_in[15:12];
    120: reg_0087 <= imem07_in[15:12];
    128: reg_0087 <= imem07_in[15:12];
    endcase
  end

  // REG#88の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0088 <= imem01_in[7:4];
    17: reg_0088 <= imem04_in[7:4];
    21: reg_0088 <= imem01_in[7:4];
    86: reg_0088 <= imem04_in[7:4];
    123: reg_0088 <= imem04_in[7:4];
    endcase
  end

  // REG#89の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0089 <= imem00_in[7:4];
    22: reg_0089 <= imem00_in[7:4];
    endcase
  end

  // REG#90の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0090 <= imem05_in[3:0];
    42: reg_0090 <= imem05_in[3:0];
    66: reg_0090 <= imem05_in[3:0];
    endcase
  end

  // REG#91の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0091 <= imem01_in[3:0];
    44: reg_0091 <= imem01_in[3:0];
    68: reg_0091 <= imem01_in[3:0];
    endcase
  end

  // REG#92の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0092 <= imem01_in[11:8];
    44: reg_0092 <= imem01_in[11:8];
    68: reg_0092 <= imem01_in[11:8];
    endcase
  end

  // REG#93の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0093 <= imem01_in[15:12];
    44: reg_0093 <= imem01_in[15:12];
    69: reg_0093 <= imem01_in[15:12];
    122: reg_0093 <= op2_00_out;
    endcase
  end

  // REG#94の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0094 <= imem04_in[7:4];
    71: reg_0094 <= imem04_in[7:4];
    82: reg_0094 <= imem04_in[7:4];
    endcase
  end

  // REG#95の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0095 <= imem04_in[15:12];
    75: reg_0095 <= imem04_in[15:12];
    endcase
  end

  // REG#96の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0096 <= imem04_in[11:8];
    78: reg_0096 <= imem04_in[11:8];
    endcase
  end

  // REG#97の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0097 <= imem04_in[3:0];
    79: reg_0097 <= imem04_in[3:0];
    endcase
  end

  // REG#98の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0098 <= op1_00_out;
    111: reg_0098 <= op2_02_out;
    endcase
  end

  // REG#99の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0099 <= op1_01_out;
    116: reg_0099 <= imem02_in[7:4];
    122: reg_0099 <= imem02_in[7:4];
    124: reg_0099 <= op1_01_out;
    126: reg_0099 <= op1_01_out;
    128: reg_0099 <= op1_01_out;
    130: reg_0099 <= op1_01_out;
    endcase
  end

  // REG#100の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0100 <= imem07_in[11:8];
    118: reg_0100 <= op2_00_out;
    125: reg_0100 <= imem07_in[11:8];
    132: reg_0100 <= op2_00_out;
    endcase
  end

  // REG#101の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0101 <= op1_02_out;
    123: reg_0101 <= op1_02_out;
    125: reg_0101 <= op1_02_out;
    127: reg_0101 <= op1_02_out;
    129: reg_0101 <= op1_02_out;
    131: reg_0101 <= op1_02_out;
    endcase
  end

  // REG#102の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0102 <= imem07_in[3:0];
    124: reg_0102 <= op2_01_out;
    endcase
  end

  // REG#103の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0103 <= imem07_in[7:4];
    128: reg_0103 <= imem07_in[7:4];
    endcase
  end

  // REG#104の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0104 <= imem03_in[15:12];
    129: reg_0104 <= imem03_in[15:12];
    endcase
  end

  // REG#105の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0105 <= imem02_in[15:12];
    130: reg_0105 <= imem02_in[15:12];
    endcase
  end

  // REG#106の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0106 <= imem02_in[11:8];
    endcase
  end

  // REG#107の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0107 <= imem03_in[7:4];
    endcase
  end

  // REG#108の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0108 <= imem03_in[3:0];
    endcase
  end

  // REG#109の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0109 <= imem06_in[15:12];
    endcase
  end

  // REG#110の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0110 <= imem06_in[11:8];
    endcase
  end

  // REG#111の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0111 <= imem02_in[3:0];
    endcase
  end

  // REG#112の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0112 <= imem02_in[7:4];
    endcase
  end

  // REG#113の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0113 <= imem03_in[11:8];
    endcase
  end

  // REG#114の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0114 <= imem07_in[15:12];
    endcase
  end

  // REG#115の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0115 <= imem06_in[3:0];
    endcase
  end

  // REG#116の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0116 <= imem06_in[7:4];
    endcase
  end

  // REG#117の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0117 <= imem04_in[3:0];
    13: reg_0117 <= imem04_in[3:0];
    76: reg_0117 <= imem04_in[3:0];
    endcase
  end

  // REG#118の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0118 <= imem05_in[11:8];
    14: reg_0118 <= imem05_in[11:8];
    endcase
  end

  // REG#119の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0119 <= imem06_in[7:4];
    14: reg_0119 <= imem06_in[7:4];
    17: reg_0119 <= imem06_in[7:4];
    endcase
  end

  // REG#120の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0120 <= imem01_in[15:12];
    17: reg_0120 <= imem01_in[15:12];
    44: reg_0120 <= imem06_in[11:8];
    46: reg_0120 <= imem06_in[11:8];
    69: reg_0120 <= imem06_in[11:8];
    84: reg_0120 <= imem01_in[15:12];
    96: reg_0120 <= imem06_in[11:8];
    101: reg_0120 <= imem01_in[15:12];
    110: reg_0120 <= imem01_in[15:12];
    113: reg_0120 <= imem06_in[11:8];
    115: reg_0120 <= imem06_in[11:8];
    117: reg_0120 <= imem06_in[11:8];
    119: reg_0120 <= imem01_in[15:12];
    127: reg_0120 <= imem01_in[15:12];
    130: reg_0120 <= imem06_in[11:8];
    endcase
  end

  // REG#121の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0121 <= imem03_in[11:8];
    21: reg_0121 <= imem00_in[7:4];
    35: reg_0121 <= imem03_in[11:8];
    72: reg_0121 <= imem00_in[7:4];
    79: reg_0121 <= imem00_in[7:4];
    84: reg_0121 <= imem03_in[11:8];
    101: reg_0121 <= imem00_in[7:4];
    106: reg_0121 <= imem03_in[11:8];
    107: reg_0121 <= op2_01_out;
    130: reg_0121 <= imem00_in[7:4];
    131: reg_0121 <= op2_01_out;
    endcase
  end

  // REG#122の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0122 <= imem00_in[3:0];
    22: reg_0122 <= imem00_in[3:0];
    endcase
  end

  // REG#123の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0123 <= imem07_in[11:8];
    28: reg_0123 <= imem07_in[11:8];
    endcase
  end

  // REG#124の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0124 <= imem07_in[15:12];
    28: reg_0124 <= imem07_in[15:12];
    121: reg_0124 <= imem07_in[15:12];
    125: reg_0124 <= imem07_in[15:12];
    129: reg_0124 <= imem07_in[15:12];
    endcase
  end

  // REG#125の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0125 <= imem02_in[11:8];
    128: reg_0125 <= imem02_in[11:8];
    130: reg_0125 <= imem02_in[11:8];
    endcase
  end

  // REG#126の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0126 <= imem02_in[15:12];
    endcase
  end

  // REG#127の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0127 <= imem02_in[7:4];
    endcase
  end

  // REG#128の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0128 <= imem02_in[3:0];
    endcase
  end

  // REG#129の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0129 <= imem04_in[7:4];
    13: reg_0129 <= imem04_in[7:4];
    74: reg_0129 <= op1_04_out;
    76: reg_0129 <= op1_04_out;
    78: reg_0129 <= op1_04_out;
    90: reg_0129 <= op1_04_out;
    93: reg_0129 <= imem04_in[7:4];
    94: reg_0129 <= op1_04_out;
    97: reg_0129 <= imem04_in[7:4];
    99: reg_0129 <= imem04_in[7:4];
    102: reg_0129 <= imem04_in[7:4];
    104: reg_0129 <= imem04_in[7:4];
    106: reg_0129 <= imem04_in[7:4];
    109: reg_0129 <= imem04_in[7:4];
    110: reg_0129 <= op1_04_out;
    113: reg_0129 <= imem04_in[7:4];
    128: reg_0129 <= imem04_in[7:4];
    endcase
  end

  // REG#130の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0130 <= imem05_in[3:0];
    14: reg_0130 <= imem05_in[3:0];
    endcase
  end

  // REG#131の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0131 <= imem05_in[15:12];
    13: reg_0131 <= imem05_in[15:12];
    56: reg_0131 <= imem05_in[15:12];
    80: reg_0131 <= imem05_in[15:12];
    endcase
  end

  // REG#132の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0132 <= imem06_in[11:8];
    14: reg_0132 <= imem06_in[11:8];
    29: reg_0132 <= imem06_in[11:8];
    endcase
  end

  // REG#133の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0133 <= imem02_in[15:12];
    18: reg_0133 <= imem02_in[15:12];
    21: reg_0133 <= imem02_in[15:12];
    37: reg_0133 <= imem02_in[15:12];
    44: reg_0133 <= imem06_in[3:0];
    47: reg_0133 <= imem06_in[3:0];
    51: reg_0133 <= imem02_in[15:12];
    61: reg_0133 <= imem06_in[3:0];
    75: reg_0133 <= imem06_in[3:0];
    94: reg_0133 <= imem02_in[15:12];
    97: reg_0133 <= imem02_in[15:12];
    100: reg_0133 <= imem06_in[3:0];
    102: reg_0133 <= imem02_in[15:12];
    120: reg_0133 <= imem06_in[3:0];
    endcase
  end

  // REG#134の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0134 <= imem00_in[3:0];
    21: reg_0134 <= op2_00_out;
    24: reg_0134 <= imem00_in[3:0];
    endcase
  end

  // REG#135の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0135 <= imem00_in[7:4];
    22: reg_0135 <= imem07_in[11:8];
    27: reg_0135 <= imem00_in[7:4];
    44: reg_0135 <= imem07_in[11:8];
    53: reg_0135 <= imem00_in[7:4];
    65: reg_0135 <= imem07_in[11:8];
    124: reg_0135 <= imem00_in[7:4];
    126: reg_0135 <= imem07_in[11:8];
    131: reg_0135 <= imem00_in[7:4];
    endcase
  end

  // REG#136の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0136 <= imem00_in[15:12];
    22: reg_0136 <= imem05_in[3:0];
    28: reg_0136 <= imem00_in[15:12];
    68: reg_0136 <= imem05_in[3:0];
    83: reg_0136 <= imem00_in[15:12];
    85: reg_0136 <= imem00_in[15:12];
    87: reg_0136 <= imem05_in[3:0];
    131: reg_0136 <= imem05_in[3:0];
    endcase
  end

  // REG#137の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0137 <= imem07_in[11:8];
    32: reg_0137 <= imem07_in[11:8];
    endcase
  end

  // REG#138の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0138 <= imem02_in[3:0];
    37: reg_0138 <= imem02_in[3:0];
    44: reg_0138 <= imem02_in[3:0];
    72: reg_0138 <= imem02_in[3:0];
    endcase
  end

  // REG#139の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0139 <= imem07_in[7:4];
    39: reg_0139 <= imem07_in[7:4];
    59: reg_0139 <= imem07_in[7:4];
    endcase
  end

  // REG#140の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0140 <= imem07_in[15:12];
    39: reg_0140 <= imem07_in[15:12];
    60: reg_0140 <= imem07_in[15:12];
    endcase
  end

  // REG#141の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0141 <= imem06_in[15:12];
    42: reg_0141 <= imem06_in[15:12];
    59: reg_0141 <= imem06_in[15:12];
    endcase
  end

  // REG#142の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0142 <= imem03_in[15:12];
    57: reg_0142 <= imem03_in[15:12];
    76: reg_0142 <= imem03_in[15:12];
    endcase
  end

  // REG#143の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0143 <= imem03_in[7:4];
    62: reg_0143 <= imem03_in[7:4];
    endcase
  end

  // REG#144の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0144 <= imem03_in[11:8];
    62: reg_0144 <= imem03_in[11:8];
    endcase
  end

  // REG#145の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0145 <= imem03_in[3:0];
    62: reg_0145 <= imem03_in[3:0];
    endcase
  end

  // REG#146の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0146 <= imem01_in[15:12];
    endcase
  end

  // REG#147の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0147 <= imem01_in[3:0];
    endcase
  end

  // REG#148の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0148 <= imem01_in[11:8];
    endcase
  end

  // REG#149の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0149 <= imem01_in[7:4];
    endcase
  end

  // REG#150の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0150 <= imem04_in[15:12];
    13: reg_0150 <= imem04_in[15:12];
    71: reg_0150 <= op1_10_out;
    73: reg_0150 <= op1_10_out;
    75: reg_0150 <= op1_10_out;
    89: reg_0150 <= op1_10_out;
    91: reg_0150 <= op1_10_out;
    93: reg_0150 <= op1_10_out;
    96: reg_0150 <= imem04_in[15:12];
    97: reg_0150 <= op1_10_out;
    99: reg_0150 <= op1_10_out;
    102: reg_0150 <= imem04_in[15:12];
    103: reg_0150 <= op1_10_out;
    106: reg_0150 <= imem04_in[15:12];
    107: reg_0150 <= op1_10_out;
    109: reg_0150 <= op1_10_out;
    111: reg_0150 <= op1_10_out;
    113: reg_0150 <= op1_10_out;
    115: reg_0150 <= op1_10_out;
    117: reg_0150 <= op1_10_out;
    119: reg_0150 <= op1_10_out;
    121: reg_0150 <= op1_10_out;
    123: reg_0150 <= op1_10_out;
    125: reg_0150 <= op1_10_out;
    127: reg_0150 <= op1_10_out;
    129: reg_0150 <= op1_10_out;
    131: reg_0150 <= op1_10_out;
    endcase
  end

  // REG#151の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0151 <= imem05_in[11:8];
    15: reg_0151 <= imem05_in[11:8];
    41: reg_0151 <= imem05_in[11:8];
    endcase
  end

  // REG#152の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0152 <= imem06_in[15:12];
    13: reg_0152 <= imem06_in[15:12];
    endcase
  end

  // REG#153の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0153 <= imem02_in[7:4];
    17: reg_0153 <= imem00_in[3:0];
    22: reg_0153 <= imem02_in[7:4];
    85: reg_0153 <= imem00_in[3:0];
    87: reg_0153 <= imem00_in[3:0];
    endcase
  end

  // REG#154の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0154 <= imem03_in[7:4];
    21: reg_0154 <= imem02_in[7:4];
    37: reg_0154 <= imem02_in[7:4];
    40: reg_0154 <= imem02_in[7:4];
    66: reg_0154 <= imem03_in[7:4];
    71: reg_0154 <= imem03_in[7:4];
    83: reg_0154 <= imem03_in[7:4];
    130: reg_0154 <= imem02_in[7:4];
    endcase
  end

  // REG#155の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0155 <= imem00_in[7:4];
    22: reg_0155 <= imem06_in[3:0];
    28: reg_0155 <= imem00_in[7:4];
    68: reg_0155 <= imem00_in[7:4];
    130: reg_0155 <= imem06_in[3:0];
    endcase
  end

  // REG#156の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0156 <= imem07_in[7:4];
    40: reg_0156 <= imem07_in[7:4];
    129: reg_0156 <= imem07_in[7:4];
    endcase
  end

  // REG#157の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0157 <= imem07_in[15:12];
    40: reg_0157 <= imem07_in[15:12];
    endcase
  end

  // REG#158の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0158 <= imem07_in[11:8];
    40: reg_0158 <= imem07_in[11:8];
    endcase
  end

  // REG#159の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0159 <= imem07_in[3:0];
    40: reg_0159 <= imem07_in[3:0];
    endcase
  end

  // REG#160の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0160 <= imem01_in[3:0];
    44: reg_0160 <= imem06_in[15:12];
    48: reg_0160 <= imem06_in[15:12];
    51: reg_0160 <= imem01_in[3:0];
    58: reg_0160 <= imem01_in[3:0];
    63: reg_0160 <= imem06_in[15:12];
    84: reg_0160 <= imem06_in[15:12];
    85: reg_0160 <= op2_01_out;
    91: reg_0160 <= op2_01_out;
    103: reg_0160 <= op2_01_out;
    115: reg_0160 <= op2_01_out;
    endcase
  end

  // REG#161の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0161 <= imem01_in[11:8];
    44: reg_0161 <= imem06_in[7:4];
    48: reg_0161 <= imem06_in[7:4];
    51: reg_0161 <= imem01_in[11:8];
    54: reg_0161 <= imem01_in[11:8];
    73: reg_0161 <= imem06_in[7:4];
    81: reg_0161 <= imem01_in[11:8];
    87: reg_0161 <= imem06_in[7:4];
    128: reg_0161 <= imem06_in[7:4];
    130: reg_0161 <= imem01_in[11:8];
    endcase
  end

  // REG#162の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0162 <= imem01_in[15:12];
    44: reg_0162 <= imem07_in[15:12];
    53: reg_0162 <= imem07_in[15:12];
    67: reg_0162 <= imem07_in[15:12];
    69: reg_0162 <= imem07_in[15:12];
    76: reg_0162 <= imem07_in[15:12];
    82: reg_0162 <= imem07_in[15:12];
    85: reg_0162 <= imem01_in[15:12];
    endcase
  end

  // REG#163の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0163 <= imem01_in[7:4];
    44: reg_0163 <= imem05_in[7:4];
    74: reg_0163 <= imem01_in[7:4];
    endcase
  end

  // REG#164の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0164 <= imem04_in[3:0];
    14: reg_0164 <= imem04_in[3:0];
    69: reg_0164 <= op1_04_out;
    71: reg_0164 <= op1_04_out;
    75: reg_0164 <= op1_04_out;
    77: reg_0164 <= op1_04_out;
    89: reg_0164 <= op1_04_out;
    92: reg_0164 <= imem04_in[3:0];
    112: reg_0164 <= imem04_in[3:0];
    114: reg_0164 <= imem04_in[3:0];
    122: reg_0164 <= imem04_in[3:0];
    125: reg_0164 <= imem04_in[3:0];
    endcase
  end

  // REG#165の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0165 <= imem06_in[15:12];
    13: reg_0165 <= imem01_in[15:12];
    17: reg_0165 <= imem06_in[15:12];
    endcase
  end

  // REG#166の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0166 <= imem01_in[3:0];
    17: reg_0166 <= imem01_in[3:0];
    56: reg_0166 <= imem01_in[3:0];
    58: reg_0166 <= imem01_in[15:12];
    64: reg_0166 <= imem01_in[15:12];
    75: reg_0166 <= imem01_in[3:0];
    94: reg_0166 <= imem01_in[3:0];
    98: reg_0166 <= imem01_in[3:0];
    100: reg_0166 <= imem01_in[3:0];
    104: reg_0166 <= imem01_in[15:12];
    112: reg_0166 <= imem01_in[3:0];
    114: reg_0166 <= imem01_in[15:12];
    endcase
  end

  // REG#167の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0167 <= imem01_in[11:8];
    17: reg_0167 <= imem01_in[11:8];
    44: reg_0167 <= imem05_in[3:0];
    76: reg_0167 <= imem01_in[11:8];
    78: reg_0167 <= imem05_in[3:0];
    80: reg_0167 <= imem05_in[3:0];
    endcase
  end

  // REG#168の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0168 <= imem02_in[7:4];
    17: reg_0168 <= imem05_in[7:4];
    58: reg_0168 <= imem05_in[7:4];
    82: reg_0168 <= imem02_in[7:4];
    endcase
  end

  // REG#169の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0169 <= imem02_in[15:12];
    19: reg_0169 <= imem02_in[15:12];
    21: reg_0169 <= imem07_in[3:0];
    39: reg_0169 <= imem07_in[3:0];
    60: reg_0169 <= imem02_in[15:12];
    79: reg_0169 <= imem02_in[15:12];
    111: reg_0169 <= imem02_in[15:12];
    117: reg_0169 <= imem02_in[15:12];
    120: reg_0169 <= imem07_in[3:0];
    129: reg_0169 <= imem02_in[15:12];
    endcase
  end

  // REG#170の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0170 <= imem07_in[3:0];
    19: reg_0170 <= imem07_in[3:0];
    41: reg_0170 <= imem07_in[3:0];
    86: reg_0170 <= imem07_in[3:0];
    endcase
  end

  // REG#171の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0171 <= imem00_in[7:4];
    22: reg_0171 <= imem06_in[7:4];
    28: reg_0171 <= imem06_in[7:4];
    129: reg_0171 <= imem00_in[7:4];
    endcase
  end

  // REG#172の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0172 <= imem00_in[11:8];
    22: reg_0172 <= imem06_in[15:12];
    28: reg_0172 <= imem00_in[11:8];
    64: reg_0172 <= imem06_in[15:12];
    74: reg_0172 <= imem06_in[15:12];
    127: reg_0172 <= imem06_in[15:12];
    endcase
  end

  // REG#173の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0173 <= imem05_in[3:0];
    48: reg_0173 <= imem05_in[3:0];
    82: reg_0173 <= imem05_in[3:0];
    endcase
  end

  // REG#174の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0174 <= imem05_in[15:12];
    48: reg_0174 <= imem05_in[15:12];
    84: reg_0174 <= imem05_in[15:12];
    123: reg_0174 <= imem05_in[15:12];
    endcase
  end

  // REG#175の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0175 <= imem05_in[7:4];
    50: reg_0175 <= imem05_in[7:4];
    58: reg_0175 <= imem01_in[7:4];
    65: reg_0175 <= imem01_in[7:4];
    79: reg_0175 <= imem05_in[7:4];
    88: reg_0175 <= imem01_in[7:4];
    endcase
  end

  // REG#176の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0176 <= imem05_in[11:8];
    50: reg_0176 <= imem05_in[11:8];
    57: reg_0176 <= imem05_in[11:8];
    endcase
  end

  // REG#177の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0177 <= imem03_in[15:12];
    53: reg_0177 <= imem03_in[15:12];
    65: reg_0177 <= imem03_in[15:12];
    81: reg_0177 <= imem03_in[15:12];
    endcase
  end

  // REG#178の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0178 <= imem03_in[11:8];
    55: reg_0178 <= imem03_in[11:8];
    endcase
  end

  // REG#179の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0179 <= imem03_in[3:0];
    57: reg_0179 <= op1_02_out;
    73: reg_0179 <= op1_02_out;
    75: reg_0179 <= op1_02_out;
    77: reg_0179 <= op1_02_out;
    79: reg_0179 <= op1_02_out;
    82: reg_0179 <= imem03_in[3:0];
    endcase
  end

  // REG#180の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0180 <= imem03_in[7:4];
    58: reg_0180 <= imem03_in[7:4];
    endcase
  end

  // REG#181の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0181 <= imem04_in[15:12];
    14: reg_0181 <= imem04_in[15:12];
    65: reg_0181 <= imem04_in[15:12];
    113: reg_0181 <= imem04_in[15:12];
    126: reg_0181 <= imem04_in[15:12];
    129: reg_0181 <= imem04_in[15:12];
    endcase
  end

  // REG#182の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0182 <= imem05_in[7:4];
    13: reg_0182 <= imem05_in[7:4];
    55: reg_0182 <= imem05_in[7:4];
    78: reg_0182 <= imem05_in[7:4];
    81: reg_0182 <= imem05_in[7:4];
    endcase
  end

  // REG#183の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0183 <= imem01_in[3:0];
    18: reg_0183 <= imem01_in[3:0];
    22: reg_0183 <= imem01_in[3:0];
    44: reg_0183 <= imem05_in[15:12];
    76: reg_0183 <= imem05_in[15:12];
    101: reg_0183 <= imem01_in[3:0];
    110: reg_0183 <= imem05_in[15:12];
    116: reg_0183 <= imem01_in[3:0];
    118: reg_0183 <= imem01_in[3:0];
    130: reg_0183 <= imem05_in[15:12];
    endcase
  end

  // REG#184の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0184 <= imem02_in[7:4];
    17: reg_0184 <= imem05_in[15:12];
    61: reg_0184 <= imem02_in[7:4];
    86: reg_0184 <= imem05_in[15:12];
    118: reg_0184 <= imem02_in[7:4];
    129: reg_0184 <= imem05_in[15:12];
    endcase
  end

  // REG#185の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0185 <= imem03_in[3:0];
    21: reg_0185 <= imem07_in[15:12];
    39: reg_0185 <= imem03_in[3:0];
    58: reg_0185 <= imem07_in[15:12];
    69: reg_0185 <= imem03_in[3:0];
    78: reg_0185 <= imem07_in[15:12];
    81: reg_0185 <= imem07_in[15:12];
    83: reg_0185 <= imem03_in[3:0];
    endcase
  end

  // REG#186の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0186 <= imem00_in[7:4];
    22: reg_0186 <= imem07_in[15:12];
    31: reg_0186 <= imem00_in[7:4];
    35: reg_0186 <= imem07_in[15:12];
    62: reg_0186 <= imem07_in[15:12];
    86: reg_0186 <= imem00_in[7:4];
    130: reg_0186 <= imem07_in[15:12];
    endcase
  end

  // REG#187の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0187 <= imem07_in[15:12];
    42: reg_0187 <= imem07_in[15:12];
    59: reg_0187 <= op2_00_out;
    61: reg_0187 <= op2_00_out;
    64: reg_0187 <= imem07_in[15:12];
    84: reg_0187 <= op2_00_out;
    86: reg_0187 <= op2_00_out;
    102: reg_0187 <= op2_00_out;
    110: reg_0187 <= op2_00_out;
    endcase
  end

  // REG#188の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0188 <= imem00_in[3:0];
    44: reg_0188 <= imem00_in[3:0];
    endcase
  end

  // REG#189の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0189 <= imem00_in[15:12];
    44: reg_0189 <= imem00_in[15:12];
    endcase
  end

  // REG#190の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0190 <= imem07_in[11:8];
    44: reg_0190 <= imem03_in[3:0];
    112: reg_0190 <= imem07_in[11:8];
    115: reg_0190 <= imem03_in[3:0];
    118: reg_0190 <= imem03_in[3:0];
    endcase
  end

  // REG#191の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0191 <= imem07_in[7:4];
    44: reg_0191 <= imem07_in[7:4];
    53: reg_0191 <= imem07_in[7:4];
    67: reg_0191 <= imem03_in[15:12];
    72: reg_0191 <= imem07_in[7:4];
    74: reg_0191 <= imem03_in[15:12];
    89: reg_0191 <= imem03_in[15:12];
    131: reg_0191 <= imem07_in[7:4];
    endcase
  end

  // REG#192の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0192 <= imem06_in[15:12];
    50: reg_0192 <= imem06_in[15:12];
    69: reg_0192 <= imem06_in[15:12];
    87: reg_0192 <= imem06_in[15:12];
    128: reg_0192 <= imem06_in[15:12];
    endcase
  end

  // REG#193の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0193 <= imem06_in[11:8];
    51: reg_0193 <= imem06_in[11:8];
    64: reg_0193 <= op1_12_out;
    67: reg_0193 <= imem06_in[11:8];
    76: reg_0193 <= op1_12_out;
    79: reg_0193 <= imem06_in[11:8];
    81: reg_0193 <= op1_12_out;
    83: reg_0193 <= op1_12_out;
    85: reg_0193 <= op1_12_out;
    87: reg_0193 <= op1_12_out;
    90: reg_0193 <= imem06_in[11:8];
    100: reg_0193 <= imem06_in[11:8];
    102: reg_0193 <= imem06_in[11:8];
    103: reg_0193 <= op1_12_out;
    106: reg_0193 <= op1_12_out;
    109: reg_0193 <= imem06_in[11:8];
    111: reg_0193 <= imem06_in[11:8];
    113: reg_0193 <= op1_12_out;
    115: reg_0193 <= op1_12_out;
    118: reg_0193 <= imem06_in[11:8];
    119: reg_0193 <= op1_12_out;
    121: reg_0193 <= op1_12_out;
    123: reg_0193 <= op1_12_out;
    125: reg_0193 <= op1_12_out;
    127: reg_0193 <= op1_12_out;
    129: reg_0193 <= op1_12_out;
    endcase
  end

  // REG#194の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0194 <= imem06_in[3:0];
    52: reg_0194 <= imem06_in[3:0];
    59: reg_0194 <= imem06_in[3:0];
    131: reg_0194 <= imem06_in[3:0];
    endcase
  end

  // REG#195の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0195 <= imem06_in[7:4];
    52: reg_0195 <= imem06_in[7:4];
    66: reg_0195 <= imem06_in[7:4];
    82: reg_0195 <= imem06_in[7:4];
    98: reg_0195 <= imem06_in[7:4];
    endcase
  end

  // REG#196の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0196 <= imem01_in[15:12];
    17: reg_0196 <= imem05_in[11:8];
    64: reg_0196 <= imem05_in[11:8];
    endcase
  end

  // REG#197の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0197 <= imem02_in[15:12];
    17: reg_0197 <= imem05_in[3:0];
    65: reg_0197 <= imem05_in[3:0];
    129: reg_0197 <= imem05_in[3:0];
    endcase
  end

  // REG#198の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0198 <= imem07_in[3:0];
    17: reg_0198 <= imem03_in[15:12];
    77: reg_0198 <= imem07_in[3:0];
    80: reg_0198 <= imem03_in[15:12];
    endcase
  end

  // REG#199の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0199 <= imem03_in[15:12];
    21: reg_0199 <= imem04_in[15:12];
    42: reg_0199 <= imem04_in[15:12];
    69: reg_0199 <= imem03_in[15:12];
    81: reg_0199 <= imem04_in[15:12];
    endcase
  end

  // REG#200の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0200 <= op1_00_out;
    22: reg_0200 <= op1_00_out;
    88: reg_0200 <= op1_00_out;
    90: reg_0200 <= op2_07_out;
    92: reg_0200 <= op2_00_out;
    114: reg_0200 <= op2_00_out;
    endcase
  end

  // REG#201の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0201 <= imem00_in[11:8];
    44: reg_0201 <= imem00_in[11:8];
    endcase
  end

  // REG#202の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0202 <= imem00_in[3:0];
    54: reg_0202 <= imem00_in[3:0];
    65: reg_0202 <= imem00_in[3:0];
    endcase
  end

  // REG#203の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0203 <= imem00_in[7:4];
    54: reg_0203 <= imem00_in[7:4];
    64: reg_0203 <= imem00_in[7:4];
    endcase
  end

  // REG#204の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0204 <= imem05_in[7:4];
    60: reg_0204 <= imem05_in[7:4];
    96: reg_0204 <= imem05_in[7:4];
    117: reg_0204 <= op2_02_out;
    123: reg_0204 <= op2_02_out;
    endcase
  end

  // REG#205の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0205 <= imem05_in[3:0];
    61: reg_0205 <= imem05_in[3:0];
    92: reg_0205 <= imem05_in[3:0];
    endcase
  end

  // REG#206の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0206 <= imem05_in[15:12];
    62: reg_0206 <= imem05_in[15:12];
    endcase
  end

  // REG#207の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0207 <= imem05_in[11:8];
    62: reg_0207 <= imem05_in[11:8];
    128: reg_0207 <= imem05_in[11:8];
    endcase
  end

  // REG#208の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0208 <= imem04_in[15:12];
    66: reg_0208 <= imem04_in[15:12];
    91: reg_0208 <= imem04_in[15:12];
    94: reg_0208 <= imem04_in[15:12];
    119: reg_0208 <= imem04_in[15:12];
    125: reg_0208 <= op2_02_out;
    endcase
  end

  // REG#209の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0209 <= imem04_in[11:8];
    71: reg_0209 <= op1_11_out;
    73: reg_0209 <= op1_11_out;
    76: reg_0209 <= imem04_in[11:8];
    131: reg_0209 <= op1_11_out;
    endcase
  end

  // REG#210の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0210 <= imem04_in[7:4];
    73: reg_0210 <= imem04_in[7:4];
    endcase
  end

  // REG#211の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0211 <= imem04_in[3:0];
    74: reg_0211 <= op1_14_out;
    77: reg_0211 <= imem04_in[3:0];
    122: reg_0211 <= op1_14_out;
    125: reg_0211 <= op1_14_out;
    127: reg_0211 <= op1_14_out;
    130: reg_0211 <= imem04_in[3:0];
    endcase
  end

  // REG#212の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0212 <= imem06_in[3:0];
    126: reg_0212 <= imem06_in[3:0];
    endcase
  end

  // REG#213の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0213 <= imem06_in[15:12];
    endcase
  end

  // REG#214の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0214 <= imem06_in[11:8];
    endcase
  end

  // REG#215の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0215 <= imem06_in[7:4];
    endcase
  end

  // REG#216の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0216 <= imem02_in[7:4];
    17: reg_0216 <= imem03_in[3:0];
    80: reg_0216 <= imem03_in[3:0];
    endcase
  end

  // REG#217の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0217 <= imem02_in[11:8];
    17: reg_0217 <= imem02_in[11:8];
    endcase
  end

  // REG#218の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0218 <= imem03_in[7:4];
    21: reg_0218 <= imem00_in[15:12];
    43: reg_0218 <= imem03_in[7:4];
    54: reg_0218 <= imem03_in[7:4];
    67: reg_0218 <= imem03_in[7:4];
    71: reg_0218 <= imem00_in[15:12];
    86: reg_0218 <= imem03_in[7:4];
    endcase
  end

  // REG#219の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0219 <= imem00_in[7:4];
    22: reg_0219 <= imem07_in[7:4];
    32: reg_0219 <= imem00_in[7:4];
    52: reg_0219 <= imem00_in[7:4];
    81: reg_0219 <= imem00_in[7:4];
    87: reg_0219 <= imem07_in[7:4];
    endcase
  end

  // REG#220の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0220 <= imem00_in[11:8];
    36: reg_0220 <= imem00_in[11:8];
    44: reg_0220 <= imem03_in[11:8];
    112: reg_0220 <= imem03_in[11:8];
    endcase
  end

  // REG#221の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0221 <= imem00_in[15:12];
    35: reg_0221 <= imem05_in[11:8];
    48: reg_0221 <= imem00_in[15:12];
    endcase
  end

  // REG#222の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0222 <= imem01_in[3:0];
    35: reg_0222 <= imem01_in[3:0];
    73: reg_0222 <= imem01_in[3:0];
    endcase
  end

  // REG#223の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0223 <= imem07_in[3:0];
    59: reg_0223 <= imem07_in[3:0];
    endcase
  end

  // REG#224の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0224 <= imem07_in[11:8];
    59: reg_0224 <= imem07_in[11:8];
    endcase
  end

  // REG#225の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0225 <= imem07_in[7:4];
    60: reg_0225 <= imem07_in[7:4];
    endcase
  end

  // REG#226の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0226 <= imem07_in[15:12];
    61: reg_0226 <= op1_01_out;
    71: reg_0226 <= imem07_in[15:12];
    75: reg_0226 <= imem07_in[15:12];
    76: reg_0226 <= op1_01_out;
    78: reg_0226 <= op1_01_out;
    80: reg_0226 <= op1_01_out;
    90: reg_0226 <= op1_01_out;
    92: reg_0226 <= op1_01_out;
    94: reg_0226 <= op1_01_out;
    97: reg_0226 <= imem07_in[15:12];
    99: reg_0226 <= imem07_in[15:12];
    102: reg_0226 <= op1_01_out;
    105: reg_0226 <= imem07_in[15:12];
    114: reg_0226 <= op1_01_out;
    116: reg_0226 <= op1_01_out;
    119: reg_0226 <= imem07_in[15:12];
    endcase
  end

  // REG#227の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0227 <= imem02_in[11:8];
    17: reg_0227 <= imem03_in[7:4];
    83: reg_0227 <= imem02_in[11:8];
    endcase
  end

  // REG#228の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0228 <= imem07_in[15:12];
    17: reg_0228 <= imem07_in[15:12];
    23: reg_0228 <= imem07_in[15:12];
    endcase
  end

  // REG#229の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0229 <= imem00_in[15:12];
    22: reg_0229 <= imem07_in[3:0];
    31: reg_0229 <= imem00_in[15:12];
    52: reg_0229 <= imem07_in[3:0];
    69: reg_0229 <= imem00_in[15:12];
    130: reg_0229 <= imem00_in[15:12];
    endcase
  end

  // REG#230の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0230 <= imem07_in[3:0];
    44: reg_0230 <= imem07_in[3:0];
    53: reg_0230 <= imem07_in[3:0];
    66: reg_0230 <= imem07_in[3:0];
    68: reg_0230 <= op1_00_out;
    70: reg_0230 <= op1_00_out;
    78: reg_0230 <= op1_00_out;
    89: reg_0230 <= op1_00_out;
    92: reg_0230 <= imem07_in[3:0];
    94: reg_0230 <= imem07_in[3:0];
    96: reg_0230 <= op2_00_out;
    endcase
  end

  // REG#231の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0231 <= imem07_in[7:4];
    43: reg_0231 <= op1_01_out;
    120: reg_0231 <= op1_01_out;
    122: reg_0231 <= op1_01_out;
    125: reg_0231 <= imem07_in[7:4];
    endcase
  end

  // REG#232の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0232 <= imem03_in[7:4];
    48: reg_0232 <= imem03_in[7:4];
    60: reg_0232 <= imem04_in[11:8];
    65: reg_0232 <= imem03_in[7:4];
    79: reg_0232 <= imem04_in[11:8];
    127: reg_0232 <= imem03_in[7:4];
    endcase
  end

  // REG#233の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0233 <= imem03_in[11:8];
    48: reg_0233 <= imem03_in[11:8];
    62: reg_0233 <= imem02_in[11:8];
    72: reg_0233 <= imem03_in[11:8];
    118: reg_0233 <= imem03_in[11:8];
    125: reg_0233 <= imem03_in[11:8];
    131: reg_0233 <= imem03_in[11:8];
    endcase
  end

  // REG#234の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0234 <= imem03_in[15:12];
    48: reg_0234 <= imem03_in[15:12];
    62: reg_0234 <= imem03_in[15:12];
    endcase
  end

  // REG#235の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0235 <= imem03_in[3:0];
    50: reg_0235 <= imem03_in[3:0];
    71: reg_0235 <= imem03_in[3:0];
    84: reg_0235 <= imem03_in[3:0];
    101: reg_0235 <= imem03_in[3:0];
    107: reg_0235 <= imem03_in[3:0];
    113: reg_0235 <= imem03_in[3:0];
    115: reg_0235 <= imem03_in[11:8];
    118: reg_0235 <= imem07_in[15:12];
    endcase
  end

  // REG#236の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0236 <= imem04_in[7:4];
    77: reg_0236 <= imem04_in[7:4];
    125: reg_0236 <= imem04_in[7:4];
    endcase
  end

  // REG#237の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0237 <= imem04_in[11:8];
    77: reg_0237 <= op2_00_out;
    79: reg_0237 <= op2_00_out;
    87: reg_0237 <= imem04_in[11:8];
    88: reg_0237 <= op2_00_out;
    91: reg_0237 <= imem04_in[11:8];
    95: reg_0237 <= op2_00_out;
    130: reg_0237 <= op2_00_out;
    endcase
  end

  // REG#238の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0238 <= imem01_in[11:8];
    125: reg_0238 <= imem01_in[11:8];
    endcase
  end

  // REG#239の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0239 <= imem01_in[7:4];
    130: reg_0239 <= imem01_in[7:4];
    endcase
  end

  // REG#240の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0240 <= imem05_in[15:12];
    endcase
  end

  // REG#241の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0241 <= imem01_in[15:12];
    endcase
  end

  // REG#242の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0242 <= imem01_in[3:0];
    130: reg_0242 <= imem01_in[3:0];
    endcase
  end

  // REG#243の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0243 <= imem05_in[7:4];
    endcase
  end

  // REG#244の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0244 <= imem06_in[11:8];
    17: reg_0244 <= imem06_in[11:8];
    endcase
  end

  // REG#245の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0245 <= imem07_in[7:4];
    17: reg_0245 <= imem07_in[7:4];
    36: reg_0245 <= imem07_in[7:4];
    64: reg_0245 <= imem07_in[7:4];
    86: reg_0245 <= op2_02_out;
    107: reg_0245 <= op2_02_out;
    130: reg_0245 <= op2_02_out;
    endcase
  end

  // REG#246の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0246 <= imem03_in[15:12];
    21: reg_0246 <= imem07_in[7:4];
    44: reg_0246 <= imem03_in[15:12];
    109: reg_0246 <= imem03_in[15:12];
    117: reg_0246 <= imem07_in[7:4];
    120: reg_0246 <= imem07_in[7:4];
    127: reg_0246 <= imem03_in[15:12];
    endcase
  end

  // REG#247の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0247 <= imem04_in[7:4];
    21: reg_0247 <= imem06_in[15:12];
    54: reg_0247 <= imem04_in[7:4];
    67: reg_0247 <= imem04_in[7:4];
    88: reg_0247 <= imem04_in[7:4];
    90: reg_0247 <= imem04_in[7:4];
    93: reg_0247 <= imem06_in[15:12];
    95: reg_0247 <= op2_01_out;
    endcase
  end

  // REG#248の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0248 <= imem00_in[3:0];
    21: reg_0248 <= op1_00_out;
    38: reg_0248 <= imem00_in[3:0];
    43: reg_0248 <= op1_00_out;
    81: reg_0248 <= op1_00_out;
    92: reg_0248 <= imem06_in[11:8];
    94: reg_0248 <= imem00_in[3:0];
    96: reg_0248 <= imem00_in[3:0];
    98: reg_0248 <= imem00_in[3:0];
    104: reg_0248 <= imem00_in[3:0];
    113: reg_0248 <= imem00_in[3:0];
    115: reg_0248 <= imem00_in[3:0];
    124: reg_0248 <= imem00_in[3:0];
    126: reg_0248 <= imem00_in[3:0];
    endcase
  end

  // REG#249の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0249 <= imem00_in[7:4];
    36: reg_0249 <= imem00_in[7:4];
    53: reg_0249 <= op2_00_out;
    56: reg_0249 <= imem00_in[7:4];
    131: reg_0249 <= op2_00_out;
    endcase
  end

  // REG#250の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0250 <= imem00_in[15:12];
    35: reg_0250 <= imem05_in[3:0];
    49: reg_0250 <= imem00_in[15:12];
    endcase
  end

  // REG#251の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0251 <= imem05_in[15:12];
    42: reg_0251 <= imem05_in[15:12];
    60: reg_0251 <= imem05_in[15:12];
    92: reg_0251 <= imem05_in[15:12];
    endcase
  end

  // REG#252の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0252 <= imem07_in[3:0];
    46: reg_0252 <= imem07_in[3:0];
    52: reg_0252 <= imem04_in[11:8];
    58: reg_0252 <= imem04_in[11:8];
    63: reg_0252 <= imem04_in[11:8];
    93: reg_0252 <= imem04_in[11:8];
    98: reg_0252 <= imem04_in[11:8];
    100: reg_0252 <= imem04_in[11:8];
    103: reg_0252 <= imem04_in[11:8];
    105: reg_0252 <= imem04_in[11:8];
    107: reg_0252 <= imem04_in[11:8];
    112: reg_0252 <= imem07_in[3:0];
    115: reg_0252 <= imem04_in[11:8];
    117: reg_0252 <= imem04_in[11:8];
    120: reg_0252 <= imem04_in[11:8];
    endcase
  end

  // REG#253の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0253 <= imem02_in[3:0];
    48: reg_0253 <= imem02_in[3:0];
    100: reg_0253 <= imem02_in[3:0];
    107: reg_0253 <= imem02_in[3:0];
    endcase
  end

  // REG#254の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0254 <= imem02_in[7:4];
    52: reg_0254 <= imem02_in[7:4];
    63: reg_0254 <= imem02_in[7:4];
    102: reg_0254 <= imem02_in[7:4];
    endcase
  end

  // REG#255の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0255 <= imem02_in[15:12];
    52: reg_0255 <= imem02_in[15:12];
    63: reg_0255 <= imem02_in[15:12];
    83: reg_0255 <= imem02_in[15:12];
    endcase
  end

  // REG#256の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0256 <= imem02_in[11:8];
    53: reg_0256 <= imem02_in[11:8];
    58: reg_0256 <= imem02_in[11:8];
    89: reg_0256 <= imem02_in[11:8];
    108: reg_0256 <= imem04_in[11:8];
    endcase
  end

  // REG#257の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0257 <= imem01_in[7:4];
    59: reg_0257 <= imem01_in[7:4];
    67: reg_0257 <= imem01_in[7:4];
    85: reg_0257 <= imem01_in[7:4];
    endcase
  end

  // REG#258の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0258 <= imem01_in[15:12];
    63: reg_0258 <= imem01_in[15:12];
    74: reg_0258 <= imem01_in[15:12];
    endcase
  end

  // REG#259の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0259 <= imem01_in[3:0];
    63: reg_0259 <= imem01_in[3:0];
    72: reg_0259 <= op1_11_out;
    74: reg_0259 <= op1_11_out;
    76: reg_0259 <= op1_11_out;
    78: reg_0259 <= op1_11_out;
    80: reg_0259 <= op1_11_out;
    82: reg_0259 <= op1_11_out;
    91: reg_0259 <= op1_11_out;
    93: reg_0259 <= op1_11_out;
    95: reg_0259 <= op1_11_out;
    97: reg_0259 <= op1_11_out;
    99: reg_0259 <= op1_11_out;
    101: reg_0259 <= op1_11_out;
    103: reg_0259 <= op1_11_out;
    105: reg_0259 <= op1_11_out;
    107: reg_0259 <= op1_11_out;
    109: reg_0259 <= op1_11_out;
    111: reg_0259 <= op1_11_out;
    113: reg_0259 <= op1_11_out;
    115: reg_0259 <= op1_11_out;
    117: reg_0259 <= op1_11_out;
    120: reg_0259 <= op1_11_out;
    122: reg_0259 <= op1_11_out;
    124: reg_0259 <= op1_11_out;
    126: reg_0259 <= op1_11_out;
    129: reg_0259 <= imem01_in[3:0];
    130: reg_0259 <= op1_11_out;
    endcase
  end

  // REG#260の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0260 <= imem01_in[11:8];
    63: reg_0260 <= imem01_in[11:8];
    73: reg_0260 <= imem01_in[11:8];
    endcase
  end

  // REG#261の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0261 <= imem03_in[3:0];
    21: reg_0261 <= imem06_in[3:0];
    57: reg_0261 <= imem03_in[3:0];
    72: reg_0261 <= imem06_in[3:0];
    78: reg_0261 <= imem06_in[3:0];
    81: reg_0261 <= imem03_in[3:0];
    127: reg_0261 <= imem06_in[3:0];
    endcase
  end

  // REG#262の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0262 <= imem04_in[3:0];
    21: reg_0262 <= imem04_in[3:0];
    41: reg_0262 <= imem04_in[3:0];
    endcase
  end

  // REG#263の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0263 <= imem04_in[7:4];
    21: reg_0263 <= imem06_in[7:4];
    59: reg_0263 <= imem04_in[7:4];
    65: reg_0263 <= imem04_in[7:4];
    111: reg_0263 <= imem06_in[7:4];
    114: reg_0263 <= imem04_in[7:4];
    122: reg_0263 <= imem04_in[7:4];
    124: reg_0263 <= imem06_in[7:4];
    126: reg_0263 <= imem06_in[7:4];
    endcase
  end

  // REG#264の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0264 <= imem04_in[11:8];
    21: reg_0264 <= imem06_in[11:8];
    59: reg_0264 <= imem04_in[11:8];
    61: reg_0264 <= imem06_in[11:8];
    75: reg_0264 <= imem06_in[11:8];
    86: reg_0264 <= imem04_in[11:8];
    123: reg_0264 <= imem06_in[11:8];
    129: reg_0264 <= imem04_in[11:8];
    endcase
  end

  // REG#265の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0265 <= op1_00_out;
    23: reg_0265 <= imem06_in[7:4];
    27: reg_0265 <= op1_00_out;
    90: reg_0265 <= op2_08_out;
    94: reg_0265 <= imem06_in[7:4];
    96: reg_0265 <= imem06_in[7:4];
    101: reg_0265 <= imem06_in[7:4];
    endcase
  end

  // REG#266の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0266 <= op1_01_out;
    22: reg_0266 <= op1_01_out;
    90: reg_0266 <= imem05_in[7:4];
    95: reg_0266 <= imem05_in[7:4];
    100: reg_0266 <= op1_01_out;
    103: reg_0266 <= imem05_in[7:4];
    130: reg_0266 <= imem05_in[7:4];
    endcase
  end

  // REG#267の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0267 <= imem00_in[7:4];
    35: reg_0267 <= imem00_in[7:4];
    43: reg_0267 <= imem00_in[7:4];
    endcase
  end

  // REG#268の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0268 <= imem06_in[3:0];
    52: reg_0268 <= imem04_in[15:12];
    60: reg_0268 <= imem04_in[15:12];
    65: reg_0268 <= imem06_in[3:0];
    69: reg_0268 <= imem06_in[3:0];
    87: reg_0268 <= imem04_in[15:12];
    89: reg_0268 <= imem04_in[15:12];
    92: reg_0268 <= imem06_in[3:0];
    95: reg_0268 <= imem04_in[15:12];
    endcase
  end

  // REG#269の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0269 <= imem06_in[11:8];
    54: reg_0269 <= imem06_in[11:8];
    99: reg_0269 <= imem06_in[11:8];
    113: reg_0269 <= imem02_in[7:4];
    115: reg_0269 <= imem01_in[3:0];
    121: reg_0269 <= imem01_in[3:0];
    124: reg_0269 <= imem01_in[3:0];
    endcase
  end

  // REG#270の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0270 <= imem06_in[7:4];
    54: reg_0270 <= imem06_in[7:4];
    99: reg_0270 <= imem06_in[7:4];
    113: reg_0270 <= imem06_in[7:4];
    117: reg_0270 <= imem06_in[7:4];
    119: reg_0270 <= imem06_in[7:4];
    123: reg_0270 <= imem06_in[7:4];
    endcase
  end

  // REG#271の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0271 <= imem06_in[15:12];
    54: reg_0271 <= imem06_in[15:12];
    95: reg_0271 <= imem06_in[15:12];
    endcase
  end

  // REG#272の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0272 <= imem05_in[15:12];
    55: reg_0272 <= imem05_in[15:12];
    79: reg_0272 <= imem05_in[15:12];
    85: reg_0272 <= imem05_in[15:12];
    endcase
  end

  // REG#273の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0273 <= imem05_in[3:0];
    59: reg_0273 <= imem05_in[3:0];
    86: reg_0273 <= op2_03_out;
    108: reg_0273 <= op2_03_out;
    endcase
  end

  // REG#274の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0274 <= imem05_in[7:4];
    64: reg_0274 <= imem05_in[7:4];
    endcase
  end

  // REG#275の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0275 <= imem05_in[11:8];
    65: reg_0275 <= imem05_in[11:8];
    129: reg_0275 <= imem05_in[11:8];
    endcase
  end

  // REG#276の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0276 <= imem02_in[11:8];
    72: reg_0276 <= imem02_in[11:8];
    129: reg_0276 <= imem02_in[11:8];
    endcase
  end

  // REG#277の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0277 <= imem01_in[3:0];
    78: reg_0277 <= imem01_in[3:0];
    99: reg_0277 <= imem01_in[3:0];
    102: reg_0277 <= imem01_in[3:0];
    108: reg_0277 <= imem01_in[3:0];
    111: reg_0277 <= imem01_in[3:0];
    115: reg_0277 <= op2_00_out;
    endcase
  end

  // REG#278の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0278 <= imem01_in[11:8];
    82: reg_0278 <= imem01_in[11:8];
    86: reg_0278 <= imem05_in[3:0];
    120: reg_0278 <= imem05_in[3:0];
    123: reg_0278 <= imem01_in[11:8];
    125: reg_0278 <= imem05_in[3:0];
    130: reg_0278 <= imem05_in[3:0];
    endcase
  end

  // REG#279の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0279 <= imem02_in[7:4];
    83: reg_0279 <= imem02_in[7:4];
    endcase
  end

  // REG#280の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0280 <= imem02_in[15:12];
    82: reg_0280 <= op2_02_out;
    131: reg_0280 <= op2_02_out;
    endcase
  end

  // REG#281の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0281 <= imem02_in[3:0];
    83: reg_0281 <= imem04_in[3:0];
    endcase
  end

  // REG#282の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0282 <= imem01_in[7:4];
    84: reg_0282 <= op2_01_out;
    87: reg_0282 <= op2_01_out;
    92: reg_0282 <= imem01_in[7:4];
    104: reg_0282 <= imem01_in[7:4];
    113: reg_0282 <= imem01_in[7:4];
    119: reg_0282 <= op2_01_out;
    128: reg_0282 <= op2_01_out;
    endcase
  end

  // REG#283の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0283 <= imem01_in[15:12];
    84: reg_0283 <= op2_02_out;
    88: reg_0283 <= op2_02_out;
    112: reg_0283 <= op2_02_out;
    endcase
  end

  // REG#284の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0284 <= imem07_in[7:4];
    endcase
  end

  // REG#285の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0285 <= imem07_in[11:8];
    endcase
  end

  // REG#286の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0286 <= imem07_in[15:12];
    endcase
  end

  // REG#287の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0287 <= imem07_in[3:0];
    endcase
  end

  // REG#288の入力
  always @ ( posedge clock ) begin
    case ( state )
    17: reg_0288 <= imem03_in[11:8];
    85: reg_0288 <= imem03_in[11:8];
    endcase
  end

  // REG#289の入力
  always @ ( posedge clock ) begin
    case ( state )
    17: reg_0289 <= imem06_in[3:0];
    128: reg_0289 <= imem06_in[3:0];
    endcase
  end

  // REG#290の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0290 <= imem03_in[7:4];
    21: reg_0290 <= imem01_in[3:0];
    84: reg_0290 <= imem01_in[3:0];
    94: reg_0290 <= imem03_in[7:4];
    96: reg_0290 <= imem01_in[3:0];
    121: reg_0290 <= imem03_in[7:4];
    endcase
  end

  // REG#291の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0291 <= imem03_in[11:8];
    21: reg_0291 <= imem01_in[15:12];
    86: reg_0291 <= imem03_in[11:8];
    endcase
  end

  // REG#292の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0292 <= imem04_in[7:4];
    21: reg_0292 <= imem01_in[11:8];
    87: reg_0292 <= imem01_in[11:8];
    endcase
  end

  // REG#293の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0293 <= imem00_in[3:0];
    22: reg_0293 <= imem03_in[3:0];
    48: reg_0293 <= imem00_in[3:0];
    endcase
  end

  // REG#294の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0294 <= imem01_in[11:8];
    22: reg_0294 <= imem02_in[15:12];
    80: reg_0294 <= imem02_in[15:12];
    endcase
  end

  // REG#295の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0295 <= imem06_in[3:0];
    28: reg_0295 <= imem06_in[3:0];
    endcase
  end

  // REG#296の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0296 <= imem06_in[15:12];
    29: reg_0296 <= imem06_in[15:12];
    endcase
  end

  // REG#297の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0297 <= imem07_in[15:12];
    41: reg_0297 <= imem07_in[15:12];
    85: reg_0297 <= imem04_in[7:4];
    endcase
  end

  // REG#298の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0298 <= imem07_in[7:4];
    42: reg_0298 <= imem07_in[7:4];
    58: reg_0298 <= op1_00_out;
    61: reg_0298 <= imem07_in[7:4];
    endcase
  end

  // REG#299の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0299 <= imem07_in[11:8];
    42: reg_0299 <= imem07_in[11:8];
    60: reg_0299 <= imem07_in[11:8];
    endcase
  end

  // REG#300の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0300 <= imem05_in[11:8];
    74: reg_0300 <= imem05_in[11:8];
    endcase
  end

  // REG#301の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0301 <= imem05_in[15:12];
    74: reg_0301 <= imem05_in[15:12];
    endcase
  end

  // REG#302の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0302 <= imem05_in[7:4];
    74: reg_0302 <= imem05_in[7:4];
    endcase
  end

  // REG#303の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0303 <= imem05_in[3:0];
    74: reg_0303 <= imem05_in[3:0];
    endcase
  end

  // REG#304の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0304 <= imem04_in[7:4];
    22: reg_0304 <= imem04_in[7:4];
    95: reg_0304 <= op2_02_out;
    132: reg_0304 <= op2_02_out;
    endcase
  end

  // REG#305の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0305 <= imem04_in[11:8];
    22: reg_0305 <= imem04_in[11:8];
    96: reg_0305 <= imem04_in[11:8];
    97: reg_0305 <= op2_00_out;
    endcase
  end

  // REG#306の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0306 <= imem00_in[15:12];
    22: reg_0306 <= imem02_in[11:8];
    86: reg_0306 <= imem02_in[11:8];
    endcase
  end

  // REG#307の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0307 <= imem01_in[11:8];
    22: reg_0307 <= imem02_in[3:0];
    86: reg_0307 <= imem02_in[3:0];
    endcase
  end

  // REG#308の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0308 <= imem06_in[15:12];
    28: reg_0308 <= imem06_in[15:12];
    endcase
  end

  // REG#309の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0309 <= imem07_in[7:4];
    41: reg_0309 <= imem07_in[7:4];
    86: reg_0309 <= imem07_in[7:4];
    endcase
  end

  // REG#310の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0310 <= imem07_in[15:12];
    43: reg_0310 <= imem07_in[15:12];
    65: reg_0310 <= imem07_in[15:12];
    126: reg_0310 <= imem07_in[15:12];
    endcase
  end

  // REG#311の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0311 <= imem03_in[7:4];
    52: reg_0311 <= imem03_in[7:4];
    89: reg_0311 <= imem03_in[7:4];
    endcase
  end

  // REG#312の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0312 <= imem03_in[11:8];
    52: reg_0312 <= imem03_in[11:8];
    89: reg_0312 <= imem03_in[11:8];
    endcase
  end

  // REG#313の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0313 <= imem03_in[15:12];
    52: reg_0313 <= imem03_in[15:12];
    86: reg_0313 <= imem03_in[15:12];
    endcase
  end

  // REG#314の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0314 <= imem03_in[3:0];
    53: reg_0314 <= imem03_in[3:0];
    61: reg_0314 <= imem03_in[3:0];
    endcase
  end

  // REG#315の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0315 <= imem05_in[11:8];
    61: reg_0315 <= imem05_in[11:8];
    96: reg_0315 <= imem05_in[11:8];
    120: reg_0315 <= imem05_in[11:8];
    125: reg_0315 <= imem05_in[11:8];
    endcase
  end

  // REG#316の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0316 <= imem05_in[3:0];
    61: reg_0316 <= imem06_in[7:4];
    68: reg_0316 <= imem06_in[7:4];
    129: reg_0316 <= imem06_in[7:4];
    endcase
  end

  // REG#317の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0317 <= imem05_in[7:4];
    62: reg_0317 <= imem05_in[7:4];
    endcase
  end

  // REG#318の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0318 <= imem05_in[15:12];
    66: reg_0318 <= imem05_in[15:12];
    endcase
  end

  // REG#319の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0319 <= imem00_in[11:8];
    22: reg_0319 <= imem04_in[15:12];
    94: reg_0319 <= imem00_in[11:8];
    97: reg_0319 <= imem04_in[15:12];
    100: reg_0319 <= imem04_in[15:12];
    103: reg_0319 <= imem00_in[11:8];
    107: reg_0319 <= imem00_in[11:8];
    110: reg_0319 <= imem00_in[11:8];
    114: reg_0319 <= imem04_in[15:12];
    120: reg_0319 <= imem00_in[11:8];
    123: reg_0319 <= imem04_in[15:12];
    128: reg_0319 <= imem00_in[11:8];
    130: reg_0319 <= imem04_in[15:12];
    endcase
  end

  // REG#320の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0320 <= imem01_in[15:12];
    22: reg_0320 <= imem01_in[15:12];
    44: reg_0320 <= imem04_in[7:4];
    129: reg_0320 <= imem01_in[15:12];
    endcase
  end

  // REG#321の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0321 <= imem07_in[3:0];
    23: reg_0321 <= imem07_in[3:0];
    endcase
  end

  // REG#322の入力
  always @ ( posedge clock ) begin
    case ( state )
    19: reg_0322 <= op1_00_out;
    23: reg_0322 <= imem02_in[11:8];
    36: reg_0322 <= op1_00_out;
    88: reg_0322 <= op2_10_out;
    90: reg_0322 <= op2_10_out;
    97: reg_0322 <= imem02_in[11:8];
    103: reg_0322 <= imem02_in[11:8];
    endcase
  end

  // REG#323の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0323 <= imem06_in[7:4];
    29: reg_0323 <= imem06_in[7:4];
    endcase
  end

  // REG#324の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0324 <= imem07_in[15:12];
    36: reg_0324 <= imem07_in[15:12];
    61: reg_0324 <= op1_04_out;
    72: reg_0324 <= imem07_in[15:12];
    74: reg_0324 <= imem07_in[15:12];
    77: reg_0324 <= imem07_in[15:12];
    80: reg_0324 <= imem07_in[15:12];
    81: reg_0324 <= op1_04_out;
    84: reg_0324 <= imem07_in[15:12];
    103: reg_0324 <= imem07_in[15:12];
    114: reg_0324 <= op1_04_out;
    116: reg_0324 <= op1_04_out;
    118: reg_0324 <= op1_04_out;
    120: reg_0324 <= op1_04_out;
    122: reg_0324 <= op1_04_out;
    124: reg_0324 <= op1_04_out;
    127: reg_0324 <= imem07_in[15:12];
    128: reg_0324 <= op1_04_out;
    130: reg_0324 <= op1_04_out;
    endcase
  end

  // REG#325の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0325 <= imem02_in[15:12];
    36: reg_0325 <= op2_00_out;
    39: reg_0325 <= imem02_in[15:12];
    83: reg_0325 <= op2_00_out;
    endcase
  end

  // REG#326の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0326 <= imem02_in[11:8];
    38: reg_0326 <= imem02_in[11:8];
    endcase
  end

  // REG#327の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0327 <= imem02_in[3:0];
    40: reg_0327 <= imem02_in[3:0];
    66: reg_0327 <= imem02_in[3:0];
    108: reg_0327 <= imem02_in[3:0];
    111: reg_0327 <= imem02_in[3:0];
    116: reg_0327 <= imem02_in[3:0];
    120: reg_0327 <= imem02_in[3:0];
    122: reg_0327 <= imem02_in[3:0];
    124: reg_0327 <= imem02_in[3:0];
    126: reg_0327 <= imem02_in[3:0];
    endcase
  end

  // REG#328の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0328 <= imem03_in[3:0];
    41: reg_0328 <= imem03_in[3:0];
    72: reg_0328 <= imem03_in[3:0];
    110: reg_0328 <= imem04_in[11:8];
    114: reg_0328 <= imem03_in[3:0];
    117: reg_0328 <= imem03_in[3:0];
    123: reg_0328 <= imem04_in[11:8];
    endcase
  end

  // REG#329の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0329 <= imem03_in[11:8];
    40: reg_0329 <= imem03_in[11:8];
    60: reg_0329 <= imem03_in[11:8];
    121: reg_0329 <= imem03_in[11:8];
    endcase
  end

  // REG#330の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0330 <= imem03_in[15:12];
    41: reg_0330 <= imem03_in[15:12];
    82: reg_0330 <= imem03_in[15:12];
    128: reg_0330 <= imem03_in[15:12];
    endcase
  end

  // REG#331の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0331 <= imem05_in[11:8];
    46: reg_0331 <= imem05_in[11:8];
    51: reg_0331 <= imem05_in[11:8];
    62: reg_0331 <= imem01_in[11:8];
    74: reg_0331 <= imem01_in[11:8];
    endcase
  end

  // REG#332の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0332 <= imem05_in[15:12];
    46: reg_0332 <= imem05_in[15:12];
    51: reg_0332 <= imem05_in[15:12];
    62: reg_0332 <= imem02_in[7:4];
    74: reg_0332 <= imem02_in[7:4];
    87: reg_0332 <= imem05_in[15:12];
    endcase
  end

  // REG#333の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0333 <= imem05_in[7:4];
    46: reg_0333 <= imem05_in[7:4];
    49: reg_0333 <= imem05_in[7:4];
    56: reg_0333 <= imem05_in[7:4];
    81: reg_0333 <= imem06_in[15:12];
    83: reg_0333 <= imem06_in[15:12];
    86: reg_0333 <= imem05_in[7:4];
    120: reg_0333 <= imem06_in[15:12];
    127: reg_0333 <= imem05_in[7:4];
    endcase
  end

  // REG#334の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0334 <= imem05_in[3:0];
    46: reg_0334 <= imem05_in[3:0];
    54: reg_0334 <= imem05_in[3:0];
    endcase
  end

  // REG#335の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0335 <= imem01_in[7:4];
    52: reg_0335 <= imem01_in[15:12];
    61: reg_0335 <= imem01_in[15:12];
    77: reg_0335 <= imem01_in[7:4];
    81: reg_0335 <= imem01_in[7:4];
    87: reg_0335 <= imem01_in[15:12];
    endcase
  end

  // REG#336の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0336 <= imem04_in[15:12];
    107: reg_0336 <= imem04_in[15:12];
    114: reg_0336 <= op2_01_out;
    endcase
  end

  // REG#337の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0337 <= imem04_in[3:0];
    109: reg_0337 <= imem04_in[3:0];
    111: reg_0337 <= imem04_in[3:0];
    endcase
  end

  // REG#338の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0338 <= imem04_in[7:4];
    109: reg_0338 <= imem05_in[7:4];
    118: reg_0338 <= imem04_in[7:4];
    121: reg_0338 <= imem04_in[7:4];
    123: reg_0338 <= imem05_in[7:4];
    endcase
  end

  // REG#339の入力
  always @ ( posedge clock ) begin
    case ( state )
    20: reg_0339 <= imem04_in[11:8];
    108: reg_0339 <= op2_00_out;
    endcase
  end

  // REG#340の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0340 <= imem04_in[3:0];
    95: reg_0340 <= imem04_in[3:0];
    118: reg_0340 <= imem04_in[3:0];
    122: reg_0340 <= imem05_in[7:4];
    endcase
  end

  // REG#341の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0341 <= imem04_in[7:4];
    42: reg_0341 <= imem04_in[7:4];
    66: reg_0341 <= imem04_in[7:4];
    91: reg_0341 <= imem04_in[7:4];
    96: reg_0341 <= op2_02_out;
    endcase
  end

  // REG#342の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0342 <= imem02_in[7:4];
    44: reg_0342 <= imem04_in[15:12];
    endcase
  end

  // REG#343の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0343 <= imem02_in[3:0];
    43: reg_0343 <= op1_02_out;
    endcase
  end

  // REG#344の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0344 <= imem05_in[3:0];
    45: reg_0344 <= op1_00_out;
    47: reg_0344 <= op1_00_out;
    91: reg_0344 <= imem05_in[3:0];
    endcase
  end

  // REG#345の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0345 <= imem05_in[15:12];
    48: reg_0345 <= imem06_in[3:0];
    50: reg_0345 <= imem05_in[15:12];
    56: reg_0345 <= imem06_in[3:0];
    endcase
  end

  // REG#346の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0346 <= imem05_in[7:4];
    48: reg_0346 <= imem05_in[7:4];
    85: reg_0346 <= imem05_in[7:4];
    endcase
  end

  // REG#347の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0347 <= imem05_in[11:8];
    49: reg_0347 <= imem05_in[11:8];
    58: reg_0347 <= imem05_in[11:8];
    86: reg_0347 <= imem05_in[11:8];
    121: reg_0347 <= imem05_in[11:8];
    127: reg_0347 <= imem05_in[11:8];
    endcase
  end

  // REG#348の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0348 <= imem03_in[15:12];
    59: reg_0348 <= imem03_in[15:12];
    endcase
  end

  // REG#349の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0349 <= imem03_in[7:4];
    61: reg_0349 <= imem03_in[7:4];
    endcase
  end

  // REG#350の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0350 <= imem00_in[3:0];
    63: reg_0350 <= imem03_in[7:4];
    72: reg_0350 <= imem00_in[3:0];
    79: reg_0350 <= imem00_in[3:0];
    81: reg_0350 <= imem00_in[3:0];
    87: reg_0350 <= imem03_in[7:4];
    endcase
  end

  // REG#351の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0351 <= imem00_in[11:8];
    65: reg_0351 <= imem00_in[11:8];
    endcase
  end

  // REG#352の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0352 <= imem00_in[15:12];
    65: reg_0352 <= imem00_in[15:12];
    endcase
  end

  // REG#353の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0353 <= imem00_in[7:4];
    65: reg_0353 <= imem00_in[7:4];
    endcase
  end

  // REG#354の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0354 <= op1_02_out;
    81: reg_0354 <= op1_02_out;
    91: reg_0354 <= op1_02_out;
    93: reg_0354 <= op1_02_out;
    95: reg_0354 <= op1_02_out;
    97: reg_0354 <= op1_02_out;
    99: reg_0354 <= op1_02_out;
    101: reg_0354 <= op1_02_out;
    103: reg_0354 <= op1_02_out;
    105: reg_0354 <= op1_02_out;
    107: reg_0354 <= op1_02_out;
    109: reg_0354 <= op1_02_out;
    111: reg_0354 <= op1_02_out;
    113: reg_0354 <= op1_02_out;
    115: reg_0354 <= op1_02_out;
    117: reg_0354 <= op1_02_out;
    119: reg_0354 <= op1_02_out;
    121: reg_0354 <= op1_02_out;
    endcase
  end

  // REG#355の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0355 <= op1_03_out;
    81: reg_0355 <= op1_03_out;
    83: reg_0355 <= op1_03_out;
    92: reg_0355 <= imem01_in[15:12];
    102: reg_0355 <= imem01_in[15:12];
    107: reg_0355 <= imem01_in[15:12];
    108: reg_0355 <= op1_03_out;
    110: reg_0355 <= op1_03_out;
    112: reg_0355 <= op1_03_out;
    114: reg_0355 <= op1_03_out;
    116: reg_0355 <= op1_03_out;
    118: reg_0355 <= op1_03_out;
    120: reg_0355 <= op1_03_out;
    122: reg_0355 <= op1_03_out;
    124: reg_0355 <= op1_03_out;
    126: reg_0355 <= op1_03_out;
    128: reg_0355 <= op1_03_out;
    130: reg_0355 <= op1_03_out;
    endcase
  end

  // REG#356の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0356 <= op1_06_out;
    85: reg_0356 <= op1_06_out;
    92: reg_0356 <= op1_06_out;
    94: reg_0356 <= op1_06_out;
    96: reg_0356 <= op1_06_out;
    98: reg_0356 <= op1_06_out;
    100: reg_0356 <= op1_06_out;
    102: reg_0356 <= op1_06_out;
    104: reg_0356 <= op1_06_out;
    106: reg_0356 <= op1_06_out;
    108: reg_0356 <= op1_06_out;
    110: reg_0356 <= op1_06_out;
    112: reg_0356 <= op1_06_out;
    114: reg_0356 <= op1_06_out;
    116: reg_0356 <= op1_06_out;
    118: reg_0356 <= op1_06_out;
    120: reg_0356 <= op1_06_out;
    122: reg_0356 <= op1_06_out;
    124: reg_0356 <= op1_06_out;
    126: reg_0356 <= op1_06_out;
    128: reg_0356 <= op1_06_out;
    130: reg_0356 <= op1_06_out;
    endcase
  end

  // REG#357の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0357 <= op1_04_out;
    91: reg_0357 <= op2_00_out;
    101: reg_0357 <= op2_00_out;
    107: reg_0357 <= op2_00_out;
    128: reg_0357 <= op2_00_out;
    endcase
  end

  // REG#358の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0358 <= op1_05_out;
    91: reg_0358 <= op1_05_out;
    93: reg_0358 <= op1_05_out;
    95: reg_0358 <= op1_05_out;
    97: reg_0358 <= op1_05_out;
    99: reg_0358 <= op1_05_out;
    101: reg_0358 <= op1_05_out;
    103: reg_0358 <= op1_05_out;
    105: reg_0358 <= op1_05_out;
    107: reg_0358 <= op1_05_out;
    109: reg_0358 <= op1_05_out;
    111: reg_0358 <= op1_05_out;
    113: reg_0358 <= op1_05_out;
    115: reg_0358 <= op1_05_out;
    117: reg_0358 <= op1_05_out;
    119: reg_0358 <= op1_05_out;
    121: reg_0358 <= op1_05_out;
    123: reg_0358 <= op1_05_out;
    125: reg_0358 <= op1_05_out;
    127: reg_0358 <= op1_05_out;
    129: reg_0358 <= op1_05_out;
    131: reg_0358 <= op1_05_out;
    endcase
  end

  // REG#359の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0359 <= op1_07_out;
    119: reg_0359 <= op1_07_out;
    121: reg_0359 <= op1_07_out;
    123: reg_0359 <= op1_07_out;
    125: reg_0359 <= op1_07_out;
    127: reg_0359 <= op1_07_out;
    129: reg_0359 <= op1_07_out;
    131: reg_0359 <= op1_07_out;
    endcase
  end

  // REG#360の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0360 <= imem01_in[7:4];
    endcase
  end

  // REG#361の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0361 <= imem07_in[11:8];
    endcase
  end

  // REG#362の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0362 <= imem01_in[3:0];
    endcase
  end

  // REG#363の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0363 <= imem01_in[15:12];
    endcase
  end

  // REG#364の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0364 <= op1_08_out;
    131: reg_0364 <= op1_08_out;
    endcase
  end

  // REG#365の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0365 <= imem01_in[11:8];
    endcase
  end

  // REG#366の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0366 <= imem07_in[7:4];
    26: reg_0366 <= imem07_in[7:4];
    endcase
  end

  // REG#367の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0367 <= imem05_in[11:8];
    28: reg_0367 <= imem05_in[11:8];
    73: reg_0367 <= op1_00_out;
    75: reg_0367 <= op1_00_out;
    77: reg_0367 <= op1_00_out;
    90: reg_0367 <= imem05_in[11:8];
    95: reg_0367 <= imem05_in[11:8];
    107: reg_0367 <= imem05_in[11:8];
    109: reg_0367 <= imem05_in[11:8];
    114: reg_0367 <= imem05_in[11:8];
    endcase
  end

  // REG#368の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0368 <= imem04_in[11:8];
    41: reg_0368 <= imem04_in[11:8];
    128: reg_0368 <= imem04_in[11:8];
    endcase
  end

  // REG#369の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0369 <= imem04_in[7:4];
    43: reg_0369 <= imem04_in[7:4];
    65: reg_0369 <= op2_00_out;
    68: reg_0369 <= imem04_in[7:4];
    endcase
  end

  // REG#370の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0370 <= imem04_in[3:0];
    45: reg_0370 <= imem04_in[3:0];
    69: reg_0370 <= op2_00_out;
    72: reg_0370 <= imem04_in[3:0];
    121: reg_0370 <= op2_00_out;
    endcase
  end

  // REG#371の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0371 <= imem06_in[15:12];
    55: reg_0371 <= imem06_in[15:12];
    endcase
  end

  // REG#372の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0372 <= imem06_in[3:0];
    56: reg_0372 <= imem01_in[11:8];
    59: reg_0372 <= imem01_in[11:8];
    65: reg_0372 <= imem01_in[11:8];
    80: reg_0372 <= imem06_in[3:0];
    101: reg_0372 <= imem01_in[11:8];
    109: reg_0372 <= imem06_in[3:0];
    112: reg_0372 <= imem01_in[11:8];
    114: reg_0372 <= imem06_in[3:0];
    127: reg_0372 <= imem01_in[11:8];
    endcase
  end

  // REG#373の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0373 <= imem06_in[7:4];
    58: reg_0373 <= imem06_in[7:4];
    endcase
  end

  // REG#374の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0374 <= imem06_in[11:8];
    59: reg_0374 <= imem06_in[11:8];
    endcase
  end

  // REG#375の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0375 <= imem03_in[3:0];
    64: reg_0375 <= imem03_in[3:0];
    77: reg_0375 <= imem03_in[3:0];
    93: reg_0375 <= imem03_in[3:0];
    endcase
  end

  // REG#376の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0376 <= imem03_in[15:12];
    64: reg_0376 <= imem03_in[15:12];
    79: reg_0376 <= op1_06_out;
    81: reg_0376 <= op1_06_out;
    83: reg_0376 <= op1_06_out;
    92: reg_0376 <= imem03_in[15:12];
    93: reg_0376 <= op1_06_out;
    96: reg_0376 <= imem03_in[15:12];
    98: reg_0376 <= imem03_in[15:12];
    99: reg_0376 <= op1_06_out;
    101: reg_0376 <= op1_06_out;
    103: reg_0376 <= op1_06_out;
    106: reg_0376 <= imem03_in[15:12];
    108: reg_0376 <= imem03_in[15:12];
    109: reg_0376 <= op1_06_out;
    111: reg_0376 <= op1_06_out;
    113: reg_0376 <= op1_06_out;
    116: reg_0376 <= imem03_in[15:12];
    121: reg_0376 <= imem03_in[15:12];
    endcase
  end

  // REG#377の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0377 <= imem03_in[11:8];
    66: reg_0377 <= imem03_in[11:8];
    72: reg_0377 <= imem06_in[11:8];
    77: reg_0377 <= imem03_in[11:8];
    93: reg_0377 <= imem06_in[11:8];
    96: reg_0377 <= imem03_in[11:8];
    98: reg_0377 <= imem03_in[11:8];
    100: reg_0377 <= imem03_in[11:8];
    109: reg_0377 <= imem03_in[11:8];
    119: reg_0377 <= imem03_in[11:8];
    122: reg_0377 <= imem03_in[11:8];
    124: reg_0377 <= imem03_in[11:8];
    endcase
  end

  // REG#378の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0378 <= imem03_in[7:4];
    66: reg_0378 <= imem07_in[15:12];
    69: reg_0378 <= imem03_in[7:4];
    78: reg_0378 <= imem03_in[7:4];
    90: reg_0378 <= imem03_in[7:4];
    124: reg_0378 <= imem03_in[7:4];
    endcase
  end

  // REG#379の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0379 <= imem02_in[7:4];
    67: reg_0379 <= imem02_in[7:4];
    85: reg_0379 <= imem02_in[7:4];
    endcase
  end

  // REG#380の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0380 <= imem02_in[11:8];
    68: reg_0380 <= imem02_in[11:8];
    endcase
  end

  // REG#381の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0381 <= imem02_in[15:12];
    68: reg_0381 <= imem02_in[15:12];
    endcase
  end

  // REG#382の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0382 <= imem02_in[3:0];
    69: reg_0382 <= imem02_in[3:0];
    endcase
  end

  // REG#383の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0383 <= imem01_in[15:12];
    122: reg_0383 <= imem01_in[15:12];
    125: reg_0383 <= imem01_in[15:12];
    endcase
  end

  // REG#384の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0384 <= imem01_in[3:0];
    125: reg_0384 <= imem01_in[3:0];
    endcase
  end

  // REG#385の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0385 <= imem01_in[11:8];
    124: reg_0385 <= imem01_in[11:8];
    endcase
  end

  // REG#386の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0386 <= imem01_in[7:4];
    125: reg_0386 <= imem01_in[7:4];
    endcase
  end

  // REG#387の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0387 <= imem00_in[11:8];
    125: reg_0387 <= imem00_in[11:8];
    endcase
  end

  // REG#388の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0388 <= imem00_in[7:4];
    endcase
  end

  // REG#389の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0389 <= imem00_in[15:12];
    endcase
  end

  // REG#390の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0390 <= imem02_in[11:8];
    37: reg_0390 <= imem02_in[11:8];
    44: reg_0390 <= imem02_in[11:8];
    77: reg_0390 <= imem02_in[11:8];
    endcase
  end

  // REG#391の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0391 <= imem05_in[7:4];
    48: reg_0391 <= imem07_in[11:8];
    52: reg_0391 <= imem05_in[7:4];
    70: reg_0391 <= imem07_in[11:8];
    82: reg_0391 <= imem05_in[7:4];
    endcase
  end

  // REG#392の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0392 <= imem05_in[11:8];
    48: reg_0392 <= imem05_in[11:8];
    83: reg_0392 <= imem05_in[11:8];
    endcase
  end

  // REG#393の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0393 <= imem05_in[15:12];
    48: reg_0393 <= imem07_in[7:4];
    52: reg_0393 <= imem05_in[15:12];
    64: reg_0393 <= imem05_in[15:12];
    endcase
  end

  // REG#394の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0394 <= op1_00_out;
    48: reg_0394 <= imem07_in[3:0];
    52: reg_0394 <= op1_00_out;
    55: reg_0394 <= imem07_in[3:0];
    59: reg_0394 <= op1_00_out;
    89: reg_0394 <= imem07_in[3:0];
    111: reg_0394 <= imem07_in[3:0];
    endcase
  end

  // REG#395の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0395 <= imem05_in[3:0];
    49: reg_0395 <= imem05_in[3:0];
    58: reg_0395 <= imem05_in[3:0];
    85: reg_0395 <= imem05_in[3:0];
    endcase
  end

  // REG#396の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0396 <= imem06_in[11:8];
    59: reg_0396 <= imem04_in[3:0];
    62: reg_0396 <= imem04_in[3:0];
    82: reg_0396 <= imem06_in[11:8];
    96: reg_0396 <= imem04_in[3:0];
    98: reg_0396 <= imem06_in[11:8];
    endcase
  end

  // REG#397の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0397 <= imem06_in[3:0];
    59: reg_0397 <= imem04_in[15:12];
    63: reg_0397 <= imem06_in[3:0];
    87: reg_0397 <= imem06_in[3:0];
    endcase
  end

  // REG#398の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0398 <= imem06_in[7:4];
    59: reg_0398 <= imem06_in[7:4];
    endcase
  end

  // REG#399の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0399 <= imem06_in[15:12];
    59: reg_0399 <= imem02_in[7:4];
    64: reg_0399 <= imem02_in[7:4];
    72: reg_0399 <= imem06_in[15:12];
    78: reg_0399 <= imem02_in[7:4];
    endcase
  end

  // REG#400の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0400 <= imem01_in[7:4];
    87: reg_0400 <= imem01_in[7:4];
    endcase
  end

  // REG#401の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0401 <= imem01_in[15:12];
    95: reg_0401 <= imem01_in[15:12];
    endcase
  end

  // REG#402の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0402 <= imem01_in[3:0];
    97: reg_0402 <= imem01_in[3:0];
    endcase
  end

  // REG#403の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0403 <= imem01_in[11:8];
    97: reg_0403 <= imem01_in[11:8];
    endcase
  end

  // REG#404の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0404 <= imem07_in[3:0];
    127: reg_0404 <= imem07_in[3:0];
    endcase
  end

  // REG#405の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0405 <= imem00_in[15:12];
    endcase
  end

  // REG#406の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0406 <= imem04_in[11:8];
    endcase
  end

  // REG#407の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0407 <= imem04_in[15:12];
    endcase
  end

  // REG#408の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0408 <= imem07_in[7:4];
    endcase
  end

  // REG#409の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0409 <= imem00_in[7:4];
    endcase
  end

  // REG#410の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0410 <= imem00_in[11:8];
    endcase
  end

  // REG#411の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0411 <= imem03_in[3:0];
    endcase
  end

  // REG#412の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0412 <= imem04_in[7:4];
    endcase
  end

  // REG#413の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0413 <= imem07_in[15:12];
    endcase
  end

  // REG#414の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0414 <= imem04_in[3:0];
    endcase
  end

  // REG#415の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0415 <= imem07_in[11:8];
    endcase
  end

  // REG#416の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0416 <= imem00_in[3:0];
    endcase
  end

  // REG#417の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0417 <= op1_01_out;
    endcase
  end

  // REG#418の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0418 <= imem05_in[15:12];
    28: reg_0418 <= imem05_in[15:12];
    75: reg_0418 <= imem05_in[15:12];
    endcase
  end

  // REG#419の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0419 <= imem06_in[11:8];
    28: reg_0419 <= imem06_in[11:8];
    endcase
  end

  // REG#420の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0420 <= imem04_in[3:0];
    34: reg_0420 <= imem04_in[3:0];
    62: reg_0420 <= imem01_in[15:12];
    74: reg_0420 <= imem04_in[3:0];
    endcase
  end

  // REG#421の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0421 <= imem04_in[15:12];
    34: reg_0421 <= imem04_in[15:12];
    62: reg_0421 <= imem04_in[15:12];
    82: reg_0421 <= imem04_in[15:12];
    endcase
  end

  // REG#422の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0422 <= op1_00_out;
    77: reg_0422 <= op2_05_out;
    79: reg_0422 <= op1_00_out;
    81: reg_0422 <= op2_05_out;
    endcase
  end

  // REG#423の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0423 <= op1_01_out;
    95: reg_0423 <= imem02_in[7:4];
    96: reg_0423 <= op1_01_out;
    99: reg_0423 <= imem02_in[7:4];
    101: reg_0423 <= imem02_in[7:4];
    endcase
  end

  // REG#424の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0424 <= op1_02_out;
    endcase
  end

  // REG#425の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0425 <= imem03_in[3:0];
    endcase
  end

  // REG#426の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0426 <= imem03_in[7:4];
    129: reg_0426 <= imem03_in[7:4];
    endcase
  end

  // REG#427の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0427 <= imem03_in[11:8];
    129: reg_0427 <= imem03_in[11:8];
    endcase
  end

  // REG#428の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0428 <= imem00_in[3:0];
    endcase
  end

  // REG#429の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0429 <= imem02_in[11:8];
    endcase
  end

  // REG#430の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0430 <= imem01_in[7:4];
    endcase
  end

  // REG#431の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0431 <= imem00_in[7:4];
    endcase
  end

  // REG#432の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0432 <= imem02_in[3:0];
    endcase
  end

  // REG#433の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0433 <= imem02_in[7:4];
    endcase
  end

  // REG#434の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0434 <= imem01_in[11:8];
    endcase
  end

  // REG#435の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0435 <= imem00_in[15:12];
    endcase
  end

  // REG#436の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0436 <= imem02_in[15:12];
    endcase
  end

  // REG#437の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0437 <= imem07_in[15:12];
    endcase
  end

  // REG#438の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0438 <= imem01_in[15:12];
    endcase
  end

  // REG#439の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0439 <= imem01_in[3:0];
    endcase
  end

  // REG#440の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0440 <= imem00_in[11:8];
    endcase
  end

  // REG#441の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0441 <= imem07_in[3:0];
    endcase
  end

  // REG#442の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0442 <= imem07_in[11:8];
    endcase
  end

  // REG#443の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0443 <= imem03_in[15:12];
    endcase
  end

  // REG#444の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0444 <= imem03_in[11:8];
    34: reg_0444 <= imem03_in[11:8];
    50: reg_0444 <= imem03_in[11:8];
    71: reg_0444 <= imem03_in[11:8];
    83: reg_0444 <= imem03_in[11:8];
    endcase
  end

  // REG#445の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0445 <= imem00_in[11:8];
    35: reg_0445 <= imem05_in[15:12];
    49: reg_0445 <= imem05_in[15:12];
    58: reg_0445 <= imem00_in[11:8];
    76: reg_0445 <= imem00_in[11:8];
    80: reg_0445 <= imem00_in[11:8];
    82: reg_0445 <= imem00_in[11:8];
    97: reg_0445 <= imem00_in[11:8];
    104: reg_0445 <= imem05_in[15:12];
    109: reg_0445 <= imem05_in[15:12];
    116: reg_0445 <= imem00_in[11:8];
    119: reg_0445 <= imem05_in[15:12];
    endcase
  end

  // REG#446の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0446 <= imem01_in[11:8];
    35: reg_0446 <= imem01_in[11:8];
    72: reg_0446 <= op1_12_out;
    74: reg_0446 <= op1_12_out;
    77: reg_0446 <= imem01_in[11:8];
    82: reg_0446 <= op1_12_out;
    91: reg_0446 <= op1_12_out;
    93: reg_0446 <= op1_12_out;
    95: reg_0446 <= op1_12_out;
    97: reg_0446 <= op1_12_out;
    100: reg_0446 <= imem01_in[11:8];
    101: reg_0446 <= op1_12_out;
    104: reg_0446 <= imem01_in[11:8];
    108: reg_0446 <= op1_12_out;
    111: reg_0446 <= imem01_in[11:8];
    116: reg_0446 <= imem01_in[11:8];
    117: reg_0446 <= op1_12_out;
    120: reg_0446 <= op1_12_out;
    122: reg_0446 <= op1_12_out;
    124: reg_0446 <= op1_12_out;
    128: reg_0446 <= op1_12_out;
    130: reg_0446 <= op1_12_out;
    endcase
  end

  // REG#447の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0447 <= op1_00_out;
    37: reg_0447 <= op1_00_out;
    71: reg_0447 <= op1_00_out;
    79: reg_0447 <= imem01_in[11:8];
    80: reg_0447 <= op1_00_out;
    83: reg_0447 <= imem01_in[11:8];
    endcase
  end

  // REG#448の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0448 <= imem03_in[3:0];
    40: reg_0448 <= imem01_in[11:8];
    43: reg_0448 <= imem03_in[3:0];
    60: reg_0448 <= imem01_in[11:8];
    87: reg_0448 <= imem03_in[3:0];
    endcase
  end

  // REG#449の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0449 <= imem05_in[7:4];
    41: reg_0449 <= imem05_in[7:4];
    endcase
  end

  // REG#450の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0450 <= imem05_in[11:8];
    41: reg_0450 <= imem01_in[15:12];
    44: reg_0450 <= imem05_in[11:8];
    73: reg_0450 <= op1_05_out;
    76: reg_0450 <= imem05_in[11:8];
    102: reg_0450 <= imem05_in[11:8];
    endcase
  end

  // REG#451の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0451 <= imem01_in[7:4];
    44: reg_0451 <= imem04_in[3:0];
    endcase
  end

  // REG#452の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0452 <= imem02_in[15:12];
    44: reg_0452 <= imem04_in[11:8];
    endcase
  end

  // REG#453の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0453 <= imem01_in[15:12];
    43: reg_0453 <= op1_03_out;
    endcase
  end

  // REG#454の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0454 <= imem04_in[11:8];
    45: reg_0454 <= imem04_in[11:8];
    70: reg_0454 <= imem04_in[11:8];
    80: reg_0454 <= imem04_in[11:8];
    endcase
  end

  // REG#455の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0455 <= imem02_in[11:8];
    48: reg_0455 <= imem02_in[11:8];
    102: reg_0455 <= imem02_in[11:8];
    endcase
  end

  // REG#456の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0456 <= imem02_in[7:4];
    48: reg_0456 <= imem02_in[7:4];
    100: reg_0456 <= imem02_in[7:4];
    108: reg_0456 <= imem02_in[7:4];
    110: reg_0456 <= imem02_in[7:4];
    114: reg_0456 <= imem02_in[7:4];
    121: reg_0456 <= imem02_in[7:4];
    125: reg_0456 <= imem02_in[7:4];
    endcase
  end

  // REG#457の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0457 <= imem02_in[3:0];
    48: reg_0457 <= imem07_in[15:12];
    54: reg_0457 <= imem02_in[3:0];
    73: reg_0457 <= imem02_in[3:0];
    86: reg_0457 <= imem07_in[15:12];
    endcase
  end

  // REG#458の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0458 <= imem06_in[7:4];
    54: reg_0458 <= imem04_in[3:0];
    67: reg_0458 <= imem06_in[7:4];
    79: reg_0458 <= imem06_in[7:4];
    84: reg_0458 <= imem06_in[7:4];
    87: reg_0458 <= imem03_in[15:12];
    endcase
  end

  // REG#459の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0459 <= imem06_in[11:8];
    54: reg_0459 <= imem00_in[15:12];
    68: reg_0459 <= imem00_in[15:12];
    endcase
  end

  // REG#460の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0460 <= imem06_in[15:12];
    54: reg_0460 <= imem00_in[11:8];
    69: reg_0460 <= imem00_in[11:8];
    endcase
  end

  // REG#461の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0461 <= imem06_in[3:0];
    56: reg_0461 <= imem07_in[7:4];
    68: reg_0461 <= imem07_in[7:4];
    113: reg_0461 <= imem06_in[3:0];
    118: reg_0461 <= imem06_in[3:0];
    121: reg_0461 <= imem06_in[3:0];
    124: reg_0461 <= imem07_in[7:4];
    129: reg_0461 <= imem06_in[3:0];
    endcase
  end

  // REG#462の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0462 <= imem04_in[15:12];
    57: reg_0462 <= imem04_in[15:12];
    endcase
  end

  // REG#463の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0463 <= imem04_in[3:0];
    58: reg_0463 <= imem04_in[3:0];
    62: reg_0463 <= imem01_in[3:0];
    74: reg_0463 <= imem01_in[3:0];
    endcase
  end

  // REG#464の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0464 <= imem04_in[7:4];
    58: reg_0464 <= imem04_in[7:4];
    62: reg_0464 <= imem04_in[7:4];
    82: reg_0464 <= imem01_in[3:0];
    87: reg_0464 <= imem01_in[3:0];
    endcase
  end

  // REG#465の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0465 <= imem07_in[7:4];
    endcase
  end

  // REG#466の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0466 <= imem04_in[3:0];
    35: reg_0466 <= imem04_in[3:0];
    72: reg_0466 <= imem06_in[7:4];
    78: reg_0466 <= imem06_in[7:4];
    87: reg_0466 <= imem05_in[11:8];
    endcase
  end

  // REG#467の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0467 <= imem04_in[7:4];
    34: reg_0467 <= imem04_in[7:4];
    57: reg_0467 <= op1_03_out;
    73: reg_0467 <= op1_03_out;
    89: reg_0467 <= imem04_in[7:4];
    94: reg_0467 <= imem04_in[7:4];
    115: reg_0467 <= op2_02_out;
    endcase
  end

  // REG#468の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0468 <= imem01_in[3:0];
    36: reg_0468 <= imem01_in[3:0];
    endcase
  end

  // REG#469の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0469 <= imem01_in[11:8];
    36: reg_0469 <= imem01_in[11:8];
    endcase
  end

  // REG#470の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0470 <= imem04_in[15:12];
    43: reg_0470 <= imem04_in[15:12];
    69: reg_0470 <= imem04_in[15:12];
    73: reg_0470 <= imem04_in[15:12];
    endcase
  end

  // REG#471の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0471 <= imem04_in[11:8];
    46: reg_0471 <= imem04_in[11:8];
    endcase
  end

  // REG#472の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0472 <= imem02_in[3:0];
    55: reg_0472 <= imem02_in[3:0];
    endcase
  end

  // REG#473の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0473 <= imem02_in[7:4];
    56: reg_0473 <= imem02_in[7:4];
    86: reg_0473 <= imem02_in[7:4];
    endcase
  end

  // REG#474の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0474 <= imem02_in[15:12];
    56: reg_0474 <= imem02_in[15:12];
    87: reg_0474 <= imem02_in[15:12];
    96: reg_0474 <= imem02_in[15:12];
    98: reg_0474 <= op2_00_out;
    endcase
  end

  // REG#475の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0475 <= imem02_in[11:8];
    56: reg_0475 <= imem02_in[11:8];
    88: reg_0475 <= op2_11_out;
    92: reg_0475 <= imem02_in[11:8];
    103: reg_0475 <= imem06_in[11:8];
    105: reg_0475 <= imem06_in[11:8];
    107: reg_0475 <= imem06_in[11:8];
    110: reg_0475 <= imem02_in[11:8];
    114: reg_0475 <= imem02_in[11:8];
    119: reg_0475 <= imem02_in[11:8];
    121: reg_0475 <= imem02_in[11:8];
    126: reg_0475 <= imem06_in[11:8];
    endcase
  end

  // REG#476の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0476 <= imem00_in[3:0];
    66: reg_0476 <= imem00_in[3:0];
    endcase
  end

  // REG#477の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0477 <= imem05_in[3:0];
    75: reg_0477 <= imem05_in[3:0];
    endcase
  end

  // REG#478の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0478 <= imem03_in[15:12];
    91: reg_0478 <= imem07_in[11:8];
    95: reg_0478 <= imem07_in[11:8];
    endcase
  end

  // REG#479の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0479 <= imem03_in[11:8];
    90: reg_0479 <= op2_09_out;
    95: reg_0479 <= imem03_in[11:8];
    97: reg_0479 <= imem03_in[11:8];
    99: reg_0479 <= imem03_in[11:8];
    101: reg_0479 <= imem03_in[11:8];
    107: reg_0479 <= imem03_in[11:8];
    116: reg_0479 <= imem03_in[11:8];
    127: reg_0479 <= imem03_in[11:8];
    endcase
  end

  // REG#480の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0480 <= imem03_in[3:0];
    91: reg_0480 <= imem03_in[3:0];
    92: reg_0480 <= op2_01_out;
    116: reg_0480 <= imem03_in[3:0];
    122: reg_0480 <= op2_01_out;
    endcase
  end

  // REG#481の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0481 <= imem03_in[7:4];
    90: reg_0481 <= op2_11_out;
    97: reg_0481 <= imem03_in[7:4];
    98: reg_0481 <= op2_01_out;
    endcase
  end

  // REG#482の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0482 <= op1_01_out;
    109: reg_0482 <= op2_00_out;
    endcase
  end

  // REG#483の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0483 <= imem07_in[3:0];
    endcase
  end

  // REG#484の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0484 <= imem07_in[7:4];
    endcase
  end

  // REG#485の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0485 <= imem00_in[3:0];
    36: reg_0485 <= imem00_in[3:0];
    53: reg_0485 <= op1_00_out;
    70: reg_0485 <= imem00_in[3:0];
    endcase
  end

  // REG#486の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0486 <= imem01_in[15:12];
    35: reg_0486 <= imem01_in[15:12];
    84: reg_0486 <= imem00_in[3:0];
    86: reg_0486 <= imem00_in[3:0];
    endcase
  end

  // REG#487の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0487 <= imem04_in[7:4];
    41: reg_0487 <= imem04_in[7:4];
    endcase
  end

  // REG#488の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0488 <= imem04_in[3:0];
    42: reg_0488 <= imem04_in[3:0];
    67: reg_0488 <= imem04_in[3:0];
    84: reg_0488 <= imem04_in[3:0];
    endcase
  end

  // REG#489の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0489 <= imem05_in[3:0];
    46: reg_0489 <= imem07_in[15:12];
    49: reg_0489 <= imem07_in[15:12];
    endcase
  end

  // REG#490の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0490 <= imem05_in[11:8];
    46: reg_0490 <= imem07_in[7:4];
    52: reg_0490 <= imem07_in[7:4];
    69: reg_0490 <= imem07_in[7:4];
    76: reg_0490 <= imem07_in[7:4];
    81: reg_0490 <= imem07_in[7:4];
    93: reg_0490 <= imem07_in[7:4];
    97: reg_0490 <= imem07_in[7:4];
    99: reg_0490 <= imem05_in[11:8];
    101: reg_0490 <= imem05_in[11:8];
    104: reg_0490 <= imem07_in[7:4];
    105: reg_0490 <= op2_01_out;
    122: reg_0490 <= imem07_in[7:4];
    123: reg_0490 <= op2_01_out;
    endcase
  end

  // REG#491の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0491 <= imem05_in[15:12];
    46: reg_0491 <= imem07_in[11:8];
    52: reg_0491 <= imem07_in[11:8];
    69: reg_0491 <= imem07_in[11:8];
    76: reg_0491 <= imem07_in[11:8];
    82: reg_0491 <= imem05_in[15:12];
    endcase
  end

  // REG#492の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0492 <= imem05_in[7:4];
    46: reg_0492 <= imem00_in[7:4];
    65: reg_0492 <= imem05_in[7:4];
    endcase
  end

  // REG#493の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0493 <= imem04_in[15:12];
    48: reg_0493 <= imem04_in[15:12];
    58: reg_0493 <= imem04_in[15:12];
    64: reg_0493 <= imem04_in[15:12];
    125: reg_0493 <= imem04_in[15:12];
    endcase
  end

  // REG#494の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0494 <= imem02_in[15:12];
    55: reg_0494 <= imem02_in[15:12];
    endcase
  end

  // REG#495の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0495 <= imem02_in[7:4];
    55: reg_0495 <= imem02_in[7:4];
    126: reg_0495 <= imem02_in[7:4];
    endcase
  end

  // REG#496の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0496 <= imem02_in[11:8];
    56: reg_0496 <= imem07_in[3:0];
    69: reg_0496 <= imem02_in[11:8];
    endcase
  end

  // REG#497の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0497 <= imem02_in[3:0];
    58: reg_0497 <= imem02_in[3:0];
    89: reg_0497 <= imem02_in[3:0];
    109: reg_0497 <= imem02_in[3:0];
    endcase
  end

  // REG#498の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0498 <= op1_00_out;
    76: reg_0498 <= op1_00_out;
    79: reg_0498 <= imem07_in[11:8];
    81: reg_0498 <= imem07_in[11:8];
    85: reg_0498 <= imem07_in[11:8];
    86: reg_0498 <= op1_00_out;
    89: reg_0498 <= imem07_in[11:8];
    114: reg_0498 <= imem07_in[11:8];
    116: reg_0498 <= imem07_in[11:8];
    123: reg_0498 <= imem07_in[11:8];
    endcase
  end

  // REG#499の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0499 <= op1_01_out;
    79: reg_0499 <= op1_01_out;
    81: reg_0499 <= op1_01_out;
    92: reg_0499 <= imem02_in[7:4];
    103: reg_0499 <= op2_02_out;
    117: reg_0499 <= imem02_in[7:4];
    119: reg_0499 <= imem02_in[7:4];
    120: reg_0499 <= op2_02_out;
    endcase
  end

  // REG#500の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0500 <= op1_03_out;
    80: reg_0500 <= op1_03_out;
    83: reg_0500 <= imem04_in[7:4];
    endcase
  end

  // REG#501の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0501 <= op1_04_out;
    82: reg_0501 <= imem00_in[15:12];
    100: reg_0501 <= imem00_in[15:12];
    endcase
  end

  // REG#502の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0502 <= op1_05_out;
    81: reg_0502 <= op1_05_out;
    83: reg_0502 <= op1_05_out;
    91: reg_0502 <= op2_02_out;
    104: reg_0502 <= op2_02_out;
    119: reg_0502 <= op2_02_out;
    129: reg_0502 <= op2_02_out;
    endcase
  end

  // REG#503の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0503 <= op1_08_out;
    85: reg_0503 <= op1_08_out;
    87: reg_0503 <= op1_08_out;
    89: reg_0503 <= op1_08_out;
    91: reg_0503 <= op1_08_out;
    93: reg_0503 <= op1_08_out;
    95: reg_0503 <= op1_08_out;
    97: reg_0503 <= op1_08_out;
    99: reg_0503 <= op1_08_out;
    101: reg_0503 <= op1_08_out;
    103: reg_0503 <= op1_08_out;
    105: reg_0503 <= op1_08_out;
    107: reg_0503 <= op1_08_out;
    109: reg_0503 <= op1_08_out;
    111: reg_0503 <= op1_08_out;
    113: reg_0503 <= op1_08_out;
    115: reg_0503 <= op1_08_out;
    117: reg_0503 <= op1_08_out;
    119: reg_0503 <= op1_08_out;
    121: reg_0503 <= op1_08_out;
    123: reg_0503 <= op1_08_out;
    125: reg_0503 <= op1_08_out;
    127: reg_0503 <= op1_08_out;
    129: reg_0503 <= op1_08_out;
    endcase
  end

  // REG#504の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0504 <= imem03_in[7:4];
    88: reg_0504 <= imem03_in[7:4];
    98: reg_0504 <= op2_02_out;
    endcase
  end

  // REG#505の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0505 <= imem03_in[3:0];
    88: reg_0505 <= imem03_in[3:0];
    100: reg_0505 <= imem03_in[3:0];
    111: reg_0505 <= imem03_in[3:0];
    endcase
  end

  // REG#506の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0506 <= imem03_in[11:8];
    88: reg_0506 <= imem03_in[11:8];
    96: reg_0506 <= op2_03_out;
    endcase
  end

  // REG#507の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0507 <= imem03_in[15:12];
    88: reg_0507 <= imem03_in[15:12];
    101: reg_0507 <= imem03_in[15:12];
    103: reg_0507 <= imem04_in[7:4];
    105: reg_0507 <= imem04_in[7:4];
    107: reg_0507 <= imem04_in[7:4];
    112: reg_0507 <= imem03_in[15:12];
    endcase
  end

  // REG#508の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0508 <= op1_02_out;
    90: reg_0508 <= op2_12_out;
    97: reg_0508 <= op2_01_out;
    endcase
  end

  // REG#509の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0509 <= op1_06_out;
    90: reg_0509 <= op1_06_out;
    94: reg_0509 <= imem07_in[15:12];
    98: reg_0509 <= imem07_in[15:12];
    99: reg_0509 <= op2_01_out;
    101: reg_0509 <= op2_01_out;
    108: reg_0509 <= op2_01_out;
    endcase
  end

  // REG#510の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0510 <= op1_07_out;
    91: reg_0510 <= op1_07_out;
    93: reg_0510 <= op1_07_out;
    95: reg_0510 <= op1_07_out;
    97: reg_0510 <= op1_07_out;
    99: reg_0510 <= op1_07_out;
    101: reg_0510 <= op1_07_out;
    103: reg_0510 <= op1_07_out;
    105: reg_0510 <= op1_07_out;
    107: reg_0510 <= op1_07_out;
    109: reg_0510 <= op1_07_out;
    111: reg_0510 <= op1_07_out;
    113: reg_0510 <= op1_07_out;
    115: reg_0510 <= op1_07_out;
    117: reg_0510 <= op1_07_out;
    120: reg_0510 <= op1_07_out;
    122: reg_0510 <= op1_07_out;
    124: reg_0510 <= op1_07_out;
    126: reg_0510 <= op1_07_out;
    128: reg_0510 <= op1_07_out;
    130: reg_0510 <= op1_07_out;
    endcase
  end

  // REG#511の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0511 <= op1_09_out;
    92: reg_0511 <= op1_09_out;
    94: reg_0511 <= op1_09_out;
    96: reg_0511 <= op1_09_out;
    98: reg_0511 <= op1_09_out;
    100: reg_0511 <= op1_09_out;
    102: reg_0511 <= op1_09_out;
    104: reg_0511 <= op1_09_out;
    106: reg_0511 <= op1_09_out;
    108: reg_0511 <= op1_09_out;
    110: reg_0511 <= op1_09_out;
    112: reg_0511 <= op1_09_out;
    114: reg_0511 <= op1_09_out;
    116: reg_0511 <= op1_09_out;
    118: reg_0511 <= op1_09_out;
    121: reg_0511 <= op1_09_out;
    123: reg_0511 <= op1_09_out;
    125: reg_0511 <= op1_09_out;
    127: reg_0511 <= op1_09_out;
    129: reg_0511 <= op1_09_out;
    131: reg_0511 <= op1_09_out;
    endcase
  end

  // REG#512の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0512 <= op1_10_out;
    94: reg_0512 <= op1_10_out;
    96: reg_0512 <= op1_10_out;
    98: reg_0512 <= op1_10_out;
    100: reg_0512 <= op1_10_out;
    102: reg_0512 <= op1_10_out;
    104: reg_0512 <= op1_10_out;
    106: reg_0512 <= op1_10_out;
    108: reg_0512 <= op1_10_out;
    110: reg_0512 <= op1_10_out;
    112: reg_0512 <= op1_10_out;
    114: reg_0512 <= op1_10_out;
    116: reg_0512 <= op1_10_out;
    118: reg_0512 <= op1_10_out;
    122: reg_0512 <= op1_10_out;
    124: reg_0512 <= op1_10_out;
    126: reg_0512 <= op1_10_out;
    128: reg_0512 <= op1_10_out;
    130: reg_0512 <= op1_10_out;
    endcase
  end

  // REG#513の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0513 <= op1_11_out;
    94: reg_0513 <= op1_11_out;
    96: reg_0513 <= op1_11_out;
    98: reg_0513 <= op1_11_out;
    100: reg_0513 <= op1_11_out;
    102: reg_0513 <= op1_11_out;
    104: reg_0513 <= op1_11_out;
    106: reg_0513 <= op1_11_out;
    108: reg_0513 <= op1_11_out;
    110: reg_0513 <= op1_11_out;
    112: reg_0513 <= op1_11_out;
    114: reg_0513 <= op1_11_out;
    116: reg_0513 <= op1_11_out;
    118: reg_0513 <= op1_11_out;
    121: reg_0513 <= op1_11_out;
    123: reg_0513 <= op1_11_out;
    125: reg_0513 <= op1_11_out;
    127: reg_0513 <= op1_11_out;
    129: reg_0513 <= op1_11_out;
    endcase
  end

  // REG#514の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0514 <= op1_12_out;
    98: reg_0514 <= op1_12_out;
    100: reg_0514 <= op1_12_out;
    102: reg_0514 <= op1_12_out;
    104: reg_0514 <= op1_12_out;
    106: reg_0514 <= op2_00_out;
    124: reg_0514 <= op2_00_out;
    endcase
  end

  // REG#515の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0515 <= op1_13_out;
    99: reg_0515 <= op1_13_out;
    101: reg_0515 <= op1_13_out;
    103: reg_0515 <= op1_13_out;
    106: reg_0515 <= op1_13_out;
    108: reg_0515 <= op1_13_out;
    110: reg_0515 <= op1_13_out;
    112: reg_0515 <= op1_13_out;
    114: reg_0515 <= op1_13_out;
    117: reg_0515 <= op1_13_out;
    120: reg_0515 <= op1_13_out;
    122: reg_0515 <= op1_13_out;
    124: reg_0515 <= op1_13_out;
    127: reg_0515 <= op1_13_out;
    129: reg_0515 <= op1_13_out;
    endcase
  end

  // REG#516の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0516 <= op1_14_out;
    102: reg_0516 <= op1_14_out;
    105: reg_0516 <= op1_14_out;
    107: reg_0516 <= op1_14_out;
    110: reg_0516 <= op1_14_out;
    113: reg_0516 <= op1_14_out;
    115: reg_0516 <= op1_14_out;
    117: reg_0516 <= op1_14_out;
    120: reg_0516 <= op1_14_out;
    123: reg_0516 <= op1_14_out;
    126: reg_0516 <= op1_14_out;
    129: reg_0516 <= op1_14_out;
    endcase
  end

  // REG#517の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0517 <= op1_15_out;
    112: reg_0517 <= op1_15_out;
    115: reg_0517 <= op1_15_out;
    117: reg_0517 <= op1_15_out;
    120: reg_0517 <= op1_15_out;
    123: reg_0517 <= op1_15_out;
    126: reg_0517 <= op1_15_out;
    129: reg_0517 <= op1_15_out;
    endcase
  end

  // REG#518の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0518 <= imem07_in[7:4];
    121: reg_0518 <= imem07_in[7:4];
    126: reg_0518 <= imem07_in[7:4];
    endcase
  end

  // REG#519の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0519 <= imem07_in[3:0];
    126: reg_0519 <= imem07_in[3:0];
    endcase
  end

  // REG#520の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0520 <= imem07_in[15:12];
    endcase
  end

  // REG#521の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0521 <= imem07_in[11:8];
    endcase
  end

  // REG#522の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0522 <= imem06_in[3:0];
    endcase
  end

  // REG#523の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0523 <= imem00_in[11:8];
    35: reg_0523 <= imem05_in[7:4];
    49: reg_0523 <= imem00_in[11:8];
    endcase
  end

  // REG#524の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0524 <= imem00_in[3:0];
    35: reg_0524 <= imem06_in[15:12];
    53: reg_0524 <= imem00_in[3:0];
    65: reg_0524 <= imem06_in[15:12];
    67: reg_0524 <= imem00_in[3:0];
    endcase
  end

  // REG#525の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0525 <= imem03_in[7:4];
    37: reg_0525 <= imem03_in[7:4];
    68: reg_0525 <= imem03_in[7:4];
    87: reg_0525 <= op2_00_out;
    89: reg_0525 <= op2_00_out;
    103: reg_0525 <= imem03_in[7:4];
    105: reg_0525 <= op2_00_out;
    120: reg_0525 <= op2_00_out;
    endcase
  end

  // REG#526の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0526 <= imem06_in[3:0];
    57: reg_0526 <= imem06_in[3:0];
    endcase
  end

  // REG#527の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0527 <= imem06_in[15:12];
    57: reg_0527 <= imem06_in[15:12];
    endcase
  end

  // REG#528の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0528 <= imem06_in[7:4];
    57: reg_0528 <= imem06_in[7:4];
    endcase
  end

  // REG#529の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0529 <= imem06_in[11:8];
    57: reg_0529 <= imem06_in[11:8];
    endcase
  end

  // REG#530の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0530 <= imem02_in[7:4];
    60: reg_0530 <= imem02_in[7:4];
    79: reg_0530 <= imem02_in[7:4];
    112: reg_0530 <= imem02_in[7:4];
    113: reg_0530 <= op2_00_out;
    endcase
  end

  // REG#531の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0531 <= imem02_in[15:12];
    60: reg_0531 <= imem04_in[3:0];
    67: reg_0531 <= imem02_in[15:12];
    85: reg_0531 <= imem04_in[3:0];
    endcase
  end

  // REG#532の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0532 <= imem02_in[3:0];
    60: reg_0532 <= imem02_in[3:0];
    77: reg_0532 <= imem02_in[3:0];
    endcase
  end

  // REG#533の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0533 <= imem02_in[11:8];
    60: reg_0533 <= imem02_in[11:8];
    72: reg_0533 <= op1_13_out;
    74: reg_0533 <= op1_13_out;
    76: reg_0533 <= op1_13_out;
    89: reg_0533 <= op1_13_out;
    91: reg_0533 <= op1_13_out;
    93: reg_0533 <= op1_13_out;
    95: reg_0533 <= op1_13_out;
    98: reg_0533 <= imem02_in[11:8];
    100: reg_0533 <= imem02_in[11:8];
    109: reg_0533 <= imem02_in[11:8];
    endcase
  end

  // REG#534の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0534 <= imem04_in[11:8];
    61: reg_0534 <= imem04_in[11:8];
    90: reg_0534 <= op2_13_out;
    99: reg_0534 <= op2_02_out;
    102: reg_0534 <= op2_02_out;
    113: reg_0534 <= imem04_in[11:8];
    127: reg_0534 <= op2_02_out;
    endcase
  end

  // REG#535の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0535 <= imem04_in[3:0];
    61: reg_0535 <= op1_11_out;
    79: reg_0535 <= op1_11_out;
    81: reg_0535 <= op1_11_out;
    83: reg_0535 <= op1_11_out;
    86: reg_0535 <= imem04_in[3:0];
    119: reg_0535 <= op1_11_out;
    123: reg_0535 <= imem04_in[3:0];
    endcase
  end

  // REG#536の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0536 <= imem04_in[15:12];
    64: reg_0536 <= imem06_in[11:8];
    76: reg_0536 <= imem04_in[15:12];
    endcase
  end

  // REG#537の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0537 <= imem04_in[7:4];
    66: reg_0537 <= imem07_in[7:4];
    69: reg_0537 <= imem04_in[7:4];
    79: reg_0537 <= imem07_in[7:4];
    81: reg_0537 <= imem04_in[7:4];
    endcase
  end

  // REG#538の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0538 <= imem05_in[7:4];
    73: reg_0538 <= op1_09_out;
    75: reg_0538 <= op1_09_out;
    77: reg_0538 <= op1_09_out;
    79: reg_0538 <= op1_09_out;
    81: reg_0538 <= op1_09_out;
    91: reg_0538 <= op1_09_out;
    94: reg_0538 <= imem05_in[7:4];
    95: reg_0538 <= op1_09_out;
    97: reg_0538 <= op1_09_out;
    100: reg_0538 <= imem05_in[7:4];
    105: reg_0538 <= imem05_in[7:4];
    108: reg_0538 <= imem05_in[7:4];
    110: reg_0538 <= imem05_in[7:4];
    117: reg_0538 <= imem05_in[7:4];
    130: reg_0538 <= op1_09_out;
    endcase
  end

  // REG#539の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0539 <= imem05_in[15:12];
    74: reg_0539 <= op1_08_out;
    78: reg_0539 <= imem05_in[15:12];
    79: reg_0539 <= op1_08_out;
    81: reg_0539 <= op1_08_out;
    91: reg_0539 <= op2_03_out;
    105: reg_0539 <= op2_03_out;
    124: reg_0539 <= op1_08_out;
    126: reg_0539 <= op1_08_out;
    128: reg_0539 <= op1_08_out;
    130: reg_0539 <= op1_08_out;
    endcase
  end

  // REG#540の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0540 <= imem05_in[3:0];
    77: reg_0540 <= op2_06_out;
    80: reg_0540 <= op2_06_out;
    113: reg_0540 <= imem05_in[3:0];
    endcase
  end

  // REG#541の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0541 <= imem05_in[11:8];
    78: reg_0541 <= imem03_in[11:8];
    90: reg_0541 <= imem03_in[11:8];
    123: reg_0541 <= imem05_in[11:8];
    126: reg_0541 <= imem03_in[11:8];
    128: reg_0541 <= imem03_in[11:8];
    endcase
  end

  // REG#542の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0542 <= op1_00_out;
    endcase
  end

  // REG#543の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0543 <= op1_01_out;
    118: reg_0543 <= op1_01_out;
    endcase
  end

  // REG#544の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0544 <= op1_02_out;
    endcase
  end

  // REG#545の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0545 <= op1_03_out;
    endcase
  end

  // REG#546の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0546 <= op1_04_out;
    126: reg_0546 <= op1_04_out;
    endcase
  end

  // REG#547の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0547 <= imem01_in[3:0];
    127: reg_0547 <= imem01_in[3:0];
    endcase
  end

  // REG#548の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0548 <= imem01_in[15:12];
    endcase
  end

  // REG#549の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0549 <= imem01_in[7:4];
    endcase
  end

  // REG#550の入力
  always @ ( posedge clock ) begin
    case ( state )
    30: reg_0550 <= imem01_in[11:8];
    endcase
  end

  // REG#551の入力
  always @ ( posedge clock ) begin
    case ( state )
    29: reg_0551 <= op1_05_out;
    endcase
  end

  // REG#552の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0552 <= imem04_in[15:12];
    35: reg_0552 <= imem04_in[15:12];
    72: reg_0552 <= imem00_in[11:8];
    79: reg_0552 <= imem00_in[11:8];
    83: reg_0552 <= imem00_in[11:8];
    85: reg_0552 <= imem04_in[15:12];
    endcase
  end

  // REG#553の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0553 <= imem01_in[11:8];
    35: reg_0553 <= imem02_in[11:8];
    53: reg_0553 <= imem01_in[11:8];
    69: reg_0553 <= imem01_in[11:8];
    124: reg_0553 <= imem02_in[11:8];
    126: reg_0553 <= imem01_in[11:8];
    endcase
  end

  // REG#554の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0554 <= imem00_in[3:0];
    52: reg_0554 <= imem00_in[3:0];
    81: reg_0554 <= imem00_in[15:12];
    87: reg_0554 <= imem00_in[15:12];
    endcase
  end

  // REG#555の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0555 <= imem00_in[11:8];
    52: reg_0555 <= imem00_in[11:8];
    81: reg_0555 <= imem00_in[11:8];
    86: reg_0555 <= imem00_in[11:8];
    endcase
  end

  // REG#556の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0556 <= imem03_in[15:12];
    54: reg_0556 <= imem03_in[15:12];
    61: reg_0556 <= op1_14_out;
    80: reg_0556 <= op1_14_out;
    90: reg_0556 <= op1_14_out;
    93: reg_0556 <= imem03_in[15:12];
    endcase
  end

  // REG#557の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0557 <= imem03_in[11:8];
    54: reg_0557 <= imem03_in[11:8];
    66: reg_0557 <= imem03_in[15:12];
    71: reg_0557 <= imem03_in[15:12];
    80: reg_0557 <= imem03_in[11:8];
    endcase
  end

  // REG#558の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0558 <= imem03_in[3:0];
    56: reg_0558 <= imem03_in[3:0];
    endcase
  end

  // REG#559の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0559 <= imem03_in[7:4];
    57: reg_0559 <= imem03_in[7:4];
    72: reg_0559 <= imem03_in[7:4];
    119: reg_0559 <= imem03_in[7:4];
    123: reg_0559 <= imem03_in[7:4];
    endcase
  end

  // REG#560の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0560 <= imem02_in[15:12];
    71: reg_0560 <= imem07_in[11:8];
    74: reg_0560 <= op1_09_out;
    78: reg_0560 <= imem07_in[11:8];
    82: reg_0560 <= imem07_in[11:8];
    85: reg_0560 <= imem02_in[15:12];
    endcase
  end

  // REG#561の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0561 <= imem02_in[11:8];
    71: reg_0561 <= imem02_in[11:8];
    endcase
  end

  // REG#562の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0562 <= imem02_in[7:4];
    72: reg_0562 <= imem00_in[15:12];
    79: reg_0562 <= imem00_in[15:12];
    83: reg_0562 <= imem05_in[15:12];
    endcase
  end

  // REG#563の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0563 <= imem02_in[3:0];
    71: reg_0563 <= op1_13_out;
    79: reg_0563 <= op1_13_out;
    82: reg_0563 <= imem02_in[3:0];
    endcase
  end

  // REG#564の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0564 <= imem05_in[11:8];
    80: reg_0564 <= imem05_in[11:8];
    endcase
  end

  // REG#565の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0565 <= imem05_in[7:4];
    80: reg_0565 <= op2_00_out;
    103: reg_0565 <= op2_00_out;
    115: reg_0565 <= imem05_in[7:4];
    endcase
  end

  // REG#566の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0566 <= imem05_in[15:12];
    81: reg_0566 <= imem05_in[15:12];
    endcase
  end

  // REG#567の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0567 <= imem05_in[3:0];
    81: reg_0567 <= op2_01_out;
    117: reg_0567 <= op2_01_out;
    123: reg_0567 <= imem05_in[3:0];
    129: reg_0567 <= op2_01_out;
    endcase
  end

  // REG#568の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0568 <= imem06_in[3:0];
    endcase
  end

  // REG#569の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0569 <= imem06_in[11:8];
    endcase
  end

  // REG#570の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0570 <= imem06_in[15:12];
    endcase
  end

  // REG#571の入力
  always @ ( posedge clock ) begin
    case ( state )
    31: reg_0571 <= imem06_in[7:4];
    endcase
  end

  // REG#572の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0572 <= imem01_in[15:12];
    36: reg_0572 <= imem01_in[15:12];
    endcase
  end

  // REG#573の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0573 <= imem03_in[15:12];
    37: reg_0573 <= imem03_in[15:12];
    68: reg_0573 <= imem03_in[15:12];
    83: reg_0573 <= imem03_in[15:12];
    endcase
  end

  // REG#574の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0574 <= imem04_in[11:8];
    48: reg_0574 <= imem04_in[11:8];
    55: reg_0574 <= imem04_in[11:8];
    endcase
  end

  // REG#575の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0575 <= imem05_in[3:0];
    48: reg_0575 <= imem01_in[11:8];
    63: reg_0575 <= imem05_in[3:0];
    endcase
  end

  // REG#576の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0576 <= imem05_in[15:12];
    48: reg_0576 <= imem01_in[7:4];
    63: reg_0576 <= imem01_in[7:4];
    73: reg_0576 <= imem05_in[15:12];
    95: reg_0576 <= imem01_in[7:4];
    endcase
  end

  // REG#577の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0577 <= imem04_in[3:0];
    49: reg_0577 <= imem04_in[3:0];
    51: reg_0577 <= imem04_in[3:0];
    56: reg_0577 <= imem04_in[3:0];
    84: reg_0577 <= imem01_in[7:4];
    90: reg_0577 <= imem04_in[3:0];
    94: reg_0577 <= imem04_in[3:0];
    118: reg_0577 <= imem01_in[7:4];
    endcase
  end

  // REG#578の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0578 <= imem05_in[7:4];
    51: reg_0578 <= imem05_in[7:4];
    61: reg_0578 <= imem05_in[7:4];
    93: reg_0578 <= op2_00_out;
    119: reg_0578 <= op2_00_out;
    127: reg_0578 <= op2_00_out;
    endcase
  end

  // REG#579の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0579 <= imem05_in[11:8];
    52: reg_0579 <= imem05_in[11:8];
    70: reg_0579 <= imem05_in[11:8];
    94: reg_0579 <= imem05_in[11:8];
    97: reg_0579 <= imem05_in[11:8];
    100: reg_0579 <= imem05_in[11:8];
    105: reg_0579 <= imem05_in[11:8];
    108: reg_0579 <= imem05_in[11:8];
    110: reg_0579 <= imem05_in[11:8];
    117: reg_0579 <= imem05_in[11:8];
    endcase
  end

  // REG#580の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0580 <= imem00_in[15:12];
    52: reg_0580 <= imem00_in[15:12];
    78: reg_0580 <= imem00_in[15:12];
    endcase
  end

  // REG#581の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0581 <= imem00_in[3:0];
    53: reg_0581 <= op1_02_out;
    70: reg_0581 <= op1_02_out;
    79: reg_0581 <= op1_10_out;
    81: reg_0581 <= op1_10_out;
    91: reg_0581 <= op2_04_out;
    110: reg_0581 <= imem00_in[3:0];
    112: reg_0581 <= imem00_in[3:0];
    117: reg_0581 <= imem00_in[3:0];
    120: reg_0581 <= op1_10_out;
    123: reg_0581 <= imem00_in[3:0];
    endcase
  end

  // REG#582の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0582 <= imem04_in[15:12];
    54: reg_0582 <= imem04_in[15:12];
    68: reg_0582 <= imem04_in[15:12];
    endcase
  end

  // REG#583の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0583 <= imem06_in[7:4];
    55: reg_0583 <= imem06_in[7:4];
    endcase
  end

  // REG#584の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0584 <= imem06_in[15:12];
    58: reg_0584 <= imem06_in[15:12];
    endcase
  end

  // REG#585の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0585 <= imem06_in[3:0];
    58: reg_0585 <= imem06_in[3:0];
    endcase
  end

  // REG#586の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0586 <= imem06_in[11:8];
    58: reg_0586 <= imem06_in[11:8];
    endcase
  end

  // REG#587の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0587 <= imem02_in[15:12];
    71: reg_0587 <= imem05_in[15:12];
    78: reg_0587 <= op2_00_out;
    81: reg_0587 <= op2_00_out;
    115: reg_0587 <= imem02_in[15:12];
    116: reg_0587 <= op2_00_out;
    endcase
  end

  // REG#588の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0588 <= imem02_in[3:0];
    71: reg_0588 <= imem02_in[3:0];
    endcase
  end

  // REG#589の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0589 <= imem02_in[11:8];
    72: reg_0589 <= imem05_in[7:4];
    89: reg_0589 <= imem05_in[7:4];
    91: reg_0589 <= imem05_in[7:4];
    endcase
  end

  // REG#590の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0590 <= imem02_in[7:4];
    73: reg_0590 <= imem02_in[7:4];
    88: reg_0590 <= imem02_in[7:4];
    94: reg_0590 <= imem02_in[7:4];
    97: reg_0590 <= imem02_in[7:4];
    105: reg_0590 <= imem02_in[7:4];
    106: reg_0590 <= op2_03_out;
    128: reg_0590 <= op2_03_out;
    endcase
  end

  // REG#591の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0591 <= imem07_in[7:4];
    endcase
  end

  // REG#592の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0592 <= imem07_in[15:12];
    endcase
  end

  // REG#593の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0593 <= imem07_in[3:0];
    endcase
  end

  // REG#594の入力
  always @ ( posedge clock ) begin
    case ( state )
    32: reg_0594 <= op1_00_out;
    38: reg_0594 <= imem04_in[7:4];
    39: reg_0594 <= op1_00_out;
    48: reg_0594 <= imem04_in[7:4];
    57: reg_0594 <= op1_00_out;
    78: reg_0594 <= op2_01_out;
    82: reg_0594 <= op2_01_out;
    129: reg_0594 <= imem04_in[7:4];
    endcase
  end

  // REG#595の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0595 <= imem04_in[7:4];
    41: reg_0595 <= imem01_in[3:0];
    52: reg_0595 <= imem04_in[7:4];
    60: reg_0595 <= imem04_in[7:4];
    66: reg_0595 <= imem01_in[3:0];
    88: reg_0595 <= imem01_in[3:0];
    endcase
  end

  // REG#596の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0596 <= imem04_in[11:8];
    42: reg_0596 <= imem04_in[11:8];
    69: reg_0596 <= imem04_in[11:8];
    78: reg_0596 <= op2_03_out;
    84: reg_0596 <= op2_03_out;
    89: reg_0596 <= op2_03_out;
    99: reg_0596 <= op2_00_out;
    endcase
  end

  // REG#597の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0597 <= imem03_in[7:4];
    44: reg_0597 <= imem03_in[7:4];
    112: reg_0597 <= imem03_in[7:4];
    endcase
  end

  // REG#598の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0598 <= imem04_in[3:0];
    46: reg_0598 <= imem04_in[3:0];
    endcase
  end

  // REG#599の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0599 <= imem04_in[15:12];
    46: reg_0599 <= imem04_in[15:12];
    endcase
  end

  // REG#600の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0600 <= imem03_in[3:0];
    48: reg_0600 <= imem03_in[3:0];
    56: reg_0600 <= imem07_in[11:8];
    68: reg_0600 <= op2_00_out;
    70: reg_0600 <= op2_00_out;
    72: reg_0600 <= op2_00_out;
    74: reg_0600 <= op2_00_out;
    76: reg_0600 <= op2_00_out;
    89: reg_0600 <= imem03_in[3:0];
    endcase
  end

  // REG#601の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0601 <= imem05_in[3:0];
    48: reg_0601 <= imem01_in[15:12];
    64: reg_0601 <= imem05_in[3:0];
    endcase
  end

  // REG#602の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0602 <= imem05_in[11:8];
    48: reg_0602 <= imem01_in[3:0];
    63: reg_0602 <= imem05_in[11:8];
    endcase
  end

  // REG#603の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0603 <= imem05_in[15:12];
    47: reg_0603 <= op1_02_out;
    76: reg_0603 <= op1_02_out;
    78: reg_0603 <= op1_02_out;
    80: reg_0603 <= op1_02_out;
    91: reg_0603 <= imem05_in[15:12];
    endcase
  end

  // REG#604の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0604 <= imem05_in[7:4];
    47: reg_0604 <= op1_03_out;
    83: reg_0604 <= imem05_in[7:4];
    endcase
  end

  // REG#605の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0605 <= imem02_in[7:4];
    50: reg_0605 <= imem02_in[7:4];
    72: reg_0605 <= op2_01_out;
    74: reg_0605 <= op2_01_out;
    77: reg_0605 <= op2_01_out;
    120: reg_0605 <= op2_01_out;
    endcase
  end

  // REG#606の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0606 <= imem02_in[3:0];
    50: reg_0606 <= imem02_in[3:0];
    76: reg_0606 <= op1_15_out;
    78: reg_0606 <= op1_15_out;
    90: reg_0606 <= op1_15_out;
    93: reg_0606 <= imem02_in[3:0];
    94: reg_0606 <= op1_15_out;
    97: reg_0606 <= op1_15_out;
    100: reg_0606 <= op1_15_out;
    103: reg_0606 <= op1_15_out;
    106: reg_0606 <= op1_15_out;
    110: reg_0606 <= imem02_in[3:0];
    114: reg_0606 <= imem02_in[3:0];
    118: reg_0606 <= imem02_in[3:0];
    130: reg_0606 <= op1_15_out;
    endcase
  end

  // REG#607の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0607 <= imem02_in[11:8];
    50: reg_0607 <= imem02_in[11:8];
    79: reg_0607 <= imem02_in[11:8];
    113: reg_0607 <= op2_01_out;
    endcase
  end

  // REG#608の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0608 <= imem02_in[15:12];
    50: reg_0608 <= imem02_in[15:12];
    72: reg_0608 <= imem02_in[15:12];
    endcase
  end

  // REG#609の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0609 <= imem01_in[15:12];
    54: reg_0609 <= imem01_in[15:12];
    73: reg_0609 <= imem01_in[15:12];
    endcase
  end

  // REG#610の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0610 <= imem01_in[11:8];
    55: reg_0610 <= imem01_in[11:8];
    endcase
  end

  // REG#611の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0611 <= imem01_in[3:0];
    59: reg_0611 <= imem01_in[3:0];
    65: reg_0611 <= imem01_in[3:0];
    72: reg_0611 <= op1_02_out;
    76: reg_0611 <= imem01_in[3:0];
    79: reg_0611 <= imem01_in[3:0];
    81: reg_0611 <= imem01_in[3:0];
    86: reg_0611 <= op1_02_out;
    88: reg_0611 <= op1_02_out;
    91: reg_0611 <= imem01_in[3:0];
    93: reg_0611 <= op2_02_out;
    121: reg_0611 <= op2_02_out;
    endcase
  end

  // REG#612の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0612 <= imem01_in[7:4];
    59: reg_0612 <= imem02_in[11:8];
    64: reg_0612 <= imem02_in[11:8];
    71: reg_0612 <= imem01_in[7:4];
    endcase
  end

  // REG#613の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0613 <= imem00_in[3:0];
    74: reg_0613 <= imem00_in[3:0];
    78: reg_0613 <= imem00_in[3:0];
    127: reg_0613 <= imem00_in[3:0];
    endcase
  end

  // REG#614の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0614 <= imem00_in[15:12];
    76: reg_0614 <= imem00_in[15:12];
    77: reg_0614 <= op1_14_out;
    90: reg_0614 <= op2_14_out;
    99: reg_0614 <= op1_14_out;
    101: reg_0614 <= op1_14_out;
    104: reg_0614 <= imem00_in[15:12];
    106: reg_0614 <= op1_14_out;
    109: reg_0614 <= op1_14_out;
    111: reg_0614 <= op1_14_out;
    113: reg_0614 <= op2_02_out;
    endcase
  end

  // REG#615の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0615 <= imem00_in[11:8];
    75: reg_0615 <= op1_08_out;
    78: reg_0615 <= imem00_in[11:8];
    endcase
  end

  // REG#616の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0616 <= imem00_in[7:4];
    77: reg_0616 <= imem00_in[7:4];
    87: reg_0616 <= imem00_in[7:4];
    endcase
  end

  // REG#617の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0617 <= imem06_in[11:8];
    127: reg_0617 <= imem06_in[11:8];
    endcase
  end

  // REG#618の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0618 <= imem07_in[11:8];
    endcase
  end

  // REG#619の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0619 <= imem06_in[7:4];
    endcase
  end

  // REG#620の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0620 <= imem07_in[15:12];
    endcase
  end

  // REG#621の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0621 <= imem07_in[7:4];
    endcase
  end

  // REG#622の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0622 <= imem06_in[3:0];
    endcase
  end

  // REG#623の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0623 <= imem07_in[3:0];
    endcase
  end

  // REG#624の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0624 <= imem06_in[15:12];
    endcase
  end

  // REG#625の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0625 <= op1_00_out;
    38: reg_0625 <= imem04_in[3:0];
    47: reg_0625 <= op1_05_out;
    86: reg_0625 <= op1_05_out;
    88: reg_0625 <= op1_05_out;
    91: reg_0625 <= imem04_in[3:0];
    92: reg_0625 <= op1_05_out;
    94: reg_0625 <= op1_05_out;
    96: reg_0625 <= op1_05_out;
    99: reg_0625 <= imem04_in[3:0];
    100: reg_0625 <= op1_05_out;
    102: reg_0625 <= op1_05_out;
    105: reg_0625 <= imem04_in[3:0];
    106: reg_0625 <= op1_05_out;
    108: reg_0625 <= op1_05_out;
    110: reg_0625 <= op1_05_out;
    112: reg_0625 <= op1_05_out;
    115: reg_0625 <= imem04_in[3:0];
    116: reg_0625 <= op1_05_out;
    118: reg_0625 <= op1_05_out;
    120: reg_0625 <= op1_05_out;
    122: reg_0625 <= op1_05_out;
    124: reg_0625 <= op1_05_out;
    126: reg_0625 <= op1_05_out;
    128: reg_0625 <= op1_05_out;
    130: reg_0625 <= op1_05_out;
    endcase
  end

  // REG#626の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0626 <= imem02_in[3:0];
    45: reg_0626 <= imem02_in[3:0];
    71: reg_0626 <= imem05_in[11:8];
    79: reg_0626 <= imem02_in[3:0];
    112: reg_0626 <= imem02_in[3:0];
    115: reg_0626 <= imem02_in[3:0];
    117: reg_0626 <= imem02_in[3:0];
    121: reg_0626 <= imem02_in[3:0];
    125: reg_0626 <= imem02_in[3:0];
    endcase
  end

  // REG#627の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0627 <= imem03_in[7:4];
    45: reg_0627 <= imem03_in[7:4];
    endcase
  end

  // REG#628の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0628 <= imem02_in[11:8];
    47: reg_0628 <= op1_01_out;
    88: reg_0628 <= op1_01_out;
    91: reg_0628 <= imem02_in[11:8];
    endcase
  end

  // REG#629の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0629 <= imem02_in[7:4];
    51: reg_0629 <= imem02_in[7:4];
    56: reg_0629 <= imem07_in[15:12];
    69: reg_0629 <= imem02_in[7:4];
    endcase
  end

  // REG#630の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0630 <= imem03_in[3:0];
    51: reg_0630 <= imem03_in[3:0];
    54: reg_0630 <= imem03_in[3:0];
    67: reg_0630 <= imem03_in[3:0];
    71: reg_0630 <= imem05_in[7:4];
    80: reg_0630 <= imem05_in[7:4];
    endcase
  end

  // REG#631の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0631 <= imem02_in[15:12];
    52: reg_0631 <= imem05_in[3:0];
    62: reg_0631 <= imem02_in[15:12];
    72: reg_0631 <= imem05_in[3:0];
    91: reg_0631 <= imem02_in[15:12];
    endcase
  end

  // REG#632の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0632 <= imem03_in[15:12];
    52: reg_0632 <= imem02_in[11:8];
    65: reg_0632 <= imem02_in[11:8];
    82: reg_0632 <= imem02_in[11:8];
    endcase
  end

  // REG#633の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0633 <= imem04_in[11:8];
    57: reg_0633 <= op1_04_out;
    74: reg_0633 <= imem04_in[11:8];
    endcase
  end

  // REG#634の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0634 <= imem06_in[3:0];
    59: reg_0634 <= imem01_in[15:12];
    68: reg_0634 <= op1_12_out;
    73: reg_0634 <= op1_12_out;
    88: reg_0634 <= op1_12_out;
    90: reg_0634 <= op1_12_out;
    92: reg_0634 <= op1_12_out;
    94: reg_0634 <= op1_12_out;
    97: reg_0634 <= imem01_in[15:12];
    endcase
  end

  // REG#635の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0635 <= imem06_in[7:4];
    58: reg_0635 <= op1_02_out;
    80: reg_0635 <= imem06_in[7:4];
    100: reg_0635 <= imem06_in[7:4];
    103: reg_0635 <= imem06_in[3:0];
    105: reg_0635 <= imem01_in[3:0];
    107: reg_0635 <= imem06_in[7:4];
    109: reg_0635 <= imem01_in[3:0];
    119: reg_0635 <= imem06_in[3:0];
    121: reg_0635 <= imem06_in[7:4];
    123: reg_0635 <= imem01_in[3:0];
    128: reg_0635 <= imem01_in[3:0];
    endcase
  end

  // REG#636の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0636 <= imem06_in[11:8];
    60: reg_0636 <= imem06_in[11:8];
    endcase
  end

  // REG#637の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0637 <= imem06_in[15:12];
    60: reg_0637 <= imem06_in[15:12];
    endcase
  end

  // REG#638の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0638 <= imem00_in[7:4];
    63: reg_0638 <= imem03_in[11:8];
    71: reg_0638 <= op1_02_out;
    89: reg_0638 <= imem00_in[7:4];
    96: reg_0638 <= imem00_in[7:4];
    99: reg_0638 <= imem00_in[7:4];
    102: reg_0638 <= imem00_in[7:4];
    123: reg_0638 <= imem03_in[11:8];
    endcase
  end

  // REG#639の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0639 <= op1_02_out;
    62: reg_0639 <= op1_02_out;
    82: reg_0639 <= op1_02_out;
    84: reg_0639 <= op1_02_out;
    91: reg_0639 <= op2_05_out;
    110: reg_0639 <= op2_01_out;
    endcase
  end

  // REG#640の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0640 <= imem00_in[15:12];
    64: reg_0640 <= imem03_in[11:8];
    77: reg_0640 <= imem00_in[15:12];
    86: reg_0640 <= imem00_in[15:12];
    endcase
  end

  // REG#641の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0641 <= imem00_in[3:0];
    64: reg_0641 <= op1_13_out;
    66: reg_0641 <= op1_13_out;
    93: reg_0641 <= op2_04_out;
    123: reg_0641 <= op1_13_out;
    125: reg_0641 <= op1_13_out;
    128: reg_0641 <= imem00_in[3:0];
    130: reg_0641 <= op1_13_out;
    endcase
  end

  // REG#642の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0642 <= imem00_in[11:8];
    64: reg_0642 <= op1_14_out;
    66: reg_0642 <= op1_14_out;
    93: reg_0642 <= op1_14_out;
    95: reg_0642 <= op1_14_out;
    97: reg_0642 <= op1_14_out;
    101: reg_0642 <= imem00_in[11:8];
    102: reg_0642 <= op2_01_out;
    111: reg_0642 <= op2_01_out;
    endcase
  end

  // REG#643の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0643 <= op1_11_out;
    66: reg_0643 <= op1_11_out;
    93: reg_0643 <= op2_05_out;
    128: reg_0643 <= op1_11_out;
    endcase
  end

  // REG#644の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0644 <= op1_04_out;
    78: reg_0644 <= op2_04_out;
    85: reg_0644 <= op1_04_out;
    92: reg_0644 <= op2_04_out;
    128: reg_0644 <= op2_04_out;
    endcase
  end

  // REG#645の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0645 <= op1_07_out;
    79: reg_0645 <= op1_07_out;
    90: reg_0645 <= op1_07_out;
    92: reg_0645 <= op1_07_out;
    94: reg_0645 <= op1_07_out;
    96: reg_0645 <= op1_07_out;
    98: reg_0645 <= op1_07_out;
    100: reg_0645 <= op1_07_out;
    102: reg_0645 <= op1_07_out;
    104: reg_0645 <= op1_07_out;
    106: reg_0645 <= op1_07_out;
    108: reg_0645 <= op1_07_out;
    110: reg_0645 <= op1_07_out;
    112: reg_0645 <= op1_07_out;
    114: reg_0645 <= op1_07_out;
    116: reg_0645 <= op1_07_out;
    118: reg_0645 <= op1_07_out;
    endcase
  end

  // REG#646の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0646 <= imem05_in[3:0];
    81: reg_0646 <= op2_03_out;
    121: reg_0646 <= imem05_in[3:0];
    126: reg_0646 <= op2_03_out;
    endcase
  end

  // REG#647の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0647 <= op1_08_out;
    82: reg_0647 <= op1_08_out;
    91: reg_0647 <= op2_06_out;
    112: reg_0647 <= op1_08_out;
    114: reg_0647 <= op1_08_out;
    116: reg_0647 <= op1_08_out;
    118: reg_0647 <= op1_08_out;
    120: reg_0647 <= op1_08_out;
    122: reg_0647 <= op1_08_out;
    endcase
  end

  // REG#648の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0648 <= imem05_in[7:4];
    84: reg_0648 <= imem05_in[7:4];
    125: reg_0648 <= imem05_in[7:4];
    endcase
  end

  // REG#649の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0649 <= imem05_in[11:8];
    84: reg_0649 <= imem05_in[11:8];
    122: reg_0649 <= imem05_in[11:8];
    endcase
  end

  // REG#650の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0650 <= imem05_in[15:12];
    83: reg_0650 <= op1_00_out;
    91: reg_0650 <= op2_07_out;
    113: reg_0650 <= imem05_in[15:12];
    120: reg_0650 <= imem05_in[15:12];
    125: reg_0650 <= imem05_in[15:12];
    endcase
  end

  // REG#651の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0651 <= op1_09_out;
    84: reg_0651 <= op1_09_out;
    91: reg_0651 <= op2_08_out;
    113: reg_0651 <= op1_09_out;
    115: reg_0651 <= op1_09_out;
    117: reg_0651 <= op1_09_out;
    119: reg_0651 <= op1_09_out;
    122: reg_0651 <= op1_09_out;
    124: reg_0651 <= op1_09_out;
    126: reg_0651 <= op1_09_out;
    128: reg_0651 <= op1_09_out;
    endcase
  end

  // REG#652の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0652 <= op1_10_out;
    85: reg_0652 <= op1_10_out;
    87: reg_0652 <= op1_10_out;
    89: reg_0652 <= op2_01_out;
    96: reg_0652 <= op2_01_out;
    endcase
  end

  // REG#653の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0653 <= op1_01_out;
    89: reg_0653 <= imem01_in[7:4];
    93: reg_0653 <= op2_06_out;
    endcase
  end

  // REG#654の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0654 <= op1_03_out;
    89: reg_0654 <= op1_03_out;
    94: reg_0654 <= op1_03_out;
    96: reg_0654 <= op1_03_out;
    98: reg_0654 <= op1_03_out;
    100: reg_0654 <= op1_03_out;
    102: reg_0654 <= op1_03_out;
    104: reg_0654 <= op1_03_out;
    106: reg_0654 <= op1_03_out;
    114: reg_0654 <= op2_02_out;
    endcase
  end

  // REG#655の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0655 <= op1_05_out;
    89: reg_0655 <= op1_05_out;
    94: reg_0655 <= op2_00_out;
    126: reg_0655 <= op2_00_out;
    endcase
  end

  // REG#656の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0656 <= op1_06_out;
    90: reg_0656 <= op2_15_out;
    101: reg_0656 <= imem04_in[11:8];
    102: reg_0656 <= op2_03_out;
    114: reg_0656 <= imem04_in[11:8];
    120: reg_0656 <= op2_03_out;
    endcase
  end

  // REG#657の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0657 <= op1_12_out;
    96: reg_0657 <= op1_12_out;
    99: reg_0657 <= op1_12_out;
    101: reg_0657 <= op2_02_out;
    109: reg_0657 <= op2_02_out;
    endcase
  end

  // REG#658の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0658 <= op1_13_out;
    96: reg_0658 <= op1_13_out;
    98: reg_0658 <= op1_13_out;
    102: reg_0658 <= op1_13_out;
    105: reg_0658 <= op1_13_out;
    107: reg_0658 <= op1_13_out;
    111: reg_0658 <= op1_13_out;
    113: reg_0658 <= op1_13_out;
    115: reg_0658 <= op1_13_out;
    118: reg_0658 <= op1_13_out;
    121: reg_0658 <= op1_13_out;
    126: reg_0658 <= op1_13_out;
    endcase
  end

  // REG#659の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0659 <= op1_14_out;
    96: reg_0659 <= op1_14_out;
    98: reg_0659 <= op1_14_out;
    103: reg_0659 <= imem02_in[15:12];
    127: reg_0659 <= imem02_in[15:12];
    130: reg_0659 <= op1_14_out;
    endcase
  end

  // REG#660の入力
  always @ ( posedge clock ) begin
    case ( state )
    33: reg_0660 <= op1_15_out;
    104: reg_0660 <= op1_15_out;
    107: reg_0660 <= op1_15_out;
    110: reg_0660 <= op1_15_out;
    113: reg_0660 <= op1_15_out;
    116: reg_0660 <= op1_15_out;
    119: reg_0660 <= op1_15_out;
    122: reg_0660 <= op1_15_out;
    125: reg_0660 <= op1_15_out;
    128: reg_0660 <= op1_15_out;
    endcase
  end

  // REG#661の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0661 <= imem07_in[7:4];
    endcase
  end

  // REG#662の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0662 <= imem01_in[3:0];
    endcase
  end

  // REG#663の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0663 <= imem07_in[11:8];
    endcase
  end

  // REG#664の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0664 <= imem07_in[15:12];
    endcase
  end

  // REG#665の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0665 <= imem07_in[3:0];
    endcase
  end

  // REG#666の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0666 <= imem02_in[3:0];
    56: reg_0666 <= imem02_in[3:0];
    87: reg_0666 <= imem02_in[3:0];
    96: reg_0666 <= imem02_in[3:0];
    99: reg_0666 <= imem02_in[3:0];
    101: reg_0666 <= imem02_in[3:0];
    endcase
  end

  // REG#667の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0667 <= imem02_in[7:4];
    55: reg_0667 <= imem07_in[11:8];
    61: reg_0667 <= imem07_in[11:8];
    endcase
  end

  // REG#668の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0668 <= imem02_in[15:12];
    55: reg_0668 <= imem07_in[15:12];
    61: reg_0668 <= op1_15_out;
    81: reg_0668 <= op1_15_out;
    84: reg_0668 <= op1_15_out;
    88: reg_0668 <= imem07_in[15:12];
    92: reg_0668 <= imem02_in[15:12];
    104: reg_0668 <= imem02_in[15:12];
    106: reg_0668 <= imem07_in[15:12];
    108: reg_0668 <= imem07_in[15:12];
    110: reg_0668 <= imem07_in[15:12];
    113: reg_0668 <= imem02_in[15:12];
    116: reg_0668 <= imem07_in[15:12];
    123: reg_0668 <= imem02_in[15:12];
    127: reg_0668 <= op1_15_out;
    endcase
  end

  // REG#669の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0669 <= imem06_in[11:8];
    57: reg_0669 <= imem02_in[11:8];
    60: reg_0669 <= imem00_in[15:12];
    73: reg_0669 <= imem06_in[11:8];
    81: reg_0669 <= imem06_in[11:8];
    83: reg_0669 <= imem06_in[11:8];
    87: reg_0669 <= imem02_in[11:8];
    96: reg_0669 <= imem00_in[15:12];
    98: reg_0669 <= imem00_in[15:12];
    104: reg_0669 <= imem02_in[11:8];
    106: reg_0669 <= imem06_in[11:8];
    108: reg_0669 <= imem06_in[11:8];
    110: reg_0669 <= imem00_in[15:12];
    114: reg_0669 <= imem06_in[11:8];
    128: reg_0669 <= imem06_in[11:8];
    endcase
  end

  // REG#670の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0670 <= imem06_in[7:4];
    58: reg_0670 <= op1_03_out;
    79: reg_0670 <= op1_03_out;
    90: reg_0670 <= op1_03_out;
    93: reg_0670 <= imem06_in[7:4];
    97: reg_0670 <= imem06_in[7:4];
    118: reg_0670 <= imem06_in[7:4];
    120: reg_0670 <= imem06_in[7:4];
    endcase
  end

  // REG#671の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0671 <= imem06_in[3:0];
    58: reg_0671 <= op1_04_out;
    79: reg_0671 <= op1_04_out;
    90: reg_0671 <= op2_01_out;
    126: reg_0671 <= op2_01_out;
    endcase
  end

  // REG#672の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0672 <= imem07_in[7:4];
    60: reg_0672 <= imem00_in[7:4];
    74: reg_0672 <= imem07_in[7:4];
    78: reg_0672 <= imem07_in[7:4];
    82: reg_0672 <= imem00_in[7:4];
    100: reg_0672 <= op2_00_out;
    104: reg_0672 <= imem00_in[7:4];
    112: reg_0672 <= op2_00_out;
    endcase
  end

  // REG#673の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0673 <= imem07_in[3:0];
    62: reg_0673 <= imem07_in[3:0];
    85: reg_0673 <= imem03_in[7:4];
    endcase
  end

  // REG#674の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0674 <= imem07_in[11:8];
    64: reg_0674 <= imem07_in[11:8];
    80: reg_0674 <= imem07_in[11:8];
    81: reg_0674 <= op2_04_out;
    121: reg_0674 <= imem07_in[11:8];
    endcase
  end

  // REG#675の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0675 <= imem03_in[15:12];
    71: reg_0675 <= imem05_in[3:0];
    79: reg_0675 <= op2_01_out;
    88: reg_0675 <= imem07_in[11:8];
    93: reg_0675 <= op2_01_out;
    122: reg_0675 <= imem07_in[11:8];
    124: reg_0675 <= imem05_in[3:0];
    126: reg_0675 <= imem03_in[15:12];
    127: reg_0675 <= op2_01_out;
    endcase
  end

  // REG#676の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0676 <= imem04_in[7:4];
    71: reg_0676 <= op1_03_out;
    88: reg_0676 <= op1_03_out;
    90: reg_0676 <= op2_02_out;
    endcase
  end

  // REG#677の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0677 <= imem03_in[3:0];
    71: reg_0677 <= op1_05_out;
    89: reg_0677 <= imem01_in[11:8];
    93: reg_0677 <= imem01_in[11:8];
    95: reg_0677 <= imem03_in[3:0];
    97: reg_0677 <= imem03_in[3:0];
    98: reg_0677 <= op1_05_out;
    100: reg_0677 <= op2_01_out;
    105: reg_0677 <= imem03_in[3:0];
    109: reg_0677 <= imem03_in[3:0];
    118: reg_0677 <= imem01_in[11:8];
    130: reg_0677 <= op2_01_out;
    endcase
  end

  // REG#678の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0678 <= imem03_in[7:4];
    71: reg_0678 <= op1_08_out;
    89: reg_0678 <= op2_02_out;
    97: reg_0678 <= op2_02_out;
    endcase
  end

  // REG#679の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0679 <= imem01_in[7:4];
    80: reg_0679 <= imem01_in[7:4];
    82: reg_0679 <= imem01_in[7:4];
    87: reg_0679 <= op2_03_out;
    93: reg_0679 <= op2_03_out;
    124: reg_0679 <= imem01_in[7:4];
    131: reg_0679 <= op2_03_out;
    endcase
  end

  // REG#680の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0680 <= op1_02_out;
    80: reg_0680 <= op2_02_out;
    106: reg_0680 <= op2_02_out;
    126: reg_0680 <= op2_02_out;
    endcase
  end

  // REG#681の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0681 <= imem04_in[11:8];
    84: reg_0681 <= imem04_in[11:8];
    endcase
  end

  // REG#682の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0682 <= op1_04_out;
    83: reg_0682 <= op1_04_out;
    92: reg_0682 <= op1_04_out;
    94: reg_0682 <= op2_01_out;
    endcase
  end

  // REG#683の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0683 <= op1_00_out;
    89: reg_0683 <= op2_04_out;
    100: reg_0683 <= op2_02_out;
    105: reg_0683 <= op2_02_out;
    122: reg_0683 <= op2_02_out;
    endcase
  end

  // REG#684の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0684 <= op1_01_out;
    91: reg_0684 <= imem02_in[7:4];
    endcase
  end

  // REG#685の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0685 <= op1_03_out;
    90: reg_0685 <= op2_03_out;
    endcase
  end

  // REG#686の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0686 <= op1_05_out;
    94: reg_0686 <= op2_02_out;
    128: reg_0686 <= op2_02_out;
    endcase
  end

  // REG#687の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0687 <= op1_06_out;
    107: reg_0687 <= op1_06_out;
    115: reg_0687 <= op1_06_out;
    117: reg_0687 <= op1_06_out;
    119: reg_0687 <= op1_06_out;
    121: reg_0687 <= op1_06_out;
    123: reg_0687 <= op1_06_out;
    125: reg_0687 <= op1_06_out;
    127: reg_0687 <= op1_06_out;
    129: reg_0687 <= op1_06_out;
    131: reg_0687 <= op1_06_out;
    endcase
  end

  // REG#688の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0688 <= op1_07_out;
    endcase
  end

  // REG#689の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0689 <= op1_08_out;
    endcase
  end

  // REG#690の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0690 <= op1_09_out;
    endcase
  end

  // REG#691の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0691 <= op1_10_out;
    endcase
  end

  // REG#692の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0692 <= op1_11_out;
    endcase
  end

  // REG#693の入力
  always @ ( posedge clock ) begin
    case ( state )
    34: reg_0693 <= op1_12_out;
    endcase
  end

  // REG#694の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0694 <= op1_00_out;
    38: reg_0694 <= imem04_in[15:12];
    48: reg_0694 <= op1_00_out;
    61: reg_0694 <= imem04_in[15:12];
    92: reg_0694 <= imem04_in[15:12];
    111: reg_0694 <= imem04_in[15:12];
    endcase
  end

  // REG#695の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0695 <= imem04_in[3:0];
    41: reg_0695 <= imem01_in[11:8];
    52: reg_0695 <= imem04_in[3:0];
    58: reg_0695 <= imem01_in[11:8];
    65: reg_0695 <= imem02_in[7:4];
    80: reg_0695 <= imem02_in[7:4];
    endcase
  end

  // REG#696の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0696 <= imem04_in[15:12];
    46: reg_0696 <= imem06_in[7:4];
    67: reg_0696 <= imem04_in[15:12];
    88: reg_0696 <= imem04_in[15:12];
    90: reg_0696 <= imem04_in[15:12];
    95: reg_0696 <= imem06_in[7:4];
    endcase
  end

  // REG#697の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0697 <= imem05_in[15:12];
    49: reg_0697 <= imem03_in[3:0];
    54: reg_0697 <= imem05_in[15:12];
    endcase
  end

  // REG#698の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0698 <= imem04_in[11:8];
    49: reg_0698 <= imem03_in[11:8];
    54: reg_0698 <= imem04_in[11:8];
    68: reg_0698 <= imem04_in[11:8];
    endcase
  end

  // REG#699の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0699 <= imem04_in[7:4];
    49: reg_0699 <= imem03_in[15:12];
    54: reg_0699 <= imem02_in[7:4];
    72: reg_0699 <= imem03_in[15:12];
    117: reg_0699 <= imem04_in[7:4];
    120: reg_0699 <= imem04_in[7:4];
    endcase
  end

  // REG#700の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0700 <= imem05_in[3:0];
    57: reg_0700 <= imem05_in[3:0];
    endcase
  end

  // REG#701の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0701 <= imem05_in[11:8];
    58: reg_0701 <= imem00_in[7:4];
    76: reg_0701 <= imem00_in[7:4];
    80: reg_0701 <= imem00_in[7:4];
    82: reg_0701 <= imem05_in[11:8];
    endcase
  end

  // REG#702の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0702 <= imem05_in[7:4];
    59: reg_0702 <= imem05_in[7:4];
    87: reg_0702 <= imem05_in[7:4];
    endcase
  end

  // REG#703の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0703 <= imem07_in[3:0];
    60: reg_0703 <= imem07_in[3:0];
    endcase
  end

  // REG#704の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0704 <= imem07_in[11:8];
    65: reg_0704 <= imem03_in[3:0];
    80: reg_0704 <= op2_03_out;
    109: reg_0704 <= imem07_in[11:8];
    110: reg_0704 <= op2_03_out;
    endcase
  end

  // REG#705の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0705 <= imem02_in[11:8];
    71: reg_0705 <= op1_09_out;
    89: reg_0705 <= op1_09_out;
    93: reg_0705 <= op1_09_out;
    99: reg_0705 <= op1_09_out;
    101: reg_0705 <= op1_09_out;
    103: reg_0705 <= op1_09_out;
    105: reg_0705 <= op1_09_out;
    107: reg_0705 <= op1_09_out;
    109: reg_0705 <= op1_09_out;
    111: reg_0705 <= op1_09_out;
    117: reg_0705 <= imem02_in[11:8];
    120: reg_0705 <= op1_09_out;
    123: reg_0705 <= imem02_in[11:8];
    endcase
  end

  // REG#706の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0706 <= imem03_in[11:8];
    77: reg_0706 <= imem07_in[7:4];
    80: reg_0706 <= imem07_in[7:4];
    82: reg_0706 <= imem03_in[11:8];
    endcase
  end

  // REG#707の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0707 <= imem03_in[3:0];
    78: reg_0707 <= imem03_in[3:0];
    90: reg_0707 <= imem03_in[3:0];
    124: reg_0707 <= imem03_in[3:0];
    endcase
  end

  // REG#708の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0708 <= imem02_in[7:4];
    79: reg_0708 <= imem05_in[3:0];
    87: reg_0708 <= op2_06_out;
    97: reg_0708 <= imem05_in[3:0];
    100: reg_0708 <= imem05_in[3:0];
    106: reg_0708 <= imem05_in[3:0];
    108: reg_0708 <= imem05_in[3:0];
    110: reg_0708 <= imem05_in[3:0];
    117: reg_0708 <= imem05_in[3:0];
    endcase
  end

  // REG#709の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0709 <= imem03_in[7:4];
    82: reg_0709 <= imem03_in[7:4];
    endcase
  end

  // REG#710の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0710 <= imem03_in[15:12];
    84: reg_0710 <= imem03_in[15:12];
    100: reg_0710 <= op2_03_out;
    107: reg_0710 <= imem03_in[15:12];
    112: reg_0710 <= op2_03_out;
    endcase
  end

  // REG#711の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0711 <= imem02_in[15:12];
    84: reg_0711 <= imem02_in[15:12];
    endcase
  end

  // REG#712の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0712 <= imem02_in[3:0];
    88: reg_0712 <= imem02_in[3:0];
    90: reg_0712 <= imem02_in[3:0];
    endcase
  end

  // REG#713の入力
  always @ ( posedge clock ) begin
    case ( state )
    35: reg_0713 <= op1_01_out;
    90: reg_0713 <= op2_04_out;
    endcase
  end

  // REG#714の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0714 <= imem06_in[15:12];
    129: reg_0714 <= imem06_in[15:12];
    endcase
  end

  // REG#715の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0715 <= imem01_in[7:4];
    endcase
  end

  // REG#716の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0716 <= imem06_in[3:0];
    endcase
  end

  // REG#717の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0717 <= imem06_in[11:8];
    endcase
  end

  // REG#718の入力
  always @ ( posedge clock ) begin
    case ( state )
    36: reg_0718 <= imem06_in[7:4];
    endcase
  end

  // REG#719の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0719 <= imem04_in[11:8];
    40: reg_0719 <= imem04_in[11:8];
    endcase
  end

  // REG#720の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0720 <= imem06_in[7:4];
    41: reg_0720 <= imem06_in[7:4];
    endcase
  end

  // REG#721の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0721 <= imem04_in[3:0];
    43: reg_0721 <= imem04_in[3:0];
    69: reg_0721 <= op1_14_out;
    73: reg_0721 <= op1_14_out;
    75: reg_0721 <= op1_14_out;
    89: reg_0721 <= op1_14_out;
    91: reg_0721 <= op1_14_out;
    94: reg_0721 <= op1_14_out;
    100: reg_0721 <= imem04_in[3:0];
    103: reg_0721 <= imem02_in[7:4];
    127: reg_0721 <= imem04_in[3:0];
    endcase
  end

  // REG#722の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0722 <= imem00_in[7:4];
    44: reg_0722 <= imem00_in[7:4];
    endcase
  end

  // REG#723の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0723 <= imem00_in[15:12];
    43: reg_0723 <= imem00_in[15:12];
    endcase
  end

  // REG#724の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0724 <= imem01_in[3:0];
    43: reg_0724 <= imem01_in[3:0];
    67: reg_0724 <= imem01_in[3:0];
    85: reg_0724 <= imem01_in[3:0];
    endcase
  end

  // REG#725の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0725 <= imem00_in[3:0];
    45: reg_0725 <= imem00_in[3:0];
    64: reg_0725 <= op1_00_out;
    85: reg_0725 <= op1_00_out;
    87: reg_0725 <= op1_00_out;
    90: reg_0725 <= imem00_in[3:0];
    95: reg_0725 <= imem00_in[3:0];
    102: reg_0725 <= imem00_in[3:0];
    125: reg_0725 <= imem00_in[3:0];
    endcase
  end

  // REG#726の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0726 <= imem01_in[11:8];
    45: reg_0726 <= imem01_in[11:8];
    67: reg_0726 <= op1_00_out;
    70: reg_0726 <= imem01_in[11:8];
    endcase
  end

  // REG#727の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0727 <= imem01_in[15:12];
    45: reg_0727 <= imem01_in[15:12];
    67: reg_0727 <= imem01_in[15:12];
    88: reg_0727 <= imem01_in[15:12];
    endcase
  end

  // REG#728の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0728 <= imem01_in[7:4];
    45: reg_0728 <= imem01_in[7:4];
    64: reg_0728 <= imem01_in[7:4];
    76: reg_0728 <= imem01_in[7:4];
    78: reg_0728 <= op1_13_out;
    91: reg_0728 <= imem01_in[7:4];
    94: reg_0728 <= op1_13_out;
    97: reg_0728 <= imem01_in[7:4];
    endcase
  end

  // REG#729の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0729 <= imem06_in[11:8];
    45: reg_0729 <= imem06_in[11:8];
    64: reg_0729 <= op1_01_out;
    85: reg_0729 <= op1_01_out;
    94: reg_0729 <= imem06_in[11:8];
    97: reg_0729 <= imem06_in[11:8];
    116: reg_0729 <= imem06_in[11:8];
    120: reg_0729 <= imem06_in[11:8];
    endcase
  end

  // REG#730の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0730 <= imem06_in[3:0];
    46: reg_0730 <= imem06_in[3:0];
    68: reg_0730 <= imem06_in[3:0];
    endcase
  end

  // REG#731の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0731 <= imem04_in[7:4];
    47: reg_0731 <= op1_04_out;
    92: reg_0731 <= imem04_in[7:4];
    111: reg_0731 <= imem04_in[7:4];
    endcase
  end

  // REG#732の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0732 <= imem03_in[3:0];
    67: reg_0732 <= imem03_in[11:8];
    71: reg_0732 <= op1_12_out;
    89: reg_0732 <= op1_12_out;
    92: reg_0732 <= imem03_in[11:8];
    94: reg_0732 <= imem03_in[11:8];
    96: reg_0732 <= imem03_in[3:0];
    102: reg_0732 <= imem03_in[3:0];
    endcase
  end

  // REG#733の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0733 <= imem05_in[11:8];
    68: reg_0733 <= imem05_in[11:8];
    85: reg_0733 <= imem05_in[11:8];
    endcase
  end

  // REG#734の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0734 <= imem03_in[11:8];
    68: reg_0734 <= imem03_in[11:8];
    84: reg_0734 <= imem01_in[11:8];
    94: reg_0734 <= imem01_in[11:8];
    99: reg_0734 <= imem01_in[11:8];
    103: reg_0734 <= imem03_in[11:8];
    105: reg_0734 <= imem03_in[11:8];
    108: reg_0734 <= imem01_in[11:8];
    110: reg_0734 <= imem03_in[11:8];
    113: reg_0734 <= imem01_in[11:8];
    120: reg_0734 <= imem03_in[11:8];
    endcase
  end

  // REG#735の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0735 <= imem05_in[15:12];
    70: reg_0735 <= imem05_in[15:12];
    95: reg_0735 <= imem05_in[15:12];
    105: reg_0735 <= imem05_in[15:12];
    112: reg_0735 <= imem05_in[15:12];
    114: reg_0735 <= imem05_in[15:12];
    endcase
  end

  // REG#736の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0736 <= imem05_in[3:0];
    70: reg_0736 <= imem05_in[3:0];
    93: reg_0736 <= imem05_in[3:0];
    102: reg_0736 <= imem05_in[3:0];
    endcase
  end

  // REG#737の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0737 <= imem05_in[7:4];
    70: reg_0737 <= imem05_in[7:4];
    94: reg_0737 <= op2_03_out;
    endcase
  end

  // REG#738の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0738 <= imem07_in[15:12];
    123: reg_0738 <= imem07_in[15:12];
    endcase
  end

  // REG#739の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0739 <= imem07_in[3:0];
    endcase
  end

  // REG#740の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0740 <= imem07_in[11:8];
    endcase
  end

  // REG#741の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0741 <= imem07_in[7:4];
    endcase
  end

  // REG#742の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0742 <= imem01_in[15:12];
    54: reg_0742 <= imem02_in[11:8];
    72: reg_0742 <= imem01_in[15:12];
    endcase
  end

  // REG#743の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0743 <= imem01_in[11:8];
    54: reg_0743 <= imem01_in[7:4];
    73: reg_0743 <= imem01_in[7:4];
    endcase
  end

  // REG#744の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0744 <= imem04_in[11:8];
    54: reg_0744 <= imem02_in[15:12];
    74: reg_0744 <= imem02_in[15:12];
    88: reg_0744 <= imem04_in[11:8];
    90: reg_0744 <= imem02_in[15:12];
    endcase
  end

  // REG#745の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0745 <= imem05_in[3:0];
    55: reg_0745 <= imem05_in[3:0];
    74: reg_0745 <= op1_15_out;
    77: reg_0745 <= op1_15_out;
    79: reg_0745 <= op1_15_out;
    82: reg_0745 <= op1_15_out;
    85: reg_0745 <= imem02_in[3:0];
    endcase
  end

  // REG#746の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0746 <= imem01_in[3:0];
    55: reg_0746 <= imem01_in[3:0];
    endcase
  end

  // REG#747の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0747 <= imem01_in[7:4];
    55: reg_0747 <= imem01_in[7:4];
    endcase
  end

  // REG#748の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0748 <= imem05_in[11:8];
    58: reg_0748 <= imem00_in[3:0];
    76: reg_0748 <= imem00_in[3:0];
    79: reg_0748 <= imem05_in[11:8];
    89: reg_0748 <= imem05_in[11:8];
    91: reg_0748 <= imem00_in[3:0];
    93: reg_0748 <= imem00_in[3:0];
    97: reg_0748 <= imem00_in[3:0];
    100: reg_0748 <= imem00_in[3:0];
    endcase
  end

  // REG#749の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0749 <= imem05_in[7:4];
    60: reg_0749 <= op1_04_out;
    73: reg_0749 <= op1_04_out;
    88: reg_0749 <= op1_04_out;
    90: reg_0749 <= op2_05_out;
    endcase
  end

  // REG#750の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0750 <= imem05_in[15:12];
    61: reg_0750 <= imem05_in[15:12];
    93: reg_0750 <= imem05_in[15:12];
    101: reg_0750 <= imem05_in[15:12];
    105: reg_0750 <= imem03_in[15:12];
    110: reg_0750 <= imem03_in[15:12];
    114: reg_0750 <= imem03_in[15:12];
    117: reg_0750 <= imem03_in[15:12];
    123: reg_0750 <= imem03_in[15:12];
    endcase
  end

  // REG#751の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0751 <= imem06_in[15:12];
    61: reg_0751 <= imem06_in[15:12];
    67: reg_0751 <= imem06_in[15:12];
    79: reg_0751 <= imem06_in[15:12];
    85: reg_0751 <= imem06_in[15:12];
    endcase
  end

  // REG#752の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0752 <= imem06_in[11:8];
    62: reg_0752 <= imem06_in[11:8];
    endcase
  end

  // REG#753の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0753 <= imem06_in[7:4];
    64: reg_0753 <= op1_02_out;
    86: reg_0753 <= imem06_in[7:4];
    92: reg_0753 <= imem06_in[7:4];
    104: reg_0753 <= op2_00_out;
    117: reg_0753 <= op2_00_out;
    122: reg_0753 <= imem06_in[7:4];
    129: reg_0753 <= op2_00_out;
    endcase
  end

  // REG#754の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0754 <= imem06_in[3:0];
    67: reg_0754 <= imem06_in[3:0];
    78: reg_0754 <= imem01_in[7:4];
    96: reg_0754 <= imem06_in[3:0];
    98: reg_0754 <= imem06_in[3:0];
    endcase
  end

  // REG#755の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0755 <= imem03_in[15:12];
    71: reg_0755 <= imem06_in[7:4];
    79: reg_0755 <= op2_02_out;
    89: reg_0755 <= imem06_in[7:4];
    108: reg_0755 <= op2_02_out;
    endcase
  end

  // REG#756の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0756 <= imem03_in[11:8];
    71: reg_0756 <= op1_14_out;
    89: reg_0756 <= op2_05_out;
    100: reg_0756 <= op1_14_out;
    103: reg_0756 <= op1_14_out;
    108: reg_0756 <= op1_14_out;
    111: reg_0756 <= imem03_in[11:8];
    endcase
  end

  // REG#757の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0757 <= imem03_in[7:4];
    71: reg_0757 <= op1_06_out;
    90: reg_0757 <= op2_06_out;
    endcase
  end

  // REG#758の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0758 <= imem03_in[3:0];
    71: reg_0758 <= op1_15_out;
    92: reg_0758 <= imem03_in[3:0];
    95: reg_0758 <= op1_15_out;
    98: reg_0758 <= op1_15_out;
    101: reg_0758 <= op1_15_out;
    105: reg_0758 <= op1_15_out;
    108: reg_0758 <= op1_15_out;
    111: reg_0758 <= op1_15_out;
    114: reg_0758 <= op1_15_out;
    118: reg_0758 <= op1_15_out;
    122: reg_0758 <= imem03_in[3:0];
    125: reg_0758 <= imem03_in[3:0];
    endcase
  end

  // REG#759の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0759 <= op1_03_out;
    84: reg_0759 <= imem03_in[7:4];
    100: reg_0759 <= imem03_in[7:4];
    109: reg_0759 <= imem03_in[7:4];
    125: reg_0759 <= imem03_in[7:4];
    endcase
  end

  // REG#760の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0760 <= op1_04_out;
    82: reg_0760 <= op1_04_out;
    96: reg_0760 <= op1_04_out;
    98: reg_0760 <= op1_04_out;
    100: reg_0760 <= op1_04_out;
    102: reg_0760 <= op1_04_out;
    104: reg_0760 <= op1_04_out;
    106: reg_0760 <= op1_04_out;
    108: reg_0760 <= op1_04_out;
    112: reg_0760 <= op1_04_out;
    endcase
  end

  // REG#761の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0761 <= op1_01_out;
    89: reg_0761 <= op2_06_out;
    104: reg_0761 <= op1_01_out;
    106: reg_0761 <= op1_01_out;
    108: reg_0761 <= op1_01_out;
    110: reg_0761 <= op1_01_out;
    112: reg_0761 <= op1_01_out;
    endcase
  end

  // REG#762の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0762 <= op1_02_out;
    89: reg_0762 <= op1_02_out;
    endcase
  end

  // REG#763の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0763 <= op1_05_out;
    104: reg_0763 <= op1_05_out;
    114: reg_0763 <= op1_05_out;
    endcase
  end

  // REG#764の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0764 <= op1_06_out;
    91: reg_0764 <= op1_06_out;
    95: reg_0764 <= op1_06_out;
    97: reg_0764 <= op1_06_out;
    105: reg_0764 <= op1_06_out;
    endcase
  end

  // REG#765の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0765 <= op1_07_out;
    endcase
  end

  // REG#766の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0766 <= op1_08_out;
    92: reg_0766 <= op1_08_out;
    94: reg_0766 <= op1_08_out;
    96: reg_0766 <= op1_08_out;
    98: reg_0766 <= op1_08_out;
    100: reg_0766 <= op1_08_out;
    102: reg_0766 <= op1_08_out;
    104: reg_0766 <= op1_08_out;
    106: reg_0766 <= op1_08_out;
    108: reg_0766 <= op1_08_out;
    110: reg_0766 <= op1_08_out;
    endcase
  end

  // REG#767の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0767 <= op1_09_out;
    endcase
  end

  // REG#768の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0768 <= op1_10_out;
    95: reg_0768 <= op1_10_out;
    101: reg_0768 <= op1_10_out;
    105: reg_0768 <= op1_10_out;
    endcase
  end

  // REG#769の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0769 <= op1_11_out;
    endcase
  end

  // REG#770の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0770 <= op1_12_out;
    105: reg_0770 <= op1_12_out;
    107: reg_0770 <= op1_12_out;
    109: reg_0770 <= op1_12_out;
    111: reg_0770 <= op1_12_out;
    114: reg_0770 <= op1_12_out;
    116: reg_0770 <= op1_12_out;
    118: reg_0770 <= op1_12_out;
    126: reg_0770 <= op1_12_out;
    endcase
  end

  // REG#771の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0771 <= op1_13_out;
    109: reg_0771 <= op1_13_out;
    116: reg_0771 <= op1_13_out;
    119: reg_0771 <= op1_13_out;
    128: reg_0771 <= op1_13_out;
    endcase
  end

  // REG#772の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0772 <= op1_14_out;
    112: reg_0772 <= op1_14_out;
    116: reg_0772 <= op1_14_out;
    119: reg_0772 <= op1_14_out;
    121: reg_0772 <= op1_14_out;
    124: reg_0772 <= op1_14_out;
    128: reg_0772 <= op1_14_out;
    endcase
  end

  // REG#773の入力
  always @ ( posedge clock ) begin
    case ( state )
    37: reg_0773 <= op1_15_out;
    121: reg_0773 <= op1_15_out;
    124: reg_0773 <= op1_15_out;
    endcase
  end

  // REG#774の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0774 <= imem07_in[15:12];
    endcase
  end

  // REG#775の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0775 <= imem07_in[11:8];
    endcase
  end

  // REG#776の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0776 <= imem02_in[7:4];
    endcase
  end

  // REG#777の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0777 <= imem07_in[3:0];
    endcase
  end

  // REG#778の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0778 <= imem02_in[15:12];
    endcase
  end

  // REG#779の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0779 <= imem07_in[7:4];
    endcase
  end

  // REG#780の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0780 <= imem06_in[11:8];
    48: reg_0780 <= imem06_in[11:8];
    52: reg_0780 <= imem06_in[11:8];
    66: reg_0780 <= imem06_in[11:8];
    80: reg_0780 <= imem06_in[11:8];
    101: reg_0780 <= imem06_in[11:8];
    endcase
  end

  // REG#781の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0781 <= op1_00_out;
    47: reg_0781 <= op1_06_out;
    endcase
  end

  // REG#782の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0782 <= imem06_in[3:0];
    50: reg_0782 <= imem06_in[3:0];
    64: reg_0782 <= op1_06_out;
    86: reg_0782 <= op1_06_out;
    88: reg_0782 <= op1_06_out;
    95: reg_0782 <= imem06_in[3:0];
    endcase
  end

  // REG#783の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0783 <= imem06_in[7:4];
    50: reg_0783 <= imem06_in[7:4];
    67: reg_0783 <= op1_01_out;
    79: reg_0783 <= imem03_in[11:8];
    endcase
  end

  // REG#784の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0784 <= imem06_in[15:12];
    51: reg_0784 <= imem06_in[15:12];
    64: reg_0784 <= op1_07_out;
    85: reg_0784 <= op1_07_out;
    97: reg_0784 <= imem06_in[15:12];
    108: reg_0784 <= imem06_in[15:12];
    112: reg_0784 <= imem06_in[15:12];
    115: reg_0784 <= imem06_in[15:12];
    119: reg_0784 <= imem06_in[15:12];
    122: reg_0784 <= imem06_in[15:12];
    endcase
  end

  // REG#785の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0785 <= imem01_in[11:8];
    52: reg_0785 <= imem01_in[11:8];
    61: reg_0785 <= imem01_in[11:8];
    78: reg_0785 <= imem01_in[11:8];
    102: reg_0785 <= imem01_in[11:8];
    106: reg_0785 <= imem01_in[11:8];
    115: reg_0785 <= imem01_in[11:8];
    122: reg_0785 <= imem01_in[11:8];
    endcase
  end

  // REG#786の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0786 <= imem01_in[3:0];
    52: reg_0786 <= imem01_in[3:0];
    61: reg_0786 <= imem01_in[3:0];
    76: reg_0786 <= imem07_in[3:0];
    83: reg_0786 <= imem07_in[3:0];
    87: reg_0786 <= imem07_in[3:0];
    endcase
  end

  // REG#787の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0787 <= imem01_in[15:12];
    55: reg_0787 <= imem01_in[15:12];
    endcase
  end

  // REG#788の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0788 <= imem01_in[7:4];
    56: reg_0788 <= imem01_in[7:4];
    60: reg_0788 <= imem01_in[7:4];
    87: reg_0788 <= op2_07_out;
    99: reg_0788 <= imem01_in[7:4];
    101: reg_0788 <= imem01_in[7:4];
    109: reg_0788 <= imem01_in[7:4];
    119: reg_0788 <= imem01_in[7:4];
    endcase
  end

  // REG#789の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0789 <= imem03_in[15:12];
    58: reg_0789 <= imem03_in[15:12];
    endcase
  end

  // REG#790の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0790 <= imem03_in[7:4];
    59: reg_0790 <= imem03_in[7:4];
    endcase
  end

  // REG#791の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0791 <= imem07_in[11:8];
    60: reg_0791 <= imem00_in[3:0];
    75: reg_0791 <= imem00_in[3:0];
    94: reg_0791 <= imem07_in[11:8];
    96: reg_0791 <= imem07_in[11:8];
    99: reg_0791 <= imem07_in[11:8];
    103: reg_0791 <= imem00_in[3:0];
    108: reg_0791 <= imem07_in[11:8];
    111: reg_0791 <= imem00_in[3:0];
    118: reg_0791 <= imem00_in[3:0];
    120: reg_0791 <= imem07_in[11:8];
    endcase
  end

  // REG#792の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0792 <= imem05_in[3:0];
    69: reg_0792 <= op1_06_out;
    74: reg_0792 <= op1_06_out;
    89: reg_0792 <= imem05_in[3:0];
    94: reg_0792 <= imem05_in[3:0];
    98: reg_0792 <= imem05_in[3:0];
    103: reg_0792 <= imem05_in[3:0];
    endcase
  end

  // REG#793の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0793 <= imem05_in[15:12];
    69: reg_0793 <= op1_07_out;
    74: reg_0793 <= op1_07_out;
    76: reg_0793 <= op1_07_out;
    78: reg_0793 <= op1_07_out;
    96: reg_0793 <= imem05_in[15:12];
    122: reg_0793 <= imem05_in[15:12];
    endcase
  end

  // REG#794の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0794 <= imem05_in[7:4];
    69: reg_0794 <= op1_05_out;
    76: reg_0794 <= imem05_in[7:4];
    102: reg_0794 <= imem05_in[7:4];
    endcase
  end

  // REG#795の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0795 <= imem04_in[15:12];
    70: reg_0795 <= imem06_in[3:0];
    77: reg_0795 <= imem06_in[3:0];
    115: reg_0795 <= imem06_in[3:0];
    122: reg_0795 <= imem06_in[3:0];
    128: reg_0795 <= imem04_in[15:12];
    endcase
  end

  // REG#796の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0796 <= imem04_in[3:0];
    71: reg_0796 <= imem04_in[3:0];
    82: reg_0796 <= imem04_in[3:0];
    endcase
  end

  // REG#797の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0797 <= imem04_in[11:8];
    72: reg_0797 <= imem05_in[15:12];
    92: reg_0797 <= imem04_in[11:8];
    111: reg_0797 <= imem04_in[11:8];
    endcase
  end

  // REG#798の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0798 <= imem04_in[7:4];
    72: reg_0798 <= imem01_in[7:4];
    endcase
  end

  // REG#799の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0799 <= imem05_in[11:8];
    72: reg_0799 <= imem05_in[11:8];
    91: reg_0799 <= imem05_in[11:8];
    endcase
  end

  // REG#800の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0800 <= imem02_in[11:8];
    80: reg_0800 <= imem02_in[11:8];
    endcase
  end

  // REG#801の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0801 <= imem02_in[3:0];
    80: reg_0801 <= imem02_in[3:0];
    endcase
  end

  // REG#802の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0802 <= imem02_in[7:4];
    84: reg_0802 <= imem02_in[7:4];
    endcase
  end

  // REG#803の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0803 <= imem00_in[15:12];
    88: reg_0803 <= imem00_in[15:12];
    endcase
  end

  // REG#804の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0804 <= imem00_in[7:4];
    88: reg_0804 <= imem00_in[7:4];
    endcase
  end

  // REG#805の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0805 <= imem00_in[11:8];
    87: reg_0805 <= imem00_in[11:8];
    endcase
  end

  // REG#806の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0806 <= imem00_in[3:0];
    88: reg_0806 <= imem00_in[3:0];
    endcase
  end

  // REG#807の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0807 <= op1_01_out;
    endcase
  end

  // REG#808の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0808 <= op1_02_out;
    endcase
  end

  // REG#809の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0809 <= op1_03_out;
    endcase
  end

  // REG#810の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0810 <= op1_04_out;
    endcase
  end

  // REG#811の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0811 <= op1_05_out;
    endcase
  end

  // REG#812の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0812 <= op1_06_out;
    endcase
  end

  // REG#813の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0813 <= op1_07_out;
    endcase
  end

  // REG#814の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0814 <= op1_08_out;
    endcase
  end

  // REG#815の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0815 <= op1_09_out;
    endcase
  end

  // REG#816の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0816 <= op1_10_out;
    endcase
  end

  // REG#817の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0817 <= op1_11_out;
    endcase
  end

  // REG#818の入力
  always @ ( posedge clock ) begin
    case ( state )
    38: reg_0818 <= op1_12_out;
    endcase
  end

  // REG#819の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0819 <= imem01_in[15:12];
    46: reg_0819 <= imem01_in[15:12];
    endcase
  end

  // REG#820の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0820 <= imem00_in[3:0];
    52: reg_0820 <= imem02_in[3:0];
    65: reg_0820 <= imem02_in[3:0];
    72: reg_0820 <= imem01_in[11:8];
    endcase
  end

  // REG#821の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0821 <= imem00_in[11:8];
    52: reg_0821 <= imem07_in[15:12];
    67: reg_0821 <= imem00_in[11:8];
    endcase
  end

  // REG#822の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0822 <= imem06_in[11:8];
    57: reg_0822 <= imem02_in[7:4];
    61: reg_0822 <= imem01_in[7:4];
    77: reg_0822 <= imem02_in[7:4];
    129: reg_0822 <= imem06_in[11:8];
    endcase
  end

  // REG#823の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0823 <= imem03_in[15:12];
    57: reg_0823 <= op1_01_out;
    79: reg_0823 <= imem03_in[15:12];
    endcase
  end

  // REG#824の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0824 <= imem00_in[15:12];
    58: reg_0824 <= imem00_in[15:12];
    74: reg_0824 <= imem00_in[15:12];
    76: reg_0824 <= imem02_in[15:12];
    88: reg_0824 <= imem02_in[15:12];
    94: reg_0824 <= imem00_in[15:12];
    97: reg_0824 <= imem00_in[15:12];
    105: reg_0824 <= imem02_in[15:12];
    107: reg_0824 <= imem02_in[15:12];
    endcase
  end

  // REG#825の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0825 <= imem06_in[7:4];
    58: reg_0825 <= op1_05_out;
    80: reg_0825 <= op1_05_out;
    83: reg_0825 <= imem06_in[7:4];
    87: reg_0825 <= op1_05_out;
    90: reg_0825 <= imem06_in[7:4];
    108: reg_0825 <= imem06_in[7:4];
    110: reg_0825 <= imem06_in[7:4];
    125: reg_0825 <= imem06_in[7:4];
    endcase
  end

  // REG#826の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0826 <= imem06_in[3:0];
    58: reg_0826 <= op1_06_out;
    80: reg_0826 <= op1_06_out;
    82: reg_0826 <= op1_06_out;
    84: reg_0826 <= op1_06_out;
    87: reg_0826 <= op1_06_out;
    89: reg_0826 <= op1_06_out;
    97: reg_0826 <= imem06_in[3:0];
    116: reg_0826 <= imem06_in[3:0];
    123: reg_0826 <= imem06_in[3:0];
    endcase
  end

  // REG#827の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0827 <= imem06_in[15:12];
    62: reg_0827 <= imem06_in[15:12];
    endcase
  end

  // REG#828の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0828 <= imem05_in[3:0];
    62: reg_0828 <= imem05_in[3:0];
    endcase
  end

  // REG#829の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0829 <= imem02_in[15:12];
    64: reg_0829 <= op1_08_out;
    86: reg_0829 <= imem02_in[15:12];
    endcase
  end

  // REG#830の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0830 <= imem02_in[11:8];
    66: reg_0830 <= imem03_in[3:0];
    72: reg_0830 <= imem01_in[3:0];
    endcase
  end

  // REG#831の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0831 <= imem05_in[11:8];
    68: reg_0831 <= imem03_in[3:0];
    84: reg_0831 <= imem05_in[3:0];
    123: reg_0831 <= imem03_in[3:0];
    endcase
  end

  // REG#832の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0832 <= imem05_in[15:12];
    69: reg_0832 <= imem05_in[15:12];
    117: reg_0832 <= imem05_in[15:12];
    endcase
  end

  // REG#833の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0833 <= imem05_in[7:4];
    69: reg_0833 <= imem05_in[7:4];
    114: reg_0833 <= imem05_in[7:4];
    endcase
  end

  // REG#834の入力
  always @ ( posedge clock ) begin
    case ( state )
    39: reg_0834 <= op1_01_out;
    86: reg_0834 <= op1_01_out;
    88: reg_0834 <= op2_12_out;
    98: reg_0834 <= op1_01_out;
    endcase
  end

  // REG#835の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0835 <= imem04_in[15:12];
    endcase
  end

  // REG#836の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0836 <= imem04_in[7:4];
    endcase
  end

  // REG#837の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0837 <= imem04_in[3:0];
    endcase
  end

  // REG#838の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0838 <= op1_03_out;
    66: reg_0838 <= op1_03_out;
    endcase
  end

  // REG#839の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0839 <= imem02_in[7:4];
    72: reg_0839 <= op1_06_out;
    76: reg_0839 <= imem02_in[7:4];
    90: reg_0839 <= imem02_in[7:4];
    endcase
  end

  // REG#840の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0840 <= imem03_in[7:4];
    73: reg_0840 <= imem03_in[7:4];
    104: reg_0840 <= imem03_in[7:4];
    114: reg_0840 <= imem03_in[7:4];
    116: reg_0840 <= imem03_in[7:4];
    endcase
  end

  // REG#841の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0841 <= imem00_in[7:4];
    74: reg_0841 <= imem00_in[7:4];
    78: reg_0841 <= imem00_in[7:4];
    125: reg_0841 <= imem00_in[7:4];
    endcase
  end

  // REG#842の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0842 <= imem00_in[11:8];
    74: reg_0842 <= imem00_in[11:8];
    75: reg_0842 <= op2_01_out;
    86: reg_0842 <= op2_01_out;
    106: reg_0842 <= op2_01_out;
    125: reg_0842 <= op2_01_out;
    endcase
  end

  // REG#843の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0843 <= imem00_in[15:12];
    73: reg_0843 <= op1_15_out;
    75: reg_0843 <= op1_15_out;
    89: reg_0843 <= op1_15_out;
    92: reg_0843 <= imem00_in[15:12];
    93: reg_0843 <= op1_15_out;
    96: reg_0843 <= op1_15_out;
    99: reg_0843 <= op1_15_out;
    102: reg_0843 <= imem00_in[15:12];
    122: reg_0843 <= imem00_in[15:12];
    endcase
  end

  // REG#844の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0844 <= imem00_in[3:0];
    73: reg_0844 <= op2_00_out;
    75: reg_0844 <= op2_00_out;
    85: reg_0844 <= op2_00_out;
    90: reg_0844 <= op2_00_out;
    125: reg_0844 <= op2_00_out;
    endcase
  end

  // REG#845の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0845 <= imem02_in[11:8];
    78: reg_0845 <= imem02_in[11:8];
    endcase
  end

  // REG#846の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0846 <= imem02_in[15:12];
    78: reg_0846 <= imem02_in[15:12];
    endcase
  end

  // REG#847の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0847 <= op1_00_out;
    79: reg_0847 <= imem03_in[3:0];
    endcase
  end

  // REG#848の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0848 <= imem02_in[3:0];
    81: reg_0848 <= imem02_in[3:0];
    endcase
  end

  // REG#849の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0849 <= imem03_in[11:8];
    83: reg_0849 <= op2_01_out;
    endcase
  end

  // REG#850の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0850 <= op1_02_out;
    83: reg_0850 <= op1_02_out;
    endcase
  end

  // REG#851の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0851 <= imem07_in[11:8];
    86: reg_0851 <= imem07_in[11:8];
    endcase
  end

  // REG#852の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0852 <= op1_05_out;
    87: reg_0852 <= op2_08_out;
    endcase
  end

  // REG#853の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0853 <= op1_01_out;
    89: reg_0853 <= op2_07_out;
    endcase
  end

  // REG#854の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0854 <= op1_04_out;
    endcase
  end

  // REG#855の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0855 <= op1_06_out;
    endcase
  end

  // REG#856の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0856 <= op1_07_out;
    endcase
  end

  // REG#857の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0857 <= op1_08_out;
    endcase
  end

  // REG#858の入力
  always @ ( posedge clock ) begin
    case ( state )
    40: reg_0858 <= op1_09_out;
    endcase
  end

  // REG#859の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0859 <= imem06_in[15:12];
    126: reg_0859 <= imem06_in[15:12];
    endcase
  end

  // REG#860の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0860 <= imem06_in[3:0];
    endcase
  end

  // REG#861の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0861 <= imem05_in[15:12];
    endcase
  end

  // REG#862の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0862 <= imem04_in[15:12];
    endcase
  end

  // REG#863の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0863 <= imem06_in[11:8];
    endcase
  end

  // REG#864の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0864 <= imem05_in[3:0];
    endcase
  end

  // REG#865の入力
  always @ ( posedge clock ) begin
    case ( state )
    41: reg_0865 <= op1_00_out;
    47: reg_0865 <= op1_07_out;
    endcase
  end

  // REG#866の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0866 <= imem06_in[11:8];
    60: reg_0866 <= imem00_in[11:8];
    75: reg_0866 <= imem00_in[11:8];
    95: reg_0866 <= imem00_in[11:8];
    98: reg_0866 <= imem00_in[11:8];
    104: reg_0866 <= imem00_in[11:8];
    112: reg_0866 <= imem00_in[11:8];
    115: reg_0866 <= imem00_in[11:8];
    endcase
  end

  // REG#867の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0867 <= imem07_in[3:0];
    59: reg_0867 <= op1_04_out;
    82: reg_0867 <= imem07_in[3:0];
    84: reg_0867 <= op1_04_out;
    93: reg_0867 <= imem07_in[3:0];
    99: reg_0867 <= imem07_in[3:0];
    101: reg_0867 <= imem07_in[3:0];
    103: reg_0867 <= imem07_in[3:0];
    114: reg_0867 <= imem07_in[3:0];
    116: reg_0867 <= imem07_in[3:0];
    123: reg_0867 <= imem07_in[3:0];
    endcase
  end

  // REG#868の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0868 <= imem01_in[7:4];
    62: reg_0868 <= imem01_in[7:4];
    73: reg_0868 <= imem07_in[3:0];
    77: reg_0868 <= imem00_in[3:0];
    88: reg_0868 <= imem07_in[3:0];
    96: reg_0868 <= imem01_in[7:4];
    121: reg_0868 <= imem01_in[7:4];
    endcase
  end

  // REG#869の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0869 <= imem06_in[3:0];
    62: reg_0869 <= imem06_in[3:0];
    endcase
  end

  // REG#870の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0870 <= imem06_in[7:4];
    64: reg_0870 <= imem06_in[7:4];
    76: reg_0870 <= imem06_in[7:4];
    endcase
  end

  // REG#871の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0871 <= imem01_in[3:0];
    64: reg_0871 <= op1_09_out;
    85: reg_0871 <= op1_09_out;
    87: reg_0871 <= op1_09_out;
    90: reg_0871 <= imem01_in[3:0];
    103: reg_0871 <= imem01_in[3:0];
    endcase
  end

  // REG#872の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0872 <= imem05_in[11:8];
    66: reg_0872 <= imem05_in[11:8];
    endcase
  end

  // REG#873の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0873 <= imem05_in[7:4];
    66: reg_0873 <= imem05_in[7:4];
    endcase
  end

  // REG#874の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0874 <= imem01_in[15:12];
    66: reg_0874 <= imem01_in[15:12];
    87: reg_0874 <= op2_09_out;
    100: reg_0874 <= imem01_in[15:12];
    103: reg_0874 <= imem01_in[15:12];
    128: reg_0874 <= imem01_in[15:12];
    endcase
  end

  // REG#875の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0875 <= imem01_in[11:8];
    67: reg_0875 <= imem01_in[11:8];
    88: reg_0875 <= imem01_in[11:8];
    endcase
  end

  // REG#876の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0876 <= imem02_in[3:0];
    68: reg_0876 <= imem02_in[3:0];
    endcase
  end

  // REG#877の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0877 <= imem02_in[15:12];
    68: reg_0877 <= imem05_in[7:4];
    87: reg_0877 <= op2_10_out;
    101: reg_0877 <= imem05_in[7:4];
    106: reg_0877 <= imem05_in[7:4];
    108: reg_0877 <= imem02_in[15:12];
    112: reg_0877 <= imem02_in[15:12];
    116: reg_0877 <= imem05_in[7:4];
    118: reg_0877 <= imem02_in[15:12];
    endcase
  end

  // REG#878の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0878 <= imem02_in[7:4];
    68: reg_0878 <= imem02_in[7:4];
    endcase
  end

  // REG#879の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0879 <= imem02_in[11:8];
    68: reg_0879 <= imem05_in[15:12];
    88: reg_0879 <= imem02_in[11:8];
    99: reg_0879 <= imem05_in[15:12];
    101: reg_0879 <= imem02_in[11:8];
    endcase
  end

  // REG#880の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0880 <= imem03_in[11:8];
    endcase
  end

  // REG#881の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0881 <= imem00_in[3:0];
    endcase
  end

  // REG#882の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0882 <= imem03_in[7:4];
    endcase
  end

  // REG#883の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0883 <= imem00_in[11:8];
    endcase
  end

  // REG#884の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0884 <= imem03_in[15:12];
    endcase
  end

  // REG#885の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0885 <= imem03_in[3:0];
    endcase
  end

  // REG#886の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0886 <= imem00_in[15:12];
    endcase
  end

  // REG#887の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0887 <= imem00_in[7:4];
    endcase
  end

  // REG#888の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0888 <= imem05_in[15:12];
    53: reg_0888 <= op1_10_out;
    74: reg_0888 <= op1_10_out;
    88: reg_0888 <= op1_10_out;
    90: reg_0888 <= op1_10_out;
    92: reg_0888 <= op1_10_out;
    100: reg_0888 <= imem05_in[15:12];
    102: reg_0888 <= imem05_in[15:12];
    endcase
  end

  // REG#889の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0889 <= imem03_in[15:12];
    57: reg_0889 <= imem02_in[3:0];
    62: reg_0889 <= imem02_in[3:0];
    73: reg_0889 <= imem03_in[15:12];
    103: reg_0889 <= imem02_in[3:0];
    endcase
  end

  // REG#890の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0890 <= imem05_in[7:4];
    57: reg_0890 <= op1_05_out;
    78: reg_0890 <= op1_05_out;
    90: reg_0890 <= op1_05_out;
    93: reg_0890 <= imem05_in[7:4];
    104: reg_0890 <= imem05_in[7:4];
    119: reg_0890 <= imem05_in[7:4];
    endcase
  end

  // REG#891の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0891 <= imem03_in[11:8];
    58: reg_0891 <= imem03_in[11:8];
    endcase
  end

  // REG#892の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0892 <= imem07_in[3:0];
    65: reg_0892 <= imem07_in[3:0];
    endcase
  end

  // REG#893の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0893 <= imem07_in[11:8];
    64: reg_0893 <= op1_10_out;
    86: reg_0893 <= op1_10_out;
    88: reg_0893 <= op2_13_out;
    97: reg_0893 <= imem07_in[11:8];
    100: reg_0893 <= imem07_in[11:8];
    103: reg_0893 <= imem07_in[11:8];
    115: reg_0893 <= imem07_in[11:8];
    endcase
  end

  // REG#894の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0894 <= imem07_in[7:4];
    65: reg_0894 <= imem07_in[7:4];
    endcase
  end

  // REG#895の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0895 <= imem05_in[11:8];
    66: reg_0895 <= imem01_in[7:4];
    83: reg_0895 <= imem01_in[7:4];
    endcase
  end

  // REG#896の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0896 <= imem05_in[3:0];
    66: reg_0896 <= imem01_in[11:8];
    85: reg_0896 <= imem01_in[11:8];
    endcase
  end

  // REG#897の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0897 <= imem02_in[3:0];
    67: reg_0897 <= imem02_in[11:8];
    85: reg_0897 <= imem02_in[11:8];
    endcase
  end

  // REG#898の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0898 <= imem02_in[7:4];
    67: reg_0898 <= imem04_in[11:8];
    87: reg_0898 <= op2_11_out;
    102: reg_0898 <= imem04_in[11:8];
    104: reg_0898 <= imem04_in[11:8];
    106: reg_0898 <= imem04_in[11:8];
    109: reg_0898 <= imem02_in[7:4];
    endcase
  end

  // REG#899の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0899 <= imem01_in[7:4];
    68: reg_0899 <= imem01_in[7:4];
    endcase
  end

  // REG#900の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0900 <= imem02_in[15:12];
    67: reg_0900 <= op1_02_out;
    100: reg_0900 <= imem02_in[15:12];
    109: reg_0900 <= imem02_in[15:12];
    endcase
  end

  // REG#901の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0901 <= imem01_in[15:12];
    68: reg_0901 <= imem01_in[15:12];
    endcase
  end

  // REG#902の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0902 <= imem01_in[11:8];
    67: reg_0902 <= op1_03_out;
    95: reg_0902 <= imem01_in[11:8];
    endcase
  end

  // REG#903の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0903 <= imem02_in[11:8];
    67: reg_0903 <= op1_04_out;
    105: reg_0903 <= imem02_in[11:8];
    107: reg_0903 <= imem02_in[11:8];
    endcase
  end

  // REG#904の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0904 <= imem04_in[11:8];
    69: reg_0904 <= op1_10_out;
    77: reg_0904 <= imem04_in[11:8];
    endcase
  end

  // REG#905の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0905 <= imem06_in[15:12];
    77: reg_0905 <= imem06_in[15:12];
    116: reg_0905 <= imem06_in[15:12];
    123: reg_0905 <= imem06_in[15:12];
    endcase
  end

  // REG#906の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0906 <= imem06_in[7:4];
    77: reg_0906 <= imem06_in[7:4];
    112: reg_0906 <= imem06_in[7:4];
    115: reg_0906 <= imem06_in[7:4];
    endcase
  end

  // REG#907の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0907 <= imem06_in[3:0];
    77: reg_0907 <= imem00_in[11:8];
    88: reg_0907 <= imem00_in[11:8];
    endcase
  end

  // REG#908の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0908 <= imem06_in[11:8];
    77: reg_0908 <= imem06_in[11:8];
    122: reg_0908 <= imem06_in[11:8];
    endcase
  end

  // REG#909の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0909 <= op1_03_out;
    85: reg_0909 <= op1_03_out;
    endcase
  end

  // REG#910の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0910 <= op1_00_out;
    89: reg_0910 <= op2_08_out;
    endcase
  end

  // REG#911の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0911 <= op1_01_out;
    endcase
  end

  // REG#912の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0912 <= op1_02_out;
    endcase
  end

  // REG#913の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0913 <= op1_04_out;
    endcase
  end

  // REG#914の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0914 <= op1_05_out;
    endcase
  end

  // REG#915の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0915 <= op1_06_out;
    endcase
  end

  // REG#916の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0916 <= op1_07_out;
    endcase
  end

  // REG#917の入力
  always @ ( posedge clock ) begin
    case ( state )
    43: reg_0917 <= imem00_in[11:8];
    endcase
  end

  // REG#918の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0918 <= op1_08_out;
    endcase
  end

  // REG#919の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0919 <= op1_09_out;
    endcase
  end

  // REG#920の入力
  always @ ( posedge clock ) begin
    case ( state )
    42: reg_0920 <= op1_10_out;
    endcase
  end

  // REG#921の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0921 <= imem07_in[3:0];
    49: reg_0921 <= imem07_in[3:0];
    endcase
  end

  // REG#922の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0922 <= imem07_in[15:12];
    49: reg_0922 <= imem02_in[7:4];
    61: reg_0922 <= imem07_in[15:12];
    endcase
  end

  // REG#923の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0923 <= imem07_in[11:8];
    49: reg_0923 <= imem07_in[11:8];
    endcase
  end

  // REG#924の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0924 <= imem07_in[7:4];
    49: reg_0924 <= imem07_in[7:4];
    endcase
  end

  // REG#925の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0925 <= imem06_in[3:0];
    64: reg_0925 <= imem06_in[3:0];
    76: reg_0925 <= imem06_in[3:0];
    endcase
  end

  // REG#926の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0926 <= imem00_in[15:12];
    64: reg_0926 <= op1_11_out;
    85: reg_0926 <= op1_11_out;
    87: reg_0926 <= op1_11_out;
    89: reg_0926 <= op1_11_out;
    92: reg_0926 <= op1_11_out;
    95: reg_0926 <= imem00_in[15:12];
    103: reg_0926 <= imem00_in[15:12];
    108: reg_0926 <= imem00_in[15:12];
    111: reg_0926 <= imem00_in[15:12];
    117: reg_0926 <= imem00_in[15:12];
    123: reg_0926 <= imem00_in[15:12];
    endcase
  end

  // REG#927の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0927 <= imem00_in[11:8];
    66: reg_0927 <= imem00_in[11:8];
    endcase
  end

  // REG#928の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0928 <= imem00_in[7:4];
    66: reg_0928 <= imem00_in[7:4];
    endcase
  end

  // REG#929の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0929 <= imem06_in[7:4];
    67: reg_0929 <= op1_05_out;
    109: reg_0929 <= imem06_in[7:4];
    114: reg_0929 <= imem06_in[7:4];
    endcase
  end

  // REG#930の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0930 <= imem01_in[3:0];
    69: reg_0930 <= imem01_in[3:0];
    endcase
  end

  // REG#931の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0931 <= imem06_in[15:12];
    68: reg_0931 <= op1_01_out;
    75: reg_0931 <= op1_01_out;
    89: reg_0931 <= imem06_in[15:12];
    109: reg_0931 <= imem06_in[15:12];
    113: reg_0931 <= imem06_in[15:12];
    117: reg_0931 <= imem06_in[15:12];
    125: reg_0931 <= imem06_in[15:12];
    endcase
  end

  // REG#932の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0932 <= imem04_in[15:12];
    69: reg_0932 <= op1_11_out;
    77: reg_0932 <= imem04_in[15:12];
    endcase
  end

  // REG#933の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0933 <= imem02_in[15:12];
    70: reg_0933 <= op1_03_out;
    79: reg_0933 <= op2_03_out;
    89: reg_0933 <= op2_09_out;
    114: reg_0933 <= imem02_in[15:12];
    116: reg_0933 <= imem02_in[15:12];
    121: reg_0933 <= op2_03_out;
    endcase
  end

  // REG#934の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0934 <= imem02_in[7:4];
    71: reg_0934 <= imem02_in[7:4];
    endcase
  end

  // REG#935の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0935 <= imem02_in[11:8];
    70: reg_0935 <= op1_05_out;
    79: reg_0935 <= op1_05_out;
    82: reg_0935 <= op1_05_out;
    122: reg_0935 <= imem02_in[11:8];
    endcase
  end

  // REG#936の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0936 <= imem04_in[7:4];
    70: reg_0936 <= op1_06_out;
    80: reg_0936 <= op2_04_out;
    110: reg_0936 <= imem04_in[7:4];
    115: reg_0936 <= imem04_in[7:4];
    127: reg_0936 <= imem04_in[7:4];
    endcase
  end

  // REG#937の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0937 <= imem05_in[7:4];
    75: reg_0937 <= imem05_in[7:4];
    endcase
  end

  // REG#938の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0938 <= imem05_in[15:12];
    77: reg_0938 <= imem05_in[15:12];
    endcase
  end

  // REG#939の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0939 <= imem05_in[11:8];
    77: reg_0939 <= imem05_in[11:8];
    endcase
  end

  // REG#940の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0940 <= imem05_in[3:0];
    77: reg_0940 <= imem05_in[3:0];
    endcase
  end

  // REG#941の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0941 <= op1_03_out;
    80: reg_0941 <= op2_05_out;
    endcase
  end

  // REG#942の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0942 <= op1_00_out;
    88: reg_0942 <= op2_14_out;
    endcase
  end

  // REG#943の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0943 <= op1_01_out;
    88: reg_0943 <= op2_15_out;
    endcase
  end

  // REG#944の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0944 <= op1_02_out;
    89: reg_0944 <= op2_10_out;
    endcase
  end

  // REG#945の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0945 <= op1_04_out;
    endcase
  end

  // REG#946の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0946 <= op1_05_out;
    endcase
  end

  // REG#947の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0947 <= op1_06_out;
    endcase
  end

  // REG#948の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0948 <= op1_07_out;
    endcase
  end

  // REG#949の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0949 <= op1_08_out;
    endcase
  end

  // REG#950の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0950 <= op1_09_out;
    endcase
  end

  // REG#951の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0951 <= op1_10_out;
    endcase
  end

  // REG#952の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0952 <= imem03_in[15:12];
    124: reg_0952 <= imem03_in[15:12];
    endcase
  end

  // REG#953の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0953 <= op1_11_out;
    endcase
  end

  // REG#954の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0954 <= imem03_in[3:0];
    endcase
  end

  // REG#955の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0955 <= op1_12_out;
    endcase
  end

  // REG#956の入力
  always @ ( posedge clock ) begin
    case ( state )
    44: reg_0956 <= op1_13_out;
    endcase
  end

  // REG#957の入力
  always @ ( posedge clock ) begin
    case ( state )
    45: reg_0957 <= imem03_in[11:8];
    endcase
  end

  // REG#958の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0958 <= imem00_in[15:12];
    67: reg_0958 <= op1_06_out;
    105: reg_0958 <= imem00_in[15:12];
    107: reg_0958 <= imem00_in[15:12];
    112: reg_0958 <= imem00_in[15:12];
    116: reg_0958 <= imem00_in[15:12];
    118: reg_0958 <= imem00_in[15:12];
    121: reg_0958 <= imem00_in[15:12];
    endcase
  end

  // REG#959の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0959 <= imem00_in[11:8];
    68: reg_0959 <= op1_02_out;
    75: reg_0959 <= op2_02_out;
    87: reg_0959 <= op2_02_out;
    92: reg_0959 <= op2_02_out;
    116: reg_0959 <= op2_02_out;
    121: reg_0959 <= imem00_in[11:8];
    endcase
  end

  // REG#960の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0960 <= imem06_in[15:12];
    68: reg_0960 <= op1_04_out;
    76: reg_0960 <= imem06_in[15:12];
    endcase
  end

  // REG#961の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0961 <= imem00_in[3:0];
    69: reg_0961 <= imem00_in[3:0];
    endcase
  end

  // REG#962の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0962 <= imem03_in[15:12];
    73: reg_0962 <= imem07_in[11:8];
    78: reg_0962 <= imem03_in[15:12];
    90: reg_0962 <= imem07_in[11:8];
    92: reg_0962 <= imem07_in[11:8];
    100: reg_0962 <= imem03_in[15:12];
    111: reg_0962 <= imem03_in[15:12];
    endcase
  end

  // REG#963の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0963 <= imem03_in[7:4];
    73: reg_0963 <= imem07_in[7:4];
    78: reg_0963 <= imem01_in[15:12];
    101: reg_0963 <= imem03_in[7:4];
    103: reg_0963 <= imem07_in[7:4];
    117: reg_0963 <= imem03_in[7:4];
    124: reg_0963 <= imem01_in[15:12];
    endcase
  end

  // REG#964の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0964 <= imem03_in[11:8];
    76: reg_0964 <= imem03_in[11:8];
    endcase
  end

  // REG#965の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0965 <= imem03_in[3:0];
    76: reg_0965 <= imem03_in[3:0];
    endcase
  end

  // REG#966の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0966 <= imem01_in[3:0];
    119: reg_0966 <= imem01_in[3:0];
    endcase
  end

  // REG#967の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0967 <= imem01_in[7:4];
    endcase
  end

  // REG#968の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0968 <= imem01_in[11:8];
    endcase
  end

  // REG#969の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0969 <= imem04_in[7:4];
    endcase
  end

  // REG#970の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0970 <= imem02_in[3:0];
    endcase
  end

  // REG#971の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0971 <= imem02_in[7:4];
    endcase
  end

  // REG#972の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0972 <= imem02_in[15:12];
    endcase
  end

  // REG#973の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0973 <= imem02_in[11:8];
    endcase
  end

  // REG#974の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0974 <= imem06_in[11:8];
    49: reg_0974 <= imem06_in[11:8];
    68: reg_0974 <= imem06_in[11:8];
    endcase
  end

  // REG#975の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0975 <= imem04_in[7:4];
    49: reg_0975 <= imem02_in[3:0];
    61: reg_0975 <= imem04_in[7:4];
    92: reg_0975 <= imem02_in[3:0];
    100: reg_0975 <= imem04_in[7:4];
    102: reg_0975 <= imem02_in[3:0];
    endcase
  end

  // REG#976の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0976 <= op2_00_out;
    49: reg_0976 <= imem02_in[15:12];
    61: reg_0976 <= imem02_in[15:12];
    82: reg_0976 <= op2_00_out;
    endcase
  end

  // REG#977の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0977 <= imem06_in[15:12];
    52: reg_0977 <= imem06_in[15:12];
    68: reg_0977 <= op1_05_out;
    76: reg_0977 <= op1_05_out;
    90: reg_0977 <= imem06_in[15:12];
    98: reg_0977 <= imem06_in[15:12];
    endcase
  end

  // REG#978の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0978 <= imem04_in[11:8];
    51: reg_0978 <= imem04_in[11:8];
    57: reg_0978 <= imem04_in[11:8];
    endcase
  end

  // REG#979の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0979 <= imem06_in[7:4];
    51: reg_0979 <= imem06_in[7:4];
    56: reg_0979 <= imem06_in[7:4];
    endcase
  end

  // REG#980の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0980 <= imem01_in[7:4];
    51: reg_0980 <= op1_01_out;
    79: reg_0980 <= op2_04_out;
    102: reg_0980 <= imem01_in[7:4];
    108: reg_0980 <= imem01_in[7:4];
    112: reg_0980 <= imem01_in[7:4];
    115: reg_0980 <= imem01_in[7:4];
    122: reg_0980 <= imem01_in[7:4];
    endcase
  end

  // REG#981の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0981 <= imem02_in[7:4];
    53: reg_0981 <= imem02_in[7:4];
    58: reg_0981 <= imem02_in[7:4];
    89: reg_0981 <= op2_11_out;
    endcase
  end

  // REG#982の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0982 <= imem01_in[15:12];
    53: reg_0982 <= imem01_in[15:12];
    68: reg_0982 <= op1_06_out;
    76: reg_0982 <= op1_06_out;
    79: reg_0982 <= imem01_in[15:12];
    81: reg_0982 <= imem01_in[15:12];
    87: reg_0982 <= op2_12_out;
    108: reg_0982 <= imem01_in[15:12];
    113: reg_0982 <= imem01_in[15:12];
    118: reg_0982 <= imem01_in[15:12];
    endcase
  end

  // REG#983の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0983 <= imem00_in[7:4];
    53: reg_0983 <= op1_11_out;
    75: reg_0983 <= imem00_in[7:4];
    92: reg_0983 <= imem00_in[7:4];
    94: reg_0983 <= imem00_in[7:4];
    97: reg_0983 <= imem00_in[7:4];
    105: reg_0983 <= imem00_in[7:4];
    107: reg_0983 <= imem00_in[7:4];
    112: reg_0983 <= imem00_in[7:4];
    115: reg_0983 <= imem00_in[7:4];
    126: reg_0983 <= imem00_in[7:4];
    endcase
  end

  // REG#984の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0984 <= imem01_in[3:0];
    54: reg_0984 <= imem01_in[3:0];
    73: reg_0984 <= imem06_in[3:0];
    79: reg_0984 <= imem06_in[3:0];
    85: reg_0984 <= imem06_in[3:0];
    endcase
  end

  // REG#985の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0985 <= imem01_in[11:8];
    53: reg_0985 <= op1_03_out;
    75: reg_0985 <= op1_03_out;
    77: reg_0985 <= op1_03_out;
    90: reg_0985 <= imem01_in[11:8];
    103: reg_0985 <= imem01_in[11:8];
    endcase
  end

  // REG#986の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0986 <= imem05_in[3:0];
    53: reg_0986 <= op1_04_out;
    76: reg_0986 <= imem05_in[3:0];
    95: reg_0986 <= imem05_in[3:0];
    107: reg_0986 <= imem05_in[3:0];
    111: reg_0986 <= imem05_in[3:0];
    114: reg_0986 <= imem05_in[3:0];
    endcase
  end

  // REG#987の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0987 <= imem00_in[3:0];
    55: reg_0987 <= imem00_in[3:0];
    endcase
  end

  // REG#988の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_0988 <= op1_00_out;
    54: reg_0988 <= op1_00_out;
    60: reg_0988 <= op1_00_out;
    69: reg_0988 <= op1_00_out;
    74: reg_0988 <= op1_00_out;
    89: reg_0988 <= op2_12_out;
    endcase
  end

  // REG#989の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0989 <= imem02_in[3:0];
    55: reg_0989 <= op1_07_out;
    71: reg_0989 <= op1_07_out;
    77: reg_0989 <= imem03_in[7:4];
    94: reg_0989 <= imem02_in[3:0];
    97: reg_0989 <= imem02_in[3:0];
    105: reg_0989 <= imem02_in[3:0];
    107: reg_0989 <= imem03_in[7:4];
    118: reg_0989 <= imem03_in[7:4];
    endcase
  end

  // REG#990の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0990 <= imem02_in[11:8];
    55: reg_0990 <= op1_02_out;
    74: reg_0990 <= op1_02_out;
    76: reg_0990 <= op2_01_out;
    109: reg_0990 <= op2_01_out;
    endcase
  end

  // REG#991の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0991 <= imem02_in[15:12];
    55: reg_0991 <= op1_03_out;
    74: reg_0991 <= op2_02_out;
    78: reg_0991 <= op2_02_out;
    83: reg_0991 <= op2_02_out;
    endcase
  end

  // REG#992の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0992 <= imem05_in[15:12];
    57: reg_0992 <= imem05_in[15:12];
    endcase
  end

  // REG#993の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0993 <= imem07_in[7:4];
    57: reg_0993 <= imem07_in[7:4];
    66: reg_0993 <= op1_00_out;
    94: reg_0993 <= imem07_in[7:4];
    98: reg_0993 <= imem07_in[7:4];
    102: reg_0993 <= imem07_in[7:4];
    107: reg_0993 <= imem07_in[7:4];
    110: reg_0993 <= imem07_in[7:4];
    113: reg_0993 <= imem07_in[7:4];
    endcase
  end

  // REG#994の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0994 <= imem07_in[3:0];
    57: reg_0994 <= imem07_in[3:0];
    66: reg_0994 <= op1_01_out;
    95: reg_0994 <= imem07_in[3:0];
    endcase
  end

  // REG#995の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0995 <= imem07_in[15:12];
    57: reg_0995 <= imem07_in[15:12];
    66: reg_0995 <= op1_02_out;
    93: reg_0995 <= imem07_in[15:12];
    102: reg_0995 <= imem07_in[15:12];
    104: reg_0995 <= imem07_in[15:12];
    112: reg_0995 <= imem07_in[15:12];
    114: reg_0995 <= imem07_in[15:12];
    117: reg_0995 <= imem07_in[15:12];
    endcase
  end

  // REG#996の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0996 <= imem05_in[7:4];
    57: reg_0996 <= imem05_in[7:4];
    endcase
  end

  // REG#997の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0997 <= imem05_in[11:8];
    57: reg_0997 <= imem02_in[15:12];
    64: reg_0997 <= imem02_in[15:12];
    74: reg_0997 <= imem07_in[11:8];
    77: reg_0997 <= op2_02_out;
    124: reg_0997 <= op2_02_out;
    endcase
  end

  // REG#998の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0998 <= imem07_in[11:8];
    57: reg_0998 <= imem07_in[11:8];
    66: reg_0998 <= op1_04_out;
    93: reg_0998 <= imem07_in[11:8];
    101: reg_0998 <= imem07_in[11:8];
    105: reg_0998 <= imem07_in[11:8];
    118: reg_0998 <= imem07_in[11:8];
    endcase
  end

  // REG#999の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_0999 <= imem03_in[11:8];
    73: reg_0999 <= imem03_in[11:8];
    104: reg_0999 <= imem03_in[11:8];
    114: reg_0999 <= imem03_in[11:8];
    117: reg_0999 <= imem03_in[11:8];
    endcase
  end

  // REG#1000の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1000 <= imem03_in[3:0];
    73: reg_1000 <= imem03_in[3:0];
    103: reg_1000 <= imem03_in[3:0];
    108: reg_1000 <= imem03_in[3:0];
    112: reg_1000 <= imem03_in[3:0];
    endcase
  end

  // REG#1001の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1001 <= imem03_in[7:4];
    72: reg_1001 <= op1_00_out;
    79: reg_1001 <= imem03_in[7:4];
    endcase
  end

  // REG#1002の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1002 <= op1_01_out;
    71: reg_1002 <= op1_01_out;
    74: reg_1002 <= op1_01_out;
    89: reg_1002 <= imem02_in[7:4];
    106: reg_1002 <= imem02_in[7:4];
    111: reg_1002 <= imem02_in[7:4];
    endcase
  end

  // REG#1003の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1003 <= imem03_in[15:12];
    77: reg_1003 <= imem03_in[15:12];
    102: reg_1003 <= imem03_in[15:12];
    endcase
  end

  // REG#1004の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1004 <= op1_04_out;
    80: reg_1004 <= imem04_in[15:12];
    endcase
  end

  // REG#1005の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1005 <= op1_05_out;
    80: reg_1005 <= op2_07_out;
    endcase
  end

  // REG#1006の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1006 <= op1_06_out;
    81: reg_1006 <= imem02_in[11:8];
    endcase
  end

  // REG#1007の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1007 <= op1_08_out;
    83: reg_1007 <= op1_08_out;
    86: reg_1007 <= op1_08_out;
    88: reg_1007 <= op1_08_out;
    90: reg_1007 <= op1_08_out;
    endcase
  end

  // REG#1008の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1008 <= op1_10_out;
    82: reg_1008 <= op1_10_out;
    endcase
  end

  // REG#1009の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1009 <= op1_13_out;
    87: reg_1009 <= op1_13_out;
    90: reg_1009 <= imem03_in[15:12];
    125: reg_1009 <= imem03_in[15:12];
    endcase
  end

  // REG#1010の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1010 <= op1_02_out;
    89: reg_1010 <= imem07_in[15:12];
    113: reg_1010 <= imem07_in[15:12];
    endcase
  end

  // REG#1011の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1011 <= op1_03_out;
    89: reg_1011 <= op2_13_out;
    endcase
  end

  // REG#1012の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1012 <= op1_07_out;
    endcase
  end

  // REG#1013の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1013 <= op1_09_out;
    90: reg_1013 <= op1_09_out;
    endcase
  end

  // REG#1014の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1014 <= op1_11_out;
    endcase
  end

  // REG#1015の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1015 <= op1_12_out;
    110: reg_1015 <= op1_12_out;
    112: reg_1015 <= op1_12_out;
    endcase
  end

  // REG#1016の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1016 <= op1_14_out;
    104: reg_1016 <= op1_14_out;
    114: reg_1016 <= op1_14_out;
    118: reg_1016 <= op1_14_out;
    endcase
  end

  // REG#1017の入力
  always @ ( posedge clock ) begin
    case ( state )
    46: reg_1017 <= op1_15_out;
    102: reg_1017 <= op1_15_out;
    109: reg_1017 <= op1_15_out;
    endcase
  end

  // REG#1018の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1018 <= imem02_in[15:12];
    101: reg_1018 <= imem02_in[15:12];
    endcase
  end

  // REG#1019の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1019 <= op1_08_out;
    endcase
  end

  // REG#1020の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1020 <= op1_09_out;
    endcase
  end

  // REG#1021の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1021 <= op1_10_out;
    endcase
  end

  // REG#1022の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1022 <= op1_11_out;
    endcase
  end

  // REG#1023の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1023 <= op1_12_out;
    endcase
  end

  // REG#1024の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1024 <= op1_13_out;
    endcase
  end

  // REG#1025の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1025 <= op1_14_out;
    endcase
  end

  // REG#1026の入力
  always @ ( posedge clock ) begin
    case ( state )
    47: reg_1026 <= op1_15_out;
    endcase
  end

  // REG#1027の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1027 <= imem00_in[11:8];
    endcase
  end

  // REG#1028の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1028 <= imem00_in[7:4];
    endcase
  end

  // REG#1029の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1029 <= imem02_in[11:8];
    61: reg_1029 <= imem02_in[11:8];
    endcase
  end

  // REG#1030の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1030 <= imem06_in[3:0];
    61: reg_1030 <= op1_02_out;
    89: reg_1030 <= imem06_in[3:0];
    108: reg_1030 <= imem06_in[3:0];
    110: reg_1030 <= imem06_in[3:0];
    125: reg_1030 <= imem06_in[3:0];
    endcase
  end

  // REG#1031の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1031 <= imem01_in[11:8];
    64: reg_1031 <= imem01_in[11:8];
    76: reg_1031 <= imem02_in[11:8];
    92: reg_1031 <= imem01_in[11:8];
    110: reg_1031 <= imem01_in[11:8];
    117: reg_1031 <= imem01_in[11:8];
    endcase
  end

  // REG#1032の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1032 <= imem01_in[3:0];
    64: reg_1032 <= imem01_in[3:0];
    76: reg_1032 <= imem02_in[3:0];
    92: reg_1032 <= imem01_in[3:0];
    104: reg_1032 <= imem01_in[3:0];
    113: reg_1032 <= imem01_in[3:0];
    120: reg_1032 <= imem01_in[3:0];
    endcase
  end

  // REG#1033の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1033 <= imem01_in[7:4];
    64: reg_1033 <= imem03_in[7:4];
    80: reg_1033 <= imem03_in[7:4];
    endcase
  end

  // REG#1034の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1034 <= imem01_in[15:12];
    65: reg_1034 <= imem01_in[15:12];
    80: reg_1034 <= imem01_in[15:12];
    82: reg_1034 <= imem01_in[15:12];
    87: reg_1034 <= op2_13_out;
    109: reg_1034 <= imem01_in[15:12];
    120: reg_1034 <= imem01_in[15:12];
    endcase
  end

  // REG#1035の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1035 <= imem06_in[15:12];
    66: reg_1035 <= imem06_in[15:12];
    80: reg_1035 <= imem06_in[15:12];
    103: reg_1035 <= imem06_in[15:12];
    105: reg_1035 <= imem06_in[15:12];
    107: reg_1035 <= imem06_in[15:12];
    110: reg_1035 <= imem06_in[15:12];
    endcase
  end

  // REG#1036の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1036 <= imem06_in[7:4];
    67: reg_1036 <= op1_07_out;
    116: reg_1036 <= imem06_in[7:4];
    endcase
  end

  // REG#1037の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1037 <= op1_02_out;
    74: reg_1037 <= op2_03_out;
    83: reg_1037 <= op2_03_out;
    85: reg_1037 <= op1_02_out;
    92: reg_1037 <= op2_03_out;
    124: reg_1037 <= op2_03_out;
    endcase
  end

  // REG#1038の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1038 <= op1_03_out;
    75: reg_1038 <= op2_03_out;
    109: reg_1038 <= op2_03_out;
    endcase
  end

  // REG#1039の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1039 <= op1_04_out;
    80: reg_1039 <= op1_04_out;
    86: reg_1039 <= op1_04_out;
    88: reg_1039 <= op2_01_out;
    112: reg_1039 <= op2_01_out;
    endcase
  end

  // REG#1040の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1040 <= op1_05_out;
    81: reg_1040 <= imem04_in[11:8];
    endcase
  end

  // REG#1041の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1041 <= op1_06_out;
    81: reg_1041 <= imem04_in[3:0];
    endcase
  end

  // REG#1042の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1042 <= op1_08_out;
    84: reg_1042 <= op1_08_out;
    87: reg_1042 <= op2_14_out;
    endcase
  end

  // REG#1043の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1043 <= op1_09_out;
    83: reg_1043 <= op1_09_out;
    86: reg_1043 <= op1_09_out;
    88: reg_1043 <= op1_09_out;
    endcase
  end

  // REG#1044の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1044 <= op1_11_out;
    86: reg_1044 <= op1_11_out;
    88: reg_1044 <= op1_11_out;
    90: reg_1044 <= op1_11_out;
    endcase
  end

  // REG#1045の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1045 <= op1_01_out;
    88: reg_1045 <= op2_03_out;
    114: reg_1045 <= op2_03_out;
    endcase
  end

  // REG#1046の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1046 <= op1_07_out;
    endcase
  end

  // REG#1047の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1047 <= op1_10_out;
    endcase
  end

  // REG#1048の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1048 <= op1_12_out;
    endcase
  end

  // REG#1049の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1049 <= op1_13_out;
    97: reg_1049 <= op1_13_out;
    100: reg_1049 <= op1_13_out;
    104: reg_1049 <= op1_13_out;
    endcase
  end

  // REG#1050の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1050 <= op1_14_out;
    endcase
  end

  // REG#1051の入力
  always @ ( posedge clock ) begin
    case ( state )
    48: reg_1051 <= op1_15_out;
    endcase
  end

  // REG#1052の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1052 <= imem00_in[7:4];
    endcase
  end

  // REG#1053の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1053 <= imem00_in[3:0];
    endcase
  end

  // REG#1054の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1054 <= op1_00_out;
    55: reg_1054 <= op1_00_out;
    70: reg_1054 <= op1_07_out;
    80: reg_1054 <= op1_07_out;
    82: reg_1054 <= op1_07_out;
    endcase
  end

  // REG#1055の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1055 <= imem07_in[7:4];
    58: reg_1055 <= imem07_in[7:4];
    67: reg_1055 <= op1_08_out;
    95: reg_1055 <= imem07_in[7:4];
    endcase
  end

  // REG#1056の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1056 <= imem07_in[11:8];
    58: reg_1056 <= imem07_in[11:8];
    68: reg_1056 <= op1_08_out;
    77: reg_1056 <= imem07_in[11:8];
    80: reg_1056 <= op1_08_out;
    83: reg_1056 <= imem07_in[11:8];
    87: reg_1056 <= imem07_in[11:8];
    endcase
  end

  // REG#1057の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1057 <= imem07_in[3:0];
    58: reg_1057 <= imem07_in[3:0];
    64: reg_1057 <= op1_03_out;
    98: reg_1057 <= imem07_in[3:0];
    102: reg_1057 <= imem07_in[3:0];
    108: reg_1057 <= imem07_in[3:0];
    110: reg_1057 <= imem07_in[3:0];
    113: reg_1057 <= imem07_in[3:0];
    endcase
  end

  // REG#1058の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1058 <= imem06_in[11:8];
    57: reg_1058 <= op1_12_out;
    79: reg_1058 <= op1_12_out;
    84: reg_1058 <= op1_12_out;
    86: reg_1058 <= op1_12_out;
    89: reg_1058 <= imem06_in[11:8];
    110: reg_1058 <= imem06_in[11:8];
    endcase
  end

  // REG#1059の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1059 <= imem05_in[3:0];
    57: reg_1059 <= op1_13_out;
    80: reg_1059 <= op1_13_out;
    90: reg_1059 <= op1_13_out;
    92: reg_1059 <= op1_13_out;
    96: reg_1059 <= imem05_in[3:0];
    122: reg_1059 <= imem05_in[3:0];
    endcase
  end

  // REG#1060の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1060 <= imem07_in[15:12];
    57: reg_1060 <= op1_15_out;
    80: reg_1060 <= op1_15_out;
    91: reg_1060 <= op1_15_out;
    95: reg_1060 <= imem07_in[15:12];
    endcase
  end

  // REG#1061の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1061 <= op1_14_out;
    62: reg_1061 <= op1_14_out;
    83: reg_1061 <= op1_14_out;
    92: reg_1061 <= op1_14_out;
    endcase
  end

  // REG#1062の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1062 <= op1_01_out;
    69: reg_1062 <= op1_01_out;
    75: reg_1062 <= op2_04_out;
    endcase
  end

  // REG#1063の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1063 <= imem03_in[7:4];
    70: reg_1063 <= op1_08_out;
    81: reg_1063 <= imem03_in[7:4];
    endcase
  end

  // REG#1064の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1064 <= imem03_in[15:12];
    71: reg_1064 <= imem06_in[15:12];
    82: reg_1064 <= imem06_in[15:12];
    99: reg_1064 <= imem06_in[15:12];
    114: reg_1064 <= imem06_in[15:12];
    endcase
  end

  // REG#1065の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1065 <= imem04_in[7:4];
    73: reg_1065 <= imem06_in[15:12];
    80: reg_1065 <= imem04_in[7:4];
    endcase
  end

  // REG#1066の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1066 <= op1_05_out;
    74: reg_1066 <= op1_05_out;
    76: reg_1066 <= op2_02_out;
    110: reg_1066 <= op2_02_out;
    endcase
  end

  // REG#1067の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1067 <= op1_07_out;
    75: reg_1067 <= op1_07_out;
    89: reg_1067 <= op1_07_out;
    endcase
  end

  // REG#1068の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1068 <= imem01_in[3:0];
    77: reg_1068 <= imem01_in[3:0];
    83: reg_1068 <= imem01_in[3:0];
    endcase
  end

  // REG#1069の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1069 <= imem01_in[11:8];
    76: reg_1069 <= op2_03_out;
    116: reg_1069 <= op2_03_out;
    endcase
  end

  // REG#1070の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1070 <= imem01_in[7:4];
    77: reg_1070 <= imem05_in[7:4];
    endcase
  end

  // REG#1071の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1071 <= imem01_in[15:12];
    77: reg_1071 <= imem01_in[15:12];
    83: reg_1071 <= imem01_in[15:12];
    endcase
  end

  // REG#1072の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1072 <= op1_08_out;
    76: reg_1072 <= op1_08_out;
    78: reg_1072 <= op1_08_out;
    endcase
  end

  // REG#1073の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1073 <= op1_09_out;
    76: reg_1073 <= op1_09_out;
    78: reg_1073 <= op1_09_out;
    80: reg_1073 <= op1_09_out;
    endcase
  end

  // REG#1074の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1074 <= op1_11_out;
    77: reg_1074 <= imem02_in[15:12];
    endcase
  end

  // REG#1075の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1075 <= op1_10_out;
    77: reg_1075 <= op1_10_out;
    endcase
  end

  // REG#1076の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1076 <= op1_13_out;
    77: reg_1076 <= op1_13_out;
    endcase
  end

  // REG#1077の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1077 <= imem04_in[3:0];
    80: reg_1077 <= imem04_in[3:0];
    endcase
  end

  // REG#1078の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1078 <= imem00_in[11:8];
    81: reg_1078 <= imem02_in[7:4];
    endcase
  end

  // REG#1079の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1079 <= imem00_in[3:0];
    82: reg_1079 <= imem00_in[3:0];
    106: reg_1079 <= imem00_in[3:0];
    108: reg_1079 <= imem00_in[3:0];
    114: reg_1079 <= imem00_in[3:0];
    121: reg_1079 <= imem00_in[3:0];
    endcase
  end

  // REG#1080の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1080 <= imem00_in[7:4];
    85: reg_1080 <= imem00_in[7:4];
    87: reg_1080 <= op2_15_out;
    109: reg_1080 <= imem00_in[7:4];
    111: reg_1080 <= imem00_in[7:4];
    116: reg_1080 <= imem00_in[7:4];
    118: reg_1080 <= imem00_in[7:4];
    120: reg_1080 <= imem00_in[7:4];
    123: reg_1080 <= imem00_in[7:4];
    endcase
  end

  // REG#1081の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1081 <= imem00_in[15:12];
    84: reg_1081 <= imem00_in[15:12];
    89: reg_1081 <= imem00_in[15:12];
    93: reg_1081 <= imem00_in[15:12];
    106: reg_1081 <= imem00_in[15:12];
    113: reg_1081 <= imem00_in[15:12];
    115: reg_1081 <= imem00_in[15:12];
    125: reg_1081 <= imem00_in[15:12];
    endcase
  end

  // REG#1082の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1082 <= imem04_in[15:12];
    83: reg_1082 <= imem04_in[15:12];
    endcase
  end

  // REG#1083の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1083 <= imem04_in[11:8];
    85: reg_1083 <= imem04_in[11:8];
    endcase
  end

  // REG#1084の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1084 <= op1_02_out;
    88: reg_1084 <= op2_04_out;
    endcase
  end

  // REG#1085の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1085 <= op1_03_out;
    88: reg_1085 <= op2_05_out;
    endcase
  end

  // REG#1086の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1086 <= op1_04_out;
    88: reg_1086 <= op2_06_out;
    endcase
  end

  // REG#1087の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1087 <= op1_06_out;
    88: reg_1087 <= op2_07_out;
    endcase
  end

  // REG#1088の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1088 <= op1_12_out;
    89: reg_1088 <= op2_14_out;
    endcase
  end

  // REG#1089の入力
  always @ ( posedge clock ) begin
    case ( state )
    49: reg_1089 <= op1_15_out;
    92: reg_1089 <= op1_15_out;
    endcase
  end

  // REG#1090の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1090 <= imem01_in[15:12];
    53: reg_1090 <= op1_13_out;
    75: reg_1090 <= op1_13_out;
    90: reg_1090 <= imem01_in[15:12];
    99: reg_1090 <= imem01_in[15:12];
    115: reg_1090 <= imem01_in[15:12];
    endcase
  end

  // REG#1091の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1091 <= imem03_in[15:12];
    53: reg_1091 <= op1_01_out;
    81: reg_1091 <= imem02_in[15:12];
    endcase
  end

  // REG#1092の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1092 <= imem03_in[7:4];
    55: reg_1092 <= imem03_in[7:4];
    endcase
  end

  // REG#1093の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1093 <= imem03_in[11:8];
    56: reg_1093 <= imem03_in[11:8];
    endcase
  end

  // REG#1094の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1094 <= imem07_in[15:12];
    59: reg_1094 <= imem07_in[15:12];
    endcase
  end

  // REG#1095の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1095 <= imem07_in[11:8];
    58: reg_1095 <= op1_07_out;
    81: reg_1095 <= op1_07_out;
    84: reg_1095 <= imem07_in[11:8];
    106: reg_1095 <= imem07_in[11:8];
    111: reg_1095 <= imem07_in[11:8];
    endcase
  end

  // REG#1096の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1096 <= imem07_in[7:4];
    58: reg_1096 <= op1_13_out;
    81: reg_1096 <= op1_13_out;
    83: reg_1096 <= op1_13_out;
    85: reg_1096 <= op1_13_out;
    88: reg_1096 <= imem07_in[7:4];
    96: reg_1096 <= imem07_in[7:4];
    99: reg_1096 <= imem07_in[7:4];
    105: reg_1096 <= imem07_in[7:4];
    115: reg_1096 <= imem07_in[7:4];
    endcase
  end

  // REG#1097の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1097 <= imem07_in[3:0];
    58: reg_1097 <= op1_14_out;
    81: reg_1097 <= op1_14_out;
    84: reg_1097 <= imem07_in[3:0];
    105: reg_1097 <= imem07_in[3:0];
    117: reg_1097 <= imem07_in[3:0];
    endcase
  end

  // REG#1098の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1098 <= imem02_in[11:8];
    59: reg_1098 <= op1_05_out;
    84: reg_1098 <= imem02_in[11:8];
    endcase
  end

  // REG#1099の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1099 <= imem00_in[7:4];
    60: reg_1099 <= op1_03_out;
    78: reg_1099 <= op1_03_out;
    91: reg_1099 <= imem00_in[7:4];
    93: reg_1099 <= imem00_in[7:4];
    100: reg_1099 <= imem00_in[7:4];
    endcase
  end

  // REG#1100の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1100 <= imem00_in[3:0];
    61: reg_1100 <= imem00_in[3:0];
    endcase
  end

  // REG#1101の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1101 <= imem00_in[11:8];
    60: reg_1101 <= op1_05_out;
    84: reg_1101 <= op1_05_out;
    89: reg_1101 <= imem00_in[11:8];
    99: reg_1101 <= imem00_in[11:8];
    102: reg_1101 <= imem00_in[11:8];
    122: reg_1101 <= imem00_in[11:8];
    endcase
  end

  // REG#1102の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1102 <= imem00_in[15:12];
    60: reg_1102 <= op1_06_out;
    78: reg_1102 <= op1_06_out;
    119: reg_1102 <= imem00_in[15:12];
    126: reg_1102 <= imem00_in[15:12];
    endcase
  end

  // REG#1103の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1103 <= imem02_in[3:0];
    61: reg_1103 <= imem02_in[3:0];
    88: reg_1103 <= op2_08_out;
    123: reg_1103 <= imem02_in[3:0];
    endcase
  end

  // REG#1104の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1104 <= imem05_in[3:0];
    60: reg_1104 <= op1_07_out;
    81: reg_1104 <= imem05_in[3:0];
    endcase
  end

  // REG#1105の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1105 <= imem06_in[3:0];
    66: reg_1105 <= imem06_in[3:0];
    82: reg_1105 <= imem06_in[3:0];
    99: reg_1105 <= imem06_in[3:0];
    endcase
  end

  // REG#1106の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1106 <= op1_11_out;
    73: reg_1106 <= op2_01_out;
    80: reg_1106 <= op2_01_out;
    104: reg_1106 <= op2_01_out;
    121: reg_1106 <= op2_01_out;
    endcase
  end

  // REG#1107の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1107 <= op1_02_out;
    76: reg_1107 <= imem04_in[7:4];
    endcase
  end

  // REG#1108の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1108 <= op1_05_out;
    75: reg_1108 <= op1_05_out;
    77: reg_1108 <= op1_05_out;
    85: reg_1108 <= op1_05_out;
    endcase
  end

  // REG#1109の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1109 <= op1_06_out;
    75: reg_1109 <= op1_06_out;
    endcase
  end

  // REG#1110の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1110 <= op1_08_out;
    77: reg_1110 <= op1_08_out;
    88: reg_1110 <= op2_09_out;
    endcase
  end

  // REG#1111の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1111 <= op1_12_out;
    78: reg_1111 <= op1_12_out;
    80: reg_1111 <= op1_12_out;
    endcase
  end

  // REG#1112の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1112 <= op1_14_out;
    78: reg_1112 <= op1_14_out;
    endcase
  end

  // REG#1113の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1113 <= op1_15_out;
    83: reg_1113 <= op1_15_out;
    endcase
  end

  // REG#1114の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1114 <= op1_00_out;
    endcase
  end

  // REG#1115の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1115 <= op1_01_out;
    endcase
  end

  // REG#1116の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1116 <= op1_03_out;
    endcase
  end

  // REG#1117の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1117 <= op1_04_out;
    endcase
  end

  // REG#1118の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1118 <= op1_07_out;
    88: reg_1118 <= op1_07_out;
    endcase
  end

  // REG#1119の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1119 <= op1_09_out;
    endcase
  end

  // REG#1120の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1120 <= op1_10_out;
    endcase
  end

  // REG#1121の入力
  always @ ( posedge clock ) begin
    case ( state )
    50: reg_1121 <= op1_13_out;
    endcase
  end

  // REG#1122の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1122 <= op1_03_out;
    86: reg_1122 <= op1_03_out;
    endcase
  end

  // REG#1123の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1123 <= op1_04_out;
    87: reg_1123 <= op1_04_out;
    endcase
  end

  // REG#1124の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1124 <= op1_05_out;
    endcase
  end

  // REG#1125の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1125 <= op1_07_out;
    83: reg_1125 <= op1_07_out;
    86: reg_1125 <= op1_07_out;
    endcase
  end

  // REG#1126の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1126 <= op1_08_out;
    endcase
  end

  // REG#1127の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1127 <= op1_10_out;
    83: reg_1127 <= op1_10_out;
    endcase
  end

  // REG#1128の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1128 <= op1_11_out;
    84: reg_1128 <= op1_11_out;
    endcase
  end

  // REG#1129の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1129 <= op1_12_out;
    endcase
  end

  // REG#1130の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1130 <= op1_14_out;
    82: reg_1130 <= op1_14_out;
    84: reg_1130 <= op1_14_out;
    endcase
  end

  // REG#1131の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1131 <= op1_15_out;
    85: reg_1131 <= op1_15_out;
    87: reg_1131 <= op1_15_out;
    endcase
  end

  // REG#1132の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1132 <= imem03_in[3:0];
    120: reg_1132 <= imem03_in[3:0];
    endcase
  end

  // REG#1133の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1133 <= op1_00_out;
    endcase
  end

  // REG#1134の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1134 <= op1_02_out;
    endcase
  end

  // REG#1135の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1135 <= op1_06_out;
    endcase
  end

  // REG#1136の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1136 <= op1_09_out;
    endcase
  end

  // REG#1137の入力
  always @ ( posedge clock ) begin
    case ( state )
    51: reg_1137 <= op1_13_out;
    endcase
  end

  // REG#1138の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1138 <= op1_01_out;
    54: reg_1138 <= op1_01_out;
    70: reg_1138 <= op1_01_out;
    endcase
  end

  // REG#1139の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1139 <= imem02_in[15:12];
    59: reg_1139 <= imem02_in[15:12];
    63: reg_1139 <= imem03_in[3:0];
    73: reg_1139 <= imem02_in[15:12];
    85: reg_1139 <= imem03_in[3:0];
    endcase
  end

  // REG#1140の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1140 <= imem02_in[3:0];
    59: reg_1140 <= imem02_in[3:0];
    64: reg_1140 <= imem02_in[3:0];
    72: reg_1140 <= op1_04_out;
    91: reg_1140 <= imem02_in[3:0];
    endcase
  end

  // REG#1141の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1141 <= imem00_in[11:8];
    60: reg_1141 <= op1_08_out;
    90: reg_1141 <= imem00_in[11:8];
    100: reg_1141 <= imem00_in[11:8];
    endcase
  end

  // REG#1142の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1142 <= op1_02_out;
    60: reg_1142 <= op1_02_out;
    63: reg_1142 <= op1_02_out;
    endcase
  end

  // REG#1143の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1143 <= imem04_in[7:4];
    61: reg_1143 <= op1_03_out;
    95: reg_1143 <= imem04_in[7:4];
    endcase
  end

  // REG#1144の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1144 <= imem04_in[3:0];
    61: reg_1144 <= op1_05_out;
    89: reg_1144 <= imem04_in[3:0];
    93: reg_1144 <= imem04_in[3:0];
    101: reg_1144 <= imem04_in[3:0];
    107: reg_1144 <= imem04_in[3:0];
    116: reg_1144 <= imem04_in[3:0];
    119: reg_1144 <= imem04_in[3:0];
    129: reg_1144 <= imem04_in[3:0];
    endcase
  end

  // REG#1145の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1145 <= imem03_in[7:4];
    61: reg_1145 <= op1_06_out;
    92: reg_1145 <= imem03_in[7:4];
    102: reg_1145 <= imem03_in[7:4];
    endcase
  end

  // REG#1146の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1146 <= imem04_in[15:12];
    61: reg_1146 <= op1_07_out;
    93: reg_1146 <= imem04_in[15:12];
    101: reg_1146 <= imem04_in[15:12];
    108: reg_1146 <= imem04_in[15:12];
    endcase
  end

  // REG#1147の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1147 <= imem04_in[11:8];
    62: reg_1147 <= imem04_in[11:8];
    82: reg_1147 <= imem04_in[11:8];
    endcase
  end

  // REG#1148の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1148 <= imem00_in[15:12];
    64: reg_1148 <= op1_04_out;
    endcase
  end

  // REG#1149の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1149 <= imem03_in[11:8];
    65: reg_1149 <= imem03_in[11:8];
    87: reg_1149 <= imem03_in[11:8];
    endcase
  end

  // REG#1150の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1150 <= imem07_in[11:8];
    66: reg_1150 <= op1_05_out;
    endcase
  end

  // REG#1151の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1151 <= imem01_in[3:0];
    69: reg_1151 <= imem04_in[3:0];
    78: reg_1151 <= imem04_in[3:0];
    endcase
  end

  // REG#1152の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1152 <= imem01_in[7:4];
    68: reg_1152 <= op1_07_out;
    77: reg_1152 <= op1_07_out;
    90: reg_1152 <= imem01_in[7:4];
    103: reg_1152 <= imem01_in[7:4];
    endcase
  end

  // REG#1153の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1153 <= op1_03_out;
    76: reg_1153 <= op1_03_out;
    endcase
  end

  // REG#1154の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1154 <= op1_04_out;
    endcase
  end

  // REG#1155の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1155 <= op1_05_out;
    endcase
  end

  // REG#1156の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1156 <= op1_08_out;
    endcase
  end

  // REG#1157の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1157 <= op1_09_out;
    endcase
  end

  // REG#1158の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1158 <= op1_10_out;
    84: reg_1158 <= op1_10_out;
    endcase
  end

  // REG#1159の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1159 <= op1_11_out;
    endcase
  end

  // REG#1160の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1160 <= op1_12_out;
    endcase
  end

  // REG#1161の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1161 <= op1_14_out;
    85: reg_1161 <= op1_14_out;
    87: reg_1161 <= op1_14_out;
    endcase
  end

  // REG#1162の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1162 <= op1_15_out;
    86: reg_1162 <= op1_15_out;
    88: reg_1162 <= op1_15_out;
    endcase
  end

  // REG#1163の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1163 <= imem05_in[15:12];
    103: reg_1163 <= imem05_in[15:12];
    endcase
  end

  // REG#1164の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1164 <= imem05_in[7:4];
    92: reg_1164 <= imem05_in[7:4];
    endcase
  end

  // REG#1165の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1165 <= op1_06_out;
    endcase
  end

  // REG#1166の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1166 <= op1_07_out;
    endcase
  end

  // REG#1167の入力
  always @ ( posedge clock ) begin
    case ( state )
    52: reg_1167 <= op1_13_out;
    endcase
  end

  // REG#1168の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1168 <= imem05_in[3:0];
    104: reg_1168 <= imem05_in[3:0];
    116: reg_1168 <= imem05_in[3:0];
    119: reg_1168 <= imem05_in[3:0];
    endcase
  end

  // REG#1169の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1169 <= imem05_in[11:8];
    93: reg_1169 <= imem05_in[11:8];
    98: reg_1169 <= imem05_in[11:8];
    103: reg_1169 <= imem05_in[11:8];
    endcase
  end

  // REG#1170の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1170 <= imem06_in[3:0];
    endcase
  end

  // REG#1171の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1171 <= op1_05_out;
    endcase
  end

  // REG#1172の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1172 <= op1_06_out;
    endcase
  end

  // REG#1173の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1173 <= op1_07_out;
    endcase
  end

  // REG#1174の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1174 <= op1_08_out;
    endcase
  end

  // REG#1175の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1175 <= op1_09_out;
    endcase
  end

  // REG#1176の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1176 <= op1_12_out;
    endcase
  end

  // REG#1177の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1177 <= op1_15_out;
    endcase
  end

  // REG#1178の入力
  always @ ( posedge clock ) begin
    case ( state )
    53: reg_1178 <= op1_14_out;
    endcase
  end

  // REG#1179の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1179 <= imem06_in[3:0];
    101: reg_1179 <= imem06_in[3:0];
    endcase
  end

  // REG#1180の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1180 <= imem05_in[11:8];
    endcase
  end

  // REG#1181の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1181 <= imem05_in[7:4];
    endcase
  end

  // REG#1182の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1182 <= imem07_in[3:0];
    endcase
  end

  // REG#1183の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1183 <= imem07_in[7:4];
    62: reg_1183 <= imem07_in[7:4];
    89: reg_1183 <= imem07_in[7:4];
    111: reg_1183 <= imem07_in[7:4];
    endcase
  end

  // REG#1184の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1184 <= op1_04_out;
    76: reg_1184 <= imem03_in[7:4];
    endcase
  end

  // REG#1185の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1185 <= op1_06_out;
    77: reg_1185 <= op1_06_out;
    endcase
  end

  // REG#1186の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1186 <= op1_09_out;
    77: reg_1186 <= op2_03_out;
    endcase
  end

  // REG#1187の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1187 <= op1_10_out;
    76: reg_1187 <= op1_10_out;
    endcase
  end

  // REG#1188の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1188 <= op1_11_out;
    77: reg_1188 <= op1_11_out;
    endcase
  end

  // REG#1189の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1189 <= op1_13_out;
    78: reg_1189 <= imem04_in[15:12];
    endcase
  end

  // REG#1190の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1190 <= op1_02_out;
    endcase
  end

  // REG#1191の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1191 <= op1_03_out;
    endcase
  end

  // REG#1192の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1192 <= op1_05_out;
    endcase
  end

  // REG#1193の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1193 <= op1_07_out;
    endcase
  end

  // REG#1194の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1194 <= op1_08_out;
    endcase
  end

  // REG#1195の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1195 <= op1_12_out;
    endcase
  end

  // REG#1196の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1196 <= op1_14_out;
    endcase
  end

  // REG#1197の入力
  always @ ( posedge clock ) begin
    case ( state )
    54: reg_1197 <= op1_15_out;
    endcase
  end

  // REG#1198の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1198 <= imem04_in[7:4];
    endcase
  end

  // REG#1199の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1199 <= imem03_in[3:0];
    endcase
  end

  // REG#1200の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1200 <= imem04_in[15:12];
    endcase
  end

  // REG#1201の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1201 <= imem00_in[7:4];
    endcase
  end

  // REG#1202の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1202 <= imem06_in[11:8];
    endcase
  end

  // REG#1203の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1203 <= imem04_in[3:0];
    endcase
  end

  // REG#1204の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1204 <= imem06_in[3:0];
    endcase
  end

  // REG#1205の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1205 <= imem00_in[11:8];
    endcase
  end

  // REG#1206の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1206 <= imem00_in[15:12];
    endcase
  end

  // REG#1207の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1207 <= imem02_in[11:8];
    endcase
  end

  // REG#1208の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1208 <= imem03_in[15:12];
    endcase
  end

  // REG#1209の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1209 <= op1_05_out;
    76: reg_1209 <= imem06_in[11:8];
    endcase
  end

  // REG#1210の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1210 <= op1_11_out;
    75: reg_1210 <= op1_11_out;
    endcase
  end

  // REG#1211の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1211 <= op1_12_out;
    75: reg_1211 <= op1_12_out;
    endcase
  end

  // REG#1212の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1212 <= imem05_in[11:8];
    77: reg_1212 <= op2_04_out;
    endcase
  end

  // REG#1213の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1213 <= op1_14_out;
    76: reg_1213 <= op1_14_out;
    79: reg_1213 <= op1_14_out;
    86: reg_1213 <= op1_14_out;
    88: reg_1213 <= op1_14_out;
    endcase
  end

  // REG#1214の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1214 <= imem04_in[11:8];
    83: reg_1214 <= imem04_in[11:8];
    endcase
  end

  // REG#1215の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1215 <= imem04_in[7:4];
    84: reg_1215 <= imem04_in[7:4];
    endcase
  end

  // REG#1216の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1216 <= imem04_in[15:12];
    109: reg_1216 <= imem04_in[15:12];
    117: reg_1216 <= imem04_in[15:12];
    120: reg_1216 <= imem04_in[15:12];
    endcase
  end

  // REG#1217の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1217 <= op1_01_out;
    endcase
  end

  // REG#1218の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1218 <= op1_04_out;
    endcase
  end

  // REG#1219の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1219 <= op1_06_out;
    endcase
  end

  // REG#1220の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1220 <= op1_08_out;
    endcase
  end

  // REG#1221の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1221 <= op1_09_out;
    endcase
  end

  // REG#1222の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1222 <= op1_10_out;
    endcase
  end

  // REG#1223の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1223 <= op1_13_out;
    88: reg_1223 <= op1_13_out;
    endcase
  end

  // REG#1224の入力
  always @ ( posedge clock ) begin
    case ( state )
    55: reg_1224 <= op1_15_out;
    endcase
  end

  // REG#1225の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1225 <= imem06_in[15:12];
    endcase
  end

  // REG#1226の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1226 <= imem03_in[15:12];
    endcase
  end

  // REG#1227の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1227 <= imem00_in[3:0];
    endcase
  end

  // REG#1228の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1228 <= imem06_in[11:8];
    endcase
  end

  // REG#1229の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1229 <= imem00_in[15:12];
    endcase
  end

  // REG#1230の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1230 <= imem00_in[11:8];
    endcase
  end

  // REG#1231の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1231 <= imem03_in[7:4];
    endcase
  end

  // REG#1232の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1232 <= op1_08_out;
    62: reg_1232 <= op1_08_out;
    endcase
  end

  // REG#1233の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1233 <= imem03_in[11:8];
    71: reg_1233 <= imem04_in[15:12];
    84: reg_1233 <= imem04_in[15:12];
    endcase
  end

  // REG#1234の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1234 <= op1_11_out;
    73: reg_1234 <= op2_02_out;
    81: reg_1234 <= op2_02_out;
    118: reg_1234 <= op2_02_out;
    endcase
  end

  // REG#1235の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1235 <= op1_00_out;
    78: reg_1235 <= imem02_in[3:0];
    endcase
  end

  // REG#1236の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1236 <= op1_01_out;
    77: reg_1236 <= op1_01_out;
    82: reg_1236 <= op1_01_out;
    84: reg_1236 <= op1_01_out;
    endcase
  end

  // REG#1237の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1237 <= op1_02_out;
    78: reg_1237 <= imem04_in[7:4];
    endcase
  end

  // REG#1238の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1238 <= op1_09_out;
    82: reg_1238 <= op1_09_out;
    endcase
  end

  // REG#1239の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1239 <= op1_12_out;
    endcase
  end

  // REG#1240の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1240 <= op1_14_out;
    endcase
  end

  // REG#1241の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1241 <= imem00_in[15:12];
    90: reg_1241 <= imem00_in[15:12];
    endcase
  end

  // REG#1242の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1242 <= imem00_in[11:8];
    91: reg_1242 <= imem00_in[11:8];
    111: reg_1242 <= imem00_in[11:8];
    123: reg_1242 <= imem00_in[11:8];
    endcase
  end

  // REG#1243の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1243 <= imem00_in[3:0];
    89: reg_1243 <= imem00_in[3:0];
    107: reg_1243 <= imem00_in[3:0];
    122: reg_1243 <= imem00_in[3:0];
    endcase
  end

  // REG#1244の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1244 <= imem00_in[7:4];
    90: reg_1244 <= imem00_in[7:4];
    103: reg_1244 <= imem00_in[7:4];
    106: reg_1244 <= imem00_in[7:4];
    114: reg_1244 <= imem00_in[7:4];
    117: reg_1244 <= imem00_in[7:4];
    122: reg_1244 <= imem00_in[7:4];
    endcase
  end

  // REG#1245の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1245 <= op1_03_out;
    endcase
  end

  // REG#1246の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1246 <= op1_04_out;
    endcase
  end

  // REG#1247の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1247 <= op1_05_out;
    endcase
  end

  // REG#1248の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1248 <= op1_06_out;
    endcase
  end

  // REG#1249の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1249 <= op1_07_out;
    endcase
  end

  // REG#1250の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1250 <= op1_10_out;
    endcase
  end

  // REG#1251の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1251 <= op1_13_out;
    endcase
  end

  // REG#1252の入力
  always @ ( posedge clock ) begin
    case ( state )
    56: reg_1252 <= op1_15_out;
    endcase
  end

  // REG#1253の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1253 <= imem01_in[7:4];
    110: reg_1253 <= imem01_in[7:4];
    116: reg_1253 <= imem01_in[7:4];
    120: reg_1253 <= imem01_in[7:4];
    endcase
  end

  // REG#1254の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1254 <= imem01_in[11:8];
    119: reg_1254 <= imem01_in[11:8];
    endcase
  end

  // REG#1255の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1255 <= imem01_in[3:0];
    110: reg_1255 <= imem01_in[3:0];
    117: reg_1255 <= imem01_in[3:0];
    126: reg_1255 <= imem01_in[3:0];
    endcase
  end

  // REG#1256の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1256 <= imem01_in[15:12];
    endcase
  end

  // REG#1257の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1257 <= imem04_in[3:0];
    endcase
  end

  // REG#1258の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1258 <= imem04_in[7:4];
    endcase
  end

  // REG#1259の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1259 <= imem05_in[15:12];
    90: reg_1259 <= imem05_in[15:12];
    107: reg_1259 <= imem05_in[15:12];
    121: reg_1259 <= imem05_in[15:12];
    127: reg_1259 <= imem05_in[15:12];
    endcase
  end

  // REG#1260の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1260 <= imem02_in[15:12];
    89: reg_1260 <= imem02_in[15:12];
    110: reg_1260 <= imem02_in[15:12];
    121: reg_1260 <= imem02_in[15:12];
    125: reg_1260 <= imem02_in[15:12];
    endcase
  end

  // REG#1261の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1261 <= op1_06_out;
    endcase
  end

  // REG#1262の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1262 <= op1_07_out;
    endcase
  end

  // REG#1263の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1263 <= op1_08_out;
    endcase
  end

  // REG#1264の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1264 <= op1_09_out;
    endcase
  end

  // REG#1265の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1265 <= op1_10_out;
    endcase
  end

  // REG#1266の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1266 <= op1_11_out;
    endcase
  end

  // REG#1267の入力
  always @ ( posedge clock ) begin
    case ( state )
    57: reg_1267 <= op1_14_out;
    endcase
  end

  // REG#1268の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1268 <= imem05_in[11:8];
    88: reg_1268 <= imem05_in[11:8];
    92: reg_1268 <= imem05_in[11:8];
    endcase
  end

  // REG#1269の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1269 <= imem05_in[15:12];
    endcase
  end

  // REG#1270の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1270 <= op1_01_out;
    endcase
  end

  // REG#1271の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1271 <= op1_08_out;
    endcase
  end

  // REG#1272の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1272 <= op1_09_out;
    endcase
  end

  // REG#1273の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1273 <= op1_10_out;
    endcase
  end

  // REG#1274の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1274 <= op1_11_out;
    endcase
  end

  // REG#1275の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1275 <= op1_12_out;
    endcase
  end

  // REG#1276の入力
  always @ ( posedge clock ) begin
    case ( state )
    58: reg_1276 <= op1_15_out;
    endcase
  end

  // REG#1277の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1277 <= imem00_in[11:8];
    endcase
  end

  // REG#1278の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1278 <= imem00_in[7:4];
    endcase
  end

  // REG#1279の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1279 <= imem00_in[15:12];
    endcase
  end

  // REG#1280の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1280 <= imem03_in[11:8];
    endcase
  end

  // REG#1281の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1281 <= imem00_in[3:0];
    endcase
  end

  // REG#1282の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1282 <= imem03_in[3:0];
    endcase
  end

  // REG#1283の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1283 <= op1_08_out;
    endcase
  end

  // REG#1284の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1284 <= op1_09_out;
    endcase
  end

  // REG#1285の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1285 <= op1_10_out;
    endcase
  end

  // REG#1286の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1286 <= op1_11_out;
    endcase
  end

  // REG#1287の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1287 <= op1_12_out;
    endcase
  end

  // REG#1288の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1288 <= op1_13_out;
    82: reg_1288 <= op1_13_out;
    84: reg_1288 <= op1_13_out;
    endcase
  end

  // REG#1289の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1289 <= op1_14_out;
    endcase
  end

  // REG#1290の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1290 <= imem01_in[3:0];
    89: reg_1290 <= imem01_in[3:0];
    93: reg_1290 <= imem01_in[3:0];
    95: reg_1290 <= imem01_in[3:0];
    endcase
  end

  // REG#1291の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1291 <= imem01_in[15:12];
    89: reg_1291 <= imem01_in[15:12];
    94: reg_1291 <= imem01_in[15:12];
    endcase
  end

  // REG#1292の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1292 <= op1_01_out;
    endcase
  end

  // REG#1293の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1293 <= op1_02_out;
    endcase
  end

  // REG#1294の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1294 <= op1_03_out;
    endcase
  end

  // REG#1295の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1295 <= op1_06_out;
    endcase
  end

  // REG#1296の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1296 <= op1_07_out;
    endcase
  end

  // REG#1297の入力
  always @ ( posedge clock ) begin
    case ( state )
    59: reg_1297 <= op1_15_out;
    endcase
  end

  // REG#1298の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1298 <= imem05_in[11:8];
    104: reg_1298 <= imem05_in[11:8];
    111: reg_1298 <= imem05_in[11:8];
    113: reg_1298 <= imem05_in[11:8];
    endcase
  end

  // REG#1299の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1299 <= imem05_in[3:0];
    118: reg_1299 <= imem05_in[3:0];
    endcase
  end

  // REG#1300の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1300 <= imem03_in[3:0];
    121: reg_1300 <= imem03_in[3:0];
    endcase
  end

  // REG#1301の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1301 <= imem03_in[15:12];
    122: reg_1301 <= imem03_in[15:12];
    endcase
  end

  // REG#1302の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1302 <= imem06_in[3:0];
    endcase
  end

  // REG#1303の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1303 <= imem06_in[7:4];
    endcase
  end

  // REG#1304の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1304 <= op1_09_out;
    endcase
  end

  // REG#1305の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1305 <= op1_14_out;
    endcase
  end

  // REG#1306の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1306 <= op1_15_out;
    endcase
  end

  // REG#1307の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1307 <= op1_01_out;
    endcase
  end

  // REG#1308の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1308 <= op1_10_out;
    endcase
  end

  // REG#1309の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1309 <= op1_11_out;
    endcase
  end

  // REG#1310の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1310 <= op1_12_out;
    endcase
  end

  // REG#1311の入力
  always @ ( posedge clock ) begin
    case ( state )
    60: reg_1311 <= op1_13_out;
    endcase
  end

  // REG#1312の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1312 <= imem04_in[3:0];
    97: reg_1312 <= imem04_in[3:0];
    104: reg_1312 <= imem04_in[3:0];
    108: reg_1312 <= imem04_in[3:0];
    endcase
  end

  // REG#1313の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1313 <= imem03_in[15:12];
    endcase
  end

  // REG#1314の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1314 <= imem03_in[11:8];
    endcase
  end

  // REG#1315の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1315 <= imem07_in[3:0];
    endcase
  end

  // REG#1316の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1316 <= op1_08_out;
    endcase
  end

  // REG#1317の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1317 <= op1_09_out;
    endcase
  end

  // REG#1318の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1318 <= op1_10_out;
    endcase
  end

  // REG#1319の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1319 <= op1_12_out;
    endcase
  end

  // REG#1320の入力
  always @ ( posedge clock ) begin
    case ( state )
    61: reg_1320 <= op1_13_out;
    endcase
  end

  // REG#1321の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1321 <= imem00_in[3:0];
    endcase
  end

  // REG#1322の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1322 <= imem00_in[15:12];
    endcase
  end

  // REG#1323の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1323 <= imem06_in[7:4];
    endcase
  end

  // REG#1324の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1324 <= imem00_in[11:8];
    endcase
  end

  // REG#1325の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1325 <= imem03_in[15:12];
    85: reg_1325 <= imem03_in[15:12];
    endcase
  end

  // REG#1326の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1326 <= imem06_in[7:4];
    85: reg_1326 <= imem06_in[7:4];
    endcase
  end

  // REG#1327の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1327 <= op1_01_out;
    83: reg_1327 <= op1_01_out;
    endcase
  end

  // REG#1328の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1328 <= op1_03_out;
    87: reg_1328 <= op1_03_out;
    endcase
  end

  // REG#1329の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1329 <= op1_04_out;
    endcase
  end

  // REG#1330の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1330 <= op1_05_out;
    endcase
  end

  // REG#1331の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1331 <= op1_06_out;
    endcase
  end

  // REG#1332の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1332 <= op1_07_out;
    84: reg_1332 <= op1_07_out;
    87: reg_1332 <= op1_07_out;
    endcase
  end

  // REG#1333の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1333 <= op1_15_out;
    endcase
  end

  // REG#1334の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1334 <= imem06_in[11:8];
    87: reg_1334 <= imem06_in[11:8];
    endcase
  end

  // REG#1335の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1335 <= op1_09_out;
    endcase
  end

  // REG#1336の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1336 <= op1_10_out;
    endcase
  end

  // REG#1337の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1337 <= op1_11_out;
    endcase
  end

  // REG#1338の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1338 <= imem04_in[15:12];
    110: reg_1338 <= imem04_in[15:12];
    124: reg_1338 <= imem04_in[15:12];
    endcase
  end

  // REG#1339の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1339 <= imem04_in[3:0];
    110: reg_1339 <= imem04_in[3:0];
    117: reg_1339 <= imem04_in[3:0];
    120: reg_1339 <= imem04_in[3:0];
    endcase
  end

  // REG#1340の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1340 <= imem04_in[7:4];
    98: reg_1340 <= imem04_in[7:4];
    101: reg_1340 <= imem04_in[7:4];
    108: reg_1340 <= imem04_in[7:4];
    endcase
  end

  // REG#1341の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1341 <= op1_12_out;
    endcase
  end

  // REG#1342の入力
  always @ ( posedge clock ) begin
    case ( state )
    62: reg_1342 <= op1_13_out;
    endcase
  end

  // REG#1343の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1343 <= imem02_in[11:8];
    endcase
  end

  // REG#1344の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1344 <= imem02_in[3:0];
    106: reg_1344 <= imem02_in[3:0];
    113: reg_1344 <= imem02_in[3:0];
    endcase
  end

  // REG#1345の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1345 <= imem07_in[11:8];
    endcase
  end

  // REG#1346の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1346 <= imem05_in[15:12];
    endcase
  end

  // REG#1347の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1347 <= imem07_in[7:4];
    endcase
  end

  // REG#1348の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1348 <= imem05_in[7:4];
    endcase
  end

  // REG#1349の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1349 <= imem07_in[15:12];
    endcase
  end

  // REG#1350の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1350 <= imem07_in[3:0];
    endcase
  end

  // REG#1351の入力
  always @ ( posedge clock ) begin
    case ( state )
    64: reg_1351 <= imem07_in[3:0];
    91: reg_1351 <= imem07_in[3:0];
    109: reg_1351 <= imem07_in[3:0];
    118: reg_1351 <= imem07_in[3:0];
    endcase
  end

  // REG#1352の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1352 <= op1_01_out;
    87: reg_1352 <= op1_01_out;
    endcase
  end

  // REG#1353の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1353 <= op1_04_out;
    endcase
  end

  // REG#1354の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1354 <= op1_05_out;
    endcase
  end

  // REG#1355の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1355 <= op1_06_out;
    endcase
  end

  // REG#1356の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1356 <= op1_08_out;
    endcase
  end

  // REG#1357の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1357 <= op1_00_out;
    endcase
  end

  // REG#1358の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1358 <= op1_03_out;
    endcase
  end

  // REG#1359の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1359 <= op1_07_out;
    endcase
  end

  // REG#1360の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1360 <= op1_09_out;
    endcase
  end

  // REG#1361の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1361 <= op1_10_out;
    endcase
  end

  // REG#1362の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1362 <= op1_11_out;
    endcase
  end

  // REG#1363の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1363 <= op1_12_out;
    endcase
  end

  // REG#1364の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1364 <= op1_13_out;
    endcase
  end

  // REG#1365の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1365 <= op1_14_out;
    endcase
  end

  // REG#1366の入力
  always @ ( posedge clock ) begin
    case ( state )
    63: reg_1366 <= op1_15_out;
    endcase
  end

  // REG#1367の入力
  always @ ( posedge clock ) begin
    case ( state )
    64: reg_1367 <= imem04_in[11:8];
    127: reg_1367 <= imem04_in[11:8];
    endcase
  end

  // REG#1368の入力
  always @ ( posedge clock ) begin
    case ( state )
    64: reg_1368 <= imem04_in[7:4];
    endcase
  end

  // REG#1369の入力
  always @ ( posedge clock ) begin
    case ( state )
    64: reg_1369 <= imem04_in[3:0];
    126: reg_1369 <= imem04_in[3:0];
    endcase
  end

  // REG#1370の入力
  always @ ( posedge clock ) begin
    case ( state )
    64: reg_1370 <= op1_05_out;
    endcase
  end

  // REG#1371の入力
  always @ ( posedge clock ) begin
    case ( state )
    64: reg_1371 <= op1_15_out;
    endcase
  end

  // REG#1372の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1372 <= imem04_in[11:8];
    116: reg_1372 <= imem04_in[11:8];
    118: reg_1372 <= imem04_in[11:8];
    122: reg_1372 <= imem04_in[11:8];
    124: reg_1372 <= imem04_in[11:8];
    endcase
  end

  // REG#1373の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1373 <= imem05_in[15:12];
    endcase
  end

  // REG#1374の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1374 <= op1_02_out;
    87: reg_1374 <= op1_02_out;
    endcase
  end

  // REG#1375の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1375 <= op1_03_out;
    endcase
  end

  // REG#1376の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1376 <= op1_05_out;
    endcase
  end

  // REG#1377の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1377 <= op1_09_out;
    endcase
  end

  // REG#1378の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1378 <= op1_10_out;
    endcase
  end

  // REG#1379の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1379 <= op1_11_out;
    endcase
  end

  // REG#1380の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1380 <= op1_12_out;
    endcase
  end

  // REG#1381の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1381 <= op1_13_out;
    endcase
  end

  // REG#1382の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1382 <= op1_14_out;
    endcase
  end

  // REG#1383の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1383 <= imem04_in[11:8];
    94: reg_1383 <= imem04_in[11:8];
    119: reg_1383 <= imem04_in[11:8];
    125: reg_1383 <= imem04_in[11:8];
    endcase
  end

  // REG#1384の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1384 <= imem04_in[3:0];
    124: reg_1384 <= imem04_in[3:0];
    endcase
  end

  // REG#1385の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1385 <= op1_00_out;
    endcase
  end

  // REG#1386の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1386 <= op1_01_out;
    endcase
  end

  // REG#1387の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1387 <= op1_04_out;
    endcase
  end

  // REG#1388の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1388 <= op1_06_out;
    endcase
  end

  // REG#1389の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1389 <= op1_07_out;
    endcase
  end

  // REG#1390の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1390 <= op1_08_out;
    endcase
  end

  // REG#1391の入力
  always @ ( posedge clock ) begin
    case ( state )
    65: reg_1391 <= op1_15_out;
    endcase
  end

  // REG#1392の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1392 <= imem02_in[15:12];
    106: reg_1392 <= imem02_in[15:12];
    endcase
  end

  // REG#1393の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1393 <= imem00_in[15:12];
    endcase
  end

  // REG#1394の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1394 <= op1_06_out;
    endcase
  end

  // REG#1395の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1395 <= op1_07_out;
    endcase
  end

  // REG#1396の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1396 <= op1_08_out;
    endcase
  end

  // REG#1397の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1397 <= op1_09_out;
    endcase
  end

  // REG#1398の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1398 <= op1_10_out;
    endcase
  end

  // REG#1399の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1399 <= op1_12_out;
    endcase
  end

  // REG#1400の入力
  always @ ( posedge clock ) begin
    case ( state )
    66: reg_1400 <= op1_15_out;
    endcase
  end

  // REG#1401の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1401 <= imem05_in[11:8];
    endcase
  end

  // REG#1402の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1402 <= imem05_in[7:4];
    endcase
  end

  // REG#1403の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1403 <= imem05_in[3:0];
    endcase
  end

  // REG#1404の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1404 <= imem05_in[15:12];
    endcase
  end

  // REG#1405の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1405 <= imem00_in[15:12];
    endcase
  end

  // REG#1406の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1406 <= imem00_in[7:4];
    endcase
  end

  // REG#1407の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1407 <= op1_09_out;
    endcase
  end

  // REG#1408の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1408 <= op1_10_out;
    endcase
  end

  // REG#1409の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1409 <= op1_11_out;
    endcase
  end

  // REG#1410の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1410 <= op1_12_out;
    endcase
  end

  // REG#1411の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1411 <= op1_13_out;
    endcase
  end

  // REG#1412の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1412 <= op1_14_out;
    endcase
  end

  // REG#1413の入力
  always @ ( posedge clock ) begin
    case ( state )
    67: reg_1413 <= op1_15_out;
    endcase
  end

  // REG#1414の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1414 <= imem07_in[3:0];
    endcase
  end

  // REG#1415の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1415 <= imem07_in[15:12];
    115: reg_1415 <= imem07_in[15:12];
    endcase
  end

  // REG#1416の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1416 <= imem07_in[11:8];
    endcase
  end

  // REG#1417の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1417 <= imem00_in[3:0];
    endcase
  end

  // REG#1418の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1418 <= imem00_in[11:8];
    endcase
  end

  // REG#1419の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1419 <= imem04_in[3:0];
    endcase
  end

  // REG#1420の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1420 <= imem06_in[15:12];
    endcase
  end

  // REG#1421の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1421 <= op1_09_out;
    endcase
  end

  // REG#1422の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1422 <= op1_10_out;
    78: reg_1422 <= op1_10_out;
    80: reg_1422 <= op1_10_out;
    endcase
  end

  // REG#1423の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1423 <= op1_13_out;
    86: reg_1423 <= op1_13_out;
    endcase
  end

  // REG#1424の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1424 <= op1_15_out;
    endcase
  end

  // REG#1425の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1425 <= imem03_in[11:8];
    81: reg_1425 <= imem03_in[11:8];
    endcase
  end

  // REG#1426の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1426 <= imem06_in[7:4];
    endcase
  end

  // REG#1427の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1427 <= op1_11_out;
    endcase
  end

  // REG#1428の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1428 <= op1_03_out;
    endcase
  end

  // REG#1429の入力
  always @ ( posedge clock ) begin
    case ( state )
    68: reg_1429 <= op1_14_out;
    endcase
  end

  // REG#1430の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1430 <= imem05_in[3:0];
    endcase
  end

  // REG#1431の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1431 <= imem05_in[11:8];
    115: reg_1431 <= imem05_in[11:8];
    endcase
  end

  // REG#1432の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1432 <= imem00_in[7:4];
    endcase
  end

  // REG#1433の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1433 <= imem02_in[15:12];
    endcase
  end

  // REG#1434の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1434 <= op1_12_out;
    77: reg_1434 <= op1_12_out;
    endcase
  end

  // REG#1435の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1435 <= imem06_in[15:12];
    78: reg_1435 <= imem06_in[15:12];
    91: reg_1435 <= imem06_in[15:12];
    100: reg_1435 <= imem06_in[15:12];
    104: reg_1435 <= imem06_in[15:12];
    118: reg_1435 <= imem06_in[15:12];
    endcase
  end

  // REG#1436の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1436 <= imem06_in[7:4];
    81: reg_1436 <= imem06_in[7:4];
    endcase
  end

  // REG#1437の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1437 <= imem06_in[11:8];
    78: reg_1437 <= imem06_in[11:8];
    88: reg_1437 <= imem06_in[11:8];
    91: reg_1437 <= imem06_in[11:8];
    95: reg_1437 <= imem06_in[11:8];
    endcase
  end

  // REG#1438の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1438 <= op1_15_out;
    endcase
  end

  // REG#1439の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1439 <= imem07_in[7:4];
    84: reg_1439 <= imem07_in[7:4];
    118: reg_1439 <= imem07_in[7:4];
    endcase
  end

  // REG#1440の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1440 <= imem07_in[15:12];
    83: reg_1440 <= imem07_in[15:12];
    87: reg_1440 <= imem07_in[15:12];
    endcase
  end

  // REG#1441の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1441 <= imem07_in[3:0];
    endcase
  end

  // REG#1442の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1442 <= op1_02_out;
    endcase
  end

  // REG#1443の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1443 <= op1_03_out;
    endcase
  end

  // REG#1444の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1444 <= op1_08_out;
    endcase
  end

  // REG#1445の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1445 <= op1_09_out;
    endcase
  end

  // REG#1446の入力
  always @ ( posedge clock ) begin
    case ( state )
    69: reg_1446 <= op1_13_out;
    endcase
  end

  // REG#1447の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1447 <= imem03_in[7:4];
    108: reg_1447 <= imem03_in[7:4];
    111: reg_1447 <= imem03_in[7:4];
    endcase
  end

  // REG#1448の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1448 <= imem03_in[15:12];
    104: reg_1448 <= imem03_in[15:12];
    115: reg_1448 <= imem03_in[15:12];
    118: reg_1448 <= imem03_in[15:12];
    endcase
  end

  // REG#1449の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1449 <= imem03_in[3:0];
    endcase
  end

  // REG#1450の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1450 <= imem02_in[11:8];
    endcase
  end

  // REG#1451の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1451 <= imem02_in[7:4];
    endcase
  end

  // REG#1452の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1452 <= imem01_in[3:0];
    endcase
  end

  // REG#1453の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1453 <= imem00_in[11:8];
    endcase
  end

  // REG#1454の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1454 <= imem00_in[7:4];
    endcase
  end

  // REG#1455の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1455 <= imem02_in[15:12];
    endcase
  end

  // REG#1456の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1456 <= imem01_in[15:12];
    endcase
  end

  // REG#1457の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1457 <= imem01_in[7:4];
    endcase
  end

  // REG#1458の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1458 <= imem02_in[3:0];
    endcase
  end

  // REG#1459の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1459 <= imem00_in[15:12];
    endcase
  end

  // REG#1460の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1460 <= op1_09_out;
    endcase
  end

  // REG#1461の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1461 <= op1_10_out;
    endcase
  end

  // REG#1462の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1462 <= op1_11_out;
    endcase
  end

  // REG#1463の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1463 <= op1_12_out;
    endcase
  end

  // REG#1464の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1464 <= op1_13_out;
    endcase
  end

  // REG#1465の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1465 <= op1_14_out;
    endcase
  end

  // REG#1466の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1466 <= op1_15_out;
    endcase
  end

  // REG#1467の入力
  always @ ( posedge clock ) begin
    case ( state )
    71: reg_1467 <= imem06_in[11:8];
    85: reg_1467 <= imem06_in[11:8];
    endcase
  end

  // REG#1468の入力
  always @ ( posedge clock ) begin
    case ( state )
    71: reg_1468 <= imem06_in[3:0];
    84: reg_1468 <= imem06_in[3:0];
    90: reg_1468 <= imem06_in[3:0];
    102: reg_1468 <= imem06_in[3:0];
    104: reg_1468 <= imem06_in[3:0];
    endcase
  end

  // REG#1469の入力
  always @ ( posedge clock ) begin
    case ( state )
    71: reg_1469 <= imem00_in[7:4];
    95: reg_1469 <= imem00_in[7:4];
    119: reg_1469 <= imem00_in[7:4];
    121: reg_1469 <= imem00_in[7:4];
    endcase
  end

  // REG#1470の入力
  always @ ( posedge clock ) begin
    case ( state )
    71: reg_1470 <= imem00_in[11:8];
    92: reg_1470 <= imem00_in[11:8];
    117: reg_1470 <= imem00_in[11:8];
    endcase
  end

  // REG#1471の入力
  always @ ( posedge clock ) begin
    case ( state )
    71: reg_1471 <= imem00_in[3:0];
    endcase
  end

  // REG#1472の入力
  always @ ( posedge clock ) begin
    case ( state )
    70: reg_1472 <= op1_04_out;
    endcase
  end

  // REG#1473の入力
  always @ ( posedge clock ) begin
    case ( state )
    71: reg_1473 <= imem01_in[3:0];
    endcase
  end

  // REG#1474の入力
  always @ ( posedge clock ) begin
    case ( state )
    71: reg_1474 <= imem01_in[15:12];
    endcase
  end

  // REG#1475の入力
  always @ ( posedge clock ) begin
    case ( state )
    71: reg_1475 <= imem01_in[11:8];
    endcase
  end

  // REG#1476の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_1476 <= op1_05_out;
    endcase
  end

  // REG#1477の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_1477 <= op1_07_out;
    endcase
  end

  // REG#1478の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_1478 <= op1_08_out;
    endcase
  end

  // REG#1479の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_1479 <= op1_09_out;
    endcase
  end

  // REG#1480の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_1480 <= op1_10_out;
    endcase
  end

  // REG#1481の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_1481 <= op1_14_out;
    endcase
  end

  // REG#1482の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_1482 <= op1_15_out;
    endcase
  end

  // REG#1483の入力
  always @ ( posedge clock ) begin
    case ( state )
    72: reg_1483 <= op1_01_out;
    endcase
  end

  // REG#1484の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1484 <= imem05_in[11:8];
    endcase
  end

  // REG#1485の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1485 <= imem05_in[7:4];
    107: reg_1485 <= imem05_in[7:4];
    121: reg_1485 <= imem05_in[7:4];
    endcase
  end

  // REG#1486の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1486 <= imem05_in[3:0];
    endcase
  end

  // REG#1487の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1487 <= imem00_in[11:8];
    endcase
  end

  // REG#1488の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1488 <= imem04_in[3:0];
    endcase
  end

  // REG#1489の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1489 <= imem00_in[7:4];
    endcase
  end

  // REG#1490の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1490 <= imem00_in[3:0];
    endcase
  end

  // REG#1491の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1491 <= imem00_in[15:12];
    endcase
  end

  // REG#1492の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1492 <= imem02_in[3:0];
    84: reg_1492 <= imem02_in[3:0];
    endcase
  end

  // REG#1493の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1493 <= imem02_in[11:8];
    90: reg_1493 <= imem02_in[11:8];
    endcase
  end

  // REG#1494の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1494 <= imem03_in[7:4];
    93: reg_1494 <= imem03_in[7:4];
    endcase
  end

  // REG#1495の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1495 <= imem03_in[11:8];
    93: reg_1495 <= imem03_in[11:8];
    endcase
  end

  // REG#1496の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1496 <= op1_01_out;
    endcase
  end

  // REG#1497の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1497 <= op1_06_out;
    endcase
  end

  // REG#1498の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1498 <= op1_07_out;
    endcase
  end

  // REG#1499の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1499 <= op1_08_out;
    endcase
  end

  // REG#1500の入力
  always @ ( posedge clock ) begin
    case ( state )
    73: reg_1500 <= op1_13_out;
    endcase
  end

  // REG#1501の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1501 <= imem06_in[7:4];
    endcase
  end

  // REG#1502の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1502 <= imem04_in[7:4];
    endcase
  end

  // REG#1503の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1503 <= imem04_in[15:12];
    endcase
  end

  // REG#1504の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1504 <= imem06_in[11:8];
    endcase
  end

  // REG#1505の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1505 <= imem06_in[3:0];
    endcase
  end

  // REG#1506の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1506 <= op2_04_out;
    87: reg_1506 <= op2_04_out;
    endcase
  end

  // REG#1507の入力
  always @ ( posedge clock ) begin
    case ( state )
    74: reg_1507 <= op2_05_out;
    87: reg_1507 <= op2_05_out;
    endcase
  end

  // REG#1508の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1508 <= imem06_in[15:12];
    92: reg_1508 <= imem06_in[15:12];
    101: reg_1508 <= imem06_in[15:12];
    endcase
  end

  // REG#1509の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1509 <= imem06_in[7:4];
    endcase
  end

  // REG#1510の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1510 <= imem00_in[15:12];
    endcase
  end

  // REG#1511の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1511 <= imem01_in[11:8];
    96: reg_1511 <= imem01_in[11:8];
    120: reg_1511 <= imem01_in[11:8];
    endcase
  end

  // REG#1512の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1512 <= imem01_in[7:4];
    100: reg_1512 <= imem01_in[7:4];
    105: reg_1512 <= imem01_in[7:4];
    117: reg_1512 <= imem01_in[7:4];
    endcase
  end

  // REG#1513の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1513 <= imem01_in[15:12];
    96: reg_1513 <= imem01_in[15:12];
    endcase
  end

  // REG#1514の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1514 <= imem05_in[11:8];
    endcase
  end

  // REG#1515の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1515 <= imem02_in[3:0];
    endcase
  end

  // REG#1516の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1516 <= imem03_in[7:4];
    endcase
  end

  // REG#1517の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1517 <= imem03_in[15:12];
    endcase
  end

  // REG#1518の入力
  always @ ( posedge clock ) begin
    case ( state )
    75: reg_1518 <= imem03_in[11:8];
    endcase
  end
endmodule
