module affine3(
  input clock,
  input reset,
  input start,
  output busy,
  output [5:0] imem00_bank,
  output imem00_rd,
  input [8:0] imem00_in,
  output [5:0] imem01_bank,
  output imem01_rd,
  input [8:0] imem01_in,
  output [5:0] imem02_bank,
  output imem02_rd,
  input [8:0] imem02_in,
  output [5:0] imem03_bank,
  output imem03_rd,
  input [8:0] imem03_in,
  output [5:0] imem04_bank,
  output imem04_rd,
  input [8:0] imem04_in,
  output omem00_wr,
  output [14:0] omem00_out);


  // 0 番目の OP1
  reg [8:0] op1_00_in00;
  reg       op1_00_inv00;
  reg [8:0] op1_00_in01;
  reg       op1_00_inv01;
  reg [8:0] op1_00_in02;
  reg       op1_00_inv02;
  reg [8:0] op1_00_in03;
  reg       op1_00_inv03;
  reg [8:0] op1_00_in04;
  reg       op1_00_inv04;
  reg [8:0] op1_00_in05;
  reg       op1_00_inv05;
  reg [8:0] op1_00_in06;
  reg       op1_00_inv06;
  reg [8:0] op1_00_in07;
  reg       op1_00_inv07;
  reg [8:0] op1_00_in08;
  reg       op1_00_inv08;
  reg [8:0] op1_00_in09;
  reg       op1_00_inv09;
  reg [8:0] op1_00_in10;
  reg       op1_00_inv10;
  reg [8:0] op1_00_in11;
  reg       op1_00_inv11;
  reg [8:0] op1_00_in12;
  reg       op1_00_inv12;
  reg [8:0] op1_00_in13;
  reg       op1_00_inv13;
  reg [8:0] op1_00_in14;
  reg       op1_00_inv14;
  reg [8:0] op1_00_in15;
  reg       op1_00_inv15;
  reg [8:0] op1_00_in16;
  reg       op1_00_inv16;
  reg [8:0] op1_00_in17;
  reg       op1_00_inv17;
  reg [8:0] op1_00_in18;
  reg       op1_00_inv18;
  reg [8:0] op1_00_in19;
  reg       op1_00_inv19;
  reg [8:0] op1_00_in20;
  reg       op1_00_inv20;
  reg [8:0] op1_00_in21;
  reg       op1_00_inv21;
  reg [8:0] op1_00_in22;
  reg       op1_00_inv22;
  reg [8:0] op1_00_in23;
  reg       op1_00_inv23;
  reg [8:0] op1_00_in24;
  reg       op1_00_inv24;
  reg [8:0] op1_00_in25;
  reg       op1_00_inv25;
  reg [8:0] op1_00_in26;
  reg       op1_00_inv26;
  reg [8:0] op1_00_in27;
  reg       op1_00_inv27;
  reg [8:0] op1_00_in28;
  reg       op1_00_inv28;
  reg [8:0] op1_00_in29;
  reg       op1_00_inv29;
  reg [8:0] op1_00_in30;
  reg       op1_00_inv30;
  reg [8:0] op1_00_in31;
  reg       op1_00_inv31;
  wire [13:0] op1_00_out;
  op1 op1_00(
    .data0_in(op1_00_in00),
    .inv0_in(op1_00_inv00),
    .data1_in(op1_00_in01),
    .inv1_in(op1_00_inv01),
    .data2_in(op1_00_in02),
    .inv2_in(op1_00_inv02),
    .data3_in(op1_00_in03),
    .inv3_in(op1_00_inv03),
    .data4_in(op1_00_in04),
    .inv4_in(op1_00_inv04),
    .data5_in(op1_00_in05),
    .inv5_in(op1_00_inv05),
    .data6_in(op1_00_in06),
    .inv6_in(op1_00_inv06),
    .data7_in(op1_00_in07),
    .inv7_in(op1_00_inv07),
    .data8_in(op1_00_in08),
    .inv8_in(op1_00_inv08),
    .data9_in(op1_00_in09),
    .inv9_in(op1_00_inv09),
    .data10_in(op1_00_in10),
    .inv10_in(op1_00_inv10),
    .data11_in(op1_00_in11),
    .inv11_in(op1_00_inv11),
    .data12_in(op1_00_in12),
    .inv12_in(op1_00_inv12),
    .data13_in(op1_00_in13),
    .inv13_in(op1_00_inv13),
    .data14_in(op1_00_in14),
    .inv14_in(op1_00_inv14),
    .data15_in(op1_00_in15),
    .inv15_in(op1_00_inv15),
    .data16_in(op1_00_in16),
    .inv16_in(op1_00_inv16),
    .data17_in(op1_00_in17),
    .inv17_in(op1_00_inv17),
    .data18_in(op1_00_in18),
    .inv18_in(op1_00_inv18),
    .data19_in(op1_00_in19),
    .inv19_in(op1_00_inv19),
    .data20_in(op1_00_in20),
    .inv20_in(op1_00_inv20),
    .data21_in(op1_00_in21),
    .inv21_in(op1_00_inv21),
    .data22_in(op1_00_in22),
    .inv22_in(op1_00_inv22),
    .data23_in(op1_00_in23),
    .inv23_in(op1_00_inv23),
    .data24_in(op1_00_in24),
    .inv24_in(op1_00_inv24),
    .data25_in(op1_00_in25),
    .inv25_in(op1_00_inv25),
    .data26_in(op1_00_in26),
    .inv26_in(op1_00_inv26),
    .data27_in(op1_00_in27),
    .inv27_in(op1_00_inv27),
    .data28_in(op1_00_in28),
    .inv28_in(op1_00_inv28),
    .data29_in(op1_00_in29),
    .inv29_in(op1_00_inv29),
    .data30_in(op1_00_in30),
    .inv30_in(op1_00_inv30),
    .data31_in(op1_00_in31),
    .inv31_in(op1_00_inv31),
    .data_out(op1_00_out));

  // 1 番目の OP1
  reg [8:0] op1_01_in00;
  reg       op1_01_inv00;
  reg [8:0] op1_01_in01;
  reg       op1_01_inv01;
  reg [8:0] op1_01_in02;
  reg       op1_01_inv02;
  reg [8:0] op1_01_in03;
  reg       op1_01_inv03;
  reg [8:0] op1_01_in04;
  reg       op1_01_inv04;
  reg [8:0] op1_01_in05;
  reg       op1_01_inv05;
  reg [8:0] op1_01_in06;
  reg       op1_01_inv06;
  reg [8:0] op1_01_in07;
  reg       op1_01_inv07;
  reg [8:0] op1_01_in08;
  reg       op1_01_inv08;
  reg [8:0] op1_01_in09;
  reg       op1_01_inv09;
  reg [8:0] op1_01_in10;
  reg       op1_01_inv10;
  reg [8:0] op1_01_in11;
  reg       op1_01_inv11;
  reg [8:0] op1_01_in12;
  reg       op1_01_inv12;
  reg [8:0] op1_01_in13;
  reg       op1_01_inv13;
  reg [8:0] op1_01_in14;
  reg       op1_01_inv14;
  reg [8:0] op1_01_in15;
  reg       op1_01_inv15;
  reg [8:0] op1_01_in16;
  reg       op1_01_inv16;
  reg [8:0] op1_01_in17;
  reg       op1_01_inv17;
  reg [8:0] op1_01_in18;
  reg       op1_01_inv18;
  reg [8:0] op1_01_in19;
  reg       op1_01_inv19;
  reg [8:0] op1_01_in20;
  reg       op1_01_inv20;
  reg [8:0] op1_01_in21;
  reg       op1_01_inv21;
  reg [8:0] op1_01_in22;
  reg       op1_01_inv22;
  reg [8:0] op1_01_in23;
  reg       op1_01_inv23;
  reg [8:0] op1_01_in24;
  reg       op1_01_inv24;
  reg [8:0] op1_01_in25;
  reg       op1_01_inv25;
  reg [8:0] op1_01_in26;
  reg       op1_01_inv26;
  reg [8:0] op1_01_in27;
  reg       op1_01_inv27;
  reg [8:0] op1_01_in28;
  reg       op1_01_inv28;
  reg [8:0] op1_01_in29;
  reg       op1_01_inv29;
  reg [8:0] op1_01_in30;
  reg       op1_01_inv30;
  reg [8:0] op1_01_in31;
  reg       op1_01_inv31;
  wire [13:0] op1_01_out;
  op1 op1_01(
    .data0_in(op1_01_in00),
    .inv0_in(op1_01_inv00),
    .data1_in(op1_01_in01),
    .inv1_in(op1_01_inv01),
    .data2_in(op1_01_in02),
    .inv2_in(op1_01_inv02),
    .data3_in(op1_01_in03),
    .inv3_in(op1_01_inv03),
    .data4_in(op1_01_in04),
    .inv4_in(op1_01_inv04),
    .data5_in(op1_01_in05),
    .inv5_in(op1_01_inv05),
    .data6_in(op1_01_in06),
    .inv6_in(op1_01_inv06),
    .data7_in(op1_01_in07),
    .inv7_in(op1_01_inv07),
    .data8_in(op1_01_in08),
    .inv8_in(op1_01_inv08),
    .data9_in(op1_01_in09),
    .inv9_in(op1_01_inv09),
    .data10_in(op1_01_in10),
    .inv10_in(op1_01_inv10),
    .data11_in(op1_01_in11),
    .inv11_in(op1_01_inv11),
    .data12_in(op1_01_in12),
    .inv12_in(op1_01_inv12),
    .data13_in(op1_01_in13),
    .inv13_in(op1_01_inv13),
    .data14_in(op1_01_in14),
    .inv14_in(op1_01_inv14),
    .data15_in(op1_01_in15),
    .inv15_in(op1_01_inv15),
    .data16_in(op1_01_in16),
    .inv16_in(op1_01_inv16),
    .data17_in(op1_01_in17),
    .inv17_in(op1_01_inv17),
    .data18_in(op1_01_in18),
    .inv18_in(op1_01_inv18),
    .data19_in(op1_01_in19),
    .inv19_in(op1_01_inv19),
    .data20_in(op1_01_in20),
    .inv20_in(op1_01_inv20),
    .data21_in(op1_01_in21),
    .inv21_in(op1_01_inv21),
    .data22_in(op1_01_in22),
    .inv22_in(op1_01_inv22),
    .data23_in(op1_01_in23),
    .inv23_in(op1_01_inv23),
    .data24_in(op1_01_in24),
    .inv24_in(op1_01_inv24),
    .data25_in(op1_01_in25),
    .inv25_in(op1_01_inv25),
    .data26_in(op1_01_in26),
    .inv26_in(op1_01_inv26),
    .data27_in(op1_01_in27),
    .inv27_in(op1_01_inv27),
    .data28_in(op1_01_in28),
    .inv28_in(op1_01_inv28),
    .data29_in(op1_01_in29),
    .inv29_in(op1_01_inv29),
    .data30_in(op1_01_in30),
    .inv30_in(op1_01_inv30),
    .data31_in(op1_01_in31),
    .inv31_in(op1_01_inv31),
    .data_out(op1_01_out));

  // 0 番目の OP2
  reg [13:0] op2_00_in00;
  reg [13:0] op2_00_in01;
  reg [13:0] op2_00_in02;
  reg [13:0] op2_00_in03;
  reg [13:0] op2_00_in04;
  reg [13:0] op2_00_in05;
  reg [13:0] op2_00_in06;
  reg [13:0] op2_00_in07;
  reg [13:0] op2_00_in08;
  reg [13:0] op2_00_in09;
  reg [13:0] op2_00_in10;
  reg [13:0] op2_00_in11;
  reg [13:0] op2_00_in12;
  reg [13:0] op2_00_in13;
  reg [13:0] op2_00_in14;
  reg [13:0] op2_00_bias;
  wire [14:0] op2_00_out;
  op2 op2_00(
    .data0_in(op2_00_in00),
    .data1_in(op2_00_in01),
    .data2_in(op2_00_in02),
    .data3_in(op2_00_in03),
    .data4_in(op2_00_in04),
    .data5_in(op2_00_in05),
    .data6_in(op2_00_in06),
    .data7_in(op2_00_in07),
    .data8_in(op2_00_in08),
    .data9_in(op2_00_in09),
    .data10_in(op2_00_in10),
    .data11_in(op2_00_in11),
    .data12_in(op2_00_in12),
    .data13_in(op2_00_in13),
    .data14_in(op2_00_in14),
    .data15_in(op2_00_bias),
    .data_out(op2_00_out));

  // 中間レジスタ
  reg [13:0] reg_0000;
  reg [13:0] reg_0001;
  reg [13:0] reg_0002;
  reg [13:0] reg_0003;
  reg [13:0] reg_0004;
  reg [13:0] reg_0005;
  reg [13:0] reg_0006;
  reg [13:0] reg_0007;
  reg [13:0] reg_0008;
  reg [13:0] reg_0009;
  reg [13:0] reg_0010;
  reg [13:0] reg_0011;
  reg [13:0] reg_0012;
  reg [13:0] reg_0013;
  reg [13:0] reg_0014;
  reg [13:0] reg_0015;
  reg [13:0] reg_0016;
  reg [13:0] reg_0017;
  reg [13:0] reg_0018;
  reg [13:0] reg_0019;
  reg [13:0] reg_0020;
  reg [13:0] reg_0021;
  reg [13:0] reg_0022;
  reg [13:0] reg_0023;
  reg [13:0] reg_0024;
  reg [13:0] reg_0025;
  reg [13:0] reg_0026;
  reg [13:0] reg_0027;
  reg [13:0] reg_0028;
  reg [13:0] reg_0029;
  reg [13:0] reg_0030;
  reg [13:0] reg_0031;
  reg [13:0] reg_0032;
  reg [13:0] reg_0033;
  reg [13:0] reg_0034;
  reg [13:0] reg_0035;
  reg [13:0] reg_0036;
  reg [13:0] reg_0037;
  reg [13:0] reg_0038;
  reg [13:0] reg_0039;
  reg [13:0] reg_0040;
  reg [13:0] reg_0041;
  reg [13:0] reg_0042;
  reg [13:0] reg_0043;
  reg [13:0] reg_0044;
  reg [13:0] reg_0045;
  reg [13:0] reg_0046;
  reg [13:0] reg_0047;
  reg [13:0] reg_0048;
  reg [13:0] reg_0049;
  reg [13:0] reg_0050;
  reg [13:0] reg_0051;
  reg [13:0] reg_0052;
  reg [13:0] reg_0053;
  reg [13:0] reg_0054;
  reg [13:0] reg_0055;
  reg [13:0] reg_0056;
  reg [13:0] reg_0057;
  reg [13:0] reg_0058;
  reg [13:0] reg_0059;
  reg [13:0] reg_0060;
  reg [13:0] reg_0061;
  reg [13:0] reg_0062;
  reg [13:0] reg_0063;
  reg [13:0] reg_0064;
  reg [13:0] reg_0065;
  reg [13:0] reg_0066;
  reg [13:0] reg_0067;
  reg [13:0] reg_0068;
  reg [13:0] reg_0069;
  reg [13:0] reg_0070;
  reg [13:0] reg_0071;
  reg [13:0] reg_0072;
  reg [13:0] reg_0073;
  reg [13:0] reg_0074;
  reg [13:0] reg_0075;
  reg [13:0] reg_0076;
  reg [13:0] reg_0077;
  reg [13:0] reg_0078;
  reg [13:0] reg_0079;
  reg [13:0] reg_0080;
  reg [13:0] reg_0081;
  reg [13:0] reg_0082;
  reg [13:0] reg_0083;
  reg [13:0] reg_0084;
  reg [13:0] reg_0085;
  reg [13:0] reg_0086;
  reg [13:0] reg_0087;
  reg [13:0] reg_0088;
  reg [13:0] reg_0089;
  reg [13:0] reg_0090;
  reg [13:0] reg_0091;
  reg [13:0] reg_0092;
  reg [13:0] reg_0093;
  reg [13:0] reg_0094;
  reg [13:0] reg_0095;
  reg [13:0] reg_0096;
  reg [13:0] reg_0097;
  reg [13:0] reg_0098;
  reg [13:0] reg_0099;
  reg [13:0] reg_0100;
  reg [13:0] reg_0101;
  reg [13:0] reg_0102;
  reg [13:0] reg_0103;
  reg [13:0] reg_0104;
  reg [13:0] reg_0105;
  reg [13:0] reg_0106;
  reg [13:0] reg_0107;
  reg [13:0] reg_0108;
  reg [13:0] reg_0109;

  // 制御マシンの状態
  reg [5:0] state;
  reg _busy;
  assign busy = _busy;
  // 制御マシンの動作
  always @ ( posedge clock or negedge reset ) begin
    if ( !reset ) begin
      _busy <= 0;
      state <= 0;
    end
    else if ( _busy ) begin
      if ( state < 37 ) begin
        state <= state + 1;
      end
      else begin
        _busy <= 0;
        state <= 0;
      end
    end
    else if ( start ) begin
      _busy <= 1;
    end
  end

  // 0番目の入力用メモリブロックの制御
  reg [5:0] _imem00_bank;
  always @ ( * ) begin
    case ( state )
    27: _imem00_bank = 0;
    26: _imem00_bank = 1;
    25: _imem00_bank = 5;
    24: _imem00_bank = 6;
    23: _imem00_bank = 10;
    22: _imem00_bank = 14;
    21: _imem00_bank = 16;
    20: _imem00_bank = 18;
    19: _imem00_bank = 19;
    18: _imem00_bank = 21;
    17: _imem00_bank = 22;
    16: _imem00_bank = 26;
    15: _imem00_bank = 27;
    14: _imem00_bank = 29;
    13: _imem00_bank = 30;
    12: _imem00_bank = 33;
    11: _imem00_bank = 35;
    10: _imem00_bank = 36;
    9: _imem00_bank = 37;
    8: _imem00_bank = 38;
    7: _imem00_bank = 39;
    6: _imem00_bank = 41;
    5: _imem00_bank = 46;
    4: _imem00_bank = 50;
    3: _imem00_bank = 52;
    2: _imem00_bank = 55;
    1: _imem00_bank = 56;
    0: _imem00_bank = 57;
    default: _imem00_bank = 0;
    endcase
  end // always @ ( * )
  assign imem00_bank = _imem00_bank;
  reg _imem00_rd;
  always @ ( * ) begin
    case ( state )
    27: _imem00_rd = 1;
    26: _imem00_rd = 1;
    25: _imem00_rd = 1;
    24: _imem00_rd = 1;
    23: _imem00_rd = 1;
    22: _imem00_rd = 1;
    21: _imem00_rd = 1;
    20: _imem00_rd = 1;
    19: _imem00_rd = 1;
    18: _imem00_rd = 1;
    17: _imem00_rd = 1;
    16: _imem00_rd = 1;
    15: _imem00_rd = 1;
    14: _imem00_rd = 1;
    13: _imem00_rd = 1;
    12: _imem00_rd = 1;
    11: _imem00_rd = 1;
    10: _imem00_rd = 1;
    9: _imem00_rd = 1;
    8: _imem00_rd = 1;
    7: _imem00_rd = 1;
    6: _imem00_rd = 1;
    5: _imem00_rd = 1;
    4: _imem00_rd = 1;
    3: _imem00_rd = 1;
    2: _imem00_rd = 1;
    1: _imem00_rd = 1;
    0: _imem00_rd = 1;
    default: _imem00_rd = 0;
    endcase
  end // always @ ( * )
  assign imem00_rd = _imem00_rd;

  // 1番目の入力用メモリブロックの制御
  reg [5:0] _imem01_bank;
  always @ ( * ) begin
    case ( state )
    27: _imem01_bank = 0;
    26: _imem01_bank = 1;
    25: _imem01_bank = 2;
    24: _imem01_bank = 3;
    23: _imem01_bank = 7;
    22: _imem01_bank = 8;
    21: _imem01_bank = 10;
    20: _imem01_bank = 13;
    19: _imem01_bank = 14;
    18: _imem01_bank = 15;
    17: _imem01_bank = 18;
    16: _imem01_bank = 19;
    15: _imem01_bank = 21;
    14: _imem01_bank = 26;
    13: _imem01_bank = 27;
    12: _imem01_bank = 28;
    11: _imem01_bank = 30;
    10: _imem01_bank = 33;
    9: _imem01_bank = 35;
    8: _imem01_bank = 37;
    7: _imem01_bank = 39;
    6: _imem01_bank = 40;
    5: _imem01_bank = 41;
    4: _imem01_bank = 42;
    3: _imem01_bank = 43;
    2: _imem01_bank = 44;
    1: _imem01_bank = 45;
    0: _imem01_bank = 49;
    33: _imem01_bank = 52;
    32: _imem01_bank = 54;
    31: _imem01_bank = 55;
    30: _imem01_bank = 57;
    29: _imem01_bank = 58;
    28: _imem01_bank = 59;
    default: _imem01_bank = 0;
    endcase
  end // always @ ( * )
  assign imem01_bank = _imem01_bank;
  reg _imem01_rd;
  always @ ( * ) begin
    case ( state )
    27: _imem01_rd = 1;
    26: _imem01_rd = 1;
    25: _imem01_rd = 1;
    24: _imem01_rd = 1;
    23: _imem01_rd = 1;
    22: _imem01_rd = 1;
    21: _imem01_rd = 1;
    20: _imem01_rd = 1;
    19: _imem01_rd = 1;
    18: _imem01_rd = 1;
    17: _imem01_rd = 1;
    16: _imem01_rd = 1;
    15: _imem01_rd = 1;
    14: _imem01_rd = 1;
    13: _imem01_rd = 1;
    12: _imem01_rd = 1;
    11: _imem01_rd = 1;
    10: _imem01_rd = 1;
    9: _imem01_rd = 1;
    8: _imem01_rd = 1;
    7: _imem01_rd = 1;
    6: _imem01_rd = 1;
    5: _imem01_rd = 1;
    4: _imem01_rd = 1;
    3: _imem01_rd = 1;
    2: _imem01_rd = 1;
    1: _imem01_rd = 1;
    0: _imem01_rd = 1;
    33: _imem01_rd = 1;
    32: _imem01_rd = 1;
    31: _imem01_rd = 1;
    30: _imem01_rd = 1;
    29: _imem01_rd = 1;
    28: _imem01_rd = 1;
    default: _imem01_rd = 0;
    endcase
  end // always @ ( * )
  assign imem01_rd = _imem01_rd;

  // 2番目の入力用メモリブロックの制御
  reg [5:0] _imem02_bank;
  always @ ( * ) begin
    case ( state )
    33: _imem02_bank = 4;
    32: _imem02_bank = 6;
    31: _imem02_bank = 7;
    30: _imem02_bank = 11;
    29: _imem02_bank = 14;
    28: _imem02_bank = 16;
    27: _imem02_bank = 17;
    26: _imem02_bank = 18;
    25: _imem02_bank = 20;
    24: _imem02_bank = 21;
    23: _imem02_bank = 22;
    22: _imem02_bank = 23;
    21: _imem02_bank = 24;
    20: _imem02_bank = 26;
    19: _imem02_bank = 27;
    18: _imem02_bank = 29;
    17: _imem02_bank = 30;
    16: _imem02_bank = 31;
    15: _imem02_bank = 32;
    14: _imem02_bank = 33;
    13: _imem02_bank = 35;
    12: _imem02_bank = 36;
    11: _imem02_bank = 39;
    10: _imem02_bank = 42;
    9: _imem02_bank = 43;
    8: _imem02_bank = 47;
    7: _imem02_bank = 50;
    6: _imem02_bank = 51;
    5: _imem02_bank = 55;
    4: _imem02_bank = 56;
    3: _imem02_bank = 57;
    2: _imem02_bank = 59;
    default: _imem02_bank = 0;
    endcase
  end // always @ ( * )
  assign imem02_bank = _imem02_bank;
  reg _imem02_rd;
  always @ ( * ) begin
    case ( state )
    33: _imem02_rd = 1;
    32: _imem02_rd = 1;
    31: _imem02_rd = 1;
    30: _imem02_rd = 1;
    29: _imem02_rd = 1;
    28: _imem02_rd = 1;
    27: _imem02_rd = 1;
    26: _imem02_rd = 1;
    25: _imem02_rd = 1;
    24: _imem02_rd = 1;
    23: _imem02_rd = 1;
    22: _imem02_rd = 1;
    21: _imem02_rd = 1;
    20: _imem02_rd = 1;
    19: _imem02_rd = 1;
    18: _imem02_rd = 1;
    17: _imem02_rd = 1;
    16: _imem02_rd = 1;
    15: _imem02_rd = 1;
    14: _imem02_rd = 1;
    13: _imem02_rd = 1;
    12: _imem02_rd = 1;
    11: _imem02_rd = 1;
    10: _imem02_rd = 1;
    9: _imem02_rd = 1;
    8: _imem02_rd = 1;
    7: _imem02_rd = 1;
    6: _imem02_rd = 1;
    5: _imem02_rd = 1;
    4: _imem02_rd = 1;
    3: _imem02_rd = 1;
    2: _imem02_rd = 1;
    default: _imem02_rd = 0;
    endcase
  end // always @ ( * )
  assign imem02_rd = _imem02_rd;

  // 3番目の入力用メモリブロックの制御
  reg [5:0] _imem03_bank;
  always @ ( * ) begin
    case ( state )
    17: _imem03_bank = 0;
    16: _imem03_bank = 1;
    15: _imem03_bank = 2;
    14: _imem03_bank = 6;
    13: _imem03_bank = 7;
    12: _imem03_bank = 9;
    11: _imem03_bank = 10;
    10: _imem03_bank = 11;
    9: _imem03_bank = 12;
    8: _imem03_bank = 13;
    7: _imem03_bank = 15;
    6: _imem03_bank = 16;
    5: _imem03_bank = 17;
    4: _imem03_bank = 19;
    3: _imem03_bank = 20;
    2: _imem03_bank = 23;
    1: _imem03_bank = 28;
    0: _imem03_bank = 30;
    32: _imem03_bank = 31;
    31: _imem03_bank = 39;
    30: _imem03_bank = 40;
    29: _imem03_bank = 41;
    28: _imem03_bank = 44;
    27: _imem03_bank = 45;
    26: _imem03_bank = 46;
    25: _imem03_bank = 48;
    24: _imem03_bank = 50;
    23: _imem03_bank = 51;
    22: _imem03_bank = 55;
    21: _imem03_bank = 56;
    20: _imem03_bank = 57;
    19: _imem03_bank = 58;
    18: _imem03_bank = 59;
    default: _imem03_bank = 0;
    endcase
  end // always @ ( * )
  assign imem03_bank = _imem03_bank;
  reg _imem03_rd;
  always @ ( * ) begin
    case ( state )
    17: _imem03_rd = 1;
    16: _imem03_rd = 1;
    15: _imem03_rd = 1;
    14: _imem03_rd = 1;
    13: _imem03_rd = 1;
    12: _imem03_rd = 1;
    11: _imem03_rd = 1;
    10: _imem03_rd = 1;
    9: _imem03_rd = 1;
    8: _imem03_rd = 1;
    7: _imem03_rd = 1;
    6: _imem03_rd = 1;
    5: _imem03_rd = 1;
    4: _imem03_rd = 1;
    3: _imem03_rd = 1;
    2: _imem03_rd = 1;
    1: _imem03_rd = 1;
    0: _imem03_rd = 1;
    32: _imem03_rd = 1;
    31: _imem03_rd = 1;
    30: _imem03_rd = 1;
    29: _imem03_rd = 1;
    28: _imem03_rd = 1;
    27: _imem03_rd = 1;
    26: _imem03_rd = 1;
    25: _imem03_rd = 1;
    24: _imem03_rd = 1;
    23: _imem03_rd = 1;
    22: _imem03_rd = 1;
    21: _imem03_rd = 1;
    20: _imem03_rd = 1;
    19: _imem03_rd = 1;
    18: _imem03_rd = 1;
    default: _imem03_rd = 0;
    endcase
  end // always @ ( * )
  assign imem03_rd = _imem03_rd;

  // 4番目の入力用メモリブロックの制御
  reg [5:0] _imem04_bank;
  always @ ( * ) begin
    case ( state )
    32: _imem04_bank = 1;
    31: _imem04_bank = 2;
    30: _imem04_bank = 4;
    29: _imem04_bank = 5;
    28: _imem04_bank = 7;
    27: _imem04_bank = 8;
    26: _imem04_bank = 9;
    25: _imem04_bank = 11;
    24: _imem04_bank = 14;
    23: _imem04_bank = 16;
    22: _imem04_bank = 17;
    21: _imem04_bank = 19;
    20: _imem04_bank = 21;
    34: _imem04_bank = 22;
    33: _imem04_bank = 25;
    19: _imem04_bank = 26;
    18: _imem04_bank = 28;
    17: _imem04_bank = 30;
    16: _imem04_bank = 31;
    15: _imem04_bank = 33;
    14: _imem04_bank = 34;
    13: _imem04_bank = 35;
    12: _imem04_bank = 36;
    11: _imem04_bank = 38;
    10: _imem04_bank = 39;
    9: _imem04_bank = 40;
    8: _imem04_bank = 41;
    7: _imem04_bank = 43;
    6: _imem04_bank = 45;
    5: _imem04_bank = 48;
    4: _imem04_bank = 50;
    3: _imem04_bank = 52;
    2: _imem04_bank = 53;
    1: _imem04_bank = 56;
    0: _imem04_bank = 57;
    default: _imem04_bank = 0;
    endcase
  end // always @ ( * )
  assign imem04_bank = _imem04_bank;
  reg _imem04_rd;
  always @ ( * ) begin
    case ( state )
    32: _imem04_rd = 1;
    31: _imem04_rd = 1;
    30: _imem04_rd = 1;
    29: _imem04_rd = 1;
    28: _imem04_rd = 1;
    27: _imem04_rd = 1;
    26: _imem04_rd = 1;
    25: _imem04_rd = 1;
    24: _imem04_rd = 1;
    23: _imem04_rd = 1;
    22: _imem04_rd = 1;
    21: _imem04_rd = 1;
    20: _imem04_rd = 1;
    34: _imem04_rd = 1;
    33: _imem04_rd = 1;
    19: _imem04_rd = 1;
    18: _imem04_rd = 1;
    17: _imem04_rd = 1;
    16: _imem04_rd = 1;
    15: _imem04_rd = 1;
    14: _imem04_rd = 1;
    13: _imem04_rd = 1;
    12: _imem04_rd = 1;
    11: _imem04_rd = 1;
    10: _imem04_rd = 1;
    9: _imem04_rd = 1;
    8: _imem04_rd = 1;
    7: _imem04_rd = 1;
    6: _imem04_rd = 1;
    5: _imem04_rd = 1;
    4: _imem04_rd = 1;
    3: _imem04_rd = 1;
    2: _imem04_rd = 1;
    1: _imem04_rd = 1;
    0: _imem04_rd = 1;
    default: _imem04_rd = 0;
    endcase
  end // always @ ( * )
  assign imem04_rd = _imem04_rd;

  // 0番目の出力用メモリブロックの制御
  reg [-1:0] _omem00_bank;
  always @ ( * ) begin
    case ( state )
    37: _omem00_bank = 0;
    default: _omem00_bank = 0;
    endcase
  end // always @ ( * )
  assign omem00_bank = _omem00_bank;
  reg _omem00_wr;
  always @ ( * ) begin
    case ( state )
    37: _omem00_wr = 1;
    default: _omem00_wr = 0;
    endcase
  end // always @ ( * )
  assign omem00_wr = _omem00_wr;
  reg [13:0] _omem00_out;
  always @ ( * ) begin
    case ( state )
    37: _omem00_out = reg_0000;
    default: _omem00_out = 0;
    endcase
  end // always @ ( * )
  assign omem00_out = _omem00_out[14:0];

  // OP1#0の0番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in00 = imem00_in[8:0];
    34: op1_00_in00 = imem01_in[8:0];
    18: op1_00_in00 = reg_0048;
    33: op1_00_in00 = imem03_in[8:0];
    35: op1_00_in00 = imem04_in[8:0];
    default: op1_00_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv00 = 1;
    34: op1_00_inv00 = 1;
    default: op1_00_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の1番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in01 = reg_0105;
    34: op1_00_in01 = reg_0021;
    18: op1_00_in01 = reg_0043;
    33: op1_00_in01 = reg_0073;
    35: op1_00_in01 = reg_0001;
    default: op1_00_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv01 = 1;
    33: op1_00_inv01 = 1;
    35: op1_00_inv01 = 1;
    default: op1_00_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の2番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in02 = reg_0102;
    34: op1_00_in02 = reg_0016;
    18: op1_00_in02 = reg_0038;
    33: op1_00_in02 = reg_0068;
    35: op1_00_in02 = reg_0078;
    default: op1_00_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv02 = 1;
    35: op1_00_inv02 = 1;
    default: op1_00_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の3番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in03 = reg_0099;
    34: op1_00_in03 = reg_0011;
    18: op1_00_in03 = reg_0033;
    33: op1_00_in03 = reg_0053;
    35: op1_00_in03 = reg_0058;
    default: op1_00_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv03 = 1;
    34: op1_00_inv03 = 1;
    18: op1_00_inv03 = 1;
    default: op1_00_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の4番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in04 = reg_0096;
    34: op1_00_in04 = reg_0006;
    18: op1_00_in04 = reg_0028;
    33: op1_00_in04 = reg_0049;
    35: op1_00_in04 = reg_0086;
    default: op1_00_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    33: op1_00_inv04 = 1;
    default: op1_00_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の5番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in05 = reg_0093;
    34: op1_00_in05 = reg_0002;
    18: op1_00_in05 = reg_0023;
    33: op1_00_in05 = reg_0044;
    35: op1_00_in05 = reg_0082;
    default: op1_00_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    18: op1_00_inv05 = 1;
    33: op1_00_inv05 = 1;
    default: op1_00_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の6番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in06 = reg_0090;
    34: op1_00_in06 = imem02_in[8:0];
    18: op1_00_in06 = reg_0018;
    33: op1_00_in06 = reg_0039;
    35: op1_00_in06 = reg_0077;
    default: op1_00_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv06 = 1;
    default: op1_00_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の7番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in07 = reg_0087;
    34: op1_00_in07 = reg_0036;
    18: op1_00_in07 = reg_0013;
    33: op1_00_in07 = reg_0034;
    35: op1_00_in07 = reg_0072;
    default: op1_00_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv07 = 1;
    default: op1_00_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の8番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in08 = reg_0068;
    34: op1_00_in08 = reg_0035;
    18: op1_00_in08 = reg_0008;
    33: op1_00_in08 = reg_0029;
    35: op1_00_in08 = reg_0067;
    default: op1_00_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv08 = 1;
    18: op1_00_inv08 = 1;
    33: op1_00_inv08 = 1;
    default: op1_00_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の9番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in09 = reg_0049;
    34: op1_00_in09 = reg_0030;
    18: op1_00_in09 = imem03_in[8:0];
    33: op1_00_in09 = reg_0024;
    35: op1_00_in09 = reg_0062;
    default: op1_00_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv09 = 1;
    34: op1_00_inv09 = 1;
    18: op1_00_inv09 = 1;
    33: op1_00_inv09 = 1;
    default: op1_00_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の10番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in10 = reg_0083;
    34: op1_00_in10 = reg_0025;
    18: op1_00_in10 = reg_0078;
    33: op1_00_in10 = reg_0019;
    35: op1_00_in10 = reg_0057;
    default: op1_00_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv10 = 1;
    33: op1_00_inv10 = 1;
    default: op1_00_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の11番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in11 = reg_0079;
    34: op1_00_in11 = reg_0005;
    18: op1_00_in11 = reg_0073;
    33: op1_00_in11 = reg_0014;
    35: op1_00_in11 = reg_0052;
    default: op1_00_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    33: op1_00_inv11 = 1;
    35: op1_00_inv11 = 1;
    default: op1_00_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の12番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in12 = reg_0074;
    34: op1_00_in12 = reg_0109;
    18: op1_00_in12 = reg_0068;
    33: op1_00_in12 = reg_0009;
    35: op1_00_in12 = reg_0047;
    default: op1_00_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv12 = 1;
    35: op1_00_inv12 = 1;
    default: op1_00_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の13番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in13 = reg_0069;
    34: op1_00_in13 = reg_0048;
    18: op1_00_in13 = reg_0063;
    33: op1_00_in13 = reg_0004;
    35: op1_00_in13 = reg_0042;
    default: op1_00_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv13 = 1;
    33: op1_00_inv13 = 1;
    35: op1_00_inv13 = 1;
    default: op1_00_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の14番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in14 = reg_0064;
    34: op1_00_in14 = reg_0043;
    18: op1_00_in14 = reg_0058;
    33: op1_00_in14 = reg_0000;
    35: op1_00_in14 = reg_0037;
    default: op1_00_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv14 = 1;
    34: op1_00_inv14 = 1;
    33: op1_00_inv14 = 1;
    default: op1_00_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の15番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in15 = reg_0059;
    34: op1_00_in15 = reg_0038;
    18: op1_00_in15 = reg_0053;
    33: op1_00_in15 = imem04_in[8:0];
    35: op1_00_in15 = reg_0032;
    default: op1_00_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv15 = 1;
    18: op1_00_inv15 = 1;
    35: op1_00_inv15 = 1;
    default: op1_00_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の16番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in16 = reg_0054;
    34: op1_00_in16 = reg_0033;
    18: op1_00_in16 = reg_0049;
    33: op1_00_in16 = reg_0031;
    35: op1_00_in16 = reg_0027;
    default: op1_00_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv16 = 1;
    18: op1_00_inv16 = 1;
    default: op1_00_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の17番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in17 = reg_0050;
    34: op1_00_in17 = reg_0028;
    18: op1_00_in17 = reg_0044;
    33: op1_00_in17 = reg_0026;
    35: op1_00_in17 = reg_0022;
    default: op1_00_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv17 = 1;
    34: op1_00_inv17 = 1;
    35: op1_00_inv17 = 1;
    default: op1_00_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の18番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in18 = reg_0045;
    34: op1_00_in18 = reg_0023;
    18: op1_00_in18 = reg_0039;
    33: op1_00_in18 = reg_0020;
    35: op1_00_in18 = reg_0017;
    default: op1_00_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv18 = 1;
    33: op1_00_inv18 = 1;
    35: op1_00_inv18 = 1;
    default: op1_00_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の19番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in19 = reg_0040;
    34: op1_00_in19 = reg_0018;
    18: op1_00_in19 = reg_0034;
    33: op1_00_in19 = reg_0001;
    35: op1_00_in19 = reg_0012;
    default: op1_00_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv19 = 1;
    18: op1_00_inv19 = 1;
    default: op1_00_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の20番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in20 = reg_0035;
    34: op1_00_in20 = reg_0013;
    18: op1_00_in20 = reg_0029;
    33: op1_00_in20 = reg_0108;
    35: op1_00_in20 = reg_0007;
    default: op1_00_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv20 = 1;
    18: op1_00_inv20 = 1;
    33: op1_00_inv20 = 1;
    35: op1_00_inv20 = 1;
    default: op1_00_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の21番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in21 = reg_0030;
    34: op1_00_in21 = reg_0008;
    18: op1_00_in21 = reg_0024;
    33: op1_00_in21 = reg_0107;
    35: op1_00_in21 = reg_0003;
    default: op1_00_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv21 = 1;
    34: op1_00_inv21 = 1;
    18: op1_00_inv21 = 1;
    default: op1_00_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の22番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in22 = reg_0025;
    34: op1_00_in22 = reg_0085;
    18: op1_00_in22 = reg_0019;
    33: op1_00_in22 = reg_0104;
    35: op1_00_in22 = imem04_in[8:0];
    default: op1_00_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv22 = 1;
    33: op1_00_inv22 = 1;
    default: op1_00_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の23番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in23 = reg_0020;
    34: op1_00_in23 = reg_0081;
    18: op1_00_in23 = reg_0014;
    33: op1_00_in23 = reg_0101;
    default: op1_00_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv23 = 1;
    default: op1_00_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の24番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in24 = reg_0015;
    34: op1_00_in24 = reg_0076;
    18: op1_00_in24 = reg_0009;
    33: op1_00_in24 = reg_0098;
    default: op1_00_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv24 = 1;
    33: op1_00_inv24 = 1;
    default: op1_00_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の25番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in25 = reg_0010;
    34: op1_00_in25 = reg_0071;
    18: op1_00_in25 = reg_0004;
    33: op1_00_in25 = reg_0095;
    default: op1_00_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    18: op1_00_inv25 = 1;
    default: op1_00_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の26番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in26 = reg_0005;
    34: op1_00_in26 = reg_0066;
    18: op1_00_in26 = reg_0000;
    33: op1_00_in26 = reg_0092;
    default: op1_00_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv26 = 1;
    34: op1_00_inv26 = 1;
    33: op1_00_inv26 = 1;
    default: op1_00_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の27番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in27 = reg_0001;
    34: op1_00_in27 = reg_0061;
    18: op1_00_in27 = reg_0033;
    33: op1_00_in27 = reg_0089;
    default: op1_00_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv27 = 1;
    18: op1_00_inv27 = 1;
    33: op1_00_inv27 = 1;
    default: op1_00_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の28番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in28 = reg_0093;
    34: op1_00_in28 = reg_0056;
    18: op1_00_in28 = reg_0028;
    33: op1_00_in28 = reg_0049;
    default: op1_00_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    34: op1_00_inv28 = 1;
    33: op1_00_inv28 = 1;
    default: op1_00_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の29番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in29 = reg_0064;
    34: op1_00_in29 = reg_0002;
    18: op1_00_in29 = reg_0004;
    33: op1_00_in29 = reg_0004;
    default: op1_00_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv29 = 1;
    18: op1_00_inv29 = 1;
    33: op1_00_inv29 = 1;
    default: op1_00_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の30番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_00_in30 = reg_0030;
    34: op1_00_in30 = reg_0002;
    18: op1_00_in30 = reg_0000;
    default: op1_00_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_00_inv30 = 1;
    default: op1_00_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#0の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_00_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_00_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の0番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in00 = imem01_in[8:0];
    default: op1_01_in00 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv00 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の1番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in01 = reg_0106;
    default: op1_01_in01 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv01 = 1;
    default: op1_01_inv01 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の2番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in02 = reg_0103;
    default: op1_01_in02 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv02 = 1;
    default: op1_01_inv02 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の3番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in03 = reg_0100;
    default: op1_01_in03 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv03 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の4番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in04 = reg_0097;
    default: op1_01_in04 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv04 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の5番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in05 = reg_0094;
    default: op1_01_in05 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv05 = 1;
    default: op1_01_inv05 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の6番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in06 = reg_0091;
    default: op1_01_in06 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv06 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の7番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in07 = reg_0088;
    default: op1_01_in07 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv07 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の8番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in08 = reg_0073;
    default: op1_01_in08 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv08 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の9番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in09 = reg_0053;
    default: op1_01_in09 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv09 = 1;
    default: op1_01_inv09 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の10番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in10 = reg_0084;
    default: op1_01_in10 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv10 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の11番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in11 = reg_0080;
    default: op1_01_in11 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv11 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の12番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in12 = reg_0075;
    default: op1_01_in12 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv12 = 1;
    default: op1_01_inv12 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の13番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in13 = reg_0070;
    default: op1_01_in13 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv13 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の14番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in14 = reg_0065;
    default: op1_01_in14 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv14 = 1;
    default: op1_01_inv14 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の15番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in15 = reg_0060;
    default: op1_01_in15 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv15 = 1;
    default: op1_01_inv15 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の16番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in16 = reg_0055;
    default: op1_01_in16 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv16 = 1;
    default: op1_01_inv16 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の17番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in17 = reg_0051;
    default: op1_01_in17 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv17 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の18番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in18 = reg_0046;
    default: op1_01_in18 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv18 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の19番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in19 = reg_0041;
    default: op1_01_in19 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv19 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の20番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in20 = reg_0036;
    default: op1_01_in20 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv20 = 1;
    default: op1_01_inv20 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の21番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in21 = reg_0031;
    default: op1_01_in21 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv21 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の22番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in22 = reg_0026;
    default: op1_01_in22 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv22 = 1;
    default: op1_01_inv22 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の23番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in23 = reg_0021;
    default: op1_01_in23 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv23 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の24番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in24 = reg_0016;
    default: op1_01_in24 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv24 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の25番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in25 = reg_0011;
    default: op1_01_in25 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv25 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の26番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in26 = reg_0006;
    default: op1_01_in26 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv26 = 1;
    default: op1_01_inv26 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の27番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in27 = reg_0002;
    default: op1_01_in27 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv27 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の28番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in28 = reg_0094;
    default: op1_01_in28 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    28: op1_01_inv28 = 1;
    default: op1_01_inv28 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の29番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in29 = reg_0073;
    default: op1_01_in29 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv29 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の30番目の入力
  always @ ( * ) begin
    case ( state )
    28: op1_01_in30 = reg_0002;
    default: op1_01_in30 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv30 = 0;
    endcase
  end // always @ ( * )

  // OP1#1の31番目の入力
  always @ ( * ) begin
    case ( state )
    default: op1_01_in31 = 0;
    endcase
  end // always @ ( * )

  // OP1#{}の{}番目の入力反転
  always @ ( * ) begin
    case ( state )
    default: op1_01_inv31 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の0番目の入力
  always @ ( * ) begin
    case ( state )
    36: op2_00_in00 = reg_0010;
    default: op2_00_in00 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の1番目の入力
  always @ ( * ) begin
    case ( state )
    36: op2_00_in01 = reg_0015;
    default: op2_00_in01 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の2番目の入力
  always @ ( * ) begin
    case ( state )
    36: op2_00_in02 = reg_0002;
    default: op2_00_in02 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の3番目の入力
  always @ ( * ) begin
    case ( state )
    36: op2_00_in03 = reg_0063;
    default: op2_00_in03 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の4番目の入力
  always @ ( * ) begin
    case ( state )
    36: op2_00_in04 = reg_0000;
    default: op2_00_in04 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の5番目の入力
  always @ ( * ) begin
    case ( state )
    36: op2_00_in05 = reg_0001;
    default: op2_00_in05 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の6番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in06 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の7番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in07 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の8番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in08 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の9番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in09 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の10番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in10 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の11番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in11 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の12番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in12 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の13番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in13 = 0;
    endcase
  end // always @ ( * )

  // OP2#0の14番目の入力
  always @ ( * ) begin
    case ( state )
    default: op2_00_in14 = 0;
    endcase
  end // always @ ( * )

  // OP2#0のバイアス入力
  always @ ( * ) begin
    case ( state )
    36: op2_00_bias = 84;
    default: op2_00_bias = 0;
    endcase
  end // always @ ( * )

  // REG#0の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0000 <= imem03_in[8:0];
    19: reg_0000 <= imem03_in[8:0];
    33: reg_0000 <= op1_00_out;
    36: reg_0000 <= op2_00_out;
    endcase
  end

  // REG#1の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0001 <= imem00_in[8:0];
    29: reg_0001 <= imem04_in[8:0];
    34: reg_0001 <= imem04_in[8:0];
    35: reg_0001 <= op1_00_out;
    endcase
  end

  // REG#2の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0002 <= imem01_in[8:0];
    29: reg_0002 <= imem01_in[8:0];
    34: reg_0002 <= op1_00_out;
    endcase
  end

  // REG#3の入力
  always @ ( posedge clock ) begin
    case ( state )
    1: reg_0003 <= imem04_in[8:0];
    endcase
  end

  // REG#4の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0004 <= imem03_in[8:0];
    20: reg_0004 <= imem03_in[8:0];
    endcase
  end

  // REG#5の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0005 <= imem00_in[8:0];
    29: reg_0005 <= imem02_in[8:0];
    endcase
  end

  // REG#6の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0006 <= imem01_in[8:0];
    30: reg_0006 <= imem01_in[8:0];
    endcase
  end

  // REG#7の入力
  always @ ( posedge clock ) begin
    case ( state )
    2: reg_0007 <= imem04_in[8:0];
    endcase
  end

  // REG#8の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0008 <= imem02_in[8:0];
    19: reg_0008 <= imem02_in[8:0];
    endcase
  end

  // REG#9の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0009 <= imem03_in[8:0];
    21: reg_0009 <= imem03_in[8:0];
    endcase
  end

  // REG#10の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0010 <= imem00_in[8:0];
    28: reg_0010 <= op1_00_out;
    endcase
  end

  // REG#11の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0011 <= imem01_in[8:0];
    31: reg_0011 <= imem01_in[8:0];
    endcase
  end

  // REG#12の入力
  always @ ( posedge clock ) begin
    case ( state )
    3: reg_0012 <= imem04_in[8:0];
    endcase
  end

  // REG#13の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0013 <= imem02_in[8:0];
    20: reg_0013 <= imem02_in[8:0];
    endcase
  end

  // REG#14の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0014 <= imem03_in[8:0];
    22: reg_0014 <= imem03_in[8:0];
    endcase
  end

  // REG#15の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0015 <= imem00_in[8:0];
    28: reg_0015 <= op1_01_out;
    endcase
  end

  // REG#16の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0016 <= imem01_in[8:0];
    32: reg_0016 <= imem01_in[8:0];
    endcase
  end

  // REG#17の入力
  always @ ( posedge clock ) begin
    case ( state )
    4: reg_0017 <= imem04_in[8:0];
    endcase
  end

  // REG#18の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0018 <= imem02_in[8:0];
    21: reg_0018 <= imem02_in[8:0];
    endcase
  end

  // REG#19の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0019 <= imem03_in[8:0];
    23: reg_0019 <= imem03_in[8:0];
    endcase
  end

  // REG#20の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0020 <= imem00_in[8:0];
    30: reg_0020 <= imem04_in[8:0];
    endcase
  end

  // REG#21の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0021 <= imem01_in[8:0];
    33: reg_0021 <= imem01_in[8:0];
    endcase
  end

  // REG#22の入力
  always @ ( posedge clock ) begin
    case ( state )
    5: reg_0022 <= imem04_in[8:0];
    endcase
  end

  // REG#23の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0023 <= imem02_in[8:0];
    22: reg_0023 <= imem02_in[8:0];
    endcase
  end

  // REG#24の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0024 <= imem03_in[8:0];
    24: reg_0024 <= imem03_in[8:0];
    endcase
  end

  // REG#25の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0025 <= imem00_in[8:0];
    30: reg_0025 <= imem02_in[8:0];
    endcase
  end

  // REG#26の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0026 <= imem01_in[8:0];
    31: reg_0026 <= imem04_in[8:0];
    endcase
  end

  // REG#27の入力
  always @ ( posedge clock ) begin
    case ( state )
    6: reg_0027 <= imem04_in[8:0];
    endcase
  end

  // REG#28の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0028 <= imem02_in[8:0];
    23: reg_0028 <= imem02_in[8:0];
    endcase
  end

  // REG#29の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0029 <= imem03_in[8:0];
    25: reg_0029 <= imem03_in[8:0];
    endcase
  end

  // REG#30の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0030 <= imem00_in[8:0];
    31: reg_0030 <= imem02_in[8:0];
    endcase
  end

  // REG#31の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0031 <= imem01_in[8:0];
    32: reg_0031 <= imem04_in[8:0];
    endcase
  end

  // REG#32の入力
  always @ ( posedge clock ) begin
    case ( state )
    7: reg_0032 <= imem04_in[8:0];
    endcase
  end

  // REG#33の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0033 <= imem02_in[8:0];
    24: reg_0033 <= imem02_in[8:0];
    endcase
  end

  // REG#34の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0034 <= imem03_in[8:0];
    26: reg_0034 <= imem03_in[8:0];
    endcase
  end

  // REG#35の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0035 <= imem00_in[8:0];
    32: reg_0035 <= imem02_in[8:0];
    endcase
  end

  // REG#36の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0036 <= imem01_in[8:0];
    33: reg_0036 <= imem02_in[8:0];
    endcase
  end

  // REG#37の入力
  always @ ( posedge clock ) begin
    case ( state )
    8: reg_0037 <= imem04_in[8:0];
    endcase
  end

  // REG#38の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0038 <= imem02_in[8:0];
    25: reg_0038 <= imem02_in[8:0];
    endcase
  end

  // REG#39の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0039 <= imem03_in[8:0];
    27: reg_0039 <= imem03_in[8:0];
    endcase
  end

  // REG#40の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0040 <= imem00_in[8:0];
    endcase
  end

  // REG#41の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0041 <= imem01_in[8:0];
    endcase
  end

  // REG#42の入力
  always @ ( posedge clock ) begin
    case ( state )
    9: reg_0042 <= imem04_in[8:0];
    endcase
  end

  // REG#43の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0043 <= imem02_in[8:0];
    26: reg_0043 <= imem02_in[8:0];
    endcase
  end

  // REG#44の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0044 <= imem03_in[8:0];
    28: reg_0044 <= imem03_in[8:0];
    endcase
  end

  // REG#45の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0045 <= imem00_in[8:0];
    endcase
  end

  // REG#46の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0046 <= imem01_in[8:0];
    endcase
  end

  // REG#47の入力
  always @ ( posedge clock ) begin
    case ( state )
    10: reg_0047 <= imem04_in[8:0];
    endcase
  end

  // REG#48の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0048 <= imem02_in[8:0];
    27: reg_0048 <= imem02_in[8:0];
    endcase
  end

  // REG#49の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0049 <= imem03_in[8:0];
    19: reg_0049 <= imem00_in[8:0];
    29: reg_0049 <= imem03_in[8:0];
    endcase
  end

  // REG#50の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0050 <= imem00_in[8:0];
    endcase
  end

  // REG#51の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0051 <= imem01_in[8:0];
    endcase
  end

  // REG#52の入力
  always @ ( posedge clock ) begin
    case ( state )
    11: reg_0052 <= imem04_in[8:0];
    endcase
  end

  // REG#53の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0053 <= imem03_in[8:0];
    19: reg_0053 <= imem01_in[8:0];
    30: reg_0053 <= imem03_in[8:0];
    endcase
  end

  // REG#54の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0054 <= imem00_in[8:0];
    endcase
  end

  // REG#55の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0055 <= imem01_in[8:0];
    endcase
  end

  // REG#56の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0056 <= imem02_in[8:0];
    endcase
  end

  // REG#57の入力
  always @ ( posedge clock ) begin
    case ( state )
    12: reg_0057 <= imem04_in[8:0];
    endcase
  end

  // REG#58の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0058 <= imem03_in[8:0];
    19: reg_0058 <= imem04_in[8:0];
    endcase
  end

  // REG#59の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0059 <= imem00_in[8:0];
    endcase
  end

  // REG#60の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0060 <= imem01_in[8:0];
    endcase
  end

  // REG#61の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0061 <= imem02_in[8:0];
    endcase
  end

  // REG#62の入力
  always @ ( posedge clock ) begin
    case ( state )
    13: reg_0062 <= imem04_in[8:0];
    endcase
  end

  // REG#63の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0063 <= imem03_in[8:0];
    18: reg_0063 <= op1_00_out;
    endcase
  end

  // REG#64の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0064 <= imem00_in[8:0];
    endcase
  end

  // REG#65の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0065 <= imem01_in[8:0];
    endcase
  end

  // REG#66の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0066 <= imem02_in[8:0];
    endcase
  end

  // REG#67の入力
  always @ ( posedge clock ) begin
    case ( state )
    14: reg_0067 <= imem04_in[8:0];
    endcase
  end

  // REG#68の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0068 <= imem03_in[8:0];
    20: reg_0068 <= imem00_in[8:0];
    31: reg_0068 <= imem03_in[8:0];
    endcase
  end

  // REG#69の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0069 <= imem00_in[8:0];
    endcase
  end

  // REG#70の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0070 <= imem01_in[8:0];
    endcase
  end

  // REG#71の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0071 <= imem02_in[8:0];
    endcase
  end

  // REG#72の入力
  always @ ( posedge clock ) begin
    case ( state )
    15: reg_0072 <= imem04_in[8:0];
    endcase
  end

  // REG#73の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0073 <= imem03_in[8:0];
    20: reg_0073 <= imem01_in[8:0];
    32: reg_0073 <= imem03_in[8:0];
    endcase
  end

  // REG#74の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0074 <= imem00_in[8:0];
    endcase
  end

  // REG#75の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0075 <= imem01_in[8:0];
    endcase
  end

  // REG#76の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0076 <= imem02_in[8:0];
    endcase
  end

  // REG#77の入力
  always @ ( posedge clock ) begin
    case ( state )
    16: reg_0077 <= imem04_in[8:0];
    endcase
  end

  // REG#78の入力
  always @ ( posedge clock ) begin
    case ( state )
    17: reg_0078 <= imem03_in[8:0];
    20: reg_0078 <= imem04_in[8:0];
    endcase
  end

  // REG#79の入力
  always @ ( posedge clock ) begin
    case ( state )
    17: reg_0079 <= imem00_in[8:0];
    endcase
  end

  // REG#80の入力
  always @ ( posedge clock ) begin
    case ( state )
    17: reg_0080 <= imem01_in[8:0];
    endcase
  end

  // REG#81の入力
  always @ ( posedge clock ) begin
    case ( state )
    17: reg_0081 <= imem02_in[8:0];
    endcase
  end

  // REG#82の入力
  always @ ( posedge clock ) begin
    case ( state )
    17: reg_0082 <= imem04_in[8:0];
    endcase
  end

  // REG#83の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0083 <= imem00_in[8:0];
    endcase
  end

  // REG#84の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0084 <= imem01_in[8:0];
    endcase
  end

  // REG#85の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0085 <= imem02_in[8:0];
    endcase
  end

  // REG#86の入力
  always @ ( posedge clock ) begin
    case ( state )
    18: reg_0086 <= imem04_in[8:0];
    endcase
  end

  // REG#87の入力
  always @ ( posedge clock ) begin
    case ( state )
    21: reg_0087 <= imem00_in[8:0];
    endcase
  end

  // REG#88の入力
  always @ ( posedge clock ) begin
    case ( state )
    21: reg_0088 <= imem01_in[8:0];
    endcase
  end

  // REG#89の入力
  always @ ( posedge clock ) begin
    case ( state )
    21: reg_0089 <= imem04_in[8:0];
    endcase
  end

  // REG#90の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0090 <= imem00_in[8:0];
    endcase
  end

  // REG#91の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0091 <= imem01_in[8:0];
    endcase
  end

  // REG#92の入力
  always @ ( posedge clock ) begin
    case ( state )
    22: reg_0092 <= imem04_in[8:0];
    endcase
  end

  // REG#93の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0093 <= imem00_in[8:0];
    endcase
  end

  // REG#94の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0094 <= imem01_in[8:0];
    endcase
  end

  // REG#95の入力
  always @ ( posedge clock ) begin
    case ( state )
    23: reg_0095 <= imem04_in[8:0];
    endcase
  end

  // REG#96の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0096 <= imem00_in[8:0];
    endcase
  end

  // REG#97の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0097 <= imem01_in[8:0];
    endcase
  end

  // REG#98の入力
  always @ ( posedge clock ) begin
    case ( state )
    24: reg_0098 <= imem04_in[8:0];
    endcase
  end

  // REG#99の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0099 <= imem00_in[8:0];
    endcase
  end

  // REG#100の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0100 <= imem01_in[8:0];
    endcase
  end

  // REG#101の入力
  always @ ( posedge clock ) begin
    case ( state )
    25: reg_0101 <= imem04_in[8:0];
    endcase
  end

  // REG#102の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0102 <= imem00_in[8:0];
    endcase
  end

  // REG#103の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0103 <= imem01_in[8:0];
    endcase
  end

  // REG#104の入力
  always @ ( posedge clock ) begin
    case ( state )
    26: reg_0104 <= imem04_in[8:0];
    endcase
  end

  // REG#105の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0105 <= imem00_in[8:0];
    endcase
  end

  // REG#106の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0106 <= imem01_in[8:0];
    endcase
  end

  // REG#107の入力
  always @ ( posedge clock ) begin
    case ( state )
    27: reg_0107 <= imem04_in[8:0];
    endcase
  end

  // REG#108の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0108 <= imem04_in[8:0];
    endcase
  end

  // REG#109の入力
  always @ ( posedge clock ) begin
    case ( state )
    28: reg_0109 <= imem02_in[8:0];
    endcase
  end
endmodule
